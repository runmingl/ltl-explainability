module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, jx0_n, jx1_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844f9f;
  wire v870222;
  wire v870225;
  wire v87048e;
  wire v8705c8;
  wire v86608f;
  wire v85a15e;
  wire v8702f6;
  wire v869783;
  wire v8660ef;
  wire v87045b;
  wire v870501;
  wire v84ff79;
  wire v870286;
  wire v870234;
  wire v865660;
  wire v865c3f;
  wire v866122;
  wire v865df6;
  wire v865f18;
  wire v87028c;
  wire v865cf1;
  wire v844fb3;
  wire v87055d;
  wire v865b09;
  wire v865ba1;
  wire v8656f8;
  wire v865faa;
  wire v8702c8;
  wire v8702fd;
  wire v8702bf;
  wire v8702a3;
  wire v844f99;
  wire v859e32;
  wire v865b7c;
  wire v866192;
  wire v8659c0;
  wire v865985;
  wire v86c31f;
  wire v865db0;
  wire v8659de;
  wire v85dbde;
  wire v865fcf;
  wire v8657e8;
  wire v865b52;
  wire v870333;
  wire v844fb5;
  wire v8660f2;
  wire v870235;
  wire v86596b;
  wire v854981;
  wire v8540cb;
  wire v865a3e;
  wire v8701ff;
  wire v865c02;
  wire v87021b;
  wire v865dd5;
  wire v870246;
  wire v870300;
  wire v8702a6;
  wire v870356;
  wire v865981;
  wire v865860;
  wire v865d5a;
  wire v85dc04;
  wire v844fa9;
  wire v844fab;
  wire v865ee5;
  wire v8694e4;
  wire v865f3c;
  wire v859b38;
  wire v865701;
  wire v8657f0;
  wire v8659f1;
  wire v85984b;
  wire v8657ee;
  wire v865857;
  wire v8702ed;
  wire v859822;
  wire v865c6a;
  wire v866044;
  wire v86c34e;
  wire v8658c7;
  wire v865884;
  wire v86b5b5;
  wire v85dbed;
  wire v8703f4;
  wire v865bf0;
  wire v870283;
  wire v87029f;
  wire v870245;
  wire v854cf5;
  wire v8694ff;
  wire v865858;
  wire v865ff1;
  wire v8702ce;
  wire v8702d4;
  wire v869509;
  wire v85dc00;
  wire v870229;
  wire v8587be;
  wire v865aff;
  wire v870277;
  wire v865f98;
  wire v8659dc;
  wire v865be6;
  wire v87023f;
  wire v8656be;
  wire v850277;
  wire v870271;
  wire v858899;
  wire v8661ce;
  wire v8659c8;
  wire v870281;
  wire v870259;
  wire v865992;
  wire v8599b0;
  wire v8704fd;
  wire v8702bc;
  wire v865f25;
  wire v865c64;
  wire v8658dc;
  wire v86c352;
  wire v865d41;
  wire v870297;
  wire v865d52;
  wire v8702f2;
  wire v87034b;
  wire v865c69;
  wire v865698;
  wire v870218;
  wire v865eef;
  wire v850b88;
  wire v865a28;
  wire v865c5b;
  wire v870278;
  wire v865908;
  wire v865ae5;
  wire v8703e0;
  wire v865da4;
  wire v858431;
  wire v865dd3;
  wire v865af5;
  wire v85445c;
  wire v8657b3;
  wire v850ad2;
  wire v86597b;
  wire v8702d1;
  wire v87029a;
  wire v865fa1;
  wire v865cd9;
  wire v865bed;
  wire v850173;
  wire v865eee;
  wire v8702a2;
  wire v865817;
  wire v86c325;
  wire v8702e1;
  wire v8702cb;
  wire v858630;
  wire v86564e;
  wire v8510be;
  wire v86c356;
  wire v865678;
  wire v8659bf;
  wire v865894;
  wire v8656cf;
  wire v865c20;
  wire v844f97;
  wire v865b94;
  wire v865c91;
  wire v87023b;
  wire v8702d9;
  wire v866158;
  wire v865f6f;
  wire v86594c;
  wire v865f3b;
  wire v8705b3;
  wire v8658b3;
  wire v865cb0;
  wire v870295;
  wire v86f0aa;
  wire v84fc72;
  wire v870476;
  wire v865623;
  wire v865f4b;
  wire v865944;
  wire v870491;
  wire v865644;
  wire v865673;
  wire v865b61;
  wire v87054a;
  wire v865c17;
  wire v8660d6;
  wire v87056c;
  wire v85a72b;
  wire v8705c0;
  wire v85a5c4;
  wire v86575b;
  wire v850fb5;
  wire v865fbb;
  wire v865b98;
  wire v86587c;
  wire v865f92;
  wire v865833;
  wire v85dbd8;
  wire v865632;
  wire v865da6;
  wire v86587f;
  wire v865622;
  wire v865a51;
  wire v867fda;
  wire v86571d;
  wire v865d63;
  wire v8659c5;
  wire v8702f8;
  wire v87026a;
  wire v8703a0;
  wire v870214;
  wire v865c46;
  wire v86c319;
  wire v84ffd7;
  wire v865863;
  wire v870381;
  wire v8701fb;
  wire v866139;
  wire v86c316;
  wire v865821;
  wire v86c35a;
  wire v865c92;
  wire v86f080;
  wire v8661c8;
  wire v865c36;
  wire v870321;
  wire v84fc5e;
  wire v870269;
  wire v865633;
  wire v8659d6;
  wire v87031c;
  wire v866204;
  wire v865989;
  wire v87020c;
  wire v859f24;
  wire v865791;
  wire v865972;
  wire v865620;
  wire v86b5d8;
  wire v8702aa;
  wire v865ff5;
  wire v8661da;
  wire v86581a;
  wire v8702d0;
  wire v865d20;
  wire v859aa5;
  wire v866128;
  wire v865c8f;
  wire v865d0e;
  wire v866137;
  wire v870348;
  wire v865d46;
  wire v8660b3;
  wire v87021c;
  wire v85a1b8;
  wire v865849;
  wire v8656a0;
  wire v870531;
  wire v8703e9;
  wire v8658a3;
  wire v865fa0;
  wire v86577a;
  wire v8585dc;
  wire v870200;
  wire v870209;
  wire v86c353;
  wire v850031;
  wire v8656bf;
  wire v87029c;
  wire v85a24a;
  wire v865cc1;
  wire v865f60;
  wire v870341;
  wire v866121;
  wire v86575e;
  wire v850aee;
  wire v866093;
  wire v8657d5;
  wire v86f0bf;
  wire v844f95;
  wire v866364;
  wire v8702a8;
  wire v87026f;
  wire v86573e;
  wire v87031a;
  wire v87024a;
  wire v86586d;
  wire v8661e8;
  wire v8660c2;
  wire v8702dc;
  wire v865ce6;
  wire v865ba9;
  wire v865eff;
  wire v85dbe2;
  wire v8704d4;
  wire v870257;
  wire v865cf3;
  wire v870210;
  wire v86dd82;
  wire v8659c3;
  wire v870292;
  wire v870484;
  wire v85dbe6;
  wire v8702a4;
  wire v865920;
  wire v8703ec;
  wire v8694ed;
  wire v87025e;
  wire v865caa;
  wire v87020f;
  wire v8659bb;
  wire v85a738;
  wire v86596e;
  wire v865beb;
  wire v850b89;
  wire v865cbd;
  wire v870284;
  wire v870467;
  wire v8660d5;
  wire v865efd;
  wire v851192;
  wire v870384;
  wire v87022b;
  wire v86b5d5;
  wire v870299;
  wire v851f5b;
  wire v865730;
  wire v865b07;
  wire v86b5e3;
  wire v866108;
  wire v853599;
  wire v870403;
  wire v8703e2;
  wire v865fd7;
  wire v865f0c;
  wire v85dbf9;
  wire v870207;
  wire v870526;
  wire v8656cd;
  wire v865ccf;
  wire v870290;
  wire v8702ca;
  wire v858042;
  wire v850819;
  wire v865d79;
  wire v87030a;
  wire v85162c;
  wire v865b8c;
  wire v8656ea;
  wire v865f8c;
  wire v86600c;
  wire v8702fe;
  wire v869795;
  wire v8584ca;
  wire v8657b4;
  wire v86584f;
  wire v86f0ad;
  wire v87022d;
  wire v8660c0;
  wire v865896;
  wire v867fdc;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  wire SLC0_n;
  wire ENQ_n;

assign v8702f6 = RtoB_ACK0_p & v870225 | !RtoB_ACK0_p & !v85a15e;
assign v8705c8 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v844f9f;
assign v8657b4 = jx1_p & v8584ca | !jx1_p & v853599;
assign v865d63 = BtoS_ACK1_p & v85a5c4 | !BtoS_ACK1_p & v86571d;
assign v865f18 = RtoB_ACK0_p & v87045b | !RtoB_ACK0_p & v865df6;
assign v865efd = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & v8660d5;
assign v866204 = BtoR_REQ1_p & v844fa9 | !BtoR_REQ1_p & v87031c;
assign v865fcf = BtoS_ACK2_p & v844f99 | !BtoS_ACK2_p & v87028c;
assign DEQ_n = !v869509;
assign v870300 = jx0_p & v870246 | !jx0_p & v8657e8;
assign v865b98 = StoB_REQ2_n & v850fb5 | !StoB_REQ2_n & !v865fbb;
assign v865f4b = jx1_p & v86f0aa | !jx1_p & v865623;
assign v8702a8 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8702f6;
assign v866158 = StoB_REQ2_n & v869783 | !StoB_REQ2_n & !v844f91;
assign v8659c3 = StoB_REQ1_p & v8702f6 | !StoB_REQ1_p & !v844f91;
assign v8660c2 = StoB_REQ2_n & v8702f6 | !StoB_REQ2_n & !v844f91;
assign v87021c = jx1_p & v870348 | !jx1_p & v8660b3;
assign v8702ed = RtoB_ACK1_p & v865857 | !RtoB_ACK1_p & !v844f91;
assign BtoR_REQ1_n = v86f0bf;
assign v87034b = StoB_REQ2_p & v865c64 | !StoB_REQ2_p & v865d41;
assign v8702d4 = StoB_REQ0_p & v8694e4 | !StoB_REQ0_p & v8702ce;
assign v87021b = BtoS_ACK2_p & v844f99 | !BtoS_ACK2_p & v865c02;
assign v8660d5 = StoB_REQ1_p & v870467 | !StoB_REQ1_p & !v844f91;
assign v8660f2 = DEQ_p & v844f91 | !DEQ_p & !v844fb5;
assign v85dbd8 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v865f92;
assign v8656f8 = RtoB_ACK0_p & v870225 | !RtoB_ACK0_p & !v865ba1;
assign v8656be = jx0_p & v8659dc | !jx0_p & v87023f;
assign v870209 = jx0_p & v8703e9 | !jx0_p & !v870200;
assign v865857 = BtoR_REQ1_p & v844fa9 | !BtoR_REQ1_p & v844f91;
assign v8702d0 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v86581a;
assign BtoS_ACK2_n = !v85dc04;
assign v8701fb = BtoS_ACK1_p & v85a5c4 | !BtoS_ACK1_p & v870381;
assign v870235 = BtoR_REQ0_p & v8660f2 | !BtoR_REQ0_p & !v844fb5;
assign v865f0c = BtoR_REQ0_p & v844fb5 | !BtoR_REQ0_p & !v844f91;
assign v870531 = StoB_REQ1_p & v8659d6 | !StoB_REQ1_p & !v8656a0;
assign v85dc04 = BtoS_ACK0_p & v8702a3 | !BtoS_ACK0_p & v865d5a;
assign v870278 = StoB_REQ2_p & v865c5b | !StoB_REQ2_p & v858899;
assign v865860 = jx1_p & v870300 | !jx1_p & v865981;
assign v865833 = BtoR_REQ0_p & v865f92 | !BtoR_REQ0_p & !v86587c;
assign v8694e4 = RtoB_ACK0_p & v844fa9 | !RtoB_ACK0_p & v865ee5;
assign v870269 = jx1_p & v870321 | !jx1_p & v84fc5e;
assign v8659f1 = StoB_REQ1_p & v8694e4 | !StoB_REQ1_p & v8657f0;
assign v86608f = BtoR_REQ1_p & v87048e | !BtoR_REQ1_p & v8705c8;
assign v866044 = StoB_REQ1_p & v8694e4 | !StoB_REQ1_p & v865c6a;
assign v8657d5 = StoB_REQ0_p & v87021c | !StoB_REQ0_p & v866093;
assign v86584f = jx0_p & v844f97 | !jx0_p & v844f91;
assign v865730 = jx1_p & v87022b | !jx1_p & v851f5b;
assign v865caa = StoB_REQ1_p & v865c17 | !StoB_REQ1_p & !v844f91;
assign v8656cd = RtoB_ACK0_p & v844fb5 | !RtoB_ACK0_p & v870526;
assign v8599b0 = StoB_REQ2_p & v858899 | !StoB_REQ2_p & v865992;
assign v86573e = BtoS_ACK1_p & v866364 | !BtoS_ACK1_p & !v87026f;
assign v866139 = jx0_p & v84ffd7 | !jx0_p & v8701fb;
assign v87048e = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v870222;
assign v858899 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v870271;
assign v865b09 = BtoR_REQ1_p & v87055d | !BtoR_REQ1_p & v844f91;
assign v865eef = StoB_REQ0_p & v850277 | !StoB_REQ0_p & v870218;
assign v870234 = BtoR_REQ1_p & v870222 | !BtoR_REQ1_p & v870286;
assign v865633 = RtoB_ACK0_p & v844fa9 | !RtoB_ACK0_p & v865c92;
assign v844fa9 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v844f91;
assign v844fb3 = DEQ_p & v844f91 | !DEQ_p & !v844f91;
assign v86564e = BtoS_ACK1_p & v8702e1 | !BtoS_ACK1_p & v858630;
assign v844f91 = 1;
assign v865be6 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844fa9;
assign v870295 = StoB_REQ1_p & v8658b3 | !StoB_REQ1_p & v865cb0;
assign v85a738 = jx1_p & v87025e | !jx1_p & v8659bb;
assign v8694ff = jx0_p & v865bf0 | !jx0_p & v854cf5;
assign v8702cb = BtoS_ACK2_p & v865be6 | !BtoS_ACK2_p & v870297;
assign v859f24 = stateG7_0_p & v865989 | !stateG7_0_p & v87020c;
assign v870491 = StoB_REQ2_n & v8659de | !StoB_REQ2_n & !v844f91;
assign v869509 = BtoS_ACK0_p & v865884 | !BtoS_ACK0_p & v8702d4;
assign v870341 = BtoS_ACK2_p & v865cc1 | !BtoS_ACK2_p & v865f60;
assign v8705b3 = StoB_REQ2_p & v865f18 | !StoB_REQ2_p & !v865f3b;
assign v85a5c4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v866158;
assign v87055d = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v844fb3;
assign v86c35a = BtoS_ACK0_p & v865944 | !BtoS_ACK0_p & !v865821;
assign v8702fe = StoB_REQ0_p & v8656ea | !StoB_REQ0_p & v86600c;
assign v865ba1 = RtoB_ACK1_p & v865b09 | !RtoB_ACK1_p & v844f91;
assign v87025e = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & !v844f91;
assign v865a51 = BtoS_ACK2_p & v865b98 | !BtoS_ACK2_p & v865622;
assign v87030a = jx0_p & v8702ca | !jx0_p & v865d79;
assign v850aee = jx0_p & v850031 | !jx0_p & v86575e;
assign v865b61 = jx0_p & v844f91 | !jx0_p & v865673;
assign v87024a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v87031a;
assign v870321 = StoB_REQ1_p & v86f080 | !StoB_REQ1_p & v865c36;
assign BtoS_ACK1_n = !v86b5e3;
assign v865fa1 = BtoS_ACK1_p & v86597b | !BtoS_ACK1_p & v87029a;
assign v865faa = StoB_REQ2_p & v8656f8 | !StoB_REQ2_p & !v844f91;
assign v8705c0 = jx1_p & v865b61 | !jx1_p & v85a72b;
assign v865817 = StoB_REQ1_p & v865908 | !StoB_REQ1_p & v8702a2;
assign v8656ea = jx1_p & v87030a | !jx1_p & !v865b8c;
assign v85984b = jx0_p & v8657f0 | !jx0_p & v8659f1;
assign v865f60 = StoB_REQ2_p & v865633 | !StoB_REQ2_p & v85a24a;
assign v85dbe2 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v865f18;
assign v865ba9 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v865ce6;
assign v87029a = BtoS_ACK2_p & v8702d1 | !BtoS_ACK2_p & v87034b;
assign v865f3b = RtoB_ACK0_p & v870225 | !RtoB_ACK0_p & !v86594c;
assign v865bed = jx1_p & v865dd3 | !jx1_p & v865cd9;
assign v866364 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8702f6;
assign v8702aa = stateG7_1_p & v844f91 | !stateG7_1_p & v865857;
assign v85dc00 = stateG7_1_p & v865857 | !stateG7_1_p & v844fa9;
assign v84fc72 = StoB_REQ2_n & v865faa | !StoB_REQ2_n & !v844f91;
assign v8702d1 = StoB_REQ2_p & v8587be | !StoB_REQ2_p & v865d41;
assign v8584ca = jx0_p & v844fb5 | !jx0_p & v844f91;
assign v8702c8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v865faa;
assign v86581a = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8661da;
assign v865c92 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v865f25;
assign v86594c = RtoB_ACK1_p & v87055d | !RtoB_ACK1_p & v844f91;
assign v854981 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v844fb5;
assign v85dbf9 = stateG7_1_p & v865f0c | !stateG7_1_p & v844fb5;
assign v866137 = StoB_REQ1_p & v86f080 | !StoB_REQ1_p & v8659d6;
assign v87023f = StoB_REQ2_p & v8587be | !StoB_REQ2_p & v865be6;
assign v865b07 = StoB_REQ0_p & v85a738 | !StoB_REQ0_p & v865730;
assign v8660d6 = StoB_REQ1_p & v865c17 | !StoB_REQ1_p & v844f91;
assign v859aa5 = StoB_REQ1_p & v8659d6 | !StoB_REQ1_p & !v865d20;
assign v865d5a = StoB_REQ0_p & v870333 | !StoB_REQ0_p & v865860;
assign v84ff79 = BtoR_REQ1_p & v870501 | !BtoR_REQ1_p & v844f91;
assign v865b52 = jx0_p & v865b7c | !jx0_p & v8657e8;
assign v870257 = jx0_p & v865eff | !jx0_p & v8704d4;
assign v865660 = stateG7_1_p & v870286 | !stateG7_1_p & v870234;
assign v865896 = jx1_p & v8660c0 | !jx1_p & v865f8c;
assign jx1_n = v867fdc;
assign v865cb0 = StoB_REQ2_n & v87028c | !StoB_REQ2_n & !v844f91;
assign v865cf1 = jx0_p & v8660ef | !jx0_p & !v87028c;
assign v850173 = StoB_REQ1_p & v865f98 | !StoB_REQ1_p & v8599b0;
assign v870284 = StoB_REQ2_n & v8701ff | !StoB_REQ2_n & !v865cbd;
assign v865af5 = StoB_REQ2_p & v8587be | !StoB_REQ2_p & v865c64;
assign v8694ed = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8703ec;
assign v8661c8 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v865c92;
assign v870384 = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & !v851192;
assign v867fdc = BtoS_ACK0_p & v87022d | !BtoS_ACK0_p & v865896;
assign v86f0ad = jx1_p & v8584ca | !jx1_p & !v86584f;
assign v858042 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v85a1b8 = StoB_REQ1_p & v865c36 | !StoB_REQ1_p & !v865620;
assign v870277 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v865aff;
assign v865c3f = stateG7_1_p & v870222 | !stateG7_1_p & v870234;
assign v870290 = BtoS_ACK2_p & v865ccf | !BtoS_ACK2_p & v844fb5;
assign v870484 = StoB_REQ1_p & v870292 | !StoB_REQ1_p & v844f91;
assign v8661da = stateG7_0_p & v8702aa | !stateG7_0_p & v865ff5;
assign v85445c = BtoS_ACK2_p & v865af5 | !BtoS_ACK2_p & v865c64;
assign v865ee5 = RtoB_ACK1_p & v844fab | !RtoB_ACK1_p & v844f91;
assign v8658b3 = StoB_REQ2_n & v8705b3 | !StoB_REQ2_n & !v865f3b;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v865c46 = jx0_p & v865d63 | !jx0_p & v870214;
assign v85a15e = RtoB_ACK1_p & v86608f | !RtoB_ACK1_p & v844f91;
assign v870476 = StoB_REQ1_p & v865db0 | !StoB_REQ1_p & !v84fc72;
assign v86586d = BtoS_ACK1_p & v87024a | !BtoS_ACK1_p & v8702a8;
assign v87026a = StoB_REQ2_n & v8659c5 | !StoB_REQ2_n & !v8702f8;
assign v870271 = RtoB_ACK1_p & v865857 | !RtoB_ACK1_p & v85dc00;
assign v870229 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v85dc00;
assign v8657b3 = StoB_REQ1_p & v85445c | !StoB_REQ1_p & v865be6;
assign v870283 = StoB_REQ1_p & v865701 | !StoB_REQ1_p & v8657f0;
assign v84ffd7 = BtoS_ACK1_p & v85a5c4 | !BtoS_ACK1_p & v86c319;
assign v8703e2 = jx1_p & v866108 | !jx1_p & v865b94;
assign v865858 = BtoS_ACK1_p & v865c6a | !BtoS_ACK1_p & v8703f4;
assign v865dd5 = StoB_REQ1_p & v859e32 | !StoB_REQ1_p & v87021b;
assign v844fab = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v844f91;
assign v8656bf = stateG7_0_p & v8702aa | !stateG7_0_p & v865857;
assign v8660b3 = jx0_p & v865d46 | !jx0_p & v870348;
assign v8659c5 = StoB_REQ2_p & v865f18 | !StoB_REQ2_p & !v8702d9;
assign v865c20 = BtoS_ACK0_p & v865eef | !BtoS_ACK0_p & v8656cf;
assign v865a28 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v844fa9;
assign v8659de = StoB_REQ2_p & v865db0 | !StoB_REQ2_p & !v844f91;
assign v865aff = RtoB_ACK1_p & v844fa9 | !RtoB_ACK1_p & v85dc00;
assign v865bf0 = BtoS_ACK1_p & v86b5b5 | !BtoS_ACK1_p & v8703f4;
assign v87031c = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8660f2;
assign v869795 = BtoS_ACK0_p & v865fd7 | !BtoS_ACK0_p & v8702fe;
assign v850b88 = StoB_REQ1_p & v8587be | !StoB_REQ1_p & v8661ce;
assign v850ad2 = BtoS_ACK1_p & v865be6 | !BtoS_ACK1_p & v8657b3;
assign v870218 = jx1_p & v8702f2 | !jx1_p & v865698;
assign v8510be = jx0_p & v86c325 | !jx0_p & v86564e;
assign v86596b = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v8660f2;
assign v850819 = BtoS_ACK2_p & v844f99 | !BtoS_ACK2_p & !v844f99;
assign v87026f = StoB_REQ2_n & v8701ff | !StoB_REQ2_n & !v8702a8;
assign v865622 = StoB_REQ2_n & v850fb5 | !StoB_REQ2_n & !v86587f;
assign v865d46 = BtoS_ACK1_p & v86f080 | !BtoS_ACK1_p & v866137;
assign v8702d9 = RtoB_ACK0_p & v870225 | !RtoB_ACK0_p & !v87023b;
assign v865df6 = RtoB_ACK1_p & v84ff79 | !RtoB_ACK1_p & v866122;
assign v865644 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v870491;
assign jx0_n = v869795;
assign v870281 = stateG7_1_p & v8659c8 | !stateG7_1_p & v844fa9;
assign v865ae5 = BtoS_ACK1_p & v850b88 | !BtoS_ACK1_p & v865908;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v86b5d8 = StoB_REQ1_p & v8659d6 | !StoB_REQ1_p & !v865620;
assign BtoS_ACK0_n = v86dd82;
assign v870222 = DEQ_p & v844f91 | !DEQ_p & !v844f9f;
assign v851f5b = jx0_p & v87020f | !jx0_p & v870299;
assign v865623 = jx0_p & v870476 | !jx0_p & v865f6f;
assign v870333 = jx1_p & v865b52 | !jx1_p & v865b7c;
assign v865c36 = StoB_REQ2_p & v86f080 | !StoB_REQ2_p & !v8661c8;
assign v87022d = StoB_REQ0_p & v8657b4 | !StoB_REQ0_p & v86f0ad;
assign v865cbd = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v850b89;
assign v859822 = RtoB_ACK0_p & v844fa9 | !RtoB_ACK0_p & !v8702ed;
assign v8658a3 = StoB_REQ1_p & v8661c8 | !StoB_REQ1_p & v865d20;
assign v866122 = stateG7_0_p & v865660 | !stateG7_0_p & v865c3f;
assign v8659c8 = BtoR_REQ1_p & v844fa9 | !BtoR_REQ1_p & v86596b;
assign v8703f4 = StoB_REQ1_p & v8694e4 | !StoB_REQ1_p & v85dbed;
assign v865eee = StoB_REQ2_p & v865be6 | !StoB_REQ2_p & v865992;
assign v866108 = jx0_p & v844fb5 | !jx0_p & !v844f99;
assign v87022b = jx0_p & v865efd | !jx0_p & v870384;
assign v866093 = jx1_p & v870209 | !jx1_p & v850aee;
assign v8703ec = jx1_p & v85dbe6 | !jx1_p & v865920;
assign v865972 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v865791;
assign v87020f = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & v865caa;
assign v870259 = RtoB_ACK1_p & v844fa9 | !RtoB_ACK1_p & v870281;
assign v86c353 = StoB_REQ1_p & v865c36 | !StoB_REQ1_p & !v865d20;
assign v865d52 = StoB_REQ1_p & v8658dc | !StoB_REQ1_p & v870297;
assign v865dd3 = jx0_p & v865ae5 | !jx0_p & v858431;
assign v8702a3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8702bf;
assign v870299 = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & v86b5d5;
assign v865da4 = BtoS_ACK2_p & v865be6 | !BtoS_ACK2_p & v8658dc;
assign v865c6a = StoB_REQ2_p & v859822 | !StoB_REQ2_p & v865701;
assign v858630 = StoB_REQ1_p & v865da4 | !StoB_REQ1_p & v8702cb;
assign v870210 = StoB_REQ0_p & v865cf3 | !StoB_REQ0_p & v844f91;
assign v86dd82 = BtoS_ACK0_p & v844f95 | !BtoS_ACK0_p & !v870210;
assign v870526 = RtoB_ACK1_p & v844fb5 | !RtoB_ACK1_p & v870207;
assign v865920 = jx0_p & v8702a4 | !jx0_p & v8659c3;
assign v8702fd = jx0_p & v8702c8 | !jx0_p & v8660ef;
assign v85dbde = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8659de;
assign v850fb5 = RtoB_ACK0_p & v870235 | !RtoB_ACK0_p & !v86575b;
assign v85dbe6 = jx0_p & v8659c3 | !jx0_p & !v870484;
assign v8659bf = jx0_p & v865678 | !jx0_p & v865be6;
assign v853599 = jx0_p & v844f91 | !jx0_p & !v844f91;
assign v865c5b = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v865a28;
assign v86587c = stateG12_p & v844f9f | !stateG12_p & !v844f91;
assign v869783 = StoB_REQ2_p & v8702f6 | !StoB_REQ2_p & !v844f91;
assign v8703e0 = StoB_REQ1_p & v865be6 | !StoB_REQ1_p & v8658dc;
assign v8659c0 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v844fb3;
assign v865f6f = StoB_REQ1_p & v8702d9 | !StoB_REQ1_p & !v866158;
assign v865ce6 = StoB_REQ2_n & v8702f6 | !StoB_REQ2_n & !v8702a8;
assign v8702f8 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8702d9;
assign v8660c0 = jx0_p & v8702ca | !jx0_p & v844f91;
assign v865a3e = RtoB_ACK1_p & v8540cb | !RtoB_ACK1_p & v844f91;
assign v85a72b = jx0_p & v87056c | !jx0_p & v844f91;
assign v86575b = RtoB_ACK1_p & v86596b | !RtoB_ACK1_p & v844f91;
assign v865c02 = StoB_REQ2_p & v8701ff | !StoB_REQ2_p & !v844f91;
assign v865620 = StoB_REQ2_p & v865633 | !StoB_REQ2_p & v865972;
assign v865d41 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v86c352;
assign v8657e8 = BtoS_ACK1_p & v85dbde | !BtoS_ACK1_p & !v865fcf;
assign v86600c = jx1_p & v87030a | !jx1_p & !v865f8c;
assign v87045b = BtoR_REQ0_p & v870222 | !BtoR_REQ0_p & v844f91;
assign v8659bb = jx0_p & v87020f | !jx0_p & v87025e;
assign v8702a4 = StoB_REQ1_p & v865db0 | !StoB_REQ1_p & !v844f91;
assign v86f0bf = BtoS_ACK0_p & v865d0e | !BtoS_ACK0_p & v8657d5;
assign v8703a0 = StoB_REQ1_p & v87026a | !StoB_REQ1_p & v865cb0;
assign v87054a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v865f18;
assign v870225 = BtoR_REQ0_p & v870222 | !BtoR_REQ0_p & !v844f9f;
assign v865fbb = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8702d9;
assign v87056c = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8660d6;
assign v870207 = stateG7_0_p & v85dbf9 | !stateG7_0_p & v844fb5;
assign v859e32 = BtoS_ACK2_p & v844f99 | !BtoS_ACK2_p & !v844f91;
assign v854cf5 = BtoS_ACK1_p & v870283 | !BtoS_ACK1_p & v870245;
assign v85a24a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v87029c;
assign v866192 = BtoR_REQ0_p & v844fb3 | !BtoR_REQ0_p & v844f91;
assign v850277 = jx1_p & v8656be | !jx1_p & v865be6;
assign SLC1_n = v86c35a;
assign v86c352 = RtoB_ACK1_p & v844fa9 | !RtoB_ACK1_p & v865f25;
assign v865b94 = jx0_p & v844f97 | !jx0_p & !v844f91;
assign v858431 = BtoS_ACK1_p & v8703e0 | !BtoS_ACK1_p & v865da4;
assign v865d20 = StoB_REQ2_p & v865633 | !StoB_REQ2_p & v8702d0;
assign v8661ce = StoB_REQ2_p & v8587be | !StoB_REQ2_p & v858899;
assign v865c8f = jx1_p & v866128 | !jx1_p & v859aa5;
assign v865ff5 = stateG7_1_p & v844fa9 | !stateG7_1_p & v865857;
assign v8661e8 = jx0_p & v86573e | !jx0_p & v86586d;
assign v86c34e = jx0_p & v866044 | !jx0_p & v8659f1;
assign v8659d6 = StoB_REQ2_p & v86f080 | !StoB_REQ2_p & !v865633;
assign v865c64 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v865f25;
assign v86c31f = RtoB_ACK1_p & v865985 | !RtoB_ACK1_p & v866122;
assign v87029c = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8656bf;
assign v84fc5e = jx0_p & v865c36 | !jx0_p & v870321;
assign v865ccf = StoB_REQ2_p & v8656cd | !StoB_REQ2_p & v844fb5;
assign v8704d4 = BtoS_ACK1_p & v85dbe2 | !BtoS_ACK1_p & !v865c17;
assign v86575e = BtoS_ACK1_p & v86c353 | !BtoS_ACK1_p & v866121;
assign v865c69 = StoB_REQ1_p & v87034b | !StoB_REQ1_p & v865be6;
assign v865944 = StoB_REQ0_p & v865c91 | !StoB_REQ0_p & !v865f4b;
assign v865beb = RtoB_ACK1_p & v86596e | !RtoB_ACK1_p & v844f91;
assign v866121 = StoB_REQ1_p & v8659d6 | !StoB_REQ1_p & !v870341;
assign v8656a0 = BtoS_ACK2_p & v865849 | !BtoS_ACK2_p & v865620;
assign v865c17 = StoB_REQ2_n & v865f18 | !StoB_REQ2_n & !v87054a;
assign v865eff = BtoS_ACK1_p & v8702dc | !BtoS_ACK1_p & v865ba9;
assign v865908 = BtoS_ACK2_p & v870278 | !BtoS_ACK2_p & v8661ce;
assign v870246 = BtoS_ACK1_p & v8660ef | !BtoS_ACK1_p & !v865dd5;
assign v87031a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v865f3b;
assign v8540cb = BtoR_REQ1_p & v86596b | !BtoR_REQ1_p & v854981;
assign v8660ef = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v869783;
assign v8701ff = RtoB_ACK0_p & v870235 | !RtoB_ACK0_p & !v865a3e;
assign v8702bf = jx1_p & v865cf1 | !jx1_p & v8702fd;
assign v865f92 = DEQ_p & v844f91 | !DEQ_p & !v86587c;
assign v87029f = BtoS_ACK2_p & v865701 | !BtoS_ACK2_p & v8657f0;
assign v865821 = StoB_REQ0_p & v8705c0 | !StoB_REQ0_p & v86c316;
assign v865673 = BtoS_ACK1_p & v865644 | !BtoS_ACK1_p & !v865cb0;
assign v865992 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v870259;
assign v865701 = RtoB_ACK0_p & v844fa9 | !RtoB_ACK0_p & v859b38;
assign v865678 = BtoS_ACK1_p & v865be6 | !BtoS_ACK1_p & v86c356;
assign v86c356 = StoB_REQ1_p & v87029a | !StoB_REQ1_p & v865be6;
assign v865b8c = jx0_p & v85162c | !jx0_p & v844f91;
assign v865b7c = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v859e32;
assign v86f0aa = jx0_p & v865f6f | !jx0_p & !v870295;
assign v86596e = BtoR_REQ1_p & v85dbd8 | !BtoR_REQ1_p & v8705c8;
assign v851192 = StoB_REQ1_p & v8702a8 | !StoB_REQ1_p & v844f91;
assign v850b89 = RtoB_ACK0_p & v865833 | !RtoB_ACK0_p & !v865beb;
assign v86597b = StoB_REQ1_p & v8587be | !StoB_REQ1_p & v87034b;
assign v86571d = StoB_REQ1_p & v865a51 | !StoB_REQ1_p & !v867fda;
assign v85162c = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & !v844f97;
assign v865849 = StoB_REQ2_p & v8661c8 | !StoB_REQ2_p & v865972;
assign v865f25 = stateG7_0_p & v8702bc | !stateG7_0_p & v844fa9;
assign v870381 = StoB_REQ1_p & v865863 | !StoB_REQ1_p & !v866158;
assign v867fda = StoB_REQ2_n & v865c02 | !StoB_REQ2_n & !v844f91;
assign v865cd9 = jx0_p & v850ad2 | !jx0_p & v865fa1;
assign v870286 = BtoR_REQ0_p & v870222 | !BtoR_REQ0_p & !v844f91;
assign v8657f0 = StoB_REQ2_p & v8694e4 | !StoB_REQ2_p & v865701;
assign v8659dc = StoB_REQ1_p & v8587be | !StoB_REQ1_p & v865f98;
assign v8702f2 = jx0_p & v8704fd | !jx0_p & v865d52;
assign v865fa0 = StoB_REQ2_p & v8661c8 | !StoB_REQ2_p & v8702d0;
assign v85dbed = BtoS_ACK2_p & v865701 | !BtoS_ACK2_p & v865c6a;
assign v8585dc = StoB_REQ1_p & v8659d6 | !StoB_REQ1_p & !v86577a;
assign v865863 = StoB_REQ2_n & v8702d9 | !StoB_REQ2_n & !v865fbb;
assign v8702a2 = BtoS_ACK2_p & v865eee | !BtoS_ACK2_p & v8599b0;
assign v8658c7 = jx1_p & v86c34e | !jx1_p & v866044;
assign v87023b = RtoB_ACK1_p & v87048e | !RtoB_ACK1_p & v844f91;
assign BtoR_REQ0_n = !v865c20;
assign v870501 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v870222;
assign v865da6 = RtoB_ACK0_p & v865833 | !RtoB_ACK0_p & !v865632;
assign v865ff1 = jx0_p & v865bf0 | !jx0_p & v865858;
assign v8704fd = StoB_REQ1_p & v8661ce | !StoB_REQ1_p & v8599b0;
assign v865fd7 = StoB_REQ0_p & v870403 | !StoB_REQ0_p & v8703e2;
assign v8656cf = StoB_REQ0_p & v865bed | !StoB_REQ0_p & v865894;
assign v865cc1 = StoB_REQ2_p & v8661c8 | !StoB_REQ2_p & v85a24a;
assign v865698 = jx0_p & v865c69 | !jx0_p & v865be6;
assign v8702ca = BtoS_ACK1_p & v844fb5 | !BtoS_ACK1_p & v870290;
assign v865c91 = jx1_p & v865b94 | !jx1_p & !v844f91;
assign v865d0e = StoB_REQ0_p & v870269 | !StoB_REQ0_p & v865c8f;
assign v8702a6 = BtoS_ACK2_p & v844f99 | !BtoS_ACK2_p & v869783;
assign v87028c = StoB_REQ2_p & v865f18 | !StoB_REQ2_p & !v844f91;
assign v844fb5 = stateG12_p & v844f91 | !stateG12_p & !v844f91;
assign v865894 = jx1_p & v8510be | !jx1_p & v8659bf;
assign v865632 = RtoB_ACK1_p & v85dbd8 | !RtoB_ACK1_p & v844f91;
assign v865f98 = StoB_REQ2_p & v8587be | !StoB_REQ2_p & v870277;
assign v8702e1 = StoB_REQ1_p & v865be6 | !StoB_REQ1_p & v870297;
assign v8702bc = stateG7_1_p & v844f91 | !stateG7_1_p & v844fa9;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v8702ce = jx1_p & v8694ff | !jx1_p & v865ff1;
assign v870356 = StoB_REQ1_p & v859e32 | !StoB_REQ1_p & v8702a6;
assign v870245 = StoB_REQ1_p & v8694e4 | !StoB_REQ1_p & v87029f;
assign v844f9f = FULL_p & v844f91 | !FULL_p & !v844f91;
assign v870200 = BtoS_ACK1_p & v8658a3 | !BtoS_ACK1_p & !v8585dc;
assign v87020c = stateG7_1_p & v844fa9 | !stateG7_1_p & v866204;
assign v8587be = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v870229;
assign v86b5d5 = StoB_REQ1_p & v865ce6 | !StoB_REQ1_p & !v844f91;
assign v86b5b5 = StoB_REQ1_p & v8657f0 | !StoB_REQ1_p & v865c6a;
assign v865f3c = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v844fa9;
assign v866128 = jx0_p & v86b5d8 | !jx0_p & v859aa5;
assign v865985 = BtoR_REQ1_p & v8659c0 | !BtoR_REQ1_p & v844f91;
assign v86c325 = BtoS_ACK1_p & v850173 | !BtoS_ACK1_p & v865817;
assign v86587f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v865da6;
assign v870467 = BtoS_ACK2_p & v87026f | !BtoS_ACK2_p & v870284;
assign v86577a = BtoS_ACK2_p & v865fa0 | !BtoS_ACK2_p & v865d20;
assign v870348 = BtoS_ACK1_p & v866137 | !BtoS_ACK1_p & v8659d6;
assign v870214 = BtoS_ACK1_p & v865644 | !BtoS_ACK1_p & !v8703a0;
assign v865989 = stateG7_1_p & v844f91 | !stateG7_1_p & v866204;
assign v870292 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8656f8;
assign v865791 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v859f24;
assign v86b5e3 = BtoS_ACK0_p & v8694ed | !BtoS_ACK0_p & !v865b07;
assign v8657ee = jx1_p & v8659f1 | !jx1_p & v85984b;
assign v865981 = BtoS_ACK1_p & v8660ef | !BtoS_ACK1_p & !v870356;
assign v865d79 = BtoS_ACK1_p & v858042 | !BtoS_ACK1_p & v850819;
assign v850031 = BtoS_ACK1_p & v86c353 | !BtoS_ACK1_p & v8585dc;
assign v86c316 = jx1_p & v865c46 | !jx1_p & v866139;
assign v8658dc = StoB_REQ2_p & v865c64 | !StoB_REQ2_p & v865be6;
assign v865db0 = RtoB_ACK0_p & v866192 | !RtoB_ACK0_p & v86c31f;
assign v86c319 = StoB_REQ1_p & v865c17 | !StoB_REQ1_p & !v866158;
assign v870403 = jx1_p & v866108 | !jx1_p & !v853599;
assign v865f8c = jx0_p & v85162c | !jx0_p & !v844f91;
assign v8702dc = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8660c2;
assign v8703e9 = BtoS_ACK1_p & v85a1b8 | !BtoS_ACK1_p & v870531;
assign v86f080 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v865c92;
assign v865cf3 = jx1_p & v8661e8 | !jx1_p & v870257;
assign v865884 = StoB_REQ0_p & v8657ee | !StoB_REQ0_p & v8658c7;
assign v870297 = StoB_REQ2_p & v865d41 | !StoB_REQ2_p & v865be6;
assign v859b38 = RtoB_ACK1_p & v865f3c | !RtoB_ACK1_p & v844f91;
assign SLC0_n = (BtoS_ACK0_n & ((SLC1_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n))) | (!StoB_REQ2_n)))))));
assign ENQ_n = (BtoS_ACK0_n & ((StoB_REQ0_n & ((!SLC1_n))))) | (!BtoS_ACK0_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((SLC1_n)))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  jx0_p = 0;
  jx1_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
