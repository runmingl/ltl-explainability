module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hbusreq2, hlock2, hbusreq3, hlock3, hburst0, hburst1, hmaster0, hmaster1, hmastlock, start, decide, locked, hgrant0, hgrant1, hgrant2, hgrant3, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, stateG10_2, stateG10_3, jx0, jx1, jx2);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v84563c;
  wire v845654;
  wire v8e1935;
  wire b26692;
  wire b26693;
  wire v84566c;
  wire b26694;
  wire b26695;
  wire b26696;
  wire b26697;
  wire b26698;
  wire b26699;
  wire b2669a;
  wire b2669b;
  wire b2669c;
  wire b2669d;
  wire b2669e;
  wire b2669f;
  wire b266a0;
  wire b266a1;
  wire b266a2;
  wire b266a3;
  wire b266a4;
  wire b266a5;
  wire b266a6;
  wire b266a7;
  wire b266a8;
  wire b266a9;
  wire b266aa;
  wire b266ab;
  wire b266ac;
  wire b266ad;
  wire b266ae;
  wire b266af;
  wire b266b0;
  wire b266b1;
  wire b266b2;
  wire b266b3;
  wire b266b4;
  wire b266b5;
  wire b266b6;
  wire b266b7;
  wire b266b8;
  wire b266b9;
  wire b266ba;
  wire b266bb;
  wire b266bc;
  wire b266bd;
  wire b266be;
  wire b266bf;
  wire b266c0;
  wire b266c1;
  wire b266c2;
  wire b266c3;
  wire b266c4;
  wire b266ca;
  wire b266cb;
  wire b266cc;
  wire b266cd;
  wire b266d2;
  wire b266d3;
  wire b266d4;
  wire b266d5;
  wire b266d6;
  wire b266da;
  wire b266db;
  wire b266dc;
  wire b266df;
  wire b266e0;
  wire b266e1;
  wire b266e2;
  wire b266e3;
  wire b266e4;
  wire b266e5;
  wire b266e6;
  wire b266e7;
  wire b266ed;
  wire b266ee;
  wire b266ef;
  wire b266f0;
  wire b266f1;
  wire b266f2;
  wire b266fa;
  wire b266fb;
  wire b266fc;
  wire b266fd;
  wire b266fe;
  wire b266ff;
  wire b26700;
  wire b26701;
  wire b26702;
  wire b26703;
  wire b26704;
  wire b26705;
  wire b26706;
  wire b26707;
  wire b26708;
  wire b26709;
  wire b2670a;
  wire b2670b;
  wire b2670c;
  wire b2670d;
  wire b2670e;
  wire b2670f;
  wire b26710;
  wire b26711;
  wire b26712;
  wire b26713;
  wire b26714;
  wire b26715;
  wire b26716;
  wire b26717;
  wire b26718;
  wire b26719;
  wire b2671a;
  wire b2671b;
  wire b2671c;
  wire b2671d;
  wire b2671e;
  wire b2671f;
  wire b26720;
  wire b26721;
  wire b26722;
  wire b26723;
  wire b26724;
  wire b26725;
  wire b26726;
  wire b26727;
  wire b26728;
  wire b26729;
  wire b2672a;
  wire b2672b;
  wire b2672c;
  wire b2672d;
  wire b2672e;
  wire b2672f;
  wire b26730;
  wire b26731;
  wire b26732;
  wire b26733;
  wire b26734;
  wire b26735;
  wire b26736;
  wire b26737;
  wire b26738;
  wire b26739;
  wire b2673a;
  wire b2673b;
  wire b2673c;
  wire b2673d;
  wire b2673e;
  wire b2673f;
  wire b26740;
  wire b26741;
  wire b26742;
  wire b26743;
  wire b26744;
  wire b26745;
  wire b26746;
  wire b26747;
  wire b26748;
  wire b26749;
  wire b2674a;
  wire b2674b;
  wire b2674c;
  wire b2674d;
  wire b2674e;
  wire b2674f;
  wire b26750;
  wire b26751;
  wire b26752;
  wire b26753;
  wire b26754;
  wire b26755;
  wire b26756;
  wire b26757;
  wire b26758;
  wire b26759;
  wire b2675a;
  wire b2675b;
  wire b2675c;
  wire b2675d;
  wire b2675e;
  wire b2675f;
  wire b26760;
  wire b26761;
  wire b26762;
  wire b26763;
  wire b26764;
  wire b26765;
  wire b26766;
  wire b26767;
  wire b26768;
  wire b26769;
  wire b2676a;
  wire b2676b;
  wire b2676c;
  wire b2676d;
  wire b2676e;
  wire b2676f;
  wire b26770;
  wire b26771;
  wire b26772;
  wire b26773;
  wire b26774;
  wire b26775;
  wire b26776;
  wire b26777;
  wire b26778;
  wire b26779;
  wire b2677a;
  wire b2677b;
  wire b2677c;
  wire b2677d;
  wire b2677e;
  wire b2677f;
  wire b26780;
  wire b26781;
  wire b26782;
  wire b26783;
  wire b26784;
  wire b26785;
  wire b26786;
  wire b26787;
  wire b26788;
  wire b26789;
  wire b2678a;
  wire b2678b;
  wire b2678c;
  wire b2678d;
  wire b2678e;
  wire v84564a;
  wire be34df;
  wire be34e5;
  wire be34e6;
  wire be34e7;
  wire be34e8;
  wire be34e9;
  wire be34ea;
  wire v845646;
  wire v8c6711;
  wire c98b95;
  wire c98b96;
  wire c98b9e;
  wire c98b9f;
  wire c98ba0;
  wire c98ba1;
  wire c98ba2;
  wire c98ba3;
  wire c98ba4;
  wire v845658;
  wire v9269ad;
  wire v8565cf;
  wire b8acd7;
  wire b8acd8;
  wire b8acd9;
  wire b8acda;
  wire b8acdb;
  wire b8acdc;
  wire b8acdf;
  wire b8ace0;
  wire b8ace1;
  wire b8ace2;
  wire b8ace3;
  wire b8ace4;
  wire b8ace5;
  wire b8ace6;
  wire b8ace7;
  wire b8ace8;
  wire b8ace9;
  wire b8acea;
  wire b8aceb;
  wire b8acec;
  wire b8aced;
  wire b8acee;
  wire b8acef;
  wire b8acf0;
  wire b8acf1;
  wire b8acf2;
  wire b8acf3;
  wire b8acf4;
  wire a81ca6;
  wire v845670;
  wire c07311;
  wire a81ca7;
  wire a81ca8;
  wire a81ca9;
  wire a81caa;
  wire a81cab;
  wire a81cac;
  wire a81cad;
  wire a81cae;
  wire v845672;
  wire a81caf;
  wire a81cb0;
  wire a81cb1;
  wire a81cb2;
  wire a81cb3;
  wire a81cb4;
  wire a81cb5;
  wire a81cb6;
  wire a81cc0;
  wire a81cc1;
  wire a81cc2;
  wire a81cc3;
  wire a81cc4;
  wire a81cc5;
  wire a81cc6;
  wire a81cc7;
  wire a81cc8;
  wire a81cc9;
  wire a81cca;
  wire a81ccb;
  wire a81ccc;
  wire a81ccd;
  wire a81cce;
  wire a81ccf;
  wire a81cd0;
  wire a81cd1;
  wire a81cd2;
  wire a81cd3;
  wire a81cd4;
  wire a81cd5;
  wire a81cd6;
  wire a81cd7;
  wire a81cd8;
  wire a81cd9;
  wire a81cda;
  wire a81cdb;
  wire a81cdc;
  wire a81cdd;
  wire a81cde;
  wire a81cdf;
  wire a81ce0;
  wire a81ce1;
  wire a81ce2;
  wire a81ce3;
  wire a81ce4;
  wire a81ce5;
  wire a81ce6;
  wire a81ce7;
  wire a81ce8;
  wire a81ce9;
  wire a81cea;
  wire a81ceb;
  wire a81cec;
  wire a81ced;
  wire a81cee;
  wire a81cef;
  wire a81cf0;
  wire a81cf1;
  wire a81cf2;
  wire a81cf3;
  wire a81cf4;
  wire a81cf5;
  wire a81cf6;
  wire a81cf7;
  wire a81cf8;
  wire a81cf9;
  wire a81cfa;
  wire a81cfb;
  wire a81cfc;
  wire a81cfd;
  wire a81cfe;
  wire a81cff;
  wire a81d00;
  wire a81d01;
  wire a81d02;
  wire a81d03;
  wire a81d04;
  wire a81d05;
  wire a81d06;
  wire a81d07;
  wire a81d08;
  wire a81d09;
  wire a81d0a;
  wire a81d0b;
  wire a81d0c;
  wire a81d0d;
  wire v845656;
  wire a57858;
  wire v845666;
  wire a57859;
  wire a5785a;
  wire a5785b;
  wire v84566e;
  wire v9703fa;
  wire v9703fb;
  wire v9703fc;
  wire v9703fd;
  wire v9703fe;
  wire v9703ff;
  wire v970400;
  wire v970401;
  wire v970407;
  wire v970408;
  wire v970409;
  wire v97040a;
  wire v97040b;
  wire v970413;
  wire v970416;
  wire v970420;
  wire v970421;
  wire v970429;
  wire v97042a;
  wire v97042b;
  wire v97042c;
  wire v97042d;
  wire v97042e;
  wire v97042f;
  wire v970430;
  wire v970431;
  wire v970432;
  wire v970433;
  wire v970434;
  wire v970435;
  wire v970436;
  wire v970437;
  wire v970438;
  wire v970439;
  wire v97043a;
  wire v97043b;
  wire v97043c;
  wire v97043d;
  wire v97043e;
  wire v97043f;
  wire v970440;
  wire v970441;
  wire v970442;
  wire v970443;
  wire v970444;
  wire v970445;
  wire v970446;
  wire v970447;
  wire v970448;
  wire v970449;
  wire v97044a;
  wire v97044b;
  wire v97044c;
  wire v97044d;
  wire v97044e;
  wire v97044f;
  wire v970450;
  wire v970451;
  wire v970452;
  wire v970453;
  wire v970454;
  wire v970455;
  wire v970456;
  wire v970457;
  wire v970458;
  wire v970459;
  wire v97045a;
  wire v97045b;
  wire v97045c;
  wire v97045d;
  wire c06d34;
  wire d40d29;
  wire d40d2a;
  wire d40d2b;
  wire d40d2c;
  wire d40d2d;
  wire d40d2e;
  wire v845674;
  wire bfbd18;
  wire bfbd19;
  wire d40d2f;
  wire d40d30;
  wire d40d31;
  wire d40d32;
  wire d40d33;
  wire d40d34;
  wire d40d35;
  wire d40d36;
  wire d40d3a;
  wire d40d3b;
  wire d40d3c;
  wire d40d3d;
  wire d40d3e;
  wire d40d41;
  wire d40d42;
  wire d40d43;
  wire d40d44;
  wire d40d45;
  wire d40d46;
  wire d40d47;
  wire d40d48;
  wire d40d4e;
  wire d40d4f;
  wire d40d50;
  wire d40d51;
  wire d40d52;
  wire d40d53;
  wire d40d54;
  wire d40d55;
  wire d40d56;
  wire d40d57;
  wire d40d58;
  wire d40d59;
  wire d40d5a;
  wire d40d5b;
  wire d40d5c;
  wire d40d60;
  wire d40d61;
  wire d40d62;
  wire d40d63;
  wire d40d64;
  wire d40d66;
  wire d40d67;
  wire d40d68;
  wire d40d69;
  wire d40d6a;
  wire d40d6b;
  wire d40d6c;
  wire d40d6d;
  wire d40d6e;
  wire d40d6f;
  wire d40d70;
  wire d40d71;
  wire d40d72;
  wire d40d73;
  wire d40d74;
  wire d40d75;
  wire d40d76;
  wire d40d77;
  wire d40d78;
  wire d40d79;
  wire d40d7a;
  wire d40d7b;
  wire d40d7c;
  wire d40d7d;
  wire d40d7e;
  wire d40d7f;
  wire d40d80;
  wire d40d81;
  wire d40d82;
  wire d40d83;
  wire d40d84;
  wire d40d85;
  wire d40d86;
  wire d40d87;
  wire d40d88;
  wire d40d89;
  wire d40d8a;
  wire d40d8b;
  wire d40d8c;
  wire d40d8d;
  wire d40d8e;
  wire d40d8f;
  wire d40d90;
  wire d40d91;
  wire d40d92;
  wire d40d93;
  wire d40d94;
  wire d40d95;
  wire d40d96;
  wire d40d97;
  wire d40d98;
  wire d40d99;
  wire d40d9a;
  wire d40d9b;
  wire d40d9c;
  wire d40d9d;
  wire v845660;
  wire deac0f;
  wire deac10;
  wire deac11;
  wire v84565a;
  wire deac17;
  wire deac18;
  wire deac19;
  wire deac1e;
  wire deac1f;
  wire deac20;
  wire deac2a;
  wire deac34;
  wire deac3e;
  wire deac3f;
  wire v845652;
  wire deac4a;
  wire v8c6449;
  wire deac4b;
  wire deac4c;
  wire deac4d;
  wire deac4e;
  wire deac4f;
  wire deac50;
  wire deac51;
  wire deac52;
  wire deac53;
  wire deac54;
  wire deac55;
  wire deac56;
  wire deac57;
  wire deac5a;
  wire deac5b;
  wire deac5c;
  wire deac5d;
  wire deac5f;
  wire deac60;
  wire deac61;
  wire deac62;
  wire deac63;
  wire deac64;
  wire deac6a;
  wire deac6b;
  wire deac6c;
  wire deac71;
  wire deac72;
  wire deac78;
  wire deac79;
  wire deac7a;
  wire deac7b;
  wire deac7c;
  wire deac7d;
  wire deac7e;
  wire deac86;
  wire deac87;
  wire deac88;
  wire deac89;
  wire deac99;
  wire deac9a;
  wire deac9b;
  wire deac9c;
  wire deac9d;
  wire deac9e;
  wire deac9f;
  wire v8c607d;
  wire deaca0;
  wire deaca1;
  wire deaca2;
  wire deacaa;
  wire deacab;
  wire deacac;
  wire deacad;
  wire deacae;
  wire deacaf;
  wire deacb0;
  wire deacb1;
  wire deacb2;
  wire deacb3;
  wire deacb4;
  wire deacb5;
  wire deacb6;
  wire deacb7;
  wire deacb8;
  wire deacbc;
  wire deacbd;
  wire deacbe;
  wire deacbf;
  wire deacc0;
  wire deacc1;
  wire deacc2;
  wire deacc3;
  wire deacc4;
  wire deacc5;
  wire deacd2;
  wire deacd3;
  wire deacd4;
  wire deacd5;
  wire deacd6;
  wire deacd7;
  wire deacd8;
  wire deacd9;
  wire deacda;
  wire deacdb;
  wire deacdc;
  wire deacdd;
  wire deacde;
  wire deacdf;
  wire deace0;
  wire deace1;
  wire deace2;
  wire deace3;
  wire deace4;
  wire deace5;
  wire deace6;
  wire deace7;
  wire deace8;
  wire deace9;
  wire deacea;
  wire deaceb;
  wire deacec;
  wire deaced;
  wire deacee;
  wire deacef;
  wire deacf0;
  wire deacf1;
  wire deacf2;
  wire deacf3;
  wire deacf4;
  wire deacf5;
  wire deacf6;
  wire deacf7;
  wire deacf8;
  wire deacf9;
  wire deacfa;
  wire deacfb;
  wire deacfc;
  wire deacfd;
  wire deacfe;
  wire deacff;
  wire dead00;
  wire dead01;
  wire dead02;
  wire dead03;
  wire dead04;
  wire dead05;
  wire dead06;
  wire dead07;
  wire dead08;
  wire dead09;
  wire dead0a;
  wire dead0b;
  wire dead0c;
  wire dead0d;
  wire dead0e;
  wire dead0f;
  wire dead10;
  wire dead11;
  wire dead12;
  wire dead13;
  wire dead14;
  wire dead15;
  wire dead16;
  wire dead17;
  wire dead18;
  wire dead19;
  wire dead1a;
  wire dead1b;
  wire dead1c;
  wire dead1d;
  wire dead20;
  wire dead21;
  wire dead22;
  wire dead23;
  wire dead24;
  wire dead25;
  wire dead26;
  wire dead27;
  wire dead28;
  wire dead29;
  wire dead2a;
  wire dead2b;
  wire dead2c;
  wire dead2d;
  wire dead2e;
  wire dead2f;
  wire dead30;
  wire dead31;
  wire dead32;
  wire dead33;
  wire dead34;
  wire dead35;
  wire dead36;
  wire dead37;
  wire dead38;
  wire dead39;
  wire dead3a;
  wire dead3b;
  wire dead3c;
  wire dead3d;
  wire dead3e;
  wire dead3f;
  wire dead40;
  wire dead41;
  wire dead42;
  wire dead43;
  wire dead44;
  wire dead45;
  wire dead46;
  wire dead47;
  wire dead48;
  wire dead49;
  wire dead4a;
  wire dead4b;
  wire dead4c;
  wire dead4d;
  wire dead4e;
  wire dead4f;
  wire dead50;
  wire dead51;
  wire dead52;
  wire v845644;
  wire dead53;
  wire dead54;
  wire dead55;
  wire dead56;
  wire dead57;
  wire dead5e;
  wire dead5f;
  wire dead60;
  wire dead61;
  wire dead62;
  wire dead63;
  wire dead64;
  wire dead65;
  wire dead66;
  wire dead67;
  wire dead68;
  wire dead69;
  wire dead6a;
  wire dead6b;
  wire dead6c;
  wire dead6d;
  wire dead6e;
  wire dead6f;
  wire dead70;
  wire dead71;
  wire dead72;
  wire dead73;
  wire dead74;
  wire dead75;
  wire dead76;
  wire dead77;
  wire dead78;
  wire dead79;
  wire dead7a;
  wire dead7b;
  wire dead7c;
  wire dead7d;
  wire dead7e;
  wire dead7f;
  wire dead80;
  wire dead81;
  wire dead82;
  wire dead83;
  wire dead84;
  wire dead85;
  wire dead86;
  wire dead87;
  wire dead88;
  wire dead89;
  wire dead8a;
  wire dead8b;
  wire dead8c;
  wire dead8d;
  wire dead8e;
  wire dead8f;
  wire dead90;
  wire dead91;
  wire dead92;
  wire dead93;
  wire dead94;
  wire dead95;
  wire dead96;
  wire dead97;
  wire dead98;
  wire dead99;
  wire dead9a;
  wire dead9b;
  wire dead9c;
  wire dead9d;
  wire dead9e;
  wire dead9f;
  wire deada0;
  wire deada6;
  wire deada7;
  wire deada8;
  wire deada9;
  wire deadaa;
  wire deadab;
  wire deadac;
  wire deadb1;
  wire deadb2;
  wire deadb3;
  wire deadb4;
  wire deadb5;
  wire deadb9;
  wire deadba;
  wire deadbb;
  wire deadbc;
  wire deadbd;
  wire deadbe;
  wire deadc3;
  wire deadc4;
  wire deadc5;
  wire deadc6;
  wire deadc7;
  wire deadc8;
  wire deadc9;
  wire deadca;
  wire deadcb;
  wire deadcc;
  wire deadcd;
  wire deadce;
  wire deadcf;
  wire deadd0;
  wire deadd1;
  wire deadd2;
  wire deadd3;
  wire deadd4;
  wire deadd5;
  wire deadd6;
  wire deadd7;
  wire deadd8;
  wire deadd9;
  wire deadda;
  wire deaddb;
  wire deaddc;
  wire deadde;
  wire deaddf;
  wire deade0;
  wire deade1;
  wire deade2;
  wire deade3;
  wire deade4;
  wire deade5;
  wire deadea;
  wire deadeb;
  wire deadec;
  wire deaded;
  wire deadee;
  wire deadef;
  wire deadf0;
  wire deadf1;
  wire deadf2;
  wire deadf3;
  wire deadf4;
  wire deadf5;
  wire deadf6;
  wire deadf7;
  wire deadf8;
  wire deadf9;
  wire deadfa;
  wire deadfb;
  wire deadfc;
  wire deadfd;
  wire deadfe;
  wire deadff;
  wire deae00;
  wire deae01;
  wire deae02;
  wire deae03;
  wire deae04;
  wire deae05;
  wire deae06;
  wire deae07;
  wire deae08;
  wire deae09;
  wire deae0a;
  wire deae0b;
  wire deae0c;
  wire deae0d;
  wire deae0e;
  wire deae0f;
  wire deae10;
  wire deae11;
  wire deae12;
  wire deae13;
  wire deae14;
  wire deae15;
  wire deae16;
  wire deae17;
  wire deae18;
  wire deae19;
  wire deae1a;
  wire deae1b;
  wire deae1c;
  wire deae1d;
  wire deae1e;
  wire deae1f;
  wire deae20;
  wire deae21;
  wire deae22;
  wire deae23;
  wire deae24;
  wire deae25;
  wire deae26;
  wire deae27;
  wire deae28;
  wire deae29;
  wire deae2a;
  wire deae2b;
  wire deae2c;
  wire deae2d;
  wire deae2e;
  wire deae2f;
  wire deae30;
  wire deae31;
  wire deae32;
  wire deae33;
  wire deae34;
  wire deae35;
  wire deae36;
  wire deae37;
  wire deae38;
  wire deae39;
  wire deae3a;
  wire deae3b;
  wire deae3c;
  wire deae3d;
  wire deae3e;
  wire deae40;
  wire deae41;
  wire deae42;
  wire deae43;
  wire deae44;
  wire deae45;
  wire deae46;
  wire deae47;
  wire deae48;
  wire deae49;
  wire deae4a;
  wire deae4b;
  wire deae4c;
  wire deae4d;
  wire deae4e;
  wire deae4f;
  wire deae50;
  wire deae51;
  wire deae52;
  wire deae53;
  wire deae54;
  wire deae55;
  wire deae56;
  wire deae57;
  wire deae58;
  wire deae59;
  wire deae5a;
  wire deae5b;
  wire deae5c;
  wire deae5d;
  wire deae5e;
  wire deae5f;
  wire deae60;
  wire deae61;
  wire deae62;
  wire deae63;
  wire deae64;
  wire deae65;
  wire deae66;
  wire deae67;
  wire deae68;
  wire deae69;
  wire deae6a;
  wire deae6b;
  wire deae6c;
  wire deae6d;
  wire deae6e;
  wire deae6f;
  wire deae70;
  wire deae74;
  wire deae75;
  wire deae76;
  wire deae79;
  wire deae7a;
  wire deae7b;
  wire deae7f;
  wire deae80;
  wire deae81;
  wire deae86;
  wire deae87;
  wire deae88;
  wire deae89;
  wire deae8a;
  wire deae8b;
  wire deae8c;
  wire deae8d;
  wire deae8e;
  wire deae8f;
  wire deae90;
  wire deae91;
  wire deae92;
  wire deae93;
  wire deae94;
  wire deae95;
  wire deae96;
  wire deae97;
  wire deae98;
  wire deae99;
  wire deae9a;
  wire deae9b;
  wire deae9c;
  wire deae9d;
  wire deaea1;
  wire deaea2;
  wire deaea3;
  wire deaea4;
  wire deaea5;
  wire deaea6;
  wire deaea7;
  wire deaea8;
  wire deaea9;
  wire deaeaa;
  wire deaeab;
  wire deaeac;
  wire deaead;
  wire deaeae;
  wire deaeaf;
  wire deaeb0;
  wire deaeb1;
  wire deaeb2;
  wire deaeb3;
  wire deaeb4;
  wire deaeb5;
  wire deaeb6;
  wire dea6b9;
  wire dea6ba;
  wire dea6bb;
  wire dea6bc;
  wire dea6bd;
  wire dea6be;
  wire dea6bf;
  wire dea6c0;
  wire dea6c1;
  wire dea6c2;
  wire dea6c3;
  wire dea6c4;
  wire dea6c5;
  wire dea6c6;
  wire dea6c7;
  wire dea6c8;
  wire dea6c9;
  wire dea6ca;
  wire dea6cb;
  wire dea6cc;
  wire dea6cd;
  wire dea6ce;
  wire dea6cf;
  wire dea6d0;
  wire dea6d1;
  wire dea6d2;
  wire dea6d3;
  wire dea6d4;
  wire dea6d5;
  wire dea6d6;
  wire dea6d7;
  wire dea6d8;
  wire dea6d9;
  wire dea6da;
  wire dea6db;
  wire dea6dc;
  wire dea6dd;
  wire dea6de;
  wire dea6df;
  wire dea6e0;
  wire dea6e1;
  wire dea6e2;
  wire dea6e3;
  wire dea6e4;
  wire dea6e5;
  wire dea6ea;
  wire dea6eb;
  wire dea6ec;
  wire dea6ed;
  wire dea6ee;
  wire dea6ef;
  wire dea6f0;
  wire dea6f1;
  wire dea6f2;
  wire dea6f3;
  wire dea6f4;
  wire dea6f5;
  wire dea6f6;
  wire dea6f7;
  wire dea6f8;
  wire dea6f9;
  wire dea6fa;
  wire dea6fb;
  wire dea6fc;
  wire dea6fd;
  wire dea6fe;
  wire dea6ff;
  wire dea700;
  wire dea701;
  wire dea724;
  wire dea725;
  wire dea726;
  wire dea727;
  wire dea728;
  wire dea729;
  wire dea72b;
  wire dea72c;
  wire dea72d;
  wire dea72e;
  wire dea72f;
  wire dea730;
  wire dea731;
  wire dea732;
  wire dea733;
  wire dea734;
  wire dea735;
  wire dea736;
  wire dea737;
  wire dea738;
  wire dea739;
  wire dea73d;
  wire dea743;
  wire dea744;
  wire dea745;
  wire dea746;
  wire dea747;
  wire dea748;
  wire dea749;
  wire dea74a;
  wire dea74b;
  wire dea74c;
  wire dea74d;
  wire dea74e;
  wire dea74f;
  wire dea750;
  wire dea751;
  wire dea752;
  wire dea753;
  wire dea757;
  wire dea758;
  wire dea759;
  wire dea75a;
  wire dea75b;
  wire dea75c;
  wire dea75d;
  wire dea75e;
  wire dea75f;
  wire dea760;
  wire dea761;
  wire dea762;
  wire dea763;
  wire dea764;
  wire dea765;
  wire dea766;
  wire dea767;
  wire dea768;
  wire dea769;
  wire dea76a;
  wire dea76b;
  wire dea76c;
  wire dea76d;
  wire dea76e;
  wire dea76f;
  wire dea782;
  wire dea784;
  wire dea785;
  wire dea786;
  wire dea787;
  wire dea788;
  wire dea789;
  wire dea78a;
  wire dea78b;
  wire dea79b;
  wire dea79c;
  wire dea79d;
  wire dea79e;
  wire dea79f;
  wire dea7a0;
  wire dea7a1;
  wire dea7a2;
  wire dea7a3;
  wire dea7a6;
  wire dea7a7;
  wire dea7a8;
  wire dea7a9;
  wire dea7aa;
  wire dea7ab;
  wire dea7ac;
  wire dea7ad;
  wire dea7ae;
  wire dea7b3;
  wire dea7b4;
  wire dea7b5;
  wire cea85c;
  wire cea85d;
  wire cea85e;
  wire cea85f;
  wire cea860;
  wire cea861;
  wire cea862;
  wire cea86c;
  wire cea86d;
  wire cea86e;
  wire cea86f;
  wire cea877;
  wire cea878;
  wire cea879;
  wire cea883;
  wire cea884;
  wire cea887;
  wire cea888;
  wire cea889;
  wire cea88d;
  wire cea89c;
  wire cea89d;
  wire cea89e;
  wire cea89f;
  wire cea8a0;
  wire cea8a1;
  wire cea8a2;
  wire cea8a3;
  wire cea8a4;
  wire cea8a7;
  wire cea8a8;
  wire cea8a9;
  wire cea8aa;
  wire cea8ab;
  wire cea8ac;
  wire cea8ad;
  wire cea8ae;
  wire cea0b5;
  wire cea0b6;
  wire cea0b7;
  wire cea0b8;
  wire cea0b9;
  wire cea0ba;
  wire cea0bb;
  wire cea0bc;
  wire cea0bd;
  wire cea0be;
  wire cea0bf;
  wire cea0c0;
  wire cea0c1;
  wire cea0c2;
  wire cea0ca;
  wire cea0d2;
  wire cea0d3;
  wire cea0d4;
  wire cea0d5;
  wire cea0d6;
  wire cea0d7;
  wire cea0e7;
  wire cea0e8;
  wire cea0e9;
  wire cea0ee;
  wire cea0ef;
  wire cea0f0;
  wire cea0f1;
  wire cea0f2;
  wire cea0f3;
  wire cea0f4;
  wire cea148;
  wire cea149;
  wire cea14a;
  wire cea14b;
  wire cea14c;
  wire cea14d;
  wire cea14e;
  wire cea14f;
  wire cea150;
  wire cea151;
  wire cea152;
  wire cea153;
  wire cea154;
  wire cea155;
  wire cea156;
  wire cea157;
  wire cea158;
  wire cea159;
  wire cea15a;
  wire cea15b;
  wire cea15c;
  wire cea15d;
  wire cea15e;
  wire cea15f;
  wire cea160;
  wire cea161;
  wire cea162;
  wire cea163;
  wire cea164;
  wire cea165;
  wire cea166;
  wire cea167;
  wire cea168;
  wire cea169;
  wire cea16a;
  wire cea16b;
  wire cea16c;
  wire cea16d;
  wire cea16e;
  wire cea16f;
  wire cea170;
  wire cea171;
  wire cea172;
  wire cea173;
  wire cea174;
  wire cea175;
  wire cea176;
  wire cea177;
  wire cea178;
  wire cea179;
  wire cea17a;
  wire cea17b;
  wire cea17c;
  wire cea17d;
  wire cea17e;
  wire cea17f;
  wire cea180;
  wire cea181;
  wire cea182;
  wire cea183;
  wire cea184;
  wire cea187;
  wire cea188;
  wire cea189;
  wire cea18a;
  wire cea18b;
  wire cea18c;
  wire v845648;
  wire cea18d;
  wire cea18e;
  wire cea18f;
  wire cea190;
  wire cea191;
  wire cea192;
  wire cea193;
  wire cea194;
  wire cea195;
  wire cea196;
  wire cea197;
  wire cea198;
  wire cea199;
  wire cea19a;
  wire cea19b;
  wire cea19c;
  wire cea19d;
  wire cea19e;
  wire cea19f;
  wire cea1a0;
  wire cea1a1;
  wire cea1a2;
  wire cea1a3;
  wire cea1a4;
  wire cea1a5;
  wire cea1a6;
  wire cea1a7;
  wire cea1a8;
  wire cea1a9;
  wire cea1aa;
  wire cea1ab;
  wire cea1ac;
  wire cea1ad;
  wire cea1ae;
  wire cea1af;
  wire cea1b0;
  wire cea1b1;
  wire cea1b2;
  wire cea1b3;
  wire cea1b4;
  wire cea1b5;
  wire cea1b6;
  wire cea1b7;
  wire cea1b8;
  wire cea1b9;
  wire cea1ba;
  wire cea1bb;
  wire cea1bc;
  wire cea1bd;
  wire cea1be;
  wire cea1bf;
  wire cea1c0;
  wire cea1c1;
  wire cea1c2;
  wire cea1c3;
  wire cea1c4;
  wire cea1c5;
  wire cea1c6;
  wire cea1c7;
  wire cea1c8;
  wire cea234;
  wire cea235;
  wire cea236;
  wire cea237;
  wire cea238;
  wire cea239;
  wire cea23a;
  wire cea23b;
  wire cea23c;
  wire cea246;
  wire cea247;
  wire cea248;
  wire cea249;
  wire cea24a;
  wire cea24b;
  wire cea24c;
  wire cea24d;
  wire cea24e;
  wire cea24f;
  wire cea250;
  wire cea251;
  wire cea252;
  wire cea253;
  wire cea254;
  wire cea255;
  wire cea256;
  wire cea257;
  wire cea258;
  wire cea259;
  wire cea25a;
  wire cea25b;
  wire cea265;
  wire cea266;
  wire cea267;
  wire cea268;
  wire cea269;
  wire cea26a;
  wire cea26b;
  wire cea26c;
  wire cea26d;
  wire cea26e;
  wire cea26f;
  wire cea270;
  wire cea271;
  wire cea272;
  wire cea273;
  wire cea274;
  wire cea275;
  wire cea276;
  wire cea277;
  wire cea278;
  wire cea279;
  wire cea27a;
  wire cea27b;
  wire cea280;
  wire cea283;
  wire cea286;
  wire cea287;
  wire cea288;
  wire cea289;
  wire cea28a;
  wire cea291;
  wire cea292;
  wire cea293;
  wire cea294;
  wire cea295;
  wire cea296;
  wire cea297;
  wire cea298;
  wire cea299;
  wire cea29a;
  wire cea29b;
  wire cea29c;
  wire cea29d;
  wire cea29e;
  wire cea29f;
  wire cea2a0;
  wire cea2a1;
  wire cea2a2;
  wire cea2a3;
  wire cea2a4;
  wire cea2a5;
  wire cea2a6;
  wire cea2a7;
  wire cea2a8;
  wire cea2ac;
  wire cea2ad;
  wire cea2ae;
  wire cea2af;
  wire cea2b0;
  wire cea2b1;
  wire cea2b2;
  wire cea2b3;
  wire cea2b4;
  wire cea2b5;
  wire cea2b6;
  wire cea2b7;
  wire cea2e2;
  wire cea2e3;
  wire cea2e4;
  wire cea2e5;
  wire cea2e6;
  wire cea2e7;
  wire cea2e8;
  wire cea2e9;
  wire cea2ea;
  wire cea2eb;
  wire cea2ec;
  wire cea2ed;
  wire cea2ee;
  wire cea2ef;
  wire cea2f0;
  wire cea2f1;
  wire cea2f2;
  wire cea2f3;
  wire cea2f4;
  wire cea2f5;
  wire cea2f6;
  wire cea2f7;
  wire cea2f8;
  wire cea2f9;
  wire cea31a;
  wire cea31b;
  wire cea31c;
  wire cea31d;
  wire cea31e;
  wire cea31f;
  wire cea320;
  wire cea321;
  wire cea322;
  wire cea323;
  wire cea324;
  wire cea325;
  wire cea326;
  wire cea327;
  wire cea328;
  wire cea329;
  wire cea32a;
  wire cea32b;
  wire cea32c;
  wire cea32d;
  wire cea32e;
  wire cea32f;
  wire cea330;
  wire cea331;
  wire cea332;
  wire cea333;
  wire cea334;
  wire cea335;
  wire cea336;
  wire cea337;
  wire cea338;
  wire cea339;
  wire cea33a;
  wire cea33b;
  wire cea33c;
  wire cea33d;
  wire cea33e;
  wire cea33f;
  wire cea340;
  wire cea341;
  wire cea342;
  wire cea343;
  wire cea344;
  wire cea345;
  wire cea346;
  wire cea347;
  wire cea348;
  wire cea354;
  wire cea355;
  wire cea356;
  wire cea357;
  wire cea358;
  wire cea359;
  wire cea35a;
  wire cea35b;
  wire cea35c;
  wire cea35d;
  wire cea35e;
  wire cea35f;
  wire cea360;
  wire cea361;
  wire cea362;
  wire cea363;
  wire cea364;
  wire cea365;
  wire cea366;
  wire cea367;
  wire cea368;
  wire cea369;
  wire cea36a;
  wire cea36b;
  wire cea36c;
  wire cea36d;
  wire cea36e;
  wire cea36f;
  wire cea370;
  wire cea371;
  wire cea372;
  wire cea373;
  wire cea374;
  wire cea375;
  wire cea376;
  wire cea377;
  wire cea378;
  wire cea379;
  wire cea37a;
  wire cea37b;
  wire cea37c;
  wire cea37d;
  wire cea37e;
  wire cea37f;
  wire cea380;
  wire cea381;
  wire cea382;
  wire cea383;
  wire cea384;
  wire cea385;
  wire cea386;
  wire cea387;
  wire cea388;
  wire cea389;
  wire cea38a;
  wire cea38b;
  wire cea38c;
  wire cea38d;
  wire cea38e;
  wire cea38f;
  wire cea390;
  wire cea391;
  wire cea392;
  wire cea393;
  wire cea394;
  wire cea395;
  wire cea396;
  wire cea397;
  wire cea398;
  wire cea399;
  wire cea39a;
  wire cea39b;
  wire cea39c;
  wire cea39d;
  wire cea39e;
  wire cea39f;
  wire cea3a0;
  wire cea3a1;
  wire cea3a2;
  wire cea3a3;
  wire cea3a4;
  wire cea3a5;
  wire cea3a6;
  wire cea3a7;
  wire cea3a8;
  wire cea3a9;
  wire cea3aa;
  wire cea3ab;
  wire cea3ac;
  wire cea3ad;
  wire cea3ae;
  wire cea3af;
  wire cea3b7;
  wire cea3b8;
  wire cea3b9;
  wire cea3ba;
  wire cea3bb;
  wire cea3bc;
  wire cea3bd;
  wire cea3be;
  wire cea3bf;
  wire cea3c0;
  wire cea3cb;
  wire cea3cc;
  wire cea3cd;
  wire cea3ce;
  wire cea3cf;
  wire cea3d0;
  wire cea3d8;
  wire cea3d9;
  wire cea3da;
  wire cea3db;
  wire cea3dc;
  wire cea3e8;
  wire cea3e9;
  wire cea3ea;
  wire cea3eb;
  wire cea3ec;
  wire cea3ed;
  wire cea3ee;
  wire cea3ef;
  wire cea3f0;
  wire cea3f1;
  wire cea3f2;
  wire cea3f3;
  wire cea3f7;
  wire cea3f8;
  wire cea3f9;
  wire cea3fa;
  wire cea3fb;
  wire cea3fc;
  wire cea404;
  wire cea405;
  wire cea406;
  wire cea407;
  wire cea408;
  wire cea409;
  wire cea40a;
  wire cea40b;
  wire cea40c;
  wire cea40d;
  wire cea40e;
  wire cea40f;
  wire cea410;
  wire cea411;
  wire cea412;
  wire cea413;
  wire cea414;
  wire cea415;
  wire cea416;
  wire cea417;
  wire cea418;
  wire cea419;
  wire cea41a;
  wire cea41b;
  wire cea41c;
  wire cea41d;
  wire cea41e;
  wire cea41f;
  wire cea420;
  wire cea421;
  wire cea422;
  wire cea423;
  wire cea424;
  wire cea425;
  wire cea426;
  wire cea427;
  wire cea428;
  wire cea42e;
  wire cea42f;
  wire cea430;
  wire cea431;
  wire cea432;
  wire cea433;
  wire cea434;
  wire cea435;
  wire cea436;
  wire cea437;
  wire cea438;
  wire cea439;
  wire cea43a;
  wire cea43b;
  wire cea43c;
  wire cea43d;
  wire cea43e;
  wire cea43f;
  wire cea440;
  wire cea441;
  wire cea442;
  wire cea443;
  wire cea444;
  wire cea445;
  wire cea446;
  wire cea447;
  wire cea448;
  wire cea449;
  wire cea44a;
  wire cea44b;
  wire cea44c;
  wire cea44d;
  wire cea44e;
  wire cea44f;
  wire cea450;
  wire cea451;
  wire cea452;
  wire cea453;
  wire cea454;
  wire cea455;
  wire cea456;
  wire cea457;
  wire cea458;
  wire cea459;
  wire cea45a;
  wire cea45b;
  wire cea45c;
  wire cea45d;
  wire cea45e;
  wire cea45f;
  wire cea460;
  wire cea461;
  wire cea462;
  wire cea463;
  wire cea464;
  wire cea465;
  wire cea466;
  wire cea467;
  wire cea468;
  wire cea469;
  wire cea46a;
  wire cea46b;
  wire cea46c;
  wire cea46d;
  wire cea46e;
  wire cea46f;
  wire cea470;
  wire cea471;
  wire cea472;
  wire cea473;
  wire cea474;
  wire cea475;
  wire cea476;
  wire cea477;
  wire cea478;
  wire cea479;
  wire cea47a;
  wire cea47b;
  wire cea47c;
  wire cea47d;
  wire cea47e;
  wire cea47f;
  wire cea480;
  wire cea481;
  wire cea482;
  wire cea483;
  wire cea484;
  wire cea485;
  wire cea486;
  wire cea487;
  wire cea488;
  wire cea489;
  wire cea48a;
  wire cea48b;
  wire cea48c;
  wire cea48d;
  wire cea48e;
  wire cea48f;
  wire cea490;
  wire cea491;
  wire cea492;
  wire cea493;
  wire cea494;
  wire cea499;
  wire cea49a;
  wire cea49b;
  wire cea49e;
  wire cea4a9;
  wire cea4aa;
  wire cea4ab;
  wire cea4ac;
  wire cea4ad;
  wire cea4ae;
  wire cea4af;
  wire ce9cb3;
  wire ce9cb4;
  wire ce9cb5;
  wire ce9cb6;
  wire ce9cb7;
  wire ce9cb8;
  wire ce9cb9;
  wire ce9cba;
  wire ce9cbb;
  wire ce9cbc;
  wire ce9cbd;
  wire ce9cbe;
  wire ce9cbf;
  wire ce9cc0;
  wire ce9cc1;
  wire ce9cc2;
  wire ce9cc3;
  wire ce9cc4;
  wire ce9cc5;
  wire ce9cc6;
  wire ce9cc7;
  wire ce9cc8;
  wire ce9cc9;
  wire ce9cca;
  wire ce9ccb;
  wire ce9ccc;
  wire ce9ccd;
  wire ce9cce;
  wire ce9ccf;
  wire ce9cd0;
  wire ce9cd1;
  wire ce9cd2;
  wire ce9cd3;
  wire ce9cd4;
  wire ce9cd7;
  wire ce9cd8;
  wire ce9cd9;
  wire ce9cda;
  wire ce9cdb;
  wire ce9cdc;
  wire ce9cdd;
  wire ce9cde;
  wire ce9cdf;
  wire ce9cf5;
  wire ce9cf6;
  wire ce9cf7;
  wire ce9cf8;
  wire ce9cf9;
  wire ce9cfa;
  wire ce9cfb;
  wire ce9cfc;
  wire ce9cfd;
  wire ce9d10;
  wire ce9d11;
  wire ce9d12;
  wire ce9d13;
  wire ce9d14;
  wire ce9d15;
  wire ce9d16;
  wire ce9d1f;
  wire ce9d20;
  wire ce9d21;
  wire ce9d22;
  wire ce9d26;
  wire ce9d27;
  wire ce9d28;
  wire ce9d29;
  wire ce9d2c;
  wire ce9d2d;
  wire ce9d2e;
  wire ce9d2f;
  wire ce9d30;
  wire ce9d31;
  wire ce9d32;
  wire ce9d33;
  wire ce9d34;
  wire ce9d35;
  wire ce9d36;
  wire ce9d37;
  wire ce9d3d;
  wire ce9d3e;
  wire ce9d3f;
  wire ce9d40;
  wire ce9d41;
  wire ce9d42;
  wire ce9d43;
  wire ce9d45;
  wire ce9d46;
  wire ce9d47;
  wire ce9d48;
  wire ce9d49;
  wire ce9d4a;
  wire ce9d4b;
  wire ce9d4d;
  wire ce9d4e;
  wire ce9d4f;
  wire ce9d50;
  wire ce9d51;
  wire ce9d52;
  wire ce9d53;
  wire ce9d54;
  wire ce9d55;
  wire ce9d56;
  wire ce9d57;
  wire ce9d58;
  wire ce9d59;
  wire ce9d5a;
  wire ce9d5b;
  wire ce9d6e;
  wire ce9d6f;
  wire ce9d70;
  wire ce9d71;
  wire ce9d72;
  wire ce9d79;
  wire ce9da5;
  wire ce9da6;
  wire ce9daf;
  wire ce9db0;
  wire ce9db5;
  wire ce9db6;
  wire ce9db7;
  wire ce9db8;
  wire ce9db9;
  wire ce9dba;
  wire ce9dbb;
  wire ce9dc6;
  wire ce9dc7;
  wire ce9dc8;
  wire ce9dd3;
  wire ce9dd4;
  wire ce9dda;
  wire ce9ddb;
  wire ce9ddc;
  wire ce9ddd;
  wire ce9def;
  wire ce9df0;
  wire ce9df1;
  wire ce9dfc;
  wire ce9dfd;
  wire ce9dfe;
  wire ce9e09;
  wire ce9e0a;
  wire ce9e0b;
  wire ce9e0c;
  wire ce9e1f;
  wire ce9e20;
  wire ce9e21;
  wire ce9e22;
  wire ce9e23;
  wire ce9e24;
  wire ce9e25;
  wire ce9e26;
  wire ce9e27;
  wire ce9e28;
  wire ce9e29;
  wire ce9e5e;
  wire ce9e5f;
  wire ce9e60;
  wire c3bbba;
  wire c3bbbb;
  wire c3bbbc;
  wire c3bbbd;
  wire c3bbbe;
  wire c3bbbf;
  wire c3bbc0;
  wire c3bbc1;
  wire c3bbd1;
  wire c3bbd2;
  wire c3bbd3;
  wire c3bbd4;
  wire c3bbd5;
  wire c3bbd6;
  wire c3bbe2;
  wire c3bbe8;
  wire c3bbea;
  wire c3bbef;
  wire c3bbf0;
  wire c3bbf1;
  wire c3bbf2;
  wire c3bbf3;
  wire c3bbf4;
  wire c3bbf5;
  wire c3bbf6;
  wire c3bbf7;
  wire c3bbf8;
  wire c3bbf9;
  wire c3bbfa;
  wire c3bbfb;
  wire c3bbfc;
  wire c3bbfd;
  wire c3bbfe;
  wire c3bc02;
  wire c3bc03;
  wire c3bc04;
  wire c3bc05;
  wire c3bc06;
  wire c3bc07;
  wire c3bc08;
  wire c3bc09;
  wire c3bc0a;
  wire c3bc0b;
  wire c3bc0c;
  wire c3bc0d;
  wire c3bc0e;
  wire c3bc0f;
  wire c3bc10;
  wire c3bc15;
  wire c3bc16;
  wire c3bc17;
  wire c3bc18;
  wire c3bc20;
  wire c3bc21;
  wire c3bc22;
  wire c3bc28;
  wire c3bc29;
  wire c3bc2a;
  wire c3bc2b;
  wire c3bc2c;
  wire c3bc2d;
  wire c3bc2e;
  wire c3bc2f;
  wire c3bc33;
  wire c3bc34;
  wire c3bc35;
  wire c3bc36;
  wire c3bc37;
  wire c3bc38;
  wire c3bc39;
  wire c3bc3a;
  wire c3bc3b;
  wire c3bc3c;
  wire c3bc41;
  wire c3bc42;
  wire c3bc43;
  wire c3bc44;
  wire c3bc45;
  wire c3bc46;
  wire c3bc47;
  wire c3bc48;
  wire c3bc49;
  wire c3bc4a;
  wire c3bc4b;
  wire c3bc4c;
  wire c3bc4d;
  wire c3bc4e;
  wire c3bc4f;
  wire c3bc50;
  wire c3bc51;
  wire c3bc52;
  wire c3bc53;
  wire c3bc54;
  wire c3bc55;
  wire c3bc56;
  wire c3bc57;
  wire c3bc58;
  wire c3bc59;
  wire c3bc5a;
  wire c3bc5b;
  wire c3bc5c;
  wire c3bc5d;
  wire c3bc5e;
  wire c3bc5f;
  wire c3bc60;
  wire c3bc61;
  wire c3bc62;
  wire c3bc63;
  wire c3bc64;
  wire c3bc65;
  wire c3bc66;
  wire c3bc67;
  wire c3bc68;
  wire c3bc69;
  wire c3bc6a;
  wire c3bc6b;
  wire c3bc6c;
  wire c3bc6d;
  wire c3bc6e;
  wire c3bc6f;
  wire c3bc70;
  wire c3bc71;
  wire c3bc72;
  wire c3bc73;
  wire c3bc74;
  wire c3bc75;
  wire c3bc76;
  wire c3bc77;
  wire c3bc78;
  wire c3bc79;
  wire c3bc7a;
  wire c3bc7b;
  wire c3bc7c;
  wire c3bc7d;
  wire c3bc7e;
  wire c3bc7f;
  wire c3bc80;
  wire c3bc81;
  wire c3bc82;
  wire c3bc83;
  wire c3bc84;
  wire c3bc85;
  wire c3bc86;
  wire c3bc87;
  wire c3bc88;
  wire c3bc89;
  wire c3bc8a;
  wire c3bc8b;
  wire c3bc8c;
  wire c3bc8d;
  wire c3bc8e;
  wire c3bc8f;
  wire c3bc90;
  wire c3bc91;
  wire c3bc92;
  wire c3bc93;
  wire c3bc94;
  wire c3bc95;
  wire c3bc96;
  wire c3bc97;
  wire c3bc98;
  wire c3bc99;
  wire c3bc9a;
  wire c3bc9b;
  wire c3bc9c;
  wire c3bc9d;
  wire c3bc9e;
  wire c3bc9f;
  wire c3bca0;
  wire c3bca1;
  wire c3bca2;
  wire c3bca3;
  wire c3bca4;
  wire c3bca5;
  wire c3bca6;
  wire c3bca7;
  wire c3bca8;
  wire c3bca9;
  wire c3bcaa;
  wire c3bcab;
  wire c3bcac;
  wire c3bcad;
  wire c3bcae;
  wire c3bcaf;
  wire c3bcb0;
  wire c3bcb1;
  wire c3bcb2;
  wire v84564c;
  wire c3bcb3;
  wire c3bcb4;
  wire c3bcb5;
  wire c3bcb6;
  wire c3bcb7;
  wire c3bcbc;
  wire c3bcbd;
  wire c3bcbe;
  wire c3bcbf;
  wire c3bcc0;
  wire c3bcc1;
  wire c3bcc2;
  wire c3bcc3;
  wire c3bcc4;
  wire c3bcc5;
  wire c3bcc6;
  wire c3bcc7;
  wire c3bcc8;
  wire c3bcc9;
  wire c3bcca;
  wire c3bccb;
  wire c3bccc;
  wire c3bccd;
  wire c3bcce;
  wire c3bccf;
  wire c3bcd0;
  wire c3bcd1;
  wire c3bcd2;
  wire c3bcd3;
  wire c3bcd4;
  wire c3bcd5;
  wire c3bcd6;
  wire c3bcd7;
  wire c3bcd8;
  wire c3bcd9;
  wire c3bcda;
  wire c3bcdb;
  wire c3bcdc;
  wire c3bcdd;
  wire c3bcde;
  wire c3bcdf;
  wire c3bce0;
  wire c3bce1;
  wire c3bce2;
  wire c3bce3;
  wire c3bce4;
  wire c3bce5;
  wire c3bce6;
  wire c3bce7;
  wire c3bce8;
  wire c3bce9;
  wire c3bcea;
  wire c3bceb;
  wire c3bcec;
  wire c3bced;
  wire c3bcee;
  wire c3bcef;
  wire c3bcf0;
  wire c3bcf1;
  wire c3bcf2;
  wire c3bcf3;
  wire c3bcf4;
  wire c3bcf5;
  wire c3bcf6;
  wire c3bcf7;
  wire c3bcf8;
  wire c3bcf9;
  wire c3bcfa;
  wire c3bcfb;
  wire c3bcfc;
  wire c3bcfd;
  wire c3bcfe;
  wire c3bcff;
  wire c3bd00;
  wire c3bd01;
  wire c3bd02;
  wire c3bd03;
  wire c3bd04;
  wire c3bd05;
  wire c3bd06;
  wire c3bd07;
  wire c3bd08;
  wire c3bd09;
  wire c3bd0f;
  wire c3bd10;
  wire c3bd11;
  wire c3bd12;
  wire c3bd13;
  wire c3bd14;
  wire c3bd15;
  wire c3bd16;
  wire c3bd17;
  wire c3bd21;
  wire c3bd22;
  wire c3bd24;
  wire c3bd25;
  wire c3bd2c;
  wire c3bd2d;
  wire c3bd35;
  wire c3bd36;
  wire c3bd37;
  wire c3bd38;
  wire c3bd39;
  wire c3bd3a;
  wire c3bd3b;
  wire c3bd3c;
  wire c3bd3d;
  wire c3bd3e;
  wire c3bd3f;
  wire c3bd41;
  wire c3bd42;
  wire c3bd43;
  wire c3bd44;
  wire c3bd45;
  wire c3bd46;
  wire c3bd47;
  wire c3bd4b;
  wire c3bd4c;
  wire c3bd4d;
  wire c3bd4e;
  wire c3bd4f;
  wire c3bd50;
  wire c3bd51;
  wire c3bd5b;
  wire c3bd5c;
  wire c3bd5d;
  wire c3bd5e;
  wire c3bd5f;
  wire c3bd60;
  wire c3bd61;
  wire c3bd62;
  wire c3bd63;
  wire c3bd64;
  wire c3bd65;
  wire c3bd66;
  wire c3bd67;
  wire c3bd68;
  wire c3bd69;
  wire c3bd6a;
  wire c3bd6b;
  wire c3bd6c;
  wire c3bd6d;
  wire c3bd71;
  wire c3bd72;
  wire c3bd73;
  wire c3bd77;
  wire c3bd78;
  wire c3bd79;
  wire c3bd7a;
  wire c3bd7b;
  wire c3bd7c;
  wire c3bd7d;
  wire c3bd7e;
  wire c3bd7f;
  wire c3bd80;
  wire c3bd81;
  wire c3bd82;
  wire c3bd83;
  wire c3bd84;
  wire c3bd85;
  wire c3bd86;
  wire c3bd87;
  wire c3bd88;
  wire c3bd89;
  wire c3bd8a;
  wire c3bd8b;
  wire c3bd8c;
  wire c3bd8d;
  wire c3bd8e;
  wire c3bd8f;
  wire c3bd90;
  wire c3bd91;
  wire c3bd92;
  wire c3bd93;
  wire c3bd94;
  wire c3bd95;
  wire c3bd96;
  wire c3bd97;
  wire c3bd98;
  wire c3bd99;
  wire c3bd9a;
  wire c3bd9b;
  wire c3bd9c;
  wire c3bd9d;
  wire c3bd9e;
  wire c3bd9f;
  wire c3bda0;
  wire c3bda1;
  wire c3bda2;
  wire c3bda3;
  wire c3bda4;
  wire c3bda5;
  wire c3bda6;
  wire c3bda7;
  wire c3bda8;
  wire c3bda9;
  wire c3bdaa;
  wire c3bdab;
  wire c3bdac;
  wire c3bdad;
  wire c3bdae;
  wire c3bdaf;
  wire c3bdb0;
  wire c3bdb1;
  wire c3bdb2;
  wire c3bdb3;
  wire c3bdb4;
  wire c3bdb5;
  wire c3bdb6;
  wire c3bdb7;
  wire c3bdb8;
  wire c3bdb9;
  wire c3bdba;
  wire c3bdbb;
  wire c3bdbc;
  wire c3bdbd;
  wire c3bdbe;
  wire c3bdbf;
  wire c3bdc0;
  wire c3bdc1;
  wire c3bdc2;
  wire c3bdc3;
  wire c3bdc4;
  wire c3bdc5;
  wire c3bdc6;
  wire c3bdc7;
  wire c3bdc8;
  wire c3bdc9;
  wire c3bdca;
  wire c3bdcb;
  wire c3bdcc;
  wire c3bdcd;
  wire c3bdce;
  wire c3bdcf;
  wire c3bdd0;
  wire c3bdd1;
  wire c3bdd2;
  wire c3bdd3;
  wire c3bdd4;
  wire c3bdd5;
  wire c3bdd6;
  wire c3bdd7;
  wire c3bdd8;
  wire c3bdd9;
  wire c3bdda;
  wire c3bddb;
  wire c3bddc;
  wire c3bddd;
  wire c3bdde;
  wire c3bddf;
  wire c3bde0;
  wire c3bde1;
  wire c3bde2;
  wire c3bde3;
  wire c3bde4;
  wire c3bde5;
  wire c3bde6;
  wire c3bde7;
  wire c3bde8;
  wire c3bde9;
  wire c3bdea;
  wire c3bdf4;
  wire c3bdf5;
  wire c3bdf6;
  wire c3bdf7;
  wire c3bdf8;
  wire c3bdf9;
  wire c3bdfa;
  wire c3bdfb;
  wire c3bdfc;
  wire c3bdfd;
  wire c3bdfe;
  wire c3bdff;
  wire c3be00;
  wire c3be01;
  wire c3be02;
  wire c3be03;
  wire c3be04;
  wire c3be05;
  wire c3be06;
  wire c3b60a;
  wire c3b60b;
  wire c3b613;
  wire c3b614;
  wire c3b615;
  wire c3b616;
  wire c3b617;
  wire c3b618;
  wire c3b619;
  wire c3b61a;
  wire c3b61b;
  wire c3b61c;
  wire c3b61d;
  wire c3b61e;
  wire c3b61f;
  wire c3b620;
  wire c3b621;
  wire c3b622;
  wire c3b623;
  wire c3b624;
  wire c3b625;
  wire c3b626;
  wire c3b627;
  wire c3b628;
  wire c3b629;
  wire c3b62a;
  wire c3b62b;
  wire c3b62c;
  wire c3b62d;
  wire c3b62e;
  wire c3b62f;
  wire c3b630;
  wire c3b631;
  wire c3b632;
  wire c3b633;
  wire c3b634;
  wire c3b635;
  wire c3b636;
  wire c3b637;
  wire c3b638;
  wire c3b639;
  wire c3b63a;
  wire c3b63b;
  wire c3b63c;
  wire c3b63d;
  wire c3b63e;
  wire c3b63f;
  wire c3b640;
  wire c3b641;
  wire c3b642;
  wire c3b643;
  wire c3b644;
  wire c3b645;
  wire c3b646;
  wire c3b647;
  wire c3b648;
  wire c3b649;
  wire c3b64a;
  wire c3b64b;
  wire c3b64c;
  wire c3b64d;
  wire c3b64e;
  wire c3b650;
  wire c3b651;
  wire c3b652;
  wire c3b653;
  wire c3b654;
  wire c3b655;
  wire c3b656;
  wire c3b657;
  wire c3b658;
  wire c3b659;
  wire c3b65a;
  wire c3b65b;
  wire c3b660;
  wire c3b661;
  wire c3b662;
  wire c3b663;
  wire c3b664;
  wire c3b665;
  wire c3b66a;
  wire c3b66b;
  wire c3b66c;
  wire c3b66e;
  wire c3b66f;
  wire c3b674;
  wire c3b675;
  wire c3b676;
  wire c3b677;
  wire c3b678;
  wire c3b679;
  wire c3b67a;
  wire c3b67b;
  wire c3b67c;
  wire c3b683;
  wire c3b684;
  wire c3b685;
  wire c3b686;
  wire c3b687;
  wire c3b689;
  wire c3b68a;
  wire c3b68b;
  wire c3b68c;
  wire c3b68d;
  wire c3b68e;
  wire c3b68f;
  wire c3b690;
  wire c3b691;
  wire c3b692;
  wire c3b693;
  wire c3b694;
  wire c3b696;
  wire c3b697;
  wire c3b698;
  wire c3b699;
  wire c3b6a0;
  wire c3b6a1;
  wire c3b6a3;
  wire c3b6a4;
  wire c3b6a5;
  wire c3b6a6;
  wire c3b6a7;
  wire c3b6a8;
  wire c3b6a9;
  wire c3b6aa;
  wire c3b6ab;
  wire c3b6ac;
  wire c3b6ad;
  wire c3b6ae;
  wire c3b6af;
  wire c3b6b0;
  wire c3b6b1;
  wire c3b6b2;
  wire c3b6b3;
  wire c3b6b4;
  wire c3b6b5;
  wire c3b6b6;
  wire c3b6b7;
  wire c3b6b8;
  wire c3b6b9;
  wire c3b6bc;
  wire c3b6bd;
  wire c3b6be;
  wire c3b6bf;
  wire c3b6c0;
  wire c3b6c1;
  wire c3b6c2;
  wire c3b6c3;
  wire c3b6c4;
  wire c3b6c5;
  wire c3b6c6;
  wire c3b6c7;
  wire c3b6c8;
  wire c3b6c9;
  wire c3b6ca;
  wire c3b6cb;
  wire c3b6cc;
  wire c3b6cd;
  wire c3b6ce;
  wire c3b6cf;
  wire c3b6d0;
  wire c3b6d1;
  wire c3b6d2;
  wire c3b6d3;
  wire c3b6d4;
  wire c3b6d5;
  wire c3b6d6;
  wire c3b6d7;
  wire c3b6d8;
  wire c3b6d9;
  wire c3b6da;
  wire c3b6db;
  wire c3b6dc;
  wire c3b6dd;
  wire c3b6de;
  wire c3b6df;
  wire c3b6e0;
  wire c3b6e1;
  wire c3b6e2;
  wire c3b6e3;
  wire c3b6e4;
  wire c3b6e5;
  wire c3b6e6;
  wire c3b6e7;
  wire c3b6e8;
  wire c3b6e9;
  wire c3b6ea;
  wire c3b6eb;
  wire c3b6ec;
  wire c3b6ed;
  wire c3b6ee;
  wire c3b6ef;
  wire c3b6f0;
  wire c3b6f1;
  wire c3b6f2;
  wire c3b6f3;
  wire c3b6f4;
  wire c3b6f5;
  wire c3b6f6;
  wire c3b6f7;
  wire c3b6f8;
  wire c3b6f9;
  wire c3b6fa;
  wire c3b6fb;
  wire c3b6fc;
  wire c3b6fd;
  wire c3b6fe;
  wire c3b6ff;
  wire c3b700;
  wire c3b701;
  wire c3b702;
  wire c3b703;
  wire c3b704;
  wire c3b705;
  wire c3b706;
  wire c3b707;
  wire c3b708;
  wire c3b709;
  wire c3b70a;
  wire c3b70b;
  wire c3b70c;
  wire c3b70d;
  wire c3b70e;
  wire c3b70f;
  wire c3b710;
  wire c3b711;
  wire c3b712;
  wire c3b713;
  wire c3b714;
  wire c3b715;
  wire c3b716;
  wire c3b717;
  wire c3b718;
  wire c3b719;
  wire c3b71a;
  wire c3b71b;
  wire c3b71c;
  wire c3b71d;
  wire c3b71e;
  wire c3b71f;
  wire c3b720;
  wire c3b721;
  wire c3b722;
  wire c3b723;
  wire c3b724;
  wire c3b725;
  wire c3b726;
  wire c3b727;
  wire c3b728;
  wire c3b729;
  wire c3b72a;
  wire c3b72b;
  wire c3b72c;
  wire c3b72d;
  wire c3b72f;
  wire c3b730;
  wire c3b731;
  wire c3b732;
  wire c3b733;
  wire c3b734;
  wire c3b735;
  wire c3b736;
  wire c3b737;
  wire c3b738;
  wire c3b739;
  wire c3b73a;
  wire c3b73b;
  wire c3b73c;
  wire c3b73d;
  wire c3b73e;
  wire c3b749;
  wire c3b74a;
  wire c3b74b;
  wire c3b74c;
  wire c3b74d;
  wire c3b74e;
  wire c3b74f;
  wire c3b750;
  wire c3b751;
  wire c3b752;
  wire c3b753;
  wire c3b754;
  wire c3b755;
  wire c3b756;
  wire c3b757;
  wire c3b768;
  wire c3b769;
  wire c3b76b;
  wire c3b76c;
  wire c3b76d;
  wire c3b76e;
  wire c3b76f;
  wire c3b770;
  wire c3b771;
  wire c3b772;
  wire c3b773;
  wire c3b774;
  wire c3b775;
  wire c3b776;
  wire c3b777;
  wire c3b778;
  wire c3b779;
  wire c3b77a;
  wire c3b77b;
  wire c3b77c;
  wire c3b77d;
  wire c3b77e;
  wire c3b77f;
  wire c3b780;
  wire c3b797;
  wire c3b798;
  wire c3b799;
  wire c3b79a;
  wire c3b79b;
  wire c3b79c;
  wire c3b79d;
  wire c3b79e;
  wire c3b79f;
  wire c3b7a0;
  wire c3b7a1;
  wire c3b7a2;
  wire c3b7a3;
  wire c3b7a4;
  wire c3b7a5;
  wire c3b7a6;
  wire c3b7a7;
  wire c3b7a8;
  wire c3b7a9;
  wire c3b7aa;
  wire c3b7ab;
  wire c3b7ac;
  wire c3b7ad;
  wire c3b7ae;
  wire c3b7af;
  wire c3b7b0;
  wire c3b7b1;
  wire c3b7b2;
  wire c3b7b3;
  wire c3b7b4;
  wire c3b7b5;
  wire c3b7b6;
  wire c3b7b7;
  wire c3b7bd;
  wire c3b7c1;
  wire c3b7c2;
  wire c3b7c3;
  wire c3b7cc;
  wire c3b7d0;
  wire c3b7d1;
  wire c3b7d2;
  wire c3b7d3;
  wire c3b7d4;
  wire c3b7d5;
  wire c3b7d6;
  wire c3b7d7;
  wire c3b7db;
  wire c3b7dc;
  wire c3b7dd;
  wire c3b7de;
  wire c3b7df;
  wire c3b7e0;
  wire c3b7e1;
  wire c3b7e4;
  wire c3b7e5;
  wire c3b7e6;
  wire c3b7e7;
  wire c3b7e8;
  wire c3b7e9;
  wire c3b7ea;
  wire c3b7eb;
  wire c3b7ec;
  wire c3b7ed;
  wire c3b7ee;
  wire c3b7ef;
  wire c3b7f0;
  wire c3b7f4;
  wire c3b7f5;
  wire c3b7f6;
  wire c3b7f7;
  wire c3b7f8;
  wire c3b7f9;
  wire c3b7fa;
  wire c3b7fb;
  wire c3b7fc;
  wire c3b7fd;
  wire c3b7fe;
  wire c3b7ff;
  wire c3b800;
  wire c3b801;
  wire c3b802;
  wire c3b803;
  wire c3b804;
  wire c3b805;
  wire c3b806;
  wire c3b807;
  wire c3b808;
  wire c3b809;
  wire c3b80a;
  wire c3b80b;
  wire c3b80c;
  wire c3b80d;
  wire c3b80e;
  wire c3b80f;
  wire c3b810;
  wire c3b811;
  wire c3b812;
  wire c3b813;
  wire c3b814;
  wire c3b815;
  wire c3b816;
  wire c3b817;
  wire c3b818;
  wire c3b819;
  wire c3b81a;
  wire c3b81b;
  wire c3b81c;
  wire c3b81d;
  wire c3b81e;
  wire c3b81f;
  wire c3b820;
  wire c3b821;
  wire c3b822;
  wire c3b823;
  wire c3b824;
  wire c3b825;
  wire c3b826;
  wire c3b827;
  wire c3b828;
  wire c3b829;
  wire c3b82a;
  wire c3b82b;
  wire c3b82c;
  wire c3b82d;
  wire c3b82e;
  wire c3b82f;
  wire c3b830;
  wire c3b844;
  wire c3b845;
  wire c3b846;
  wire c3b849;
  wire c3b84a;
  wire c3b84b;
  wire c3b84c;
  wire c3b84d;
  wire c3b84e;
  wire c3b84f;
  wire c3b850;
  wire c3b851;
  wire c3b852;
  wire c3b85b;
  wire c3b870;
  wire c3b871;
  wire c3b872;
  wire c3b873;
  wire c3b874;
  wire c3b875;
  wire c3b876;
  wire c3b877;
  wire c3b878;
  wire c3b883;
  wire c3b884;
  wire c3b885;
  wire c3b886;
  wire c3b887;
  wire c3b888;
  wire c3b889;
  wire c3b88b;
  wire c3b88c;
  wire c3b88d;
  wire c3b88e;
  wire c3b88f;
  wire c3b890;
  wire c3b891;
  wire c3b892;
  wire c3b893;
  wire c3b894;
  wire c3b895;
  wire c3b896;
  wire c3b8ab;
  wire c3b8ac;
  wire c3b8ae;
  wire c3b8af;
  wire c3b8b0;
  wire c3b8b1;
  wire c3b8b2;
  wire c3b8b3;
  wire c3b8b4;
  wire c3b8b5;
  wire c3b8b6;
  wire c3b8b7;
  wire c3b8b8;
  wire c3b8ca;
  wire c3b8cb;
  wire c3b8cc;
  wire bdb580;
  wire bdb581;
  wire bdb582;
  wire bdb583;
  wire bdb584;
  wire bdb585;
  wire bdb586;
  wire bdb587;
  wire bdb588;
  wire bdb589;
  wire bdb58a;
  wire bdb58b;
  wire bdb58c;
  wire bdb58d;
  wire bdb595;
  wire bdb596;
  wire bdb597;
  wire bdb598;
  wire bdb599;
  wire bdb59a;
  wire bdb59b;
  wire bdb59c;
  wire bdb59d;
  wire bdb59e;
  wire bdb59f;
  wire bdb5a0;
  wire bdb5a1;
  wire bdb5a2;
  wire bdb5a3;
  wire bdb5a4;
  wire bdb5a5;
  wire bdb5a6;
  wire bdb5a7;
  wire bdb5a8;
  wire bdb5a9;
  wire bdb5aa;
  wire bdb5ab;
  wire bdb5ac;
  wire bdb5ad;
  wire bdb5ae;
  wire bdb5af;
  wire bdb5b0;
  wire bdb5b1;
  wire bdb5b2;
  wire bdb5b3;
  wire bdb5b4;
  wire bdb5b5;
  wire bdb5b6;
  wire bdb5b7;
  wire bdb5b8;
  wire bdb5b9;
  wire bdb5ba;
  wire v84564f;
  wire v845647;
  wire b840ac;
  wire v84564b;
  wire v845643;
  wire b840ad;
  wire b840ae;
  wire b840af;
  wire b840b0;
  wire b840b1;
  wire b840b2;
  wire b840b3;
  wire b29c3b;
  wire b29c3c;
  wire b29c3d;
  wire b29cb9;
  wire b29cba;
  wire b29cbb;
  wire b29cbc;
  wire b29cbd;
  wire b29cbe;
  wire b29cbf;
  wire b29cc0;
  wire b29cc1;
  wire b29cc8;
  wire b29cc9;
  wire b29cca;
  wire b29ccb;
  wire b29cd4;
  wire b29cd5;
  wire b29cd6;
  wire b29cd7;
  wire b29cd8;
  wire b29cd9;
  wire b29cda;
  wire b29cdb;
  wire b29cdd;
  wire b29cdf;
  wire b29ce0;
  wire b29ce4;
  wire b29ce5;
  wire b29ce6;
  wire b29ce7;
  wire b29ce8;
  wire b29ce9;
  wire b29cea;
  wire b29ceb;
  wire b29cec;
  wire b29cf0;
  wire b29cf2;
  wire b29cf3;
  wire b29cf6;
  wire b29cf7;
  wire b29cf8;
  wire b29cfb;
  wire b29cfc;
  wire b29cfd;
  wire b29cfe;
  wire b29cff;
  wire b29d00;
  wire b29d01;
  wire b29d02;
  wire b29d03;
  wire b29d04;
  wire b29d05;
  wire b29d06;
  wire b29d07;
  wire b29d0d;
  wire b29d0e;
  wire b29d0f;
  wire b29d17;
  wire b29d1e;
  wire b29d1f;
  wire b29d20;
  wire b29d21;
  wire b29d22;
  wire b29d23;
  wire b29d24;
  wire b29d25;
  wire b29d29;
  wire b29d2a;
  wire b29d2b;
  wire b29d2c;
  wire b29d2e;
  wire b29d2f;
  wire b29d30;
  wire b29d33;
  wire b29d34;
  wire b29d35;
  wire b29d36;
  wire b29d37;
  wire b29d38;
  wire b29d39;
  wire b29d3a;
  wire b29d3b;
  wire b29d3c;
  wire b29d3d;
  wire b29d3e;
  wire b29d49;
  wire b29d4a;
  wire b29d4b;
  wire b29d4c;
  wire b29d4d;
  wire b29d4e;
  wire b29d4f;
  wire b29d50;
  wire b29d51;
  wire b29d52;
  wire b29d53;
  wire b29d54;
  wire b29d55;
  wire b29d56;
  wire b29d57;
  wire b29d58;
  wire b29d59;
  wire b29d5a;
  wire b29d5b;
  wire b29d5c;
  wire b29d5d;
  wire b29d5e;
  wire b29d5f;
  wire b29d60;
  wire b29d61;
  wire b29d62;
  wire b29d63;
  wire b29d64;
  wire b29d65;
  wire b29d66;
  wire b29d67;
  wire b29d68;
  wire b29d69;
  wire b29d6a;
  wire b29d6b;
  wire b29d6c;
  wire b29d6d;
  wire b29d6e;
  wire b29d6f;
  wire b29d70;
  wire b29d71;
  wire b29d72;
  wire b29d73;
  wire b29d74;
  wire b29d75;
  wire b29d76;
  wire b29d77;
  wire b29d78;
  wire b29d79;
  wire b29d7a;
  wire b29d7b;
  wire b29d7c;
  wire b29d7d;
  wire b29d7e;
  wire b29d7f;
  wire b29d80;
  wire b29d81;
  wire b29d82;
  wire b29d83;
  wire b29d84;
  wire b29d85;
  wire b29d86;
  wire b29d87;
  wire b29d88;
  wire b29d89;
  wire b29d8a;
  wire b29d8b;
  wire b29d8c;
  wire b29d8d;
  wire b29d8e;
  wire b29d8f;
  wire b29d90;
  wire b29d91;
  wire b29d92;
  wire b29d93;
  wire b29d94;
  wire b29d95;
  wire b29d96;
  wire b29d97;
  wire b29d98;
  wire b29d99;
  wire b29d9a;
  wire b29d9b;
  wire b29d9c;
  wire b29d9d;
  wire b29e47;
  wire b29e48;
  wire b29e49;
  wire b29e4a;
  wire b29e4b;
  wire b29e4c;
  wire b29e4d;
  wire b29e4e;
  wire b29e4f;
  wire b29e50;
  wire b29e51;
  wire b29e52;
  wire b29e53;
  wire b29e54;
  wire b29e55;
  wire b29e56;
  wire b29e57;
  wire b29e58;
  wire b29e59;
  wire b29e5a;
  wire b29e5b;
  wire b29e5c;
  wire b29e5d;
  wire b29e5e;
  wire b29e5f;
  wire b29e60;
  wire b29e61;
  wire b29e65;
  wire b29e66;
  wire b29e67;
  wire b29e68;
  wire b29e69;
  wire b29e6a;
  wire b29e6b;
  wire b29e6c;
  wire b29e6d;
  wire b29e6e;
  wire b29e6f;
  wire b29e70;
  wire b29e71;
  wire b29e72;
  wire b29e95;
  wire b29e96;
  wire b29e97;
  wire b29e98;
  wire b29e99;
  wire b29e9a;
  wire b29e9b;
  wire b29e9c;
  wire b29e9d;
  wire b29e9e;
  wire b29e9f;
  wire b29ea0;
  wire b29ea1;
  wire b29ea2;
  wire b29ea3;
  wire b29ea4;
  wire b29ea5;
  wire b29ea6;
  wire b29ea7;
  wire b29ea8;
  wire b29ea9;
  wire b29eaa;
  wire b29eab;
  wire b29eac;
  wire b29ead;
  wire b29eae;
  wire b29eaf;
  wire b29eb0;
  wire b29eb1;
  wire b29eb2;
  wire b29eb3;
  wire b29eb4;
  wire b29eb5;
  wire b29eb6;
  wire b29eb7;
  wire b29eb8;
  wire b29eb9;
  wire b29eba;
  wire b29ebb;
  wire b29ebc;
  wire b29ebd;
  wire b29ebe;
  wire b29ebf;
  wire b29ec0;
  wire b29ec1;
  wire b29ec2;
  wire b29ec3;
  wire b29ec4;
  wire b29ec5;
  wire b29ec6;
  wire b29ec7;
  wire b29ec8;
  wire b29ec9;
  wire b29eca;
  wire b29ecb;
  wire b29ecc;
  wire b29ecd;
  wire b29ece;
  wire b29ecf;
  wire b29ed0;
  wire b29ed1;
  wire b29ed2;
  wire b29ed3;
  wire b29ed4;
  wire b29ed5;
  wire b29ed6;
  wire b29ed7;
  wire b29ed8;
  wire b29ed9;
  wire b29eda;
  wire b29edb;
  wire b29edc;
  wire b29edd;
  wire b29ede;
  wire b29edf;
  wire b29ee0;
  wire b29ee1;
  wire b29ee5;
  wire b29ee6;
  wire b29ee7;
  wire b29ee8;
  wire b29ee9;
  wire b29eea;
  wire b29eeb;
  wire b29eec;
  wire b29eed;
  wire b29eee;
  wire b29ef5;
  wire b29efa;
  wire b29efb;
  wire b29efc;
  wire b29efd;
  wire b29efe;
  wire b29f03;
  wire b29f04;
  wire b29f05;
  wire b29f06;
  wire b29f07;
  wire b29f08;
  wire b29f09;
  wire b29f0a;
  wire b29f0b;
  wire b29f0c;
  wire b29f0d;
  wire b29f0e;
  wire b29f0f;
  wire b29f10;
  wire b29f17;
  wire b29f18;
  wire b29f19;
  wire b29f1a;
  wire b29f1b;
  wire b29f1c;
  wire b29f1d;
  wire b29f1e;
  wire b29f1f;
  wire b29f31;
  wire b29f32;
  wire b29f33;
  wire b29f34;
  wire b29f35;
  wire b29f36;
  wire b29f37;
  wire b29f38;
  wire b29f39;
  wire b29f3c;
  wire b29f3d;
  wire b29f3e;
  wire b29f40;
  wire b29f41;
  wire b29f42;
  wire b29f43;
  wire b29f44;
  wire b29f45;
  wire b29f46;
  wire b29f47;
  wire b29f4f;
  wire b29f50;
  wire b29f51;
  wire b29f52;
  wire b29f53;
  wire b29f54;
  wire b29f55;
  wire b29f56;
  wire b29f57;
  wire b29f58;
  wire b29f59;
  wire b29f5a;
  wire b29f5b;
  wire b29f5c;
  wire b29f5d;
  wire b29f5e;
  wire b29f5f;
  wire b29f60;
  wire b29f61;
  wire b29f62;
  wire b29f63;
  wire b29f64;
  wire b29f65;
  wire b29f66;
  wire b29f67;
  wire b29f68;
  wire b29f69;
  wire b29f6a;
  wire b29f6b;
  wire b29f6c;
  wire b29f6d;
  wire b29f74;
  wire b29f75;
  wire b29f76;
  wire b29f77;
  wire b29f78;
  wire b29f79;
  wire b29f7a;
  wire b29f7b;
  wire b29f7c;
  wire b29f7d;
  wire b29f7e;
  wire b29f7f;
  wire b29f80;
  wire b29f81;
  wire b29f82;
  wire b29f83;
  wire b29f84;
  wire b29f85;
  wire b29f86;
  wire b29f87;
  wire b29f88;
  wire b29f89;
  wire b29f8a;
  wire b29f8b;
  wire b29f8c;
  wire b29f8d;
  wire b29f8e;
  wire b29f8f;
  wire b29f90;
  wire b29f91;
  wire b29f92;
  wire b29f93;
  wire b29f94;
  wire b29f95;
  wire b29f96;
  wire b29f97;
  wire b29f98;
  wire b29f99;
  wire b29f9a;
  wire b29f9b;
  wire b29f9c;
  wire b29f9d;
  wire b29f9e;
  wire b29f9f;
  wire b29fa0;
  wire b29fa1;
  wire b29fa2;
  wire b29fa3;
  wire b29fa4;
  wire b29fa5;
  wire b29fa6;
  wire b29fa7;
  wire b29fa8;
  wire b29fa9;
  wire b29faa;
  wire b29fab;
  wire b29fac;
  wire b29fad;
  wire b29fae;
  wire b29faf;
  wire b29fb0;
  wire b29fb1;
  wire b29fb2;
  wire b29fb3;
  wire b29fb4;
  wire b29fb5;
  wire b29fb6;
  wire b29fb7;
  wire b29fb8;
  wire b29fb9;
  wire b29fba;
  wire b29fbb;
  wire b29fbc;
  wire b29fbd;
  wire b29fbe;
  wire b29fbf;
  wire b29fc0;
  wire b29fc1;
  wire b29fc2;
  wire b29fc3;
  wire b29fc4;
  wire b29fc5;
  wire b29fc6;
  wire b29fc7;
  wire b29fc8;
  wire b29fc9;
  wire b29fca;
  wire b29fcb;
  wire b29fcc;
  wire b29fcd;
  wire b29fce;
  wire b29fcf;
  wire b29fd0;
  wire b29fd1;
  wire b29fd2;
  wire b29fd3;
  wire b29fd4;
  wire b29fd5;
  wire b29fd6;
  wire b29fd7;
  wire b29fd8;
  wire b29fd9;
  wire b29fda;
  wire b29fdb;
  wire b29fdc;
  wire b29fdd;
  wire b29fde;
  wire b29fdf;
  wire b29fe0;
  wire b29fe1;
  wire b29fe2;
  wire b29fe3;
  wire b29fe4;
  wire b29fe5;
  wire b29fe6;
  wire b29fe7;
  wire b29fe8;
  wire b29fe9;
  wire b29fea;
  wire b29feb;
  wire b29fec;
  wire b29fed;
  wire b29fee;
  wire b29fef;
  wire b29ff0;
  wire b29ff1;
  wire b29ff2;
  wire b29ff3;
  wire b29ff4;
  wire b29ff5;
  wire b29ff6;
  wire b29ff7;
  wire b29ff8;
  wire b29ff9;
  wire b29ffa;
  wire b29ffb;
  wire b29ffc;
  wire b29ffd;
  wire b29ffe;
  wire b29fff;
  wire b2a000;
  wire b2a001;
  wire b2a002;
  wire b2a003;
  wire b2a004;
  wire b2a005;
  wire b2a006;
  wire b2a007;
  wire b2a008;
  wire b2a009;
  wire b2a00a;
  wire b2a00b;
  wire b2a00c;
  wire b2a00d;
  wire b2a00e;
  wire b2a00f;
  wire b2a010;
  wire b2a011;
  wire b2a012;
  wire b2a013;
  wire b2a014;
  wire b2a015;
  wire b2a016;
  wire b2a017;
  wire b2a018;
  wire b2a019;
  wire b2a01a;
  wire b2a01b;
  wire b2a01c;
  wire b2a01d;
  wire b2a01e;
  wire b2a01f;
  wire b2a020;
  wire b29823;
  wire b29824;
  wire b29825;
  wire b29826;
  wire b29827;
  wire b29828;
  wire b29829;
  wire b2982a;
  wire b2982b;
  wire b2982c;
  wire b2982d;
  wire b2982e;
  wire b2982f;
  wire b29830;
  wire b29831;
  wire b29832;
  wire b29833;
  wire b29834;
  wire b29835;
  wire b29836;
  wire b29837;
  wire b29838;
  wire b298a0;
  wire b298a1;
  wire b298a2;
  wire b298a3;
  wire b298a4;
  wire b298a5;
  wire b298a6;
  wire b298a7;
  wire b298a8;
  wire b298a9;
  wire b298aa;
  wire b298ab;
  wire b298ac;
  wire b298ad;
  wire b298ae;
  wire b298af;
  wire b298b0;
  wire b298b1;
  wire b298b2;
  wire b298b3;
  wire b29907;
  wire b29908;
  wire b29909;
  wire b2990a;
  wire b2990b;
  wire b2990c;
  wire b2990d;
  wire b2990e;
  wire b2990f;
  wire b29910;
  wire b29914;
  wire b29915;
  wire b29916;
  wire b29917;
  wire b29918;
  wire b29919;
  wire b2991a;
  wire b2991b;
  wire b2991c;
  wire b2991d;
  wire b2991e;
  wire b29923;
  wire b29924;
  wire b29925;
  wire b29926;
  wire b29927;
  wire b29928;
  wire b29929;
  wire b2992a;
  wire b2992b;
  wire b2992c;
  wire b2992d;
  wire b2992e;
  wire b2992f;
  wire b29930;
  wire b29931;
  wire b29932;
  wire b29933;
  wire b29934;
  wire b29939;
  wire b2993a;
  wire b2993b;
  wire b2993d;
  wire b2993e;
  wire b2993f;
  wire b29940;
  wire b29941;
  wire b29942;
  wire b29943;
  wire b29944;
  wire b29946;
  wire b29947;
  wire b29948;
  wire b29949;
  wire b2994a;
  wire b2994b;
  wire b2994c;
  wire b2994d;
  wire b2994e;
  wire b2994f;
  wire b29950;
  wire b29951;
  wire b29952;
  wire b29953;
  wire b29954;
  wire b29955;
  wire b29956;
  wire b29957;
  wire b29958;
  wire b29959;
  wire b2995a;
  wire b2995b;
  wire b2995c;
  wire b2995d;
  wire b2995e;
  wire b2995f;
  wire b29960;
  wire b29961;
  wire b29962;
  wire b29966;
  wire b29967;
  wire b29969;
  wire b2996a;
  wire b2996b;
  wire b2996c;
  wire b2996d;
  wire b2996e;
  wire b2996f;
  wire b29970;
  wire b29971;
  wire b29972;
  wire b29973;
  wire b29974;
  wire b29975;
  wire b29976;
  wire b29977;
  wire b29978;
  wire b29979;
  wire b2997a;
  wire b2997b;
  wire b2997c;
  wire b2997d;
  wire b2997e;
  wire b2997f;
  wire b29980;
  wire b29981;
  wire b29982;
  wire b29983;
  wire b29984;
  wire b29985;
  wire b29986;
  wire b29987;
  wire b29988;
  wire b29989;
  wire b2998a;
  wire b2998b;
  wire b2998c;
  wire b2998d;
  wire b2998e;
  wire b2998f;
  wire b29990;
  wire b29991;
  wire b29992;
  wire b29993;
  wire b29994;
  wire b29995;
  wire b29996;
  wire b29997;
  wire b29998;
  wire b29999;
  wire b2999a;
  wire b2999b;
  wire b2999c;
  wire b2999d;
  wire b2999e;
  wire b2999f;
  wire b299a0;
  wire b299a1;
  wire b299a2;
  wire b299a3;
  wire b299a4;
  wire b299a5;
  wire b299a6;
  wire b299a7;
  wire b299a8;
  wire b299a9;
  wire b299aa;
  wire b299ab;
  wire b299ac;
  wire b299ad;
  wire b299ae;
  wire b299af;
  wire b299b0;
  wire b299cb;
  wire b299cc;
  wire b299cd;
  wire b299ce;
  wire b299cf;
  wire b299d0;
  wire b299d1;
  wire b299d2;
  wire b299d3;
  wire b299d4;
  wire b299d5;
  wire b299d6;
  wire b299d7;
  wire b299d8;
  wire b299d9;
  wire b299da;
  wire b299db;
  wire b299dc;
  wire b299dd;
  wire b299de;
  wire b299df;
  wire b299e0;
  wire b299e1;
  wire b299e2;
  wire b299e3;
  wire b299e4;
  wire b299e5;
  wire b299e6;
  wire b299e7;
  wire b299e8;
  wire b299e9;
  wire b299ea;
  wire b299eb;
  wire b299ec;
  wire b299ed;
  wire b299ee;
  wire b299ef;
  wire b299f0;
  wire b299f1;
  wire b299f2;
  wire b299f3;
  wire b299f4;
  wire b299f5;
  wire b299ff;
  wire b29a19;
  wire b29a1a;
  wire b29a1b;
  wire b29a1c;
  wire b29a1d;
  wire b29a1e;
  wire b29a1f;
  wire b29a20;
  wire b29a21;
  wire b29a22;
  wire b29a3c;
  wire b29a3d;
  wire b29a3e;
  wire b29a3f;
  wire b29a40;
  wire b29a41;
  wire b29a42;
  wire b29a43;
  wire b29a44;
  wire b29a45;
  wire b29a46;
  wire b29a47;
  wire b29a48;
  wire b29a49;
  wire b29a4a;
  wire b29a4b;
  wire b29a4c;
  wire b29a4d;
  wire b29a4e;
  wire b29a4f;
  wire b29a50;
  wire b29a51;
  wire b29a52;
  wire b29a53;
  wire b29a54;
  wire b29a55;
  wire b29a56;
  wire b29a57;
  wire b29a58;
  wire b29a59;
  wire b29a5a;
  wire b29a5b;
  wire b29a5c;
  wire b29a5d;
  wire b29a62;
  wire b29a63;
  wire b29a64;
  wire b29a65;
  wire b29a66;
  wire b29a67;
  wire b29a68;
  wire b29a69;
  wire b29a6a;
  wire b29a6b;
  wire b29a6c;
  wire b29a6d;
  wire b29a6e;
  wire b29a6f;
  wire b29a76;
  wire b29a77;
  wire b29a78;
  wire b29a79;
  wire b29a7a;
  wire b29a7b;
  wire b29a7c;
  wire b29a7d;
  wire b29a7e;
  wire b29a82;
  wire b29a83;
  wire b29a84;
  wire b29a85;
  wire b29a86;
  wire b29a87;
  wire b29a88;
  wire b29a89;
  wire b29a8a;
  wire b29a8b;
  wire b29a8c;
  wire b29a8d;
  wire b29a8e;
  wire b29a8f;
  wire b29a90;
  wire b29a91;
  wire b29a92;
  wire b29a93;
  wire b29a94;
  wire b29a95;
  wire b29a96;
  wire b29a97;
  wire b29a98;
  wire b29a99;
  wire b29a9a;
  wire b29a9b;
  wire b29a9c;
  wire b29a9d;
  wire b29a9e;
  wire b29a9f;
  wire b29aa0;
  wire b29aa1;
  wire b29aa2;
  wire b29aa3;
  wire b29aa4;
  wire b29aa5;
  wire b29aa6;
  wire b29aa7;
  wire b29aa8;
  wire b29aa9;
  wire b29aaa;
  wire b29aab;
  wire b29aac;
  wire b29aad;
  wire b29aae;
  wire b29aaf;
  wire b29ab0;
  wire b29ab1;
  wire b29ab2;
  wire b29ab3;
  wire b29ab4;
  wire b29ab5;
  wire b29ab6;
  wire b29ab7;
  wire b29ab8;
  wire b29ab9;
  wire b29aba;
  wire b29abb;
  wire b29abc;
  wire b29abd;
  wire b29abe;
  wire b29abf;
  wire b29ac0;
  wire b29ac1;
  wire b29ac2;
  wire b29ac3;
  wire b29ac4;
  wire b29ac5;
  wire b29ac6;
  wire b29ac7;
  wire b29ae2;
  wire b29ae3;
  wire b29ae4;
  wire b29ae5;
  wire b29ae6;
  wire b29ae7;
  wire b29ae8;
  wire b29ae9;
  wire b29aea;
  wire b29aef;
  wire b29b08;
  wire b29b09;
  wire b29b0a;
  wire b29b0b;
  wire b29b0c;
  wire b29b0d;
  wire b29b0e;
  wire b29b0f;
  wire b29b10;
  wire b29b11;
  wire b29b12;
  wire b29b16;
  wire b29b17;
  wire b29b18;
  wire b29b19;
  wire b29b1a;
  wire b29b1b;
  wire b29b1c;
  wire b29b1d;
  wire b29b1e;
  wire b29b1f;
  wire b29b20;
  wire b29b21;
  wire b29b22;
  wire b29b23;
  wire b29b24;
  wire b29b25;
  wire b29b26;
  wire b29b27;
  wire b29b28;
  wire b29b29;
  wire b29b31;
  wire b29b32;
  wire b29b33;
  wire b29b34;
  wire b29b35;
  wire b29b36;
  wire b29b5f;
  wire b29b60;
  wire b29b61;
  wire v845668;
  wire b0d8fd;
  wire b0c0fd;
  wire b0c0fe;
  wire b0c0ff;
  wire d5edb8;
  wire adaeba;
  wire adaebb;
  wire adaebc;
  wire adaebd;
  wire adaebe;
  wire adaebf;
  wire adaec0;
  wire adaec1;
  wire adaec2;
  wire adaec3;
  wire adaec4;
  wire adaec5;
  wire adaec6;
  wire adaec7;
  wire adaec8;
  wire adaec9;
  wire adaeca;
  wire adaecb;
  wire adaecc;
  wire adaecd;
  wire adaece;
  wire adaecf;
  wire adaed0;
  wire adaed1;
  wire adaed2;
  wire adaed3;
  wire adaed4;
  wire adaed5;
  wire adaed6;
  wire adaed7;
  wire adaed8;
  wire adaed9;
  wire adaeda;
  wire adaedb;
  wire adaedc;
  wire adaedd;
  wire adaede;
  wire adaedf;
  wire adaee0;
  wire adaee1;
  wire adaee2;
  wire adaee3;
  wire adaee4;
  wire adaee5;
  wire adaee6;
  wire adaee7;
  wire adaee8;
  wire adaee9;
  wire adaeea;
  wire adaeeb;
  wire adaeec;
  wire adaeed;
  wire adaeee;
  wire adaeef;
  wire adaef0;
  wire adaef1;
  wire adaef2;
  wire adaef3;
  wire adaef4;
  wire adaef5;
  wire adaef6;
  wire adaef7;
  wire adaef8;
  wire adaef9;
  wire adaefa;
  wire adaefb;
  wire adaefc;
  wire adaefd;
  wire adaefe;
  wire adaeff;
  wire adaf00;
  wire adaf01;
  wire adaf02;
  wire adaf03;
  wire adaf04;
  wire adaf05;
  wire adaf06;
  wire adaf07;
  wire adaf08;
  wire adaf09;
  wire adaf0a;
  wire adaf0b;
  wire adaf0c;
  wire adaf0d;
  wire adaf0e;
  wire adaf0f;
  wire adaf10;
  wire adaf11;
  wire adaf12;
  wire adaf13;
  wire adaf14;
  wire adaf15;
  wire adaf16;
  wire adaf17;
  wire adaf18;
  wire adaf19;
  wire adaf1a;
  wire adaf1b;
  wire adaf1c;
  wire v94aab7;
  wire v856555;
  wire af3c10;
  wire af3c11;
  wire af3c12;
  wire af3c13;
  wire af3c14;
  wire af3c15;
  wire af3c16;
  wire v877992;
  wire v8567b4;
  wire af3c17;
  wire af3c18;
  wire af3c19;
  wire af3c1a;
  wire af3c1c;
  wire af3c1d;
  wire af3c1f;
  wire af3c20;
  wire af3c21;
  wire af3c22;
  wire af3c23;
  wire af3c24;
  wire af3c25;
  wire af3c26;
  wire af3c27;
  wire af3c28;
  wire af3c29;
  wire af3c2a;
  wire af3c2b;
  wire af3c2c;
  wire af3c2d;
  wire af3c2e;
  wire af3c2f;
  wire af3c30;
  wire af3c31;
  wire af3c32;
  wire af3c33;
  wire af3c34;
  wire af3c35;
  wire af3c36;
  wire af3c37;
  wire af3c38;
  wire af3c39;
  wire af3c3a;
  wire af3c3b;
  wire af3c3c;
  wire af3c3d;
  wire af3c3e;
  wire af3c3f;
  wire af3c40;
  wire af3c41;
  wire af3c42;
  wire af3c43;
  wire af3c44;
  wire af3c45;
  wire af3c46;
  wire af3c47;
  wire v85f3c3;
  wire v856b00;
  wire af3c48;
  wire af3c49;
  wire af3c4a;
  wire af3c4b;
  wire af3c4c;
  wire af3c4d;
  wire af3c4e;
  wire af3c4f;
  wire af3c50;
  wire af3c51;
  wire af3c52;
  wire af3c53;
  wire af3c54;
  wire af3c55;
  wire af3c56;
  wire af3c57;
  wire af3c58;
  wire af3c59;
  wire af3c5a;
  wire af3c5b;
  wire af3c5c;
  wire af3c5d;
  wire af3c5e;
  wire af3c5f;
  wire af3c60;
  wire af3c61;
  wire af3c62;
  wire af3c63;
  wire af3c64;
  wire af3c65;
  wire af3c66;
  wire af3c67;
  wire af3c68;
  wire c0730a;
  wire af3c69;
  wire af3c6a;
  wire af3c6b;
  wire af3c6c;
  wire af3c6d;
  wire af3c6e;
  wire af3c6f;
  wire af3c70;
  wire af3c71;
  wire af3c72;
  wire af3c73;
  wire af3c79;
  wire af3c7a;
  wire af3c7b;
  wire af3c7d;
  wire af3c7f;
  wire af3c80;
  wire af3c81;
  wire af3485;
  wire af3486;
  wire af3487;
  wire af3488;
  wire af3489;
  wire af348a;
  wire af348b;
  wire af348c;
  wire af348d;
  wire af348e;
  wire af348f;
  wire af3490;
  wire af3491;
  wire af3492;
  wire af3493;
  wire af3494;
  wire af3495;
  wire af3496;
  wire af3497;
  wire af3498;
  wire af3499;
  wire af349a;
  wire af349b;
  wire af349c;
  wire af349d;
  wire af349e;
  wire af349f;
  wire af34a0;
  wire af34a1;
  wire af34a2;
  wire af34a3;
  wire af34a4;
  wire af34a5;
  wire af34a6;
  wire af34a7;
  wire af34a8;
  wire af34a9;
  wire af34aa;
  wire af34ab;
  wire af34ac;
  wire af34ad;
  wire af34ae;
  wire af34af;
  wire af34b0;
  wire af34b1;
  wire af34b2;
  wire af34b3;
  wire af34b4;
  wire af34b5;
  wire af34b6;
  wire af34b7;
  wire af34b8;
  wire af34b9;
  wire af34ba;
  wire af34bb;
  wire af34bc;
  wire af34bd;
  wire af34be;
  wire af34bf;
  wire af34c0;
  wire af34c1;
  wire af34c2;
  wire af34c3;
  wire af34c4;
  wire af34c5;
  wire af34c6;
  wire af34c7;
  wire af34c8;
  wire af34c9;
  wire af34ca;
  wire af34cb;
  wire af34cc;
  wire af34cd;
  wire af34ce;
  wire af34cf;
  wire af34d0;
  wire af34d1;
  wire af34d2;
  wire af34d3;
  wire af34d4;
  wire af34d5;
  wire af34d6;
  wire af34d7;
  wire af34d8;
  wire af34d9;
  wire af34da;
  wire af34db;
  wire af34dc;
  wire af34dd;
  wire af34de;
  wire af34df;
  wire af34e0;
  wire af34e1;
  wire af34e2;
  wire af34e3;
  wire af34e4;
  wire af34e5;
  wire af34e6;
  wire af34e7;
  wire af34e8;
  wire af34e9;
  wire af34ea;
  wire af34eb;
  wire af34ec;
  wire af34ed;
  wire af34ee;
  wire af34ef;
  wire af34f0;
  wire af34f1;
  wire af34f2;
  wire af34f3;
  wire af34f4;
  wire af34f5;
  wire af34f6;
  wire af34f7;
  wire af34f8;
  wire af34f9;
  wire af34fa;
  wire af34fb;
  wire af34fc;
  wire af34fd;
  wire af34fe;
  wire af34ff;
  wire af3500;
  wire af3501;
  wire af3502;
  wire af3503;
  wire af3504;
  wire af3505;
  wire af3506;
  wire af3507;
  wire af3508;
  wire af3509;
  wire af350a;
  wire af350b;
  wire af350c;
  wire af350d;
  wire af350e;
  wire af350f;
  wire af3510;
  wire af3511;
  wire v845642;
  wire af3518;
  wire af3519;
  wire af351a;
  wire af352c;
  wire af352d;
  wire af352e;
  wire af352f;
  wire af3530;
  wire af3531;
  wire af3532;
  wire af3533;
  wire af3534;
  wire af3535;
  wire af3536;
  wire af3537;
  wire af3538;
  wire af3539;
  wire af353f;
  wire af3540;
  wire af3541;
  wire af3546;
  wire af3547;
  wire af3548;
  wire af354b;
  wire af354c;
  wire af354d;
  wire af354e;
  wire af354f;
  wire af3550;
  wire af3551;
  wire af3552;
  wire af3558;
  wire af355e;
  wire af355f;
  wire af3560;
  wire af3561;
  wire af3562;
  wire af3563;
  wire af3564;
  wire af3565;
  wire af3566;
  wire af3567;
  wire af3568;
  wire af3569;
  wire af356a;
  wire af356b;
  wire af356c;
  wire af356d;
  wire af356e;
  wire af356f;
  wire af3570;
  wire af3571;
  wire af3572;
  wire af3573;
  wire af3574;
  wire af3575;
  wire af3576;
  wire af3577;
  wire af3578;
  wire af3579;
  wire af357a;
  wire af357b;
  wire af357c;
  wire af357d;
  wire af357e;
  wire af357f;
  wire af3580;
  wire af3581;
  wire af3582;
  wire af3583;
  wire af3584;
  wire af3585;
  wire af3586;
  wire af3587;
  wire af3588;
  wire af3589;
  wire af358a;
  wire af358b;
  wire af358c;
  wire af358d;
  wire af358e;
  wire af358f;
  wire af3590;
  wire af3591;
  wire af3594;
  wire af3595;
  wire af3596;
  wire af3597;
  wire af3598;
  wire af3599;
  wire af359a;
  wire af359b;
  wire af359c;
  wire af359d;
  wire af359e;
  wire af359f;
  wire af35a0;
  wire af35a1;
  wire af35a2;
  wire af35a3;
  wire af35a4;
  wire af35a5;
  wire af35a6;
  wire af35a7;
  wire af35a8;
  wire af35a9;
  wire af35aa;
  wire af35ab;
  wire af35ac;
  wire af35ad;
  wire af35ae;
  wire af35af;
  wire af35b0;
  wire af35b1;
  wire af35b2;
  wire af35b3;
  wire af35b4;
  wire af35b5;
  wire af35b6;
  wire af35b7;
  wire af35b8;
  wire af35b9;
  wire af35ba;
  wire af35bb;
  wire af35bc;
  wire af35bd;
  wire af35be;
  wire af35bf;
  wire af35c0;
  wire af35c1;
  wire af35c2;
  wire af35c3;
  wire af35c4;
  wire af35c5;
  wire ab0acb;
  wire ab0acc;
  wire ab0acd;
  wire ab0ace;
  wire ab0acf;
  wire ab0ad0;
  wire ab0ad1;
  wire ab0ad2;
  wire ab0ad6;
  wire ab0adc;
  wire ab0add;
  wire ab0ade;
  wire ab0adf;
  wire ab0ae0;
  wire ab0ae1;
  wire ab0ae2;
  wire ab0ae3;
  wire ab0ae4;
  wire ab0ae5;
  wire ab0ae6;
  wire ab0aeb;
  wire ab0aec;
  wire ab0aed;
  wire ab0aee;
  wire ab0aef;
  wire ab0af0;
  wire ab0af1;
  wire ab0af2;
  wire ab0af3;
  wire ab0af4;
  wire ab0af5;
  wire ab0af6;
  wire ab0af7;
  wire ab0af9;
  wire ab0afa;
  wire ab0afb;
  wire ab0b00;
  wire ab0b01;
  wire ab0b02;
  wire ab0b03;
  wire ab0b04;
  wire ab0b09;
  wire ab0b0a;
  wire ab0b0b;
  wire ab0b0c;
  wire ab0b0d;
  wire ab0b0e;
  wire ab0b0f;
  wire ab0b10;
  wire ab0b11;
  wire ab0b15;
  wire ab0b16;
  wire ab0b17;
  wire ab0b18;
  wire ab0b19;
  wire ab0b21;
  wire ab0b22;
  wire ab0b23;
  wire ab0b24;
  wire ab0b2d;
  wire ab0b2e;
  wire ab0b2f;
  wire ab0b30;
  wire ab0b31;
  wire ab0b32;
  wire ab0b33;
  wire ab0b34;
  wire ab0b35;
  wire ab0b36;
  wire ab0b37;
  wire ab0b38;
  wire ab0b39;
  wire ab0b3a;
  wire ab0b3b;
  wire ab0b3c;
  wire ab0b3d;
  wire ab0b3e;
  wire ab0b3f;
  wire ab0b40;
  wire ab0b44;
  wire ab0b45;
  wire ab0b46;
  wire ab0b48;
  wire ab0b49;
  wire ab0b4a;
  wire ab0b4b;
  wire ab0b4c;
  wire ab0b4d;
  wire ab0b4e;
  wire ab0b4f;
  wire ab0b50;
  wire ab0b51;
  wire ab0b52;
  wire ab0b53;
  wire ab0b54;
  wire ab0b55;
  wire ab0b56;
  wire ab0b57;
  wire ab0b58;
  wire ab0b59;
  wire ab0b5a;
  wire ab0b5b;
  wire ab0b5c;
  wire ab0b5d;
  wire ab0b5e;
  wire ab0b5f;
  wire ab0b60;
  wire ab0b61;
  wire ab0b62;
  wire ab0b63;
  wire ab0b64;
  wire ab0b65;
  wire ab0b66;
  wire ab0b67;
  wire ab0b68;
  wire ab0b69;
  wire ab0b6a;
  wire ab0b6b;
  wire ab0b6c;
  wire ab0b6d;
  wire ab0b6e;
  wire ab0b6f;
  wire ab0b70;
  wire ab0b71;
  wire ab0b78;
  wire ab0b79;
  wire ab0b7a;
  wire ab0b7b;
  wire ab0b7c;
  wire ab0b7d;
  wire ab0b7e;
  wire ab0b7f;
  wire ab0b80;
  wire ab0b81;
  wire ab0b82;
  wire ab0b83;
  wire ab0b84;
  wire ab0b85;
  wire ab0b86;
  wire ab0b87;
  wire ab0b88;
  wire ab0b89;
  wire ab0b8a;
  wire ab0b8b;
  wire ab0b8c;
  wire ab0b8d;
  wire ab0b8e;
  wire ab0b8f;
  wire ab0b90;
  wire ab0b91;
  wire ab0b92;
  wire ab0b93;
  wire ab0b94;
  wire ab0b95;
  wire ab0b96;
  wire ab0b97;
  wire ab0b98;
  wire ab0b99;
  wire ab0b9a;
  wire ab0ba1;
  wire ab0ba2;
  wire ab0ba3;
  wire ab0ba4;
  wire ab0ba5;
  wire ab0ba6;
  wire ab0ba7;
  wire ab0ba8;
  wire ab0ba9;
  wire ab0baa;
  wire ab0bab;
  wire ab0bac;
  wire ab0bad;
  wire ab0bae;
  wire ab0baf;
  wire ab0bb0;
  wire ab0bb1;
  wire ab0bb2;
  wire ab0bb3;
  wire ab0bb4;
  wire ab0bb5;
  wire ab0bb6;
  wire ab0bb7;
  wire ab0bb8;
  wire ab0bb9;
  wire ab0bba;
  wire ab0bbb;
  wire ab0bbc;
  wire ab0bbd;
  wire ab0bbe;
  wire ab0bbf;
  wire ab0bc2;
  wire ab0bc3;
  wire ab0bc4;
  wire ab0bc5;
  wire v845662;
  wire ab0bc6;
  wire ab0bc7;
  wire ab0bc8;
  wire ab0bc9;
  wire ab0bca;
  wire ab0bcb;
  wire ab0bcc;
  wire ab0bcd;
  wire ab0bd3;
  wire ab0bd4;
  wire ab0bd5;
  wire ab0bd6;
  wire ab0bd7;
  wire ab0bd8;
  wire ab0bd9;
  wire ab0bda;
  wire ab0bdb;
  wire ab0bdc;
  wire ab0bdd;
  wire ab0bde;
  wire ab0bdf;
  wire ab0be0;
  wire ab0be1;
  wire ab0be2;
  wire ab0be3;
  wire ab0be4;
  wire ab0be5;
  wire ab0be6;
  wire ab0be7;
  wire ab0be8;
  wire ab0be9;
  wire ab0bea;
  wire ab0beb;
  wire ab0bec;
  wire ab0bed;
  wire ab0bee;
  wire ab0bef;
  wire ab0bf0;
  wire ab0bf1;
  wire ab0bf2;
  wire ab0bf3;
  wire ab0bf4;
  wire ab0bf5;
  wire ab0bf6;
  wire ab0bf7;
  wire ab0bf8;
  wire ab0bf9;
  wire ab0bfa;
  wire ab0bfb;
  wire ab0bfc;
  wire ab0bfd;
  wire ab0bfe;
  wire ab0bff;
  wire ab0c00;
  wire ab0c01;
  wire ab0c02;
  wire ab0c03;
  wire ab0c04;
  wire ab0c05;
  wire ab0c06;
  wire ab0c07;
  wire ab0c08;
  wire ab0c09;
  wire ab0c0a;
  wire ab0c0b;
  wire ab0c0c;
  wire ab0c0d;
  wire ab0c0e;
  wire ab0c0f;
  wire ab0c10;
  wire ab0c11;
  wire ab0c12;
  wire ab0c13;
  wire ab0c14;
  wire ab0c15;
  wire ab0c16;
  wire ab0c17;
  wire ab0c18;
  wire ab0c19;
  wire ab0c1a;
  wire ab0c1b;
  wire ab0c1c;
  wire ab0c1d;
  wire ab0c1e;
  wire ab0c1f;
  wire ab0c20;
  wire ab0c21;
  wire ab0c22;
  wire ab0c23;
  wire ab0c24;
  wire ab0c25;
  wire ab0c26;
  wire ab0c27;
  wire ab0c28;
  wire ab0c29;
  wire ab0c2a;
  wire ab0c2b;
  wire ab0c2c;
  wire ab0c2d;
  wire ab0c2e;
  wire ab0c2f;
  wire ab0c30;
  wire ab0c31;
  wire ab0c32;
  wire ab0c33;
  wire ab0c34;
  wire ab0c35;
  wire ab0c3c;
  wire ab0c3d;
  wire ab0c3e;
  wire ab0c3f;
  wire ab0c40;
  wire ab0c41;
  wire ab0c42;
  wire ab0c43;
  wire ab0c44;
  wire ab0c45;
  wire ab0c46;
  wire ab0c47;
  wire ab0c48;
  wire ab0c49;
  wire ab0c4a;
  wire ab0c58;
  wire ab0c59;
  wire ab0c5a;
  wire ab0c5b;
  wire ab0c5c;
  wire ab0c5d;
  wire ab0c5e;
  wire ab0c5f;
  wire ab0c60;
  wire ab0c61;
  wire ab0c62;
  wire ab0c63;
  wire ab0c64;
  wire ab0c65;
  wire ab0c69;
  wire ab0c6a;
  wire ab0c6b;
  wire ab0c6c;
  wire ab0c6d;
  wire ab0c6e;
  wire ab0c6f;
  wire ab0c70;
  wire ab0c71;
  wire ab0c72;
  wire ab0c73;
  wire ab0c74;
  wire ab0c75;
  wire ab0c76;
  wire ab0c77;
  wire ab0c78;
  wire ab0c79;
  wire ab0c7a;
  wire ab0c7b;
  wire ab0c7c;
  wire ab0c7d;
  wire ab0c7e;
  wire ab0c7f;
  wire ab0c80;
  wire ab0c81;
  wire ab0c82;
  wire ab0c83;
  wire ab0c84;
  wire ab0c85;
  wire ab0c86;
  wire ab0c87;
  wire ab0c88;
  wire ab0c89;
  wire ab0c8a;
  wire ab0c8b;
  wire ab0c8c;
  wire ab0c8d;
  wire ab0c8e;
  wire ab0c8f;
  wire ab0c90;
  wire ab0c91;
  wire ab0c92;
  wire ab0c93;
  wire ab0c94;
  wire ab0c95;
  wire ab0c96;
  wire ab0c97;
  wire ab0c98;
  wire ab0c99;
  wire ab0c9a;
  wire ab0c9b;
  wire ab0c9c;
  wire ab0c9d;
  wire ab0c9e;
  wire ab0c9f;
  wire ab0ca0;
  wire ab0ca1;
  wire ab0ca2;
  wire ab0ca3;
  wire ab0ca4;
  wire ab0ca5;
  wire ab0ca6;
  wire ab0ca7;
  wire ab0ca8;
  wire ab0ca9;
  wire ab0caa;
  wire ab0cab;
  wire ab0cac;
  wire ab0cad;
  wire ab0cae;
  wire ab0caf;
  wire ab0cb0;
  wire ab0cb1;
  wire ab0cb2;
  wire ab0cb3;
  wire ab0cb4;
  wire ab0cb5;
  wire ab0cb6;
  wire ab0cb7;
  wire ab0cb8;
  wire ab0cb9;
  wire ab0cba;
  wire ab0cbb;
  wire ab0cbc;
  wire ab0cbd;
  wire ab0cbe;
  wire ab0cbf;
  wire ab0cc0;
  wire ab0cc1;
  wire ab0cc2;
  wire ab0cc3;
  wire ab0cc4;
  wire ab0cc5;
  wire ab0cc6;
  wire ab0cc7;
  wire ab0cc8;
  wire ab0cc9;
  wire ab0cca;
  wire ab0cce;
  wire ab0ccf;
  wire ab0cd0;
  wire ab0cd1;
  wire ab0cd2;
  wire ab0cd3;
  wire ab0cd4;
  wire ab0cd5;
  wire ab0cd6;
  wire ab0cd7;
  wire ab0cd8;
  wire ab0cd9;
  wire ab0cda;
  wire ab0cdb;
  wire ab0cdc;
  wire ab0cdd;
  wire ab0cde;
  wire ab0cdf;
  wire ab0ce0;
  wire ab0ce1;
  wire ab0ce2;
  wire ab0ce3;
  wire ab0ce4;
  wire ab0ce5;
  wire ab0ce6;
  wire ab0ce7;
  wire ab0ce8;
  wire ab0ce9;
  wire ab0cea;
  wire ab0ceb;
  wire ab0cec;
  wire ab0ced;
  wire ab0cee;
  wire ab0cef;
  wire ab0cf0;
  wire ab0cf1;
  wire ab0cf2;
  wire ab0cf3;
  wire ab0cf4;
  wire ab0cf5;
  wire ab0cf6;
  wire ab0cf7;
  wire ab0cf8;
  wire ab0cf9;
  wire ab0cfa;
  wire ab0cfb;
  wire ab0cfc;
  wire ab0cfd;
  wire ab0cfe;
  wire ab0cff;
  wire ab0d00;
  wire ab0d01;
  wire ab0d02;
  wire ab0d03;
  wire ab0d04;
  wire ab0d05;
  wire ab0d06;
  wire ab0d07;
  wire ab050b;
  wire ab050c;
  wire ab050d;
  wire ab050e;
  wire ab050f;
  wire ab0510;
  wire ab0511;
  wire ab0512;
  wire ab0513;
  wire ab0514;
  wire ab0515;
  wire ab0516;
  wire ab0517;
  wire ab0518;
  wire ab0519;
  wire ab051a;
  wire ab051b;
  wire ab051c;
  wire ab051d;
  wire ab051e;
  wire ab051f;
  wire ab0520;
  wire ab0521;
  wire ab0522;
  wire ab0523;
  wire ab0524;
  wire ab0525;
  wire ab0526;
  wire ab0527;
  wire ab0528;
  wire ab0529;
  wire ab052a;
  wire ab052b;
  wire ab052c;
  wire ab052d;
  wire ab052e;
  wire ab052f;
  wire ab0530;
  wire ab0531;
  wire ab0532;
  wire ab0533;
  wire ab0534;
  wire ab0538;
  wire ab0539;
  wire ab053a;
  wire ab053b;
  wire ab053c;
  wire ab053d;
  wire ab053e;
  wire ab053f;
  wire ab0540;
  wire ab0541;
  wire ab0546;
  wire ab0547;
  wire ab0548;
  wire ab0549;
  wire ab054a;
  wire ab054b;
  wire ab054c;
  wire ab054d;
  wire ab054e;
  wire ab054f;
  wire ab0550;
  wire ab0551;
  wire ab0552;
  wire ab0553;
  wire ab0554;
  wire ab0555;
  wire ab055a;
  wire ab055b;
  wire ab055c;
  wire ab055d;
  wire ab055e;
  wire ab055f;
  wire ab0560;
  wire ab0561;
  wire ab0562;
  wire ab0563;
  wire ab0564;
  wire ab0565;
  wire ab0566;
  wire ab056a;
  wire ab056b;
  wire ab056c;
  wire ab056d;
  wire ab056e;
  wire ab056f;
  wire ab0570;
  wire ab0571;
  wire ab0572;
  wire ab0573;
  wire ab0574;
  wire ab0575;
  wire ab0576;
  wire ab0577;
  wire ab0578;
  wire ab0579;
  wire ab057a;
  wire ab057b;
  wire ab057c;
  wire ab057d;
  wire ab057e;
  wire ab057f;
  wire ab0580;
  wire ab0581;
  wire ab0582;
  wire ab0583;
  wire ab0584;
  wire ab0585;
  wire ab0586;
  wire ab0587;
  wire ab0588;
  wire ab0589;
  wire ab058a;
  wire ab058b;
  wire ab058c;
  wire ab058d;
  wire ab058e;
  wire ab058f;
  wire ab0590;
  wire ab0591;
  wire ab0592;
  wire ab0593;
  wire ab0594;
  wire ab0595;
  wire ab0596;
  wire ab0597;
  wire ab0598;
  wire ab0599;
  wire ab059a;
  wire ab059b;
  wire ab059c;
  wire ab059d;
  wire ab059e;
  wire ab059f;
  wire ab05a0;
  wire ab05a1;
  wire ab05a2;
  wire ab05a3;
  wire ab05a4;
  wire ab05a5;
  wire ab05a6;
  wire ab05a7;
  wire ab05a8;
  wire ab05a9;
  wire ab05aa;
  wire ab05ab;
  wire ab05ac;
  wire ab05ad;
  wire ab05ae;
  wire ab05af;
  wire ab05b0;
  wire ab05b1;
  wire ab05b2;
  wire ab05b3;
  wire ab05b4;
  wire ab05b5;
  wire ab05b6;
  wire ab05b7;
  wire ab05b8;
  wire ab05b9;
  wire ab05ba;
  wire ab05bb;
  wire ab05bc;
  wire ab05bd;
  wire ab05be;
  wire ab05bf;
  wire ab05c0;
  wire ab05c1;
  wire ab05c2;
  wire ab05c3;
  wire ab05c4;
  wire ab05c5;
  wire ab05c6;
  wire ab05c7;
  wire ab05c8;
  wire ab05c9;
  wire ab05ca;
  wire ab05cb;
  wire ab05cc;
  wire ab05cd;
  wire ab05ce;
  wire ab05cf;
  wire ab05d0;
  wire ab05d1;
  wire ab05d2;
  wire ab05d3;
  wire ab05d4;
  wire ab05d5;
  wire ab05d6;
  wire ab05d7;
  wire ab05d8;
  wire ab05d9;
  wire ab05da;
  wire ab05db;
  wire ab05dc;
  wire ab05dd;
  wire ab05de;
  wire ab05df;
  wire ab05e0;
  wire ab05e1;
  wire ab05e2;
  wire ab05e3;
  wire ab05e4;
  wire ab05e5;
  wire ab05e6;
  wire ab05e7;
  wire ab05e8;
  wire ab05e9;
  wire ab05ea;
  wire ab05eb;
  wire ab05ec;
  wire ab05ed;
  wire ab05ee;
  wire ab05ef;
  wire ab05f0;
  wire ab05f1;
  wire ab05f2;
  wire ab05f3;
  wire ab05f4;
  wire ab05f5;
  wire ab05f6;
  wire ab05f7;
  wire ab05f8;
  wire ab05f9;
  wire ab05fa;
  wire ab05fb;
  wire ab05fc;
  wire ab05fd;
  wire ab05fe;
  wire ab05ff;
  wire ab0600;
  wire ab0601;
  wire ab0602;
  wire ab0603;
  wire ab0604;
  wire ab0605;
  wire ab0606;
  wire ab0607;
  wire ab0608;
  wire ab0609;
  wire ab060a;
  wire ab060b;
  wire ab060c;
  wire ab060d;
  wire ab060e;
  wire ab060f;
  wire ab0610;
  wire ab0611;
  wire ab0612;
  wire ab0613;
  wire ab0614;
  wire ab0615;
  wire ab0616;
  wire ab0617;
  wire ab0618;
  wire ab0619;
  wire ab061a;
  wire ab061b;
  wire ab061c;
  wire ab061d;
  wire ab061e;
  wire ab061f;
  wire ab0620;
  wire ab0621;
  wire ab0622;
  wire ab0623;
  wire ab0624;
  wire ab0625;
  wire ab0626;
  wire ab0627;
  wire ab0628;
  wire ab0629;
  wire ab062a;
  wire ab062b;
  wire ab062c;
  wire ab062d;
  wire ab062e;
  wire ab062f;
  wire ab0630;
  wire ab0631;
  wire ab0632;
  wire ab0633;
  wire ab0634;
  wire ab0635;
  wire ab0636;
  wire ab0637;
  wire ab0638;
  wire ab0639;
  wire ab063a;
  wire ab063b;
  wire ab063c;
  wire ab063d;
  wire ab063e;
  wire ab063f;
  wire ab0640;
  wire ab0641;
  wire ab0642;
  wire ab0643;
  wire ab0644;
  wire ab0645;
  wire ab0646;
  wire ab0647;
  wire ab0648;
  wire ab0649;
  wire ab064a;
  wire ab064b;
  wire ab064c;
  wire ab064d;
  wire ab064e;
  wire ab064f;
  wire ab0650;
  wire ab0651;
  wire ab0652;
  wire ab0653;
  wire ab0654;
  wire ab0655;
  wire ab0656;
  wire ab066a;
  wire ab066b;
  wire ab066c;
  wire ab066d;
  wire ab066e;
  wire ab066f;
  wire ab0670;
  wire ab0671;
  wire ab0672;
  wire ab0673;
  wire ab0674;
  wire ab0675;
  wire ab0676;
  wire ab0677;
  wire ab0678;
  wire ab0679;
  wire ab067a;
  wire ab067b;
  wire ab067c;
  wire ab067d;
  wire ab067e;
  wire ab067f;
  wire ab0680;
  wire ab0681;
  wire ab0682;
  wire ab0683;
  wire ab0684;
  wire ab0685;
  wire ab0686;
  wire ab0687;
  wire ab0688;
  wire ab0689;
  wire ab068c;
  wire ab068d;
  wire ab068e;
  wire ab068f;
  wire ab0690;
  wire ab0692;
  wire ab0699;
  wire ab069a;
  wire ab069b;
  wire ab069c;
  wire ab069d;
  wire ab069e;
  wire ab069f;
  wire ab06a0;
  wire ab06a2;
  wire ab06a3;
  wire ab06a4;
  wire ab06a5;
  wire ab06a6;
  wire ab06a7;
  wire ab06a8;
  wire ab06a9;
  wire ab06aa;
  wire ab06ab;
  wire ab06ac;
  wire ab06ad;
  wire ab06ae;
  wire ab06af;
  wire ab06b0;
  wire ab06b1;
  wire ab06b2;
  wire ab06b3;
  wire ab06b4;
  wire ab06b5;
  wire ab06b6;
  wire ab06b7;
  wire ab06b8;
  wire ab06b9;
  wire ab06ba;
  wire ab06bb;
  wire ab06bc;
  wire ab06bd;
  wire ab06be;
  wire ab06bf;
  wire ab06c0;
  wire ab06c1;
  wire ab06c2;
  wire ab06c3;
  wire ab06c4;
  wire ab06c5;
  wire ab06c6;
  wire ab06c7;
  wire ab06c8;
  wire ab06c9;
  wire ab06ca;
  wire ab06cb;
  wire ab06cc;
  wire ab06cd;
  wire ab06ce;
  wire ab06cf;
  wire ab06d0;
  wire ab06d1;
  wire ab06d2;
  wire ab06d3;
  wire ab06d4;
  wire ab06d5;
  wire ab06d6;
  wire ab06d7;
  wire ab06d8;
  wire ab06d9;
  wire ab06da;
  wire ab06db;
  wire ab06dc;
  wire ab06dd;
  wire ab06de;
  wire ab06df;
  wire ab06e0;
  wire ab06e1;
  wire ab06e2;
  wire ab06e3;
  wire ab06e4;
  wire ab06e5;
  wire ab06e6;
  wire ab06e7;
  wire ab06e8;
  wire ab06e9;
  wire ab06ea;
  wire ab06eb;
  wire ab06ec;
  wire ab06ed;
  wire ab06ee;
  wire ab06ef;
  wire ab06f0;
  wire ab06f1;
  wire ab06f2;
  wire ab06f3;
  wire ab06f4;
  wire ab06f5;
  wire ab06f6;
  wire ab06f7;
  wire ab06f8;
  wire ab06f9;
  wire ab06fa;
  wire ab06fb;
  wire ab06fc;
  wire ab06fd;
  wire ab06fe;
  wire ab06ff;
  wire ab0700;
  wire ab0701;
  wire ab0702;
  wire ab0703;
  wire ab0704;
  wire ab0712;
  wire ab0713;
  wire ab0714;
  wire ab0715;
  wire ab0716;
  wire ab0717;
  wire ab0718;
  wire ab0719;
  wire ab071a;
  wire ab071b;
  wire ab071c;
  wire ab071d;
  wire ab071e;
  wire ab0722;
  wire ab072e;
  wire ab072f;
  wire ab0730;
  wire ab0731;
  wire ab0732;
  wire ab0733;
  wire ab0734;
  wire ab0735;
  wire ab0736;
  wire ab0737;
  wire ab0738;
  wire ab0739;
  wire ab073a;
  wire ab073b;
  wire ab073c;
  wire ab073d;
  wire ab073e;
  wire ab073f;
  wire ab0740;
  wire ab0741;
  wire ab0742;
  wire ab0743;
  wire ab0744;
  wire ab0745;
  wire ab0746;
  wire ab0747;
  wire ab0748;
  wire ab0749;
  wire ab074a;
  wire ab074b;
  wire ab074c;
  wire ab074d;
  wire ab0754;
  wire ab0755;
  wire ab0756;
  wire ab0757;
  wire ab0758;
  wire ab0759;
  wire ab075a;
  wire ab075b;
  wire ab075c;
  wire ab075d;
  wire ab075e;
  wire ab075f;
  wire ab076a;
  wire ab076b;
  wire ab076c;
  wire aa0e0a;
  wire v868347;
  wire aa0e0b;
  wire aa0e0c;
  wire a60140;
  wire a60141;
  wire a60142;
  wire a60143;
  wire a60144;
  wire a60145;
  wire a60146;
  wire a60147;
  wire a60164;
  wire a60165;
  wire a60166;
  wire a60167;
  wire a60168;
  wire a60169;
  wire a6016a;
  wire a6016b;
  wire a6016c;
  wire a6016d;
  wire a6016e;
  wire a6016f;
  wire a60170;
  wire a60171;
  wire a60172;
  wire a60173;
  wire a60174;
  wire a60175;
  wire a60176;
  wire a60177;
  wire a60178;
  wire a60179;
  wire a60184;
  wire a60185;
  wire a60186;
  wire a60187;
  wire a60188;
  wire a60189;
  wire a6018a;
  wire a6018b;
  wire a6018c;
  wire a6018d;
  wire a60192;
  wire a60193;
  wire a60194;
  wire a60195;
  wire a60196;
  wire a60197;
  wire a60198;
  wire a60199;
  wire a6019a;
  wire a6019b;
  wire a601a6;
  wire a5f9c2;
  wire a5f9c3;
  wire a5f9c4;
  wire a5f9c5;
  wire a5f9c6;
  wire a5f9c7;
  wire a5f9c8;
  wire a5f9c9;
  wire a5f9ca;
  wire a5f9cb;
  wire a5f9d9;
  wire a5f9da;
  wire a5f9db;
  wire a5f9dc;
  wire a5f9dd;
  wire a5f9de;
  wire a5f9df;
  wire a5f9e0;
  wire a5f9e1;
  wire a5f9e7;
  wire a5f9e8;
  wire a5f9e9;
  wire a5f9f4;
  wire a5f9f5;
  wire a5f9f6;
  wire a5f9f7;
  wire a5f9f8;
  wire a5f9f9;
  wire a5f9fa;
  wire a5fa00;
  wire a5fa01;
  wire a5fa02;
  wire a5fa0e;
  wire a5fa0f;
  wire a5fa10;
  wire a5fa11;
  wire a5fa12;
  wire a5fa13;
  wire a5fa14;
  wire a5fa15;
  wire a5fa16;
  wire a5fa1a;
  wire a5fa1b;
  wire a5fa1c;
  wire a5fa1d;
  wire a5fa1e;
  wire a5fa1f;
  wire a5fa20;
  wire a5fa21;
  wire a5fa22;
  wire a5fa23;
  wire v845641;
  wire a5fa25;
  wire a5fa26;
  wire a5fa27;
  wire a5fa28;
  wire a5fa2b;
  wire a5fa2d;
  wire a5fa2e;
  wire a5fa37;
  wire a5fa41;
  wire a5fa42;
  wire a5fa55;
  wire a5fa56;
  wire a5fa57;
  wire a5fa58;
  wire a5fa59;
  wire a5fa5a;
  wire a5fa5b;
  wire a5fa5c;
  wire a5fa5d;
  wire a5fa5e;
  wire a5fa5f;
  wire a5fa60;
  wire a5fa61;
  wire a5fa62;
  wire a5fa63;
  wire a5fa64;
  wire a5fa65;
  wire a5fa66;
  wire a5fa67;
  wire a5fa68;
  wire a5fa69;
  wire a5fa6a;
  wire a5fa6b;
  wire a5fa6c;
  wire a5fa6d;
  wire a5fa6e;
  wire a5fa6f;
  wire a5fa70;
  wire a5fa71;
  wire a5fa86;
  wire a5fa87;
  wire a5fa88;
  wire a5fa89;
  wire a5fa8a;
  wire a5fa8b;
  wire a5fa8c;
  wire a5fa9e;
  wire a5faaa;
  wire a5faab;
  wire a5faac;
  wire a5faad;
  wire a5faae;
  wire a5faaf;
  wire a5fab0;
  wire a5fab1;
  wire a5fab2;
  wire a5fab3;
  wire a5fab4;
  wire a5fabb;
  wire a5fabc;
  wire a5fad1;
  wire a5fad2;
  wire a5fad3;
  wire a5fad4;
  wire a5fad5;
  wire a5fad6;
  wire a5fad7;
  wire a5fae2;
  wire a5fae3;
  wire a5fae4;
  wire a5fae5;
  wire a5fae6;
  wire a5fae7;
  wire a5fae8;
  wire a5fae9;
  wire a5faea;
  wire a5faeb;
  wire a5fafb;
  wire a5fafc;
  wire a5fafd;
  wire a5fb02;
  wire a5fb03;
  wire a5fb10;
  wire a5fb11;
  wire a5fb12;
  wire a5fb13;
  wire a5fb14;
  wire a5fb1b;
  wire a5fb1c;
  wire a5fb1d;
  wire a5fb1e;
  wire a5fb1f;
  wire a5fb20;
  wire a5fb21;
  wire a5fb22;
  wire a5fb23;
  wire a5fb26;
  wire a5fb27;
  wire a5fb28;
  wire a5fb29;
  wire a5fb2a;
  wire a5fb2b;
  wire a5fb2c;
  wire a5fb2d;
  wire v84564d;
  wire a5fb2e;
  wire a5fb2f;
  wire a5fb30;
  wire a5fb31;
  wire a5fb32;
  wire a5fb33;
  wire a5fb34;
  wire a5fb35;
  wire a5fb36;
  wire a5fb37;
  wire a5fb4c;
  wire a5fb4d;
  wire a5fb54;
  wire a5fb5d;
  wire a5fb5e;
  wire a5fb5f;
  wire a5fb60;
  wire a5fb61;
  wire a5fb62;
  wire a5fb63;
  wire a5fb64;
  wire a5fb65;
  wire a5fb66;
  wire a5fb67;
  wire a5fb68;
  wire a5fb69;
  wire a5fb6a;
  wire a5fb6b;
  wire a5fb6c;
  wire a5fb6d;
  wire a5fb6e;
  wire a5fb6f;
  wire a5fb70;
  wire a5fb71;
  wire a5fb72;
  wire a5fb73;
  wire a5fb74;
  wire a5fb75;
  wire a5fb76;
  wire a5fb77;
  wire a5fb78;
  wire a5fb79;
  wire a5fb7a;
  wire a5fb7b;
  wire a5fb7c;
  wire a5fb7d;
  wire a5fb7e;
  wire a5fb7f;
  wire a5fb80;
  wire a5fb81;
  wire a5fb82;
  wire a5fb83;
  wire a5fb84;
  wire a5fb85;
  wire a5fb86;
  wire a5fb87;
  wire a5fb88;
  wire a5fb89;
  wire a5fb8a;
  wire a5fb8b;
  wire a5fb8c;
  wire a5fb8d;
  wire a5fb8e;
  wire a5fb8f;
  wire a5fb90;
  wire a5fb91;
  wire a5fb92;
  wire a5fb93;
  wire a5fb94;
  wire a5fb95;
  wire a5fb96;
  wire a5fb97;
  wire a5fb98;
  wire a5fb99;
  wire a5fb9a;
  wire a5fb9b;
  wire a5fb9c;
  wire d615cf;
  wire a5fb9d;
  wire a5fb9e;
  wire a5fb9f;
  wire a5fba0;
  wire a5fba1;
  wire a5fba2;
  wire a5fba3;
  wire a5fba4;
  wire a5fba5;
  wire a5fba6;
  wire a5fba7;
  wire a5fba8;
  wire a5fba9;
  wire a5fbaa;
  wire a5fbab;
  wire a5fbac;
  wire a5fbad;
  wire a5fbae;
  wire a5fbaf;
  wire a5fbb0;
  wire a5fbb1;
  wire a5fbb2;
  wire a5fbb3;
  wire a5fbb4;
  wire a5fbb5;
  wire a5fbb6;
  wire a5fbb7;
  wire a5fbb8;
  wire a5fbb9;
  wire a5fbba;
  wire a5fbbb;
  wire a5fbbc;
  wire a5fbbd;
  wire a5fbbe;
  wire a5fbbf;
  wire a5fbc0;
  wire a5fbc1;
  wire a5fbc2;
  wire a5fbc3;
  wire a5fbc4;
  wire a5fbc5;
  wire a5fbc6;
  wire a5fbc7;
  wire a5fbc8;
  wire a5fbc9;
  wire a5fbca;
  wire a5fbcb;
  wire a5fbcc;
  wire a5fbcd;
  wire a5fbce;
  wire a5fbd3;
  wire a5fbd4;
  wire a5fbd5;
  wire a5fbd6;
  wire a5fbd7;
  wire a5fbd8;
  wire a5fbd9;
  wire a5fbda;
  wire a5fbdb;
  wire a5fbdc;
  wire a5fbdd;
  wire a5fbde;
  wire a5fbdf;
  wire a5fbe0;
  wire a5fbe1;
  wire a5fbe2;
  wire a5fbe3;
  wire a5fbe4;
  wire a5fbe5;
  wire a5fbe6;
  wire a5fbe7;
  wire a5fbe8;
  wire a5fbe9;
  wire a5fbea;
  wire a5fbeb;
  wire a5fbec;
  wire a5fbed;
  wire a5fbee;
  wire a5fbef;
  wire a5fbf0;
  wire a5fbf1;
  wire a5fbf2;
  wire a5fbf3;
  wire a5fbf4;
  wire a5fbf5;
  wire a5fbf6;
  wire a5fbf7;
  wire a5fbf8;
  wire a5fbf9;
  wire a5fbfa;
  wire a5fbfb;
  wire a5fbfc;
  wire a5fbfd;
  wire a5fbfe;
  wire a5fbff;
  wire a5fc00;
  wire a5fc01;
  wire a5fc02;
  wire a5fc03;
  wire a5fc04;
  wire a5fc05;
  wire a5fc06;
  wire a5fc07;
  wire a5fc08;
  wire a5fc09;
  wire a5fc0a;
  wire a5fc0b;
  wire a5fc0c;
  wire a5fc0d;
  wire a5fc0e;
  wire a5fc0f;
  wire a5fc10;
  wire a5fc11;
  wire a5fc12;
  wire a5fc13;
  wire a5fc14;
  wire a5fc15;
  wire a5fc17;
  wire a5fc18;
  wire a5fc19;
  wire a5fc1a;
  wire a5fc1b;
  wire a5fc1c;
  wire a5fc1d;
  wire a5fc1e;
  wire a5fc1f;
  wire a5fc20;
  wire a5fc21;
  wire a5fc22;
  wire a5fc23;
  wire a5fc24;
  wire a5fc25;
  wire a5fc26;
  wire a5fc27;
  wire a5fc28;
  wire a5fc29;
  wire a5fc2a;
  wire a5fc2b;
  wire a5fc2c;
  wire a5fc2d;
  wire a5fc2e;
  wire a5fc2f;
  wire a5fc30;
  wire a5fc31;
  wire a5fc38;
  wire a5fc39;
  wire a5fc3a;
  wire a5fc3b;
  wire a5fc3d;
  wire a5fc3e;
  wire a5fc3f;
  wire a5fc40;
  wire a5fc41;
  wire a5fc42;
  wire a5fc43;
  wire a5fc44;
  wire a5fc45;
  wire a5fc46;
  wire a5fc47;
  wire a5fc48;
  wire a5fc49;
  wire a5fc4a;
  wire a5fc4b;
  wire a5fc4c;
  wire a5fc4d;
  wire a5fc4e;
  wire a5fc4f;
  wire a5fc50;
  wire a5fc51;
  wire a5fc52;
  wire a5fc53;
  wire a5fc54;
  wire a5fc55;
  wire a5fc56;
  wire a5fc57;
  wire a5fc58;
  wire a5fc59;
  wire a5fc5a;
  wire a5fc5b;
  wire a5fc5c;
  wire a5fc5d;
  wire a5fc5e;
  wire a5fc5f;
  wire a5fc60;
  wire a5fc61;
  wire a5fc62;
  wire a5fc63;
  wire a5fc64;
  wire a5fc65;
  wire a5fc66;
  wire a5fc67;
  wire a5fc68;
  wire a5fc69;
  wire a5fc6a;
  wire a5fc6b;
  wire a5fc6c;
  wire a5fc6d;
  wire a5fc6e;
  wire a5fc6f;
  wire a5fc70;
  wire a5fc71;
  wire a5fc72;
  wire a5fc73;
  wire a5fc74;
  wire a5fc75;
  wire a5fc76;
  wire a5fc77;
  wire a5fc78;
  wire a5fc79;
  wire a5fc7a;
  wire a5fc7b;
  wire a5fc7c;
  wire a5fc7d;
  wire a5fc7e;
  wire a5fc7f;
  wire a5fc80;
  wire a5fc81;
  wire a5fc82;
  wire a5fc83;
  wire a5fc84;
  wire a5fc85;
  wire a5fc86;
  wire a5fc87;
  wire a5fc88;
  wire a5fc89;
  wire a5fc8a;
  wire a5fc8b;
  wire a5fc8c;
  wire a5fc8d;
  wire a5fc8e;
  wire a5fc8f;
  wire a5fc90;
  wire a5fc91;
  wire a5fc92;
  wire a5fc93;
  wire a5fc94;
  wire a5fc95;
  wire a5fc96;
  wire a5fc97;
  wire a5fc9b;
  wire a5fc9c;
  wire a5fc9d;
  wire a5fc9e;
  wire a5fc9f;
  wire a5fca0;
  wire a5fca1;
  wire a5fca2;
  wire a5fca3;
  wire a5fca4;
  wire a5fca5;
  wire a5fca6;
  wire a5fca7;
  wire a5fca8;
  wire a5fca9;
  wire a5fcaa;
  wire a5fcab;
  wire a5fcac;
  wire a5fcad;
  wire a5fcae;
  wire a5fcb0;
  wire a5fcb3;
  wire a5fcb4;
  wire a5fcb5;
  wire a5fcb6;
  wire a5fcbb;
  wire a5fcbc;
  wire a5fcbd;
  wire a5fcbe;
  wire a5fcbf;
  wire a5fcc0;
  wire a5fcc1;
  wire a5fcc2;
  wire a5fcc3;
  wire a5fcc4;
  wire a5fcc5;
  wire a5fcc6;
  wire a5fcc7;
  wire a5fcc8;
  wire a5fcc9;
  wire a5fcca;
  wire a5fccb;
  wire a5fccc;
  wire a5fccd;
  wire a5fcce;
  wire a5fccf;
  wire a5fcd0;
  wire a5fcd1;
  wire a5fcd2;
  wire a5fcd3;
  wire a5fcd4;
  wire a5fcd5;
  wire a5fcd6;
  wire a5fcd7;
  wire a5fcd8;
  wire a5fcd9;
  wire a5fcda;
  wire a5fcdb;
  wire a5fcdc;
  wire a5fcdd;
  wire a5fcde;
  wire a5fcdf;
  wire a5fce0;
  wire a5fce1;
  wire a5fce2;
  wire a5fce3;
  wire a5fce4;
  wire a5fce5;
  wire a5fce6;
  wire a5fce7;
  wire a5fce8;
  wire a5fce9;
  wire a5fcea;
  wire a5fceb;
  wire a5fcef;
  wire a5fcf0;
  wire a5fcf1;
  wire a5fcf2;
  wire a5fcf3;
  wire a5fcf4;
  wire a5fcf5;
  wire a5fcf6;
  wire a5fcf7;
  wire a5fcf8;
  wire a5fcf9;
  wire a5fcfa;
  wire a5fcfb;
  wire a5fcfc;
  wire a5fcfd;
  wire a5fcfe;
  wire a5fcff;
  wire a5fd00;
  wire a5fd01;
  wire a5fd02;
  wire a5fd03;
  wire a5fd05;
  wire a5fd08;
  wire a5fd09;
  wire a5fd0a;
  wire a5fd0b;
  wire a5fd0f;
  wire a5fd10;
  wire a5fd11;
  wire a5fd12;
  wire a5fd13;
  wire a5fd14;
  wire a5fd15;
  wire a5fd16;
  wire a5fd17;
  wire a5fd18;
  wire a5fd19;
  wire a5fd1a;
  wire a5fd1b;
  wire a5fd1c;
  wire a5fd21;
  wire a5fd22;
  wire a5fd23;
  wire a5fd24;
  wire a5fd25;
  wire a5fd26;
  wire a5fd27;
  wire a5fd28;
  wire a5fd34;
  wire a5fd35;
  wire a5fd36;
  wire a5fd37;
  wire a5fd38;
  wire a5fd39;
  wire a5fd3a;
  wire a5fd3b;
  wire a5f6ce;
  wire a5f6cf;
  wire a5f6d0;
  wire a5f6d1;
  wire a5f6d2;
  wire a5f6d3;
  wire a5f6d4;
  wire a5f6d5;
  wire a5f6d6;
  wire a5f6d7;
  wire a5f6d8;
  wire a5f6d9;
  wire a5f6da;
  wire a5f6db;
  wire a5f6dc;
  wire a5f6dd;
  wire a5f6de;
  wire a5f6df;
  wire a5f6e0;
  wire a5f6e1;
  wire a5f6e2;
  wire a5f6e3;
  wire a5f6e4;
  wire a5f6e5;
  wire a5f6e6;
  wire a5f6e7;
  wire a5f6e8;
  wire a5f6e9;
  wire a5f6ea;
  wire a5f6eb;
  wire a5f6ec;
  wire a5f6ed;
  wire a5f6ee;
  wire a5f6ef;
  wire a5f6f0;
  wire a5f6f1;
  wire a5f6f2;
  wire a5f6f3;
  wire a5f6f4;
  wire a5f6f5;
  wire a5f6f6;
  wire a5f6f7;
  wire a5f6f8;
  wire a5f6f9;
  wire a5f6fa;
  wire a5f6fb;
  wire a5f6fc;
  wire a5f6fd;
  wire a5f703;
  wire a5f704;
  wire a5f705;
  wire a5f706;
  wire a5f707;
  wire a5f708;
  wire a5f709;
  wire a5f70a;
  wire a5f70b;
  wire a5f70c;
  wire a5f70d;
  wire a5f70e;
  wire a5f70f;
  wire a5f710;
  wire a5f711;
  wire a5f712;
  wire a5f713;
  wire a5f714;
  wire a5f715;
  wire a5f716;
  wire a5f717;
  wire a5f718;
  wire a5f719;
  wire a5f71a;
  wire a5f71b;
  wire a5f71d;
  wire a5f71e;
  wire a5f71f;
  wire a5f720;
  wire a5f721;
  wire a5f722;
  wire a5f723;
  wire a5f724;
  wire a5f726;
  wire a5f727;
  wire a5f728;
  wire a5f729;
  wire a5f72a;
  wire a5f72b;
  wire a5f72c;
  wire a5f72d;
  wire a5f72e;
  wire a5f72f;
  wire a5f730;
  wire a5f731;
  wire a5f733;
  wire a5f734;
  wire a5f735;
  wire a5f739;
  wire a5f73a;
  wire a5f73b;
  wire a5f73c;
  wire a5f73d;
  wire a5f73e;
  wire a5f73f;
  wire a5f741;
  wire a5f742;
  wire a5f743;
  wire a5f744;
  wire a5f745;
  wire a5f746;
  wire a5f747;
  wire a5f748;
  wire a5f749;
  wire a5f74a;
  wire a5f74b;
  wire a5f74c;
  wire a5f74d;
  wire a5f74e;
  wire a5f74f;
  wire a5f750;
  wire a5f751;
  wire a5f752;
  wire a5f753;
  wire a5f754;
  wire a5f755;
  wire a5f756;
  wire a5f757;
  wire a5f783;
  wire a5f784;
  wire a5f785;
  wire a5f786;
  wire a5f787;
  wire a5f78d;
  wire a5f78e;
  wire a5f795;
  wire a5f796;
  wire a5f797;
  wire a5f798;
  wire a5f7a2;
  wire a5f7a3;
  wire a5f7a4;
  wire a5f7b4;
  wire a5f7ba;
  wire a5f7bb;
  wire a5f7bc;
  wire a5f7be;
  wire a5f7c0;
  wire a5f7c2;
  wire a5f7c3;
  wire a5f7c4;
  wire a5f7cb;
  wire a5f7cd;
  wire a5f7ce;
  wire a5f7cf;
  wire a5f7d0;
  wire a5f7f3;
  wire a5f7f4;
  wire a5f7f5;
  wire a5f7f6;
  wire a5f7f7;
  wire a5f7f8;
  wire a5f7f9;
  wire a5f7fa;
  wire a5f7fb;
  wire a5f7fc;
  wire a5f7fd;
  wire a5f804;
  wire a5f805;
  wire a5f806;
  wire a5f807;
  wire a5f821;
  wire a5f828;
  wire a5f829;
  wire a5f82a;
  wire a5f82b;
  wire a5f82c;
  wire a5f833;
  wire a5f834;
  wire a5f835;
  wire a5f836;
  wire a5f837;
  wire a5f838;
  wire a5f839;
  wire a5f83a;
  wire a5f83b;
  wire a5f83c;
  wire a5f83e;
  wire a5f83f;
  wire a5f840;
  wire a5f841;
  wire a5f842;
  wire a5f843;
  wire a5f844;
  wire a5f845;
  wire a5f855;
  wire a5f856;
  wire a5f857;
  wire a5f858;
  wire a5f861;
  wire a5f862;
  wire a5f863;
  wire a5f864;
  wire a5f86a;
  wire a5f86b;
  wire a5f86c;
  wire a5f86d;
  wire a5f879;
  wire a5f87a;
  wire a5f87b;
  wire a5f87c;
  wire a5f87d;
  wire a5f87f;
  wire a5f880;
  wire a5f881;
  wire a5f882;
  wire a5f883;
  wire a5f884;
  wire a5f885;
  wire a5f886;
  wire a5f887;
  wire a5f888;
  wire a5f8b4;
  wire a5f8b5;
  wire a5f8b6;
  wire a5f8b7;
  wire a5f8b8;
  wire a5f8b9;
  wire a5f8ba;
  wire a5f8bb;
  wire a5f8bc;
  wire a5f8bd;
  wire a5f8be;
  wire a5f8bf;
  wire a5f8c0;
  wire a5f8c1;
  wire a5f8c2;
  wire a5f8c3;
  wire a5f8c4;
  wire a5f8c5;
  wire a5f8c6;
  wire a5f8c7;
  wire a5f8c8;
  wire a5f8c9;
  wire a5f8ca;
  wire a5f8cb;
  wire a5f8cc;
  wire a5f8cd;
  wire a5f8ce;
  wire a5f8cf;
  wire a5f8d0;
  wire a5f8d1;
  wire a5f8d2;
  wire a5f8d3;
  wire a5f8d4;
  wire a5f8d5;
  wire a5f8d6;
  wire a5f8d7;
  wire a5f8d8;
  wire a5f8d9;
  wire a5f8da;
  wire a5f8db;
  wire a5f8dc;
  wire a5f8dd;
  wire a5f8de;
  wire a5f8df;
  wire a5f8e0;
  wire a5f8e1;
  wire a5f8e2;
  wire a5f8e3;
  wire a5f8e4;
  wire a5f8e5;
  wire a5f8e6;
  wire a5f8e7;
  wire a5f8e8;
  wire a5f8e9;
  wire a5f8ea;
  wire a5f8eb;
  wire a5f8ec;
  wire a5f8ed;
  wire a5f8ee;
  wire a5f8ef;
  wire a5f8f0;
  wire a5f8f1;
  wire a5f8f2;
  wire a5f8f3;
  wire a5f8f4;
  wire a5f8f5;
  wire a5f8f6;
  wire a5f8f7;
  wire a5f8f8;
  wire a5f8fd;
  wire a5f8fe;
  wire a5f8ff;
  wire a5f900;
  wire a5f901;
  wire a5f902;
  wire a5f903;
  wire a5f904;
  wire a5f906;
  wire a5f907;
  wire a5f908;
  wire a5f909;
  wire a5f90a;
  wire a5f90b;
  wire a5f90c;
  wire a5f917;
  wire a5f918;
  wire a5f919;
  wire a5f91a;
  wire a5f921;
  wire a5f922;
  wire a5f923;
  wire a5f924;
  wire a5f925;
  wire a5f926;
  wire a5f927;
  wire a5f92c;
  wire a5f92d;
  wire a5f92e;
  wire a5f92f;
  wire a5f930;
  wire a5f931;
  wire a5f932;
  wire a5f933;
  wire a5f934;
  wire a5f935;
  wire a5f936;
  wire a5f937;
  wire a5f938;
  wire a5f939;
  wire a5f93a;
  wire a5f93b;
  wire a5f93c;
  wire a5f93d;
  wire a5f93e;
  wire a5f93f;
  wire a5f940;
  wire a5f941;
  wire a5f942;
  wire a5f943;
  wire a5f944;
  wire a5f945;
  wire a5f946;
  wire a5f947;
  wire a5f948;
  wire a5f949;
  wire a5f94a;
  wire a5f94b;
  wire a5f94c;
  wire a5f94d;
  wire a5f94e;
  wire a5f94f;
  wire a5f950;
  wire a5f951;
  wire a5f952;
  wire a5f953;
  wire a5f954;
  wire a5f955;
  wire a5f956;
  wire a5f957;
  wire a5f958;
  wire a5f959;
  wire a5f95a;
  wire a5f95b;
  wire a5f95c;
  wire a5f95d;
  wire a5f95e;
  wire a5f95f;
  wire a5f960;
  wire a5f961;
  wire a5f962;
  wire a5f964;
  wire a5f965;
  wire a5f966;
  wire a5f967;
  wire a5f968;
  wire a5f969;
  wire a5f96a;
  wire a5f96b;
  wire a5f96c;
  wire a5f96d;
  wire a5f96e;
  wire a5f96f;
  wire a5f970;
  wire a5f971;
  wire a5f972;
  wire a5f973;
  wire a5f974;
  wire a5f975;
  wire a5f976;
  wire a5f977;
  wire a5f978;
  wire a5f979;
  wire a5f97a;
  wire a5f97b;
  wire a5f97c;
  wire a5f97d;
  wire a5f97e;
  wire a5f97f;
  wire a5f980;
  wire a5f981;
  wire a5f982;
  wire a5f983;
  wire a5f984;
  wire a5f985;
  wire a5f986;
  wire a5f987;
  wire a5f988;
  wire a5f989;
  wire a5f98a;
  wire a5f98b;
  wire a5f98c;
  wire a5f98d;
  wire a5f98e;
  wire a5f98f;
  wire a5f990;
  wire a5f991;
  wire a5f992;
  wire a5f993;
  wire a5f994;
  wire a5f995;
  wire a5f996;
  wire a5f997;
  wire a5f998;
  wire a5f999;
  wire a5f99a;
  wire a5f99b;
  wire a5f99c;
  wire a5f99d;
  wire a5f99e;
  wire a5f9a0;
  wire a5f9a1;
  wire a5f9a2;
  wire a5f9a3;
  wire a5f9a4;
  wire a5f9a5;
  wire a5f9a6;
  wire a5f9a7;
  wire a5f9a8;
  wire a5f1ac;
  wire a5f1ad;
  wire a5f1ae;
  wire a5f1af;
  wire a5f1b0;
  wire a5f1b1;
  wire a5f1b2;
  wire a5f1b3;
  wire a5f1b4;
  wire a5f1b5;
  wire a5f1b6;
  wire a5f1b7;
  wire a5f1b8;
  wire a5f1b9;
  wire a5f1bd;
  wire a5f1be;
  wire a5f1bf;
  wire a5f1c0;
  wire a5f1c1;
  wire a5f1c2;
  wire a5f1c3;
  wire a5f1c4;
  wire a5f1c8;
  wire a5f1c9;
  wire a5f1ca;
  wire a5f1cb;
  wire a5f1cc;
  wire a5f1cd;
  wire a5f1ce;
  wire a5f1cf;
  wire a5f1d0;
  wire a5f1d1;
  wire a5f1d2;
  wire a5f1d3;
  wire a5f1d4;
  wire a5f1d5;
  wire a5f1d6;
  wire a5f1d7;
  wire a5f1d8;
  wire a5f1d9;
  wire a5f1da;
  wire a5f1db;
  wire a5f1dc;
  wire a5f1dd;
  wire a5f1de;
  wire a5f1df;
  wire a5f1e0;
  wire a5f1e1;
  wire a5f1e2;
  wire a5f1e3;
  wire a5f1e4;
  wire a5f1e5;
  wire a5f1e6;
  wire a5f1e7;
  wire a5f1e8;
  wire a5f1e9;
  wire a5f1ea;
  wire a5f1eb;
  wire a5f1ec;
  wire a5f1ed;
  wire a5f1ef;
  wire a5f1f0;
  wire a5f1f1;
  wire a5f1f2;
  wire a5f1f3;
  wire a5f1f4;
  wire a5f1f5;
  wire a5f1f6;
  wire a5f1f7;
  wire a5f1f8;
  wire a5f1f9;
  wire a5f1fa;
  wire a5f1fb;
  wire a5f1fc;
  wire a5f1fd;
  wire a5f1ff;
  wire a5f200;
  wire a5f201;
  wire a5f202;
  wire a5f203;
  wire a5f204;
  wire a5f205;
  wire a5f206;
  wire a5f207;
  wire a5f208;
  wire a5f209;
  wire a5f20a;
  wire a5f20b;
  wire a5f20c;
  wire a5f20d;
  wire a5f20e;
  wire a5f20f;
  wire a5f210;
  wire a5f211;
  wire a5f212;
  wire a5f213;
  wire a5f214;
  wire a5f215;
  wire a5f216;
  wire a5f217;
  wire a5f218;
  wire a5f219;
  wire a5f21a;
  wire a5f21b;
  wire a5f22d;
  wire a5f22e;
  wire a5f22f;
  wire a5f230;
  wire a5f231;
  wire a5f232;
  wire a5f233;
  wire a5f234;
  wire a5f235;
  wire a5f236;
  wire a5f237;
  wire a5f238;
  wire a5f239;
  wire a5f23a;
  wire a5f23b;
  wire a5f23c;
  wire a5f246;
  wire a5f247;
  wire a5f248;
  wire a5f249;
  wire a5f24a;
  wire a5f24b;
  wire a5f24c;
  wire a5f24d;
  wire a5f24e;
  wire a5f24f;
  wire a5f250;
  wire a5f251;
  wire a5f252;
  wire a5f253;
  wire a5f254;
  wire a5f255;
  wire a5f256;
  wire a5f25a;
  wire a5f268;
  wire a5f269;
  wire a5f26a;
  wire a5f26b;
  wire a5f26c;
  wire a5f26d;
  wire a5f26e;
  wire a5f26f;
  wire a5f270;
  wire a5f271;
  wire a5f282;
  wire a5f283;
  wire a5f284;
  wire a5f285;
  wire a5f286;
  wire a5f287;
  wire a5f288;
  wire a5f289;
  wire a5f28a;
  wire a5f28b;
  wire a5f28c;
  wire a5f28d;
  wire a5f28f;
  wire a5f290;
  wire a5f291;
  wire a5f292;
  wire a5f293;
  wire a5f294;
  wire a5f295;
  wire a5f296;
  wire a5f297;
  wire a5f298;
  wire a5f299;
  wire a5f29a;
  wire a5f29b;
  wire a5f29c;
  wire a5f29d;
  wire a5f29e;
  wire a5f29f;
  wire a5f2c7;
  wire a5f2c8;
  wire a5f2c9;
  wire a5f2ca;
  wire a5f2d2;
  wire a5f2d3;
  wire a5f2d4;
  wire a5f2d5;
  wire a5f2d6;
  wire a5f2d7;
  wire a5f2d8;
  wire a5f2d9;
  wire a5f2da;
  wire a5f2db;
  wire a5f2dc;
  wire a5f2dd;
  wire a5f2de;
  wire a5f2df;
  wire a5f2e3;
  wire a5f2e4;
  wire a5f2e5;
  wire a5f2e6;
  wire a5f2e7;
  wire a5f2e8;
  wire a5f2e9;
  wire a5f2ea;
  wire a5f2eb;
  wire a5f2ec;
  wire a5f2ed;
  wire a5f2f1;
  wire a5f2f2;
  wire a5f2f3;
  wire a5f2f4;
  wire a5f2f5;
  wire a5f2f6;
  wire a5f2f7;
  wire a5f2f8;
  wire a5f2f9;
  wire a5f2fa;
  wire a5f2fb;
  wire a5f2fc;
  wire a5f2fd;
  wire a5f2fe;
  wire a5f2ff;
  wire a5f300;
  wire a5f301;
  wire a5f302;
  wire a5f303;
  wire a5f304;
  wire a5f305;
  wire a5f306;
  wire a5f320;
  wire a5f321;
  wire a5f323;
  wire a5f324;
  wire a5f325;
  wire a5f326;
  wire a5f328;
  wire a5f329;
  wire a5f32a;
  wire a5f32c;
  wire a5f32d;
  wire a5f32e;
  wire a5f32f;
  wire a5f330;
  wire a5f331;
  wire a5f332;
  wire a5f333;
  wire a5f334;
  wire a5f335;
  wire a5f343;
  wire a5f344;
  wire a5f345;
  wire a5f346;
  wire a5f35b;
  wire a5f35c;
  wire a5f35d;
  wire a5f35e;
  wire a5f35f;
  wire a5f360;
  wire a5f361;
  wire a5f362;
  wire a5f363;
  wire a5f364;
  wire a5f365;
  wire a5f366;
  wire a5f367;
  wire a5f368;
  wire a5f369;
  wire a5f36a;
  wire a5f36b;
  wire a5f36c;
  wire a5f36d;
  wire a5f36e;
  wire a5f36f;
  wire a5f370;
  wire a5f371;
  wire a5f372;
  wire a5f373;
  wire a5f374;
  wire a5f375;
  wire a5f376;
  wire a5f377;
  wire a5f378;
  wire a5f379;
  wire a5f37a;
  wire a5f37b;
  wire a5f37c;
  wire a5f37d;
  wire a5f37e;
  wire a5f37f;
  wire a5f380;
  wire a5f381;
  wire a5f382;
  wire a5f383;
  wire a5f384;
  wire a5f385;
  wire a5f386;
  wire a5f387;
  wire a5f388;
  wire a5f389;
  wire a5f38a;
  wire a5f38b;
  wire a5f38c;
  wire a5f38d;
  wire a5f38e;
  wire a5f38f;
  wire a5f390;
  wire a5f391;
  wire a5f392;
  wire a5f393;
  wire a5f394;
  wire a5f395;
  wire a5f396;
  wire a5f397;
  wire a5f398;
  wire a5f399;
  wire a5f39a;
  wire a5f39b;
  wire a5f39c;
  wire a5f39d;
  wire a5f39e;
  wire a5f39f;
  wire a5f3a0;
  wire a5f3a1;
  wire a5f3a2;
  wire a5f3a3;
  wire a5f3a4;
  wire a5f3a5;
  wire a5f3a6;
  wire a5f3a7;
  wire a5f3ad;
  wire a5f3ae;
  wire a5f3af;
  wire a5f3b0;
  wire a5f3b1;
  wire a5f3b2;
  wire a5f3b3;
  wire a5f3b4;
  wire a5f3b5;
  wire a5f3b6;
  wire a5f3b7;
  wire a5f3b8;
  wire a5f3b9;
  wire a5f3ba;
  wire a5f3bb;
  wire a5f3bc;
  wire a5f3bd;
  wire a5f3be;
  wire a5f3bf;
  wire a5f3c0;
  wire a5f3c1;
  wire a5f3c2;
  wire a5f3c3;
  wire a5f3c4;
  wire a5f3c5;
  wire a5f3c6;
  wire a5f3c7;
  wire a5f3c8;
  wire a5f3c9;
  wire a5f3ca;
  wire a5f3cb;
  wire a5f3cc;
  wire a5f3cd;
  wire a5f3ce;
  wire a5f3cf;
  wire a5f3d0;
  wire a5f3d1;
  wire a5f3d2;
  wire a5f3d3;
  wire a5f3d4;
  wire a5f3d5;
  wire a5f3d6;
  wire a5f3d7;
  wire a5f3d8;
  wire a5f3d9;
  wire a5f3da;
  wire a5f3db;
  wire a5f3dc;
  wire a5f3dd;
  wire a5f3de;
  wire a5f3ef;
  wire a5f3f0;
  wire a5f3f1;
  wire a5f3f2;
  wire a5f3f3;
  wire a5f3f4;
  wire a5f3f5;
  wire a5f3f6;
  wire a5f3f7;
  wire a5f3f8;
  wire a5f409;
  wire a5f40a;
  wire a5f40b;
  wire a5f40c;
  wire a5f40d;
  wire a5f40e;
  wire a5f41b;
  wire a5f41c;
  wire a5f41d;
  wire a5f41e;
  wire a5f41f;
  wire a5f420;
  wire a5f421;
  wire a5f422;
  wire a5f434;
  wire a5f435;
  wire a5f436;
  wire a5f437;
  wire a5f438;
  wire a5f439;
  wire a5f43a;
  wire a5f43b;
  wire a5f43c;
  wire a5f43d;
  wire a5f43e;
  wire a5f43f;
  wire a5f440;
  wire a5f455;
  wire a5f456;
  wire a5f457;
  wire a5f458;
  wire a5f459;
  wire a5f45a;
  wire a5f45b;
  wire a5f45c;
  wire a5f46d;
  wire a5f46e;
  wire a5f46f;
  wire a5f470;
  wire a5f471;
  wire a5f472;
  wire a5f473;
  wire a5f474;
  wire a5f475;
  wire a5f476;
  wire a5f477;
  wire a5f478;
  wire a5f479;
  wire a5f47a;
  wire a5f47b;
  wire a5f47c;
  wire a5f485;
  wire a5f486;
  wire a5f487;
  wire a5f488;
  wire a5f489;
  wire a5f48a;
  wire a5f490;
  wire a5f491;
  wire a5f492;
  wire a5f493;
  wire a5f494;
  wire a5f495;
  wire a5f496;
  wire a5f4a2;
  wire a5f4a3;
  wire a5f4a4;
  wire a5f4a5;
  wire a5f4a6;
  wire a5f4a7;
  wire a5f4a8;
  wire a5f4b8;
  wire a5f4b9;
  wire a5f4ba;
  wire a5f4c7;
  wire a5f4c8;
  wire a5f4c9;
  wire a5f4ca;
  wire a5f4cb;
  wire a5f4cc;
  wire a5f4cd;
  wire a5f4ce;
  wire a5f4cf;
  wire a5f4d0;
  wire a5f4d1;
  wire a5f4e3;
  wire a5f4e4;
  wire a5f4e5;
  wire a5f4e6;
  wire a5f4e7;
  wire a5f4e8;
  wire a5f4e9;
  wire a5f4ea;
  wire a5f4eb;
  wire a5f4ec;
  wire a5f4ed;
  wire a5f4ee;
  wire a5f4ef;
  wire a5f4f0;
  wire a5f4f1;
  wire a5f4f2;
  wire a5f4f3;
  wire a5f4fa;
  wire a5f4fb;
  wire a5f4fc;
  wire a5f500;
  wire a5f510;
  wire a5f511;
  wire a5f515;
  wire a5f516;
  wire a5f51a;
  wire a5f51b;
  wire a5f51c;
  wire a5f520;
  wire a5f521;
  wire a5f525;
  wire a5f526;
  wire a5f527;
  wire a5f528;
  wire a5f529;
  wire a5f52a;
  wire a5f52b;
  wire a5f52c;
  wire a5f530;
  wire a5f531;
  wire a5f532;
  wire a5f533;
  wire a5f534;
  wire a5f535;
  wire a5f536;
  wire a5f537;
  wire a5f538;
  wire a5f539;
  wire a5f53a;
  wire a5f53b;
  wire a5f53c;
  wire a5f53d;
  wire a5f53e;
  wire a5f53f;
  wire a5f540;
  wire a5f541;
  wire a5f542;
  wire a5f543;
  wire a5f544;
  wire a5f545;
  wire a5f546;
  wire a5f547;
  wire a5f548;
  wire a5f549;
  wire a5f54a;
  wire a5f54b;
  wire a5f54c;
  wire a5f54d;
  wire a5f54e;
  wire a5f555;
  wire a5f556;
  wire a5f557;
  wire a5f558;
  wire a5f559;
  wire a5f55a;
  wire a5f55b;
  wire a5f55c;
  wire a5f560;
  wire a5f561;
  wire a5f565;
  wire a5f566;
  wire a5f567;
  wire a5f568;
  wire a5f569;
  wire a5f56a;
  wire a5f56b;
  wire a5f56c;
  wire a5f56d;
  wire a5f56e;
  wire a5f56f;
  wire a5f570;
  wire a5f571;
  wire a5f572;
  wire a5f573;
  wire a5f574;
  wire a5f575;
  wire a5f576;
  wire a5f577;
  wire a5f57b;
  wire a5f57c;
  wire a5f57d;
  wire a5f57e;
  wire a5f57f;
  wire a5f580;
  wire a5f581;
  wire a5f582;
  wire a5f583;
  wire a5f584;
  wire a5f585;
  wire a5f586;
  wire a5f587;
  wire a5f588;
  wire a5f589;
  wire a5f58a;
  wire a5f58b;
  wire a5f58c;
  wire a5f58d;
  wire a5f58e;
  wire a5f58f;
  wire a5f590;
  wire a5f591;
  wire a5f592;
  wire a5f593;
  wire a5f594;
  wire a5f595;
  wire a5f596;
  wire a5f597;
  wire a5f598;
  wire a5f599;
  wire a5f59a;
  wire a5f5a2;
  wire a5f5a3;
  wire a5f5a8;
  wire a5f5a9;
  wire a5edac;
  wire a5edb6;
  wire a5edb7;
  wire a5edb8;
  wire a5edb9;
  wire a5edba;
  wire a5edbb;
  wire a5edbc;
  wire a5edbe;
  wire a5edbf;
  wire a5edc0;
  wire a5edc1;
  wire a5edc2;
  wire a5edc6;
  wire a5edc7;
  wire a5edc8;
  wire a5edc9;
  wire a5edca;
  wire a5edcb;
  wire a5edcc;
  wire a5edcd;
  wire a5edce;
  wire a5edcf;
  wire a5edd0;
  wire a5edd1;
  wire a5edd2;
  wire a5edd4;
  wire a5edd5;
  wire a5edd6;
  wire a5edd7;
  wire a5edd8;
  wire a5edd9;
  wire a5edda;
  wire a5eddb;
  wire a5eddc;
  wire a5eddd;
  wire a5edde;
  wire a5eddf;
  wire a5ede0;
  wire a5ede1;
  wire a5ede2;
  wire a5ede3;
  wire a5ede4;
  wire a5ede5;
  wire a5ede6;
  wire a5ede7;
  wire a5ede8;
  wire a5ede9;
  wire a5edea;
  wire a5edeb;
  wire a5edec;
  wire a5eded;
  wire a5edee;
  wire a5edef;
  wire a5edf0;
  wire a5edf1;
  wire a5edf2;
  wire a5edf3;
  wire a5edf4;
  wire a5edf5;
  wire a5edf6;
  wire a5edf7;
  wire a5edf8;
  wire a5edf9;
  wire a5edfa;
  wire a5edfb;
  wire a5edfc;
  wire a5edfd;
  wire a5edfe;
  wire a5edff;
  wire a5ee00;
  wire a5ee01;
  wire a5ee02;
  wire a5ee03;
  wire a5ee04;
  wire a5ee05;
  wire a5ee06;
  wire a5ee07;
  wire a5ee08;
  wire a5ee09;
  wire a5ee0a;
  wire a5ee0b;
  wire a5ee0c;
  wire a5ee0d;
  wire a5ee0e;
  wire a5ee0f;
  wire a5ee10;
  wire a5ee11;
  wire a5ee12;
  wire a5ee13;
  wire a5ee14;
  wire a5ee15;
  wire a5ee16;
  wire a5ee17;
  wire a5ee18;
  wire a5ee19;
  wire a5ee1a;
  wire a5ee1b;
  wire a5ee1c;
  wire a5ee1d;
  wire a5ee1e;
  wire a5ee1f;
  wire a5ee20;
  wire a5ee21;
  wire a5ee22;
  wire a5ee23;
  wire a5ee24;
  wire a5ee25;
  wire a5ee26;
  wire a5ee27;
  wire a5ee28;
  wire a5ee29;
  wire a5ee2a;
  wire a5ee2b;
  wire a5ee2c;
  wire a5ee2d;
  wire a5ee2e;
  wire a5ee2f;
  wire a5ee30;
  wire a5ee31;
  wire a5ee32;
  wire a5ee33;
  wire a5ee34;
  wire a5ee35;
  wire a5ee36;
  wire a5ee37;
  wire a5ee38;
  wire a5ee39;
  wire a5ee3a;
  wire a5ee3b;
  wire a5ee3c;
  wire a5ee3d;
  wire a5ee3e;
  wire a5ee3f;
  wire a5ee40;
  wire a5ee41;
  wire a5ee42;
  wire a5ee43;
  wire a5ee44;
  wire a5ee45;
  wire a5ee46;
  wire a5ee47;
  wire a5ee48;
  wire a5ee49;
  wire a5ee4a;
  wire a5ee4b;
  wire a5ee4c;
  wire a5ee4d;
  wire a5ee4e;
  wire a5ee4f;
  wire a5ee50;
  wire a5ee51;
  wire a5ee52;
  wire a5ee53;
  wire a5ee54;
  wire a5ee55;
  wire a5ee56;
  wire a5ee57;
  wire a5ee58;
  wire a5ee59;
  wire a5ee5a;
  wire a5ee5b;
  wire a5ee5c;
  wire a5ee5d;
  wire a5ee5e;
  wire a5ee5f;
  wire a5ee60;
  wire a5ee61;
  wire a5ee62;
  wire a5ee63;
  wire a5ee64;
  wire a5ee65;
  wire a5ee66;
  wire a5ee67;
  wire a5ee68;
  wire a5ee69;
  wire a5ee6a;
  wire a5ee6b;
  wire a5ee6c;
  wire a5ee6d;
  wire a5ee6e;
  wire a5ee6f;
  wire a5ee70;
  wire a5ee71;
  wire a5ee72;
  wire a5ee73;
  wire a5ee74;
  wire a5ee75;
  wire a5ee76;
  wire a5ee77;
  wire a5ee78;
  wire a5ee79;
  wire a5ee7a;
  wire a5ee7b;
  wire a5ee7c;
  wire a5ee7d;
  wire a5ee7e;
  wire a5ee7f;
  wire a5ee80;
  wire a5ee81;
  wire a5ee82;
  wire a5ee83;
  wire a5ee84;
  wire a5ee85;
  wire a5ee86;
  wire a5ee87;
  wire a5ee88;
  wire a5ee89;
  wire a5ee8a;
  wire a5ee8b;
  wire a5ee8c;
  wire a5ee8d;
  wire a5ee8e;
  wire a5ee8f;
  wire a5ee90;
  wire a5ee91;
  wire a5ee92;
  wire a5ee93;
  wire a5ee94;
  wire a5ee95;
  wire a5ee96;
  wire a5ee97;
  wire a5ee98;
  wire a5ee99;
  wire a5ee9a;
  wire a5ee9b;
  wire a5ee9c;
  wire a5ee9d;
  wire a5ee9e;
  wire a5ee9f;
  wire a5eea0;
  wire a5eea1;
  wire a5eea2;
  wire a5eea3;
  wire a5eea4;
  wire a5eea5;
  wire a5eea6;
  wire a5eea7;
  wire a5eea8;
  wire a5eea9;
  wire a5eeaa;
  wire a5eeab;
  wire a5eeac;
  wire a5eead;
  wire a5eeae;
  wire a5eeaf;
  wire a5eeb0;
  wire a5eeb1;
  wire a5eeb2;
  wire a5eeb3;
  wire a5eeb4;
  wire a5eeb5;
  wire a5eeb6;
  wire a5eeb7;
  wire a5eeb8;
  wire a5eeb9;
  wire a5eeba;
  wire a5eebb;
  wire a5eebc;
  wire a5eebd;
  wire a5eebe;
  wire a5eebf;
  wire a5eec0;
  wire a5eec1;
  wire a5eec2;
  wire a5eec3;
  wire a5eec4;
  wire a5eec5;
  wire a5eec6;
  wire a5eec7;
  wire a5eec8;
  wire a5eec9;
  wire a5eeca;
  wire a5eecb;
  wire a5eecc;
  wire a5eecd;
  wire a5eece;
  wire a5eecf;
  wire a5eed0;
  wire a5eed1;
  wire a5eed2;
  wire a5eed3;
  wire a5eed4;
  wire a5eed5;
  wire a5eed6;
  wire a5eeda;
  wire a5eedb;
  wire a5eedc;
  wire a5eedd;
  wire a5eede;
  wire a5eedf;
  wire a5eee1;
  wire a5eee2;
  wire a5eee3;
  wire a5eee7;
  wire a5eee8;
  wire a5eee9;
  wire a5eeea;
  wire a5eeee;
  wire a5eeef;
  wire a5eef0;
  wire a5eef1;
  wire a5eef2;
  wire a5eef3;
  wire a5eef4;
  wire a5eef5;
  wire a5eef6;
  wire a5eef7;
  wire a5eef8;
  wire a5eef9;
  wire a5eefa;
  wire a5ef05;
  wire a5ef06;
  wire a5ef07;
  wire a5ef08;
  wire a5ef09;
  wire a5ef0a;
  wire a5ef0b;
  wire a5ef0c;
  wire a5ef0d;
  wire a5ef0e;
  wire a5ef0f;
  wire a5ef10;
  wire a5ef11;
  wire a5ef12;
  wire a5ef13;
  wire a5ef14;
  wire a5ef15;
  wire a5ef16;
  wire a5ef17;
  wire a5ef18;
  wire a5ef25;
  wire a5ef26;
  wire a5ef27;
  wire a5ef28;
  wire a5ef29;
  wire a5ef2a;
  wire a5ef2b;
  wire a5ef2c;
  wire a5ef2d;
  wire a5ef2e;
  wire a5ef2f;
  wire a5ef30;
  wire a5ef31;
  wire a5ef32;
  wire a5ef33;
  wire a5ef34;
  wire a5ef35;
  wire a5ef36;
  wire a5ef37;
  wire a5ef38;
  wire a5ef39;
  wire a5ef3a;
  wire a5ef3b;
  wire a5ef3c;
  wire a5ef42;
  wire a5ef43;
  wire a5ef44;
  wire a5ef45;
  wire a5ef46;
  wire a5ef47;
  wire a5ef48;
  wire a5ef50;
  wire a5ef51;
  wire a5ef52;
  wire a5ef53;
  wire a5ef58;
  wire a5ef59;
  wire a5ef5a;
  wire a5ef5e;
  wire a5ef5f;
  wire a5ef60;
  wire a5ef61;
  wire a5ef62;
  wire a5ef6b;
  wire a5ef6c;
  wire a5ef6d;
  wire a5ef6e;
  wire a5ef6f;
  wire a5ef70;
  wire a5ef71;
  wire a5ef72;
  wire a5ef73;
  wire a5ef74;
  wire a5ef75;
  wire a5ef76;
  wire a5ef78;
  wire a5ef79;
  wire a5ef7a;
  wire a5ef7b;
  wire a5ef7c;
  wire a5ef7d;
  wire a5ef7e;
  wire a5ef7f;
  wire a5ef80;
  wire a5ef81;
  wire a5ef82;
  wire a5ef83;
  wire a5ef84;
  wire a5ef85;
  wire a5ef86;
  wire a5ef87;
  wire a5ef88;
  wire a5ef89;
  wire a5ef8a;
  wire a5ef8b;
  wire a5ef8c;
  wire a5ef8d;
  wire a5ef8e;
  wire a5ef8f;
  wire a5ef90;
  wire a5ef91;
  wire a5ef92;
  wire a5ef93;
  wire a5ef94;
  wire a5ef95;
  wire a5ef96;
  wire a5ef97;
  wire a5ef98;
  wire a5ef99;
  wire a5ef9a;
  wire a5ef9b;
  wire a5ef9c;
  wire a5ef9d;
  wire a5ef9e;
  wire a5ef9f;
  wire a5efa0;
  wire a5efa1;
  wire a5efa2;
  wire a5efa3;
  wire a5efa4;
  wire a5efa5;
  wire a5efa6;
  wire a5efa7;
  wire a5efa8;
  wire a5efa9;
  wire a5efaa;
  wire a5efab;
  wire a5efac;
  wire a5efad;
  wire a5efae;
  wire a5efaf;
  wire a5efb0;
  wire a5efb1;
  wire a5efb2;
  wire a5efb3;
  wire a5efb4;
  wire a5efb5;
  wire a5efb6;
  wire a5efb7;
  wire a5efb8;
  wire a5efb9;
  wire a5efba;
  wire a5efbb;
  wire a5efbc;
  wire a5efbd;
  wire a5efbe;
  wire a5efbf;
  wire a5efc0;
  wire a5efc1;
  wire a5efc2;
  wire a5efc3;
  wire a5efc4;
  wire a5efc5;
  wire a5efc6;
  wire a5efc7;
  wire a5efc8;
  wire a5efc9;
  wire a5efca;
  wire a5efcb;
  wire a5efcc;
  wire a5efcd;
  wire a5efce;
  wire a5efcf;
  wire a5efd0;
  wire a5efd1;
  wire a5efd2;
  wire a5efd3;
  wire a5efd4;
  wire a5efd5;
  wire a5efd6;
  wire a5efd7;
  wire a5efd8;
  wire a5efd9;
  wire a5efda;
  wire a5efdb;
  wire a5efdc;
  wire a5efdd;
  wire a5efde;
  wire a5efdf;
  wire a5efe0;
  wire a5efe1;
  wire a5efe2;
  wire a5efe3;
  wire a5efe4;
  wire a5efe5;
  wire a5efe6;
  wire a5efe7;
  wire a5efe8;
  wire a5efe9;
  wire a5efea;
  wire a5efeb;
  wire a5efec;
  wire a5efed;
  wire a5eff8;
  wire a5eff9;
  wire a5f00c;
  wire a5f00d;
  wire a5f00e;
  wire a5f00f;
  wire a5f010;
  wire a5f011;
  wire a5f012;
  wire a5f013;
  wire a5f014;
  wire a5f01b;
  wire a5f01c;
  wire a5f01d;
  wire a5f01e;
  wire a5f01f;
  wire a5f020;
  wire a5f021;
  wire a5f022;
  wire a5f023;
  wire a5f024;
  wire a5f025;
  wire a5f026;
  wire a5f027;
  wire a5f028;
  wire a5f029;
  wire a5f02a;
  wire a5f02b;
  wire a5f02c;
  wire a5f02d;
  wire a5f034;
  wire a5f035;
  wire a5f036;
  wire a5f037;
  wire a5f038;
  wire a5f039;
  wire a5f03a;
  wire a5f03b;
  wire a5f03c;
  wire a5f03d;
  wire a5f03e;
  wire a5f03f;
  wire a5f040;
  wire a5f041;
  wire a5f042;
  wire a5f043;
  wire a5f044;
  wire a5f045;
  wire a5f046;
  wire a5f047;
  wire a5f065;
  wire a5f066;
  wire a5f067;
  wire a5f068;
  wire a5f069;
  wire a5f06a;
  wire a5f06b;
  wire a5f06c;
  wire a5f06d;
  wire a5f06e;
  wire a5f06f;
  wire a5f070;
  wire a5f071;
  wire a5f072;
  wire a5f073;
  wire a5f074;
  wire a5f075;
  wire a5f076;
  wire a5f077;
  wire a5f079;
  wire a5f07a;
  wire a5f07b;
  wire a5f07c;
  wire a5f07d;
  wire a5f07e;
  wire a5f07f;
  wire a5f080;
  wire a5f081;
  wire a5f082;
  wire a5f083;
  wire a5f084;
  wire a5f085;
  wire a5f086;
  wire a5f087;
  wire a5f089;
  wire a5f08a;
  wire a5f08b;
  wire a5f08c;
  wire a5f08d;
  wire a5f08e;
  wire a5f08f;
  wire a5f090;
  wire a5f092;
  wire a5f094;
  wire a5f095;
  wire a5f096;
  wire a5f097;
  wire a5f098;
  wire a5f099;
  wire a5f09b;
  wire a5f09c;
  wire a5f09d;
  wire a5f09e;
  wire a5f09f;
  wire a5f0a0;
  wire a5f0a1;
  wire a5f0a2;
  wire a5f0a3;
  wire a5f0a4;
  wire a5f0a5;
  wire a5f0a6;
  wire a5f0a7;
  wire a5f0a8;
  wire a5f0a9;
  wire a5f0aa;
  wire a5f0ab;
  wire a5f0ac;
  wire a5f0ad;
  wire a5f0ae;
  wire a5f0af;
  wire a5f0b0;
  wire a5f0b1;
  wire a5f0c3;
  wire a5f0d0;
  wire a5f0d1;
  wire a5f0d5;
  wire a5f0d9;
  wire a5f0da;
  wire a5f0db;
  wire a5f0dc;
  wire a5f0e5;
  wire a5f0e6;
  wire a5f0eb;
  wire a5f0ec;
  wire a5f0ed;
  wire a5f0ee;
  wire a5f108;
  wire a5f109;
  wire a5f110;
  wire a5f11a;
  wire a5f11b;
  wire a5f11c;
  wire a5f11d;
  wire a5f11e;
  wire a5f11f;
  wire a5f120;
  wire a5f121;
  wire a5f122;
  wire a5f123;
  wire a5f124;
  wire a5f135;
  wire a5f136;
  wire a5f137;
  wire a5f138;
  wire a5f139;
  wire a5f13a;
  wire a5f13b;
  wire a5f13c;
  wire a5f13d;
  wire a5f144;
  wire a5f145;
  wire a5f146;
  wire a5f148;
  wire a5f149;
  wire a5f14a;
  wire a5f14b;
  wire a5f14c;
  wire a5f14d;
  wire a5f14e;
  wire a5f153;
  wire a5f154;
  wire a5f15b;
  wire a5f15c;
  wire a5f15d;
  wire a5f15e;
  wire a5f15f;
  wire a5f160;
  wire a5f161;
  wire a5f162;
  wire a5f163;
  wire a5f164;
  wire a5f16f;
  wire a5f171;
  wire a5f172;
  wire a5f174;
  wire a5f175;
  wire a5f176;
  wire a5f177;
  wire a5f17c;
  wire a5f17d;
  wire a5f17e;
  wire a5f187;
  wire a5f188;
  wire a5f189;
  wire a5f18a;
  wire a5f18b;
  wire a5f18c;
  wire a5f18d;
  wire a5f192;
  wire a5f193;
  wire a5f194;
  wire a5f195;
  wire a5f196;
  wire a5f197;
  wire a5f198;
  wire a5f199;
  wire a5f19a;
  wire a5f1a2;
  wire a5f1a3;
  wire a5f1a4;
  wire a5f1a5;
  wire a5f1a6;
  wire a5f1a7;
  wire a5f1a8;
  wire a5f1a9;
  wire a5e9ad;
  wire a5e9ae;
  wire a5e9b3;
  wire a5e9b4;
  wire a5e9b5;
  wire a5e9b9;
  wire a5e9ba;
  wire a5e9bb;
  wire a5e9bc;
  wire a5e9bd;
  wire a5e9be;
  wire a5e9c0;
  wire a5e9c1;
  wire a5e9c2;
  wire a5e9c3;
  wire a5e9c4;
  wire a5e9c5;
  wire a5e9c6;
  wire a5e9c7;
  wire a5e9c8;
  wire a5e9c9;
  wire a5e9ca;
  wire a5e9cc;
  wire a5e9cd;
  wire a5e9ce;
  wire a5e9cf;
  wire a5e9d0;
  wire a5e9d2;
  wire a5e9d3;
  wire a5e9d4;
  wire a5e9d5;
  wire a5e9d6;
  wire a5e9d7;
  wire a5e9d8;
  wire a5e9d9;
  wire a5e9da;
  wire a5e9db;
  wire a5e9dc;
  wire a5e9dd;
  wire a5e9df;
  wire a5e9e0;
  wire a5e9e1;
  wire a5e9e6;
  wire a5e9e8;
  wire a5e9e9;
  wire a5e9ea;
  wire a5e9eb;
  wire a5e9f1;
  wire a5e9f2;
  wire a5e9f6;
  wire a5e9f7;
  wire a5e9fd;
  wire a5e9fe;
  wire a5e9ff;
  wire a5ea00;
  wire a5ea06;
  wire a5ea07;
  wire a5ea0d;
  wire a5ea0e;
  wire a5ea0f;
  wire a5ea10;
  wire a5ea11;
  wire a5ea12;
  wire a5ea13;
  wire a5ea14;
  wire a5ea15;
  wire a5ea16;
  wire a5ea17;
  wire a5ea18;
  wire a5ea19;
  wire a5ea1a;
  wire a5ea1b;
  wire a5ea1c;
  wire a5ea1d;
  wire a5ea1e;
  wire a5ea1f;
  wire a5ea20;
  wire a5ea21;
  wire a5ea22;
  wire a5ea23;
  wire a5ea24;
  wire a5ea25;
  wire a5ea26;
  wire a5ea27;
  wire a5ea28;
  wire a5ea29;
  wire a5ea2a;
  wire a5ea2b;
  wire a5ea2c;
  wire a5ea2d;
  wire a5ea2e;
  wire a5ea2f;
  wire a5ea30;
  wire a5ea33;
  wire a5ea34;
  wire a5ea35;
  wire a5ea37;
  wire a5ea38;
  wire a5ea39;
  wire a5ea3a;
  wire a5ea3b;
  wire a5ea3c;
  wire a5ea3d;
  wire a5ea3e;
  wire a5ea3f;
  wire a5ea40;
  wire a5ea41;
  wire a5ea42;
  wire a5ea43;
  wire a5ea44;
  wire a5ea45;
  wire a5ea46;
  wire a5ea47;
  wire a5ea48;
  wire a5ea49;
  wire a5ea4a;
  wire a5ea4b;
  wire a5ea4c;
  wire a5ea4d;
  wire a5ea4e;
  wire a5ea4f;
  wire a5ea50;
  wire a5ea51;
  wire a5ea52;
  wire a5ea53;
  wire a5ea54;
  wire a5ea55;
  wire a5ea56;
  wire a5ea57;
  wire a5ea58;
  wire a5ea59;
  wire a5ea5a;
  wire a5ea5b;
  wire a5ea5c;
  wire a5ea5d;
  wire a5ea5e;
  wire a5ea5f;
  wire a5ea60;
  wire a5ea61;
  wire a5ea62;
  wire a5ea63;
  wire a5ea64;
  wire a5ea65;
  wire a5ea66;
  wire a5ea67;
  wire a5ea68;
  wire a5ea69;
  wire a5ea6a;
  wire a5ea6b;
  wire a5ea6c;
  wire a5ea6d;
  wire a5ea6e;
  wire a5ea6f;
  wire a5ea70;
  wire a5ea73;
  wire a5ea74;
  wire a5ea75;
  wire a5ea76;
  wire a5ea77;
  wire a5ea78;
  wire a5ea79;
  wire a5ea7a;
  wire a5ea7b;
  wire a5ea7c;
  wire a5ea7d;
  wire a5ea7e;
  wire a5ea7f;
  wire a5ea80;
  wire a5ea81;
  wire a5ea82;
  wire a5ea83;
  wire a5ea84;
  wire a5ea85;
  wire a5ea86;
  wire a5ea87;
  wire a5ea88;
  wire a5ea89;
  wire a5ea8a;
  wire a5ea8b;
  wire a5ea8c;
  wire a5ea8d;
  wire a5ea8e;
  wire a5ea8f;
  wire a5ea90;
  wire a5ea91;
  wire a5ea92;
  wire a5ea93;
  wire a5ea94;
  wire a5ea95;
  wire a5ea96;
  wire a5ea97;
  wire a5ea98;
  wire a5ea99;
  wire a5ea9a;
  wire a5ea9b;
  wire a5ea9c;
  wire a5ea9d;
  wire a5ea9e;
  wire a5ea9f;
  wire a5eaa0;
  wire a5eaa1;
  wire a5eaa2;
  wire a5eaa3;
  wire a5eaa4;
  wire a5ead0;
  wire a5ead1;
  wire a5ead2;
  wire a5ead3;
  wire a5ead4;
  wire a5ead5;
  wire a5ead6;
  wire a5ead7;
  wire a5eada;
  wire a5eadb;
  wire a5eadc;
  wire a5eadd;
  wire a5eade;
  wire a5eadf;
  wire a5eae4;
  wire a5eae5;
  wire a5eae6;
  wire a5eae7;
  wire a5eae8;
  wire a5eae9;
  wire a5eaea;
  wire a5eaeb;
  wire a5eaec;
  wire a5eaed;
  wire a5eaee;
  wire a5eaef;
  wire a5eaf0;
  wire a5eaf1;
  wire a5eaf2;
  wire a5eaf3;
  wire a5eaf4;
  wire a5eaf5;
  wire a5eafc;
  wire a5eb1c;
  wire a5eb2a;
  wire a5eb2b;
  wire a5eb34;
  wire a5eb35;
  wire a5eb36;
  wire a5eb37;
  wire a5eb38;
  wire a5eb39;
  wire a5eb3a;
  wire a5eb3b;
  wire a5eb3c;
  wire a5eb3d;
  wire a5eb3e;
  wire a5eb3f;
  wire a5eb40;
  wire a5eb41;
  wire a5eb42;
  wire a5eb43;
  wire a5eb44;
  wire a5eb45;
  wire a5eb46;
  wire a5eb47;
  wire a5eb48;
  wire a5eb49;
  wire a5eb4b;
  wire a5eb4c;
  wire a5eb4d;
  wire a5eb4e;
  wire a5eb4f;
  wire a5eb50;
  wire a5eb51;
  wire a5eb52;
  wire a5eb53;
  wire a5eb54;
  wire a5eb6f;
  wire a5eb70;
  wire a5eb74;
  wire a5eb75;
  wire a5eb76;
  wire a5eb82;
  wire a5eb83;
  wire a5eb84;
  wire a5eb85;
  wire a5eb86;
  wire a5eb87;
  wire a5eb88;
  wire a5eb89;
  wire a5eb8a;
  wire a5eb8b;
  wire a5eb8c;
  wire a5eb8d;
  wire a5eb8e;
  wire a5eb8f;
  wire a5eb90;
  wire a5eb91;
  wire a5eb92;
  wire a5eb93;
  wire a5eb94;
  wire a5eb95;
  wire a5eb96;
  wire a5eb97;
  wire a5eb98;
  wire a5eb99;
  wire a5eb9a;
  wire a5eb9b;
  wire a5eb9c;
  wire a5eb9d;
  wire a5eb9e;
  wire a5eb9f;
  wire a5eba0;
  wire a5eba1;
  wire a5eba2;
  wire a5eba3;
  wire a5ebc1;
  wire a5ebc2;
  wire a5ebc3;
  wire a5ebc7;
  wire a5ebc8;
  wire a5ebc9;
  wire a5ebca;
  wire a5ebcb;
  wire a5ebcc;
  wire a5ebdc;
  wire a5ebdd;
  wire a5ebe6;
  wire a5ebe7;
  wire a5ebe8;
  wire a5ebe9;
  wire a5ebea;
  wire a5ebeb;
  wire a5ebec;
  wire a5ebed;
  wire a5ebee;
  wire a5ec18;
  wire a5ec19;
  wire a5ec1e;
  wire a5ec1f;
  wire a5ec20;
  wire a5ec21;
  wire a5ec22;
  wire a5ec23;
  wire a5ec24;
  wire a5ec30;
  wire a5ec31;
  wire a5ec32;
  wire a5ec33;
  wire a9b9d0;
  wire a9b9d1;
  wire a9b9d2;
  wire a9b9d3;
  wire a9b9d4;
  wire a9b9d5;
  wire a9b9d6;
  wire a9b9d7;
  wire a9b9d8;
  wire a9b9d9;
  wire a9b9da;
  wire a9b9db;
  wire a9b9dc;
  wire a9b9dd;
  wire a9b9de;
  wire a9b9df;
  wire a9b9e0;
  wire a9b9e1;
  wire a9b9e2;
  wire a9b9e3;
  wire a9b9e4;
  wire a9b9e5;
  wire a9b9e6;
  wire a9b9e7;
  wire a9b9e8;
  wire a9b9e9;
  wire a9b9ea;
  wire a9b9eb;
  wire a9b9ec;
  wire a9b9ed;
  wire a9b9ee;
  wire a9b9ef;
  wire a9b9f0;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hbusreq2_p;
  input hbusreq2;
  reg hlock2_p;
  input hlock2;
  reg hbusreq3_p;
  input hbusreq3;
  reg hlock3_p;
  input hlock3;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmaster1_p;
  output hmaster1;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg hgrant2_p;
  output hgrant2;
  reg hgrant3_p;
  output hgrant3;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg stateG10_2_p;
  output stateG10_2;
  reg stateG10_3_p;
  output stateG10_3;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;
  reg jx2_p;
  output jx2;

assign a5f044 = hready_p & a5f6cf | !hready_p & a5f043;
assign ab05a7 = hlock0_p & v84563c | !hlock0_p & !b2998c;
assign deac78 = hbusreq2_p & deac72 | !hbusreq2_p & v84565a;
assign cea189 = hmaster1_p & cea86e | !hmaster1_p & cea188;
assign a5f0a3 = hbusreq0_p & a5fc7a | !hbusreq0_p & v84563c;
assign b29970 = hlock2 & b2996e | !hlock2 & b2996f;
assign b29fa7 = hgrant2_p & c3bcfb | !hgrant2_p & !b29ecf;
assign ab05b5 = hlock2 & ab052f | !hlock2 & ab05b4;
assign b8acf1 = hgrant3_p & b8ace2 | !hgrant3_p & b8acf0;
assign a5f0af = hmaster1_p & a5f0ae | !hmaster1_p & v84563c;
assign b2999f = locked_p & c3b6f8 | !locked_p & !v84563c;
assign a5eae4 = hbusreq0_p & a5f24c | !hbusreq0_p & ab0c31;
assign a5f595 = hbusreq3 & a5f591 | !hbusreq3 & a5f594;
assign c3bd9e = hbusreq2_p & c3bd9d | !hbusreq2_p & c3bc7f;
assign a5fc06 = hlock0_p & a5fc03 | !hlock0_p & a5fc05;
assign a5edea = hbusreq1 & a5ede9 | !hbusreq1 & v84563c;
assign ab0638 = hgrant2_p & ab0635 | !hgrant2_p & ab0637;
assign a5f1fa = hlock2_p & a5f1f9 | !hlock2_p & a5f1b5;
assign b2997e = hlock2 & b29907 | !hlock2 & b2997d;
assign b29ec2 = hlock2_p & b29ebc | !hlock2_p & !b29ec1;
assign c3b80c = hbusreq2_p & c3b80b | !hbusreq2_p & c3b809;
assign cea36a = hbusreq2_p & cea367 | !hbusreq2_p & !cea0bf;
assign cea42e = hlock1_p & deac52 | !hlock1_p & !cea3be;
assign ab0538 = hmastlock_p & deac50 | !hmastlock_p & v84563c;
assign a5fb27 = hlock0_p & a5fb26 | !hlock0_p & a5fa2d;
assign cea1c8 = hmaster0_p & cea1c6 | !hmaster0_p & cea1c7;
assign ab06fe = hbusreq2_p & ab0679 | !hbusreq2_p & ab06fd;
assign c3bddf = hmaster0_p & c3bdde | !hmaster0_p & c3bd67;
assign cea1c7 = hmaster1_p & cea860 | !hmaster1_p & cea1c5;
assign a5ee51 = hlock2 & a5ee4a | !hlock2 & a5ee50;
assign a5fbf8 = hmaster1_p & a5fbc5 | !hmaster1_p & a5fbf7;
assign cea23a = hmaster0_p & cea234 | !hmaster0_p & cea239;
assign af34b9 = locked_p & af34b5 | !locked_p & af34b8;
assign b29d60 = hbusreq2_p & b29d5f | !hbusreq2_p & v84563c;
assign b29fc9 = hlock2_p & b29fb7 | !hlock2_p & v845660;
assign af3c2f = hlock2_p & af3c2e | !hlock2_p & af3c2d;
assign cea0b6 = hgrant1_p & deadde | !hgrant1_p & cea8a9;
assign b26782 = hmaster0_p & b26781 | !hmaster0_p & !b26763;
assign deae2e = hready_p & deae1b | !hready_p & !deae2d;
assign c3bbd2 = hmastlock_p & deada7 | !hmastlock_p & v84566c;
assign a5f2ea = hlock2_p & a5f2e9 | !hlock2_p & v84563c;
assign a5f19a = hbusreq2_p & a5f197 | !hbusreq2_p & a5f199;
assign a5fc4f = stateA1_p & v84566e | !stateA1_p & !a5fb87;
assign ab0c7a = hlock2_p & ab0c79 | !hlock2_p & c3bc3c;
assign b29b26 = hmaster1_p & b29ab6 | !hmaster1_p & b29e96;
assign c3bbfe = hbusreq2_p & c3bbfd | !hbusreq2_p & !v84565a;
assign ab0cdc = hmaster1_p & ab0bca | !hmaster1_p & ab0cdb;
assign a5f1cc = hlock2_p & a5f1cb | !hlock2_p & v84563c;
assign cea862 = decide_p & cea861 | !decide_p & v84563c;
assign a5fc3a = hbusreq2_p & a5fc39 | !hbusreq2_p & v84563c;
assign deae1c = hgrant1_p & deada8 | !hgrant1_p & deadaa;
assign b29f93 = hmaster1_p & c3bceb | !hmaster1_p & b29f92;
assign c3b6a7 = hlock1_p & c3bbd2 | !hlock1_p & deada8;
assign a5f333 = hgrant2_p & a5f332 | !hgrant2_p & a5f8f5;
assign ab0c95 = hlock0_p & v84563c | !hlock0_p & !b29aa7;
assign a5eebc = locked_p & a5eebb | !locked_p & a5f3d7;
assign a5f8e1 = stateG10_1_p & a5f8dd | !stateG10_1_p & !a5f8e0;
assign ab073f = hready_p & ab0736 | !hready_p & ab073e;
assign b29b34 = hready_p & b29b29 | !hready_p & b29b33;
assign b29f92 = hbusreq2_p & b29f91 | !hbusreq2_p & v84563c;
assign cea0e9 = hbusreq3 & v84563c | !hbusreq3 & cea86e;
assign b29977 = decide_p & b29976 | !decide_p & v84563c;
assign a5eb3a = hbusreq0 & a5eb39 | !hbusreq0 & v84563c;
assign a5f35c = hmaster1_p & a5f35b | !hmaster1_p & a5f285;
assign d40d74 = hmaster1_p & d40d73 | !hmaster1_p & v84563c;
assign a5ef39 = hlock2_p & a5ef34 | !hlock2_p & a5ef38;
assign a5f45b = hready & a5f457 | !hready & a5f45a;
assign dea6cc = hlock2_p & dea6cb | !hlock2_p & !deada8;
assign b29d00 = hready & deae1d | !hready & c3bdce;
assign a5f07d = hbusreq3 & a5f075 | !hbusreq3 & !a5f07c;
assign ab0bab = hlock0_p & v84563c | !hlock0_p & !ab0baa;
assign ab0c1b = hbusreq2_p & ab0c1a | !hbusreq2_p & v84563c;
assign a5f32f = hmaster1_p & a5f32e | !hmaster1_p & a5f887;
assign b29958 = hmaster0_p & b29934 | !hmaster0_p & !b29957;
assign a5ee2d = hlock1_p & a5fb8c | !hlock1_p & !b2982f;
assign b29f42 = hlock2 & deaca2 | !hlock2 & b29f41;
assign b29ede = hmaster1_p & v84563c | !hmaster1_p & b29edd;
assign ab0625 = decide_p & ab0624 | !decide_p & v845662;
assign ab0c15 = hlock2_p & ab0c14 | !hlock2_p & v84563c;
assign cea0c2 = hgrant2_p & cea0b5 | !hgrant2_p & cea0c1;
assign ab0c25 = hbusreq0_p & b26695 | !hbusreq0_p & !c3bcef;
assign ce9e24 = hmaster1_p & ce9e20 | !hmaster1_p & !ce9e23;
assign a5f8d1 = hlock1_p & a5f8ce | !hlock1_p & !a5f8d0;
assign a5ef9a = hlock2_p & a5ee0c | !hlock2_p & a5ef99;
assign cea466 = hmaster1_p & cea461 | !hmaster1_p & cea465;
assign ab05c0 = hlock0_p & ab05bf | !hlock0_p & ab0591;
assign ab0ad2 = hbusreq3 & ab0ad1 | !hbusreq3 & v84563c;
assign a60141 = locked_p & v84563c | !locked_p & a60140;
assign c3bc6c = hlock2_p & c3bbbc | !hlock2_p & !v84563c;
assign ce9d51 = hgrant0_p & cea85f | !hgrant0_p & ce9d50;
assign a5f51a = hbusreq1 & c3b6c4 | !hbusreq1 & !a5f493;
assign cea434 = hready & cea433 | !hready & cea40a;
assign b29a97 = hbusreq2_p & b29a96 | !hbusreq2_p & !c3bc21;
assign bdb5b4 = hgrant2_p & bdb5b2 | !hgrant2_p & bdb5b3;
assign c3b6b1 = hlock0_p & c3b6a8 | !hlock0_p & c3b6af;
assign a5fc5a = hready & a5fb89 | !hready & dead76;
assign deae6d = hmaster1_p & deae6a | !hmaster1_p & deae6c;
assign d40d48 = hmaster1_p & d40d36 | !hmaster1_p & d40d47;
assign b29f85 = hready_p & b29ee1 | !hready_p & b29f84;
assign a5f535 = hbusreq1 & a5f534 | !hbusreq1 & a5f493;
assign ab05bd = hlock0_p & v845660 | !hlock0_p & !cea38d;
assign a5f7c2 = hready & a5fb12 | !hready & !deacb7;
assign a5f2d4 = hbusreq0 & a5f2d2 | !hbusreq0 & a5f2d3;
assign ab0cb5 = hgrant2_p & ab0bba | !hgrant2_p & ab0c9f;
assign a5f1fc = hgrant2_p & v84563c | !hgrant2_p & a5f1fb;
assign a5f58b = hmaster0_p & a5f47c | !hmaster0_p & a5f58a;
assign a5f069 = hlock0_p & a5f6ea | !hlock0_p & a5f067;
assign a5eea7 = hlock0_p & a5eea6 | !hlock0_p & !a5ee5f;
assign a5faae = hgrant1_p & a60196 | !hgrant1_p & a5faad;
assign cea3ac = hmaster1_p & cea3a8 | !hmaster1_p & cea3ab;
assign a60199 = hlock0_p & a60198 | !hlock0_p & a6018c;
assign b266db = hgrant1_p & b266da | !hgrant1_p & b26696;
assign a81cd0 = hlock1_p & a81ca9 | !hlock1_p & v84563c;
assign af353f = stateG10_1_p & v84563c | !stateG10_1_p & af352c;
assign a5ef29 = hbusreq2 & a5ef0b | !hbusreq2 & a5ef13;
assign cea38d = hready & deae67 | !hready & !deae59;
assign ab067d = hmaster1_p & ab067c | !hmaster1_p & ab0ace;
assign dea6f7 = hlock3_p & dea6f2 | !hlock3_p & dea6f6;
assign dea6d3 = hbusreq3 & dea6cd | !hbusreq3 & dea6d2;
assign deae3e = decide_p & deae3d | !decide_p & v84563c;
assign c3b724 = hbusreq2_p & c3b717 | !hbusreq2_p & c3b716;
assign stateG3_0 = !adaf1c;
assign cea89c = hlock0_p & c98b96 | !hlock0_p & deacaa;
assign dea752 = hgrant2_p & deade2 | !hgrant2_p & dea751;
assign b26746 = hmaster0_p & b26742 | !hmaster0_p & b26745;
assign b29916 = hgrant1_p & b29915 | !hgrant1_p & b29914;
assign c3bbd6 = hbusreq2_p & c3bbd5 | !hbusreq2_p & !c3bbd3;
assign a81cf3 = hlock0_p & a81cc8 | !hlock0_p & a81cf2;
assign a5f8b6 = hgrant1_p & deac52 | !hgrant1_p & a5f8b5;
assign cea392 = hbusreq3 & cea390 | !hbusreq3 & cea391;
assign a5ef8b = hlock0_p & a5edda | !hlock0_p & a5f36e;
assign a5ea3b = hbusreq2_p & a5ea3a | !hbusreq2_p & a5ea39;
assign dea6d4 = hbusreq2_p & dea6cc | !hbusreq2_p & dea6cb;
assign a5f1de = hlock0_p & a5f1dd | !hlock0_p & v84563c;
assign b299ce = hbusreq2_p & b299cd | !hbusreq2_p & !b29948;
assign b266ca = hmastlock_p & b26692 | !hmastlock_p & v84566c;
assign cea0f1 = hmaster0_p & cea0e8 | !hmaster0_p & cea0f0;
assign ab0c99 = hlock0_p & v84563c | !hlock0_p & !ab0c98;
assign a5f982 = hlock1_p & a5f980 | !hlock1_p & a5f981;
assign a5fc75 = hburst0_p & d615cf | !hburst0_p & a5fc74;
assign a5ea93 = hgrant2_p & a5ea91 | !hgrant2_p & a5ea92;
assign a5fb93 = hlock0_p & a5fb90 | !hlock0_p & a5fb92;
assign v97045b = hready_p & v97044e | !hready_p & v97045a;
assign a5ea46 = hbusreq2 & a5ea42 | !hbusreq2 & a5ea45;
assign ab0b53 = hlock2_p & ab0b52 | !hlock2_p & dead2e;
assign ab0561 = hlock0_p & v84563c | !hlock0_p & !b29942;
assign a5eeb4 = hgrant0_p & a5ee93 | !hgrant0_p & a5eeb3;
assign a5ea4a = hgrant2_p & a5ea3f | !hgrant2_p & a5ea49;
assign a5ede7 = hbusreq1 & a5ede6 | !hbusreq1 & v84563c;
assign a5fc2e = hlock2 & a5fc27 | !hlock2 & a5fc2d;
assign c3b7d0 = hlock0_p & c3bd3e | !hlock0_p & deadc4;
assign a5f39b = hbusreq3 & a5f39a | !hbusreq3 & a5fbc0;
assign b29f6c = hgrant2_p & b29f6a | !hgrant2_p & b29f6b;
assign a9b9e2 = hmaster1_p & v84563c | !hmaster1_p & !a9b9d0;
assign ab0515 = hlock0_p & v84563c | !hlock0_p & b298a4;
assign a5f8fd = hbusreq1_p & v84563c | !hbusreq1_p & v84566c;
assign c3bc16 = hlock0_p & c3bbd2 | !hlock0_p & deac86;
assign a5f9a5 = hready & v84563c | !hready & !dead0a;
assign stateG2 = !v97045d;
assign cea43e = hmaster1_p & cea438 | !hmaster1_p & cea43d;
assign b266f0 = hlock0_p & b266ef | !hlock0_p & b266a0;
assign a5f542 = hlock2 & a5f53e | !hlock2 & a5f541;
assign ab0c33 = hlock2 & v84563c | !hlock2 & ab0c32;
assign a5ea6f = hgrant0_p & a60144 | !hgrant0_p & a5ea6e;
assign a5f41d = hbusreq1 & a5f41b | !hbusreq1 & a5f41c;
assign a5fcb0 = hbusreq2 & a5fc7a | !hbusreq2 & !a5fc89;
assign a5efa8 = hlock2 & a5efa6 | !hlock2 & a5efa7;
assign cea2e8 = hready & cea2e7 | !hready & cea151;
assign a5ee5b = hbusreq1 & a5ee5a | !hbusreq1 & v84563c;
assign a5ea18 = hbusreq2_p & a5ea17 | !hbusreq2_p & a5f198;
assign dead38 = hmaster0_p & dead30 | !hmaster0_p & dead37;
assign a5f496 = hlock0_p & a5f48a | !hlock0_p & a5f495;
assign c3b887 = hmaster0_p & c3b886 | !hmaster0_p & c3b7fe;
assign hgrant3 = dea7b5;
assign c3b7e5 = hlock2_p & c3b7bd | !hlock2_p & !c3b7e4;
assign a5efe0 = hbusreq2 & a5efdf | !hbusreq2 & a5efd8;
assign c3b891 = hbusreq2_p & c3b80b | !hbusreq2_p & c3b890;
assign b0c0fd = hready_p & v84563c | !hready_p & v845658;
assign dead86 = hmaster1_p & dead83 | !hmaster1_p & dead85;
assign a5f14e = hbusreq2_p & a5f14d | !hbusreq2_p & a5f14c;
assign af3c5b = hbusreq2_p & af3c5a | !hbusreq2_p & af3c59;
assign ab0b63 = hready & b29d77 | !hready & c3bd8a;
assign a5f96f = hready & a5fc78 | !hready & a5fb8e;
assign a5f00d = hgrant2_p & a5f00c | !hgrant2_p & v84563c;
assign a5fa66 = hready & a60187 | !hready & a5fa1c;
assign a5fd11 = hbusreq0_p & v845660 | !hbusreq0_p & a5fcef;
assign b29cd8 = hbusreq2_p & b29cd4 | !hbusreq2_p & v84563c;
assign b299a9 = decide_p & b299a8 | !decide_p & b29e57;
assign a5ee8a = hlock1_p & a5fba6 | !hlock1_p & !a5ee1b;
assign a5ea89 = hbusreq0 & a5ea88 | !hbusreq0 & a5fbc1;
assign bdb582 = hlock3_p & v845660 | !hlock3_p & bdb581;
assign b2a004 = hlock2_p & b2a003 | !hlock2_p & v845660;
assign a5f4fc = hready & v84563c | !hready & a5f4fb;
assign a5f458 = hgrant1_p & a5f43a | !hgrant1_p & a5f439;
assign af34cd = hgrant0_p & af34ab | !hgrant0_p & af34cc;
assign a5edd4 = hready & a5f520 | !hready & a5f40a;
assign a5fbc1 = hlock0_p & a5fbc0 | !hlock0_p & v84563c;
assign ab051a = hlock0_p & b298a4 | !hlock0_p & ab0519;
assign b29a8c = hlock2_p & v84563c | !hlock2_p & !b29ce7;
assign b29a46 = hmaster1_p & b29a45 | !hmaster1_p & b29c3d;
assign b29f57 = hready & deaca1 | !hready & !v84565a;
assign a5f989 = hbusreq1_p & a5f988 | !hbusreq1_p & a5fc84;
assign a5f969 = hready & a5f6e4 | !hready & a5fb8e;
assign a5f2e7 = locked_p & v84563c | !locked_p & a5f2e6;
assign b29ff3 = hbusreq2_p & b29f62 | !hbusreq2_p & !v845644;
assign ab0b68 = hlock2_p & ab0b66 | !hlock2_p & !ab0b67;
assign a5fb6c = hlock0_p & a5fb6b | !hlock0_p & v84563c;
assign a5edd0 = hbusreq2 & a5edce | !hbusreq2 & a5edcf;
assign a5edcd = hlock0_p & a5edcc | !hlock0_p & a5f4fc;
assign a5f2fd = hgrant0_p & a5f2ed | !hgrant0_p & a5f2fc;
assign a5f1ec = hmaster0_p & a5f1ce | !hmaster0_p & a5f1eb;
assign b29f9c = hready & c3bdbd | !hready & !dead40;
assign a5ef30 = hgrant0_p & a5ef18 | !hgrant0_p & a5ef2f;
assign cea180 = hlock3_p & cea177 | !hlock3_p & cea17f;
assign ab0ca2 = hbusreq2_p & ab0c15 | !hbusreq2_p & cea15a;
assign busreq = b840b3;
assign a5f99d = hbusreq2_p & a5f99c | !hbusreq2_p & v84563c;
assign adaedb = hready_p & adaec1 | !hready_p & adaeda;
assign a5eead = hlock2 & a5f3b9 | !hlock2 & a5eeac;
assign a5ead1 = hbusreq0_p & a5fa8a | !hbusreq0_p & a5f233;
assign a5f6de = hmaster1_p & a5f6db | !hmaster1_p & a5f6dd;
assign ce9db9 = hmaster1_p & ce9db6 | !hmaster1_p & ce9db8;
assign cea277 = hbusreq2_p & cea276 | !hbusreq2_p & v84563c;
assign a5edb9 = hlock0_p & a5edb8 | !hlock0_p & a5f4ea;
assign a5fb2f = hbusreq3 & a5fb23 | !hbusreq3 & a5fb2e;
assign c3b731 = hlock0_p & c3b648 | !hlock0_p & c3b730;
assign a5f23b = hlock2_p & a5f235 | !hlock2_p & a5f23a;
assign a5f91a = hlock0_p & a5f919 | !hlock0_p & a5f86c;
assign a5fc64 = hmaster1_p & a5fc63 | !hmaster1_p & v84563c;
assign ab06b4 = hlock2_p & ab06b3 | !hlock2_p & b29a7b;
assign cea18f = hlock0_p & v84563c | !hlock0_p & cea18e;
assign b2998f = hlock2_p & b2998b | !hlock2_p & b2998e;
assign dea6c6 = hgrant0_p & dea6be | !hgrant0_p & dea6c5;
assign af3534 = hmaster1_p & af3531 | !hmaster1_p & af3533;
assign a5ee3d = hlock2 & a5f36b | !hlock2 & a5ee38;
assign b29eae = locked_p & b29ead | !locked_p & !v84563c;
assign cea3a2 = hbusreq3 & cea39b | !hbusreq3 & cea3a1;
assign adaeee = hmaster1_p & v84563c | !hmaster1_p & adaeed;
assign ab054b = hready & ab054a | !hready & v84563c;
assign c3bd37 = hmastlock_p & c3bd36 | !hmastlock_p & !v84563c;
assign a5eef1 = hlock2_p & a5eeea | !hlock2_p & !a5eef0;
assign a5ee76 = hbusreq0_p & v845641 | !hbusreq0_p & a5ee26;
assign bdb59b = decide_p & bdb597 | !decide_p & bdb59a;
assign ab05ca = hlock0_p & v84563c | !hlock0_p & !ab05a4;
assign cea17a = locked_p & cea179 | !locked_p & v84563c;
assign cea19d = hbusreq2_p & cea198 | !hbusreq2_p & cea197;
assign aa0e0a = jx1_p & af3c47 | !jx1_p & af3510;
assign ab059e = hbusreq2_p & ab059d | !hbusreq2_p & ab059c;
assign b29e51 = hbusreq3 & b29e50 | !hbusreq3 & !v845660;
assign a5ee83 = locked_p & v84563c | !locked_p & a5f3b4;
assign a5ee2b = hbusreq1 & a5ee2a | !hbusreq1 & v84563c;
assign af355e = hbusreq2_p & af3558 | !hbusreq2_p & af3541;
assign a5ee58 = hready & a5ee54 | !hready & a5ee57;
assign a5f476 = hbusreq2_p & a5f475 | !hbusreq2_p & !a5f474;
assign a5f548 = hlock0_p & a5fa6c | !hlock0_p & a5f4fc;
assign b29b1f = hlock2_p & v845660 | !hlock2_p & !b29b1e;
assign a5f925 = hlock2_p & a5f924 | !hlock2_p & a5f883;
assign ab063a = hmaster0_p & ab0631 | !hmaster0_p & ab0639;
assign dea724 = hlock0_p & dead71 | !hlock0_p & !dead77;
assign ab0613 = hlock2 & ab0529 | !hlock2 & ab0612;
assign b29fa4 = hbusreq2_p & b29fa3 | !hbusreq2_p & v84563c;
assign a5eb53 = hmaster0_p & a5eb52 | !hmaster0_p & !a5f0af;
assign a5ea80 = hlock2 & a5ea7c | !hlock2 & a5ea7f;
assign cea2f0 = hgrant2_p & cea159 | !hgrant2_p & !cea2ef;
assign deac53 = hbusreq1_p & deac52 | !hbusreq1_p & v84565a;
assign c3bd51 = hmaster1_p & c3bd46 | !hmaster1_p & c3bd50;
assign deac4c = hburst0_p & v8c6449 | !hburst0_p & deac4b;
assign c3bdb1 = hlock0_p & c3bdb0 | !hlock0_p & !c3bd8e;
assign a5ee4a = hlock0_p & a5ee45 | !hlock0_p & a5ee49;
assign c3b81a = hlock2_p & c3b7a5 | !hlock2_p & !c3b7b0;
assign a5f250 = hlock2 & a5f24c | !hlock2 & a5f24f;
assign a5ee37 = hlock0_p & a60140 | !hlock0_p & a5f36b;
assign ab0745 = hbusreq0_p & dead41 | !hbusreq0_p & !cea18d;
assign b29b10 = hmaster1_p & b29a54 | !hmaster1_p & b29e5c;
assign a5eb91 = hbusreq2_p & a5eb90 | !hbusreq2_p & a5eb8f;
assign cea415 = hlock2_p & cea413 | !hlock2_p & cea414;
assign b29d89 = hlock0_p & b29d88 | !hlock0_p & !v84563c;
assign dea6f0 = hbusreq3_p & dea6dd | !hbusreq3_p & dea6ef;
assign a5ee30 = locked_p & a5ee2f | !locked_p & v845641;
assign a5fc45 = hlock0_p & a5fc44 | !hlock0_p & v84563c;
assign a9b9d4 = decide_p & a9b9d3 | !decide_p & a9b9d2;
assign ab0c03 = hlock0_p & v84563c | !hlock0_p & !c3bce0;
assign c3b76d = hmaster1_p & c3b76c | !hmaster1_p & c3bccf;
assign c3bd6d = hbusreq3 & c3bd6a | !hbusreq3 & c3bd6c;
assign dea7a6 = decide_p & dea7a3 | !decide_p & v84563c;
assign a5eb43 = hgrant2_p & a5eb42 | !hgrant2_p & a5ea2c;
assign a5ee42 = hmaster1_p & a5ee41 | !hmaster1_p & a5fbc5;
assign a5edc9 = hlock0_p & a5edc8 | !hlock0_p & a5f536;
assign a5efd9 = hbusreq2_p & a5efd3 | !hbusreq2_p & a5efd8;
assign af3c36 = hmaster1_p & af3c35 | !hmaster1_p & !v84563c;
assign a5f93e = hready & a60192 | !hready & a5f8d2;
assign af34dd = hbusreq2_p & af34dc | !hbusreq2_p & af3c4c;
assign a5ebe6 = hbusreq0 & a5ea2a | !hbusreq0 & v84563c;
assign ab0b79 = locked_p & v84563c | !locked_p & !b29d66;
assign ab0585 = hlock3_p & ab0578 | !hlock3_p & ab0584;
assign a5fc86 = start_p & a5fba3 | !start_p & a5fc85;
assign cea151 = hlock1_p & v84563c | !hlock1_p & cea150;
assign ab0b7f = hbusreq2_p & ab0b7b | !hbusreq2_p & ab0b7e;
assign a5fc62 = hbusreq3 & a5fc61 | !hbusreq3 & v84563c;
assign a5fd18 = hmaster0_p & a5fd03 | !hmaster0_p & a5fd17;
assign a5ef84 = hbusreq2 & a5ef82 | !hbusreq2 & a5ef83;
assign a5f571 = hlock1_p & a60177 | !hlock1_p & !a5f570;
assign c3b74b = decide_p & c3b74a | !decide_p & !v845660;
assign a5f728 = locked_p & v84563c | !locked_p & a5f727;
assign c3bd14 = hgrant1_p & c3bd12 | !hgrant1_p & c3bd13;
assign deacb6 = hgrant1_p & deacb5 | !hgrant1_p & deaca1;
assign af34d5 = hlock2_p & af3c58 | !hlock2_p & af3c4c;
assign ab0646 = hgrant2_p & ab0644 | !hgrant2_p & ab0645;
assign a5e9ea = hgrant2_p & a5e9e6 | !hgrant2_p & a5e9e9;
assign a5fccb = locked_p & v84563c | !locked_p & c3bd5f;
assign c3bc0d = hlock0_p & c3bbe2 | !hlock0_p & !v84563c;
assign ab0c9b = locked_p & ab0c9a | !locked_p & !v84563c;
assign b29ea0 = hmaster0_p & b29e9c | !hmaster0_p & !b29e9f;
assign dea7a9 = hmaster1_p & dea758 | !hmaster1_p & !dead65;
assign a5f55a = hready & a5f520 | !hready & a5f559;
assign af34b0 = hlock2_p & af34af | !hlock2_p & af3c5e;
assign c3bde5 = hbusreq2_p & c3bde4 | !hbusreq2_p & v84563c;
assign b29957 = hmaster1_p & b29955 | !hmaster1_p & !b29956;
assign c3bc02 = hlock1_p & v84563c | !hlock1_p & v84565a;
assign cea2ac = hlock1_p & deada8 | !hlock1_p & !deac56;
assign a5f3a5 = hbusreq2 & a5f3a1 | !hbusreq2 & a5f3a4;
assign a5f302 = hgrant2_p & v84563c | !hgrant2_p & a5f2ff;
assign ce9cb6 = hmaster1_p & ce9cb5 | !hmaster1_p & cea85f;
assign a5fc69 = hmastlock_p & a5fc68 | !hmastlock_p & v84563c;
assign ce9d41 = hlock3_p & ce9d2f | !hlock3_p & ce9d40;
assign cea358 = hbusreq2_p & cea343 | !hbusreq2_p & cea85d;
assign ab058b = hbusreq2_p & ab058a | !hbusreq2_p & ab0588;
assign b29ea6 = locked_p & b29ea5 | !locked_p & !c3bc47;
assign a5f4d1 = hready & a5f4cb | !hready & a5f4d0;
assign c3bc7e = hbusreq2_p & c3bc7d | !hbusreq2_p & c3bc7c;
assign a5f320 = hready & v84563c | !hready & !deac7a;
assign b29fcf = hlock3_p & b29faa | !hlock3_p & b29fce;
assign cea8a4 = hmaster1_p & cea879 | !hmaster1_p & !cea8a3;
assign b29cb9 = hlock3_p & b29c3d | !hlock3_p & v84563c;
assign ab0683 = hlock0_p & c3bcdb | !hlock0_p & !v84563c;
assign a5f4eb = hlock0_p & a5f4d1 | !hlock0_p & !a5f4ea;
assign a5ea65 = hbusreq2 & a5ea64 | !hbusreq2 & a5fbc1;
assign bdb59e = hmaster0_p & dead2e | !hmaster0_p & bdb59d;
assign b29f69 = hlock2_p & b29f3d | !hlock2_p & !b29f42;
assign af35a5 = decide_p & af35a4 | !decide_p & af3535;
assign ab0c16 = hbusreq2_p & ab0c15 | !hbusreq2_p & ab0acb;
assign a81cb4 = hlock1_p & a81cb1 | !hlock1_p & a81cb3;
assign a5eaa4 = decide_p & a5ea8e | !decide_p & a5eaa3;
assign a5fcf9 = hbusreq1_p & a5fcdd | !hbusreq1_p & a5fce3;
assign adaed1 = hlock0_p & adaec4 | !hlock0_p & v84563c;
assign b29a90 = hbusreq3 & b29a8d | !hbusreq3 & b29a8f;
assign b2990c = hbusreq2_p & b2990b | !hbusreq2_p & v84563c;
assign c3b660 = hmastlock_p & c3bd10 | !hmastlock_p & v84563c;
assign cea174 = hgrant2_p & cea15e | !hgrant2_p & !cea173;
assign a5fbfc = locked_p & a5fbfb | !locked_p & v84563c;
assign b0d8fd = hbusreq3_p & v84563c | !hbusreq3_p & v845668;
assign a5fb7f = hmaster1_p & a5fb6e | !hmaster1_p & a5fb7e;
assign b29f8f = hlock0_p & b29eac | !hlock0_p & v84563c;
assign b29fe2 = hbusreq3 & b29fd6 | !hbusreq3 & b29fe1;
assign dead6c = stateA1_p & v84563c | !stateA1_p & !c07311;
assign b266f1 = hbusreq2_p & b266e7 | !hbusreq2_p & !b266f0;
assign a5fb61 = hbusreq3 & a5fb54 | !hbusreq3 & a5fb60;
assign a5fc54 = hbusreq1 & v84563c | !hbusreq1 & v970413;
assign c3b6d5 = hready_p & c3b65b | !hready_p & c3b6d4;
assign a5ee61 = hbusreq2 & a5ee51 | !hbusreq2 & !a5ee60;
assign c3bca7 = hmaster1_p & c3bca4 | !hmaster1_p & c3bca6;
assign ab0c6f = hbusreq3 & ab0c6c | !hbusreq3 & ab0c6e;
assign ab062d = hlock0_p & ab0adc | !hlock0_p & !ab05f0;
assign ab0bfb = locked_p & ab0bfa | !locked_p & b26695;
assign c3b756 = hgrant0_p & c3b750 | !hgrant0_p & c3b755;
assign c3b729 = hmaster0_p & c3b728 | !hmaster0_p & c3b6b6;
assign cea32b = hmaster1_p & cea178 | !hmaster1_p & cea31e;
assign a5e9c7 = hbusreq2 & a5e9be | !hbusreq2 & !a5e9c6;
assign c3bc62 = hready & cea151 | !hready & c3bc61;
assign ab0bc9 = hgrant3_p & ab0b51 | !hgrant3_p & !ab0bc8;
assign b29fb3 = hlock1_p & v84563c | !hlock1_p & b29fb2;
assign b299ea = hgrant3_p & b299d6 | !hgrant3_p & b299e9;
assign ab0522 = hlock0_p & b298a4 | !hlock0_p & !b298ae;
assign adaebb = start_p & v84563c | !start_p & adaeba;
assign v970440 = hbusreq0_p & v9703fd | !hbusreq0_p & v97043f;
assign a5ea5c = hlock0_p & a5ea5a | !hlock0_p & !a5ea5b;
assign ab05af = locked_p & v84563c | !locked_p & b29992;
assign a5eb86 = hbusreq3 & a5eb84 | !hbusreq3 & a5eb85;
assign a5f4a6 = hbusreq1 & a5f4a5 | !hbusreq1 & v84563c;
assign a5f1d6 = hready & v84563c | !hready & !a5fb8c;
assign a5eec0 = hbusreq1 & a5eebf | !hbusreq1 & !v84563c;
assign deaded = hlock1_p & deadde | !hlock1_p & !deadec;
assign ce9cf9 = hmaster1_p & ce9cf7 | !hmaster1_p & ce9cf8;
assign c3b883 = hlock0_p & c3bd4b | !hlock0_p & ce9dc7;
assign b29f37 = hbusreq2_p & b29efd | !hbusreq2_p & v84563c;
assign a5f1ed = hgrant2_p & v84563c | !hgrant2_p & a5f734;
assign a5f99b = hlock0_p & a5fb6b | !hlock0_p & a5f726;
assign ab0531 = hmaster1_p & ab052e | !hmaster1_p & ab0530;
assign a5ebc2 = hbusreq2_p & a5ebc1 | !hbusreq2_p & a5f199;
assign a5f971 = hlock0_p & a5f970 | !hlock0_p & a5fc2c;
assign ab06c9 = hlock1_p & deac52 | !hlock1_p & ab06c8;
assign c3b713 = hgrant1_p & c3b712 | !hgrant1_p & deae74;
assign c3bc4d = locked_p & v84563c | !locked_p & !deace1;
assign af3495 = hmaster0_p & af3491 | !hmaster0_p & af3494;
assign a5f97e = stateA1_p & a5fb9d | !stateA1_p & a5f97d;
assign a5f070 = hbusreq0_p & v84563c | !hbusreq0_p & a5f6fa;
assign adaee5 = hgrant2_p & adaee4 | !hgrant2_p & v84563c;
assign a5f54a = hlock2 & a5f548 | !hlock2 & a5f549;
assign c3bcf5 = hbusreq3 & c3bcf4 | !hbusreq3 & c3bceb;
assign cea43c = hbusreq2_p & cea43a | !hbusreq2_p & cea439;
assign a5f724 = hmaster1_p & a5f71b | !hmaster1_p & a5f723;
assign deadd2 = hlock2_p & deadd1 | !hlock2_p & !v84563c;
assign b29d55 = hbusreq2_p & b29d54 | !hbusreq2_p & v84563c;
assign d40d4f = hgrant1_p & d40d33 | !hgrant1_p & d40d3c;
assign b29a4c = hbusreq3 & b29a49 | !hbusreq3 & b29a4b;
assign d40d8e = hmaster1_p & d40d68 | !hmaster1_p & v84563c;
assign adaefe = start_p & a81ca6 | !start_p & !v845670;
assign c3b824 = hready & c3bdae | !hready & deae02;
assign d40d52 = hbusreq2_p & d40d31 | !hbusreq2_p & d40d51;
assign deac52 = hmastlock_p & v84563c | !hmastlock_p & v84566c;
assign b29d17 = hlock2_p & v84563c | !hlock2_p & v84565a;
assign a5ee6a = hbusreq2_p & a5ee64 | !hbusreq2_p & a5ee69;
assign deaca1 = hmastlock_p & deaca0 | !hmastlock_p & v84563c;
assign af34c6 = hbusreq2_p & af34c5 | !hbusreq2_p & af3c4c;
assign a5f6d2 = hlock2_p & a5fa6d | !hlock2_p & v84563c;
assign a5f6ed = locked_p & a5f6ec | !locked_p & v845641;
assign dea74b = hbusreq2_p & deadd2 | !hbusreq2_p & !v84563c;
assign cea46a = hgrant2_p & cea469 | !hgrant2_p & !v845660;
assign ab061b = hbusreq2_p & ab05a9 | !hbusreq2_p & ab061a;
assign a5f8c4 = hready & v84563c | !hready & a5f8c3;
assign c3b67b = hlock1_p & v84563c | !hlock1_p & !c3b67a;
assign a5f833 = start_p & v845654 | !start_p & !c06d34;
assign b29eca = hbusreq3 & b29ec9 | !hbusreq3 & dead84;
assign a5fab2 = hready & a60193 | !hready & a60196;
assign b29cff = hlock0_p & b29cfd | !hlock0_p & !b29cfe;
assign deae74 = hbusreq1_p & deada8 | !hbusreq1_p & !v84563c;
assign ab0607 = hlock0_p & ab0590 | !hlock0_p & ab0606;
assign bdb595 = hmaster1_p & bdb58d | !hmaster1_p & v84565a;
assign c3bd7d = hbusreq2_p & c3bd7c | !hbusreq2_p & !c3bc21;
assign cea487 = hbusreq2_p & cea47d | !hbusreq2_p & cea47c;
assign a5fbb7 = hready & a5fbb6 | !hready & !a5fbae;
assign ab0b3d = hbusreq3 & v84563c | !hbusreq3 & ab0b3c;
assign a5ee68 = locked_p & v84563c | !locked_p & a5ee26;
assign af34e3 = hmaster1_p & af3c5e | !hmaster1_p & af3c58;
assign cea3ed = hbusreq2_p & cea3ec | !hbusreq2_p & cea3ea;
assign ab0c84 = hbusreq2_p & ab0c83 | !hbusreq2_p & ab0b5f;
assign ab0ba1 = hbusreq0_p & b266a8 | !hbusreq0_p & ab0b96;
assign ab0b97 = hlock0_p & v84563c | !hlock0_p & ab0b96;
assign cea346 = hmaster1_p & cea345 | !hmaster1_p & cea238;
assign a5f950 = hmaster0_p & a5f927 | !hmaster0_p & a5f94f;
assign deacac = hlock2_p & deacab | !hlock2_p & v84563c;
assign b26744 = hbusreq2_p & b2670b | !hbusreq2_p & b26743;
assign b29ac7 = decide_p & b29ac6 | !decide_p & b29e57;
assign af358b = hgrant2_p & af352f | !hgrant2_p & af352d;
assign c3b85b = hmaster0_p & c3b852 | !hmaster0_p & c3b7ed;
assign b2992b = hready & b29926 | !hready & b2992a;
assign ab0c69 = hlock0_p & v84563c | !hlock0_p & !c3bd5f;
assign dead78 = hlock2_p & dead73 | !hlock2_p & !dead77;
assign a5eeb2 = hmaster1_p & a5eeab | !hmaster1_p & a5eeb1;
assign a5f6d9 = hgrant2_p & a5f9c5 | !hgrant2_p & a5f9c8;
assign a5f956 = hbusreq3 & a5f953 | !hbusreq3 & !a5f955;
assign b29f08 = start_p & cea1aa | !start_p & !b29f07;
assign cea2f9 = hgrant0_p & cea2ee | !hgrant0_p & cea2f8;
assign a5f74f = hbusreq3 & a5f74c | !hbusreq3 & !a5f74e;
assign a5ea16 = hbusreq2 & a5ea14 | !hbusreq2 & a5ea15;
assign c3bc48 = locked_p & v84563c | !locked_p & c3bc47;
assign cea31e = hgrant2_p & v84563c | !hgrant2_p & !cea31d;
assign a5ee1e = hbusreq1_p & v9703fc | !hbusreq1_p & !dead7b;
assign a5f06a = locked_p & a5fb97 | !locked_p & v845641;
assign a5ebc7 = hbusreq2_p & a5ebc1 | !hbusreq2_p & a5e9c9;
assign a5f366 = hready & a5f365 | !hready & a5fbd9;
assign a5f18a = hbusreq1_p & a5fa1c | !hbusreq1_p & !a60177;
assign ab0577 = hmaster1_p & ab056e | !hmaster1_p & !ab0576;
assign b29aa4 = hlock2 & b29a4d | !hlock2 & b29aa3;
assign a5f798 = hready & a5f9f6 | !hready & a5f797;
assign deae8e = hmaster1_p & deae8d | !hmaster1_p & !v84563c;
assign a57858 = hready_p & v84563c | !hready_p & v845656;
assign ab0be6 = hmaster1_p & ab0be3 | !hmaster1_p & ab0be5;
assign a5fbbc = hbusreq0 & a5fb9c | !hbusreq0 & !a5fbbb;
assign c3bc55 = hbusreq2_p & c3bc54 | !hbusreq2_p & c3bc53;
assign b29f78 = hlock1_p & deac52 | !hlock1_p & b29f77;
assign cea235 = hlock0_p & b26697 | !hlock0_p & v84563c;
assign af35c0 = hready_p & af35b3 | !hready_p & af35bf;
assign d40d59 = hgrant2_p & d40d4e | !hgrant2_p & d40d58;
assign c3bc98 = hlock0_p & b266a8 | !hlock0_p & c3bc90;
assign deace8 = hmaster1_p & v84563c | !hmaster1_p & deace7;
assign a5ef48 = decide_p & a5ef44 | !decide_p & !a5ef47;
assign b29fac = hlock2_p & b29fab | !hlock2_p & dead2e;
assign a5f03f = hbusreq0 & a5f6dc | !hbusreq0 & a5f03e;
assign a5fb20 = hready & a5fb1d | !hready & a5fb1f;
assign deae40 = hbusreq2_p & deadd7 | !hbusreq2_p & !v84563c;
assign deace4 = hlock0_p & deace3 | !hlock0_p & deace1;
assign a5fcbd = hbusreq2 & a5fcbc | !hbusreq2 & v845660;
assign cea2b4 = hmaster0_p & cea2b2 | !hmaster0_p & cea2b3;
assign a5f9ca = hgrant2_p & a5f9c6 | !hgrant2_p & a5f9c9;
assign ab073a = hgrant2_p & ab06a3 | !hgrant2_p & ab0739;
assign c3b63b = hlock0_p & c3b639 | !hlock0_p & c3b63a;
assign dea784 = hbusreq2_p & deae24 | !hbusreq2_p & !deadba;
assign a5fc1a = hready & a5fb71 | !hready & !v84563c;
assign b29fcc = hmaster1_p & b29fc8 | !hmaster1_p & b29fcb;
assign a5f079 = hbusreq0_p & a5f70c | !hbusreq0_p & v84563c;
assign a5eeab = hgrant2_p & a5eeaa | !hgrant2_p & v84563c;
assign b29931 = hbusreq2_p & b2992d | !hbusreq2_p & v84563c;
assign a5f719 = hlock2_p & a5f70e | !hlock2_p & !a5f718;
assign dea6e0 = hlock2_p & dea6df | !hlock2_p & !v84563c;
assign a5f7a3 = hlock0_p & a5f798 | !hlock0_p & a5f7a2;
assign a5f172 = hlock0_p & a5f16f | !hlock0_p & a5f171;
assign cea160 = hready & dead0a | !hready & !b266da;
assign ab0549 = hgrant1_p & ab0548 | !hgrant1_p & v84563c;
assign af3c4d = hbusreq1_p & af3c4c | !hbusreq1_p & d40d33;
assign ce9dba = hmaster0_p & ce9db9 | !hmaster0_p & ce9d13;
assign d40d2b = hmastlock_p & d40d2a | !hmastlock_p & v84563c;
assign a5f3f4 = hbusreq1_p & v84563c | !hbusreq1_p & !ab0aeb;
assign cea2a7 = hbusreq2_p & cea2a6 | !hbusreq2_p & v84563c;
assign af3589 = hmaster1_p & af3531 | !hmaster1_p & af352d;
assign a5eb9c = hbusreq2 & a5f0ac | !hbusreq2 & a5ea8f;
assign b29948 = hlock0_p & b29947 | !hlock0_p & !v84563c;
assign ce9def = hbusreq2_p & cea35c | !hbusreq2_p & cea35b;
assign c3bc8e = hbusreq3 & c3bc8d | !hbusreq3 & c3bc70;
assign a5e9d2 = hbusreq2_p & a5f195 | !hbusreq2_p & a5f196;
assign deae5b = locked_p & deae59 | !locked_p & deae5a;
assign v9269ad = hmaster0_p & v845658 | !hmaster0_p & !v84563c;
assign deade0 = hlock0_p & deaddf | !hlock0_p & !v84563c;
assign b29aac = hmaster1_p & b29aa2 | !hmaster1_p & b29aab;
assign c3bbf3 = hbusreq3 & c3bbf1 | !hbusreq3 & c3bbf2;
assign a60171 = hbusreq1 & a60169 | !hbusreq1 & !a60170;
assign af3562 = hlock1_p & v84563c | !hlock1_p & af3561;
assign ab0629 = hbusreq2_p & ab0628 | !hbusreq2_p & ab05f1;
assign a5fb83 = hlock0_p & a5fb82 | !hlock0_p & a5fb71;
assign b29d80 = hlock2 & b29d7c | !hlock2 & b29d7f;
assign hgrant1 = !ce9e60;
assign ab05d0 = hlock2 & ab051b | !hlock2 & ab05cf;
assign dead9b = hbusreq2_p & dead9a | !hbusreq2_p & v84563c;
assign a5eb98 = hgrant2_p & a5eb92 | !hgrant2_p & a5eb97;
assign deacc3 = hbusreq3 & deacc1 | !hbusreq3 & !deacc2;
assign v845674 = stateG3_2_p & v84563c | !stateG3_2_p & !v84563c;
assign a5f0c3 = hready & a5f9f6 | !hready & a5f786;
assign deace1 = hlock1_p & b26695 | !hlock1_p & deace0;
assign b29d6e = hready & dead0c | !hready & b2672b;
assign a5fcf6 = hbusreq1 & a5fcf3 | !hbusreq1 & !a5fcf5;
assign ab056c = hlock2 & ab056a | !hlock2 & ab056b;
assign b29e4c = hready & dead76 | !hready & v84563c;
assign a81cf7 = hlock1_p & a81cb1 | !hlock1_p & a81cf6;
assign deadbc = hbusreq1_p & deadba | !hbusreq1_p & !v84565a;
assign cea8ac = hlock0_p & cea8ab | !hlock0_p & v84563c;
assign a5f86b = hbusreq1 & deac5b | !hbusreq1 & a5f86a;
assign deadb2 = hlock1_p & deada8 | !hlock1_p & deadb1;
assign b29d5d = locked_p & b29d5c | !locked_p & b26695;
assign c3b849 = hlock0_p & c3bdd5 | !hlock0_p & !deadba;
assign b2675b = hmaster0_p & b26755 | !hmaster0_p & b2675a;
assign b266d6 = hgrant2_p & b266d4 | !hgrant2_p & b266d5;
assign a5fd24 = hlock0_p & a5fd23 | !hlock0_p & v84563c;
assign ab05d7 = decide_p & ab05d6 | !decide_p & v845662;
assign a81ccf = hmaster0_p & v84563c | !hmaster0_p & a81cce;
assign ab05de = locked_p & deae59 | !locked_p & !v8c6711;
assign a5fabb = hbusreq2_p & a5fab4 | !hbusreq2_p & !a5fab3;
assign c3b7f0 = hmaster1_p & c3b7ef | !hmaster1_p & c3b7dc;
assign a5fba2 = hmastlock_p & a5fba1 | !hmastlock_p & !v84563c;
assign af34cb = hmaster1_p & af34c4 | !hmaster1_p & af34ca;
assign cea4ae = hmaster0_p & cea4ad | !hmaster0_p & cea43e;
assign a5f43c = hgrant1_p & a5f43a | !hgrant1_p & a5f43b;
assign a5ef2d = hgrant2_p & a5ef2c | !hgrant2_p & v84563c;
assign adaec2 = stateG2_p & v84563c | !stateG2_p & !v845670;
assign c3bc73 = hlock2_p & c3bc72 | !hlock2_p & !deace1;
assign a5f386 = hlock0_p & a60141 | !hlock0_p & a5f385;
assign ab075a = hmaster1_p & ab06c3 | !hmaster1_p & !ab0bf3;
assign c3bc0b = hlock2_p & c3bc0a | !hlock2_p & !deac52;
assign b29942 = hready & b29940 | !hready & b29941;
assign ce9cb4 = hlock2_p & cea448 | !hlock2_p & cea460;
assign c3b7a2 = hbusreq2_p & c3b7a1 | !hbusreq2_p & c3bc75;
assign c3bc76 = hlock2_p & c3bc75 | !hlock2_p & !v84563c;
assign bdb5a2 = decide_p & bdb5a1 | !decide_p & v845660;
assign a5fb63 = hbusreq3 & a5fb54 | !hbusreq3 & a5fb62;
assign b29e59 = decide_p & b29d4e | !decide_p & b29e57;
assign a5f1ef = hlock1_p & a5fc09 | !hlock1_p & !v84563c;
assign a5f1e9 = hbusreq2_p & a5f1e8 | !hbusreq2_p & !v84563c;
assign b2672e = hlock2_p & b2672d | !hlock2_p & b2672c;
assign ab0b30 = hbusreq2_p & ab0b24 | !hbusreq2_p & ab0b21;
assign a5ee95 = hlock2 & a5f3af | !hlock2 & a5ee94;
assign a5f368 = hlock1_p & a5fb8c | !hlock1_p & !ab05a1;
assign a5ea59 = hready & a5ea58 | !hready & a5fc0f;
assign af3500 = hmaster1_p & af3c4c | !hmaster1_p & af34a3;
assign ce9dfd = hbusreq2_p & ce9d48 | !hbusreq2_p & ce9dfc;
assign cea456 = hlock2_p & cea37d | !hlock2_p & cea39b;
assign a5f26c = hbusreq2_p & a5f26b | !hbusreq2_p & v84563c;
assign a5f87f = hbusreq1 & deaca2 | !hbusreq1 & a5f862;
assign b29fc4 = hlock2_p & b29fc3 | !hlock2_p & !b29fa2;
assign c3b770 = hready_p & c3b757 | !hready_p & c3b76f;
assign cea3f7 = hlock1_p & deac51 | !hlock1_p & !cea3be;
assign b29d7a = hready & dead6e | !hready & v84563c;
assign a81ca8 = start_p & a81ca6 | !start_p & a81ca7;
assign ab0b6b = hbusreq2_p & ab0b6a | !hbusreq2_p & ab0b5f;
assign a5f37c = hbusreq1 & a5f374 | !hbusreq1 & v84563c;
assign af354c = hlock1_p & af352c | !hlock1_p & af354b;
assign deadd4 = hgrant1_p & v84563c | !hgrant1_p & deadd3;
assign af3508 = hmaster0_p & af3507 | !hmaster0_p & af34ea;
assign c3bdc9 = hmaster1_p & c3bca4 | !hmaster1_p & c3bdc8;
assign b2995b = hlock2_p & v84563c | !hlock2_p & !b2994a;
assign a5f02d = hready_p & a60147 | !hready_p & a5f02c;
assign a5ef14 = hbusreq0_p & a5edf2 | !hbusreq0_p & a5ef13;
assign dead93 = hlock1_p & b26695 | !hlock1_p & !dead92;
assign b0c0ff = hgrant3_p & b0c0fd | !hgrant3_p & !b0c0fe;
assign d40d34 = stateG10_1_p & d40d33 | !stateG10_1_p & d40d31;
assign a5ef72 = hbusreq2_p & a5ef5a | !hbusreq2_p & a5ef71;
assign a5f3ba = hlock0_p & a5f36b | !hlock0_p & a5f3b8;
assign b29a69 = hbusreq3 & b29a5d | !hbusreq3 & b29a68;
assign b2670c = hlock2_p & b2670a | !hlock2_p & b2670b;
assign a5fbad = start_p & a5fba3 | !start_p & a5fbac;
assign ab06b3 = hlock2 & ab068d | !hlock2 & ab06b2;
assign a5f980 = hmastlock_p & a5f97f | !hmastlock_p & !v84563c;
assign a5f36f = locked_p & a5f369 | !locked_p & a5f36e;
assign b26705 = hmaster1_p & b26704 | !hmaster1_p & b266fb;
assign a5ef79 = hbusreq2 & a5ef78 | !hbusreq2 & a5ef6d;
assign a5f796 = hgrant1_p & v84565a | !hgrant1_p & a5f795;
assign c3b6d3 = hlock3_p & c3b6b7 | !hlock3_p & !c3b6d2;
assign ab0ba8 = hbusreq0_p & b26695 | !hbusreq0_p & !b29d87;
assign c3b6db = hlock0_p & c3bbbb | !hlock0_p & c3b635;
assign deaeac = decide_p & deaeab | !decide_p & v84563c;
assign ab0bf7 = hready_p & ab0be9 | !hready_p & !ab0bf6;
assign a5f01d = hbusreq2_p & a5f01c | !hbusreq2_p & v845644;
assign adaef9 = hgrant0_p & adaeef | !hgrant0_p & adaef8;
assign a5f9e0 = hlock1_p & a81cf0 | !hlock1_p & a5f9df;
assign a5ef98 = hlock0_p & a5ef97 | !hlock0_p & a5f38f;
assign b29a1b = hgrant0_p & c3bceb | !hgrant0_p & !b29a1a;
assign c3b719 = stateG10_1_p & deadba | !stateG10_1_p & c3b678;
assign b266cd = hlock1_p & b26693 | !hlock1_p & b266cc;
assign b26702 = hmaster1_p & b26695 | !hmaster1_p & b266e0;
assign b29cf7 = hlock2 & b29cf3 | !hlock2 & b29cf6;
assign c3b7f7 = hlock0_p & c3b7f6 | !hlock0_p & deadb2;
assign deacde = start_p & v84563c | !start_p & v8e1935;
assign c3b66f = hbusreq2_p & c3b66e | !hbusreq2_p & !c3b66b;
assign b8acea = hgrant2_p & v8c6711 | !hgrant2_p & b8ace9;
assign af3c3e = decide_p & af3c3d | !decide_p & v8567b4;
assign ab06d9 = decide_p & ab06d8 | !decide_p & v84563c;
assign af3594 = hmaster1_p & af352c | !hmaster1_p & af3551;
assign adaef3 = hgrant2_p & v84563c | !hgrant2_p & adaef2;
assign cea324 = hready & cea322 | !hready & cea323;
assign c3bce8 = hlock2_p & c3bce7 | !hlock2_p & v845660;
assign a5fb77 = hlock2_p & a5fb74 | !hlock2_p & a5fb76;
assign v845642 = hbusreq0_p & v84563c | !hbusreq0_p & !v84563c;
assign b29fd6 = hbusreq2_p & b29fd5 | !hbusreq2_p & b29cbb;
assign c3bda7 = hlock2_p & c3bda6 | !hlock2_p & dead2e;
assign a5f489 = hbusreq1 & a5f488 | !hbusreq1 & v84563c;
assign ab06f3 = hlock0_p & b29fc2 | !hlock0_p & !dead41;
assign af3c73 = decide_p & af3c6e | !decide_p & af3c72;
assign a5f73a = hlock0_p & a5f739 | !hlock0_p & v84563c;
assign a5fbef = hbusreq1 & v84563c | !hbusreq1 & a5fbee;
assign af3577 = decide_p & af356e | !decide_p & af3576;
assign a5f7fb = hgrant1_p & a5fa1d | !hgrant1_p & a5f7fa;
assign adaecc = hlock2_p & adaec9 | !hlock2_p & v84563c;
assign c3bdb3 = hbusreq2_p & c3bdb2 | !hbusreq2_p & dead2e;
assign ab05f1 = hlock0_p & v84563c | !hlock0_p & !ab05f0;
assign a81cfd = hmaster1_p & a81cfc | !hmaster1_p & v84563c;
assign b29eeb = hgrant1_p & b29eea | !hgrant1_p & b29ee9;
assign a5f2f6 = hlock0_p & a5f2f5 | !hlock0_p & v84563c;
assign a5fcc4 = decide_p & a5fc67 | !decide_p & a5fcc3;
assign c3bd78 = hgrant1_p & c3bd11 | !hgrant1_p & c3bd77;
assign deae81 = hlock1_p & v84565a | !hlock1_p & !deae80;
assign ab0cfe = decide_p & ab0cfd | !decide_p & !v845662;
assign ab06dc = hbusreq2_p & ab0679 | !hbusreq2_p & ab0bae;
assign ab056e = hgrant2_p & ab0566 | !hgrant2_p & ab056d;
assign a5f57b = hbusreq1_p & a60193 | !hbusreq1_p & v84563c;
assign a5ea9f = hbusreq0 & a5ea9e | !hbusreq0 & v84563c;
assign b29ab4 = hlock2 & b29ab2 | !hlock2 & b29ab3;
assign a5fa13 = hbusreq1_p & v9703fb | !hbusreq1_p & !a60177;
assign a5f731 = hmaster0_p & a5f724 | !hmaster0_p & a5f730;
assign ce9d3f = hmaster1_p & ce9d3e | !hmaster1_p & cea188;
assign c3bcb6 = hmaster0_p & c3bcb5 | !hmaster0_p & c3bcb4;
assign a5efd0 = hlock0_p & a5efcf | !hlock0_p & a5f4fc;
assign a5f1e0 = hlock1_p & a5fba6 | !hlock1_p & a5f1df;
assign c3b88f = hgrant2_p & c3b88c | !hgrant2_p & c3b88e;
assign af350a = decide_p & af3504 | !decide_p & af3509;
assign b2677e = hgrant0_p & b26776 | !hgrant0_p & b2677d;
assign cea344 = hbusreq2_p & cea343 | !hbusreq2_p & v84563c;
assign cea1b0 = hburst0 & cea1ae | !hburst0 & cea1af;
assign a5f3bf = hbusreq3 & a5f3be | !hbusreq3 & v845641;
assign a5f53c = hbusreq1 & a5f53b | !hbusreq1 & deac7a;
assign af3c39 = hlock3_p & af3c34 | !hlock3_p & af3c38;
assign a5edf6 = hbusreq1 & deac17 | !hbusreq1 & v84563c;
assign b266c3 = hmaster0_p & b266c0 | !hmaster0_p & !b266c2;
assign ce9d16 = decide_p & ce9d15 | !decide_p & v84563c;
assign b266a8 = locked_p & v84563c | !locked_p & !b26695;
assign a5f390 = locked_p & v84563c | !locked_p & a5f38f;
assign adaf06 = hlock1_p & adaec4 | !hlock1_p & adaf05;
assign a5f077 = hlock0_p & a5f70a | !hlock0_p & !a5f076;
assign a5e9fe = hbusreq2 & a5e9f7 | !hbusreq2 & a5e9fd;
assign c3b74d = hlock2_p & c3b6db | !hlock2_p & c3b6f6;
assign b29fbd = hlock2_p & c3bcf8 | !hlock2_p & v845660;
assign c3b7a9 = hmaster1_p & c3b7a8 | !hmaster1_p & c3bbbf;
assign ab05d5 = hgrant0_p & ab05c4 | !hgrant0_p & !ab05d4;
assign cea382 = hready & cea151 | !hready & dead7d;
assign a5eb4d = hmaster1_p & a5eb4c | !hmaster1_p & a5f098;
assign a5f3c0 = hmaster1_p & a5f3b7 | !hmaster1_p & a5f3bf;
assign b2a009 = hgrant2_p & b29e95 | !hgrant2_p & !b29ecf;
assign dea7ae = hbusreq3_p & dea79e | !hbusreq3_p & dea7ad;
assign a5f026 = hbusreq2_p & a5fd36 | !hbusreq2_p & a5fd35;
assign af3c17 = hlock3_p & af3c16 | !hlock3_p & v8567b4;
assign c3b65a = hlock3_p & c3b646 | !hlock3_p & !c3b659;
assign ab0cc1 = hbusreq2_p & ab0cc0 | !hbusreq2_p & ab0ad1;
assign ab0673 = hbusreq3 & ab066e | !hbusreq3 & ab0672;
assign ab0ae1 = hbusreq3 & ab0ad6 | !hbusreq3 & ab0ae0;
assign c3b62e = hbusreq2_p & c3b62d | !hbusreq2_p & c3b62c;
assign a5f1c2 = hlock0_p & a5f726 | !hlock0_p & a5f6e9;
assign a81d09 = hready_p & a81d05 | !hready_p & a81d08;
assign a5f2d2 = hbusreq2_p & a5f93c | !hbusreq2_p & v84563c;
assign b29fbc = hmaster0_p & b29fb1 | !hmaster0_p & b29fbb;
assign b29d96 = hbusreq2_p & b29d95 | !hbusreq2_p & b29d94;
assign ab06e4 = hgrant2_p & ab06df | !hgrant2_p & ab06e3;
assign ab0bc4 = hgrant0_p & ab0bb9 | !hgrant0_p & !ab0bc3;
assign dead62 = hbusreq2_p & deacbf | !hbusreq2_p & !v845644;
assign a5efed = hmaster0_p & a5efdc | !hmaster0_p & a5efec;
assign c3b84e = hbusreq2_p & c3b845 | !hbusreq2_p & c3b7e8;
assign c3b6c9 = hbusreq2_p & c3b6c8 | !hbusreq2_p & c3b6a1;
assign a5f207 = hlock3_p & a5f1c1 | !hlock3_p & a5f206;
assign c3b648 = locked_p & v84563c | !locked_p & !deae59;
assign a5f4f2 = hbusreq2 & a5f4ee | !hbusreq2 & a5f4f1;
assign b29edb = hlock2_p & c3bd02 | !hlock2_p & !v84563c;
assign ab0702 = hgrant0_p & bdb59e | !hgrant0_p & !ab0701;
assign b2a00c = hgrant0_p & b2a001 | !hgrant0_p & !b2a00b;
assign b29fec = hlock2_p & c3bd8d | !hlock2_p & !v84563c;
assign a5f285 = hgrant2_p & v84563c | !hgrant2_p & a5f284;
assign b29b33 = decide_p & b29b32 | !decide_p & b29e57;
assign b29ac2 = hgrant2_p & b29ac1 | !hgrant2_p & !b29d5a;
assign b29aa1 = hbusreq2_p & b29aa0 | !hbusreq2_p & b29d92;
assign a5f3c9 = locked_p & a5f3c5 | !locked_p & a5f3c8;
assign ab0759 = hmaster1_p & ab0755 | !hmaster1_p & ab0758;
assign a5fc7c = start_p & v845652 | !start_p & a5fc7b;
assign b29ce6 = hlock2 & b29ce0 | !hlock2 & b29ce5;
assign c3b6c1 = hlock2_p & c3b6c0 | !hlock2_p & c3b698;
assign b29faf = hlock2_p & b29fae | !hlock2_p & dead2e;
assign b29d7f = hlock0_p & b29d7e | !hlock0_p & !dead72;
assign deac6c = hlock1_p & deac51 | !hlock1_p & deac6b;
assign a5f8ca = hready & v84563c | !hready & !deaca0;
assign cea297 = hlock2_p & cea296 | !hlock2_p & v84563c;
assign dead3e = hbusreq2_p & dead3d | !hbusreq2_p & !v84563c;
assign a5f995 = hbusreq2 & a5f993 | !hbusreq2 & a5f994;
assign c3bde7 = hmaster1_p & c3bde6 | !hmaster1_p & c3bcff;
assign deae60 = hlock0_p & deae5f | !hlock0_p & !v84563c;
assign ab0cf8 = hgrant2_p & ab0cdf | !hgrant2_p & ab0cf7;
assign d40d61 = hmaster1_p & d40d31 | !hmaster1_p & d40d60;
assign a5f15b = hready & v84563c | !hready & deacaa;
assign a60184 = stateG2_p & v84563c | !stateG2_p & c06d34;
assign a5f235 = hbusreq2 & a5f232 | !hbusreq2 & a5f234;
assign ab061d = hbusreq0_p & b2997c | !hbusreq0_p & !ab0610;
assign ab0648 = hmaster0_p & ab0643 | !hmaster0_p & ab0647;
assign adaee7 = hmaster0_p & adaee2 | !hmaster0_p & adaee6;
assign a5fbe5 = hmastlock_p & a5fbe4 | !hmastlock_p & v84563c;
assign a5fb1d = hlock1_p & a60186 | !hlock1_p & a5fb1c;
assign deae88 = hbusreq2_p & deae87 | !hbusreq2_p & !deadc4;
assign ab055a = hbusreq1_p & v84563c | !hbusreq1_p & !deaca0;
assign cea26f = hlock1_p & v84563c | !hlock1_p & cea26e;
assign adaed3 = hmaster0_p & adaecb | !hmaster0_p & adaed2;
assign cea1af = hburst1 & cea1ae | !hburst1 & dead6d;
assign c3bde0 = hlock3_p & c3bddf | !hlock3_p & !c3bd7f;
assign c3b6be = hlock1_p & deada8 | !hlock1_p & c3b6bc;
assign dead13 = hmaster1_p & v84563c | !hmaster1_p & dead12;
assign cea1b9 = hburst1 & v84563c | !hburst1 & deacf4;
assign a5ea8c = hmaster0_p & a5ea7a | !hmaster0_p & a5ea8b;
assign a5f3b5 = hlock0_p & a5f3b4 | !hlock0_p & a5f38f;
assign a5eded = hbusreq1_p & a5fbab | !hbusreq1_p & !v84563c;
assign c3b6a5 = hgrant1_p & c3b6a4 | !hgrant1_p & deae74;
assign a5e9c0 = hgrant1_p & a60187 | !hgrant1_p & a5f187;
assign ab0cce = hlock3_p & ab0cca | !hlock3_p & ab0c7f;
assign v9703ff = hmaster0_p & v9703fe | !hmaster0_p & v84563c;
assign b29e9a = hbusreq2_p & v84564c | !hbusreq2_p & v84563c;
assign a81cc7 = hlock3_p & a81cc4 | !hlock3_p & a81cc6;
assign a5f72b = hbusreq0_p & a5f726 | !hbusreq0_p & v84563c;
assign d40d69 = hbusreq0_p & d40d2c | !hbusreq0_p & d40d68;
assign a5f919 = hready & a60189 | !hready & a5f918;
assign af34a1 = hlock0_p & af3c58 | !hlock0_p & af3c4c;
assign a5fa2b = hready & v84563c | !hready & !deac19;
assign b29949 = hready & b29946 | !hready & b29941;
assign a81d0b = hready_p & a81ceb | !hready_p & a81d0a;
assign deaea4 = hbusreq2_p & deaea3 | !hbusreq2_p & !v84563c;
assign b29d8d = hlock2 & b29d89 | !hlock2 & b29d8c;
assign ab0b39 = hlock0_p & v84563c | !hlock0_p & b29d34;
assign a5f987 = start_p & a81ca6 | !start_p & a5f986;
assign c3bc64 = hlock0_p & c3bc63 | !hlock0_p & !deacfc;
assign dead4b = hmaster1_p & dead49 | !hmaster1_p & !dead4a;
assign cea1a4 = hmaster1_p & cea1a3 | !hmaster1_p & cea188;
assign a5ef0e = hbusreq1_p & a5fce1 | !hbusreq1_p & !v84563c;
assign ab0b86 = hgrant2_p & ab0b83 | !hgrant2_p & ab0b85;
assign dead27 = hbusreq3 & dead26 | !hbusreq3 & v84563c;
assign a5ea7e = locked_p & a5ea7d | !locked_p & v845641;
assign ab051b = hlock0_p & v84563c | !hlock0_p & ab0519;
assign c3b7c1 = hlock0_p & c3bd21 | !hlock0_p & deadb2;
assign c3b6e1 = hbusreq0_p & c3b647 | !hbusreq0_p & c3b6e0;
assign v970442 = hmaster1_p & v84563c | !hmaster1_p & v970441;
assign b2a01e = stateA1_p & dead31 | !stateA1_p & v84563c;
assign d40d97 = hgrant2_p & d40d95 | !hgrant2_p & d40d96;
assign a5f9f6 = hlock1_p & a60168 | !hlock1_p & a5f9f5;
assign dead23 = hbusreq3 & dead22 | !hbusreq3 & v84563c;
assign a5f139 = hbusreq0 & a5f137 | !hbusreq0 & a5f138;
assign a5f038 = hbusreq2_p & v845644 | !hbusreq2_p & v84563c;
assign b29b09 = decide_p & b29b08 | !decide_p & b29e57;
assign a5fc30 = hlock2_p & a5fc2b | !hlock2_p & a5fc2f;
assign cea85d = hlock0_p & cea85c | !hlock0_p & v84563c;
assign ab0c4a = hmaster1_p & ab0c42 | !hmaster1_p & ab0c49;
assign b29cf3 = hlock0_p & b29cf0 | !hlock0_p & b29cf2;
assign a5efe6 = hlock0_p & a5f55a | !hlock0_p & a5ef81;
assign cea31c = hmaster0_p & cea15e | !hmaster0_p & cea31b;
assign cea443 = hlock0_p & cea389 | !hlock0_p & cea37b;
assign a5f0d9 = hlock0_p & a5fa00 | !hlock0_p & a5f0d0;
assign c3b626 = locked_p & deae50 | !locked_p & c3b625;
assign ab0be1 = hmaster0_p & ab0b61 | !hmaster0_p & ab0be0;
assign b298a2 = hlock2_p & v84563c | !hlock2_p & b298a1;
assign c3b694 = hlock1_p & v84563c | !hlock1_p & !c3b693;
assign ab0aeb = hmastlock_p & deaca0 | !hmastlock_p & !v84563c;
assign a5f0ed = hbusreq2_p & a5f0ec | !hbusreq2_p & a5f0eb;
assign b29d3d = hbusreq3 & b29d3b | !hbusreq3 & !b29d3c;
assign a5f856 = hlock2_p & a5f821 | !hlock2_p & !a5f855;
assign c3bcaa = hbusreq3 & c3bca9 | !hbusreq3 & !dead3e;
assign cea250 = hmastlock_p & cea24f | !hmastlock_p & v84566c;
assign bdb5ab = decide_p & bdb597 | !decide_p & !bdb5aa;
assign cea257 = hlock1_p & v84563c | !hlock1_p & !cea256;
assign c3bbbd = hlock2_p & c3bbbc | !hlock2_p & v845660;
assign a5f149 = hbusreq1 & deacaa | !hbusreq1 & a5f148;
assign a5f747 = hbusreq3 & a5f746 | !hbusreq3 & v84563c;
assign ab0b6d = hmaster1_p & ab0b62 | !hmaster1_p & ab0b6c;
assign ce9dd4 = hgrant2_p & ce9d34 | !hgrant2_p & ce9dd3;
assign b26699 = locked_p & b26693 | !locked_p & b26695;
assign ab0d05 = hlock2_p & ab0d03 | !hlock2_p & ab0d04;
assign ab0b81 = hlock2_p & ab0b80 | !hlock2_p & v84563c;
assign a5eedd = hbusreq2 & a5f560 | !hbusreq2 & a5eedc;
assign af34f6 = hgrant2_p & af3497 | !hgrant2_p & d40d60;
assign b299aa = decide_p & b29976 | !decide_p & b29e57;
assign c3b633 = hlock2_p & c3b632 | !hlock2_p & c3b631;
assign a5fc20 = hbusreq3 & a5fc1f | !hbusreq3 & a5fbc4;
assign a5f146 = hlock0_p & a5f86c | !hlock0_p & a5f144;
assign a5f41b = hlock1_p & v84565a | !hlock1_p & ab055c;
assign a5fa5e = hready & a60168 | !hready & v84565a;
assign cea49a = hlock0_p & cea499 | !hlock0_p & cea405;
assign ab0cee = hgrant2_p & ab0be2 | !hgrant2_p & ab0ced;
assign a5f249 = hready & a5f7f5 | !hready & a5fa1d;
assign b29e5d = hmaster1_p & v84563c | !hmaster1_p & b29e5c;
assign a5f9e7 = hlock1_p & a5f9dd | !hlock1_p & a5f9df;
assign a5ee23 = locked_p & a5ee22 | !locked_p & !v845641;
assign c3bdf5 = hmaster0_p & c3bdf4 | !hmaster0_p & !c3bd7e;
assign c3b641 = hlock0_p & c3b631 | !hlock0_p & c3b63f;
assign b266aa = hlock2_p & b266a9 | !hlock2_p & b266a8;
assign ab050d = hbusreq2_p & ab050c | !hbusreq2_p & ab0d07;
assign af356d = hmaster0_p & af3569 | !hmaster0_p & af356c;
assign a5f3ca = hbusreq1_p & a5fc84 | !hbusreq1_p & !v84563c;
assign a5ee29 = hlock0_p & a5ee23 | !hlock0_p & !a5ee28;
assign a5fbfb = hready & a5fbfa | !hready & !cea151;
assign a5ea22 = hbusreq0 & a5ea21 | !hbusreq0 & !v84563c;
assign ab0bb3 = hgrant2_p & ab0bb1 | !hgrant2_p & ab0bb2;
assign ab05e4 = hbusreq2_p & ab052c | !hbusreq2_p & ab05e3;
assign ce9d4b = hmaster1_p & ce9d45 | !hmaster1_p & ce9d4a;
assign a5ee1a = hbusreq2_p & a5ee19 | !hbusreq2_p & a5ee15;
assign cea2ed = hmaster1_p & cea85f | !hmaster1_p & cea2ec;
assign ab0ce5 = hready_p & ab0cde | !hready_p & ab0ce4;
assign b266c2 = hmaster1_p & b266c1 | !hmaster1_p & b266b3;
assign ce9cdf = jx1_p & ce9ccf | !jx1_p & ce9cde;
assign b29d0e = hlock2_p & v84563c | !hlock2_p & !b29d0d;
assign a5f92d = hgrant2_p & a5f92c | !hgrant2_p & a5fd28;
assign a5f752 = hmaster1_p & a5f74f | !hmaster1_p & a5f751;
assign af3499 = hmaster0_p & af3498 | !hmaster0_p & d40d60;
assign c3b7b5 = hmaster0_p & c3b7af | !hmaster0_p & c3b7b4;
assign cea3cd = hready & cea3cb | !hready & cea3cc;
assign c3bdcd = decide_p & c3bdcc | !decide_p & v845660;
assign c3bcef = hready & deacdf | !hready & !v84563c;
assign c3bcd4 = hmaster0_p & c3bcd0 | !hmaster0_p & c3bcd3;
assign c3bbfd = hlock2_p & c3bbfc | !hlock2_p & !deac52;
assign dea6b9 = locked_p & deaeb6 | !locked_p & !deae5a;
assign a5fc6c = hready & b266a2 | !hready & a5fc6b;
assign c3b79e = hbusreq2_p & c3b79d | !hbusreq2_p & c3b79b;
assign c3bcf3 = hlock2_p & c3bcf2 | !hlock2_p & v845660;
assign ab0596 = hmaster1_p & ab058e | !hmaster1_p & ab0595;
assign a5ef92 = hmaster1_p & a5ef91 | !hmaster1_p & !v84563c;
assign a5fa1e = stateG10_1_p & a5fa1d | !stateG10_1_p & a5fa1c;
assign b26726 = hbusreq2_p & b26725 | !hbusreq2_p & !b266a2;
assign cea48e = decide_p & cea48d | !decide_p & a57859;
assign b29f6a = hbusreq2_p & b29f69 | !hbusreq2_p & deacab;
assign a5f28c = hready_p & a5f21b | !hready_p & a5f28b;
assign a5f585 = hbusreq0 & a5f569 | !hbusreq0 & !a5f584;
assign b29f9e = hlock0_p & dead41 | !hlock0_p & !b29f9d;
assign b26769 = hgrant3_p & b26709 | !hgrant3_p & !b26768;
assign ab0bf0 = hbusreq2_p & ab0b02 | !hbusreq2_p & v845644;
assign v84564c = hlock2_p & v84563c | !hlock2_p & !v84563c;
assign d40d81 = hlock1_p & d40d31 | !hlock1_p & d40d80;
assign a5ec30 = hbusreq3_p & a5ec24 | !hbusreq3_p & a5f6e2;
assign ab075f = hbusreq3_p & ab0731 | !hbusreq3_p & ab075e;
assign a5f1b6 = hlock2_p & a5f9a8 | !hlock2_p & a5f1b5;
assign af3c65 = hlock2_p & af3c63 | !hlock2_p & af3c64;
assign c3bc37 = hbusreq3 & c3bc34 | !hbusreq3 & !c3bc36;
assign b2982d = hbusreq1_p & b2982c | !hbusreq1_p & dead7b;
assign dead00 = hbusreq2_p & deacff | !hbusreq2_p & deacfd;
assign a5f399 = hlock2_p & a5f395 | !hlock2_p & a5f398;
assign ab0b59 = hbusreq3 & ab0b55 | !hbusreq3 & ab0b58;
assign a5f56c = hbusreq1 & a5f56b | !hbusreq1 & !v84563c;
assign a5ee90 = hbusreq2_p & a5ee8f | !hbusreq2_p & a5ee8e;
assign a5eb1c = hlock3_p & a5eafc | !hlock3_p & a5ea1d;
assign c3bc7a = hlock1_p & dead6e | !hlock1_p & v84563c;
assign deacf3 = stateA1_p & v84563c | !stateA1_p & !deacf2;
assign c3b7fb = hlock2_p & c3b7fa | !hlock2_p & c3b7e4;
assign c3b6d0 = hgrant2_p & c3b6ce | !hgrant2_p & c3b6cf;
assign cea361 = hmaster1_p & cea35e | !hmaster1_p & cea360;
assign ab0b92 = hlock2 & ab0b90 | !hlock2 & ab0b91;
assign ab0c7c = hbusreq2_p & ab0c7a | !hbusreq2_p & !ab0bd9;
assign c3b64d = hbusreq3 & c3b647 | !hbusreq3 & c3b64c;
assign a5f202 = hbusreq2_p & a5f201 | !hbusreq2_p & v84563c;
assign cea288 = hbusreq2_p & cea286 | !hbusreq2_p & cea89c;
assign ab06bd = hbusreq0_p & deaca1 | !hbusreq0_p & ab06bc;
assign a5fbc6 = hready & a5fb73 | !hready & !v84563c;
assign ab0c2d = decide_p & ab0c2c | !decide_p & v84563c;
assign b29ee8 = hmastlock_p & b29ee7 | !hmastlock_p & v84566c;
assign ab0ca9 = hmaster1_p & ab0ca7 | !hmaster1_p & ab0ca8;
assign a5f437 = hlock1_p & a5fbab | !hlock1_p & !a5f436;
assign a5f8f0 = hlock2_p & a5f8ec | !hlock2_p & !a5f8ef;
assign a5f6f1 = hlock2 & a5f6eb | !hlock2 & a5f6f0;
assign ab063e = hbusreq3_p & ab05da | !hbusreq3_p & ab063d;
assign a5fa87 = hlock1_p & a60172 | !hlock1_p & a5fa86;
assign b29d33 = hlock2 & b29cf2 | !hlock2 & v84565a;
assign b29d57 = hmaster1_p & c3bceb | !hmaster1_p & b29d56;
assign a5ea50 = hbusreq1_p & a5fb8a | !hbusreq1_p & a5fc78;
assign deae69 = hbusreq2_p & deae66 | !hbusreq2_p & !deae68;
assign cea39c = hready & v845646 | !hready & !v84563c;
assign a5f87a = hlock0_p & a5f9c2 | !hlock0_p & a5f879;
assign b29ed9 = hbusreq3 & b29ed8 | !hbusreq3 & !v84564a;
assign d40d71 = hmaster1_p & v84563c | !hmaster1_p & d40d70;
assign cea432 = hbusreq2_p & cea431 | !hbusreq2_p & cea405;
assign a5f097 = hbusreq0 & a5f094 | !hbusreq0 & a5f096;
assign ab05cc = hlock2_p & ab05cb | !hlock2_p & ab05a8;
assign b26751 = hmaster1_p & b2674e | !hmaster1_p & !b26750;
assign b29eec = hlock1_p & deac51 | !hlock1_p & b29eeb;
assign a5ede9 = hbusreq1_p & deac52 | !hbusreq1_p & v84563c;
assign ab06f8 = hlock0_p & b29fb5 | !hlock0_p & !ab066a;
assign deae57 = hmaster1_p & deae56 | !hmaster1_p & deac0f;
assign b29d1f = hbusreq3 & b29d0f | !hbusreq3 & b29d1e;
assign ab0654 = hgrant3_p & ab064b | !hgrant3_p & !ab0653;
assign deacb4 = hmastlock_p & deacb3 | !hmastlock_p & v84563c;
assign a5f081 = hlock2_p & a5fb7b | !hlock2_p & a5f080;
assign v970400 = hlock3_p & v9703ff | !hlock3_p & v84563c;
assign c3b7e7 = hbusreq2_p & c3b7e5 | !hbusreq2_p & !c3b7e6;
assign a81d02 = hgrant3_p & a81ccc | !hgrant3_p & a81d01;
assign cea17f = hgrant0_p & v84563c | !hgrant0_p & cea17e;
assign cea439 = hlock0_p & cea434 | !hlock0_p & cea412;
assign ce9cf6 = hbusreq2_p & cea1c1 | !hbusreq2_p & cea1c0;
assign cea463 = hlock0_p & cea462 | !hlock0_p & cea44b;
assign deae19 = hgrant0_p & deae0a | !hgrant0_p & deae18;
assign a5f29d = hmaster1_p & a5f29c | !hmaster1_p & !a5f751;
assign ab0615 = hgrant2_p & ab0614 | !hgrant2_p & cea15a;
assign a5fad7 = hlock2_p & a5fad1 | !hlock2_p & a5fad6;
assign ab06cf = hbusreq2_p & ab06ce | !hbusreq2_p & ab06b5;
assign b29ceb = hlock2_p & b29ce6 | !hlock2_p & b29cea;
assign ab0b16 = hlock0_p & ab0b15 | !hlock0_p & deac86;
assign ab0acd = hbusreq2_p & ab0acc | !hbusreq2_p & ab0acb;
assign a5fc72 = hbusreq2_p & c3bcf8 | !hbusreq2_p & a5fc71;
assign a5f83a = hgrant1_p & a5f839 | !hgrant1_p & a5f837;
assign a5fca6 = hbusreq1 & a5fca3 | !hbusreq1 & !a5fca5;
assign af34ff = hready_p & af34fd | !hready_p & af34fe;
assign b29e70 = hmaster0_p & b29e66 | !hmaster0_p & !b29e6f;
assign a5fc89 = locked_p & a5fc88 | !locked_p & v84563c;
assign af35b8 = hmaster1_p & af35b7 | !hmaster1_p & af3551;
assign cea45a = hbusreq2_p & cea459 | !hbusreq2_p & cea3aa;
assign deadf9 = hlock0_p & deadf8 | !hlock0_p & v84563c;
assign b29a19 = hmaster1_p & b29fc8 | !hmaster1_p & b29e48;
assign b266a1 = hbusreq1_p & b26695 | !hbusreq1_p & !b266a0;
assign c3b81d = hlock2_p & c3b7a0 | !hlock2_p & !c3b7ad;
assign b29d22 = hbusreq3 & b29d20 | !hbusreq3 & b29d21;
assign deacd2 = hlock2_p & deacbe | !hlock2_p & v84563c;
assign a5ea8d = hgrant0_p & v84563c | !hgrant0_p & a5ea8c;
assign a5ef6e = hbusreq2 & a5ef6c | !hbusreq2 & a5ef6d;
assign cea333 = hlock1_p & v84563c | !hlock1_p & !cea332;
assign a5fafd = hready & a5fafc | !hready & a6018b;
assign c3bd94 = hlock0_p & c3bc48 | !hlock0_p & c3bcee;
assign deadf1 = hbusreq2_p & deadef | !hbusreq2_p & !deacbe;
assign dead16 = hbusreq2_p & dead15 | !hbusreq2_p & deacfb;
assign cea44b = hbusreq0_p & cea39b | !hbusreq0_p & cea44a;
assign af34d7 = hgrant2_p & af34d6 | !hgrant2_p & af34bb;
assign ab0cd5 = hbusreq2_p & ab0c1d | !hbusreq2_p & v845644;
assign d40d6f = locked_p & d40d6e | !locked_p & v84563c;
assign a5efdb = hgrant2_p & a5efd5 | !hgrant2_p & a5efda;
assign b29c3d = hbusreq3 & b29c3c | !hbusreq3 & v84563c;
assign af3c45 = hready_p & af3c43 | !hready_p & af3c44;
assign a5f6e2 = hgrant3_p & a5fd3b | !hgrant3_p & a5f6e1;
assign c3b61e = hready_p & c3b60b | !hready_p & c3b61d;
assign c3bccd = hbusreq3 & c3bccb | !hbusreq3 & c3bccc;
assign cea373 = jx0_p & cea1a9 | !jx0_p & cea372;
assign a5efc2 = hbusreq2_p & a5ee79 | !hbusreq2_p & a5efc1;
assign c3b752 = hbusreq2_p & c3b751 | !hbusreq2_p & c3b635;
assign c3b809 = hlock0_p & c3bd99 | !hlock0_p & !cea17a;
assign c3b77b = hlock3_p & c3bcc3 | !hlock3_p & c3b77a;
assign d5edb8 = stateG3_1_p & v845670 | !stateG3_1_p & v84563c;
assign b29d9c = hbusreq3 & v84563c | !hbusreq3 & c3bceb;
assign a81cec = hmaster1_p & a81cb1 | !hmaster1_p & a81cb5;
assign a5ee3f = hlock2_p & a5ee3c | !hlock2_p & a5ee3e;
assign ce9d4e = hgrant2_p & cea31a | !hgrant2_p & !ce9d4d;
assign ab06d2 = hlock2 & ab06d0 | !hlock2 & ab06d1;
assign d40d89 = hmaster0_p & d40d85 | !hmaster0_p & d40d88;
assign b26692 = stateA1_p & v84563c | !stateA1_p & !v8e1935;
assign a5eb9b = hgrant0_p & a60144 | !hgrant0_p & a5eb9a;
assign a5fbd7 = hlock1_p & a5fb8a | !hlock1_p & v84563c;
assign ab0620 = hbusreq2_p & ab05b6 | !hbusreq2_p & ab061f;
assign a5ee88 = hlock2_p & a5ee87 | !hlock2_p & a5ee18;
assign ab05ed = hbusreq0_p & b29947 | !hbusreq0_p & b29946;
assign ab0bd5 = hlock2 & ab0bd4 | !hlock2 & ab0b3b;
assign v94aab7 = hmaster1_p & v84563c | !hmaster1_p & !v84564a;
assign af3487 = hgrant2_p & af3485 | !hgrant2_p & af3486;
assign b29f7d = hlock2_p & b29f7c | !hlock2_p & !b29f59;
assign c3bc58 = hlock0_p & b26720 | !hlock0_p & !b26695;
assign b26760 = hmaster1_p & b266a8 | !hmaster1_p & b2675f;
assign b29f75 = hgrant2_p & b29f74 | !hgrant2_p & b29e6b;
assign c3b80f = locked_p & cea2e8 | !locked_p & c3bc47;
assign b29ff1 = hmaster0_p & b29fef | !hmaster0_p & b29ff0;
assign b29e9d = hbusreq2_p & b29cf8 | !hbusreq2_p & v845644;
assign a5f269 = hbusreq2_p & a5f268 | !hbusreq2_p & v84563c;
assign a5f706 = hlock1_p & a5fc84 | !hlock1_p & !a5f705;
assign a5ee12 = locked_p & a5ee11 | !locked_p & a60140;
assign af3581 = hgrant2_p & af352f | !hgrant2_p & af3580;
assign b29b0a = hready_p & b29ac7 | !hready_p & b29b09;
assign b299f0 = hmaster1_p & v84563c | !hmaster1_p & b29e65;
assign dead1d = hgrant2_p & dead17 | !hgrant2_p & dead1c;
assign c3bd41 = hlock2_p & c3bd3f | !hlock2_p & !deadc4;
assign a5ee16 = hlock0_p & a5f36c | !hlock0_p & a5ee14;
assign ab053a = stateG10_1_p & v84563c | !stateG10_1_p & ab0539;
assign c3bc3b = hgrant2_p & c3bc37 | !hgrant2_p & c3bc3a;
assign a60168 = hmastlock_p & a60167 | !hmastlock_p & v84563c;
assign cea270 = stateG10_1_p & deacb3 | !stateG10_1_p & deadb9;
assign a5fb34 = hlock2_p & a5fb33 | !hlock2_p & v84563c;
assign ce9d3d = hbusreq2_p & cea297 | !hbusreq2_p & cea2a5;
assign b29e6c = hgrant2_p & b29e6a | !hgrant2_p & b29e6b;
assign a5eba3 = decide_p & a5eb9b | !decide_p & a5eba2;
assign a5ebed = hgrant3_p & a5eb8a | !hgrant3_p & a5ebec;
assign a5e9dd = hgrant2_p & a5e9d8 | !hgrant2_p & a5e9dc;
assign adaf16 = hmaster0_p & adaf15 | !hmaster0_p & v84563c;
assign deadac = hlock1_p & deac51 | !hlock1_p & !deadab;
assign b840b3 = hgrant3_p & b840af | !hgrant3_p & b840b2;
assign c3bcc6 = hlock2_p & c3bcc5 | !hlock2_p & !v84563c;
assign adaf14 = decide_p & v84563c | !decide_p & adaf13;
assign a5ee7f = hlock0_p & a5f39f | !hlock0_p & a5f36b;
assign v8c6449 = stateG3_1_p & v84563c | !stateG3_1_p & v845670;
assign a5ee74 = hlock0_p & a5ee38 | !hlock0_p & a5ee73;
assign b29a54 = hbusreq3 & b29a53 | !hbusreq3 & v84563c;
assign b8ace1 = decide_p & b8ace0 | !decide_p & b8acd9;
assign a5efac = hbusreq2 & a5efab | !hbusreq2 & a5ee26;
assign a5f565 = hready & a5f520 | !hready & a5f41d;
assign a5ee05 = hlock0_p & a60141 | !hlock0_p & a5f36b;
assign a5ee46 = hbusreq1_p & a5fb89 | !hbusreq1_p & v84563c;
assign deae27 = hbusreq2_p & deae1f | !hbusreq2_p & deac1e;
assign b2674e = hgrant2_p & b2674d | !hgrant2_p & !b266c1;
assign a5fba4 = stateA1_p & a5fb9d | !stateA1_p & a5f9da;
assign ab060f = hlock2_p & ab060c | !hlock2_p & ab060e;
assign c3b872 = hready_p & c3b830 | !hready_p & c3b871;
assign ab0cbc = decide_p & ab0cbb | !decide_p & v845662;
assign cea158 = hmaster0_p & cea14a | !hmaster0_p & cea157;
assign deaeb3 = locked_p & v84563c | !locked_p & deae67;
assign b299e5 = hgrant0_p & b299dc | !hgrant0_p & !b299e4;
assign deacd6 = hbusreq3 & deacc5 | !hbusreq3 & !deacd5;
assign c3bcbd = hmaster0_p & cea187 | !hmaster0_p & !c3bcbc;
assign a5fce6 = hbusreq0_p & a5fcdf | !hbusreq0_p & a5fce5;
assign c3bc2c = hbusreq3 & c3bc2a | !hbusreq3 & c3bc2b;
assign a5fcea = hmaster1_p & a5fcd0 | !hmaster1_p & a5fce9;
assign a5ee4e = hready & a5f515 | !hready & v84563c;
assign ab0b8f = hlock2_p & ab0b8b | !hlock2_p & ab0b8e;
assign b2671b = hmaster1_p & b26714 | !hmaster1_p & !b2671a;
assign ab0c5f = hlock2 & ab0b16 | !hlock2 & ab0c5e;
assign a5e9bb = hready & a5e9ba | !hready & a5f797;
assign c3b7e0 = hgrant2_p & c3b7de | !hgrant2_p & c3b7df;
assign a5efab = hlock2 & a5f38f | !hlock2 & a5ee65;
assign dead88 = hmaster0_p & dead86 | !hmaster0_p & dead87;
assign dea6fe = hready_p & dea6fc | !hready_p & !dea6fd;
assign a5ef9c = hmaster1_p & a5ef9b | !hmaster1_p & a60144;
assign b29ec3 = hbusreq2_p & b29ec2 | !hbusreq2_p & v84563c;
assign b29efd = hlock2_p & b29eee | !hlock2_p & !b29efc;
assign ce9d56 = hmaster1_p & ce9d45 | !hmaster1_p & ce9d55;
assign a5e9b4 = hbusreq0_p & a5fa5b | !hbusreq0_p & a5fa2d;
assign c3bd99 = locked_p & v845648 | !locked_p & c3bd98;
assign ab0ca8 = hbusreq2_p & ab0c86 | !hbusreq2_p & dead2e;
assign a5f6f6 = hlock0_p & a5f6f3 | !hlock0_p & a5f6f5;
assign a5f9a3 = locked_p & a5fbe8 | !locked_p & a5f9a2;
assign cea23b = hlock3_p & cea1c8 | !hlock3_p & cea23a;
assign af3c30 = hbusreq2_p & af3c2f | !hbusreq2_p & af3c2e;
assign a5efd6 = hlock0_p & a5efcf | !hlock0_p & a5ef5e;
assign a5ea6d = hmaster1_p & a5ea6c | !hmaster1_p & a5fbc5;
assign a5f2ff = hbusreq2_p & a5f2fe | !hbusreq2_p & v84563c;
assign a5f478 = hbusreq2_p & a5f421 | !hbusreq2_p & a5f40e;
assign b29d64 = hgrant2_p & c3bcfb | !hgrant2_p & !b29c3c;
assign ce9dc7 = hbusreq0_p & cea887 | !hbusreq0_p & !deacaa;
assign a5f270 = hmaster1_p & v84563c | !hmaster1_p & a5f26f;
assign a5f923 = hlock0_p & a5f922 | !hlock0_p & a5f879;
assign a5fc70 = hready & b266a0 | !hready & a5fc69;
assign a5f941 = hgrant1_p & a5f8e1 | !hgrant1_p & a5f940;
assign c3b8b7 = hgrant3_p & c3b889 | !hgrant3_p & !c3b8b6;
assign ab0c86 = hlock2_p & ab0c85 | !hlock2_p & dead2e;
assign b2a006 = hgrant2_p & b29e95 | !hgrant2_p & !b2a005;
assign ab0c3f = hlock2 & v84563c | !hlock2 & ab0c3e;
assign dead84 = hbusreq2_p & v845660 | !hbusreq2_p & v84563c;
assign cea46c = hlock0_p & cea462 | !hlock0_p & cea37c;
assign b29951 = hlock0_p & b29950 | !hlock0_p & !deada8;
assign a5f2e5 = hlock0_p & a5f2e4 | !hlock0_p & a5f727;
assign a5ee6f = hlock2 & a5ee6c | !hlock2 & a5ee6e;
assign a5f4fa = hlock1_p & v84565a | !hlock1_p & b8acdb;
assign cea3bb = hlock1_p & deac51 | !hlock1_p & !cea3ba;
assign c3bc09 = hlock1_p & v84563c | !hlock1_p & !c3bc08;
assign ab0af3 = hlock0_p & v84563c | !hlock0_p & !b29ce8;
assign a5edd2 = hgrant2_p & a5edbc | !hgrant2_p & a5edd1;
assign b29a88 = hbusreq2_p & b29a87 | !hbusreq2_p & !v84563c;
assign a5efcb = hmaster1_p & a5efca | !hmaster1_p & v84563c;
assign c3b7d2 = hbusreq2_p & c3b7d1 | !hbusreq2_p & !c3b7d0;
assign a5f40b = hlock1_p & v84563c | !hlock1_p & a5f409;
assign a5fc2c = hbusreq0_p & v845641 | !hbusreq0_p & a5fc1a;
assign c3bdfa = hlock0_p & c3bdf9 | !hlock0_p & c3bcef;
assign d40d5b = hmaster0_p & d40d57 | !hmaster0_p & d40d5a;
assign ab05ef = hbusreq2_p & ab0563 | !hbusreq2_p & ab05ee;
assign af3579 = locked_p & b29d6c | !locked_p & v84563c;
assign bdb584 = hlock1_p & v84565a | !hlock1_p & cea0bb;
assign ce9db7 = hbusreq2_p & cea236 | !hbusreq2_p & cea235;
assign b29eac = locked_p & b29eab | !locked_p & v84563c;
assign c3b662 = stateG10_1_p & deacb4 | !stateG10_1_p & c3b661;
assign cea8a2 = hbusreq3 & cea8a0 | !hbusreq3 & cea8a1;
assign cea3ba = hgrant1_p & cea3b9 | !hgrant1_p & cea255;
assign af357e = hbusreq1_p & v84563c | !hbusreq1_p & b29d6c;
assign a5f1cd = hbusreq2_p & a5f1cc | !hbusreq2_p & v84563c;
assign cea279 = hbusreq2_p & cea25a | !hbusreq2_p & cea86c;
assign a5fd13 = hbusreq2 & a5fd10 | !hbusreq2 & a5fd12;
assign ce9cdb = decide_p & ce9cd2 | !decide_p & a57859;
assign b2990e = hmaster0_p & b298b3 | !hmaster0_p & b2990d;
assign dead60 = hmaster1_p & dead5e | !hmaster1_p & !dead5f;
assign b29ef5 = hready & deacb7 | !hready & !v84565a;
assign a5f3a0 = hready & v84563c | !hready & v8c6711;
assign a5ef32 = hready_p & a5eed6 | !hready_p & a5ef31;
assign a5edd6 = hlock2_p & a5edd5 | !hlock2_p & a5f567;
assign ab072e = hlock3_p & ab0722 | !hlock3_p & ab06d7;
assign c3bccb = hbusreq2_p & c3bcc6 | !hbusreq2_p & c3bcc5;
assign a5fcbf = hbusreq3 & a5fcbc | !hbusreq3 & v84563c;
assign b29ff8 = hmaster1_p & b29e6c | !hmaster1_p & !b29ff7;
assign deae76 = hlock1_p & deac51 | !hlock1_p & !deae75;
assign a5edcf = hlock0_p & a5edcc | !hlock0_p & a5f4f0;
assign dea734 = hbusreq2_p & dead9a | !hbusreq2_p & !dea733;
assign b29f04 = hburst1 & deacb3 | !hburst1 & b29f03;
assign v97042e = hlock3_p & v97042b | !hlock3_p & v97042d;
assign a5f90b = hbusreq2_p & a5f90a | !hbusreq2_p & v84563c;
assign a5f967 = hbusreq2_p & a5f966 | !hbusreq2_p & a60142;
assign ab0c72 = hbusreq2_p & ab0bd6 | !hbusreq2_p & v84563c;
assign cea36f = decide_p & cea36e | !decide_p & a57859;
assign b29b12 = decide_p & b29b11 | !decide_p & v84563c;
assign a5f6dc = hbusreq2_p & a5fad7 | !hbusreq2_p & v84563c;
assign c3bdce = hlock1_p & v84563c | !hlock1_p & !dea6c9;
assign be34e5 = decide_p & be34df | !decide_p & v84564a;
assign a5ef7e = hbusreq2 & a5ef7c | !hbusreq2 & a5ef7d;
assign a5f43a = stateG10_1_p & a5fa1d | !stateG10_1_p & a5f439;
assign deac55 = hbusreq1_p & deac52 | !hbusreq1_p & !v84563c;
assign a5ec19 = hmaster0_p & a5f01b | !hmaster0_p & a5ec18;
assign cea3cf = hlock2_p & cea3ce | !hlock2_p & cea3cd;
assign c3bdf8 = hready & deacec | !hready & !v84563c;
assign deae00 = hmaster1_p & deadfb | !hmaster1_p & deadff;
assign ab076a = jx1_p & ab075f | !jx1_p & ab0655;
assign cea1ad = stateA1_p & v84563c | !stateA1_p & cea1ac;
assign bdb597 = hlock3_p & bdb596 | !hlock3_p & v84565a;
assign cea8aa = hgrant1_p & cea8a8 | !hgrant1_p & cea8a9;
assign a5ee48 = hready & a5ee47 | !hready & !c3b6f8;
assign b2994a = hlock0_p & b29949 | !hlock0_p & !v84563c;
assign dead49 = hgrant2_p & dead47 | !hgrant2_p & !dead48;
assign a5eef5 = hbusreq2_p & a5eef1 | !hbusreq2_p & a5eeea;
assign ab059c = hlock2 & ab0528 | !hlock2 & ab059b;
assign b298ac = hlock2_p & v84563c | !hlock2_p & !b298ab;
assign deada6 = stateA1_p & v8c607d | !stateA1_p & v8c6449;
assign ab0b61 = hbusreq2_p & ab0b60 | !hbusreq2_p & ab0b5f;
assign a5ee81 = hbusreq2_p & a5ee80 | !hbusreq2_p & a5ee7f;
assign a5fcf4 = hbusreq1_p & a5fbab | !hbusreq1_p & a5fce1;
assign a5fb6a = hready & v84563c | !hready & !b2671f;
assign a5f557 = hgrant1_p & ab055b | !hgrant1_p & b29914;
assign b8ace3 = hlock1_p & v84563c | !hlock1_p & b8acda;
assign a5fb6e = hbusreq2_p & a5fb6d | !hbusreq2_p & a5fb6c;
assign c3b84b = hlock2_p & c3b849 | !hlock2_p & !c3b84a;
assign b26771 = decide_p & b26770 | !decide_p & b2676d;
assign b2a00d = decide_p & b2a00c | !decide_p & b29e57;
assign cea182 = decide_p & cea0f2 | !decide_p & a57859;
assign c3bd35 = stateA1_p & v84563c | !stateA1_p & v8c6449;
assign deac4e = start_p & deac4a | !start_p & deac4d;
assign a5f881 = hlock0_p & a5f87d | !hlock0_p & a5f880;
assign a5eef3 = hbusreq3 & a5eedf | !hbusreq3 & !a5eef2;
assign cea153 = hlock0_p & cea152 | !hlock0_p & v84563c;
assign cea386 = hbusreq2_p & cea385 | !hbusreq2_p & cea384;
assign b29ee5 = start_p & deac4a | !start_p & v84563c;
assign deacda = hlock3_p & deac9f | !hlock3_p & deacd9;
assign a5ea33 = hbusreq2 & a5f089 | !hbusreq2 & a5fbc1;
assign b29fa2 = hlock2 & b29f9e | !hlock2 & b29fa1;
assign deac4a = stateA1_p & v84563c | !stateA1_p & !v845652;
assign ab0681 = hbusreq3 & b29a4d | !hbusreq3 & !v84563c;
assign af3c10 = jx0_p & v8565cf | !jx0_p & v856555;
assign dea6e5 = decide_p & dea6e4 | !decide_p & v84563c;
assign b29f55 = hlock0_p & b29f54 | !hlock0_p & c3bd61;
assign cea19f = hbusreq3 & cea19d | !hbusreq3 & cea19e;
assign a5fc25 = hbusreq3 & a5fc24 | !hbusreq3 & v84563c;
assign ab0747 = hbusreq2_p & ab06e2 | !hbusreq2_p & ab0746;
assign v970432 = hmaster1_p & v84563c | !hmaster1_p & v970431;
assign a5f962 = hbusreq2_p & a5f961 | !hbusreq2_p & a60142;
assign c3bd66 = hgrant2_p & c3bd64 | !hgrant2_p & c3bd65;
assign ab05c6 = hlock2 & ab0511 | !hlock2 & ab05c5;
assign dea729 = hmaster1_p & dea728 | !hmaster1_p & v845660;
assign c3b68d = hbusreq2_p & c3b689 | !hbusreq2_p & c3b687;
assign a5f335 = hmaster0_p & a5f32f | !hmaster0_p & a5f334;
assign deae34 = hbusreq2_p & deae33 | !hbusreq2_p & v845644;
assign c3b70a = hlock2_p & c3b641 | !hlock2_p & !c3b656;
assign ab05bb = hgrant0_p & ab0597 | !hgrant0_p & !ab05ba;
assign a5f0ad = hbusreq2_p & a5f0ab | !hbusreq2_p & a5f0ac;
assign a5edfa = hready & a5edf6 | !hready & v84565a;
assign c3bcda = locked_p & c3bcd9 | !locked_p & c3bc47;
assign af34df = hmaster1_p & af34db | !hmaster1_p & af34de;
assign b29ecf = hbusreq2_p & b29ece | !hbusreq2_p & v84563c;
assign deae95 = hlock0_p & deae94 | !hlock0_p & !v84563c;
assign cea239 = hmaster1_p & v84563c | !hmaster1_p & cea238;
assign a6018a = hlock1_p & v9703fb | !hlock1_p & v84563c;
assign deae5e = hbusreq2_p & deae5d | !hbusreq2_p & deae5c;
assign a5fb91 = locked_p & v84563c | !locked_p & a5fb71;
assign a5eae6 = hlock0_p & a5f249 | !hlock0_p & a5eae4;
assign adaec5 = start_p & a81ca6 | !start_p & v84563c;
assign c3bc8c = hlock0_p & c3bc8a | !hlock0_p & c3bc8b;
assign b2993e = hlock0_p & b2993d | !hlock0_p & !deadb2;
assign dead42 = hbusreq3 & dead41 | !hbusreq3 & !dead3b;
assign adaede = hmaster0_p & v84563c | !hmaster0_p & adaedd;
assign ab05b3 = hbusreq0_p & b2997c | !hbusreq0_p & !b29992;
assign a5ea44 = locked_p & a5fbf0 | !locked_p & a5ea43;
assign a5ee2f = hready & a5ee2b | !hready & !a5ee2e;
assign a5f1dc = hready & a5fba6 | !hready & a5fbae;
assign af3c2d = locked_p & v84563c | !locked_p & v845646;
assign a5f0a1 = hmaster0_p & a5f099 | !hmaster0_p & a5f0a0;
assign a5f3dd = hmaster0_p & a5f3d1 | !hmaster0_p & a5f3dc;
assign ab05e2 = hmaster1_p & ab05e1 | !hmaster1_p & ab0bca;
assign b29f44 = hbusreq2_p & b29f43 | !hbusreq2_p & deacab;
assign v97044b = hmaster1_p & v97044a | !hmaster1_p & v84563c;
assign cea1c5 = hbusreq3 & cea1c4 | !hbusreq3 & v84563c;
assign a5f046 = hbusreq3_p & a5f037 | !hbusreq3_p & a5f045;
assign b29d62 = hmaster1_p & b29d5b | !hmaster1_p & b29d61;
assign ab0b50 = decide_p & ab0b4f | !decide_p & v84563c;
assign c3be01 = hlock0_p & c3be00 | !hlock0_p & c3bcf0;
assign b2669f = start_p & v84563c | !start_p & b2669e;
assign af34b7 = stateG10_1_p & af34b6 | !stateG10_1_p & !af3c4c;
assign c3bdfd = hmaster1_p & c3bdfc | !hmaster1_p & c3bd88;
assign deacbe = hlock1_p & v84565a | !hlock1_p & deacbd;
assign a5eeca = hbusreq2 & a5f3d2 | !hbusreq2 & v845660;
assign ab0caf = hlock2 & ab0cac | !hlock2 & ab0cae;
assign a5ebdd = hbusreq0 & a5ebdc | !hbusreq0 & v84563c;
assign ab0ad6 = hlock0_p & v84563c | !hlock0_p & !b29cc8;
assign b29b28 = hgrant0_p & c3bceb | !hgrant0_p & !b29b27;
assign ab0c97 = hready & ab0c96 | !hready & !v84563c;
assign b29930 = hbusreq2_p & b2991d | !hbusreq2_p & v84563c;
assign dea75f = hbusreq2_p & deae0e | !hbusreq2_p & deae0d;
assign a5eb3c = hmaster1_p & a5eb35 | !hmaster1_p & a5eb3b;
assign b29f99 = locked_p & cea15f | !locked_p & !c3bd98;
assign c3bd2c = hlock1_p & v84563c | !hlock1_p & !deae80;
assign cea3ae = hlock3_p & cea39a | !hlock3_p & cea3ad;
assign a5ede2 = hgrant2_p & a5edde | !hgrant2_p & a5ede1;
assign dea6f9 = hready_p & deac11 | !hready_p & dea6f8;
assign c3bd09 = decide_p & c3bd08 | !decide_p & v845660;
assign cea18a = hmaster0_p & cea187 | !hmaster0_p & cea189;
assign b29fc7 = hmaster1_p & b29fbf | !hmaster1_p & b29fc6;
assign c3bbd4 = hlock0_p & c3bbd1 | !hlock0_p & !c3bbd3;
assign a5ee71 = hlock0_p & a5fbc0 | !hlock0_p & a5ee70;
assign a5edcb = hlock2_p & a5edca | !hlock2_p & a5f546;
assign a5f70f = start_p & v845654 | !start_p & a5f9db;
assign a5ea2d = hmaster1_p & a5ea2c | !hmaster1_p & v84563c;
assign c3b6e8 = hlock2_p & c3b632 | !hlock2_p & !c3b625;
assign a5fc43 = hready & a5fb8a | !hready & v84563c;
assign a5f08b = hlock0_p & a5f2e4 | !hlock0_p & v84563c;
assign a5fc04 = hready & a5f9dd | !hready & v84563c;
assign b29b60 = jx0_p & b29a22 | !jx0_p & b29b5f;
assign b29f95 = hlock0_p & b29ecc | !hlock0_p & c3bcf8;
assign ab05f8 = hgrant2_p & ab05f6 | !hgrant2_p & ab05f7;
assign a5eaf4 = hgrant2_p & a5eaed | !hgrant2_p & a5eaf3;
assign ab0c1d = hlock2_p & ab0c1c | !hlock2_p & v84563c;
assign dea6ca = hlock1_p & deac51 | !hlock1_p & !dea6c9;
assign a5f36d = hlock0_p & a5f367 | !hlock0_p & a5f36c;
assign a60192 = start_p & v845654 | !start_p & !a60185;
assign c3b80a = hlock0_p & c3bd9b | !hlock0_p & cea17a;
assign a5edfd = hbusreq2 & a5edfb | !hbusreq2 & a5edfc;
assign b29f5e = hmaster1_p & b29f4f | !hmaster1_p & !b29f5d;
assign a5f8d4 = hgrant1_p & a5f8d2 | !hgrant1_p & a5f8d3;
assign adaf08 = hgrant2_p & v84563c | !hgrant2_p & adaf07;
assign cea468 = hlock2_p & cea38a | !hlock2_p & cea37b;
assign a5fbbe = hmaster1_p & a5fb85 | !hmaster1_p & a5fbbd;
assign dea6d6 = hbusreq3 & dea6d4 | !hbusreq3 & dea6d5;
assign dea757 = hbusreq2_p & deadef | !hbusreq2_p & deadd6;
assign a5eaf3 = hbusreq3 & a5eaf0 | !hbusreq3 & !a5eaf2;
assign a5fc96 = hmaster1_p & a5fc73 | !hmaster1_p & a5fc95;
assign b29fb6 = hlock0_p & b29fb5 | !hlock0_p & c3bd8e;
assign b2991e = hbusreq2_p & b2991d | !hbusreq2_p & !b2991c;
assign cea41a = hmaster0_p & cea3f3 | !hmaster0_p & cea419;
assign ab0c23 = hbusreq3 & ab0c22 | !hbusreq3 & v84564a;
assign a5fce2 = start_p & a5fc8d | !start_p & !b29f07;
assign af34e8 = hmaster1_p & af3c5e | !hmaster1_p & af34e7;
assign c3b6df = locked_p & c3b6de | !locked_p & c3bbba;
assign a60164 = hburst1_p & c06d34 | !hburst1_p & !v84563c;
assign c3b7f6 = hready & c3b7f5 | !hready & deadb2;
assign ab0b4c = hgrant2_p & ab0b49 | !hgrant2_p & ab0b4b;
assign c3bbf0 = hbusreq3 & c3bbd6 | !hbusreq3 & c3bbef;
assign a6019a = hbusreq2 & a6018c | !hbusreq2 & a60199;
assign c3bdd4 = hlock1_p & v84563c | !hlock1_p & !dea6ce;
assign a81cd7 = hmaster1_p & a81cd6 | !hmaster1_p & v84563c;
assign dead65 = hgrant2_p & deacd3 | !hgrant2_p & dead64;
assign b29f18 = start_p & v84563c | !start_p & b29f17;
assign a5eddc = hlock2_p & a5eddb | !hlock2_p & a5f582;
assign b299a5 = hmaster1_p & b299a4 | !hmaster1_p & b29981;
assign a5ea5a = locked_p & a5ea59 | !locked_p & !v845641;
assign ab0627 = hbusreq2_p & ab0626 | !hbusreq2_p & ab05ee;
assign a5ef47 = hmaster0_p & a5ef46 | !hmaster0_p & !a5f3dc;
assign a5fb9a = hbusreq2 & a5fb96 | !hbusreq2 & a5fb99;
assign ab057c = hgrant2_p & ab0566 | !hgrant2_p & ab057b;
assign b29f17 = stateA1_p & v8c6449 | !stateA1_p & v84563c;
assign a5eeba = hbusreq1 & a5eeb9 | !hbusreq1 & !v84563c;
assign ce9e22 = hbusreq2_p & cea286 | !hbusreq2_p & ce9e21;
assign ab0cb3 = hmaster0_p & ab0ca9 | !hmaster0_p & ab0cb2;
assign a5ee53 = hlock1_p & a5fba2 | !hlock1_p & !a5ee52;
assign a5ea91 = hbusreq0 & a5ea90 | !hbusreq0 & v84563c;
assign b29f88 = hbusreq2_p & b29f87 | !hbusreq2_p & v84563c;
assign a5fcfe = hlock1_p & v84563c | !hlock1_p & b29918;
assign dea74d = hbusreq2_p & deadd2 | !hbusreq2_p & deadd1;
assign ab0c87 = hbusreq2_p & ab0c86 | !hbusreq2_p & ab0b5f;
assign a5ec1e = hmaster1_p & a5f92d | !hmaster1_p & a5ea1b;
assign b29d2e = hlock2 & b29cdf | !hlock2 & deadb2;
assign a5f3b7 = hbusreq3 & a5f3b6 | !hbusreq3 & v845641;
assign a5f541 = hlock0_p & a5f36e | !hlock0_p & a5f540;
assign ab0c13 = hbusreq0_p & b266a8 | !hbusreq0_p & c3bcf0;
assign a5f537 = hlock0_p & a5f52c | !hlock0_p & !a5f536;
assign a5edda = hready & a5f57c | !hready & a5edd9;
assign c3b777 = hready_p & c3bbc1 | !hready_p & c3b776;
assign dea6f5 = hmaster1_p & deadea | !hmaster1_p & dea6f4;
assign cea348 = decide_p & cea347 | !decide_p & v84563c;
assign a5f1ea = hbusreq0 & a5f1db | !hbusreq0 & !a5f1e9;
assign b29d53 = hlock0_p & b29d52 | !hlock0_p & v84563c;
assign b299cc = decide_p & b299cb | !decide_p & v84563c;
assign dea75b = hlock3_p & dea74a | !hlock3_p & dea75a;
assign b29ffb = hready_p & b29ff2 | !hready_p & b29ffa;
assign a5ea56 = hlock2 & a5ea4f | !hlock2 & a5ea55;
assign a9b9e9 = hgrant0_p & a9b9e3 | !hgrant0_p & a9b9e8;
assign c3b7a3 = hbusreq3 & c3b7a2 | !hbusreq3 & cea15a;
assign dea79c = decide_p & dea79b | !decide_p & !v84563c;
assign a5f98f = locked_p & a5f974 | !locked_p & v845641;
assign c3b722 = hbusreq2_p & c3b721 | !hbusreq2_p & !c3b71f;
assign v970443 = hmaster0_p & v84563c | !hmaster0_p & v970442;
assign c3bd7b = hlock0_p & c3bd7a | !hlock0_p & c3bd61;
assign c3bc10 = hgrant2_p & c3bc07 | !hgrant2_p & c3bc0f;
assign a5f74d = hbusreq2 & a5fc89 | !hbusreq2 & !v84563c;
assign c3bdc8 = hgrant2_p & dead3e | !hgrant2_p & c3bdc7;
assign a5f301 = hmaster0_p & a5f300 | !hmaster0_p & a5f210;
assign a5f8e3 = hgrant1_p & a5f8e1 | !hgrant1_p & a5f8e2;
assign a60177 = hmastlock_p & a60176 | !hmastlock_p & v84563c;
assign c3bd10 = hburst0 & cea24d | !hburst0 & c3bd0f;
assign deadda = hbusreq2_p & deadd7 | !hbusreq2_p & v84563c;
assign a5ea4c = locked_p & a5fbfb | !locked_p & a5fb6a;
assign a5ea14 = hlock2 & a5ea12 | !hlock2 & a5ea13;
assign b29ab2 = hlock0_p & c3bd8d | !hlock0_p & !v84563c;
assign ab05fe = hgrant2_p & ab05fb | !hgrant2_p & ab05fd;
assign b299e9 = hready_p & b299e6 | !hready_p & b299e8;
assign cea45e = hgrant0_p & cea451 | !hgrant0_p & cea45d;
assign a5fbaa = start_p & a81ca6 | !start_p & a5fba9;
assign a5f6cf = decide_p & a5f6ce | !decide_p & v84563c;
assign a5fc48 = hmastlock_p & a5fc47 | !hmastlock_p & v84563c;
assign b29b1b = hready_p & b29b12 | !hready_p & b29b1a;
assign dead36 = hbusreq3 & dead35 | !hbusreq3 & !dead2d;
assign a5fb1b = stateG10_1_p & v970407 | !stateG10_1_p & a60186;
assign cea48c = hmaster0_p & cea48b | !hmaster0_p & cea419;
assign ab0cbb = hlock3_p & ab0ca6 | !hlock3_p & ab0cba;
assign deae49 = hready_p & deae3e | !hready_p & deae48;
assign cea394 = hlock0_p & cea389 | !hlock0_p & cea393;
assign deadb5 = hbusreq2_p & deadb4 | !hbusreq2_p & v84565a;
assign deae47 = hmaster0_p & deae43 | !hmaster0_p & !deae46;
assign ce9ddd = hready_p & ce9dbb | !hready_p & ce9ddc;
assign a5f3d1 = hmaster1_p & a5f3d0 | !hmaster1_p & v84563c;
assign deac5c = hlock0_p & deac57 | !hlock0_p & deac5b;
assign bdb5a0 = hmaster0_p & c3bca4 | !hmaster0_p & bdb59f;
assign a5f807 = hlock0_p & a5f7fd | !hlock0_p & !a5f806;
assign a5f174 = hbusreq1_p & a60168 | !hbusreq1_p & a5fb8b;
assign dea743 = hbusreq2_p & deadc6 | !hbusreq2_p & !deadc4;
assign b29d82 = hready & b26695 | !hready & !v84563c;
assign c3b7ab = hlock0_p & c3bcf8 | !hlock0_p & v84563c;
assign a5eb2b = hbusreq0 & a5eb2a | !hbusreq0 & v84563c;
assign a5eed0 = hgrant2_p & a5eecf | !hgrant2_p & v84563c;
assign be34e9 = hready_p & be34e7 | !hready_p & be34e8;
assign a5f2f4 = hready & v84563c | !hready & !dead18;
assign a5f8c6 = hlock0_p & a5f8c4 | !hlock0_p & a5f8c5;
assign d40d46 = hbusreq2_p & d40d44 | !hbusreq2_p & d40d43;
assign a81cfb = hbusreq2_p & a81cc8 | !hbusreq2_p & a81cf1;
assign a5faea = hmaster1_p & a5fa71 | !hmaster1_p & a5fae9;
assign b29f60 = hlock2_p & c3bd5f | !hlock2_p & !v84563c;
assign ab0c63 = hgrant2_p & ab0c61 | !hgrant2_p & ab0c62;
assign a5eea3 = hlock1_p & a5fc0d | !hlock1_p & !a5ee55;
assign v97043e = hmastlock_p & v97043d | !hmastlock_p & v84563c;
assign deadbe = hlock1_p & v84565a | !hlock1_p & !deadbd;
assign bdb5b7 = decide_p & bdb5b6 | !decide_p & bdb5aa;
assign deae6f = hlock3_p & deae58 | !hlock3_p & deae6e;
assign b29ea7 = hlock0_p & b29ea6 | !hlock0_p & c3bcf8;
assign c3bc57 = hmaster1_p & c3bc4b | !hmaster1_p & c3bc56;
assign c3b655 = hbusreq0_p & c3b625 | !hbusreq0_p & !c3b635;
assign cea473 = hmaster1_p & cea46f | !hmaster1_p & cea472;
assign ab06e6 = locked_p & b29fb4 | !locked_p & !c3bc47;
assign dead6f = hbusreq1_p & dead6e | !hbusreq1_p & !deacf7;
assign cea2f2 = hlock0_p & cea2f1 | !hlock0_p & !dead72;
assign a5e9d0 = hmaster0_p & a5f164 | !hmaster0_p & a5e9cf;
assign ab0cda = hbusreq2_p & ab0c27 | !hbusreq2_p & v845644;
assign a5f576 = hbusreq0_p & a5f36e | !hbusreq0_p & a5f540;
assign af3488 = hmaster1_p & af3c7b | !hmaster1_p & af3487;
assign a5f4b8 = hready & a5f4a6 | !hready & a5f493;
assign ab0b2e = hbusreq3 & ab0b19 | !hbusreq3 & ab0b2d;
assign c3bc20 = hlock0_p & c3bc03 | !hlock0_p & !v84563c;
assign ab0605 = hmaster1_p & ab0604 | !hmaster1_p & ab0b61;
assign a5f952 = hbusreq2 & a5fcd2 | !hbusreq2 & v84563c;
assign a5e9db = hbusreq0 & a5e9da | !hbusreq0 & v845641;
assign a5f2d6 = hmaster0_p & a5f2ca | !hmaster0_p & a5f2d5;
assign a5fd38 = hmaster1_p & a5fd28 | !hmaster1_p & a5fd37;
assign c3bd3b = hlock1_p & c3bd37 | !hlock1_p & c3bd3a;
assign ab0cde = decide_p & ab0cdd | !decide_p & v84563c;
assign deae0e = hlock2_p & deae0d | !hlock2_p & v84563c;
assign b29ec0 = hlock0_p & dead7f | !hlock0_p & !b29eae;
assign c3b773 = hmaster1_p & deac3f | !hmaster1_p & c3bccf;
assign b266bf = hlock3_p & b266b7 | !hlock3_p & b266be;
assign a5f03d = hready_p & v84563c | !hready_p & a5f03c;
assign ab0c9d = hlock2 & ab0c99 | !hlock2 & ab0c9c;
assign c3b6ee = hgrant2_p & c3b6ed | !hgrant2_p & c3bc70;
assign b29aae = locked_p & cea151 | !locked_p & !v84563c;
assign a5f292 = hbusreq2 & a5f728 | !hbusreq2 & a5f291;
assign a5efdc = hmaster1_p & a5efdb | !hmaster1_p & a5f6d9;
assign af3547 = hgrant1_p & af3546 | !hgrant1_p & v84563c;
assign b29d02 = hlock2 & b29cff | !hlock2 & b29d01;
assign a5f957 = hbusreq2 & a5fcc8 | !hbusreq2 & v84563c;
assign ab069b = hbusreq2_p & ab069a | !hbusreq2_p & ab0699;
assign cea184 = hgrant3_p & cea0f4 | !hgrant3_p & cea183;
assign a5eedb = hlock0_p & a5eeda | !hlock0_p & a5f560;
assign b29ae7 = hbusreq2_p & b29ae4 | !hbusreq2_p & v84563c;
assign c3bbf1 = hbusreq2_p & c3bbd5 | !hbusreq2_p & c3bbd4;
assign cea162 = hlock0_p & cea161 | !hlock0_p & !dead72;
assign af3c4f = locked_p & af3c49 | !locked_p & af3c4e;
assign a5f13c = hbusreq3 & a5f139 | !hbusreq3 & !a5f13b;
assign c3bc28 = hbusreq2_p & c3bc22 | !hbusreq2_p & c3bc21;
assign cea15c = hbusreq2_p & cea15b | !hbusreq2_p & cea15a;
assign a5f329 = hlock2_p & a5f328 | !hlock2_p & v84563c;
assign a5f07f = hlock0_p & a5fbc7 | !hlock0_p & v84563c;
assign dea786 = hbusreq2_p & deae1f | !hbusreq2_p & deae1e;
assign c3bd21 = hready & c3bbfb | !hready & deadb2;
assign a5ee4c = hready & a5f365 | !hready & a5ee4b;
assign ab0579 = hbusreq3 & ab0561 | !hbusreq3 & ab0564;
assign b2676a = hmaster1_p & b26715 | !hmaster1_p & !b266a2;
assign af3564 = hbusreq2_p & af355f | !hbusreq2_p & af3563;
assign a5f8df = start_p & a5f8de | !start_p & a5f8db;
assign a5fa68 = hbusreq2 & a5fa60 | !hbusreq2 & !a5fa67;
assign c3bca9 = hbusreq2_p & c3bca8 | !hbusreq2_p & v84563c;
assign d40d7e = hmaster1_p & d40d60 | !hmaster1_p & d40d7d;
assign c3bc45 = decide_p & c3bc44 | !decide_p & v845660;
assign a5edbb = hlock2_p & a5edba | !hlock2_p & a5f4f2;
assign ab0bc7 = decide_p & ab0b4f | !decide_p & !v845662;
assign ab0ade = hlock0_p & v84563c | !hlock0_p & deacaa;
assign b298a4 = locked_p & v84563c | !locked_p & b29832;
assign cea14f = hbusreq3 & cea14e | !hbusreq3 & cea85f;
assign a5efbe = hbusreq0_p & a5ee38 | !hbusreq0_p & a5efae;
assign c3bd82 = hready_p & c3bd09 | !hready_p & c3bd81;
assign dea763 = hgrant2_p & dea761 | !hgrant2_p & dea762;
assign cea3e9 = hlock1_p & v84563c | !hlock1_p & !cea271;
assign a5fb81 = hlock1_p & v84563c | !hlock1_p & a5fb80;
assign cea2b2 = hmaster1_p & cea2a8 | !hmaster1_p & cea2b1;
assign a81cf9 = hgrant2_p & v84563c | !hgrant2_p & a81cf8;
assign adaee2 = hmaster1_p & v84563c | !hmaster1_p & adaee1;
assign af34cf = hbusreq2_p & af349d | !hbusreq2_p & af3c4c;
assign a5f546 = hbusreq2 & a5f542 | !hbusreq2 & a5f545;
assign ab0540 = hlock2_p & ab053e | !hlock2_p & ab053f;
assign a5f8f6 = hgrant2_p & a5f8f2 | !hgrant2_p & a5f8f5;
assign c3b6b2 = hlock2_p & c3b6b0 | !hlock2_p & !c3b6b1;
assign cea485 = hbusreq2_p & cea484 | !hbusreq2_p & cea3ea;
assign a5f82a = hgrant1_p & a5f829 | !hgrant1_p & a5f828;
assign af3c55 = hlock1_p & d40d33 | !hlock1_p & af3c54;
assign ce9d2d = hgrant2_p & cea25b | !hgrant2_p & ce9d2c;
assign a5f372 = hlock2_p & a5f36d | !hlock2_p & a5f371;
assign ab0b11 = hgrant2_p & ab0b04 | !hgrant2_p & ab0b10;
assign ab0c2a = hmaster1_p & v84563c | !hmaster1_p & ab0c29;
assign c3b6f3 = hmaster0_p & c3b6eb | !hmaster0_p & c3b6f2;
assign dead9d = hmaster1_p & v84563c | !hmaster1_p & dead9c;
assign a5ea38 = hgrant2_p & a5ea35 | !hgrant2_p & a5ea37;
assign ab0cfa = hbusreq2_p & ab0c60 | !hbusreq2_p & b29cbb;
assign ab069e = hbusreq2_p & ab069a | !hbusreq2_p & ab0692;
assign af34d3 = hbusreq2_p & af34d2 | !hbusreq2_p & af3c4c;
assign a5fa61 = hgrant1_p & a60187 | !hgrant1_p & a5fa0f;
assign cea326 = hlock0_p & cea325 | !hlock0_p & !dead72;
assign a5f098 = hbusreq3 & a5f097 | !hbusreq3 & v84563c;
assign a5fb70 = start_p & v84563c | !start_p & a5fb6f;
assign c3b806 = hgrant2_p & c3b804 | !hgrant2_p & c3b805;
assign cea410 = hbusreq2_p & cea40d | !hbusreq2_p & !cea40f;
assign a5fc84 = hmastlock_p & a5fc83 | !hmastlock_p & !v84563c;
assign cea3ea = hready & cea3e8 | !hready & cea3e9;
assign c3b6a1 = hready & c3b6a0 | !hready & v84563c;
assign af3511 = jx1_p & af3c47 | !jx1_p & !af3510;
assign af34bf = hgrant2_p & af34b4 | !hgrant2_p & af34be;
assign a5f527 = hlock2 & a5f51c | !hlock2 & a5f526;
assign a5f486 = stateG10_1_p & v84563c | !stateG10_1_p & a5f485;
assign cea0d3 = hbusreq2_p & cea0b9 | !hbusreq2_p & cea0b8;
assign c3bca2 = hmaster1_p & dead2e | !hmaster1_p & !c3bca1;
assign c3bd16 = hlock1_p & v84563c | !hlock1_p & !deae75;
assign adaed4 = hmaster1_p & v84563c | !hmaster1_p & adaeca;
assign c3b6fd = hbusreq2_p & c3b6fc | !hbusreq2_p & c3b6fb;
assign b29ea2 = hready_p & b29e98 | !hready_p & b29ea1;
assign c3bdbf = locked_p & c3bdbe | !locked_p & !c3bd9a;
assign b29a4a = hlock2_p & v84563c | !hlock2_p & !dead2e;
assign dea6c0 = hgrant2_p & dea6bf | !hgrant2_p & dead3b;
assign b29a43 = hbusreq3 & b29a42 | !hbusreq3 & v84563c;
assign ce9cfc = hmaster1_p & ce9cfb | !hmaster1_p & cea860;
assign b29fdb = hlock0_p & b29fd9 | !hlock0_p & b29fda;
assign cea417 = hbusreq2_p & cea415 | !hbusreq2_p & cea413;
assign a5fbca = hbusreq2 & a5fbc9 | !hbusreq2 & a5fbc8;
assign a6016c = hburst0_p & c06d34 | !hburst0_p & a6016b;
assign a5ee39 = locked_p & v84563c | !locked_p & a5ee38;
assign a5f97c = hburst1_p & v845672 | !hburst1_p & d615cf;
assign a5fc50 = start_p & v8e1935 | !start_p & !a5fc4f;
assign cea29c = hmaster0_p & cea28a | !hmaster0_p & cea29b;
assign ab0c59 = hbusreq1_p & c3b660 | !hbusreq1_p & !v84565a;
assign a5ef85 = hbusreq2_p & a5edd6 | !hbusreq2_p & a5ef84;
assign cea49e = hbusreq2_p & cea49b | !hbusreq2_p & cea405;
assign dea6fc = decide_p & dea6fb | !decide_p & v84563c;
assign a5ef08 = hbusreq1_p & a5fcd7 | !hbusreq1_p & !v84563c;
assign a5f598 = hbusreq3 & a5f596 | !hbusreq3 & a5f597;
assign ab0754 = hbusreq2_p & ab06b5 | !hbusreq2_p & !ab06c1;
assign a5eea5 = hready & a5eea2 | !hready & a5eea4;
assign dead7b = hmastlock_p & dead7a | !hmastlock_p & !v84563c;
assign a5eb45 = hmaster0_p & a5eb3c | !hmaster0_p & a5eb44;
assign a5f304 = hmaster0_p & a5f303 | !hmaster0_p & a5f218;
assign ce9d35 = hbusreq2_p & cea2b0 | !hbusreq2_p & cea2af;
assign ce9cca = hmaster1_p & ce9cc9 | !hmaster1_p & cea1a1;
assign ab0c6a = hlock2 & ab0af2 | !hlock2 & ab0c69;
assign c3bc95 = hlock2_p & c3bc94 | !hlock2_p & !v84563c;
assign a5f164 = hmaster1_p & a5f13d | !hmaster1_p & a5f163;
assign c3b79d = hlock2_p & c3b79b | !hlock2_p & !c3b79c;
assign a5f566 = hlock0_p & a5f565 | !hlock0_p & a5f55b;
assign cea287 = hbusreq2_p & cea286 | !hbusreq2_p & deacaa;
assign b29992 = hready & deae67 | !hready & v84563c;
assign a5f1f7 = locked_p & v84563c | !locked_p & a5f1f6;
assign a5f4e8 = hlock1_p & a5fa1c | !hlock1_p & a5f4e7;
assign a5f1d5 = hlock2 & a5f1cf | !hlock2 & a5f1d4;
assign a5f01b = hmaster1_p & v84563c | !hmaster1_p & a5f6d9;
assign c3b614 = hlock0_p & c3b613 | !hlock0_p & !c3bd60;
assign deadef = hlock2_p & deadee | !hlock2_p & !v84563c;
assign ab06a4 = hlock2_p & ab06a2 | !hlock2_p & ab06a3;
assign af3c6b = locked_p & af3c6a | !locked_p & af3c4c;
assign a5fb1e = hgrant1_p & a5fa12 | !hgrant1_p & v9703fb;
assign deac62 = hbusreq3 & deac61 | !hbusreq3 & v84563c;
assign a5fc55 = hready & a5fc53 | !hready & a5fc54;
assign cea441 = decide_p & cea440 | !decide_p & v84563c;
assign a5fc66 = hgrant0_p & a5fc4e | !hgrant0_p & a5fc65;
assign deae20 = hbusreq2_p & deae1f | !hbusreq2_p & v84565a;
assign cea356 = decide_p & cea355 | !decide_p & v84563c;
assign ab0c60 = hlock2_p & ab0c5f | !hlock2_p & !c3bc3c;
assign ab0570 = hbusreq0_p & b29942 | !hbusreq0_p & b29947;
assign a5eb84 = hbusreq0 & a5eb3e | !hbusreq0 & !v84563c;
assign ab0c7f = hmaster0_p & ab0c70 | !hmaster0_p & ab0c7e;
assign af358e = hmaster1_p & af358d | !hmaster1_p & af3533;
assign dead6a = hgrant3_p & dead69 | !hgrant3_p & !v84563c;
assign ab0528 = hlock0_p & v84563c | !hlock0_p & !cea37b;
assign deac9a = hbusreq3 & deac99 | !hbusreq3 & v84563c;
assign ab0c90 = hmaster1_p & ab0b61 | !hmaster1_p & ab0c8f;
assign c3b619 = hbusreq3 & c3b617 | !hbusreq3 & c3b618;
assign a5eec2 = hbusreq1 & a5eec1 | !hbusreq1 & !v84563c;
assign ab0bee = hgrant2_p & ab0ae0 | !hgrant2_p & ab0ae2;
assign a5f3a7 = hbusreq2_p & a5f3a6 | !hbusreq2_p & a5f3a2;
assign dea7a7 = hgrant2_p & deae40 | !hgrant2_p & dea74e;
assign cea176 = hmaster0_p & cea167 | !hmaster0_p & cea175;
assign b299e0 = hlock2_p & v845660 | !hlock2_p & !b299df;
assign c3b874 = hbusreq3 & c3b812 | !hbusreq3 & dead39;
assign ab062f = hbusreq3 & ab062c | !hbusreq3 & ab062e;
assign af35ab = hmaster0_p & af35aa | !hmaster0_p & af357c;
assign d40d29 = stateG2_p & v84563c | !stateG2_p & !c06d34;
assign a5f55c = hlock0_p & a5f55a | !hlock0_p & a5f55b;
assign a5eee2 = hbusreq1 & a5eee1 | !hbusreq1 & !v84563c;
assign a5edef = hbusreq1_p & a5fcdd | !hbusreq1_p & !v84563c;
assign c3b727 = hgrant2_p & c3b723 | !hgrant2_p & c3b726;
assign a5e9c9 = hlock0_p & a5f320 | !hlock0_p & v84563c;
assign a5efb4 = hgrant2_p & a5efb3 | !hgrant2_p & v84563c;
assign a5f456 = hlock1_p & a5f455 | !hlock1_p & a5f436;
assign a5f9a1 = locked_p & a5fbdb | !locked_p & a5f9a0;
assign b29925 = hgrant1_p & b29924 | !hgrant1_p & b29923;
assign ab0520 = hmaster0_p & ab050f | !hmaster0_p & ab051f;
assign c3b61c = hmaster0_p & c3b61b | !hmaster0_p & c3bd67;
assign deadca = hbusreq3 & deadc9 | !hbusreq3 & deadc7;
assign c3bcc4 = decide_p & c3bcc3 | !decide_p & v845660;
assign a5ea8a = hgrant2_p & a5ea87 | !hgrant2_p & a5ea89;
assign b299a7 = hgrant0_p & b2997b | !hgrant0_p & !b299a6;
assign dea7a0 = hbusreq3 & dea79f | !hbusreq3 & dea72e;
assign ce9da6 = decide_p & ce9da5 | !decide_p & a57859;
assign a5e9cc = hbusreq0 & a5e9ca | !hbusreq0 & a5e9ad;
assign b29cca = hlock2_p & v84563c | !hlock2_p & !b29cc9;
assign c3bd8e = hbusreq0_p & c3bcf8 | !hbusreq0_p & c3bd8d;
assign a5f733 = hlock2_p & a5f726 | !hlock2_p & v84563c;
assign b26707 = hlock3_p & b26701 | !hlock3_p & b26706;
assign a5f189 = hlock1_p & a5fbab | !hlock1_p & !a5f188;
assign a5f717 = hlock2 & a5f70b | !hlock2 & a5f716;
assign cea3fc = hlock2_p & cea3f9 | !hlock2_p & cea3fb;
assign a5fb7c = hlock2_p & a5fb7b | !hlock2_p & v84563c;
assign deadfd = hlock0_p & deadfc | !hlock0_p & v84563c;
assign a5f974 = hready & v84563c | !hready & a5f973;
assign c3b829 = hlock0_p & c3bcf0 | !hlock0_p & v845660;
assign a5f93c = hlock2_p & a5f93b | !hlock2_p & a5f8cb;
assign a5f8bc = hbusreq1_p & v84565a | !hbusreq1_p & !deaca1;
assign a5fab4 = hlock2_p & a5fab1 | !hlock2_p & !a5fab3;
assign ab0675 = hlock2_p & ab0b80 | !hlock2_p & ab0674;
assign deaddb = hbusreq3 & deadd9 | !hbusreq3 & deadda;
assign c3b6c7 = hlock0_p & c3b6c6 | !hlock0_p & c3b6a8;
assign cea452 = hlock2_p & cea38b | !hlock2_p & cea37b;
assign c3b82e = hgrant0_p & dead2e | !hgrant0_p & c3b82d;
assign c3bde4 = hlock2_p & c3bd8d | !hlock2_p & v84563c;
assign deacfd = hlock0_p & deacfa | !hlock0_p & deacfc;
assign a5ee27 = locked_p & v845646 | !locked_p & a5ee26;
assign ce9cf7 = hbusreq3 & ce9cf5 | !hbusreq3 & ce9cf6;
assign ab0583 = hmaster1_p & ab057c | !hmaster1_p & ab0582;
assign a5f4a4 = hgrant1_p & a5f4a3 | !hgrant1_p & a5f4a2;
assign deae29 = hgrant2_p & deae26 | !hgrant2_p & deae28;
assign a9b9d2 = hmaster0_p & a9b9d1 | !hmaster0_p & !v84563c;
assign a5fc8e = start_p & a5fc8d | !start_p & b29eb3;
assign ab06ae = hgrant1_p & ab06ad | !hgrant1_p & deaca0;
assign dead0f = hlock2_p & dead0e | !hlock2_p & dead0d;
assign ce9cc0 = hlock0_p & ce9cbf | !hlock0_p & !cea405;
assign a5ef58 = hlock0_p & a5f540 | !hlock0_p & a5f4fc;
assign a5f726 = locked_p & v84563c | !locked_p & a5f6e9;
assign ab0601 = decide_p & ab0600 | !decide_p & v84563c;
assign c3b826 = hlock0_p & c3b825 | !hlock0_p & !dead77;
assign deac7b = hlock0_p & deac7a | !hlock0_p & !v84565a;
assign ce9cc7 = hbusreq2_p & ce9cc3 | !hbusreq2_p & cea40f;
assign cea89e = hbusreq2_p & cea89d | !hbusreq2_p & deacaa;
assign deac5b = hlock1_p & deac52 | !hlock1_p & deac5a;
assign b29d5b = hbusreq3 & b29d5a | !hbusreq3 & c3bceb;
assign ab0bcc = hmaster0_p & ab0bcb | !hmaster0_p & ab0bca;
assign b29d98 = hgrant2_p & b29d97 | !hgrant2_p & !b29d90;
assign c3bd5b = hgrant1_p & c3bd11 | !hgrant1_p & c3bd13;
assign c3b637 = hlock0_p & c3bbbb | !hlock0_p & c3b636;
assign a5f370 = hlock0_p & a5f36f | !hlock0_p & a5f36c;
assign af34c4 = hgrant2_p & af34c2 | !hgrant2_p & af34c3;
assign a5f8ba = hbusreq0_p & a5f8b9 | !hbusreq0_p & ab0c31;
assign cea384 = hlock0_p & cea381 | !hlock0_p & cea383;
assign a5f041 = hmaster1_p & a5f6db | !hmaster1_p & a5f040;
assign b29b31 = hmaster1_p & b29a89 | !hmaster1_p & !b29e6e;
assign d40d54 = hlock0_p & d40d31 | !hlock0_p & d40d33;
assign a5fc82 = stateA1_p & a5fb9d | !stateA1_p & d615cf;
assign a5f908 = hlock0_p & a5fb2a | !hlock0_p & ab0c31;
assign cea26d = hbusreq1_p & cea26b | !hbusreq1_p & v84563c;
assign a5efc9 = hbusreq2 & a5f3d8 | !hbusreq2 & v845660;
assign cea37c = locked_p & cea37a | !locked_p & cea37b;
assign a5eb4f = hbusreq0 & a5ea9b | !hbusreq0 & !v84563c;
assign a5f4d0 = hbusreq1 & a5f4cf | !hbusreq1 & !v84563c;
assign dead96 = hbusreq2_p & dead95 | !hbusreq2_p & v84563c;
assign a5f209 = hbusreq2_p & a5f208 | !hbusreq2_p & v84563c;
assign ab0ce7 = hlock2_p & ab0ce6 | !hlock2_p & dead2e;
assign a5f993 = hlock2 & a5fc4a | !hlock2 & a5f992;
assign cea259 = hlock0_p & cea258 | !hlock0_p & v84563c;
assign ab06d0 = hlock0_p & b29f79 | !hlock0_p & !ab06b7;
assign a5f3c7 = hbusreq1 & a5f3c6 | !hbusreq1 & v84563c;
assign a5f2c8 = hlock2_p & a5f2c7 | !hlock2_p & v84563c;
assign a5f1d3 = locked_p & a5f1d2 | !locked_p & v845641;
assign c3b72d = hgrant3_p & c3b6d5 | !hgrant3_p & c3b72c;
assign ce9ccc = decide_p & ce9ccb | !decide_p & !a57859;
assign dead21 = hlock0_p & b26695 | !hlock0_p & dead20;
assign a5ea73 = hbusreq2_p & a5f080 | !hbusreq2_p & a5ea39;
assign dead76 = hmastlock_p & dead75 | !hmastlock_p & !v84563c;
assign b29ac0 = hlock2_p & b29abf | !hlock2_p & b29d81;
assign a5f283 = hbusreq2 & a5fd00 | !hbusreq2 & v84563c;
assign a81d04 = hmaster0_p & a81d03 | !hmaster0_p & v84563c;
assign a5ead7 = hbusreq2_p & a5ead6 | !hbusreq2_p & a5ead5;
assign cea85f = hbusreq2_p & cea85e | !hbusreq2_p & cea85d;
assign b29e95 = hbusreq2_p & dead2c | !hbusreq2_p & v845644;
assign v9703fd = locked_p & v9703fc | !locked_p & v84563c;
assign ab0b57 = hlock2_p & ab0b56 | !hlock2_p & dead2e;
assign af35b3 = decide_p & af35ae | !decide_p & af35b2;
assign b26762 = hgrant2_p & b26761 | !hgrant2_p & !b266c1;
assign a5fa57 = hbusreq2_p & a5fa56 | !hbusreq2_p & v84563c;
assign b29e5b = hgrant3_p & b29d50 | !hgrant3_p & b29e5a;
assign a5ea29 = hbusreq2 & a5ea27 | !hbusreq2 & a5ea28;
assign a5fae3 = hbusreq3 & a5fabc | !hbusreq3 & a5fae2;
assign a5f491 = hlock1_p & a5f9dd | !hlock1_p & a5f490;
assign a81cc9 = hmaster1_p & a81cc8 | !hmaster1_p & v84563c;
assign a5efe4 = hbusreq2_p & a5f583 | !hbusreq2_p & !a5ef86;
assign a5f379 = hbusreq1 & a5f378 | !hbusreq1 & !v84563c;
assign a5f252 = hlock2_p & a5f24b | !hlock2_p & !a5f251;
assign ab0bbd = hbusreq3 & v84563c | !hbusreq3 & cea15a;
assign af35bf = decide_p & af35b9 | !decide_p & af35be;
assign a5fbe3 = hbusreq1 & a5fbd7 | !hbusreq1 & a5fbe2;
assign a5f8cc = hlock2_p & a5f8c7 | !hlock2_p & a5f8cb;
assign ab0518 = hbusreq3 & ab0514 | !hbusreq3 & ab0517;
assign a5efb0 = hlock0_p & a5ee65 | !hlock0_p & a5efaf;
assign a5ef87 = hbusreq2_p & a5eddc | !hbusreq2_p & a5ef86;
assign bdb58d = hgrant2_p & v84565a | !hgrant2_p & bdb58c;
assign cea32d = hgrant0_p & cea31c | !hgrant0_p & cea32c;
assign v84565a = hmastlock_p & v84563c | !hmastlock_p & !v84563c;
assign a5f87c = hbusreq1 & a60167 | !hbusreq1 & a60192;
assign c3b62c = hlock0_p & c3b62a | !hlock0_p & !c3b62b;
assign cea475 = hgrant0_p & cea467 | !hgrant0_p & cea474;
assign dead3c = hgrant2_p & dead39 | !hgrant2_p & dead3b;
assign cea28a = hmaster1_p & cea27b | !hmaster1_p & !cea289;
assign a5f568 = hlock2_p & a5f55c | !hlock2_p & a5f567;
assign c3b819 = hgrant0_p & c3bc5e | !hgrant0_p & c3b818;
assign a5e9f6 = hlock0_p & a5fa00 | !hlock0_p & a5f17c;
assign a5f841 = hgrant1_p & a5f840 | !hgrant1_p & a5f83f;
assign c3b6fb = hlock0_p & c3b6fa | !hlock0_p & !c3b6e1;
assign c3bdc3 = hgrant2_p & dead3e | !hgrant2_p & c3bdc2;
assign a5f198 = hlock0_p & ab0c31 | !hlock0_p & v84563c;
assign a5f901 = hlock0_p & a5f900 | !hlock0_p & v84563c;
assign b29d8f = hbusreq3 & b29d8e | !hbusreq3 & c3bcfb;
assign b2a01c = hbusreq3_p & b29feb | !hbusreq3_p & b2a01b;
assign c3bd68 = hmaster0_p & c3bd51 | !hmaster0_p & c3bd67;
assign cea454 = hgrant2_p & cea453 | !hgrant2_p & !cea15c;
assign a5f067 = hbusreq0_p & a5fc44 | !hbusreq0_p & a5f066;
assign a5f9e9 = hlock0_p & a5f9e1 | !hlock0_p & a5f9e8;
assign cea299 = hbusreq2_p & cea297 | !hbusreq2_p & cea86c;
assign ab0603 = hlock2_p & ab058d | !hlock2_p & ab05bd;
assign a5fc22 = locked_p & v84563c | !locked_p & a5fc21;
assign c3b894 = hmaster0_p & c3b893 | !hmaster0_p & c3b817;
assign b29d85 = hlock2 & b29d81 | !hlock2 & b29d84;
assign dead4d = hgrant0_p & dead38 | !hgrant0_p & dead4c;
assign dead25 = hlock0_p & dead24 | !hlock0_p & deacfc;
assign a5fb8f = hready & a5fb8a | !hready & a5fb8e;
assign b26697 = hlock1_p & v84563c | !hlock1_p & !b26696;
assign a5f710 = hmastlock_p & a5f70f | !hmastlock_p & v84563c;
assign af35a7 = hmaster0_p & af35a6 | !hmaster0_p & af356c;
assign deac6a = hbusreq1_p & deac52 | !hbusreq1_p & deac51;
assign a5fa5c = hlock0_p & a5fa5a | !hlock0_p & a5fa5b;
assign a5f144 = hbusreq0_p & a5fafd | !hbusreq0_p & v84563c;
assign a5f3f6 = hgrant1_p & a5f3f5 | !hgrant1_p & v84563c;
assign cea0e8 = hmaster1_p & v84563c | !hmaster1_p & cea0e7;
assign a5f15d = hlock2_p & a5f154 | !hlock2_p & a5f15c;
assign b29967 = hlock0_p & b29966 | !hlock0_p & b29cdf;
assign ab0b6f = hlock2_p & ab0acb | !hlock2_p & v84563c;
assign c3b725 = hbusreq2_p & c3b721 | !hbusreq2_p & c3b720;
assign a5f745 = hlock2_p & a5f744 | !hlock2_p & v84563c;
assign af34f8 = hmaster0_p & af34f5 | !hmaster0_p & af34f7;
assign cea1a6 = decide_p & cea1a5 | !decide_p & !a57859;
assign a60178 = hbusreq1 & a60173 | !hbusreq1 & !a60177;
assign dea7ac = hready_p & dea7a6 | !hready_p & dea7ab;
assign a5f1b8 = hgrant2_p & a5fbc4 | !hgrant2_p & a5f1b7;
assign cea247 = hburst1 & cea246 | !hburst1 & deacb3;
assign b299d2 = hgrant2_p & b299cf | !hgrant2_p & b299d1;
assign a5f0eb = hlock0_p & ab0c31 | !hlock0_p & a5f0e5;
assign ab0be3 = hgrant2_p & ab0be2 | !hgrant2_p & cea15a;
assign d40d99 = hmaster0_p & d40d98 | !hmaster0_p & d40d55;
assign deaea6 = hgrant2_p & deaea4 | !hgrant2_p & deaea5;
assign b26784 = decide_p & b2677e | !decide_p & b26783;
assign ce9d43 = hready_p & ce9d16 | !hready_p & ce9d42;
assign b299dd = hlock0_p & cea38d | !hlock0_p & v84563c;
assign af3587 = hmaster0_p & af3582 | !hmaster0_p & af3586;
assign c3b696 = hlock0_p & c3b694 | !hlock0_p & !c3b66b;
assign a5efd7 = hbusreq2_p & a5efd1 | !hbusreq2_p & a5efd6;
assign ab051d = hbusreq2_p & ab051c | !hbusreq2_p & ab051a;
assign b266e3 = hbusreq2_p & b266e2 | !hbusreq2_p & b266e0;
assign c3bd0f = hburst1 & cea24d | !hburst1 & deada7;
assign c3bbbe = hbusreq2_p & c3bbbd | !hbusreq2_p & c3bbbc;
assign dead0d = locked_p & v84563c | !locked_p & dead0c;
assign a5f38a = hlock2_p & a5f386 | !hlock2_p & a5f389;
assign a5f247 = hlock1_p & a5fbab | !hlock1_p & !a5f246;
assign af3532 = hbusreq0_p & v84563c | !hbusreq0_p & af352c;
assign b29e48 = hgrant2_p & dead3e | !hgrant2_p & !b29c3c;
assign b29d3b = hbusreq2_p & b29d3a | !hbusreq2_p & v84563c;
assign a5f56e = stateG10_1_p & v9703fb | !stateG10_1_p & a5f56d;
assign ce9d2f = hmaster0_p & ce9d29 | !hmaster0_p & ce9d2e;
assign c3b631 = locked_p & v84563c | !locked_p & !c3b625;
assign cea448 = hlock0_p & cea389 | !hlock0_p & !cea38d;
assign b26738 = hgrant2_p & b26733 | !hgrant2_p & !b26737;
assign c3bdcb = hgrant0_p & c3bdb5 | !hgrant0_p & c3bdca;
assign b29e61 = hgrant2_p & b29e60 | !hgrant2_p & v84563c;
assign ab0712 = hlock0_p & c3bd5f | !hlock0_p & !ab06b7;
assign c3bcfb = hbusreq2_p & dead2c | !hbusreq2_p & v84563c;
assign a5efba = hlock2 & a5efb6 | !hlock2 & a5efb9;
assign a5f6e6 = hlock1_p & a5fb8b | !hlock1_p & !a5f6e5;
assign cea3cb = hlock1_p & deac52 | !hlock1_p & !cea255;
assign a5eba0 = hmaster1_p & a5eb9f | !hmaster1_p & a5ea98;
assign cea419 = hmaster1_p & cea411 | !hmaster1_p & cea418;
assign ab0749 = hmaster1_p & ab0744 | !hmaster1_p & ab0748;
assign af351a = hmaster0_p & af3518 | !hmaster0_p & af3519;
assign cea266 = hburst1 & v84563c | !hburst1 & cea265;
assign af34a3 = hbusreq2_p & af34a2 | !hbusreq2_p & af34a0;
assign ab0d07 = hlock0_p & b298a4 | !hlock0_p & !b29833;
assign deacfb = locked_p & v84563c | !locked_p & !deacdf;
assign b266ee = hgrant1_p & b266a0 | !hgrant1_p & b266ab;
assign a5fa16 = hready & a5fa11 | !hready & a5fa15;
assign d40d63 = decide_p & d40d5c | !decide_p & d40d62;
assign af3c62 = hbusreq0_p & af3c5e | !hbusreq0_p & af3c4c;
assign a5f9f4 = stateG10_1_p & v84563c | !stateG10_1_p & a60168;
assign af350c = hmaster0_p & af350b | !hmaster0_p & af348f;
assign a5ea9a = hbusreq2 & a5f0a3 | !hbusreq2 & !a5f0a5;
assign b26715 = locked_p & b2669f | !locked_p & b266a0;
assign deae91 = hlock0_p & deae90 | !hlock0_p & !v84563c;
assign cea368 = hbusreq2_p & cea367 | !hbusreq2_p & v84563c;
assign ab06ea = hbusreq2_p & ab06e9 | !hbusreq2_p & b29ab2;
assign deaeaa = hmaster0_p & deae9d | !hmaster0_p & deaea9;
assign b29a67 = hlock2_p & v84563c | !hlock2_p & !b29a66;
assign a5f234 = hlock0_p & a5f7b4 | !hlock0_p & a5f233;
assign a5f47b = hgrant2_p & a5f477 | !hgrant2_p & a5f47a;
assign a5f3f1 = hgrant1_p & a5f3f0 | !hgrant1_p & a5f3ef;
assign a5f73f = hmaster1_p & a5f735 | !hmaster1_p & a5f73e;
assign d40d32 = start_p & v84563c | !start_p & !v845674;
assign ab0550 = hbusreq3 & ab0541 | !hbusreq3 & ab054f;
assign deaceb = hbusreq1_p & deacdf | !hbusreq1_p & v84563c;
assign c3b657 = hbusreq3 & c3b656 | !hbusreq3 & !c3b653;
assign a5f8eb = hlock0_p & a5f8ea | !hlock0_p & a5f8c5;
assign deae4d = hbusreq1_p & dead76 | !hbusreq1_p & !v84563c;
assign ab0594 = hlock2_p & ab0592 | !hlock2_p & !ab0593;
assign b2672c = locked_p & b26728 | !locked_p & b2672b;
assign cea1ac = hburst0_p & v84563c | !hburst0_p & cea1ab;
assign b29d91 = hgrant2_p & b29d8f | !hgrant2_p & !b29d90;
assign c3b630 = hmaster1_p & c3b62f | !hmaster1_p & c3bbbf;
assign c3bc2f = hmaster0_p & c3bbf5 | !hmaster0_p & c3bc2e;
assign b2a01f = start_p & cea1aa | !start_p & !b2a01e;
assign b2670a = hlock0_p & b2669d | !hlock0_p & !b26695;
assign ab0bd3 = hmaster1_p & dead53 | !hmaster1_p & ab0ade;
assign b29a5a = hlock1_p & deadde | !hlock1_p & b29a59;
assign af34db = hgrant2_p & af34da | !hgrant2_p & af3c70;
assign ab0ced = hbusreq2_p & ab0cec | !hbusreq2_p & cea15a;
assign a5ef16 = hbusreq0 & a5ef0d | !hbusreq0 & !a5ef15;
assign af3539 = decide_p & af3538 | !decide_p & af3535;
assign dead07 = hbusreq3 & dead06 | !hbusreq3 & v84563c;
assign v970429 = hlock0_p & v9703fc | !hlock0_p & v84563c;
assign a5f37a = hready & a5f376 | !hready & a5f379;
assign c3bc71 = hgrant2_p & c3bc6d | !hgrant2_p & c3bc70;
assign b26724 = hgrant2_p & b2671e | !hgrant2_p & b26723;
assign a5fb75 = locked_p & v84563c | !locked_p & a5fb73;
assign b8acec = hmaster0_p & b8aceb | !hmaster0_p & b8acea;
assign c3b6a9 = hlock0_p & c3b6a6 | !hlock0_p & !c3b6a8;
assign b29fc2 = locked_p & b29fc1 | !locked_p & c3bd9a;
assign ce9d70 = hbusreq3 & ce9d6e | !hbusreq3 & ce9d6f;
assign a5f24f = hlock0_p & a5f24d | !hlock0_p & a5f24e;
assign d40d8b = decide_p & d40d79 | !decide_p & d40d8a;
assign a5fc9b = hbusreq2 & a5fc6d | !hbusreq2 & v845660;
assign bdb5b9 = hgrant3_p & bdb5b0 | !hgrant3_p & bdb5b8;
assign a5ef25 = hbusreq2 & a5edf5 | !hbusreq2 & v845660;
assign b29a76 = hgrant1_p & deada9 | !hgrant1_p & c3b691;
assign c3b63f = hbusreq0_p & c3b631 | !hbusreq0_p & c3b636;
assign af354e = hlock2_p & af354d | !hlock2_p & af354c;
assign c3b735 = hlock0_p & deae59 | !hlock0_p & c3b72f;
assign c3bc9a = hbusreq2_p & c3bc98 | !hbusreq2_p & c3bc99;
assign a5f397 = hlock0_p & a5f387 | !hlock0_p & a5f394;
assign a5f8c8 = hready & a60167 | !hready & !deaca0;
assign a5f703 = start_p & v8e1935 | !start_p & a5fb88;
assign a81ce1 = hbusreq1_p & a81ca9 | !hbusreq1_p & a81cdb;
assign ab0b70 = hbusreq2_p & ab0b6f | !hbusreq2_p & v84563c;
assign c3b6f8 = hlock1_p & deae02 | !hlock1_p & !deae4d;
assign v845644 = hlock0_p & v84563c | !hlock0_p & !v84563c;
assign c3bc88 = hbusreq2_p & c3bc87 | !hbusreq2_p & !deacfb;
assign c3bc74 = hbusreq2_p & c3bc73 | !hbusreq2_p & !deace1;
assign a81ce8 = hmaster1_p & a81ce7 | !hmaster1_p & v84563c;
assign af348b = hlock2_p & af3c49 | !hlock2_p & d40d33;
assign b299da = hbusreq2_p & b299d9 | !hbusreq2_p & v84563c;
assign b2991d = hlock2_p & v84563c | !hlock2_p & !b2991c;
assign a5ef80 = hgrant2_p & a5ef7a | !hgrant2_p & a5ef7f;
assign c3b7de = hbusreq2_p & c3b7dd | !hbusreq2_p & !c3b7dc;
assign b29a6b = hbusreq2_p & b29a67 | !hbusreq2_p & v84563c;
assign af3502 = hmaster1_p & af3c4c | !hmaster1_p & af34bf;
assign ab0bad = hbusreq2_p & ab0ba7 | !hbusreq2_p & ab0bac;
assign b2673c = hlock2_p & b2673b | !hlock2_p & b266b3;
assign a5f388 = hlock0_p & a5f387 | !hlock0_p & a5f385;
assign b29d77 = hlock1_p & deacf7 | !hlock1_p & b29d76;
assign a5ef2f = hmaster0_p & a5ef27 | !hmaster0_p & a5ef2e;
assign d40d92 = decide_p & d40d5b | !decide_p & d40d91;
assign cea24e = hburst1 & cea24d | !hburst1 & deaca0;
assign ab060a = hmaster0_p & ab0605 | !hmaster0_p & ab0609;
assign ab0534 = decide_p & ab0533 | !decide_p & v84563c;
assign b29cc9 = hlock0_p & b29cc8 | !hlock0_p & !v84563c;
assign b29fd4 = hlock2 & deaca1 | !hlock2 & b29fd3;
assign a81cff = hgrant0_p & a81cf5 | !hgrant0_p & a81cfe;
assign a5f5a2 = hready & a5f492 | !hready & c3b6bd;
assign a5785b = hgrant3_p & a57858 | !hgrant3_p & !a5785a;
assign ab0bf5 = hmaster0_p & ab0bef | !hmaster0_p & ab0bf4;
assign b29fe4 = hbusreq3 & b29fe3 | !hbusreq3 & b29fe1;
assign af3c71 = hmaster1_p & af3c70 | !hmaster1_p & af3c64;
assign a5f593 = hlock2_p & a5f4f1 | !hlock2_p & a5f592;
assign dead2f = hbusreq3 & dead2e | !hbusreq3 & dead2d;
assign adaeca = hlock1_p & adaec4 | !hlock1_p & v84563c;
assign ab0cd8 = hbusreq3 & ab0cd7 | !hbusreq3 & v84564a;
assign b2670e = hlock0_p & b2669d | !hlock0_p & !b266a2;
assign a5fcfb = hbusreq1 & a5fcf8 | !hbusreq1 & !a5fcfa;
assign cea2a2 = hlock2_p & cea2a1 | !hlock2_p & v84563c;
assign b29fbf = hgrant2_p & dead3e | !hgrant2_p & !b29fbe;
assign b298b0 = hlock2_p & v84563c | !hlock2_p & !b298af;
assign a5f559 = hbusreq1 & a5f556 | !hbusreq1 & a5f558;
assign b2996b = hlock2_p & b2996a | !hlock2_p & !b29943;
assign b298a9 = hmaster0_p & b29838 | !hmaster0_p & b298a8;
assign ab06da = hready_p & ab0689 | !hready_p & ab06d9;
assign a5f72e = hbusreq2_p & a5f72d | !hbusreq2_p & a60142;
assign deac7d = hbusreq3 & deac7c | !hbusreq3 & v84563c;
assign a5f38e = hbusreq1 & a5f38d | !hbusreq1 & !v84563c;
assign cea3f0 = hbusreq2_p & cea3ec | !hbusreq2_p & cea3eb;
assign c3bda5 = hgrant0_p & c3bd93 | !hgrant0_p & c3bda4;
assign adaef1 = hlock1_p & adaebc | !hlock1_p & adaef0;
assign a5edf4 = hmaster1_p & a5edf3 | !hmaster1_p & v84563c;
assign a5fbf5 = hbusreq2_p & a5fbf4 | !hbusreq2_p & a5fbea;
assign a5f71a = hbusreq2_p & a5f719 | !hbusreq2_p & !v84563c;
assign b2669d = locked_p & v84563c | !locked_p & b26697;
assign c3bcb4 = hbusreq3 & v84563c | !hbusreq3 & !c3bcb3;
assign b29971 = hlock2_p & b29970 | !hlock2_p & !b29943;
assign ab0732 = hbusreq3 & b29ab2 | !hbusreq3 & dead2e;
assign a5f6f8 = hready & a5f9dd | !hready & !dead33;
assign af349b = hready_p & af3c73 | !hready_p & af349a;
assign ab0562 = hlock2_p & ab0560 | !hlock2_p & ab0561;
assign c3bc4b = hbusreq2_p & c3bc4a | !hbusreq2_p & c3bc49;
assign c3bdae = hlock1_p & deae02 | !hlock1_p & c3bdad;
assign b266b3 = hlock0_p & b266a8 | !hlock0_p & b266b1;
assign c3b644 = hbusreq3 & c3b643 | !hbusreq3 & c3b63d;
assign a5f22e = hlock0_p & a5f22d | !hlock0_p & a5f92e;
assign ce9d14 = hmaster0_p & ce9cf8 | !hmaster0_p & ce9d13;
assign c3b6f1 = hgrant2_p & c3b6f0 | !hgrant2_p & c3bc70;
assign cea15e = hbusreq2_p & cea149 | !hbusreq2_p & v84563c;
assign b29c3b = hlock2_p & v84563c | !hlock2_p & dead39;
assign b29cc1 = hgrant2_p & b29cbe | !hgrant2_p & b29cc0;
assign b29944 = hlock2_p & b2993f | !hlock2_p & b29943;
assign dea761 = hbusreq2_p & deadfe | !hbusreq2_p & v84563c;
assign af34e1 = hgrant0_p & af34d1 | !hgrant0_p & af34e0;
assign b266a5 = hlock2_p & b266a4 | !hlock2_p & b266a3;
assign cea16a = hlock0_p & dead24 | !hlock0_p & v845660;
assign cea375 = hlock1_p & deacf7 | !hlock1_p & !cea374;
assign a5eb82 = hmaster1_p & a5ea1a | !hmaster1_p & a5fd37;
assign b2982a = stateA1_p & c07311 | !stateA1_p & !v84563c;
assign a5f53d = hready & v84563c | !hready & a5f53c;
assign ab0ba3 = locked_p & v84563c | !locked_p & !b29d82;
assign c3b650 = hbusreq2_p & c3b625 | !hbusreq2_p & !c3b635;
assign a5f219 = hmaster0_p & a5f216 | !hmaster0_p & a5f218;
assign a5fae7 = hbusreq2_p & a5fad7 | !hbusreq2_p & a5fad1;
assign c3bc46 = hready_p & c3bbc1 | !hready_p & c3bc45;
assign ab05ad = hbusreq2_p & ab05a9 | !hbusreq2_p & ab05ac;
assign c3b6d9 = hbusreq2_p & c3b6d8 | !hbusreq2_p & c3b6d6;
assign dead5e = hgrant2_p & v84564a | !hgrant2_p & dead53;
assign a5f20e = hbusreq2_p & a5f20d | !hbusreq2_p & !v84563c;
assign d40d6d = hbusreq1_p & d40d2b | !hbusreq1_p & d40d67;
assign a5eadb = hlock0_p & a5f7b4 | !hlock0_p & a5eada;
assign a5f26b = hbusreq2 & a5fcdb | !hbusreq2 & v84563c;
assign c3b7d4 = hbusreq2_p & c3b7c2 | !hbusreq2_p & c3b7bd;
assign b29d04 = hbusreq2_p & b29d03 | !hbusreq2_p & !v84563c;
assign ab06f4 = hlock2_p & ab06f3 | !hlock2_p & ab06e1;
assign c3b6ef = hlock2_p & c3b640 | !hlock2_p & !c3b656;
assign deacd8 = hmaster1_p & deacc4 | !hmaster1_p & deacd7;
assign adaf18 = hready_p & adaf14 | !hready_p & adaf17;
assign c3bc2a = hbusreq2_p & c3bc17 | !hbusreq2_p & c3bc15;
assign a5f29b = hbusreq2_p & a5f29a | !hbusreq2_p & !v84563c;
assign c3b80d = hgrant2_p & c3b808 | !hgrant2_p & c3b80c;
assign c3bd07 = hmaster0_p & c3bd00 | !hmaster0_p & c3bd06;
assign af3c15 = hmaster1_p & af3c14 | !hmaster1_p & !v84563c;
assign ce9e09 = hmaster1_p & ce9df0 | !hmaster1_p & ce9dfe;
assign af3c47 = hbusreq3_p & af3c40 | !hbusreq3_p & af3c46;
assign ab0bba = hbusreq2_p & cea15a | !hbusreq2_p & v845644;
assign a5fb21 = hbusreq2 & a5fb14 | !hbusreq2 & a5fb20;
assign c3b750 = hmaster0_p & c3b74f | !hmaster0_p & c3b6e6;
assign b29d6c = start_p & v84563c | !start_p & !v84566c;
assign a5fbd9 = hlock1_p & a5fb8b | !hlock1_p & v84563c;
assign a5fc15 = hbusreq2 & a5fc07 | !hbusreq2 & !a5fc14;
assign ab0b33 = hmaster1_p & ab0b11 | !hmaster1_p & !ab0b32;
assign c3bc84 = hmaster1_p & c3bc71 | !hmaster1_p & c3bc83;
assign b29d20 = hbusreq2_p & b29d0e | !hbusreq2_p & v84563c;
assign ce9dda = hmaster1_p & ce9dc6 | !hmaster1_p & ce9dd4;
assign a5f51c = hlock0_p & a5f516 | !hlock0_p & a5f51b;
assign a81d0d = hbusreq3_p & a81d02 | !hbusreq3_p & a81d0c;
assign a5fba6 = hmastlock_p & a5fba5 | !hmastlock_p & !v84563c;
assign a5efc0 = hlock2 & a5f3ba | !hlock2 & a5efbf;
assign deadf7 = hready_p & deada0 | !hready_p & deadf6;
assign ab0b00 = hlock0_p & ab0afa | !hlock0_p & c3bd60;
assign a5ea78 = hbusreq0 & a5ea77 | !hbusreq0 & a5f084;
assign dead1b = hbusreq2_p & deace9 | !hbusreq2_p & dead1a;
assign b29b0c = hlock2_p & v84563c | !hlock2_p & !b29ab2;
assign c3b624 = hlock1_p & b26695 | !hlock1_p & v84563c;
assign a5ebeb = decide_p & a5ebcc | !decide_p & a5ebea;
assign c3b77d = hready_p & c3b77c | !hready_p & c3b776;
assign b29f7f = hbusreq2_p & b29f7d | !hbusreq2_p & v84563c;
assign a5edbf = hlock0_p & a5edbe | !hlock0_p & a5f51b;
assign c3b6e6 = hmaster1_p & c3b6dc | !hmaster1_p & c3b6e5;
assign deacd4 = hbusreq3 & deacc5 | !hbusreq3 & !deacd3;
assign a5f6e4 = hlock1_p & a5f9dd | !hlock1_p & a5fb8a;
assign a5eb34 = hbusreq0 & a5ea27 | !hbusreq0 & v84563c;
assign a5fb80 = hbusreq1_p & a5fb71 | !hbusreq1_p & v84563c;
assign b29aef = hmaster0_p & b29aea | !hmaster0_p & !b29a8a;
assign ab05ce = hgrant2_p & ab05cd | !hgrant2_p & cea15a;
assign ab0cc3 = hready & v84563c | !hready & !deadb9;
assign c3bddb = hbusreq2_p & c3bdd2 | !hbusreq2_p & deac1e;
assign a5ebcc = hmaster0_p & a5ebca | !hmaster0_p & a5ebcb;
assign ab0b0b = hlock0_p & v84563c | !hlock0_p & !ab0b0a;
assign b29ff7 = hgrant2_p & b29ff6 | !hgrant2_p & b29f7f;
assign b29eb9 = hlock1_p & v84563c | !hlock1_p & !b29eb8;
assign a5eecc = hmaster1_p & a5eecb | !hmaster1_p & v84563c;
assign c3b797 = hlock0_p & c3bcda | !hlock0_p & !dead77;
assign a5fcd3 = stateA1_p & c07311 | !stateA1_p & deacf2;
assign c3b70e = hmaster0_p & c3b704 | !hmaster0_p & c3b70d;
assign c3bc8f = hgrant2_p & c3bc89 | !hgrant2_p & c3bc8e;
assign a5ea42 = hlock0_p & a5f9a3 | !hlock0_p & a5ea40;
assign b29aba = hready & deae02 | !hready & !v84563c;
assign adaef6 = hgrant2_p & adaef5 | !hgrant2_p & v84563c;
assign a5fc7a = locked_p & a5fc79 | !locked_p & c3bcdb;
assign c3b7eb = hbusreq2_p & c3b7e9 | !hbusreq2_p & c3b7ea;
assign a5fa27 = hlock2_p & a5fa23 | !hlock2_p & a5fa26;
assign cea335 = hlock0_p & cea334 | !hlock0_p & v84563c;
assign b29ebe = locked_p & b29ebd | !locked_p & !v84563c;
assign c98ba0 = hgrant2_p & v8c6711 | !hgrant2_p & v84563c;
assign a81cea = hgrant0_p & a81ce0 | !hgrant0_p & a81ce9;
assign a5fcc3 = hgrant0_p & a5fc97 | !hgrant0_p & a5fcc2;
assign cea883 = hlock1_p & v84563c | !hlock1_p & deac56;
assign a5f1e6 = hlock0_p & a5f1e5 | !hlock0_p & a5fad4;
assign cea44f = hbusreq2_p & cea44e | !hbusreq2_p & cea44c;
assign cea18c = hready_p & v84563c | !hready_p & cea18b;
assign af3c28 = hlock3_p & af3c24 | !hlock3_p & af3c27;
assign a5ef45 = hbusreq3 & a5eebc | !hbusreq3 & a5eec4;
assign ab057e = hlock0_p & ab057d | !hlock0_p & !ab0570;
assign v856b00 = stateG3_1_p & v84563c | !stateG3_1_p & v85f3c3;
assign a5fbaf = hbusreq1_p & a5fbae | !hbusreq1_p & a5fbab;
assign a5fbe2 = hlock1_p & a5fbe1 | !hlock1_p & v84563c;
assign a5f9dc = start_p & v84563c | !start_p & a5f9db;
assign b29ce4 = hready & deadac | !hready & c3bd16;
assign a5f8e0 = hmastlock_p & a5f8df | !hmastlock_p & !v84563c;
assign ab0b84 = hlock0_p & v84563c | !hlock0_p & !b29d6f;
assign a5f212 = hgrant2_p & v84563c | !hgrant2_p & a5f209;
assign b29e6a = hbusreq2_p & b29e69 | !hbusreq2_p & v845644;
assign b26753 = hgrant0_p & b26746 | !hgrant0_p & b26752;
assign b29d66 = hready & deace1 | !hready & !v84563c;
assign b29ed2 = hmaster0_p & b29ecb | !hmaster0_p & b29ed1;
assign c3bbfb = hlock1_p & c3bbd2 | !hlock1_p & c3bbfa;
assign v970453 = hready_p & v97044e | !hready_p & v970452;
assign af3570 = hmaster1_p & af352d | !hmaster1_p & af356f;
assign ab0b8d = hlock0_p & v84563c | !hlock0_p & !b29d83;
assign a5f704 = hmastlock_p & a5f703 | !hmastlock_p & v84563c;
assign ce9cbb = hmaster1_p & ce9cba | !hmaster1_p & cea191;
assign deac3e = hbusreq3 & deac34 | !hbusreq3 & v84563c;
assign ce9d37 = hmaster1_p & ce9d33 | !hmaster1_p & ce9d36;
assign b29982 = hmaster1_p & b29981 | !hmaster1_p & b29d64;
assign a5ede4 = hmaster0_p & a5f59a | !hmaster0_p & a5ede3;
assign a5f137 = hbusreq2_p & a5f0db | !hbusreq2_p & a5f0d1;
assign a5e9bd = hlock0_p & a5e9bb | !hlock0_p & a5e9bc;
assign dea6bc = hbusreq2_p & dea6bb | !hbusreq2_p & dea6ba;
assign b29efb = hlock0_p & b29ef5 | !hlock0_p & b29efa;
assign a5f14b = hlock0_p & a5f14a | !hlock0_p & a5f144;
assign a5f1a9 = hlock2_p & a5f1a6 | !hlock2_p & a5f1a8;
assign dead09 = stateG10_1_p & b26693 | !stateG10_1_p & deace0;
assign c3b675 = hburst1 & v84563c | !hburst1 & c3b674;
assign a5eaea = hlock2_p & a5eae5 | !hlock2_p & !a5eae9;
assign c3bd96 = hbusreq2_p & c3bd95 | !hbusreq2_p & c3bc6e;
assign a5f3b0 = hlock0_p & a5f36e | !hlock0_p & a5f36b;
assign b2674c = hlock2_p & b26699 | !hlock2_p & b266b8;
assign ab0cf1 = hmaster1_p & ab0cee | !hmaster1_p & ab0cf0;
assign a5fa1c = hmastlock_p & v9703fb | !hmastlock_p & !v84563c;
assign c3b802 = hready_p & c3b7b7 | !hready_p & c3b801;
assign a5f4b9 = hlock0_p & a5f4a8 | !hlock0_p & a5f4b8;
assign b2a018 = hmaster0_p & b2a014 | !hmaster0_p & b2a017;
assign a5f1a6 = hbusreq2 & a5f1a5 | !hbusreq2 & a5f1a4;
assign cea248 = hburst0 & cea246 | !hburst0 & cea247;
assign a5f03b = hmaster0_p & v84563c | !hmaster0_p & a5f03a;
assign ab0c8e = hlock2_p & ab0c8d | !hlock2_p & !c3bca0;
assign a5f7f7 = hbusreq1_p & a5f7f5 | !hbusreq1_p & !a5fbab;
assign cea2ef = hbusreq2_p & cea16b | !hbusreq2_p & cea15a;
assign cea2ea = hlock0_p & cea2e9 | !hlock0_p & v84563c;
assign a5fb60 = hbusreq2_p & a5fb5f | !hbusreq2_p & a5fad6;
assign v845666 = hgrant2_p & v84563c | !hgrant2_p & !v84563c;
assign af34ab = hmaster0_p & af34a4 | !hmaster0_p & af34aa;
assign a5fc6e = hbusreq3 & a5fc6d | !hbusreq3 & v84563c;
assign deacf1 = hburst1_p & c07311 | !hburst1_p & !v84563c;
assign a5f583 = hlock2_p & a5f577 | !hlock2_p & !a5f582;
assign ab071b = hbusreq2_p & ab0717 | !hbusreq2_p & ab0715;
assign a5ee7d = hmaster0_p & a5ee42 | !hmaster0_p & a5ee7c;
assign b26780 = hmaster0_p & b2677f | !hmaster0_p & b2675a;
assign ab0b7e = hlock2 & ab0b7c | !hlock2 & ab0b7d;
assign b29e57 = hgrant0_p & v84563c | !hgrant0_p & !v845666;
assign a5ef74 = hbusreq3 & a5ef72 | !hbusreq3 & a5ef73;
assign a5f083 = hlock2_p & a5fbc1 | !hlock2_p & v84563c;
assign a5fad1 = hlock0_p & a5fa37 | !hlock0_p & v84563c;
assign af356b = hgrant2_p & af355e | !hgrant2_p & af356a;
assign a5fd01 = hbusreq3 & a5fd00 | !hbusreq3 & v84563c;
assign c3b7e9 = hlock2_p & c3b7e8 | !hlock2_p & !c3b7e4;
assign a5f9c9 = hbusreq3 & a5f9c7 | !hbusreq3 & a5f9c8;
assign c3bce1 = hlock0_p & cea1bf | !hlock0_p & !c3bce0;
assign a5fce0 = start_p & a5fc8a | !start_p & c07311;
assign b29fe7 = hmaster0_p & b29fe6 | !hmaster0_p & !b29f5e;
assign ab0c5e = hlock0_p & ab0c5c | !hlock0_p & ab0c5d;
assign c3bdea = decide_p & c3bde9 | !decide_p & !v845660;
assign a5f28a = hgrant0_p & a5f271 | !hgrant0_p & a5f289;
assign ab054d = hlock0_p & v84563c | !hlock0_p & !b2992b;
assign a5ee18 = hbusreq2 & a5ee16 | !hbusreq2 & a5ee17;
assign ab05a5 = hlock0_p & b298a4 | !hlock0_p & !ab05a4;
assign a5f109 = hlock0_p & a5f7fd | !hlock0_p & !a5f108;
assign ab0c49 = hgrant2_p & ab0c47 | !hgrant2_p & ab0c48;
assign b29fb4 = hready & b29fb3 | !hready & v84563c;
assign cea412 = hbusreq0_p & cea3fb | !hbusreq0_p & cea405;
assign cea44d = hlock0_p & cea37c | !hlock0_p & cea44b;
assign ab0c40 = hlock2_p & ab0c3c | !hlock2_p & ab0c3f;
assign a5f510 = hbusreq2 & a5f500 | !hbusreq2 & a5f4f1;
assign a5ef96 = hlock0_p & a5f390 | !hlock0_p & a5f38f;
assign ab06c2 = hbusreq2_p & ab06c0 | !hbusreq2_p & !ab06c1;
assign ab0c2b = hmaster0_p & ab0c24 | !hmaster0_p & ab0c2a;
assign v877992 = hmaster1_p & v845646 | !hmaster1_p & !v84563c;
assign deae02 = hmastlock_p & deae01 | !hmastlock_p & v84563c;
assign cea26c = stateG10_1_p & cea268 | !stateG10_1_p & cea26b;
assign ce9d29 = hmaster1_p & ce9d22 | !hmaster1_p & !ce9d28;
assign ab0656 = jx1_p & ab063e | !jx1_p & ab0655;
assign b266fe = hbusreq2_p & b266fc | !hbusreq2_p & b266fa;
assign a5f095 = hlock2_p & v845641 | !hlock2_p & v84563c;
assign a5fbed = start_p & v845654 | !start_p & !a5fbac;
assign b8acdb = hgrant1_p & b8acda | !hgrant1_p & v845646;
assign a5f4c8 = stateG10_1_p & v970407 | !stateG10_1_p & a5f4c7;
assign af35b6 = hbusreq2_p & af35b4 | !hbusreq2_p & af3563;
assign a5f0dc = hbusreq2_p & a5f0db | !hbusreq2_p & a5f0da;
assign b29d38 = hbusreq3 & b29d30 | !hbusreq3 & !b29d37;
assign c3bcd6 = hready_p & c3bcc4 | !hready_p & c3bcd5;
assign af3485 = hbusreq2_p & af3c81 | !hbusreq2_p & af3c7f;
assign b2982f = hbusreq1_p & v84563c | !hbusreq1_p & !dead7b;
assign a5fb13 = hready & a5fb12 | !hready & v84563c;
assign deacdc = hready_p & deac11 | !hready_p & deacdb;
assign ab0b40 = hgrant2_p & ab0b3d | !hgrant2_p & ab0b3f;
assign cea33b = hmaster1_p & cea33a | !hmaster1_p & !cea289;
assign cea461 = hbusreq2_p & cea444 | !hbusreq2_p & cea460;
assign b29eaa = hlock0_p & dead34 | !hlock0_p & !b29ea9;
assign b29cfc = hbusreq3 & b29cec | !hbusreq3 & b29cfb;
assign a5edc1 = hlock0_p & a5edc0 | !hlock0_p & a5f525;
assign ab0b0f = hbusreq2_p & ab0b02 | !hbusreq2_p & ab0b0e;
assign a5f439 = hbusreq1_p & a5fa1d | !hbusreq1_p & v84565a;
assign c3bcea = hlock2_p & v84563c | !hlock2_p & v845660;
assign af359c = hgrant2_p & af352d | !hgrant2_p & af3572;
assign cea35e = hgrant2_p & cea159 | !hgrant2_p & !cea35d;
assign deacaa = hlock1_p & v84565a | !hlock1_p & !v84563c;
assign a5fc0e = hbusreq1_p & a5fc0d | !hbusreq1_p & a5fbab;
assign b29997 = hgrant2_p & b29996 | !hgrant2_p & !b29c3c;
assign a5f708 = hlock1_p & a5fbab | !hlock1_p & !a5f707;
assign dea739 = decide_p & dea738 | !decide_p & v84563c;
assign a5f948 = hbusreq2 & a5f945 | !hbusreq2 & a5f947;
assign a5fbc4 = hbusreq2_p & a5fbc3 | !hbusreq2_p & v84563c;
assign deacb2 = hmaster1_p & v84563c | !hmaster1_p & deacb1;
assign deadc9 = hbusreq2_p & deadb4 | !hbusreq2_p & deac1e;
assign a5f421 = hlock2_p & a5f40e | !hlock2_p & a5f420;
assign b29f1b = hgrant1_p & b29f1a | !hgrant1_p & b29f19;
assign dea732 = hmaster1_p & dea72f | !hmaster1_p & dea731;
assign a5ee1c = hlock1_p & a5fba2 | !hlock1_p & !a5ee1b;
assign ab0bc2 = hmaster1_p & ab0bbd | !hmaster1_p & ab0bbe;
assign cea268 = hmastlock_p & cea267 | !hmastlock_p & v84563c;
assign b266c0 = hmaster1_p & b26699 | !hmaster1_p & !b266a3;
assign a5f83c = hready & a5f836 | !hready & a5f83b;
assign b26748 = hgrant2_p & b26747 | !hgrant2_p & b266a8;
assign a5f4e6 = stateG10_1_p & v970407 | !stateG10_1_p & a5f4e5;
assign a5fd17 = hmaster1_p & a5fd0b | !hmaster1_p & a5fd16;
assign c3bbef = hbusreq2_p & c3bbea | !hbusreq2_p & deacaa;
assign cea17d = hmaster1_p & cea178 | !hmaster1_p & cea17c;
assign a5ebe9 = hmaster0_p & a5ebe8 | !hmaster0_p & a5eb44;
assign a5ea20 = hbusreq0 & a5ea1f | !hbusreq0 & v84563c;
assign b2a014 = hmaster1_p & b2a013 | !hmaster1_p & !b29f46;
assign a5f938 = hlock1_p & deac52 | !hlock1_p & a5f937;
assign a5f7f8 = hgrant1_p & a5f7f6 | !hgrant1_p & a5f7f7;
assign b29ee1 = decide_p & b29ee0 | !decide_p & v84563c;
assign a5eb89 = decide_p & a5eb83 | !decide_p & !a5eb88;
assign a5fc87 = hmastlock_p & a5fc86 | !hmastlock_p & !v84563c;
assign cea426 = hbusreq3 & cea424 | !hbusreq3 & cea425;
assign a5f29f = decide_p & a5f297 | !decide_p & !a5f29e;
assign v97042c = hmaster1_p & v84563c | !hmaster1_p & v970413;
assign c3b73d = hmaster0_p & c3b734 | !hmaster0_p & c3b73c;
assign v97043b = hmaster0_p & v970436 | !hmaster0_p & v97043a;
assign a5eb88 = hmaster0_p & a5eb87 | !hmaster0_p & !a5ea2d;
assign a5f16f = hready & a5f9e0 | !hready & !c3bbf9;
assign b29ac6 = hlock3_p & b29ab9 | !hlock3_p & b29ac5;
assign a5fc28 = hbusreq0_p & a5fbc0 | !hbusreq0_p & a5fc1c;
assign b29d2a = hbusreq3 & v84563c | !hbusreq3 & b29cd8;
assign c3bc8a = locked_p & v84563c | !locked_p & dead18;
assign a5fcb5 = hbusreq3 & a5fcb4 | !hbusreq3 & v84563c;
assign cea178 = hgrant2_p & v84563c | !hgrant2_p & !v845660;
assign c3bd3e = hready & c3bd3b | !hready & c3bd3d;
assign a9b9d0 = locked_p & v84565a | !locked_p & !v84563c;
assign cea421 = hlock2_p & cea420 | !hlock2_p & cea405;
assign d40d7c = hbusreq0_p & d40d31 | !hbusreq0_p & d40d7b;
assign cea428 = hmaster1_p & cea427 | !hmaster1_p & !deacaa;
assign c3b757 = decide_p & c3b756 | !decide_p & v845660;
assign a5f1b9 = hmaster1_p & a5f99e | !hmaster1_p & a5f1b8;
assign c3bdd6 = hready & c3bd37 | !hready & deadb9;
assign a5eb8d = hlock0_p & a5eb8c | !hlock0_p & v84563c;
assign cea45c = hmaster1_p & cea458 | !hmaster1_p & cea45b;
assign deade4 = hgrant2_p & deade2 | !hgrant2_p & deade3;
assign b299ee = hmaster1_p & b29f4f | !hmaster1_p & !b299ed;
assign a5f074 = hbusreq2_p & a5f073 | !hbusreq2_p & a5f071;
assign af35a1 = hready_p & af3591 | !hready_p & af35a0;
assign a5f558 = hlock1_p & v84563c | !hlock1_p & a5f557;
assign a5fc57 = hbusreq3 & a5fc56 | !hbusreq3 & v84563c;
assign ab06fb = hlock2_p & ab06fa | !hlock2_p & ab067f;
assign a5f306 = decide_p & a5f2fd | !decide_p & a5f305;
assign ab05d3 = hmaster1_p & ab05ce | !hmaster1_p & ab05d2;
assign d40d8a = hgrant0_p & d40d7f | !hgrant0_p & d40d89;
assign c3b828 = hbusreq2_p & c3b827 | !hbusreq2_p & !c3b812;
assign cea8a8 = stateG10_1_p & cea8a7 | !stateG10_1_p & deadde;
assign v84563c = 1;
assign c3b64b = hlock2_p & c3b64a | !hlock2_p & c3b649;
assign c3bd60 = hready & v84565a | !hready & v84563c;
assign b29d3a = hlock2_p & b29d39 | !hlock2_p & v84563c;
assign hmastlock = bdb5ba;
assign ce9db0 = hgrant3_p & ce9d43 | !hgrant3_p & ce9daf;
assign a5f575 = hready & a5f56c | !hready & a5f574;
assign a5ea69 = hlock0_p & a5f2f2 | !hlock0_p & v84563c;
assign c3bcdc = locked_p & dead6e | !locked_p & c3bcdb;
assign a5f023 = hmaster0_p & a5f01b | !hmaster0_p & a5f022;
assign c3bca4 = hgrant2_p & dead3e | !hgrant2_p & v845660;
assign cea0d6 = hmaster1_p & cea0c2 | !hmaster1_p & cea0d5;
assign b29f33 = hlock2 & b29f1f | !hlock2 & b29f32;
assign deac64 = hmaster1_p & deac3f | !hmaster1_p & !deac63;
assign ce9cc3 = hlock2_p & cea40f | !hlock2_p & !cea405;
assign c3bcf0 = locked_p & v84563c | !locked_p & c3bcef;
assign a5fcc1 = hmaster1_p & a5fcb6 | !hmaster1_p & a5fcc0;
assign b29838 = hmaster1_p & b29837 | !hmaster1_p & b29c3d;
assign b29d90 = hbusreq3 & b29d5a | !hbusreq3 & b29c3c;
assign b29ee0 = hlock3_p & b29ed2 | !hlock3_p & b29edf;
assign deadd7 = hlock2_p & deadd6 | !hlock2_p & !v84563c;
assign a5f09e = hbusreq0 & a5f09d | !hbusreq0 & v845641;
assign a5f7bb = hlock0_p & a5f7b4 | !hlock0_p & a5f7ba;
assign ab0ce1 = hbusreq2_p & ab0c7a | !hbusreq2_p & !b29cbb;
assign c3bd17 = hready & c3bd15 | !hready & c3bd16;
assign cea291 = hgrant1_p & cea250 | !hgrant1_p & cea252;
assign a5f8d8 = stateA1_p & v845654 | !stateA1_p & !a81ca6;
assign ab073e = decide_p & ab073d | !decide_p & v84563c;
assign b29834 = hlock0_p & b29833 | !hlock0_p & !v84563c;
assign a5fb7b = hlock0_p & a5fb7a | !hlock0_p & v84563c;
assign d40d3a = hmastlock_p & v845674 | !hmastlock_p & !v84563c;
assign deacc2 = hbusreq2_p & deacbf | !hbusreq2_p & !v84563c;
assign a9b9dd = hbusreq2_p & a9b9dc | !hbusreq2_p & v845660;
assign b29cbc = hlock2_p & v84563c | !hlock2_p & b29cbb;
assign ab06a9 = hbusreq1_p & b29ee9 | !hbusreq1_p & v84565a;
assign ab0bb6 = hgrant0_p & ab0b6e | !hgrant0_p & !ab0bb5;
assign b2997b = hmaster0_p & b29979 | !hmaster0_p & b2997a;
assign a5fc3d = hlock0_p & v84563c | !hlock0_p & a5fb92;
assign cea445 = hlock2_p & cea443 | !hlock2_p & cea444;
assign ce9daf = hready_p & ce9d5b | !hready_p & ce9da6;
assign a5eec4 = locked_p & a5eec3 | !locked_p & v84563c;
assign b29f62 = hlock2_p & c3bd60 | !hlock2_p & !v84563c;
assign a5fc8b = start_p & a5fc8a | !start_p & d615cf;
assign b26768 = hready_p & b26766 | !hready_p & !b26767;
assign cea2f5 = hgrant2_p & cea159 | !hgrant2_p & !cea2f4;
assign a5f74b = hbusreq2 & a5fc7a | !hbusreq2 & v84563c;
assign a5f97d = hburst0_p & v845672 | !hburst0_p & a5f97c;
assign b2672d = hlock0_p & b2672a | !hlock0_p & b2672c;
assign a60166 = stateA1_p & v84563c | !stateA1_p & !a60165;
assign a5fcf3 = hlock1_p & a5fb8b | !hlock1_p & a5fcf2;
assign c3b821 = hbusreq2_p & c3b820 | !hbusreq2_p & c3b81f;
assign ce9db5 = hbusreq2_p & cea343 | !hbusreq2_p & cea342;
assign ab0677 = hbusreq3 & ab0676 | !hbusreq3 & v845660;
assign deacea = hlock0_p & deace9 | !hlock0_p & b26695;
assign a5f3d6 = hbusreq1 & a5f3d5 | !hbusreq1 & !v84563c;
assign ab0624 = hgrant0_p & ab060a | !hgrant0_p & !ab0623;
assign b26757 = locked_p & b26756 | !locked_p & b266a0;
assign b29d7b = locked_p & b29d7a | !locked_p & v84563c;
assign b29a95 = hmaster1_p & b29a94 | !hmaster1_p & b29a6e;
assign a5ef59 = hbusreq2 & a5f4fc | !hbusreq2 & a5ef58;
assign a5f756 = hmaster0_p & a5f752 | !hmaster0_p & a5f755;
assign a5fca3 = hlock1_p & v84563c | !hlock1_p & a5fca2;
assign dea72d = hbusreq2_p & dead8d | !hbusreq2_p & dead8c;
assign af35ad = hmaster0_p & af35ac | !hmaster0_p & af3586;
assign c3b705 = locked_p & c3b6f8 | !locked_p & !c3b625;
assign ab0c46 = hlock2_p & ab0ad6 | !hlock2_p & ab0c45;
assign cea413 = hlock0_p & cea40b | !hlock0_p & cea412;
assign a5f3db = hlock0_p & a5f3d2 | !hlock0_p & a5f3da;
assign c3bd47 = hready & c3bbd1 | !hready & v845648;
assign cea478 = stateG10_1_p & deaca1 | !stateG10_1_p & cea3b8;
assign a5eed2 = hgrant2_p & a5eed1 | !hgrant2_p & v84563c;
assign c3b800 = hlock3_p & c3b7ee | !hlock3_p & !c3b7ff;
assign a9b9ec = hgrant3_p & a9b9d5 | !hgrant3_p & !a9b9eb;
assign c3bc5f = hbusreq3 & c3bc5b | !hbusreq3 & c3bc5e;
assign v970445 = hlock1_p & v9703fc | !hlock1_p & v970444;
assign a5fc68 = start_p & v84563c | !start_p & v84566c;
assign ab0c6b = hlock2_p & ab0c6a | !hlock2_p & v84563c;
assign a5f720 = hbusreq2 & a5f71f | !hbusreq2 & a5fb7b;
assign a5f888 = hmaster1_p & a5f858 | !hmaster1_p & a5f887;
assign ce9e60 = jx2_p & cea373 | !jx2_p & ce9e5f;
assign b29ce0 = hlock0_p & b29cdd | !hlock0_p & !b29cdf;
assign dead48 = hbusreq3 & v845660 | !hbusreq3 & dead3b;
assign ab0add = hlock0_p & ab0adc | !hlock0_p & deacaa;
assign adaebe = hmaster1_p & adaebd | !hmaster1_p & v84563c;
assign ab0cb0 = hlock2_p & ab0caf | !hlock2_p & !c3bca0;
assign deae31 = locked_p & v84563c | !locked_p & !deae30;
assign a5efae = hready & a5ee25 | !hready & !v845648;
assign stateG10_2 = !be34ea;
assign a5eb95 = hlock2_p & a5ea69 | !hlock2_p & a5eb94;
assign ab0526 = hbusreq3 & ab0521 | !hbusreq3 & ab0525;
assign ce9cb8 = hlock2_p & cea38f | !hlock2_p & !cea38d;
assign a5f362 = hbusreq3_p & a5f28d | !hbusreq3_p & a5f361;
assign b29a1c = hlock3_p & b299ff | !hlock3_p & b29a1b;
assign a5e9d6 = hbusreq2_p & a5e9d5 | !hbusreq2_p & a5f199;
assign a5ea87 = hbusreq0 & a5ea86 | !hbusreq0 & a5ea67;
assign a5ea43 = hready & a5fbdd | !hready & !v84563c;
assign ab062a = hbusreq3 & ab0627 | !hbusreq3 & ab0629;
assign a5f21b = decide_p & a5f207 | !decide_p & a5f21a;
assign cea471 = hbusreq2_p & cea470 | !hbusreq2_p & cea3aa;
assign a5f735 = hbusreq3 & a5f734 | !hbusreq3 & v84563c;
assign deac88 = hlock0_p & deac52 | !hlock0_p & deac86;
assign a5f8ea = hready & v84563c | !hready & a5f8e9;
assign deae22 = hlock1_p & v84565a | !hlock1_p & !deae21;
assign a5f715 = hready & a5f710 | !hready & !a5f714;
assign a5fb87 = hburst0_p & d5edb8 | !hburst0_p & a5fb86;
assign a5ee65 = hready & a5ee25 | !hready & !deae59;
assign c3bc94 = hlock0_p & c3bc48 | !hlock0_p & v845660;
assign a5ea13 = hlock0_p & a5fa5e | !hlock0_p & a5e9bc;
assign a5ec22 = hready_p & a60147 | !hready_p & a5ec21;
assign a81cdd = hbusreq0_p & a81caa | !hbusreq0_p & a81cdc;
assign cea1a7 = hready_p & cea195 | !hready_p & !cea1a6;
assign a6016a = stateA1_p & a81ca6 | !stateA1_p & !v8e1935;
assign c0730a = stateG3_1_p & v84563c | !stateG3_1_p & v845674;
assign a5fbb9 = hlock0_p & a5fbb8 | !hlock0_p & a5fbb3;
assign a5f966 = hlock2_p & a5f965 | !hlock2_p & v84563c;
assign ab0ae4 = hgrant2_p & ab0ae1 | !hgrant2_p & ab0ae3;
assign a5ef52 = hready & v84563c | !hready & a5ef51;
assign a5f187 = hbusreq1_p & a60187 | !hbusreq1_p & !a5fbab;
assign cea397 = hbusreq2_p & cea396 | !hbusreq2_p & cea394;
assign c3bcf8 = locked_p & v84563c | !locked_p & c3bcdb;
assign c3bbba = hready & deae59 | !hready & v845648;
assign bdb58a = hmaster1_p & v84565a | !hmaster1_p & bdb589;
assign a5ee20 = hlock1_p & v84563c | !hlock1_p & b2982f;
assign v845654 = hburst1_p & v84563c | !hburst1_p & !v84563c;
assign a5f86c = hready & a60189 | !hready & a5f86b;
assign c3b82b = hgrant2_p & c3b828 | !hgrant2_p & c3b82a;
assign cea33e = decide_p & cea33d | !decide_p & a57859;
assign af35c3 = jx1_p & af351a | !jx1_p & !af35c2;
assign cea48a = hgrant2_p & cea486 | !hgrant2_p & cea489;
assign c3bc22 = hlock2_p & c3bc20 | !hlock2_p & c3bc21;
assign c3bc51 = hready & b26697 | !hready & !v84563c;
assign b29f3e = hlock0_p & b29f3c | !hlock0_p & b29f3d;
assign b29929 = hgrant1_p & b29928 | !hgrant1_p & b29927;
assign a5f9dd = hmastlock_p & a5f9dc | !hmastlock_p & v84563c;
assign ab05fc = hlock0_p & ab057d | !hlock0_p & !ab05f9;
assign cea86d = hlock2_p & cea86c | !hlock2_p & v84563c;
assign a5f806 = hready & a5f805 | !hready & a5fa1d;
assign a81cad = hlock3_p & a81cac | !hlock3_p & v84563c;
assign c3bce4 = hbusreq3 & c3bcdf | !hbusreq3 & c3bce3;
assign b29f8a = hlock2_p & b29f89 | !hlock2_p & dead2e;
assign a5f7c0 = hready & a5fb12 | !hready & !ab06af;
assign b29aa7 = locked_p & b29d6d | !locked_p & c3bd9a;
assign a5f294 = hbusreq2_p & a5f293 | !hbusreq2_p & v84563c;
assign deac9c = hbusreq3 & deac9b | !hbusreq3 & v84563c;
assign dead55 = hmaster1_p & dead53 | !hmaster1_p & dead54;
assign a5f997 = hbusreq2_p & a5f996 | !hbusreq2_p & !a5fbc0;
assign deae0b = hlock1_p & b26695 | !hlock1_p & !v84563c;
assign b29a51 = hmaster1_p & b29a4c | !hmaster1_p & b29a50;
assign b26696 = hbusreq1_p & b26695 | !hbusreq1_p & !v84563c;
assign a5fc42 = hgrant0_p & a5fbbf | !hgrant0_p & a5fc41;
assign ab0c74 = hbusreq1_p & c3b660 | !hbusreq1_p & deada8;
assign a5f54e = hgrant2_p & a5f511 | !hgrant2_p & a5f54d;
assign a5f371 = hbusreq2 & a5f36c | !hbusreq2 & a5f370;
assign a5f8f4 = hbusreq2_p & a5f8f0 | !hbusreq2_p & !a5fa37;
assign cea14d = hlock0_p & cea14c | !hlock0_p & v84563c;
assign a5f8dd = hmastlock_p & a5f8dc | !hmastlock_p & v84563c;
assign a5fbe0 = start_p & v8e1935 | !start_p & !a5fbdf;
assign dea736 = hmaster1_p & dea735 | !hmaster1_p & v84563c;
assign c3bd9a = hready & dead0c | !hready & v84563c;
assign b2675f = hgrant2_p & b266a3 | !hgrant2_p & !b2675e;
assign af34e7 = hgrant2_p & af3c58 | !hgrant2_p & af34e6;
assign deace0 = hbusreq1_p & b26695 | !hbusreq1_p & !deacdf;
assign deae44 = hbusreq2_p & deadef | !hbusreq2_p & !deacbf;
assign a5edc0 = hready & a5f520 | !hready & c3b6a0;
assign c3bbc1 = decide_p & c3bbc0 | !decide_p & v845660;
assign b29aa0 = hlock2_p & v845660 | !hlock2_p & b29d92;
assign ce9e21 = hlock0_p & cea280 | !hlock0_p & !ce9dc7;
assign cea499 = hready & deae94 | !hready & deae59;
assign b29ff4 = hgrant2_p & b29ff3 | !hgrant2_p & b29f66;
assign dead2c = hlock2_p & v845660 | !hlock2_p & v84563c;
assign b29ebb = locked_p & b29eba | !locked_p & !v84563c;
assign ab0600 = hmaster0_p & ab05f4 | !hmaster0_p & ab05ff;
assign a5fa5b = hready & a5f9dd | !hready & deada8;
assign c3bbf7 = hbusreq1_p & c3bbd2 | !hbusreq1_p & !v84563c;
assign dea6ba = hlock0_p & dea6b9 | !hlock0_p & v84563c;
assign dea767 = locked_p & v84563c | !locked_p & dea766;
assign a5f960 = hlock0_p & a5fb6b | !hlock0_p & a5f6e9;
assign a5e9c2 = hgrant1_p & a5fa1c | !hgrant1_p & a5f18a;
assign dea788 = hbusreq3 & dea786 | !hbusreq3 & dea787;
assign a5fc27 = hlock0_p & v84563c | !hlock0_p & a5fbb3;
assign c3b76f = decide_p & c3b76e | !decide_p & v845660;
assign c3b818 = hmaster0_p & c3b80e | !hmaster0_p & c3b817;
assign a5ef0d = hlock0_p & a5edec | !hlock0_p & a5ef0c;
assign a5ea62 = hbusreq2 & a5ea60 | !hbusreq2 & a5ea61;
assign a5f7d0 = hbusreq2_p & a5f7cf | !hbusreq2_p & v84563c;
assign c3b664 = hlock1_p & v84563c | !hlock1_p & !c3b663;
assign a5f1b0 = hlock1_p & a5fbab | !hlock1_p & v84563c;
assign a5f0db = hlock2_p & a5f0d1 | !hlock2_p & a5f0da;
assign a5fcd0 = hbusreq3 & a5fccf | !hbusreq3 & v84563c;
assign ab074a = hmaster1_p & ab06ed | !hmaster1_p & ab0be3;
assign ab0b7c = hlock0_p & v84563c | !hlock0_p & !b29d51;
assign adaf01 = hbusreq0_p & adaed7 | !hbusreq0_p & adaf00;
assign b2676c = hmaster1_p & b26757 | !hmaster1_p & b266a3;
assign a5f00c = hbusreq2 & a5edfc | !hbusreq2 & a5fcef;
assign c3bc82 = hbusreq3 & c3bc7e | !hbusreq3 & c3bc81;
assign b2992f = hbusreq3 & b2991e | !hbusreq3 & b2992e;
assign dea6ea = hgrant2_p & deae97 | !hgrant2_p & deae9a;
assign a5e9ca = hbusreq2_p & a5e9c8 | !hbusreq2_p & a5e9c9;
assign b26755 = hmaster1_p & b266a8 | !hmaster1_p & b266a3;
assign a9b9d8 = hmaster0_p & v84563c | !hmaster0_p & a9b9d7;
assign cea274 = hready & cea26f | !hready & cea273;
assign ab05c8 = hgrant2_p & ab05c7 | !hgrant2_p & cea15a;
assign a5eaa3 = hgrant0_p & v84563c | !hgrant0_p & a5eaa2;
assign cea1ab = hburst1_p & v84563c | !hburst1_p & !c07311;
assign cea164 = hbusreq2_p & cea163 | !hbusreq2_p & cea162;
assign af3c53 = hbusreq2_p & af3c52 | !hbusreq2_p & af3c51;
assign a5f93b = hbusreq2 & a5f935 | !hbusreq2 & a5f93a;
assign c3b658 = hmaster1_p & c3b654 | !hmaster1_p & c3b657;
assign deadcd = hmaster0_p & deadcc | !hmaster0_p & !v84563c;
assign a5f014 = hbusreq3_p & a5ef33 | !hbusreq3_p & a5f013;
assign a5ee03 = decide_p & a5ede5 | !decide_p & a5ee02;
assign a5f951 = hlock3_p & a5f8f8 | !hlock3_p & a5f950;
assign ce9cd7 = hgrant0_p & cea85f | !hgrant0_p & cea15d;
assign ab0572 = hlock0_p & deada8 | !hlock0_p & !ab0570;
assign ab0739 = hbusreq2_p & ab06a3 | !hbusreq2_p & ab0738;
assign b2999b = hmaster1_p & b29981 | !hmaster1_p & b29e48;
assign af352c = hmastlock_p & b29d6c | !hmastlock_p & v84563c;
assign b29b16 = hgrant2_p & b29a8f | !hgrant2_p & b29a92;
assign ab0c11 = hbusreq3 & ab0c10 | !hbusreq3 & v84563c;
assign a5f90c = hbusreq3 & a5f904 | !hbusreq3 & a5f90b;
assign b29f89 = hlock0_p & b29ec5 | !hlock0_p & c3bce5;
assign ab05a3 = hready & b29824 | !hready & ab05a2;
assign c3b775 = hlock3_p & c3b774 | !hlock3_p & !c3bcbd;
assign a5edd7 = hbusreq2_p & a5edd6 | !hbusreq2_p & a5f567;
assign a5f53f = hbusreq1 & b29941 | !hbusreq1 & v84563c;
assign b2a00a = hmaster1_p & b29e96 | !hmaster1_p & b2a009;
assign a5f1c0 = hmaster0_p & a5f1b9 | !hmaster0_p & a5f1bf;
assign v970437 = hlock2_p & v9703fd | !hlock2_p & v84563c;
assign b2669e = stateA1_p & v84563c | !stateA1_p & v8e1935;
assign ab066f = hlock0_p & b29ebb | !hlock0_p & !dead7f;
assign b29b22 = hlock2_p & v84563c | !hlock2_p & b29b21;
assign ab05c1 = hlock2_p & ab05c0 | !hlock2_p & !ab0593;
assign c3b886 = hmaster1_p & c3b7e6 | !hmaster1_p & c3b885;
assign b2994d = hlock1_p & deac51 | !hlock1_p & !c3b6a5;
assign af3c81 = hlock2_p & af3c80 | !hlock2_p & af3c7f;
assign ce9d79 = hmaster0_p & ce9d72 | !hmaster0_p & ce9d2e;
assign deacbc = hbusreq1_p & v84563c | !hbusreq1_p & v84565a;
assign ab0b85 = hbusreq3 & ab0b84 | !hbusreq3 & cea15a;
assign d40d43 = hlock0_p & d40d3e | !hlock0_p & d40d42;
assign a5eb50 = hbusreq0 & a5ea9c | !hbusreq0 & !v84563c;
assign c3b66a = hlock1_p & c3bbd2 | !hlock1_p & deadb1;
assign a5fc73 = hbusreq3 & a5fc72 | !hbusreq3 & v84563c;
assign b29973 = hgrant2_p & b2996c | !hgrant2_p & b29972;
assign a5edfc = locked_p & v845641 | !locked_p & a5edf6;
assign a5f3a2 = hlock0_p & a5f39f | !hlock0_p & a5f3a1;
assign a5f25a = hlock3_p & a5f256 | !hlock3_p & a5f950;
assign cea341 = locked_p & v84563c | !locked_p & deacec;
assign ce9d52 = hlock0_p & cea325 | !hlock0_p & !cea17a;
assign a5fbf4 = hlock2_p & a5fbea | !hlock2_p & a5fbf3;
assign a5ee86 = locked_p & a5f369 | !locked_p & a5f39e;
assign a5efc8 = hmaster0_p & a5efc7 | !hmaster0_p & a5eec8;
assign bdb5a6 = hmaster1_p & bdb598 | !hmaster1_p & bdb5a5;
assign c3b7a5 = hlock0_p & c3bcee | !hlock0_p & v845660;
assign cea469 = hbusreq2_p & cea468 | !hbusreq2_p & cea37b;
assign cea2a3 = hbusreq2_p & cea2a2 | !hbusreq2_p & v84563c;
assign a5f8d6 = hready & a5f8d1 | !hready & a5f8d5;
assign a5fb97 = hready & a5f9dd | !hready & !a5fb8c;
assign a5fce5 = locked_p & a5fce4 | !locked_p & v84563c;
assign a5f8e5 = hready & a5f8e4 | !hready & a5f8d5;
assign a5ea2f = decide_p & a5ea1e | !decide_p & a5ea2e;
assign cea237 = hbusreq2_p & cea236 | !hbusreq2_p & v84563c;
assign b29fee = hbusreq3 & b29fed | !hbusreq3 & b29ed5;
assign a5f196 = hbusreq2 & a5f195 | !hbusreq2 & a5fa6b;
assign a5f1ac = hbusreq1 & a5f9dd | !hbusreq1 & a5fc48;
assign a5ea6c = hgrant2_p & a5ea68 | !hgrant2_p & a5ea6b;
assign bdb598 = locked_p & v84563c | !locked_p & !v84565a;
assign c3b6a3 = hbusreq2_p & c3b699 | !hbusreq2_p & !c3b6a1;
assign a5fae8 = hbusreq3 & a5fae6 | !hbusreq3 & a5fae7;
assign c3b769 = hbusreq2_p & c3b768 | !hbusreq2_p & !c3b6a1;
assign deae11 = locked_p & deae02 | !locked_p & !deae0b;
assign ab0c75 = hgrant1_p & c3b660 | !hgrant1_p & ab0c74;
assign af350e = hready_p & af350a | !hready_p & af350d;
assign a5fc2f = hbusreq2 & a5fc2e | !hbusreq2 & a5fc2d;
assign bdb5b0 = hready_p & bdb5ae | !hready_p & bdb5af;
assign a5fc88 = hready & a5fc84 | !hready & a5fc87;
assign b26776 = hmaster0_p & b26775 | !hmaster0_p & b2671b;
assign ab0b8e = hlock2 & ab0b8c | !hlock2 & ab0b8d;
assign dea759 = hmaster1_p & dea758 | !hmaster1_p & !dea6f4;
assign a5fbc8 = hlock0_p & v84563c | !hlock0_p & a5fbc7;
assign a5fbb0 = hlock1_p & a5fbab | !hlock1_p & a5fbaf;
assign b299f5 = hready_p & b29cba | !hready_p & b299f4;
assign a5faaa = hbusreq1_p & a60193 | !hbusreq1_p & !a6016f;
assign a5fc94 = hbusreq0 & a5fc81 | !hbusreq0 & !a5fc93;
assign a5f985 = hlock0_p & a5f984 | !hlock0_p & v84563c;
assign cea15a = hlock0_p & v84563c | !hlock0_p & v845660;
assign cea483 = hlock0_p & cea482 | !hlock0_p & cea3ea;
assign cea1c4 = hbusreq2_p & cea149 | !hbusreq2_p & cea85d;
assign ce9e28 = hgrant3_p & ce9ddd | !hgrant3_p & ce9e27;
assign ce9cd4 = hready_p & cea862 | !hready_p & ce9cd3;
assign c3b7cc = hlock0_p & c3bd2d | !hlock0_p & !deadc4;
assign ab058e = hbusreq2_p & ab058a | !hbusreq2_p & ab058d;
assign ab0c09 = hlock0_p & v84563c | !hlock0_p & !ab0c08;
assign c3b851 = hgrant2_p & c3b84d | !hgrant2_p & c3b850;
assign ab05b9 = hmaster1_p & ab05ae | !hmaster1_p & ab05b8;
assign c3b61a = hgrant2_p & c3b616 | !hgrant2_p & c3b619;
assign ab06b8 = hlock0_p & b29f51 | !hlock0_p & !ab06b7;
assign c3b6dd = hlock1_p & v84563c | !hlock1_p & !dead76;
assign deae58 = hmaster0_p & deae57 | !hmaster0_p & v845660;
assign c3b6d6 = hlock0_p & c3bbbb | !hlock0_p & !c3b625;
assign a5ea97 = hbusreq0 & a5ea96 | !hbusreq0 & v84563c;
assign a5f835 = hgrant1_p & a5f834 | !hgrant1_p & a5f833;
assign a5f40e = hlock0_p & a5f3f8 | !hlock0_p & a5f40d;
assign a5f8e4 = hlock1_p & a5fbab | !hlock1_p & !a5f8e3;
assign a5ef26 = hgrant2_p & a5ef25 | !hgrant2_p & v84563c;
assign b29a9e = decide_p & b29a9d | !decide_p & v84563c;
assign c3b7f9 = hbusreq2_p & c3b7f8 | !hbusreq2_p & c3b7e6;
assign a5fc6b = hlock1_p & v84563c | !hlock1_p & a5fc6a;
assign b26742 = hmaster1_p & b2670b | !hmaster1_p & b2670f;
assign a9b9df = hmaster1_p & a9b9de | !hmaster1_p & !v84563c;
assign c3bcff = hbusreq3 & c3bcfe | !hbusreq3 & !c3bcb3;
assign b29d9d = hmaster1_p & c3bceb | !hmaster1_p & b29d9c;
assign a5ee79 = hlock2_p & a5ee72 | !hlock2_p & a5ee78;
assign ab0c31 = hready & v84563c | !hready & v84565a;
assign cea1c3 = hbusreq3 & cea1b8 | !hbusreq3 & cea1c2;
assign b29ffd = hlock0_p & b29ffc | !hlock0_p & !c3bcef;
assign b2678e = hbusreq3_p & b26769 | !hbusreq3_p & !b2678d;
assign ab0630 = hgrant2_p & ab062a | !hgrant2_p & ab062f;
assign ab0c91 = hmaster0_p & ab0c88 | !hmaster0_p & ab0c90;
assign a5fa8a = hready & a60168 | !hready & v84563c;
assign b2a003 = hlock0_p & b2a002 | !hlock0_p & c3bd8d;
assign a5fd35 = hlock0_p & v84563c | !hlock0_p & a5fd34;
assign a5fc02 = hready & a5fb8a | !hready & a5fc01;
assign b29e58 = decide_p & b29e56 | !decide_p & b29e57;
assign c3b7fc = hbusreq2_p & c3b7fb | !hbusreq2_p & c3b7e6;
assign a5ea25 = hbusreq0 & a5ea24 | !hbusreq0 & v84563c;
assign a5f52c = hready & a5f529 | !hready & a5f52b;
assign a5ee96 = hbusreq2 & a5ee95 | !hbusreq2 & a5fbc0;
assign adaf0b = hgrant2_p & adaf0a | !hgrant2_p & v84563c;
assign deacff = hlock2_p & deacfd | !hlock2_p & deacfe;
assign cea459 = hlock2_p & cea394 | !hlock2_p & cea3aa;
assign a5fcae = hmaster1_p & v84563c | !hmaster1_p & a5fcad;
assign a5fa1b = hlock1_p & a60187 | !hlock1_p & a5fa1a;
assign deae93 = hbusreq2_p & deae92 | !hbusreq2_p & !v84563c;
assign dea75d = hready_p & dea739 | !hready_p & dea75c;
assign a5f3d8 = locked_p & v84563c | !locked_p & !a5f3d7;
assign ab0c79 = hlock2 & ab0b17 | !hlock2 & ab0c78;
assign deadcc = hmaster1_p & deadcb | !hmaster1_p & !v84563c;
assign b29f5c = hbusreq2_p & b29f5a | !hbusreq2_p & v84563c;
assign ab06d4 = hbusreq2_p & ab06d3 | !hbusreq2_p & ab06b5;
assign cea450 = hmaster1_p & cea449 | !hmaster1_p & cea44f;
assign a5f0a8 = hbusreq0_p & a5fc6d | !hbusreq0_p & v84563c;
assign dea6d7 = hgrant2_p & dea6d3 | !hgrant2_p & dea6d6;
assign c3bd5d = hlock1_p & v84563c | !hlock1_p & !deada8;
assign ab0634 = hgrant2_p & ab05f6 | !hgrant2_p & ab0633;
assign dea6c9 = hgrant1_p & deada8 | !hgrant1_p & deae74;
assign c3bd69 = hlock2_p & c3bd5f | !hlock2_p & v84563c;
assign c3b84a = hlock0_p & c3bdd6 | !hlock0_p & deadba;
assign af3491 = hmaster1_p & d40d33 | !hmaster1_p & af3c7f;
assign b29d86 = hlock2_p & b29d80 | !hlock2_p & b29d85;
assign b29a85 = hlock0_p & b29a84 | !hlock0_p & !deada8;
assign a81cd5 = hbusreq2_p & a81cd4 | !hbusreq2_p & v84563c;
assign b2996a = hlock2 & b29967 | !hlock2 & b29969;
assign ab05ea = hmaster1_p & ab05e5 | !hmaster1_p & ab05e9;
assign a9b9e3 = hmaster0_p & v84563c | !hmaster0_p & a9b9e2;
assign ab06e0 = hlock0_p & b29f99 | !hlock0_p & !dead41;
assign b29f80 = hgrant2_p & b29f7e | !hgrant2_p & b29f7f;
assign b299af = hbusreq3 & b299ae | !hbusreq3 & b298b1;
assign b8acf4 = jx2_p & b8acd7 | !jx2_p & b8acf3;
assign ab0bec = hbusreq2_p & ab0bea | !hbusreq2_p & ab0b0e;
assign a5f6ef = locked_p & a5f6ee | !locked_p & v845641;
assign b29cd4 = hlock2_p & v84563c | !hlock2_p & deacab;
assign cea3b8 = hbusreq1_p & deaca1 | !hbusreq1_p & cea3b7;
assign c3bdc2 = hbusreq2_p & c3bdc1 | !hbusreq2_p & cea18d;
assign c3b700 = hlock2_p & c3b631 | !hlock2_p & !c3b625;
assign c3b780 = jx1_p & c3b772 | !jx1_p & c3b77f;
assign a5fb14 = hlock2 & a5f9e8 | !hlock2 & a5fb13;
assign cea3a7 = hbusreq2_p & cea3a6 | !hbusreq2_p & cea3a5;
assign ab0714 = hbusreq2_p & ab0713 | !hbusreq2_p & ab0712;
assign a5fb90 = locked_p & a5fb8f | !locked_p & v84563c;
assign a5ea55 = hlock0_p & a5ea53 | !hlock0_p & a5ea54;
assign a5efcd = hgrant0_p & a5efc8 | !hgrant0_p & a5efcc;
assign a5fbae = hmastlock_p & a5fbad | !hmastlock_p & !v84563c;
assign ab0741 = hbusreq2_p & ab0740 | !hbusreq2_p & !b29b1c;
assign a5f2e9 = hbusreq2 & a5f2e5 | !hbusreq2 & a5f2e8;
assign deae15 = hgrant2_p & dead39 | !hgrant2_p & deae14;
assign cea41d = hlock2_p & cea41c | !hlock2_p & cea3fb;
assign b29924 = stateG10_1_p & v84563c | !stateG10_1_p & b29923;
assign ab0650 = hlock3_p & ab064c | !hlock3_p & ab064f;
assign ab0cac = hlock0_p & ab0cab | !hlock0_p & ab0c89;
assign a5eebf = hbusreq1_p & a5fc8c | !hbusreq1_p & !v84563c;
assign c3be03 = hbusreq2_p & c3be02 | !hbusreq2_p & c3bc6e;
assign af34ed = decide_p & af34e2 | !decide_p & af34ec;
assign deac57 = hlock1_p & deac51 | !hlock1_p & deac56;
assign a5ee4f = locked_p & a5ee4e | !locked_p & a5ee38;
assign a60194 = hlock1_p & a60193 | !hlock1_p & v84563c;
assign c3bc06 = hbusreq2_p & c3bc05 | !hbusreq2_p & !v84563c;
assign a5f8da = hburst0_p & c07311 | !hburst0_p & a5f8d9;
assign b266df = hgrant1_p & b266da | !hgrant1_p & b266a1;
assign af3c32 = hmaster1_p & af3c31 | !hmaster1_p & !v84563c;
assign a5f253 = hbusreq2_p & a5f252 | !hbusreq2_p & !v84563c;
assign cea40c = hlock0_p & cea40b | !hlock0_p & cea3cd;
assign a5fc2a = hlock2 & a5fc27 | !hlock2 & a5fc29;
assign ab0b64 = locked_p & ab0b63 | !locked_p & !v84563c;
assign b2673e = hgrant2_p & b2673a | !hgrant2_p & b2673d;
assign a5ede3 = hmaster1_p & a5edd2 | !hmaster1_p & a5ede2;
assign ab0598 = locked_p & v84563c | !locked_p & !b2997c;
assign b299df = hlock2 & b299dd | !hlock2 & b299de;
assign af34d1 = hmaster0_p & af34ce | !hmaster0_p & af34d0;
assign b2671d = hlock2_p & b266a9 | !hlock2_p & !b26695;
assign a5f46e = hlock1_p & a5f46d | !hlock1_p & a5f436;
assign b26727 = hbusreq1_p & b26694 | !hbusreq1_p & !b2669f;
assign c3b8b2 = hgrant2_p & c3b7de | !hgrant2_p & c3b8b1;
assign c3b68a = hbusreq2_p & c3b689 | !hbusreq2_p & !c3b686;
assign c3bc15 = hlock0_p & c3bc09 | !hlock0_p & !deac86;
assign a5f2e4 = locked_p & v84563c | !locked_p & a5f2e3;
assign cea154 = hlock2_p & cea153 | !hlock2_p & v84563c;
assign a5fb5e = hlock0_p & v84563c | !hlock0_p & a5fb5d;
assign deae37 = hbusreq2_p & dead95 | !hbusreq2_p & v845644;
assign c3b720 = hlock0_p & c3b71c | !hlock0_p & !c3b71f;
assign a5fc4a = hlock0_p & a5fc49 | !hlock0_p & v84563c;
assign b29e69 = hlock2_p & b29d33 | !hlock2_p & b29e68;
assign a5ee8e = hlock0_p & a5ee8d | !hlock0_p & !a5ee28;
assign v97044c = hmaster0_p & v970448 | !hmaster0_p & v97044b;
assign a5f1c9 = locked_p & v84563c | !locked_p & a5f739;
assign ab0c00 = hlock0_p & v84563c | !hlock0_p & !ab0bff;
assign b29d4f = decide_p & b29d4e | !decide_p & v84563c;
assign a5fc7f = locked_p & a5fc7e | !locked_p & a5fc70;
assign c3b7d3 = hbusreq3 & c3b7c3 | !hbusreq3 & c3b7d2;
assign a60145 = hbusreq3 & a60144 | !hbusreq3 & v84563c;
assign b29edc = hbusreq2_p & b29edb | !hbusreq2_p & v84563c;
assign a5f9cb = hmaster1_p & v84563c | !hmaster1_p & a5f9ca;
assign a5ea5f = hlock2_p & a5ea5d | !hlock2_p & a5ea5e;
assign a5efbb = hbusreq2 & a5efba | !hbusreq2 & a5ee68;
assign a5f07a = hlock2_p & a5f077 | !hlock2_p & !a5f079;
assign a5ee34 = hbusreq0 & a5ee1a | !hbusreq0 & !a5ee33;
assign ab06b1 = hbusreq0_p & deacb7 | !hbusreq0_p & ab06b0;
assign a5ef8f = hmaster1_p & a5ef80 | !hmaster1_p & a5ef8e;
assign b2994c = hbusreq2_p & b29944 | !hbusreq2_p & b2994b;
assign cea41f = hready & deae94 | !hready & cea29f;
assign a5f32e = hgrant2_p & a5f326 | !hgrant2_p & a5f32d;
assign ab054f = hbusreq2_p & ab054e | !hbusreq2_p & ab054d;
assign a5eaf1 = hbusreq2_p & a5eaea | !hbusreq2_p & a5eae5;
assign ab06ba = hlock1_p & v84565a | !hlock1_p & ab06b9;
assign c3b896 = decide_p & c3b895 | !decide_p & v845660;
assign ab05b2 = hlock2 & ab051a | !hlock2 & ab05b1;
assign ab064e = hmaster0_p & ab0bbb | !hmaster0_p & ab064d;
assign c3b8b8 = hbusreq3_p & c3b873 | !hbusreq3_p & !c3b8b7;
assign deacf7 = hmastlock_p & deacf6 | !hmastlock_p & v84563c;
assign c3bdd7 = hlock0_p & c3bdd5 | !hlock0_p & !c3bdd6;
assign a5f477 = hbusreq3 & a5f422 | !hbusreq3 & !a5f476;
assign a5f83e = start_p & a81ca6 | !start_p & !v8c6449;
assign cea1b2 = hbusreq1_p & cea1b1 | !hbusreq1_p & !v84563c;
assign dead98 = hmaster1_p & dead91 | !hmaster1_p & dead97;
assign cea36d = hmaster1_p & cea36c | !hmaster1_p & !cea289;
assign ab0565 = hlock2 & ab0563 | !hlock2 & ab0564;
assign af3530 = hmaster1_p & af352d | !hmaster1_p & af352f;
assign a5ee54 = hbusreq1 & a5ee53 | !hbusreq1 & !v84563c;
assign bdb5a9 = hmaster0_p & bdb5a6 | !hmaster0_p & !bdb5a8;
assign a5ea4e = hbusreq0_p & a5fc5b | !hbusreq0_p & a5ea4d;
assign a5f9a8 = hbusreq2 & a5f9a4 | !hbusreq2 & a5f9a7;
assign af34b5 = hlock1_p & af3c49 | !hlock1_p & af3c6a;
assign deae06 = hlock0_p & deae05 | !hlock0_p & v84563c;
assign a5ee9b = hready & a5ee43 | !hready & !c3b6f8;
assign a5efa0 = hbusreq0_p & a5ee24 | !hbusreq0_p & a5ee68;
assign c3bd03 = hlock2_p & c3bd02 | !hlock2_p & v84563c;
assign a5f94e = hgrant2_p & a5f94b | !hgrant2_p & a5f94d;
assign a5fd14 = hbusreq3 & a5fd13 | !hbusreq3 & v84563c;
assign deac1f = hlock2_p & deac1e | !hlock2_p & v84565a;
assign a5f6d3 = hbusreq2_p & a5f6d2 | !hbusreq2_p & v84563c;
assign af3c43 = decide_p & af3c34 | !decide_p & v8567b4;
assign a5ea48 = hbusreq2_p & a5ea47 | !hbusreq2_p & a5ea41;
assign cea194 = hgrant0_p & cea85f | !hgrant0_p & cea193;
assign a5ee9f = hlock0_p & a5ee9e | !hlock0_p & a5ee4f;
assign d40d55 = hmaster1_p & d40d53 | !hmaster1_p & d40d54;
assign ce9d1f = hbusreq2_p & cea25a | !hbusreq2_p & cea259;
assign ab0b48 = hbusreq2_p & ab0b46 | !hbusreq2_p & ab0b23;
assign b298af = hlock0_p & b298ae | !hlock0_p & !v84563c;
assign a5f493 = hlock1_p & v84565a | !hlock1_p & b29919;
assign cea3bd = stateG10_1_p & deacb4 | !stateG10_1_p & cea3bc;
assign a5f6f3 = locked_p & a5f6f2 | !locked_p & a5fb6a;
assign a5f918 = hbusreq1 & deac5b | !hbusreq1 & a5f917;
assign a5edb8 = hready & a5f4e4 | !hready & a5edb7;
assign a5ee6d = hbusreq0_p & a5ee39 | !hbusreq0_p & a5ee66;
assign v970401 = decide_p & v970400 | !decide_p & v9703ff;
assign a5fb9b = hlock2_p & a5fb93 | !hlock2_p & a5fb9a;
assign a5fc09 = hmastlock_p & a5fc08 | !hmastlock_p & !v84563c;
assign adaec8 = hgrant1_p & adaec7 | !hgrant1_p & adaec4;
assign c3bbe8 = hlock0_p & c3bbe2 | !hlock0_p & deacaa;
assign af3537 = hmaster0_p & af3536 | !hmaster0_p & af3534;
assign b29f53 = hlock1_p & v84565a | !hlock1_p & deac52;
assign c3b623 = locked_p & c3b622 | !locked_p & c3bbba;
assign c3b6b4 = hbusreq2_p & c3b6b2 | !hbusreq2_p & c3b6b0;
assign bdb586 = hlock2_p & bdb585 | !hlock2_p & v84565a;
assign cea191 = hgrant2_p & cea159 | !hgrant2_p & !cea190;
assign a5f6da = hmaster1_p & a5f6d8 | !hmaster1_p & a5f6d9;
assign b29e4f = hlock2_p & b29e4e | !hlock2_p & v84563c;
assign adaefb = hmaster1_p & adaec4 | !hmaster1_p & adaeca;
assign a5efa4 = hmaster1_p & a5ee0d | !hmaster1_p & a5efa3;
assign a5f296 = hmaster1_p & a5f295 | !hmaster1_p & a5f73e;
assign ab061e = hlock0_p & v84563c | !hlock0_p & !ab061d;
assign b2a016 = hgrant2_p & b2a015 | !hgrant2_p & b29f5c;
assign ab0cca = hmaster0_p & ab0cc9 | !hmaster0_p & ab0c64;
assign ab055b = stateG10_1_p & v84563c | !stateG10_1_p & ab055a;
assign a81d05 = decide_p & v84563c | !decide_p & a81d04;
assign b29d06 = hbusreq3 & b29d04 | !hbusreq3 & b29d05;
assign deadfc = locked_p & v84563c | !locked_p & !dead93;
assign b26722 = hlock2_p & b26721 | !hlock2_p & b266a8;
assign ab0b4f = hlock3_p & ab0b34 | !hlock3_p & ab0b4e;
assign dead05 = hlock2_p & dead04 | !hlock2_p & deace1;
assign dea6c2 = hbusreq2_p & dea6bb | !hbusreq2_p & v84563c;
assign a5f8bd = hgrant1_p & v84565a | !hgrant1_p & a5f8bc;
assign af3c24 = hmaster0_p & b8acdf | !hmaster0_p & af3c23;
assign a5f561 = hlock0_p & a5f560 | !hlock0_p & a5f55b;
assign ab0c45 = hlock2 & v84563c | !hlock2 & ab0c44;
assign c3b72f = hready & v845648 | !hready & !v84563c;
assign b29aa6 = hbusreq2_p & b29aa5 | !hbusreq2_p & b29aa4;
assign a5ea57 = hbusreq1_p & a5fc09 | !hbusreq1_p & a5fc84;
assign a5f94a = hbusreq2_p & a5f949 | !hbusreq2_p & v845644;
assign af358c = hmaster1_p & v84563c | !hmaster1_p & af358b;
assign c3b659 = hmaster0_p & c3b64e | !hmaster0_p & c3b658;
assign cea435 = hlock0_p & cea434 | !hlock0_p & cea3cd;
assign af3541 = hlock1_p & af352c | !hlock1_p & af3540;
assign b29fb7 = hlock0_p & c3bcf8 | !hlock0_p & c3bd8e;
assign c3b68c = hbusreq2_p & c3b66e | !hbusreq2_p & c3b66c;
assign ab0bdd = hmaster0_p & ab0bd3 | !hmaster0_p & ab0bdc;
assign cea39f = hlock0_p & cea39d | !hlock0_p & cea39e;
assign c3bc7f = hlock0_p & v845648 | !hlock0_p & cea18d;
assign c3b6cd = hlock2_p & c3b6cc | !hlock2_p & c3b6b1;
assign ab0ceb = hlock0_p & v84563c | !hlock0_p & c3bcf0;
assign d40d2f = stateG2_p & v84563c | !stateG2_p & bfbd19;
assign b26713 = hlock0_p & b266ad | !hlock0_p & b266a0;
assign cea38c = hlock2_p & cea38b | !hlock2_p & cea38a;
assign a5e9f7 = hlock2 & a5e9f2 | !hlock2 & a5e9f6;
assign deac99 = hbusreq2_p & deac89 | !hbusreq2_p & deac88;
assign c3bcd0 = hmaster1_p & c3bcce | !hmaster1_p & c3bccf;
assign a5f161 = hbusreq2_p & a5f15d | !hbusreq2_p & a5f154;
assign b299a2 = hlock2_p & b299a1 | !hlock2_p & b2998e;
assign d40d3d = hgrant1_p & d40d3b | !hgrant1_p & !d40d3c;
assign a5eeb0 = hbusreq2_p & a5eeaf | !hbusreq2_p & a5ee78;
assign b29917 = hlock1_p & deadde | !hlock1_p & !b29916;
assign ab071d = hgrant2_p & ab0719 | !hgrant2_p & ab071c;
assign a5f935 = hlock2 & a5f92f | !hlock2 & a5f934;
assign b2671f = hlock1_p & v84563c | !hlock1_p & !b26695;
assign b29d4d = hmaster0_p & b29d2c | !hmaster0_p & b29d4c;
assign ab0584 = hmaster0_p & ab057a | !hmaster0_p & ab0583;
assign dead7d = hlock1_p & v84563c | !hlock1_p & !dead7c;
assign b29d93 = hlock0_p & b29d82 | !hlock0_p & !v84563c;
assign a5f70c = locked_p & a5f70b | !locked_p & v84563c;
assign b29ec7 = hlock0_p & b29ec5 | !hlock0_p & b29ec6;
assign ab064b = hready_p & ab0ad0 | !hready_p & ab064a;
assign cea152 = locked_p & cea151 | !locked_p & b26697;
assign a5f975 = locked_p & a5f974 | !locked_p & a5fb6a;
assign a6016e = start_p & a6016a | !start_p & a6016d;
assign cea2ec = hbusreq2_p & cea2eb | !hbusreq2_p & cea85d;
assign cea366 = hlock0_p & cea365 | !hlock0_p & v84563c;
assign a5fc92 = hbusreq0_p & a5fc89 | !hbusreq0_p & a5fc91;
assign ce9d4f = hmaster1_p & ce9d4e | !hmaster1_p & cea15d;
assign v845668 = hgrant3_p & v84563c | !hgrant3_p & !v84563c;
assign bfbd18 = stateG3_0_p & v84563c | !stateG3_0_p & !v845674;
assign cea3a0 = hlock2_p & cea39f | !hlock2_p & cea39e;
assign b29d29 = hbusreq3 & v84563c | !hbusreq3 & b29cd5;
assign ab06ec = hbusreq2_p & ab0679 | !hbusreq2_p & ab06eb;
assign d40d93 = hready_p & d40d8f | !hready_p & d40d92;
assign v970458 = decide_p & v97042d | !decide_p & v970456;
assign c3b711 = decide_p & c3b710 | !decide_p & v845660;
assign a5f154 = hlock0_p & a5f153 | !hlock0_p & v84563c;
assign a5fd1b = hready_p & a5fcc4 | !hready_p & a5fd1a;
assign v97044e = decide_p & v97043c | !decide_p & v97044d;
assign b2998b = hlock2 & b29987 | !hlock2 & b2998a;
assign b26772 = hready_p & b2676e | !hready_p & b26771;
assign c3bcf7 = hmaster0_p & c3bced | !hmaster0_p & c3bcf6;
assign deae4a = hgrant3_p & deae49 | !hgrant3_p & !v84563c;
assign a5f70d = hlock0_p & a5f70a | !hlock0_p & !a5f70c;
assign deacdb = decide_p & deacda | !decide_p & v84563c;
assign b299e1 = hbusreq2_p & b299e0 | !hbusreq2_p & !b299df;
assign a5fad3 = hlock0_p & v84563c | !hlock0_p & a5fad2;
assign c3bceb = hbusreq2_p & c3bcea | !hbusreq2_p & v84563c;
assign a5fd0b = hgrant2_p & a5fd0a | !hgrant2_p & a5fcd0;
assign c3bd4e = hbusreq2_p & c3bd4d | !hbusreq2_p & deacaa;
assign c3b7fe = hmaster1_p & c3b7fd | !hmaster1_p & !c3bc21;
assign a5fb8c = hmastlock_p & b29f03 | !hmastlock_p & !v84563c;
assign ab0682 = hmaster1_p & ab0680 | !hmaster1_p & ab0681;
assign af3c48 = start_p & v84563c | !start_p & !v856b00;
assign a5f528 = hlock1_p & a6016f | !hlock1_p & !a5f4c7;
assign cea16c = hready & dead18 | !hready & b266a0;
assign b29991 = hlock0_p & b29990 | !hlock0_p & !v84563c;
assign a5f4e7 = hgrant1_p & a5f4e6 | !hgrant1_p & a5f4e5;
assign c3bd88 = hbusreq2_p & c3bd87 | !hbusreq2_p & c3bc5c;
assign a5f36a = hbusreq1 & c3b624 | !hbusreq1 & v84563c;
assign ab0baa = hbusreq0_p & b29d82 | !hbusreq0_p & !b29d8a;
assign a5f581 = hready & a5f57c | !hready & a5f580;
assign ab0b0d = hbusreq2_p & ab0b0c | !hbusreq2_p & ab0af6;
assign ab0bf4 = hmaster1_p & ab0bf1 | !hmaster1_p & !ab0bf3;
assign a5f4ee = hready & v84563c | !hready & a5f4ed;
assign c3b817 = hmaster1_p & c3b816 | !hmaster1_p & c3bc71;
assign c3bddc = hbusreq3 & c3bddb | !hbusreq3 & c3bdd9;
assign cea3dc = hready & cea3db | !hready & cea273;
assign cea888 = hlock0_p & cea884 | !hlock0_p & !cea887;
assign b29ed5 = hbusreq2_p & dead3d | !hbusreq2_p & v84563c;
assign c3b6bf = hready & c3b6bd | !hready & c3b6be;
assign cea46d = hlock2_p & cea46c | !hlock2_p & cea39b;
assign a5f1f0 = hbusreq1 & a5fbd7 | !hbusreq1 & !a5f1ef;
assign a5ee08 = hbusreq2 & a5ee06 | !hbusreq2 & a5ee07;
assign dea6cd = hbusreq2_p & dea6cc | !hbusreq2_p & !deada8;
assign a5ee98 = hbusreq2_p & a5ee97 | !hbusreq2_p & a5ee3e;
assign cea0bd = hlock0_p & cea0bc | !hlock0_p & v84563c;
assign ab05ab = hlock0_p & v84563c | !hlock0_p & !b29993;
assign af3c69 = stateA1_p & v84563c | !stateA1_p & c0730a;
assign b2a012 = hbusreq2_p & b2a010 | !hbusreq2_p & !v84563c;
assign a5ea7b = locked_p & a5fbfd | !locked_p & a5f6e9;
assign dea7a2 = hmaster1_p & dea735 | !hmaster1_p & dead54;
assign a5fba0 = stateA1_p & a5fb9d | !stateA1_p & !a5fb9f;
assign af3c41 = decide_p & af3c27 | !decide_p & v8567b4;
assign c3b629 = hbusreq2_p & c3b628 | !hbusreq2_p & c3b627;
assign cea17b = hbusreq3 & cea17a | !hbusreq3 & !v845660;
assign deade2 = hbusreq2_p & deade1 | !hbusreq2_p & !v84563c;
assign ab075c = decide_p & ab075b | !decide_p & !v845662;
assign a5f531 = hbusreq1 & a5f530 | !hbusreq1 & v84563c;
assign c3bc38 = hlock2_p & deada8 | !hlock2_p & v84563c;
assign a5fc0c = start_p & a6016a | !start_p & a5fbac;
assign b29f1d = hready & b29f1c | !hready & v84563c;
assign cea0ef = hgrant2_p & cea0e9 | !hgrant2_p & cea0ee;
assign c3b6ca = hgrant2_p & c3b6c2 | !hgrant2_p & c3b6c9;
assign a5f3af = hlock0_p & a5f39e | !hlock0_p & a5f36b;
assign af34ad = hbusreq2_p & af34ac | !hbusreq2_p & af3c4c;
assign cea19b = hbusreq2_p & cea19a | !hbusreq2_p & !v84563c;
assign a5f3ce = hready & a5f3cb | !hready & a5f3cd;
assign dead30 = hmaster1_p & dead2d | !hmaster1_p & dead2f;
assign deacb7 = hlock1_p & deaca1 | !hlock1_p & deacb6;
assign a5f6f5 = locked_p & a5f6f4 | !locked_p & a5f6e9;
assign cea292 = hlock1_p & v84563c | !hlock1_p & !cea291;
assign c3bd85 = hbusreq2_p & c3bd84 | !hbusreq2_p & c3bc5c;
assign a5ea3e = hbusreq2_p & a5ea3d | !hbusreq2_p & a5ea3c;
assign adaf1c = hbusreq3_p & adaf11 | !hbusreq3_p & adaf1b;
assign af35b1 = hmaster0_p & af35b0 | !hmaster0_p & af358e;
assign a5ee72 = hbusreq2 & a5ee6f | !hbusreq2 & a5ee71;
assign cea0bf = hlock0_p & c98b95 | !hlock0_p & !v84563c;
assign c3b6ec = hlock2_p & c3b627 | !hlock2_p & !c3b647;
assign a5f1f9 = hbusreq2 & a5f1f5 | !hbusreq2 & a5f1f8;
assign a5f214 = hbusreq2_p & a5f213 | !hbusreq2_p & v84563c;
assign a5f795 = hbusreq1_p & v84565a | !hbusreq1_p & a60172;
assign dea74f = hbusreq3 & dea74d | !hbusreq3 & dea74e;
assign b8ace8 = hgrant0_p & b8acd9 | !hgrant0_p & b8ace7;
assign b29ed4 = hbusreq2_p & b29ed3 | !hbusreq2_p & v84563c;
assign ab0622 = hmaster1_p & ab061c | !hmaster1_p & ab0621;
assign dead52 = hgrant3_p & deacdc | !hgrant3_p & !dead51;
assign aa0e0b = jx0_p & aa0e0a | !jx0_p & v868347;
assign ab0c29 = hbusreq3 & ab0c28 | !hbusreq3 & v84564a;
assign a5fa25 = hlock0_p & v845641 | !hlock0_p & ab0c31;
assign cea3ee = hbusreq3 & cea3d0 | !hbusreq3 & cea3ed;
assign af3548 = hlock1_p & af352c | !hlock1_p & af3547;
assign bdb596 = hmaster0_p & bdb58a | !hmaster0_p & bdb595;
assign c3b875 = hmaster1_p & c3b874 | !hmaster1_p & c3b7ae;
assign b266ae = locked_p & v84563c | !locked_p & b266a0;
assign a5f1fd = hmaster1_p & a5f1ed | !hmaster1_p & a5f1fc;
assign a5e9be = hlock2 & a5e9b5 | !hlock2 & a5e9bd;
assign a5f2dd = hmaster0_p & a5f2dc | !hmaster0_p & !a5f95c;
assign a5ef35 = hready & a5f38c | !hready & !v845648;
assign c3b686 = hready & c3b684 | !hready & c3b685;
assign b299d9 = hlock2_p & v84563c | !hlock2_p & b299d8;
assign a5ec18 = hmaster1_p & a5f6db | !hmaster1_p & a5e9ce;
assign a5efdf = hlock2 & a5efde | !hlock2 & a5f549;
assign a60165 = hburst0_p & c06d34 | !hburst0_p & a60164;
assign dead74 = stateA1_p & dead31 | !stateA1_p & !c07311;
assign a5f1d0 = hbusreq1_p & a5fc78 | !hbusreq1_p & a5f9dd;
assign ce9d27 = hbusreq2_p & cea286 | !hbusreq2_p & cea283;
assign b29e6b = hbusreq2_p & b29e69 | !hbusreq2_p & !v84563c;
assign af3566 = hlock0_p & af352c | !hlock0_p & af3532;
assign a5eea9 = hlock2_p & a5eea8 | !hlock2_p & a5ee63;
assign c3bd95 = hlock2_p & c3bd94 | !hlock2_p & v845660;
assign d40d6a = hlock0_p & d40d2c | !hlock0_p & d40d69;
assign c3b7d5 = hbusreq2_p & c3b7d1 | !hbusreq2_p & c3b7cc;
assign a5ea77 = hbusreq2_p & a5ea76 | !hbusreq2_p & a5ea75;
assign a5eaeb = hbusreq2_p & a5eaea | !hbusreq2_p & !a5eae9;
assign b266dc = hlock1_p & b26693 | !hlock1_p & b266db;
assign a5ea1b = hgrant2_p & a5f024 | !hgrant2_p & a5f026;
assign a5ea27 = hbusreq0_p & a5fccb | !hbusreq0_p & v84563c;
assign a5ef75 = hgrant2_p & a5ef70 | !hgrant2_p & a5ef74;
assign a5fad6 = hbusreq2 & a5fad3 | !hbusreq2 & a5fad5;
assign a5fbb3 = hbusreq0_p & v84563c | !hbusreq0_p & a5fb71;
assign cea47f = stateG10_1_p & deadba | !stateG10_1_p & cea3d8;
assign af34ba = hlock1_p & af3c4c | !hlock1_p & !af34b7;
assign a5eb38 = hbusreq0 & a5eb37 | !hbusreq0 & v84563c;
assign c3bcd8 = hbusreq3_p & c3bcb2 | !hbusreq3_p & !c3bcd7;
assign a5fcde = hready & a5fbab | !hready & a5fcdd;
assign a5eb36 = hbusreq0_p & a5fcef | !hbusreq0_p & v84563c;
assign a5f98d = hlock0_p & a5f98c | !hlock0_p & !a5fc2c;
assign c3bc3a = hbusreq3 & c3bc39 | !hbusreq3 & !c3bc36;
assign a5f58e = hlock0_p & a5f36e | !hlock0_p & a5f4ee;
assign ab0bca = hbusreq3 & dead53 | !hbusreq3 & v84564a;
assign deae67 = hlock1_p & deacdf | !hlock1_p & v845646;
assign a5fb26 = hready & v84563c | !hready & !c3bc02;
assign deadf5 = hlock3_p & deadcd | !hlock3_p & deadf4;
assign a5f06e = hbusreq2_p & a5f06d | !hbusreq2_p & a5f068;
assign b29e49 = hbusreq3 & v84563c | !hbusreq3 & b29c3c;
assign c3b716 = hlock0_p & c3b715 | !hlock0_p & !c3b6a8;
assign a5ebe8 = hmaster1_p & a5ebe7 | !hmaster1_p & a5eb3b;
assign a5fbd3 = hbusreq2 & a5fb7b | !hbusreq2 & a5fbc1;
assign cea88d = hbusreq2_p & cea889 | !hbusreq2_p & !cea887;
assign a5f862 = hlock1_p & a60177 | !hlock1_p & v84563c;
assign a5fd03 = hmaster1_p & v84563c | !hmaster1_p & a5fd02;
assign a60174 = stateG2_p & v84563c | !stateG2_p & !v8c6449;
assign ab0611 = hbusreq0_p & b29992 | !hbusreq0_p & ab0610;
assign cea23c = decide_p & cea23b | !decide_p & v84563c;
assign c3bc2d = hgrant2_p & c3bc29 | !hgrant2_p & c3bc2c;
assign ab0c0c = hbusreq2_p & ab0c0b | !hbusreq2_p & v84563c;
assign c3bd8c = locked_p & c3bd8b | !locked_p & c3bc47;
assign b29f58 = hlock0_p & b29f57 | !hlock0_p & v84563c;
assign cea47a = hlock1_p & deac51 | !hlock1_p & !cea479;
assign b29969 = hlock0_p & c3b6be | !hlock0_p & deadb2;
assign a5ea15 = hlock0_p & a5fa66 | !hlock0_p & a5e9c5;
assign ab0553 = hbusreq3 & ab0551 | !hbusreq3 & ab0552;
assign ab0b98 = hbusreq2_p & ab0b95 | !hbusreq2_p & ab0b97;
assign ab0be9 = decide_p & ab0be8 | !decide_p & v845662;
assign b299e8 = decide_p & b299e7 | !decide_p & b29e57;
assign ab0c65 = hmaster0_p & ab0c4a | !hmaster0_p & ab0c64;
assign a5f123 = hlock2_p & a5f109 | !hlock2_p & !a5f122;
assign a5fa41 = hlock0_p & a5fa37 | !hlock0_p & ab0c31;
assign b299d5 = decide_p & b299d4 | !decide_p & v84563c;
assign d40d45 = hbusreq2_p & d40d44 | !hbusreq2_p & d40d42;
assign a5f11c = hmastlock_p & v845654 | !hmastlock_p & v84563c;
assign a5f065 = locked_p & a5f6ec | !locked_p & a5fb6a;
assign a5e9d8 = hbusreq3 & a5e9d3 | !hbusreq3 & a5e9d7;
assign b29eb3 = stateA1_p & c07311 | !stateA1_p & !cea1ac;
assign a5fbea = hlock0_p & a5fbde | !hlock0_p & a5fbe9;
assign a5fc12 = hready & a5fbe1 | !hready & a5fbe5;
assign c3bd01 = hbusreq0_p & c3bcdb | !hbusreq0_p & !c3bcef;
assign a5f8b9 = hready & v84563c | !hready & deac52;
assign c3b7e4 = hlock0_p & c3bd5f | !hlock0_p & v84563c;
assign hmaster1 = b0c0ff;
assign b266e5 = hgrant2_p & b266e3 | !hgrant2_p & b266e4;
assign a5ee0e = hlock1_p & a5fb8b | !hlock1_p & ab05a1;
assign adaf10 = hready_p & adaefa | !hready_p & adaf0f;
assign deae01 = start_p & deac4a | !start_p & dead6c;
assign cea377 = hready & cea375 | !hready & cea376;
assign a5f072 = hlock0_p & a5f1e5 | !hlock0_p & a5f070;
assign ab06d6 = hmaster1_p & ab06d5 | !hmaster1_p & !ab0646;
assign af359e = hmaster0_p & af359b | !hmaster0_p & af359d;
assign deae51 = locked_p & deae50 | !locked_p & v84563c;
assign ab053f = hlock0_p & v84563c | !hlock0_p & !b2991b;
assign b29d70 = hlock0_p & b29d6f | !hlock0_p & !v84563c;
assign a5f2db = hbusreq3 & a5f2d8 | !hbusreq3 & a5f2da;
assign c3bcfd = hlock2_p & c3bce5 | !hlock2_p & v84563c;
assign ab05e8 = hbusreq2_p & ab052c | !hbusreq2_p & ab05e7;
assign c3bd90 = hlock2_p & c3bd8f | !hlock2_p & !c3bca0;
assign ab0b2f = hbusreq2_p & ab0b18 | !hbusreq2_p & ab0b16;
assign a5ea4b = hmaster1_p & a5ea38 | !hmaster1_p & a5ea4a;
assign d40d88 = hmaster1_p & d40d87 | !hmaster1_p & d40d60;
assign a5eade = hbusreq2_p & a5eadd | !hbusreq2_p & a5eadc;
assign a5f4cd = stateG10_1_p & v970407 | !stateG10_1_p & a5f4cc;
assign b29b0e = hbusreq3 & b29b0d | !hbusreq3 & b29a4b;
assign ab0b91 = hlock0_p & v84563c | !hlock0_p & !b29d8b;
assign c3bcc3 = hgrant0_p & c3bc5e | !hgrant0_p & c3bcc2;
assign b29e56 = hlock3_p & b29d9b | !hlock3_p & b29e55;
assign b29cfd = hready & deae1d | !hready & !v84563c;
assign c3bc8b = locked_p & v84563c | !locked_p & deacdf;
assign a5f231 = hlock0_p & a5f22f | !hlock0_p & a5f230;
assign dead70 = hlock1_p & deacf7 | !hlock1_p & !dead6f;
assign cea3f3 = hmaster1_p & cea3f2 | !hmaster1_p & !cea1a1;
assign a5f983 = hready & a5f982 | !hready & a5fbb0;
assign c3b635 = hready & c3b634 | !hready & !v84563c;
assign dead4f = decide_p & dead4e | !decide_p & v84563c;
assign ab06c7 = hmaster1_p & ab06c6 | !hmaster1_p & ab06a3;
assign ab051f = hmaster1_p & ab0518 | !hmaster1_p & ab051e;
assign c3bc61 = hlock1_p & v84563c | !hlock1_p & !c3bc60;
assign b299d0 = hbusreq2_p & b299cd | !hbusreq2_p & v84563c;
assign c3bdc5 = hlock0_p & c3bcee | !hlock0_p & c3bcf1;
assign a5ee7b = hgrant2_p & a5ee7a | !hgrant2_p & v84563c;
assign bdb5b3 = hbusreq2_p & bdb5b1 | !hbusreq2_p & bdb58b;
assign c3b8cb = jx0_p & c3b780 | !jx0_p & c3b8ca;
assign adaeef = hmaster0_p & v84563c | !hmaster0_p & adaeee;
assign d40d30 = start_p & v84563c | !start_p & d40d2f;
assign a5fb73 = hlock1_p & v84563c | !hlock1_p & a5fb72;
assign bdb5af = decide_p & v84565a | !decide_p & bdb59a;
assign b29a5c = hlock2_p & v84563c | !hlock2_p & !b29a5b;
assign v97040a = hgrant1_p & v970409 | !hgrant1_p & v9703fc;
assign cea38f = hlock0_p & cea389 | !hlock0_p & cea38e;
assign adaebc = hmastlock_p & adaebb | !hmastlock_p & v84563c;
assign ce9da5 = hlock3_p & ce9d79 | !hlock3_p & ce9d40;
assign a5ef6b = hbusreq0_p & a5f4f0 | !hbusreq0_p & a5edcc;
assign af3c2b = hbusreq2_p & af3c13 | !hbusreq2_p & v845646;
assign a5fd21 = hlock2 & a5fa2d | !hlock2 & ab0c32;
assign a5fa37 = hready & v84563c | !hready & ab0af9;
assign ab0cf3 = hmaster1_p & ab0be3 | !hmaster1_p & ab0cf2;
assign af34c1 = hlock2_p & af3c51 | !hlock2_p & af3c6b;
assign a5f7f5 = hmastlock_p & a5f7f4 | !hmastlock_p & v84563c;
assign cea15d = hgrant2_p & cea159 | !hgrant2_p & !cea15c;
assign v845652 = hburst0_p & v84563c | !hburst0_p & !v84563c;
assign b2670f = hlock0_p & b266a3 | !hlock0_p & !b266a2;
assign b29eb8 = hbusreq1_p & b29eb7 | !hbusreq1_p & !v84563c;
assign a60187 = hmastlock_p & a60186 | !hmastlock_p & v84563c;
assign b29a7d = hlock2_p & b29a7a | !hlock2_p & b29a7c;
assign a5fba8 = hlock1_p & a5fba2 | !hlock1_p & a5fba7;
assign c3bc42 = hmaster1_p & c3bc3b | !hmaster1_p & c3bc41;
assign ab0c5c = hready & ab0c5b | !hready & c3bd5d;
assign b26708 = decide_p & b26707 | !decide_p & b266c3;
assign a5f36b = hready & v84563c | !hready & a5f36a;
assign b29fe9 = decide_p & b29fe8 | !decide_p & b29e57;
assign a5ef9f = hbusreq2_p & a5ee19 | !hbusreq2_p & a5ef9e;
assign deaeb0 = hlock2_p & deaeaf | !hlock2_p & v84563c;
assign a5f3f8 = hready & a5f3f3 | !hready & a5f3f7;
assign b29cda = hgrant2_p & b29cd6 | !hgrant2_p & b29cd9;
assign c3bc9f = hgrant0_p & c3bc6b | !hgrant0_p & c3bc9e;
assign a5f24d = hready & a5f833 | !hready & a5f837;
assign c3b702 = hgrant2_p & c3b701 | !hgrant2_p & v845660;
assign dea764 = hmaster1_p & dea760 | !hmaster1_p & dea763;
assign a5f8ec = hbusreq2 & a5f8e7 | !hbusreq2 & !a5f8eb;
assign a5f9c7 = hbusreq2_p & a6019b | !hbusreq2_p & a6018d;
assign b29d79 = locked_p & b29d78 | !locked_p & !v84563c;
assign c3bd79 = hlock1_p & c3bbd2 | !hlock1_p & c3bd78;
assign a5ef10 = hbusreq1_p & a5fce3 | !hbusreq1_p & !v84563c;
assign a5f282 = hgrant2_p & v84563c | !hgrant2_p & a5f269;
assign a5fa2e = hlock0_p & a5fa2b | !hlock0_p & a5fa2d;
assign af34fb = hready_p & af34ed | !hready_p & af34fa;
assign b29d2f = hlock2_p & b29d2e | !hlock2_p & v84563c;
assign c3b6f2 = hmaster1_p & c3b6ee | !hmaster1_p & c3b6f1;
assign a5fc5f = hbusreq2 & a5fc5d | !hbusreq2 & a5fc5e;
assign b29e60 = hbusreq2_p & v84563c | !hbusreq2_p & !v845644;
assign ab0cd9 = hmaster1_p & ab0cd6 | !hmaster1_p & ab0cd8;
assign a5f906 = hready & v84563c | !hready & !cea0bc;
assign adaeff = hmastlock_p & adaefe | !hmastlock_p & v84563c;
assign a5f1be = hgrant2_p & a5fbc4 | !hgrant2_p & a5f1bd;
assign d40d78 = hmaster0_p & d40d77 | !hmaster0_p & d40d55;
assign deacd9 = hmaster0_p & deacb2 | !hmaster0_p & deacd8;
assign ab068c = hbusreq0_p & deacb7 | !hbusreq0_p & b29ef5;
assign b266a4 = hlock0_p & b2669d | !hlock0_p & b266a3;
assign a5fbf1 = locked_p & a5fbf0 | !locked_p & a5fbdd;
assign b266b1 = hbusreq0_p & b266a8 | !hbusreq0_p & b266ae;
assign ab0b21 = hlock0_p & c3bc03 | !hlock0_p & v84563c;
assign dea78b = hmaster0_p & dea78a | !hmaster0_p & !v84563c;
assign ce9e5f = jx0_p & ce9cdf | !jx0_p & ce9e5e;
assign c3b7db = hlock0_p & c3bd47 | !hlock0_p & !cea887;
assign a5f382 = hbusreq2_p & a5f381 | !hbusreq2_p & a5f380;
assign ab0b02 = hlock2_p & ab0b01 | !hlock2_p & v84563c;
assign c3b71c = hready & c3b71b | !hready & c3bdd4;
assign ab0573 = hlock2_p & ab0571 | !hlock2_p & !ab0572;
assign af356f = locked_p & v84563c | !locked_p & af352f;
assign a5f843 = hready & a5f836 | !hready & !a5f842;
assign b266b0 = hbusreq2_p & b266aa | !hbusreq2_p & b266af;
assign cea0d4 = hbusreq3 & cea0d3 | !hbusreq3 & cea877;
assign c3b7b0 = hlock0_p & c3bcdb | !hlock0_p & v84563c;
assign c3b771 = hgrant3_p & c3b74c | !hgrant3_p & !c3b770;
assign ab0cc6 = hlock2_p & ab0cc2 | !hlock2_p & ab0cc5;
assign a5fcc8 = locked_p & v845641 | !locked_p & a5fcc7;
assign b8acef = decide_p & b8ace0 | !decide_p & b8aced;
assign a5ea1e = hlock3_p & a5e9d0 | !hlock3_p & a5ea1d;
assign a5f38c = hbusreq1 & a5f38b | !hbusreq1 & v84563c;
assign af3504 = hgrant0_p & af3501 | !hgrant0_p & af3503;
assign a5fbdb = hready & a5fbd8 | !hready & a5fbda;
assign dea76a = hgrant2_p & dea765 | !hgrant2_p & dea769;
assign b2a011 = hbusreq2_p & b2a010 | !hbusreq2_p & v845644;
assign b2a01a = hready_p & b2a00d | !hready_p & !b2a019;
assign a5eb3e = hbusreq0_p & a5fcd9 | !hbusreq0_p & !v84563c;
assign af3584 = hbusreq2_p & af3583 | !hbusreq2_p & af3579;
assign v9703fb = start_p & v8e1935 | !start_p & !v9703fa;
assign cea26a = hburst0 & v84563c | !hburst0 & cea269;
assign cea494 = decide_p & cea493 | !decide_p & v84563c;
assign c3b811 = hlock2_p & c3b810 | !hlock2_p & !c3b7ab;
assign cea37e = hlock2_p & cea37d | !hlock2_p & cea37c;
assign b29989 = locked_p & b29988 | !locked_p & !v84563c;
assign dead8d = hlock2_p & dead8c | !hlock2_p & !v84563c;
assign a5fbcb = hlock2 & a5fb73 | !hlock2 & a5fbc6;
assign c3b615 = hlock2_p & c3b614 | !hlock2_p & !v84563c;
assign ab0734 = hmaster1_p & ab0685 | !hmaster1_p & ab0bca;
assign af349d = hlock0_p & af3c5e | !hlock0_p & af3c4c;
assign c3bcb3 = hbusreq2_p & v84564c | !hbusreq2_p & v845644;
assign a5ee0b = hmaster1_p & a5ee0a | !hmaster1_p & a60144;
assign ab066d = hlock2_p & ab066b | !hlock2_p & ab066c;
assign c3b72b = decide_p & c3b72a | !decide_p & v845660;
assign a5ef81 = hbusreq0_p & a5f4ee | !hbusreq0_p & a5edcc;
assign a5f588 = hbusreq0 & a5f586 | !hbusreq0 & !a5f587;
assign a5f1d9 = hbusreq2 & a5f1d5 | !hbusreq2 & a5f1d8;
assign a5f7a2 = hready & a5f9f6 | !hready & !deacb7;
assign c3bdb8 = hgrant2_p & dead3e | !hgrant2_p & c3bdb7;
assign v845647 = hbusreq1 & v84563c | !hbusreq1 & !v84563c;
assign a5f086 = hbusreq3 & a5f085 | !hbusreq3 & v84563c;
assign c3b646 = hmaster0_p & c3b630 | !hmaster0_p & c3b645;
assign ab0701 = hmaster0_p & ab06f7 | !hmaster0_p & ab0700;
assign b29fd2 = hready & deaca1 | !hready & !v84563c;
assign a81cc3 = hmaster1_p & a81cc1 | !hmaster1_p & a81cc2;
assign a5f946 = hready & v84563c | !hready & deacbe;
assign b2669a = hlock0_p & b26698 | !hlock0_p & b26699;
assign b29b21 = hlock0_p & c3bcf0 | !hlock0_p & v84563c;
assign b29fef = hmaster1_p & b29fee | !hmaster1_p & b29ed9;
assign b2a01b = hgrant3_p & b29ffb | !hgrant3_p & b2a01a;
assign deae0d = hlock0_p & deae0c | !hlock0_p & v84563c;
assign b29980 = hbusreq2_p & b2997f | !hbusreq2_p & b2997e;
assign a5f743 = hbusreq0_p & a5f6e9 | !hbusreq0_p & v84563c;
assign af3c5f = hlock0_p & af3c5d | !hlock0_p & af3c5e;
assign a5f20c = hbusreq2_p & a5f20b | !hbusreq2_p & v84563c;
assign ab0ba5 = hbusreq0_p & ab0ba3 | !hbusreq0_p & ab0ba4;
assign b298b2 = hbusreq3 & b298ad | !hbusreq3 & b298b1;
assign a5f028 = hgrant2_p & a5f025 | !hgrant2_p & a5f027;
assign af3c60 = hlock2_p & af3c5f | !hlock2_p & af3c5e;
assign adaee3 = hlock2_p & adaebd | !hlock2_p & v84563c;
assign c3bdad = hbusreq1_p & cea2e5 | !hbusreq1_p & deae02;
assign b840ad = hmaster1_p & v84564b | !hmaster1_p & v845643;
assign a5f1ad = hmastlock_p & a60196 | !hmastlock_p & v84563c;
assign a5fa69 = hlock2_p & a5fa68 | !hlock2_p & a5fa26;
assign ce9d13 = hmaster1_p & ce9d12 | !hmaster1_p & v84563c;
assign af34a5 = hbusreq2_p & af349e | !hbusreq2_p & af3c4c;
assign b26764 = hmaster0_p & b26760 | !hmaster0_p & !b26763;
assign b29f0d = hbusreq1_p & b29f0b | !hbusreq1_p & !v84565a;
assign dea7ad = hgrant3_p & dea7ac | !hgrant3_p & !v84563c;
assign c3b70d = hmaster1_p & c3b709 | !hmaster1_p & c3b70c;
assign b26719 = hlock2_p & b26717 | !hlock2_p & b26718;
assign c3b678 = hbusreq1_p & deadba | !hbusreq1_p & !c3b677;
assign a5fd08 = hbusreq2 & a5fcd9 | !hbusreq2 & a5fce5;
assign dead10 = hbusreq2_p & dead0f | !hbusreq2_p & dead0e;
assign ab0cc9 = hmaster1_p & ab0cc8 | !hmaster1_p & ab0c49;
assign cea1a1 = hgrant2_p & cea89e | !hgrant2_p & cea8a1;
assign a5ef61 = hbusreq2 & a5ef5f | !hbusreq2 & a5ef60;
assign a5f376 = hbusreq1 & a5f375 | !hbusreq1 & !v84563c;
assign a5f3c4 = hbusreq1 & a5f3c3 | !hbusreq1 & v84563c;
assign a5ef60 = hlock0_p & a5f540 | !hlock0_p & a5ef5e;
assign a5fa6e = hbusreq2 & a5fa6b | !hbusreq2 & a5fa6d;
assign ce9d11 = hbusreq2_p & cea236 | !hbusreq2_p & ce9d10;
assign a5f6e8 = locked_p & a5f6e7 | !locked_p & a5fb6a;
assign a5fbe9 = locked_p & a5fbe8 | !locked_p & a5fbdd;
assign a5f8ce = start_p & a5fba3 | !start_p & a6016d;
assign af3591 = decide_p & af3588 | !decide_p & af3590;
assign a5f24a = hlock0_p & a5f248 | !hlock0_p & !a5f249;
assign ab0aee = hlock1_p & ab0aeb | !hlock1_p & ab0aed;
assign a5eece = hbusreq2 & a5eebc | !hbusreq2 & a5eec4;
assign af3598 = hmaster1_p & af3572 | !hmaster1_p & af352d;
assign b29efe = hbusreq2_p & b29efd | !hbusreq2_p & b29cbb;
assign dea7aa = hmaster0_p & dea7a8 | !hmaster0_p & dea7a9;
assign af3572 = hbusreq2_p & v84563c | !hbusreq2_p & af3571;
assign b29a86 = hlock2 & b29cff | !hlock2 & b29a85;
assign a5efd3 = hlock2_p & a5f54b | !hlock2_p & a5f592;
assign a5ee1f = hlock1_p & a5fbab | !hlock1_p & !a5ee1e;
assign a5fa10 = hgrant1_p & a5fa0e | !hgrant1_p & a5fa0f;
assign adaeda = decide_p & adaed6 | !decide_p & adaed9;
assign c3bc68 = hbusreq2_p & c3bc67 | !hbusreq2_p & c3bc64;
assign a5f4a3 = stateG10_1_p & v84563c | !stateG10_1_p & a5f4a2;
assign c3bc0a = hlock0_p & c3bc09 | !hlock0_p & !c3bbd2;
assign a5fa59 = hlock1_p & a81cf0 | !hlock1_p & a5f9dd;
assign a81ce6 = hbusreq2_p & a81caa | !hbusreq2_p & a81cdc;
assign a5f71f = hlock0_p & a5fb7a | !hlock0_p & a5f71e;
assign a5f716 = hlock0_p & a5f713 | !hlock0_p & a5f715;
assign c3bcae = hgrant0_p & c3bca3 | !hgrant0_p & c3bcad;
assign c3b652 = hlock2_p & c3b651 | !hlock2_p & v845648;
assign ab0b35 = hbusreq3 & v84563c | !hbusreq3 & ab0ade;
assign af34f2 = hmaster0_p & d40d60 | !hmaster0_p & af34f1;
assign cea1b5 = locked_p & cea1b4 | !locked_p & b26697;
assign a5f71e = locked_p & v84563c | !locked_p & a5f71d;
assign a5f021 = hgrant2_p & a5f01e | !hgrant2_p & a5f020;
assign a5f343 = hbusreq2 & a5fcce | !hbusreq2 & v84563c;
assign b29a9f = hready_p & b29a58 | !hready_p & b29a9e;
assign a5f6dd = hgrant2_p & a5f6dc | !hgrant2_p & a5fae7;
assign a5f57f = hlock1_p & v84563c | !hlock1_p & b29929;
assign c3bde3 = hgrant3_p & c3bd82 | !hgrant3_p & c3bde2;
assign dead3a = hlock2_p & dead39 | !hlock2_p & v84563c;
assign ab0ca6 = hgrant0_p & ab0c91 | !hgrant0_p & !ab0ca5;
assign a5fa8b = hlock0_p & a5fa8a | !hlock0_p & v84563c;
assign cea3d0 = hbusreq2_p & cea3cf | !hbusreq2_p & cea3cd;
assign b29908 = hlock2_p & v84563c | !hlock2_p & !b29907;
assign a5ef2a = hbusreq2_p & a5ef28 | !hbusreq2_p & !a5ef29;
assign ab0b3c = hbusreq2_p & ab0b3a | !hbusreq2_p & ab0b3b;
assign cea252 = hbusreq1_p & cea250 | !hbusreq1_p & !v84563c;
assign ab0af1 = hlock2 & ab0ae6 | !hlock2 & ab0af0;
assign af3519 = hmaster1_p & af3518 | !hmaster1_p & !v84563c;
assign af3c21 = hbusreq2_p & af3c1d | !hbusreq2_p & v845646;
assign ce9cbd = hgrant0_p & ce9cb7 | !hgrant0_p & ce9cbc;
assign ce9d45 = hgrant2_p & cea15e | !hgrant2_p & !cea172;
assign a5f203 = hgrant2_p & v84563c | !hgrant2_p & a5f202;
assign c3b6e5 = hbusreq2_p & c3b6e4 | !hbusreq2_p & c3b6e2;
assign c3bc5d = hlock2_p & c3bc5c | !hlock2_p & dead2e;
assign c98ba4 = hgrant3_p & c98b9f | !hgrant3_p & c98ba3;
assign c3b7af = hmaster1_p & c3b7ac | !hmaster1_p & c3b7ae;
assign ab06a2 = hlock0_p & b29f3c | !hlock0_p & !deaca2;
assign a5f135 = hbusreq0 & a5f124 | !hbusreq0 & !ab0c31;
assign c3bc87 = hlock2_p & c3bc86 | !hlock2_p & !deace9;
assign b29a6e = hgrant2_p & b29ccb | !hgrant2_p & b29cd7;
assign deaea8 = hgrant2_p & deaea4 | !hgrant2_p & deaea7;
assign dea7b3 = jx1_p & dea7ae | !jx1_p & dea700;
assign af35bc = hmaster1_p & af3571 | !hmaster1_p & af359a;
assign a5f175 = hgrant1_p & a5f9f4 | !hgrant1_p & a5f174;
assign adaef4 = hmaster1_p & v84563c | !hmaster1_p & adaef3;
assign b29ae4 = hlock2_p & v84563c | !hlock2_p & !b29ae3;
assign ab0b54 = hbusreq2_p & ab0b53 | !hbusreq2_p & ab0b52;
assign b29d8a = hready & deacdf | !hready & v84563c;
assign a5ee2a = hlock1_p & a5fbb6 | !hlock1_p & a5ee1b;
assign a5fa71 = hgrant2_p & a5fa58 | !hgrant2_p & a5fa70;
assign c3b846 = hbusreq2_p & c3b845 | !hbusreq2_p & !c3b844;
assign a5f999 = hmaster1_p & a60144 | !hmaster1_p & a5f998;
assign dead79 = hbusreq2_p & dead78 | !hbusreq2_p & v845660;
assign dea744 = hbusreq3 & dea73d | !hbusreq3 & dea743;
assign d40d35 = hgrant1_p & d40d34 | !hgrant1_p & d40d31;
assign b29961 = hgrant2_p & b2995d | !hgrant2_p & b29960;
assign b29ab5 = hbusreq2_p & b29ab1 | !hbusreq2_p & b29ab4;
assign a9b9ee = hready_p & a9b9ed | !hready_p & v84563c;
assign cea2e3 = hburst1 & cea2e2 | !hburst1 & deae01;
assign cea337 = hbusreq2_p & cea336 | !hbusreq2_p & v84563c;
assign v8565cf = hbusreq3_p & v9269ad | !hbusreq3_p & v84563c;
assign c3b62a = locked_p & dead7d | !locked_p & deae59;
assign ab0b5b = hlock0_p & v845660 | !hlock0_p & b26695;
assign c3b698 = hready & c3b697 | !hready & v84563c;
assign be34e6 = hready_p & v84564a | !hready_p & be34e5;
assign a5e9d4 = hlock0_p & a5f906 | !hlock0_p & v84563c;
assign adaeea = hmastlock_p & adaee9 | !hmastlock_p & v84563c;
assign dead81 = hlock2_p & dead80 | !hlock2_p & !dead7f;
assign a5f73c = hlock2_p & a5f73b | !hlock2_p & v84563c;
assign cea476 = hlock3_p & cea45e | !hlock3_p & cea475;
assign c3b6fe = hmaster1_p & c3b6f7 | !hmaster1_p & c3b6fd;
assign cea1bf = locked_p & cea1be | !locked_p & v84563c;
assign cea18e = hbusreq0_p & v845660 | !hbusreq0_p & cea18d;
assign a5f7c4 = hlock2 & a5f7be | !hlock2 & a5f7c3;
assign ab06b7 = hbusreq0_p & deaca1 | !hbusreq0_p & b29f57;
assign a5f1b3 = hlock0_p & a5f1af | !hlock0_p & a5f1b2;
assign ab0d01 = hbusreq3_p & ab0cd1 | !hbusreq3_p & ab0d00;
assign b26736 = hlock0_p & b26735 | !hlock0_p & b266ae;
assign a5f8c1 = hlock2 & a5f8bb | !hlock2 & a5f8c0;
assign ab0cb2 = hmaster1_p & dead2e | !hmaster1_p & ab0cb1;
assign deadc6 = hlock2_p & deadc5 | !hlock2_p & !deadc4;
assign a5ea8f = hbusreq0_p & v845660 | !hbusreq0_p & v84563c;
assign af348f = hmaster1_p & af348d | !hmaster1_p & af348e;
assign c3b617 = hbusreq2_p & c3b615 | !hbusreq2_p & c3bcc5;
assign af357b = hlock0_p & af352d | !hlock0_p & af357a;
assign deadba = hmastlock_p & deadb9 | !hmastlock_p & v84563c;
assign a9b9ea = decide_p & a9b9e1 | !decide_p & a9b9e9;
assign cea166 = hgrant2_p & cea15e | !hgrant2_p & !cea165;
assign ab0512 = hlock2_p & ab0510 | !hlock2_p & ab0511;
assign af35c1 = hgrant3_p & af35a9 | !hgrant3_p & af35c0;
assign ce9cdc = hready_p & ce9cda | !hready_p & ce9cdb;
assign deae8b = hbusreq2_p & deae87 | !hbusreq2_p & deae86;
assign dea76c = hmaster0_p & dea764 | !hmaster0_p & dea76b;
assign b29aaa = hbusreq2_p & b29aa9 | !hbusreq2_p & v84563c;
assign a5f954 = hbusreq2 & a5fcdf | !hbusreq2 & !v84563c;
assign ab05fa = hlock0_p & deada8 | !hlock0_p & !ab05f9;
assign a5f034 = hlock3_p & a5f6ce | !hlock3_p & v84563c;
assign ab067f = hlock0_p & c3bcf8 | !hlock0_p & !v84563c;
assign deac9e = hmaster1_p & deac7e | !hmaster1_p & deac9d;
assign a5ef0b = locked_p & a5ef0a | !locked_p & !a5edfa;
assign a5ea85 = hlock2_p & a5ea84 | !hlock2_p & a5ea5e;
assign b29e9f = hmaster1_p & b29e9e | !hmaster1_p & !b29e6e;
assign a5fc21 = hlock1_p & v84563c | !hlock1_p & a5fb71;
assign b26750 = hgrant2_p & b2674f | !hgrant2_p & b266b3;
assign b29a59 = hgrant1_p & cea8a8 | !hgrant1_p & deadde;
assign b266fb = hlock0_p & b266ca | !hlock0_p & b266bb;
assign ab0d04 = hlock0_p & v84563c | !hlock0_p & !b29826;
assign a5ee06 = hlock0_p & a5f385 | !hlock0_p & a5f36b;
assign a5ec24 = hgrant3_p & a5ec22 | !hgrant3_p & a5ec23;
assign c3bbbc = hlock0_p & c3bbbb | !hlock0_p & v845660;
assign a5e9c4 = hready & a5e9c1 | !hready & a5e9c3;
assign a5ede5 = hlock3_p & a5f58b | !hlock3_p & a5ede4;
assign ab06e2 = hlock2_p & ab06e0 | !hlock2_p & ab06e1;
assign a5ea11 = hready & a5f9dd | !hready & c3bbd2;
assign dea728 = hbusreq3 & dea727 | !hbusreq3 & deae55;
assign cea31b = hmaster1_p & v84563c | !hmaster1_p & cea31a;
assign b29a22 = jx1_p & b299eb | !jx1_p & b29a21;
assign a5f246 = hgrant1_p & a5f7f5 | !hgrant1_p & a5f7f7;
assign a81cdb = hmastlock_p & a81cda | !hmastlock_p & v84563c;
assign a5fb4d = hlock0_p & a5fb4c | !hlock0_p & v84563c;
assign a5f324 = hbusreq2 & a5f321 | !hbusreq2 & a5f323;
assign c3b870 = hlock3_p & c3b85b | !hlock3_p & !c3b7ff;
assign ab0609 = hmaster1_p & ab058e | !hmaster1_p & ab0608;
assign c3b63c = hlock2_p & c3b63b | !hlock2_p & c3b63a;
assign ab0cbe = hlock0_p & v84563c | !hlock0_p & !ab0cbd;
assign dea6de = locked_p & deae59 | !locked_p & !deae67;
assign a5ee8c = hready & a5ee8b | !hready & a5ee2e;
assign a5e9c6 = hlock0_p & a5e9c4 | !hlock0_p & !a5e9c5;
assign b29a52 = hlock2_p & v84563c | !hlock2_p & !b29d92;
assign b29cd6 = hbusreq3 & b29ccb | !hbusreq3 & b29cd5;
assign c3b877 = hmaster0_p & c3b875 | !hmaster0_p & c3b876;
assign a5f4ca = hlock1_p & a6016f | !hlock1_p & !a5f4c9;
assign a5f921 = hlock1_p & deac52 | !hlock1_p & deacbd;
assign af3c19 = hlock2_p & b8acdc | !hlock2_p & v845646;
assign dead0b = locked_p & dead08 | !locked_p & !dead0a;
assign a5f6d7 = hbusreq3 & a5f6d5 | !hbusreq3 & a5f6d6;
assign a5fc3f = hgrant2_p & a5fc3b | !hgrant2_p & a5fc3e;
assign b29f83 = hlock3_p & b29f5f | !hlock3_p & b29f82;
assign a5fc40 = hmaster1_p & a5fc26 | !hmaster1_p & a5fc3f;
assign dead39 = hlock0_p & v845660 | !hlock0_p & v84563c;
assign c3bc53 = hlock0_p & c3bc52 | !hlock0_p & !v84563c;
assign c3bc5c = hlock0_p & c3bbbb | !hlock0_p & !v84563c;
assign ab069f = hbusreq3 & ab069d | !hbusreq3 & ab069e;
assign deadeb = hbusreq1_p & v84563c | !hbusreq1_p & !deadde;
assign b266ed = hbusreq2_p & b266e7 | !hbusreq2_p & !b266a0;
assign a5f1f3 = hready & a5f1f0 | !hready & a5f1f2;
assign ab0575 = hbusreq2_p & ab0573 | !hbusreq2_p & ab0571;
assign af34e5 = hmaster0_p & af34e3 | !hmaster0_p & af34e4;
assign a5f54c = hbusreq2 & a5f54a | !hbusreq2 & a5f54b;
assign a5f215 = hgrant2_p & v84563c | !hgrant2_p & a5f214;
assign a5f39d = hmaster0_p & a5f384 | !hmaster0_p & a5f39c;
assign a5f47c = hmaster1_p & a5f47b | !hmaster1_p & a5f6d9;
assign a5efec = hmaster1_p & a5efe2 | !hmaster1_p & a5efeb;
assign deae42 = hgrant2_p & deae40 | !hgrant2_p & deae41;
assign ab0bbb = hgrant2_p & ab0bba | !hgrant2_p & cea15a;
assign a5eba1 = hmaster0_p & a5eba0 | !hmaster0_p & a5eaa1;
assign b29aa9 = hlock2_p & v84563c | !hlock2_p & !b29aa8;
assign bdb5a4 = hmaster0_p & bdb598 | !hmaster0_p & bdb5a3;
assign cea399 = hmaster1_p & cea392 | !hmaster1_p & cea398;
assign dea6ec = hmaster0_p & dea6eb | !hmaster0_p & deaea9;
assign b2994f = hlock0_p & b2994e | !hlock0_p & !b29cfe;
assign cea86f = hbusreq3 & cea86e | !hbusreq3 & v84563c;
assign b2675d = hlock1_p & b26693 | !hlock1_p & b2675c;
assign ab0c9e = hlock2_p & ab0c95 | !hlock2_p & ab0c9d;
assign a5fa64 = hlock1_p & a60177 | !hlock1_p & !a5fa63;
assign adaf05 = hbusreq1_p & adaec4 | !hbusreq1_p & adaeff;
assign c3b8af = hgrant2_p & c3b8ac | !hgrant2_p & c3b8ae;
assign b29fae = hlock0_p & b29ec6 | !hlock0_p & c3bce5;
assign adaf03 = hmaster1_p & v84563c | !hmaster1_p & adaf02;
assign adaed6 = hlock3_p & adaed3 | !hlock3_p & adaed5;
assign a5f2c9 = hbusreq2_p & a5f2c8 | !hbusreq2_p & v84563c;
assign a5f1ca = hlock0_p & a5f1c9 | !hlock0_p & v84563c;
assign a5fcd6 = start_p & cea1aa | !start_p & !b29f17;
assign a5eaee = hbusreq2_p & a5ead6 | !hbusreq2_p & a5ead2;
assign c3b6c0 = hlock0_p & c3b6bf | !hlock0_p & c3b66b;
assign a5fcbc = hlock0_p & c3bcf8 | !hlock0_p & a5fcbb;
assign cea489 = hbusreq3 & cea487 | !hbusreq3 & cea488;
assign a5ea34 = hbusreq2 & a5f09b | !hbusreq2 & v845641;
assign deac86 = hbusreq0_p & deac52 | !hbusreq0_p & v84565a;
assign a5fb23 = hbusreq2_p & a5fb22 | !hbusreq2_p & v84563c;
assign a5f18d = hready & a5f189 | !hready & a5f18c;
assign a5f4a7 = hbusreq1 & a60173 | !hbusreq1 & v84563c;
assign a5fd26 = hbusreq2 & a5fd25 | !hbusreq2 & !v84563c;
assign a5fb85 = hbusreq3 & a5fb84 | !hbusreq3 & a60144;
assign c3bcc8 = hlock2_p & c3bc0d | !hlock2_p & !v84563c;
assign a5eaa1 = hmaster1_p & a5eaa0 | !hmaster1_p & v84563c;
assign a81cf5 = hmaster0_p & v84563c | !hmaster0_p & a81cf4;
assign c3bcc1 = hmaster1_p & c3bc71 | !hmaster1_p & c3bcc0;
assign ce9d58 = hmaster0_p & ce9d56 | !hmaster0_p & ce9d57;
assign cea2b6 = decide_p & cea2b5 | !decide_p & v84563c;
assign b29b24 = hgrant2_p & b29b20 | !hgrant2_p & !b29b23;
assign a5fb32 = hready & a60186 | !hready & v9703fb;
assign c3b753 = hgrant2_p & c3b752 | !hgrant2_p & c3bc70;
assign a5f97b = hbusreq2_p & a5f97a | !hbusreq2_p & a60142;
assign cea364 = decide_p & cea363 | !decide_p & a57859;
assign a5f43d = hlock1_p & a60177 | !hlock1_p & !a5f43c;
assign dea785 = hbusreq3 & dea782 | !hbusreq3 & dea784;
assign deace6 = hbusreq2_p & deace5 | !hbusreq2_p & deace2;
assign ab061c = hgrant2_p & ab061b | !hgrant2_p & cea15a;
assign a5fc1c = locked_p & v84563c | !locked_p & a5fc1a;
assign v970408 = hmastlock_p & v970407 | !hmastlock_p & v84563c;
assign af3c51 = hlock0_p & af3c4f | !hlock0_p & af3c50;
assign cea46f = hgrant2_p & cea46e | !hgrant2_p & !v845660;
assign a5f525 = hready & a5f520 | !hready & a5f493;
assign ab074c = hgrant0_p & ab0be1 | !hgrant0_p & !ab074b;
assign af3c58 = locked_p & af3c55 | !locked_p & af3c4c;
assign a5fc51 = hmastlock_p & a5fc50 | !hmastlock_p & v84563c;
assign a5f2f9 = hbusreq2_p & a5f2f8 | !hbusreq2_p & v84563c;
assign ab0581 = hbusreq2_p & ab057f | !hbusreq2_p & ab057e;
assign b2999d = locked_p & b2999c | !locked_p & !v84563c;
assign b2678a = hmaster0_p & b26789 | !hmaster0_p & !b26700;
assign a5ea66 = hlock2_p & a5ea65 | !hlock2_p & v845641;
assign b29fd9 = hready & b29fd8 | !hready & v84563c;
assign af35a3 = hmaster1_p & af3579 | !hmaster1_p & af352f;
assign a5f4e4 = hbusreq1 & a5f4e3 | !hbusreq1 & v84563c;
assign cea1bd = hlock1_p & v84563c | !hlock1_p & cea1bc;
assign a5e9ce = hgrant2_p & a5fae2 | !hgrant2_p & a5fae7;
assign dead40 = hlock1_p & dead33 | !hlock1_p & v84563c;
assign a5ee9d = hlock0_p & a5ee9c | !hlock0_p & a5ee49;
assign ab0737 = hbusreq0_p & deaca2 | !hbusreq0_p & !deacaa;
assign a5f9a6 = locked_p & v84563c | !locked_p & a5f9a5;
assign a5f194 = hbusreq2 & a5f17e | !hbusreq2 & !a5f193;
assign a81cca = hmaster0_p & a81cc9 | !hmaster0_p & v84563c;
assign a5ea2b = hbusreq2_p & a5ea29 | !hbusreq2_p & a5ea2a;
assign v97043d = start_p & b2669e | !start_p & v84563c;
assign b266ba = hbusreq2_p & b26695 | !hbusreq2_p & !b266a0;
assign a5eeaf = hlock2_p & a5eeae | !hlock2_p & a5ee78;
assign a5f6d0 = hlock2_p & a5fa6b | !hlock2_p & v84563c;
assign ab05d1 = hbusreq2_p & ab05d0 | !hbusreq2_p & ab05b5;
assign cea878 = hbusreq3 & cea877 | !hbusreq3 & v84563c;
assign a5f754 = hbusreq2_p & a5f753 | !hbusreq2_p & v84563c;
assign ab0679 = hlock0_p & c3bcf8 | !hlock0_p & v845660;
assign c3bca6 = hgrant2_p & dead3e | !hgrant2_p & !c3bca5;
assign a5edc7 = hbusreq1 & a5edc6 | !hbusreq1 & c3b6a0;
assign a5ee6b = hgrant2_p & a5ee6a | !hgrant2_p & v84563c;
assign ab06a7 = hgrant2_p & ab06a5 | !hgrant2_p & ab06a6;
assign cea3c0 = hready & cea3bb | !hready & cea3bf;
assign b29832 = hready & v8c6711 | !hready & v84563c;
assign c3bd6b = hlock2_p & c3bd60 | !hlock2_p & v84563c;
assign deadcf = hgrant1_p & v84563c | !hgrant1_p & deadce;
assign b29836 = hbusreq2_p & b29835 | !hbusreq2_p & v84563c;
assign a81cb1 = hmastlock_p & a81cb0 | !hmastlock_p & v84563c;
assign deadd9 = hbusreq2_p & deadd2 | !hbusreq2_p & v84563c;
assign b29cbe = hbusreq3 & b29cbd | !hbusreq3 & v84563c;
assign a5f784 = hbusreq1_p & deac52 | !hbusreq1_p & a60172;
assign ce9cc5 = hbusreq3 & ce9cc2 | !hbusreq3 & ce9cc4;
assign v97042b = hmaster0_p & v970416 | !hmaster0_p & v97042a;
assign b29995 = hlock2 & b29991 | !hlock2 & b29994;
assign af34fd = decide_p & af3c6d | !decide_p & af3c72;
assign c3bc65 = locked_p & dead6e | !locked_p & b26695;
assign a5f3d4 = hbusreq1 & a5f3d3 | !hbusreq1 & !v84563c;
assign a5eb9e = hbusreq0 & a5f0ac | !hbusreq0 & v84563c;
assign cea3f1 = hbusreq3 & cea3ef | !hbusreq3 & cea3f0;
assign dea747 = hbusreq3 & dea745 | !hbusreq3 & dea746;
assign dead7f = locked_p & dead7b | !locked_p & v84563c;
assign a5f59a = hmaster1_p & a5f599 | !hmaster1_p & v84563c;
assign a5fcd9 = locked_p & a5fcd8 | !locked_p & !v84565a;
assign ab073c = hmaster1_p & ab06d5 | !hmaster1_p & !ab0bdb;
assign b2993b = hlock0_p & b2993a | !hlock0_p & !b29cdf;
assign a5ee22 = hready & a5ee1d | !hready & a5ee21;
assign a5fcf1 = hbusreq3 & a5fcf0 | !hbusreq3 & v84563c;
assign a5edd9 = hbusreq1 & a5f57e | !hbusreq1 & a5edd8;
assign b29955 = hgrant2_p & b2994c | !hgrant2_p & b29954;
assign b29ea4 = hbusreq3_p & b29e5b | !hbusreq3_p & b29ea3;
assign ab0c6d = hlock2_p & ab0af6 | !hlock2_p & v84563c;
assign b29cc0 = hbusreq3 & b29cbf | !hbusreq3 & v84563c;
assign a5f025 = hbusreq0 & a5f024 | !hbusreq0 & v845644;
assign c3bd45 = hbusreq3 & c3bd44 | !hbusreq3 & c3bd42;
assign cea171 = hgrant2_p & cea169 | !hgrant2_p & !cea170;
assign b29a93 = hbusreq3 & b29a91 | !hbusreq3 & b29a92;
assign ab0c8c = hlock0_p & ab0c8b | !hlock0_p & ab0c89;
assign deacae = hbusreq3 & deaca2 | !hbusreq3 & !deacad;
assign c3b823 = hmaster1_p & c3b81c | !hmaster1_p & c3b822;
assign b2672a = locked_p & b26728 | !locked_p & !b26729;
assign a5fb64 = hgrant2_p & a5fb61 | !hgrant2_p & a5fb63;
assign cea2f7 = hmaster1_p & cea15d | !hmaster1_p & cea2f0;
assign ab06cd = hlock2 & ab06cb | !hlock2 & ab06cc;
assign b29f64 = hbusreq3 & b29f61 | !hbusreq3 & b29f63;
assign deacec = hlock1_p & v84563c | !hlock1_p & deaceb;
assign a5f364 = hbusreq1_p & a5fb8a | !hbusreq1_p & v84563c;
assign af3c1d = hlock2_p & af3c1c | !hlock2_p & v845646;
assign b2995e = hbusreq2_p & b29959 | !hbusreq2_p & v84563c;
assign a5f886 = hbusreq2_p & a5f884 | !hbusreq2_p & a5f9c3;
assign ce9cb3 = hready_p & cea494 | !hready_p & cea4af;
assign a5eddd = hbusreq2_p & a5eddc | !hbusreq2_p & a5f582;
assign b29eda = hmaster1_p & b29ed6 | !hmaster1_p & b29ed9;
assign b29f66 = hbusreq2_p & b29f62 | !hbusreq2_p & v84563c;
assign deae3b = hbusreq3 & deae3a | !hbusreq3 & !v84563c;
assign c3bcf2 = hlock0_p & c3bc48 | !hlock0_p & c3bcf1;
assign c3b60a = hgrant0_p & c3bdfe | !hgrant0_p & c3be06;
assign c3b74c = hready_p & c3b73e | !hready_p & c3b74b;
assign b29d35 = hlock2_p & b29d33 | !hlock2_p & b29d34;
assign b266b7 = hmaster0_p & b266a7 | !hmaster0_p & !b266b6;
assign ab0588 = hlock0_p & ab0b5e | !hlock0_p & cea37b;
assign ab050c = hlock2_p & ab0d07 | !hlock2_p & ab050b;
assign a5f722 = hbusreq2_p & a5f721 | !hbusreq2_p & a60142;
assign cea2af = hlock0_p & cea2ae | !hlock0_p & cea887;
assign b29fa9 = hmaster0_p & b29fa6 | !hmaster0_p & b29fa8;
assign a5ee84 = hlock0_p & a5ee83 | !hlock0_p & a5f38f;
assign a5eb76 = hmaster1_p & a5eb75 | !hmaster1_p & a5e9ea;
assign a5ea95 = hbusreq0 & a5ea94 | !hbusreq0 & v84563c;
assign b26759 = hlock0_p & b26699 | !hlock0_p & b26758;
assign a5ea60 = hlock0_p & a5f728 | !hlock0_p & v84563c;
assign a5ec20 = hlock3_p & a5ec19 | !hlock3_p & a5ec1f;
assign a5fa6a = hbusreq2_p & a5fa69 | !hbusreq2_p & v84563c;
assign af3c35 = hgrant2_p & v845646 | !hgrant2_p & af3c2d;
assign c3b6bd = hlock1_p & c3bbd2 | !hlock1_p & c3b6bc;
assign a5ee94 = hlock0_p & a5f387 | !hlock0_p & a5ee39;
assign ab0758 = hgrant2_p & ab06a5 | !hgrant2_p & ab0757;
assign dea72b = hmaster1_p & v845660 | !hmaster1_p & deac0f;
assign a5f713 = hready & a5f710 | !hready & a5f712;
assign a5fb12 = hlock1_p & a60167 | !hlock1_p & a5fb11;
assign b29d7d = hready & b29d77 | !hready & cea151;
assign b29d2c = hmaster1_p & v84563c | !hmaster1_p & b29d2b;
assign af3c6e = hlock3_p & af3c68 | !hlock3_p & af3c6d;
assign b29824 = hlock1_p & dead6e | !hlock1_p & b29823;
assign c3b73b = hbusreq3 & c3b656 | !hbusreq3 & !c3b73a;
assign c3b79f = hbusreq3 & c3b79a | !hbusreq3 & c3b79e;
assign ab0524 = hlock2_p & ab0522 | !hlock2_p & ab0523;
assign c3bd12 = stateG10_1_p & cea249 | !stateG10_1_p & c3bd11;
assign a5ebcb = hmaster1_p & a5e9cd | !hmaster1_p & a5f6dd;
assign cea25a = hlock2_p & cea259 | !hlock2_p & v84563c;
assign dead2a = hmaster0_p & dead13 | !hmaster0_p & dead29;
assign a5f28f = hready & v84563c | !hready & !deacdf;
assign dead32 = start_p & v845652 | !start_p & !dead31;
assign b29a4e = hlock2_p & v84563c | !hlock2_p & !b29a4d;
assign a5f879 = hready & v84563c | !hready & deac5b;
assign a5f0e6 = hlock0_p & a5f7b4 | !hlock0_p & a5f0e5;
assign b26717 = hlock0_p & b26698 | !hlock0_p & b26716;
assign a5eec6 = hlock0_p & a5f3cf | !hlock0_p & a5eec5;
assign cea390 = hbusreq2_p & cea38c | !hbusreq2_p & cea38f;
assign a6018b = hbusreq1 & v84563c | !hbusreq1 & a6018a;
assign a5f797 = hlock1_p & a60172 | !hlock1_p & a5f796;
assign deae9b = hbusreq3 & deae99 | !hbusreq3 & deae9a;
assign a9b9e8 = hmaster0_p & a9b9e5 | !hmaster0_p & !a9b9e7;
assign a5f545 = hlock0_p & a5f36e | !hlock0_p & a5f544;
assign b29f41 = hlock0_p & deaca2 | !hlock0_p & b29f40;
assign b29d68 = hlock2 & b29d65 | !hlock2 & b29d67;
assign b29f06 = hmastlock_p & b29f05 | !hmastlock_p & v84563c;
assign b29a78 = hready & b29a77 | !hready & c3bd16;
assign deae17 = hmaster1_p & dead3c | !hmaster1_p & deae10;
assign b29f76 = hbusreq1_p & b29ee9 | !hbusreq1_p & deac52;
assign a5f95c = hmaster1_p & v84563c | !hmaster1_p & a5f95b;
assign a5efcf = hready & v84563c | !hready & b8acdb;
assign cea40a = hlock1_p & v84563c | !hlock1_p & !cea408;
assign a5fc7d = hmastlock_p & a5fc7c | !hmastlock_p & !v84563c;
assign ab0bea = hlock2_p & ab0b0e | !hlock2_p & v84563c;
assign a5fbb5 = start_p & v845654 | !start_p & !a5fba4;
assign c3b7ec = hgrant2_p & c3b7e7 | !hgrant2_p & c3b7eb;
assign c3b68f = hgrant2_p & c3b68b | !hgrant2_p & c3b68e;
assign c3b622 = hlock1_p & v84563c | !hlock1_p & !deae4d;
assign a5f2f2 = locked_p & v84563c | !locked_p & a5f2f1;
assign a5eec8 = hmaster1_p & a5f3d9 | !hmaster1_p & a5eec7;
assign a5f6d5 = hbusreq2_p & a5f6d0 | !hbusreq2_p & a5fa6b;
assign cea156 = hbusreq3 & cea155 | !hbusreq3 & cea85f;
assign b29f82 = hmaster0_p & b29f6d | !hmaster0_p & !b29f81;
assign ab05a1 = hbusreq1_p & v84563c | !hbusreq1_p & !dead33;
assign a5f92e = hready & a60168 | !hready & deac52;
assign a5efa2 = hbusreq2_p & a5ee32 | !hbusreq2_p & a5efa1;
assign dead64 = hbusreq2_p & deacd2 | !hbusreq2_p & deacbf;
assign af34b3 = hlock2_p & af3c59 | !hlock2_p & af3c4c;
assign b29e67 = hready & deacbe | !hready & !cea29f;
assign c3b8b0 = hlock0_p & c3bd47 | !hlock0_p & !ce9dc7;
assign a9b9e5 = hmaster1_p & v84563c | !hmaster1_p & a9b9e4;
assign b29a49 = hbusreq2_p & b29a48 | !hbusreq2_p & v84563c;
assign deae5f = locked_p & deae59 | !locked_p & !v84563c;
assign ab0ce0 = hmaster1_p & ab0cdf | !hmaster1_p & ab0c47;
assign d40d50 = hlock1_p & v84563c | !hlock1_p & d40d4f;
assign a5ea41 = hlock0_p & a5f9a1 | !hlock0_p & a5ea40;
assign ab0619 = hlock0_p & v84563c | !hlock0_p & !ab0618;
assign cea149 = hlock2_p & cea148 | !hlock2_p & v84563c;
assign c3b6f6 = hlock0_p & c3b636 | !hlock0_p & c3b635;
assign c3bc34 = hbusreq2_p & c3bc33 | !hbusreq2_p & v84563c;
assign b29a48 = hlock2_p & v84563c | !hlock2_p & !b29d81;
assign ab0513 = hlock0_p & b298a4 | !hlock0_p & b299d7;
assign b29a83 = hlock1_p & v84565a | !hlock1_p & !b29a82;
assign jx2 = !b8acf4;
assign c3be05 = hmaster1_p & c3be04 | !hmaster1_p & c3bd9f;
assign c3b737 = hbusreq3 & c3b650 | !hbusreq3 & !c3b736;
assign a5fafc = hbusreq1 & a60169 | !hbusreq1 & a5fafb;
assign ab0743 = hbusreq2_p & ab0742 | !hbusreq2_p & ab06eb;
assign v970456 = hmaster0_p & v970455 | !hmaster0_p & v84563c;
assign a5ea99 = hmaster1_p & a5ea93 | !hmaster1_p & a5ea98;
assign ab0baf = hlock2_p & ab0bae | !hlock2_p & v84563c;
assign a5eb52 = hmaster1_p & a5eb51 | !hmaster1_p & !a5f0a9;
assign a5fc78 = hmastlock_p & a5fc77 | !hmastlock_p & v84563c;
assign deadc3 = hgrant1_p & deadbb | !hgrant1_p & deadba;
assign c3bc04 = hlock0_p & c3bc03 | !hlock0_p & v84565a;
assign cea383 = locked_p & cea382 | !locked_p & !cea380;
assign ab0caa = hready & deae02 | !hready & !dead6e;
assign a5ee36 = hmaster0_p & a5ee0b | !hmaster0_p & a5ee35;
assign ab0afb = hlock0_p & ab0afa | !hlock0_p & v84565a;
assign a5fc4c = hbusreq3 & a5fc4b | !hbusreq3 & v84563c;
assign deacc0 = hbusreq3 & deacb8 | !hbusreq3 & !deacbf;
assign ab0b4d = hmaster1_p & ab0b40 | !hmaster1_p & ab0b4c;
assign deae99 = hbusreq2_p & deae92 | !hbusreq2_p & deae91;
assign a5f298 = hbusreq2 & a5fc7f | !hbusreq2 & !v84563c;
assign dea72e = hbusreq2_p & dead8f | !hbusreq2_p & dead2e;
assign b29fb1 = hmaster1_p & b29fad | !hmaster1_p & b29fb0;
assign a5f857 = hbusreq2_p & a5f856 | !hbusreq2_p & !v84563c;
assign a5fc2d = hlock0_p & v845641 | !hlock0_p & a5fc2c;
assign b29f1a = stateG10_1_p & v84565a | !stateG10_1_p & b29f19;
assign a5e9fd = hlock0_p & a5fa21 | !hlock0_p & a5f192;
assign dead43 = hgrant2_p & dead3f | !hgrant2_p & !dead42;
assign ab0595 = hbusreq2_p & ab0594 | !hbusreq2_p & ab0592;
assign ce9ccf = hbusreq3_p & cea490 | !hbusreq3_p & ce9cce;
assign a5efc5 = hmaster0_p & a5efb5 | !hmaster0_p & a5efc4;
assign dea760 = hgrant2_p & dea75e | !hgrant2_p & dea75f;
assign a5f474 = hbusreq2 & a5f45b | !hbusreq2 & a5f473;
assign b29aa2 = hgrant2_p & b29aa1 | !hgrant2_p & !b29d5a;
assign a5ee32 = hlock2_p & a5ee29 | !hlock2_p & !a5ee31;
assign a5ec1f = hmaster0_p & v84563c | !hmaster0_p & a5ec1e;
assign a5ef7a = hbusreq2_p & a5edbb | !hbusreq2_p & a5ef79;
assign dea6db = decide_p & dea6da | !decide_p & !v84563c;
assign b29d4b = hgrant2_p & b29d49 | !hgrant2_p & b29d4a;
assign ce9d48 = hlock2_p & ce9d46 | !hlock2_p & !ce9d47;
assign c3bd62 = hlock0_p & c3bd5e | !hlock0_p & !c3bd61;
assign c3b81e = hbusreq2_p & c3b81d | !hbusreq2_p & !c3b7ad;
assign cea3a4 = hbusreq2_p & cea37b | !hbusreq2_p & !cea38d;
assign a60143 = hlock2_p & a60142 | !hlock2_p & v84563c;
assign ab06d3 = hlock2_p & ab06d2 | !hlock2_p & b29a7b;
assign a5eebd = hbusreq0_p & a5f3c9 | !hbusreq0_p & !a5eebc;
assign cea3ce = hlock0_p & cea3c0 | !hlock0_p & cea3cd;
assign ab0716 = hlock0_p & b29fda | !hlock0_p & !b29fdc;
assign b298ab = hlock0_p & b298aa | !hlock0_p & !v84563c;
assign ab0547 = hbusreq1_p & v84563c | !hbusreq1_p & !ab0546;
assign a5f94c = hbusreq2_p & a5f93c | !hbusreq2_p & a5fd35;
assign cea0b9 = hlock2_p & cea0b8 | !hlock2_p & v84563c;
assign bdb581 = hmaster0_p & bdb580 | !hmaster0_p & !v84563c;
assign cea196 = hready & c98b95 | !hready & !v84563c;
assign a5efa6 = hlock0_p & a60140 | !hlock0_p & a5f38f;
assign b298a0 = locked_p & v84563c | !locked_p & !cea37b;
assign af3c44 = decide_p & af3c3c | !decide_p & v8567b4;
assign a5f3c2 = hlock3_p & a5f39d | !hlock3_p & a5f3c1;
assign b299ec = hmaster1_p & b29cc1 | !hmaster1_p & b29e65;
assign a5f177 = hready & a5f176 | !hready & a5f797;
assign bdb588 = hbusreq2_p & bdb586 | !hbusreq2_p & bdb585;
assign a5ea82 = locked_p & a5ea81 | !locked_p & !v845641;
assign a5f479 = hbusreq2_p & a5f475 | !hbusreq2_p & a5f45c;
assign cea405 = hready & cea404 | !hready & deae59;
assign dead99 = hlock0_p & dead8a | !hlock0_p & !v84563c;
assign a5fc1e = hbusreq2 & a5fc1b | !hbusreq2 & a5fc1d;
assign a5fb67 = hlock3_p & a5faeb | !hlock3_p & a5fb66;
assign ab05dc = hlock0_p & v84563c | !hlock0_p & !ab05db;
assign deae04 = hlock1_p & deae02 | !hlock1_p & deae03;
assign a5edbc = hbusreq2_p & a5edbb | !hbusreq2_p & a5f510;
assign c3bdd9 = hbusreq2_p & c3bdd8 | !hbusreq2_p & v84563c;
assign cea8ae = hbusreq2_p & cea8ad | !hbusreq2_p & v84563c;
assign b29f51 = hready & b29f50 | !hready & v84563c;
assign a5ee56 = hlock1_p & a5fbab | !hlock1_p & !a5ee55;
assign d40d8c = hready_p & d40d76 | !hready_p & d40d8b;
assign a5fc00 = hbusreq1_p & v84563c | !hbusreq1_p & a5fb8b;
assign cea38a = locked_p & v84563c | !locked_p & cea37b;
assign a5f1e2 = locked_p & a5f1e1 | !locked_p & !v845641;
assign b266d3 = hlock2_p & b266d2 | !hlock2_p & b266ca;
assign ab05c3 = hmaster1_p & ab05be | !hmaster1_p & ab05c2;
assign dea6d1 = hlock2_p & dea6d0 | !hlock2_p & !deadba;
assign a5f96a = locked_p & a5f969 | !locked_p & a5fb6a;
assign adaec0 = hlock3_p & adaebf | !hlock3_p & v84563c;
assign a5ee40 = hbusreq2_p & a5ee3f | !hbusreq2_p & a5ee3e;
assign ab05b7 = hbusreq2_p & ab05b6 | !hbusreq2_p & ab05b5;
assign deac50 = hburst0 & deac4e | !hburst0 & deac4f;
assign ab0c77 = hready & ab0c76 | !hready & deada8;
assign deae38 = hbusreq3 & deae37 | !hbusreq3 & !v84563c;
assign b2669c = hbusreq2_p & b2669b | !hbusreq2_p & b2669a;
assign af34d8 = hmaster1_p & af34d4 | !hmaster1_p & af34d7;
assign cea36b = hbusreq3 & cea369 | !hbusreq3 & cea36a;
assign d40d41 = hgrant1_p & d40d3b | !hgrant1_p & !d40d33;
assign a5f2ec = hmaster1_p & a5f2eb | !hmaster1_p & a5f967;
assign deae1f = hlock2_p & deae1e | !hlock2_p & !deada8;
assign a5efb1 = hlock2 & a5f38f | !hlock2 & a5efb0;
assign a5ee5d = hbusreq1 & a5ee5c | !hbusreq1 & v84563c;
assign ab0bfd = hlock2 & ab0b88 | !hlock2 & ab0bfc;
assign c3bc91 = hlock0_p & b2671f | !hlock0_p & c3bc90;
assign a5eef8 = hmaster1_p & a5eef7 | !hmaster1_p & a5f6d9;
assign a5faad = hbusreq1_p & a60196 | !hbusreq1_p & !a60176;
assign cea37f = hbusreq2_p & cea37e | !hbusreq2_p & cea37d;
assign a9b9f0 = hbusreq3_p & a9b9ec | !hbusreq3_p & a9b9ef;
assign d40d86 = hbusreq2_p & d40d31 | !hbusreq2_p & d40d7b;
assign b26749 = hbusreq2_p & b266a3 | !hbusreq2_p & !b266a2;
assign c3bc81 = hbusreq2_p & c3bc80 | !hbusreq2_p & c3bc7f;
assign c3b76b = hbusreq2_p & c3b768 | !hbusreq2_p & c3b6ab;
assign a5eae8 = hlock0_p & a5eae7 | !hlock0_p & a5eae4;
assign ab05bf = locked_p & c3b6f9 | !locked_p & !v84563c;
assign a5f1a5 = hlock2 & a5f1a2 | !hlock2 & a5f1a4;
assign af3574 = hlock0_p & v84563c | !hlock0_p & af3573;
assign c3b88c = hbusreq2_p & c3b88b | !hbusreq2_p & c3b7b1;
assign a81ccd = hlock0_p & a81caa | !hlock0_p & v84563c;
assign a5f8b4 = hlock1_p & a60167 | !hlock1_p & a60168;
assign ab0636 = hlock0_p & ab056f | !hlock0_p & ab05f9;
assign a5f8e7 = hlock2 & a5f8d7 | !hlock2 & a5f8e6;
assign ab0bdb = hbusreq2_p & ab0bda | !hbusreq2_p & b29cbb;
assign b29ebd = hready & deae02 | !hready & !dead7b;
assign dea738 = hlock3_p & dea72c | !hlock3_p & dea737;
assign ce9cf5 = hbusreq2_p & cea1b7 | !hbusreq2_p & cea1b6;
assign a5ea5d = hbusreq2 & a5ea56 | !hbusreq2 & !a5ea5c;
assign a5f597 = hbusreq2_p & a5f593 | !hbusreq2_p & a5f4f1;
assign dead69 = hready_p & dead57 | !hready_p & dead68;
assign a5f8d0 = hgrant1_p & a60192 | !hgrant1_p & a5f8cf;
assign c3bdb6 = hlock2_p & c3bcee | !hlock2_p & v845660;
assign ce9e26 = decide_p & ce9e25 | !decide_p & a57859;
assign b26720 = locked_p & v84563c | !locked_p & b2671f;
assign a5fb95 = locked_p & a5fb94 | !locked_p & v84563c;
assign b29ab9 = hgrant0_p & c3bceb | !hgrant0_p & !b29ab8;
assign c3bd05 = hbusreq3 & c3bd04 | !hbusreq3 & !c3bcb3;
assign a5f35e = hgrant0_p & a5f346 | !hgrant0_p & a5f35d;
assign a5f573 = hlock1_p & v84563c | !hlock1_p & a5f572;
assign ab0c07 = hready & b2982c | !hready & dead7b;
assign deae13 = hlock2_p & deae12 | !hlock2_p & v84563c;
assign b29eb1 = hlock2_p & b29ea7 | !hlock2_p & !b29eb0;
assign c3b71f = hready & c3b71d | !hready & c3b71e;
assign a5ea6a = hbusreq2_p & a5f08a | !hbusreq2_p & a5ea69;
assign dead9f = hlock3_p & dead88 | !hlock3_p & dead9e;
assign a5eeb9 = hbusreq1_p & b2982c | !hbusreq1_p & !v84563c;
assign a5fce7 = hlock0_p & a5fcdf | !hlock0_p & a5fce6;
assign a60196 = start_p & v845654 | !start_p & !v9703fa;
assign ab058c = hmaster1_p & ab058b | !hmaster1_p & ab0b61;
assign b299a0 = hlock0_p & b2999f | !hlock0_p & !deae51;
assign c3bcfa = hbusreq2_p & c3bcf9 | !hbusreq2_p & v84563c;
assign a5f043 = decide_p & a5f042 | !decide_p & v84563c;
assign a5f1dd = locked_p & a5f1dc | !locked_p & v84563c;
assign a5f533 = hgrant1_p & a5f532 | !hgrant1_p & a5f4e5;
assign cea43a = hlock2_p & cea439 | !hlock2_p & cea414;
assign c3b707 = hlock2_p & c3b706 | !hlock2_p & !c3b647;
assign a5f96c = locked_p & v84563c | !locked_p & !a5f96b;
assign ab0616 = hmaster1_p & ab0615 | !hmaster1_p & ab0be5;
assign c3bd5f = hready & deac52 | !hready & v84563c;
assign a81cf1 = locked_p & a81cf0 | !locked_p & v84563c;
assign af3551 = hgrant2_p & af354f | !hgrant2_p & af3550;
assign a5fbb2 = locked_p & a5fbb1 | !locked_p & !v84563c;
assign cea24a = hburst1_p & v84563c | !hburst1_p & v8c6449;
assign dead57 = decide_p & dead56 | !decide_p & v84563c;
assign ab0c81 = decide_p & ab0c80 | !decide_p & v84563c;
assign a5f8ef = hbusreq2 & a5f8ee | !hbusreq2 & ab0cc3;
assign a5f538 = hbusreq2 & a5f527 | !hbusreq2 & !a5f537;
assign ab067b = hbusreq2_p & ab0679 | !hbusreq2_p & ab067a;
assign b8acf2 = jx1_p & b8acf1 | !jx1_p & v84563c;
assign a5f6fc = hlock2_p & a5f6f7 | !hlock2_p & a5f6fb;
assign cea2a5 = hlock0_p & cea2a4 | !hlock0_p & v84563c;
assign a5f829 = stateG10_1_p & v970407 | !stateG10_1_p & a5f828;
assign ab0632 = hlock2 & ab062b | !hlock2 & ab062d;
assign b29f91 = hlock2_p & b29f8e | !hlock2_p & !b29f90;
assign b2991b = hready & b29917 | !hready & b2991a;
assign b26786 = hbusreq2_p & b26785 | !hbusreq2_p & b266a0;
assign ab05f4 = hmaster1_p & ab05f3 | !hmaster1_p & ab0ade;
assign c3bdd0 = hready & c3bbd2 | !hready & deada8;
assign b29f5a = hlock2_p & b29f56 | !hlock2_p & !b29f59;
assign b29933 = hgrant2_p & b2992f | !hgrant2_p & b29932;
assign a5f837 = hmastlock_p & a5f711 | !hmastlock_p & !v84563c;
assign deae2b = hmaster0_p & deae2a | !hmaster0_p & !v84563c;
assign cea481 = hlock1_p & v84565a | !hlock1_p & !cea480;
assign cea1c1 = hlock2_p & cea1c0 | !hlock2_p & v84563c;
assign c3b7dc = hlock0_p & c3bd4b | !hlock0_p & cea887;
assign b29fff = hbusreq2_p & b29ffe | !hbusreq2_p & v84563c;
assign a5ee63 = hbusreq2 & a5ee62 | !hbusreq2 & a5fbc0;
assign deae1a = hlock3_p & v84563c | !hlock3_p & deae19;
assign b29828 = hlock2_p & v84563c | !hlock2_p & !b29827;
assign deae33 = hlock2_p & deae32 | !hlock2_p & !v84563c;
assign c3bd9c = hlock0_p & c3bd99 | !hlock0_p & !c3bd9b;
assign cea4af = decide_p & cea4ae | !decide_p & v84563c;
assign dea6d8 = hmaster1_p & dea6d7 | !hmaster1_p & !v84563c;
assign ab0c93 = hbusreq2_p & ab0c92 | !hbusreq2_p & cea15a;
assign c3bd7e = hmaster1_p & c3bc36 | !hmaster1_p & !c3bd7d;
assign deac18 = hgrant1_p & v84565a | !hgrant1_p & deac17;
assign ab0c27 = hlock2_p & ab0c26 | !hlock2_p & v84563c;
assign b29a9c = hmaster0_p & b29a95 | !hmaster0_p & b29a9b;
assign b2678c = hready_p & b26784 | !hready_p & b2678b;
assign cea457 = hbusreq2_p & cea456 | !hbusreq2_p & cea44a;
assign a5f076 = hbusreq0_p & a5f70b | !hbusreq0_p & v84563c;
assign b29a99 = hbusreq2_p & b29a98 | !hbusreq2_p & v84563c;
assign a5f40c = hbusreq1 & a5f40a | !hbusreq1 & a5f40b;
assign a5eebb = hready & a5eeb8 | !hready & a5eeba;
assign a5ef71 = hlock0_p & a5ef52 | !hlock0_p & a5ef5e;
assign b29f9a = locked_p & v84563c | !locked_p & c3bd9a;
assign a5f1bf = hmaster1_p & a5fbc5 | !hmaster1_p & a5f1be;
assign cea48f = hready_p & cea477 | !hready_p & cea48e;
assign b298a5 = hlock0_p & b298a4 | !hlock0_p & v84563c;
assign b29b1d = hlock0_p & deacdf | !hlock0_p & v84563c;
assign b29f8d = hlock0_p & b29ea6 | !hlock0_p & c3bd8e;
assign ab0c1a = hlock2_p & ab0b8c | !hlock2_p & v84563c;
assign ab060c = hlock2 & ab0513 | !hlock2 & ab060b;
assign a5edfe = hbusreq2_p & a5edf9 | !hbusreq2_p & a5edfd;
assign dea6f2 = hmaster0_p & dea6f1 | !hmaster0_p & !v84563c;
assign a5f964 = hlock0_p & a5fb7a | !hlock0_p & a5f71d;
assign dead46 = hbusreq2_p & dead45 | !hbusreq2_p & v84563c;
assign deae65 = hlock0_p & deae5a | !hlock0_p & !v84563c;
assign b840b0 = hgrant2_p & v84564b | !hgrant2_p & v845647;
assign a5eed4 = hmaster0_p & a5eecc | !hmaster0_p & a5eed3;
assign ab0b45 = hlock0_p & v84565a | !hlock0_p & ab0b44;
assign adaedc = hlock0_p & adaebd | !hlock0_p & v84563c;
assign cea0bb = hgrant1_p & v84565a | !hgrant1_p & cea0ba;
assign a5fcbe = hbusreq3 & a5fcbd | !hbusreq3 & v84563c;
assign dead18 = hlock1_p & v84563c | !hlock1_p & deacdf;
assign a5f8f1 = hbusreq2_p & a5f8f0 | !hbusreq2_p & !v845644;
assign a5eeea = hlock0_p & a5eee3 | !hlock0_p & !a5eee9;
assign a5fb2e = hbusreq2_p & a5fb2d | !hbusreq2_p & v84564d;
assign c3bcca = hbusreq3 & c3bcc7 | !hbusreq3 & c3bcc9;
assign a5f299 = hbusreq2_p & a5f298 | !hbusreq2_p & !v84563c;
assign ab057a = hmaster1_p & ab0579 | !hmaster1_p & ab0ade;
assign a5f3b3 = hbusreq1 & a5f38d | !hbusreq1 & c3b634;
assign a5f1fb = hbusreq2_p & a5f1fa | !hbusreq2_p & v84563c;
assign c3bce6 = locked_p & v84563c | !locked_p & !c3bce5;
assign a5ee3e = hbusreq2 & a5ee3d | !hbusreq2 & v845641;
assign deac11 = decide_p & deac10 | !decide_p & v84563c;
assign adaed9 = hmaster0_p & adaed8 | !hmaster0_p & v84563c;
assign b29947 = hready & b29946 | !hready & v845648;
assign a5f011 = decide_p & a5efed | !decide_p & a5f010;
assign b29e6e = hgrant2_p & b29e6d | !hgrant2_p & b29d21;
assign a5ea0e = hlock2_p & a5ea0d | !hlock2_p & a5f1a8;
assign ab05f9 = hbusreq0_p & b29942 | !hbusreq0_p & b29946;
assign ab053d = hready & ab053c | !hready & v84563c;
assign dead9a = hlock2_p & dead99 | !hlock2_p & !v84563c;
assign a5ee10 = hbusreq1 & a5ee0e | !hbusreq1 & a5ee0f;
assign a5fbfe = locked_p & a5fbfd | !locked_p & v84563c;
assign ab0704 = decide_p & ab0703 | !decide_p & v845662;
assign cea14b = hready & deacec | !hready & b266ab;
assign a81cab = hmaster1_p & a81caa | !hmaster1_p & v84563c;
assign c3bd97 = hgrant2_p & c3bc6d | !hgrant2_p & c3bd96;
assign a5ef37 = hlock0_p & a5ef36 | !hlock0_p & a5ee13;
assign dead54 = hbusreq3 & dead53 | !hbusreq3 & !v84563c;
assign c3bdab = hbusreq2_p & c3bdaa | !hbusreq2_p & dead2e;
assign c3b804 = hbusreq2_p & c3b803 | !hbusreq2_p & !c3b7b0;
assign af3c57 = locked_p & af3c55 | !locked_p & af3c56;
assign cea39e = locked_p & deae59 | !locked_p & !cea380;
assign a5ea75 = hlock0_p & a5f1f4 | !hlock0_p & a5ea40;
assign b29fea = hready_p & b29fd0 | !hready_p & b29fe9;
assign ab0cd3 = hlock2_p & ab0cd2 | !hlock2_p & v84563c;
assign deadc4 = hlock1_p & deadba | !hlock1_p & deadc3;
assign cea19c = hbusreq3 & cea199 | !hbusreq3 & cea19b;
assign c3bde1 = decide_p & c3bde0 | !decide_p & v845660;
assign b2996e = hlock0_p & b2996d | !hlock0_p & b29cfe;
assign a5ec32 = jx0_p & a5f047 | !jx0_p & a5ec31;
assign a5fc9e = hlock1_p & a5fc78 | !hlock1_p & a5fc9d;
assign ab0b52 = hlock0_p & c3bc48 | !hlock0_p & v84563c;
assign a5f237 = hlock0_p & a5f8c8 | !hlock0_p & a5f236;
assign c3bc3c = hlock0_p & deada8 | !hlock0_p & v84563c;
assign a5eb8b = hready & a5fb81 | !hready & !v84563c;
assign a5f06c = hbusreq2 & a5f069 | !hbusreq2 & a5f06b;
assign adaee1 = hgrant2_p & v84563c | !hgrant2_p & adaee0;
assign a81ca6 = hburst0_p & v84563c | !hburst0_p & !v845654;
assign a5fa23 = hbusreq2 & a5fa02 | !hbusreq2 & !a5fa22;
assign a5efc3 = hgrant2_p & a5efc2 | !hgrant2_p & v84563c;
assign b29f7b = hlock0_p & c3bd5f | !hlock0_p & c3bd61;
assign ab0cb8 = hmaster1_p & cea15a | !hmaster1_p & ab0cb7;
assign a5f345 = hmaster1_p & a5f344 | !hmaster1_p & a5f958;
assign b266ac = hlock1_p & v84563c | !hlock1_p & b266ab;
assign c3bc33 = hlock2_p & deadb2 | !hlock2_p & v84563c;
assign c3bd83 = hlock0_p & c3bc48 | !hlock0_p & !c3bcdb;
assign deada9 = stateG10_1_p & deacb4 | !stateG10_1_p & deada8;
assign c3bcbf = hready_p & c3bcb7 | !hready_p & c3bcbe;
assign ab05e6 = hbusreq0_p & b29832 | !hbusreq0_p & v8c6711;
assign c3bd92 = hmaster1_p & c3bc5e | !hmaster1_p & c3bd91;
assign c3bc41 = hbusreq3 & c3bc3c | !hbusreq3 & !c3bc21;
assign b299d3 = hmaster1_p & b299d2 | !hmaster1_p & b29e65;
assign cea47c = hlock0_p & cea47b | !hlock0_p & cea3cd;
assign ab0c3d = hready & v84563c | !hready & !c3bd3d;
assign b29ae9 = hgrant2_p & b29ae6 | !hgrant2_p & b29ae8;
assign a5fbd5 = hbusreq2_p & a5fbd4 | !hbusreq2_p & v84563c;
assign b29986 = locked_p & b29985 | !locked_p & v84563c;
assign a5f121 = hlock0_p & a5f120 | !hlock0_p & a5f108;
assign a5f6ea = locked_p & a5fb94 | !locked_p & a5f6e9;
assign a5f839 = stateG10_1_p & a5f838 | !stateG10_1_p & a5f837;
assign a60173 = hlock1_p & a60172 | !hlock1_p & v84563c;
assign c3b6ac = hbusreq2_p & c3b6aa | !hbusreq2_p & c3b6ab;
assign c3b7b3 = hbusreq3 & c3b7b2 | !hbusreq3 & !v845644;
assign b299f3 = hlock3_p & b299ef | !hlock3_p & b299f2;
assign b299e3 = hmaster1_p & b299e2 | !hmaster1_p & b29e96;
assign a5f41e = hready & a5f3f3 | !hready & a5f41d;
assign a5f834 = stateG10_1_p & v845654 | !stateG10_1_p & a5f833;
assign b29f47 = hmaster1_p & b29f39 | !hmaster1_p & b29f46;
assign a5e9df = hlock0_p & a5f919 | !hlock0_p & a5f144;
assign deae1d = hlock1_p & deac51 | !hlock1_p & !deae1c;
assign deadf3 = hmaster1_p & deadea | !hmaster1_p & !deadf2;
assign ab0b96 = locked_p & v84563c | !locked_p & b29d87;
assign c3bc2b = hbusreq2_p & c3bc22 | !hbusreq2_p & c3bc20;
assign b29abf = hlock2 & b29abc | !hlock2 & b29abe;
assign a5f95e = decide_p & a5f951 | !decide_p & a5f95d;
assign a5f1a2 = hlock0_p & v845641 | !hlock0_p & !v84563c;
assign b26694 = start_p & v84566c | !start_p & b26692;
assign a5f17d = hlock0_p & a5f177 | !hlock0_p & a5f17c;
assign c3bc66 = hlock0_p & c3bc65 | !hlock0_p & deacfc;
assign b29d51 = hready & deace1 | !hready & b266a2;
assign b26700 = hmaster1_p & b266f2 | !hmaster1_p & b266ff;
assign a5fb28 = hlock2 & a5fb27 | !hlock2 & ab0c32;
assign ab0c35 = hbusreq2_p & ab0c34 | !hbusreq2_p & ab0ad1;
assign ab0555 = hmaster1_p & ab0554 | !hmaster1_p & ab0bee;
assign b29fc1 = hready & b29fc0 | !hready & v84563c;
assign a5fc10 = hready & a5fc0b | !hready & a5fc0f;
assign ab0c2f = hlock0_p & v84563c | !hlock0_p & !ab0c2e;
assign af35ae = hgrant0_p & af35ab | !hgrant0_p & af35ad;
assign c3b82c = hmaster1_p & c3b82b | !hmaster1_p & c3bca4;
assign b29a3f = hbusreq3 & b29d60 | !hbusreq3 & b29a3e;
assign adaf12 = hmaster1_p & adaeeb | !hmaster1_p & v84563c;
assign d40d2d = hmaster1_p & d40d2c | !hmaster1_p & v84563c;
assign b29e54 = hmaster0_p & b29e4b | !hmaster0_p & !b29e53;
assign ab0c0e = hlock0_p & v84563c | !hlock0_p & c3bce6;
assign b29d8c = hlock0_p & b29d8b | !hlock0_p & !v84563c;
assign a5f11e = hgrant1_p & a5f11d | !hgrant1_p & a5f11b;
assign c3bc54 = hlock2_p & c3bc53 | !hlock2_p & dead2e;
assign a5f18b = hgrant1_p & a5fa1e | !hgrant1_p & a5f18a;
assign a5f7fd = hready & a5f7f9 | !hready & a5f7fc;
assign a5fa55 = hbusreq2 & a5fa42 | !hbusreq2 & a5fa41;
assign c3b739 = hlock0_p & deae59 | !hlock0_p & c3b738;
assign a81cee = hlock3_p & a81ced | !hlock3_p & a81cc6;
assign hmaster0 = a5785b;
assign a6016f = hmastlock_p & a6016e | !hmastlock_p & !v84563c;
assign cea331 = hlock1_p & v84563c | !hlock1_p & cea330;
assign d40d57 = hmaster1_p & d40d33 | !hmaster1_p & d40d42;
assign a5f8f8 = hmaster0_p & a5f888 | !hmaster0_p & a5f8f7;
assign a81d07 = hmaster0_p & a81d06 | !hmaster0_p & v84563c;
assign adaeec = hbusreq0_p & adaebd | !hbusreq0_p & adaeeb;
assign ab0bb1 = hbusreq3 & ab0bad | !hbusreq3 & ab0bb0;
assign cea40f = hlock0_p & cea40e | !hlock0_p & !cea405;
assign d40d60 = locked_p & v84563c | !locked_p & d40d33;
assign b2992c = hlock0_p & b2992b | !hlock0_p & !v84563c;
assign b29f1f = hready & deadc4 | !hready & c3bd3d;
assign a5f7cd = hlock0_p & a5f7cb | !hlock0_p & a5f7ba;
assign c3bcd2 = hgrant2_p & c3bc28 | !hgrant2_p & c3bc2b;
assign ce9cd9 = hlock3_p & ce9cd7 | !hlock3_p & ce9cd8;
assign dea79d = hready_p & dea76f | !hready_p & !dea79c;
assign a5f163 = hgrant2_p & a5f15f | !hgrant2_p & a5f162;
assign b29a64 = hlock1_p & c3b683 | !hlock1_p & b29a63;
assign c3bd8b = hready & cea2e7 | !hready & c3bd8a;
assign c3bc7d = hlock2_p & c3bc7c | !hlock2_p & !c3bc7b;
assign be34e8 = decide_p & be34df | !decide_p & be34e7;
assign a5f56a = hbusreq1_p & a60192 | !hbusreq1_p & v84563c;
assign b29f35 = hbusreq2_p & b29f34 | !hbusreq2_p & v84563c;
assign a5f931 = hgrant1_p & a5fb8b | !hgrant1_p & a5f930;
assign be34ea = hgrant3_p & be34e6 | !hgrant3_p & be34e9;
assign ab05cb = hlock2 & ab0d04 | !hlock2 & ab05ca;
assign b29f74 = hbusreq2_p & b29e69 | !hbusreq2_p & b29d36;
assign a5f361 = hgrant3_p & a5f2df | !hgrant3_p & a5f360;
assign ab06b5 = hlock0_p & c3bd60 | !hlock0_p & !v84563c;
assign a5fa15 = hlock1_p & a60177 | !hlock1_p & !a5fa14;
assign b2674a = hgrant2_p & b26749 | !hgrant2_p & !b2672c;
assign a5ef6d = hlock0_p & a5f36e | !hlock0_p & a5ef6b;
assign b2677a = hbusreq2_p & b26779 | !hbusreq2_p & b26736;
assign ab0c7b = hbusreq2_p & ab0c7a | !hbusreq2_p & !ab0b23;
assign c3bced = hmaster1_p & c3bce4 | !hmaster1_p & c3bcec;
assign a5f904 = hbusreq2_p & a5f903 | !hbusreq2_p & v84563c;
assign ab0b5d = hbusreq2_p & ab0b5b | !hbusreq2_p & ab0b5c;
assign cea423 = hbusreq3 & cea41e | !hbusreq3 & cea422;
assign a5f933 = hready & a5f932 | !hready & v84565a;
assign deaeb2 = hmaster1_p & deaeb1 | !hmaster1_p & dead2d;
assign a5ee14 = hbusreq0_p & a5f3a1 | !hbusreq0_p & a5ee13;
assign b29fde = hlock0_p & b29fdc | !hlock0_p & b29fdd;
assign af35b7 = hgrant2_p & af35b5 | !hgrant2_p & af35b6;
assign b26703 = hlock2_p & b266ca | !hlock2_p & b26695;
assign ab0cd1 = hgrant3_p & ab0c82 | !hgrant3_p & !ab0cd0;
assign b29915 = stateG10_1_p & v84563c | !stateG10_1_p & b29914;
assign af3497 = locked_p & af3c49 | !locked_p & d40d33;
assign deaeb5 = hbusreq2_p & deaeb0 | !hbusreq2_p & deaeb4;
assign deae4c = jx0_p & dead6b | !jx0_p & deae4b;
assign c3bd4c = hlock0_p & c3bd47 | !hlock0_p & !c3bd4b;
assign cea188 = hgrant2_p & cea86e | !hgrant2_p & cea877;
assign ab06aa = hgrant1_p & b29eea | !hgrant1_p & ab06a9;
assign af3c26 = hmaster1_p & af3c25 | !hmaster1_p & v845646;
assign b29fa0 = locked_p & b29f9f | !locked_p & !v84563c;
assign ab0641 = hmaster1_p & ab0c58 | !hmaster1_p & !ab0640;
assign b29eb6 = hburst0 & dead7a | !hburst0 & b29eb5;
assign af34e0 = hmaster0_p & af34d8 | !hmaster0_p & af34df;
assign deacf5 = hburst1 & deacf4 | !hburst1 & v84563c;
assign af3c3b = hmaster1_p & af3c22 | !hmaster1_p & !v84563c;
assign c3b620 = hbusreq3_p & c3bde3 | !hbusreq3_p & !c3b61f;
assign a5f70a = locked_p & a5f709 | !locked_p & !v84563c;
assign ab0c18 = hmaster1_p & ab0ace | !hmaster1_p & ab0c17;
assign ab064d = hmaster1_p & cea15a | !hmaster1_p & ab0bbb;
assign cea1bc = hbusreq1_p & cea1bb | !hbusreq1_p & v84563c;
assign a5ef70 = hbusreq3 & a5ef62 | !hbusreq3 & a5ef6f;
assign b29e65 = hgrant2_p & b29cd5 | !hgrant2_p & b29cd8;
assign a5f57d = hgrant1_p & a5f56e | !hgrant1_p & a5f56d;
assign b2982b = start_p & cea1aa | !start_p & b2982a;
assign a5f435 = stateG10_1_p & v970407 | !stateG10_1_p & a5f434;
assign ab0c20 = hlock0_p & v84563c | !hlock0_p & !c3bce5;
assign ce9e0b = hgrant0_p & cea85f | !hgrant0_p & ce9e0a;
assign c3bdde = hmaster1_p & c3bddd | !hmaster1_p & c3bd50;
assign ab0c04 = hready & b2982c | !hready & !v84563c;
assign cea2a0 = hready & cea29e | !hready & cea29f;
assign a5f3ad = hbusreq3 & a5f3a7 | !hbusreq3 & a5fbc0;
assign a5eeef = hlock0_p & a5eeee | !hlock0_p & a5eee9;
assign ab06f1 = hgrant2_p & ab06db | !hgrant2_p & ab0679;
assign b29f9d = locked_p & b29f9c | !locked_p & !v84563c;
assign a5f0ab = hbusreq0_p & c3bcf8 | !hbusreq0_p & v84563c;
assign a5fc0a = hbusreq1_p & a5fc09 | !hbusreq1_p & a5fba2;
assign deacb5 = stateG10_1_p & deacb4 | !stateG10_1_p & deaca1;
assign c3bdfe = hmaster0_p & c3bdfd | !hmaster0_p & c3bd92;
assign c3b7d7 = hgrant2_p & c3b7d3 | !hgrant2_p & c3b7d6;
assign a5f3bd = hlock2_p & a5f3b9 | !hlock2_p & a5f3bc;
assign a5fd3b = hready_p & v84563c | !hready_p & a5fd3a;
assign ce9cbf = hready & c98b96 | !hready & v845646;
assign b29d1e = hbusreq2_p & b29d17 | !hbusreq2_p & v84565a;
assign b29a7b = hlock0_p & c3bd5f | !hlock0_p & !v84563c;
assign a5efd2 = hbusreq2_p & a5efd1 | !hbusreq2_p & a5ef61;
assign ab06a6 = hbusreq2_p & ab06a4 | !hbusreq2_p & ab06a2;
assign a5ef2c = hbusreq2 & a5ee00 | !hbusreq2 & a5fd12;
assign cea430 = hlock0_p & cea42f | !hlock0_p & cea3cd;
assign ab052a = hbusreq2_p & ab0528 | !hbusreq2_p & ab0529;
assign a5f4e9 = hbusreq1 & a5f4e8 | !hbusreq1 & a5f493;
assign a5f200 = hbusreq2 & a5f1ff | !hbusreq2 & a5f72b;
assign a5efbc = hbusreq2_p & a5ee64 | !hbusreq2_p & a5efbb;
assign ab063c = hready_p & ab0625 | !hready_p & !ab063b;
assign b29ed7 = hlock2_p & c3bce5 | !hlock2_p & !v84563c;
assign dea6ee = hready_p & dea6e5 | !hready_p & dea6ed;
assign ab0b18 = hlock2_p & ab0b16 | !hlock2_p & !ab0b17;
assign a5f978 = hlock2 & a5fc45 | !hlock2 & a5f6f8;
assign cea437 = hbusreq2_p & cea436 | !hbusreq2_p & cea420;
assign ab0ca3 = hgrant2_p & ab0b70 | !hgrant2_p & ab0ca2;
assign af34b1 = hbusreq2_p & af34b0 | !hbusreq2_p & af34af;
assign c3b6c4 = hlock1_p & c3bbd2 | !hlock1_p & c3b6c3;
assign a5f3cc = hbusreq1_p & a5fc87 | !hbusreq1_p & !v84563c;
assign af34a0 = hlock0_p & af3c57 | !hlock0_p & af3c4c;
assign ce9d30 = hbusreq2_p & cea2a2 | !hbusreq2_p & cea2a1;
assign a5fca8 = stateG10_1_p & v84563c | !stateG10_1_p & a5fc6a;
assign ab075e = hgrant3_p & ab073f | !hgrant3_p & !ab075d;
assign b29993 = locked_p & deae59 | !locked_p & !b29992;
assign a5fb8a = hmastlock_p & a5fb89 | !hmastlock_p & v84563c;
assign ab0bb8 = hmaster1_p & dead2e | !hmaster1_p & !ab0bb7;
assign ab0652 = decide_p & ab0649 | !decide_p & !v845662;
assign c3b627 = hlock0_p & c3b623 | !hlock0_p & !c3b626;
assign a5fc19 = hlock2_p & a5fc15 | !hlock2_p & a5fc18;
assign a5fa89 = hlock0_p & a5fa88 | !hlock0_p & v84563c;
assign a5fca4 = hbusreq1_p & a5fc87 | !hbusreq1_p & a5fc8f;
assign a5f4ec = hbusreq2 & a5f4ba | !hbusreq2 & !a5f4eb;
assign a5fb2b = hlock0_p & a5fb2a | !hlock0_p & v84563c;
assign c3bdbb = hbusreq1_p & v84563c | !hbusreq1_p & !c3bdba;
assign v970420 = hlock2_p & v9703fc | !hlock2_p & v84563c;
assign a5f5a8 = hready & a5f4a6 | !hready & c3b6a0;
assign ab0c43 = hready & v84563c | !hready & !deaca2;
assign ab0bc5 = hlock3_p & ab0bb6 | !hlock3_p & ab0bc4;
assign af34af = hlock0_p & af34ae | !hlock0_p & af3c5e;
assign b2677c = hmaster1_p & b2677b | !hmaster1_p & b26730;
assign c3b79b = hlock0_p & cea1bf | !hlock0_p & !dead7f;
assign ab0af7 = hbusreq2_p & ab0af5 | !hbusreq2_p & ab0af6;
assign ab06ed = hgrant2_p & ab06ea | !hgrant2_p & ab06ec;
assign adaec7 = stateG10_1_p & adaec6 | !stateG10_1_p & adaec4;
assign dead72 = locked_p & dead6e | !locked_p & v84563c;
assign c3b6e3 = hlock0_p & c3b626 | !hlock0_p & c3b6e1;
assign a5fbdc = stateG10_1_p & v84563c | !stateG10_1_p & a5fb72;
assign a5fa6c = hready & v84563c | !hready & c98b95;
assign af34f4 = hgrant2_p & d40d60 | !hgrant2_p & af34f3;
assign a5e9e9 = hbusreq0 & a5e9e8 | !hbusreq0 & a5f15c;
assign a5f786 = hlock1_p & a60172 | !hlock1_p & a5f785;
assign ab0645 = hbusreq2_p & ab0bda | !hbusreq2_p & ab0bd9;
assign af355f = hlock2_p & af352c | !hlock2_p & v84563c;
assign deae97 = hbusreq2_p & deae96 | !hbusreq2_p & !v84563c;
assign b29a6f = hmaster1_p & b29a6d | !hmaster1_p & b29a6e;
assign a5f72a = hlock0_p & a5fb6b | !hlock0_p & a5f729;
assign b8acd9 = hmaster0_p & b8acd8 | !hmaster0_p & v8c6711;
assign b29a8d = hbusreq2_p & b29a8c | !hbusreq2_p & !b29ce7;
assign af34a7 = hlock0_p & af3c50 | !hlock0_p & af3c6b;
assign ab0ba7 = hlock2 & ab0ba2 | !hlock2 & ab0ba6;
assign dea7a3 = hmaster0_p & dea7a1 | !hmaster0_p & dea7a2;
assign a5ea7f = hlock0_p & a5ea7e | !hlock0_p & a5ea54;
assign a81cc5 = hmaster1_p & v84563c | !hmaster1_p & a81cb5;
assign b29e5f = decide_p & b29e5e | !decide_p & v84563c;
assign a5ede0 = hbusreq2_p & a5eddc | !hbusreq2_p & a5eddb;
assign af3c1f = hbusreq2_p & af3c1d | !hbusreq2_p & af3c1c;
assign a5ee3a = hlock0_p & a60141 | !hlock0_p & a5ee39;
assign ab0cfc = hmaster1_p & ab0bf1 | !hmaster1_p & !ab0cfb;
assign cea381 = locked_p & dead7d | !locked_p & !cea380;
assign a5f374 = hbusreq1_p & a5f704 | !hbusreq1_p & v84563c;
assign a5f741 = hbusreq0_p & a5f6e9 | !hbusreq0_p & a5f727;
assign b26739 = hlock2_p & b266b2 | !hlock2_p & !b266bc;
assign ab06a0 = hgrant2_p & ab069c | !hgrant2_p & ab069f;
assign af34eb = hmaster0_p & af34e8 | !hmaster0_p & af34ea;
assign dead8b = locked_p & v84563c | !locked_p & dead8a;
assign a5f148 = hlock1_p & a5f8d2 | !hlock1_p & !v84563c;
assign af3568 = hmaster0_p & af3552 | !hmaster0_p & af3567;
assign c3b815 = hbusreq2_p & c3b7a5 | !hbusreq2_p & c3b814;
assign bdb583 = decide_p & bdb582 | !decide_p & v845660;
assign a81cb3 = hgrant1_p & a81cb2 | !hgrant1_p & a81cb1;
assign b29f0b = hmastlock_p & b29f0a | !hmastlock_p & v84563c;
assign a5f992 = hready & a5fc48 | !hready & !a5fbab;
assign b26766 = decide_p & b26754 | !decide_p & b26765;
assign af34bc = hlock0_p & af34b9 | !hlock0_p & af34bb;
assign c3bd43 = hbusreq3 & c3bd25 | !hbusreq3 & c3bd42;
assign dead11 = hbusreq3 & dead10 | !hbusreq3 & v84563c;
assign c3bd64 = hbusreq2_p & c3bd63 | !hbusreq2_p & c3bc21;
assign v856555 = hmaster0_p & v84564a | !hmaster0_p & !v94aab7;
assign cea371 = hgrant3_p & cea357 | !hgrant3_p & cea370;
assign ab0bd7 = hbusreq2_p & ab0bd6 | !hbusreq2_p & v845644;
assign a5f205 = hmaster0_p & a5f1fd | !hmaster0_p & a5f204;
assign dea745 = hbusreq2_p & deadb4 | !hbusreq2_p & deadb3;
assign ab0aec = stateG10_1_p & c3bd38 | !stateG10_1_p & ab0aeb;
assign deadd1 = hlock0_p & deadd0 | !hlock0_p & !v84563c;
assign cea1b7 = hlock2_p & cea1b6 | !hlock2_p & v84563c;
assign a5fb9e = hburst1_p & d5edb8 | !hburst1_p & !d615cf;
assign d40d67 = hmastlock_p & d40d66 | !hmastlock_p & v84563c;
assign a5efb8 = hbusreq0_p & a5ee66 | !hbusreq0_p & a5efb7;
assign a5f9c5 = hbusreq2_p & a5f9c4 | !hbusreq2_p & v84563c;
assign a5f1b5 = hbusreq2 & a5f1b4 | !hbusreq2 & v84563c;
assign b29fbb = hmaster1_p & c3bceb | !hmaster1_p & b29fba;
assign dead20 = hbusreq0_p & b26695 | !hbusreq0_p & !deacdf;
assign cea388 = hmaster1_p & cea387 | !hmaster1_p & cea860;
assign c3b654 = hbusreq3 & c3b650 | !hbusreq3 & !c3b653;
assign a5ee44 = hready & a5ee43 | !hready & !c3b622;
assign cea320 = hburst0 & v84563c | !hburst0 & cea31f;
assign c3bcdd = hlock0_p & c3bcda | !hlock0_p & !c3bcdc;
assign ab0af0 = hlock0_p & v84563c | !hlock0_p & !ab0aef;
assign a5f845 = hlock2 & a5f82c | !hlock2 & a5f844;
assign b26712 = hmaster1_p & b2670d | !hmaster1_p & b26711;
assign a5e9f2 = hlock0_p & a5e9f1 | !hlock0_p & a5f171;
assign deae75 = hgrant1_p & deada9 | !hgrant1_p & deae74;
assign af35ba = hmaster1_p & af3571 | !hmaster1_p & af356f;
assign b29ae6 = hbusreq3 & b29d0f | !hbusreq3 & b29ae5;
assign a5f8c3 = hlock1_p & v84563c | !hlock1_p & a5f8c2;
assign a5f32a = hbusreq2_p & a5f329 | !hbusreq2_p & a5fa6b;
assign ab0b3e = hbusreq2_p & ab0b3a | !hbusreq2_p & v84563c;
assign ab0b83 = hbusreq3 & ab0b7f | !hbusreq3 & ab0b82;
assign cea1a3 = hgrant2_p & cea86e | !hgrant2_p & cea0c0;
assign c98ba2 = decide_p & c98b96 | !decide_p & c98ba1;
assign c3b66c = hlock0_p & c3b665 | !hlock0_p & !c3b66b;
assign c3bda4 = hmaster0_p & c3bda0 | !hmaster0_p & c3bda3;
assign a5f2d8 = hbusreq2_p & a5f2d7 | !hbusreq2_p & !v84563c;
assign a5fc31 = hbusreq2_p & a5fc30 | !hbusreq2_p & a5fc2f;
assign a5f488 = hlock1_p & a81cf0 | !hlock1_p & a5f487;
assign dea7b5 = jx2_p & deae4c | !jx2_p & dea7b4;
assign c3b6f4 = hgrant0_p & c3b6e7 | !hgrant0_p & c3b6f3;
assign ab0756 = hlock0_p & b29f3c | !hlock0_p & !ab0737;
assign cea254 = hlock1_p & v84563c | !hlock1_p & !cea253;
assign c3b704 = hmaster1_p & c3b702 | !hmaster1_p & c3b703;
assign a5eb4b = hbusreq0 & a5ea60 | !hbusreq0 & a5f096;
assign cea339 = hbusreq3 & cea299 | !hbusreq3 & cea337;
assign c3b7ad = hlock0_p & c3bce5 | !hlock0_p & v84563c;
assign a5f255 = hmaster1_p & a5f254 | !hmaster1_p & a5f887;
assign a5f884 = hlock2_p & a5f87b | !hlock2_p & a5f883;
assign deacee = hlock0_p & deaced | !hlock0_p & !deacdf;
assign c3b8b5 = decide_p & c3b8b4 | !decide_p & v845660;
assign a5eb41 = hbusreq2_p & a5eb3d | !hbusreq2_p & !a5eb40;
assign a5ead3 = hlock0_p & a5f92e | !hlock0_p & a5ead1;
assign ab0d03 = hlock0_p & b298a4 | !hlock0_p & !b29826;
assign deae53 = hlock2_p & deae52 | !hlock2_p & !deae51;
assign v970448 = hmaster1_p & v84563c | !hmaster1_p & v970447;
assign c3bd3c = hgrant1_p & cea270 | !hgrant1_p & deadb9;
assign b26732 = hlock2_p & b2669a | !hlock2_p & b266b8;
assign b2a020 = hmastlock_p & b2a01f | !hmastlock_p & !v84563c;
assign a5efe8 = hlock0_p & a5f575 | !hlock0_p & !a5f36e;
assign a5f9f8 = hgrant1_p & v84563c | !hgrant1_p & a5f9f7;
assign ce9d47 = hlock0_p & dead72 | !hlock0_p & cea17a;
assign cea343 = hlock2_p & cea342 | !hlock2_p & v84563c;
assign c3b709 = hgrant2_p & c3b708 | !hgrant2_p & v845660;
assign d40d95 = hbusreq2_p & d40d94 | !hbusreq2_p & d40d33;
assign cea2ad = hlock1_p & deada8 | !hlock1_p & !c98b95;
assign b26734 = hlock1_p & v84563c | !hlock1_p & b266a0;
assign c3b7e6 = hlock0_p & c3bd60 | !hlock0_p & v84563c;
assign c3bc6d = hbusreq2_p & c3bc6c | !hbusreq2_p & !v84563c;
assign c3b684 = hlock1_p & c3b683 | !hlock1_p & deadc3;
assign b29fe0 = hlock2_p & b29fdb | !hlock2_p & !b29fdf;
assign a5fbe7 = hbusreq1 & v84563c | !hbusreq1 & a5fbe6;
assign a5eff8 = hmaster1_p & a5edfc | !hmaster1_p & v84563c;
assign c3b6b7 = hmaster0_p & c3b690 | !hmaster0_p & c3b6b6;
assign af3c7b = hlock1_p & af3c49 | !hlock1_p & af3c7a;
assign ab0be0 = hmaster1_p & ab0b61 | !hmaster1_p & ab0b6b;
assign a5f37e = hready & a5f37c | !hready & a5f37d;
assign a5ee01 = hmaster1_p & a5edfe | !hmaster1_p & a5ee00;
assign dead29 = hmaster1_p & dead1d | !hmaster1_p & dead28;
assign ab05f6 = hbusreq2_p & ab0562 | !hbusreq2_p & ab05f5;
assign af34c8 = hlock2_p & af34c7 | !hlock2_p & af3c64;
assign cea4ac = hgrant2_p & cea4a9 | !hgrant2_p & cea4ab;
assign b29ec5 = locked_p & v84563c | !locked_p & !c3bc51;
assign a5eeb7 = hbusreq1_p & a5fc7d | !hbusreq1_p & !v84563c;
assign cea2e5 = hmastlock_p & cea2e4 | !hmastlock_p & v84563c;
assign c3b890 = hlock0_p & c3bd99 | !hlock0_p & !ce9df1;
assign dead67 = hmaster0_p & dead60 | !hmaster0_p & !dead66;
assign b29a57 = hlock3_p & b29a47 | !hlock3_p & b29a56;
assign a5f02a = hmaster0_p & v84563c | !hmaster0_p & a5f029;
assign ce9cfa = hbusreq2_p & cea149 | !hbusreq2_p & cea342;
assign c3b74e = hbusreq2_p & c3b74d | !hbusreq2_p & c3b6db;
assign a5f20b = hbusreq2 & a5fc81 | !hbusreq2 & v84563c;
assign d40d98 = hmaster1_p & d40d97 | !hmaster1_p & d40d47;
assign c3b691 = hbusreq1_p & deada8 | !hbusreq1_p & !v84565a;
assign ab076b = jx0_p & ab0656 | !jx0_p & ab076a;
assign c3bcac = hmaster1_p & c3bcab | !hmaster1_p & !c3bca4;
assign a5f0b1 = decide_p & a5f0a2 | !decide_p & a5f0b0;
assign c3b733 = hbusreq3 & c3b6e0 | !hbusreq3 & c3b732;
assign ab057f = hlock2_p & ab057e | !hlock2_p & ab0572;
assign a5eee8 = hbusreq1 & a5eee7 | !hbusreq1 & v84563c;
assign adaed0 = hgrant2_p & adaecd | !hgrant2_p & adaecf;
assign b29d01 = hlock0_p & b29d00 | !hlock0_p & !deada8;
assign c3b7b2 = hbusreq2_p & c3b7b0 | !hbusreq2_p & !c3b7b1;
assign b26788 = hgrant2_p & b26786 | !hgrant2_p & b26787;
assign a5ef42 = hbusreq3 & a5ef3c | !hbusreq3 & a5fbc0;
assign ab0ce3 = hmaster0_p & ab0ce0 | !hmaster0_p & ab0ce2;
assign ce9df0 = hgrant2_p & cea344 | !hgrant2_p & !ce9def;
assign b2675a = hmaster1_p & b266c1 | !hmaster1_p & !b26759;
assign a5f748 = hmaster1_p & v84563c | !hmaster1_p & a5f747;
assign adaefd = hlock3_p & adaefc | !hlock3_p & adaed5;
assign b266fd = hbusreq2_p & b266fc | !hbusreq2_p & b266fb;
assign cea25b = hbusreq2_p & cea25a | !hbusreq2_p & v84563c;
assign a60189 = hbusreq1 & a60169 | !hbusreq1 & a60188;
assign dead34 = locked_p & dead33 | !locked_p & v84563c;
assign a5f036 = hready_p & a5f035 | !hready_p & a5f02c;
assign ab0b88 = hlock0_p & v84563c | !hlock0_p & !b29d5d;
assign a5f981 = hbusreq1_p & a5fba6 | !hbusreq1_p & a5f980;
assign af349f = hbusreq2_p & af349e | !hbusreq2_p & af349c;
assign deae9d = hmaster1_p & deae9c | !hmaster1_p & !dead5f;
assign ab06de = hlock2_p & ab0b80 | !hlock2_p & b29a4d;
assign a5fcd4 = start_p & v845652 | !start_p & a5fcd3;
assign deae87 = hlock2_p & deae86 | !hlock2_p & !deadc4;
assign a5f586 = hbusreq2_p & a5f568 | !hbusreq2_p & a5f55c;
assign a5edf8 = locked_p & v84563c | !locked_p & a5edf7;
assign c3b63a = locked_p & v84563c | !locked_p & v845648;
assign d40d75 = hmaster0_p & d40d71 | !hmaster0_p & d40d74;
assign b29910 = decide_p & b2990f | !decide_p & v84563c;
assign bdb5b5 = hmaster1_p & bdb5b4 | !hmaster1_p & !bdb589;
assign b29d95 = hlock2_p & v845660 | !hlock2_p & b29d94;
assign a81cc1 = hbusreq2_p & a81cc0 | !hbusreq2_p & v84563c;
assign ab0bf9 = hbusreq3_p & ab0bc9 | !hbusreq3_p & ab0bf8;
assign a5f7a4 = hlock2 & a5f78e | !hlock2 & a5f7a3;
assign c3bc9d = hmaster1_p & c3bc8f | !hmaster1_p & c3bc9c;
assign ab0cf5 = hgrant0_p & ab0cea | !hgrant0_p & !ab0cf4;
assign ab06e9 = hlock2_p & ab06e8 | !hlock2_p & ab067f;
assign a5f95a = hbusreq2 & a5fd10 | !hbusreq2 & v84563c;
assign a5e9e0 = hbusreq2 & a5f146 | !hbusreq2 & a5e9df;
assign b29f43 = hlock2_p & b29f3e | !hlock2_p & !b29f42;
assign a5f230 = hready & a60168 | !hready & !deaca1;
assign af3c14 = hbusreq2_p & af3c13 | !hbusreq2_p & af3c12;
assign bdb5ad = hgrant3_p & bdb59c | !hgrant3_p & bdb5ac;
assign a9b9d6 = hlock0_p & a9b9d0 | !hlock0_p & v845660;
assign a5fb71 = hmastlock_p & a5fb70 | !hmastlock_p & v84563c;
assign a5f8fe = hgrant1_p & v84563c | !hgrant1_p & a5f8fd;
assign deae55 = hbusreq2_p & dead81 | !hbusreq2_p & dead80;
assign ab0731 = hgrant3_p & ab06da | !hgrant3_p & !ab0730;
assign ab0688 = hlock3_p & ab067e | !hlock3_p & ab0687;
assign d40d9d = hbusreq3_p & d40d8d | !hbusreq3_p & d40d9c;
assign a5ef12 = hready & a5ef0f | !hready & a5ef11;
assign ab069d = hbusreq2_p & ab068f | !hbusreq2_p & ab068d;
assign af3582 = hmaster1_p & v84563c | !hmaster1_p & af3581;
assign a5fcdb = hlock0_p & a5fcd2 | !hlock0_p & a5fcda;
assign b29fc8 = hgrant2_p & v845660 | !hgrant2_p & !b29c3c;
assign ab0bf2 = hbusreq2_p & ab0b24 | !hbusreq2_p & b29cbb;
assign cea16e = hlock0_p & cea16d | !hlock0_p & v845660;
assign b29eee = hlock0_p & b29eed | !hlock0_p & c3bd5f;
assign af3597 = hmaster1_p & v84563c | !hmaster1_p & af356f;
assign b29d73 = hbusreq3 & b29d72 | !hbusreq3 & b29c3c;
assign af3c4b = start_p & v84563c | !start_p & !af3c4a;
assign a5f39f = locked_p & v84563c | !locked_p & a5f39e;
assign c3bcb1 = hready_p & c3bcb0 | !hready_p & c3bc45;
assign ab05d8 = decide_p & ab0585 | !decide_p & !v845662;
assign a5f864 = hready & a60171 | !hready & a5f863;
assign d40d83 = locked_p & d40d81 | !locked_p & d40d82;
assign b29940 = hlock1_p & deac52 | !hlock1_p & !b8acdb;
assign c3bbf5 = hmaster1_p & deac3f | !hmaster1_p & c3bbf4;
assign af34f9 = hgrant0_p & af34f2 | !hgrant0_p & af34f8;
assign a5fd23 = hready & v84563c | !hready & !deadd5;
assign ab06c5 = hmaster0_p & ab06a8 | !hmaster0_p & ab06c4;
assign a5ef5e = hbusreq0_p & a5f4fc | !hbusreq0_p & a5edcc;
assign c3b7a8 = hbusreq3 & c3b7a7 | !hbusreq3 & cea15a;
assign deaea1 = hlock1_p & deadde | !hlock1_p & !deacbd;
assign c3b6cb = hready & c3b6c4 | !hready & deada8;
assign b29b36 = hbusreq3_p & b29b0b | !hbusreq3_p & b29b35;
assign a5fc5d = hlock2 & a5fc5b | !hlock2 & a5fc5c;
assign a5f821 = hbusreq2 & a5f807 | !hbusreq2 & !ab0c31;
assign a5fa62 = hlock1_p & a6016f | !hlock1_p & !a5fa61;
assign adaee8 = hgrant0_p & adaede | !hgrant0_p & adaee7;
assign ab054a = hlock1_p & v84563c | !hlock1_p & ab0549;
assign cea3ec = hlock2_p & cea3eb | !hlock2_p & cea3ea;
assign b26778 = hbusreq2_p & b26777 | !hbusreq2_p & b266a0;
assign c3b640 = hlock0_p & c3bbbb | !hlock0_p & c3b63f;
assign cea329 = hgrant2_p & v84563c | !hgrant2_p & !cea328;
assign a5fccc = locked_p & v84563c | !locked_p & c3bd60;
assign a5f384 = hmaster1_p & a5f383 | !hmaster1_p & a60145;
assign b29b19 = hmaster0_p & b29b17 | !hmaster0_p & b29b18;
assign ab068e = hlock0_p & c3bd5f | !hlock0_p & !ab068c;
assign ab052d = hbusreq2_p & ab052c | !hbusreq2_p & b29832;
assign cea0f3 = decide_p & cea0f2 | !decide_p & v84563c;
assign a5ef99 = hbusreq2 & a5ef96 | !hbusreq2 & a5ef98;
assign ab066b = hlock0_p & b29ea6 | !hlock0_p & !ab066a;
assign cea322 = hlock1_p & deae02 | !hlock1_p & cea321;
assign af3560 = hbusreq1_p & af352c | !hbusreq1_p & v84563c;
assign a81cd3 = hmaster1_p & v84563c | !hmaster1_p & a81cd2;
assign a5ef94 = decide_p & a5ef90 | !decide_p & !a5ef93;
assign a5f1d7 = locked_p & a5f1d6 | !locked_p & a5f6e9;
assign adaf0d = hmaster0_p & adaf09 | !hmaster0_p & adaf0c;
assign cea3fb = hready & cea3fa | !hready & deae59;
assign a5f98b = hready & a5f98a | !hready & a5fbb0;
assign a5ea52 = hready & a5ea51 | !hready & a5fc01;
assign b29a1e = decide_p & b299f3 | !decide_p & b29e57;
assign b299d7 = locked_p & v84563c | !locked_p & cea38d;
assign a5f6e1 = hready_p & a5f6cf | !hready_p & a5f6e0;
assign b29ce9 = hlock0_p & b29ce8 | !hlock0_p & !v84563c;
assign b2673a = hbusreq2_p & b26739 | !hbusreq2_p & !b266bc;
assign cea294 = hlock1_p & v84563c | !hlock1_p & !cea293;
assign a5f1af = hready & a5f1ac | !hready & a5f1ae;
assign a5fbbd = hbusreq3 & a5fbbc | !hbusreq3 & a60144;
assign ab0b23 = hlock0_p & v84565a | !hlock0_p & ab0b22;
assign a5f58c = hready & v84563c | !hready & c3b697;
assign a5f330 = hbusreq2_p & a5f8cc | !hbusreq2_p & v84563c;
assign a5ef83 = hlock0_p & a5f565 | !hlock0_p & a5ef81;
assign bdb58c = hbusreq2_p & v84565a | !hbusreq2_p & !bdb58b;
assign dea6e3 = hmaster1_p & dea6e2 | !hmaster1_p & dead54;
assign b29ac4 = hmaster0_p & b29aac | !hmaster0_p & b29ac3;
assign b840af = hready_p & v84564f | !hready_p & b840ae;
assign a5fae2 = hbusreq2_p & a5fad7 | !hbusreq2_p & a5fad6;
assign ab0bac = hlock2 & ab0ba9 | !hlock2 & ab0bab;
assign b29b08 = hlock3_p & b29aef | !hlock3_p & b29a9c;
assign b266bc = hlock0_p & b26695 | !hlock0_p & b266bb;
assign a5f43f = hbusreq1 & a5f43d | !hbusreq1 & !a5f43e;
assign c3b71a = hgrant1_p & c3b719 | !hgrant1_p & deae7f;
assign af3506 = hmaster0_p & af3505 | !hmaster0_p & af34e4;
assign a5ea9d = hbusreq2 & a5ea9b | !hbusreq2 & a5ea9c;
assign c3bc78 = hbusreq3 & c3bc74 | !hbusreq3 & c3bc77;
assign a5f8bf = hready & a5fb8b | !hready & a5f8be;
assign deaeae = locked_p & v84563c | !locked_p & !deae5a;
assign ab0566 = hbusreq2_p & ab0562 | !hbusreq2_p & ab0565;
assign ab0cc8 = hbusreq3 & ab0cc1 | !hbusreq3 & ab0cc7;
assign a5fccf = hbusreq2_p & a5fccd | !hbusreq2_p & a5fcce;
assign cea379 = locked_p & cea377 | !locked_p & !cea378;
assign a5f392 = hbusreq2_p & a5f38a | !hbusreq2_p & a5f391;
assign a5f38f = hready & a5f38c | !hready & !a5f38e;
assign a5fa01 = hlock0_p & a5f9fa | !hlock0_p & a5fa00;
assign b29fd0 = decide_p & b29fcf | !decide_p & b29e57;
assign ab055d = hlock1_p & deaca0 | !hlock1_p & !ab055c;
assign b29eea = stateG10_1_p & b29ee8 | !stateG10_1_p & b29ee9;
assign ab0548 = stateG10_1_p & v84563c | !stateG10_1_p & ab0547;
assign a5eeaa = hbusreq2_p & a5eea9 | !hbusreq2_p & a5ee69;
assign af34a9 = hbusreq2_p & af34a8 | !hbusreq2_p & af34a6;
assign c3bdb4 = hmaster1_p & dead2e | !hmaster1_p & c3bdb3;
assign a5f192 = hbusreq0_p & a5fb20 | !hbusreq0_p & ab0c31;
assign b8acd8 = hmaster1_p & v8c6711 | !hmaster1_p & !v84563c;
assign af350b = hmaster1_p & d40d97 | !hmaster1_p & af3487;
assign ab0bb9 = hmaster0_p & dead2e | !hmaster0_p & ab0bb8;
assign b29932 = hbusreq3 & b29930 | !hbusreq3 & b29931;
assign a5f72d = hlock2_p & a5f72c | !hlock2_p & v84563c;
assign decide = !a5ec33;
assign af3c12 = hlock0_p & af3c11 | !hlock0_p & v845646;
assign dea7a8 = hmaster1_p & dea7a7 | !hmaster1_p & dea752;
assign b2a01d = jx0_p & b29ea4 | !jx0_p & b2a01c;
assign dead2e = hlock0_p & v845660 | !hlock0_p & !v84563c;
assign a5f2f7 = hbusreq2 & a5f2f3 | !hbusreq2 & a5f2f6;
assign deacdf = hmastlock_p & deacde | !hmastlock_p & v84563c;
assign ab0bf1 = hgrant2_p & ab0bf0 | !hgrant2_p & ab0b0f;
assign a5f396 = hlock0_p & a5f385 | !hlock0_p & a5f394;
assign a5f902 = hbusreq2 & a5f8b9 | !hbusreq2 & a5f901;
assign a5f271 = hmaster0_p & a5f26a | !hmaster0_p & a5f270;
assign a5f346 = hmaster0_p & a5f345 | !hmaster0_p & a5f270;
assign a5f391 = hlock0_p & a60141 | !hlock0_p & a5f390;
assign c3b728 = hmaster1_p & c3b727 | !hmaster1_p & c3bccf;
assign c3b7c3 = hbusreq2_p & c3b7c2 | !hbusreq2_p & !c3b7c1;
assign a5f3f3 = hbusreq1 & a5f3f2 | !hbusreq1 & v84563c;
assign c3b736 = hbusreq2_p & c3b652 | !hbusreq2_p & c3b735;
assign c3bda8 = hbusreq2_p & c3bda7 | !hbusreq2_p & dead2e;
assign b26785 = hlock2_p & b266f0 | !hlock2_p & b266a0;
assign b29d39 = hlock2 & b29cfe | !hlock2 & deada8;
assign ab0cd2 = hlock0_p & v84563c | !hlock0_p & !c3bd8d;
assign ab05f2 = hbusreq2_p & ab0564 | !hbusreq2_p & ab05f1;
assign a5f26f = hbusreq0 & a5f26c | !hbusreq0 & !a5f26e;
assign cea35d = hbusreq2_p & cea35c | !hbusreq2_p & cea15a;
assign b266b5 = hbusreq2_p & b266b4 | !hbusreq2_p & b266b2;
assign a5f9c8 = hbusreq2_p & a5f9c4 | !hbusreq2_p & a5f9c3;
assign a5ea4f = hlock0_p & a5ea4c | !hlock0_p & a5ea4e;
assign a5f977 = hbusreq2 & a5f972 | !hbusreq2 & a5f976;
assign b26701 = hmaster0_p & b266e6 | !hmaster0_p & b26700;
assign a81ce9 = hmaster0_p & a81ce5 | !hmaster0_p & a81ce8;
assign c3b7dd = hlock2_p & c3b7db | !hlock2_p & !c3b7dc;
assign ab05d6 = hlock3_p & ab05bb | !hlock3_p & ab05d5;
assign c3b88e = hbusreq2_p & c3b88d | !hbusreq2_p & c3b814;
assign af3576 = hmaster0_p & af3570 | !hmaster0_p & af3575;
assign ab0733 = hmaster1_p & ab0732 | !hmaster1_p & ab0681;
assign a5f15c = hlock0_p & a5f15b | !hlock0_p & v84563c;
assign a5eede = hlock2_p & a5eedb | !hlock2_p & a5eedd;
assign c3bcfc = hbusreq3 & c3bcfa | !hbusreq3 & c3bcfb;
assign d40d62 = hmaster0_p & d40d61 | !hmaster0_p & d40d60;
assign cea2a8 = hbusreq3 & cea2a3 | !hbusreq3 & cea2a7;
assign adaf07 = locked_p & adaf06 | !locked_p & v84563c;
assign a5f730 = hmaster1_p & a60145 | !hmaster1_p & a5f72f;
assign c3bcb7 = decide_p & c3bcb6 | !decide_p & !v845660;
assign a5f855 = hbusreq2 & a5f845 | !hbusreq2 & ab0c31;
assign af34c7 = hlock0_p & af34ae | !hlock0_p & af3c62;
assign a5f37b = locked_p & a5f37a | !locked_p & !v845641;
assign b266a6 = hbusreq2_p & b266a5 | !hbusreq2_p & b266a4;
assign ab0cff = hready_p & ab0cf6 | !hready_p & !ab0cfe;
assign b29d75 = hmaster1_p & b29d64 | !hmaster1_p & b29d74;
assign c3b7b4 = hmaster1_p & c3b7b3 | !hmaster1_p & v84563c;
assign a5e9ff = hlock2_p & a5e9fe | !hlock2_p & a5f196;
assign b29fbe = hbusreq2_p & b29fbd | !hbusreq2_p & v84563c;
assign af3c18 = decide_p & af3c17 | !decide_p & v8567b4;
assign a5f7fc = hlock1_p & a60177 | !hlock1_p & !a5f7fb;
assign cea345 = hbusreq3 & cea344 | !hbusreq3 & v84563c;
assign af3595 = hmaster0_p & af3594 | !hmaster0_p & af3567;
assign v970430 = hready_p & v970401 | !hready_p & v97042f;
assign ce9dfc = hlock0_p & cea2f1 | !hlock0_p & !ce9df1;
assign af34a2 = hlock2_p & af34a0 | !hlock2_p & af34a1;
assign a5fae4 = hbusreq2_p & a5fa8c | !hbusreq2_p & a5fa89;
assign a5eb74 = hbusreq0 & a5f198 | !hbusreq0 & v845641;
assign a81cfc = hgrant2_p & a81cfb | !hgrant2_p & v84563c;
assign b266a7 = hmaster1_p & b2669c | !hmaster1_p & !b266a6;
assign c3bc89 = hbusreq3 & c3bc88 | !hbusreq3 & c3bc6d;
assign ab06c3 = hgrant2_p & ab06b6 | !hgrant2_p & ab06c2;
assign v84566c = stateA1_p & v84563c | !stateA1_p & !v84563c;
assign cea372 = hbusreq3_p & cea340 | !hbusreq3_p & cea371;
assign deae90 = hlock1_p & deac52 | !hlock1_p & !c98b95;
assign c3b7a1 = hlock2_p & c3bc75 | !hlock2_p & c3b7a0;
assign a5f0a9 = hbusreq0 & a5f0a8 | !hbusreq0 & v84563c;
assign b29941 = hlock1_p & v84563c | !hlock1_p & !b8acdb;
assign a5f53b = hlock1_p & deac52 | !hlock1_p & a5f53a;
assign ce9cb5 = hbusreq2_p & ce9cb4 | !hbusreq2_p & cea448;
assign ce9e1f = hbusreq2_p & cea367 | !hbusreq2_p & cea366;
assign a5fcda = hbusreq0_p & a5fcd2 | !hbusreq0_p & !a5fcd9;
assign b29e66 = hmaster1_p & b29e61 | !hmaster1_p & b29e65;
assign cea4ad = hmaster1_p & cea4ac | !hmaster1_p & !deacaa;
assign a5f387 = locked_p & v84563c | !locked_p & a5f36e;
assign b29a68 = hbusreq2_p & b29a67 | !hbusreq2_p & !b29a66;
assign deac17 = hbusreq1_p & v84565a | !hbusreq1_p & v84563c;
assign ce9ccb = hmaster0_p & ce9cca | !hmaster0_p & !cea419;
assign d40d33 = hmastlock_p & d40d32 | !hmastlock_p & v84563c;
assign b29fdc = hready & deadba | !hready & deadb9;
assign a6016b = hburst1_p & c06d34 | !hburst1_p & c07311;
assign cea258 = hready & cea254 | !hready & cea257;
assign b29a6c = hbusreq3 & b29a6a | !hbusreq3 & b29a6b;
assign dead77 = locked_p & dead76 | !locked_p & v84563c;
assign a81ca7 = stateG2_p & v84563c | !stateG2_p & c07311;
assign d40d9b = hready_p & d40d76 | !hready_p & d40d9a;
assign af354b = hgrant1_p & af3546 | !hgrant1_p & af352e;
assign a5f13d = hgrant2_p & a5f136 | !hgrant2_p & a5f13c;
assign a5f0b0 = hmaster0_p & a5f0aa | !hmaster0_p & a5f0af;
assign b266a0 = hmastlock_p & b2669f | !hmastlock_p & v84563c;
assign a5fc83 = start_p & a81ca6 | !start_p & a5fc82;
assign b29ab3 = hlock0_p & deacfb | !hlock0_p & !v84563c;
assign a5eddf = hbusreq2_p & a5edd6 | !hbusreq2_p & a5edd5;
assign cea455 = hmaster1_p & cea454 | !hmaster1_p & cea15d;
assign ab0b5f = hlock0_p & ab0b5e | !hlock0_p & v84563c;
assign a81ce0 = hmaster0_p & v84563c | !hmaster0_p & a81cdf;
assign c3bce7 = hlock0_p & c3bc52 | !hlock0_p & c3bce6;
assign bdb5ac = hready_p & bdb5a2 | !hready_p & bdb5ab;
assign a5ef95 = hready_p & a5ef48 | !hready_p & a5ef94;
assign b299d1 = hbusreq3 & b299d0 | !hbusreq3 & b2995f;
assign b29e96 = hgrant2_p & b29e95 | !hgrant2_p & !b29c3c;
assign c3bc49 = hlock0_p & c3bc48 | !hlock0_p & !v84563c;
assign a5ef15 = hlock0_p & a5edf2 | !hlock0_p & a5ef14;
assign deaeb6 = hlock1_p & deae02 | !hlock1_p & v84563c;
assign a57859 = hgrant0_p & v84563c | !hgrant0_p & v845666;
assign a5fbbb = hbusreq2_p & a5fbba | !hbusreq2_p & a5fbb4;
assign a5f996 = hlock2_p & a5f991 | !hlock2_p & !a5f995;
assign c3b6d2 = hmaster0_p & c3b6b9 | !hmaster0_p & c3b6d1;
assign af3507 = hmaster1_p & af3c4c | !hmaster1_p & af34e7;
assign c3b647 = locked_p & v84563c | !locked_p & c3b625;
assign c3b7f8 = hlock2_p & c3b7f7 | !hlock2_p & c3b7e4;
assign ab0b31 = hbusreq3 & ab0b2f | !hbusreq3 & ab0b30;
assign deae54 = hbusreq2_p & deae53 | !hbusreq2_p & deae52;
assign cea24c = stateA1_p & v8c607d | !stateA1_p & cea24b;
assign b2996d = hready & c3b6c5 | !hready & v84563c;
assign c3bcb0 = decide_p & c3bcaf | !decide_p & v845660;
assign a5fccd = hbusreq2 & a5fccb | !hbusreq2 & a5fccc;
assign ab0bf8 = hgrant3_p & ab0bdf | !hgrant3_p & !ab0bf7;
assign b29cf6 = hlock0_p & c3bc02 | !hlock0_p & v84565a;
assign a5e9ad = hbusreq2_p & a5f1a9 | !hbusreq2_p & v845641;
assign a81cd1 = locked_p & a81cd0 | !locked_p & v84563c;
assign a5f236 = hready & a60167 | !hready & !deaca1;
assign deae8d = hgrant2_p & deae89 | !hgrant2_p & deae8c;
assign b298a7 = hbusreq2_p & b298a6 | !hbusreq2_p & v84563c;
assign b8aceb = hmaster1_p & b8acea | !hmaster1_p & !v84563c;
assign c3b730 = locked_p & v84563c | !locked_p & !c3b72f;
assign a5ef2e = hmaster1_p & a5ef2b | !hmaster1_p & a5ef2d;
assign ab0bbe = hgrant2_p & ab0bbc | !hgrant2_p & ab0bbd;
assign b29d76 = hbusreq1_p & deae02 | !hbusreq1_p & deacf7;
assign a5f87d = hready & a5f87c | !hready & a60197;
assign a5f06b = hlock0_p & a5f06a | !hlock0_p & a5f067;
assign ce9d28 = hgrant2_p & ce9d26 | !hgrant2_p & ce9d27;
assign ce9dc6 = hgrant2_p & cea2a7 | !hgrant2_p & ce9d31;
assign deae80 = hgrant1_p & deadbb | !hgrant1_p & deae7f;
assign b29fe3 = hbusreq2_p & b29fd5 | !hbusreq2_p & v84563c;
assign a81cb6 = hmaster1_p & a81cb4 | !hmaster1_p & a81cb5;
assign dead24 = locked_p & v84563c | !locked_p & !b2671f;
assign ab060b = hlock0_p & b298a4 | !hlock0_p & ab05af;
assign ab0be7 = hmaster0_p & ab0be6 | !hmaster0_p & ab0be3;
assign dead3f = hbusreq3 & dead3e | !hbusreq3 & dead39;
assign b2982c = hmastlock_p & b2982b | !hmastlock_p & !v84563c;
assign ab051c = hlock2_p & ab051a | !hlock2_p & ab051b;
assign ab06d8 = hlock3_p & ab06c5 | !hlock3_p & ab06d7;
assign a5ef0f = hbusreq1 & a5ef0e | !hbusreq1 & !v84563c;
assign cea360 = hgrant2_p & cea159 | !hgrant2_p & !cea35f;
assign b2990d = hbusreq3 & b29909 | !hbusreq3 & b2990c;
assign ab0718 = hbusreq2_p & ab0717 | !hbusreq2_p & ab0716;
assign c3bcdf = hbusreq2_p & c3bcde | !hbusreq2_p & c3bbbc;
assign a5f739 = hready & v84563c | !hready & deace1;
assign a60172 = hmastlock_p & deac4e | !hmastlock_p & !v84563c;
assign ab0b9a = hgrant2_p & ab0b94 | !hgrant2_p & ab0b99;
assign a5f9f7 = hbusreq1_p & v84563c | !hbusreq1_p & a60172;
assign a5fc38 = hbusreq2 & a5fb6c | !hbusreq2 & a5fbc1;
assign b299ab = hready_p & b299a9 | !hready_p & b299aa;
assign ab0b6c = hbusreq3 & ab0b69 | !hbusreq3 & ab0b6b;
assign cea32c = hmaster0_p & cea32a | !hmaster0_p & cea32b;
assign b29e47 = hmaster0_p & b29d9d | !hmaster0_p & b29d9c;
assign b29cf2 = hready & v84565a | !hready & !v84563c;
assign a5e9c8 = hlock2_p & a5e9c7 | !hlock2_p & a5f196;
assign a5eb85 = hbusreq0 & a5eb3f | !hbusreq0 & !v84563c;
assign a5f584 = hbusreq2_p & a5f583 | !hbusreq2_p & !a5f582;
assign dead4a = hgrant2_p & dead3f | !hgrant2_p & dead48;
assign cea3f8 = hready & cea3f7 | !hready & cea3bf;
assign ab0748 = hgrant2_p & ab06df | !hgrant2_p & ab0747;
assign b2670d = hbusreq2_p & b2670c | !hbusreq2_p & b2670a;
assign a5efe5 = hbusreq0 & a5efe3 | !hbusreq0 & !a5efe4;
assign v970441 = hlock0_p & v9703fd | !hlock0_p & v970440;
assign b29ec6 = locked_p & v84563c | !locked_p & c3bce5;
assign a5f0ee = hbusreq0 & a5f0dc | !hbusreq0 & a5f0ed;
assign c3b689 = hlock2_p & c3b687 | !hlock2_p & !c3b686;
assign a5f949 = hlock2_p & a5f948 | !hlock2_p & a5f8ef;
assign cea251 = stateG10_1_p & cea249 | !stateG10_1_p & cea250;
assign c3bd24 = hlock2_p & c3bd22 | !hlock2_p & !deadb2;
assign a5eadc = hlock0_p & ab0c31 | !hlock0_p & a5eada;
assign ab0b78 = hlock0_p & v84563c | !hlock0_p & b29d52;
assign af3c46 = hgrant3_p & af3c42 | !hgrant3_p & af3c45;
assign ab0b80 = hlock0_p & b29ec5 | !hlock0_p & v845660;
assign c3b634 = hlock1_p & deacdf | !hlock1_p & !v84563c;
assign b29d8b = locked_p & v84563c | !locked_p & !b29d8a;
assign a5f136 = hbusreq3 & a5f0ee | !hbusreq3 & !a5f135;
assign deac7e = hgrant2_p & deac79 | !hgrant2_p & deac7d;
assign a5ef90 = hmaster0_p & a5ef76 | !hmaster0_p & a5ef8f;
assign c3bc36 = hbusreq2_p & c3bc35 | !hbusreq2_p & !v84563c;
assign a5f72c = hbusreq2 & a5f72a | !hbusreq2 & a5f72b;
assign a5f9d9 = hburst1_p & v845672 | !hburst1_p & !v84563c;
assign a5f746 = hbusreq2_p & a5f745 | !hbusreq2_p & v84563c;
assign b266e4 = hbusreq2_p & b266e2 | !hbusreq2_p & b266e1;
assign a81caa = locked_p & a81ca9 | !locked_p & v84563c;
assign cea416 = hbusreq2_p & cea415 | !hbusreq2_p & cea414;
assign d40d51 = hlock0_p & d40d50 | !hlock0_p & d40d33;
assign deae52 = hlock0_p & deae4f | !hlock0_p & !deae51;
assign b29983 = hready & deae4e | !hready & !v84563c;
assign b29928 = stateG10_1_p & v84563c | !stateG10_1_p & b29927;
assign ab06db = hbusreq2_p & ab0679 | !hbusreq2_p & ab0683;
assign dead28 = hgrant2_p & dead23 | !hgrant2_p & dead27;
assign cea49b = hlock2_p & cea49a | !hlock2_p & cea405;
assign c3b674 = start_p & deac4a | !start_p & b26692;
assign b29e5c = hbusreq3 & v84563c | !hbusreq3 & !v84564a;
assign ab0591 = hbusreq0_p & b298aa | !hbusreq0_p & b29990;
assign ab0cef = hbusreq2_p & ab0c9e | !hbusreq2_p & cea18f;
assign a5f1e8 = hlock2_p & a5f1e7 | !hlock2_p & !a5f995;
assign cea16b = hlock2_p & cea16a | !hlock2_p & v845660;
assign c3bdf6 = decide_p & c3bdf5 | !decide_p & !v845660;
assign a9b9d3 = hlock3_p & a9b9d2 | !hlock3_p & bdb581;
assign c3b76c = hgrant2_p & c3b769 | !hgrant2_p & c3b76b;
assign b29b32 = hmaster0_p & b29b17 | !hmaster0_p & !b29b31;
assign a5f3c1 = hmaster0_p & a5f3ae | !hmaster0_p & a5f3c0;
assign deada8 = hmastlock_p & deada7 | !hmastlock_p & v84563c;
assign b2a00b = hmaster0_p & b2a008 | !hmaster0_p & b2a00a;
assign c3bda0 = hmaster1_p & c3bd97 | !hmaster1_p & c3bd9f;
assign ab0cf9 = hmaster1_p & ab0cf8 | !hmaster1_p & ab0c49;
assign a5ee3c = hbusreq2 & a5ee3b | !hbusreq2 & a5fbc0;
assign a5eb92 = hbusreq0 & a5eb91 | !hbusreq0 & a5ea3e;
assign a5fa56 = hlock2_p & a5fa55 | !hlock2_p & v84563c;
assign ab0ce6 = hlock0_p & v845660 | !hlock0_p & !c3bcef;
assign a81d00 = decide_p & a81cee | !decide_p & a81cff;
assign a5f1c3 = hlock2_p & a5f1c2 | !hlock2_p & v84563c;
assign a5ead6 = hlock2_p & a5ead2 | !hlock2_p & a5ead5;
assign ab0647 = hmaster1_p & ab0c73 | !hmaster1_p & !ab0646;
assign c3bc77 = hbusreq2_p & c3bc76 | !hbusreq2_p & !v84563c;
assign a5edbe = hready & a5f515 | !hready & c3b6c4;
assign adaf1a = hready_p & adaefa | !hready_p & adaf19;
assign a5fbab = hmastlock_p & a5fbaa | !hmastlock_p & !v84563c;
assign c3b6c8 = hlock2_p & c3b6c7 | !hlock2_p & c3b698;
assign ab0bcd = decide_p & ab0bcc | !decide_p & v84563c;
assign c3b84d = hbusreq3 & c3b846 | !hbusreq3 & c3b84c;
assign c3bdcc = hlock3_p & c3bda5 | !hlock3_p & c3bdcb;
assign a5f286 = hmaster1_p & a5f282 | !hmaster1_p & a5f285;
assign a5edf5 = locked_p & v84563c | !locked_p & a5edeb;
assign a5f8c5 = hbusreq0_p & v84563c | !hbusreq0_p & v845641;
assign b26710 = hlock2_p & b2670e | !hlock2_p & b2670f;
assign cea296 = hlock0_p & cea295 | !hlock0_p & v84563c;
assign c3b7c2 = hlock2_p & c3b7bd | !hlock2_p & !c3b7c1;
assign a5f233 = hready & v84563c | !hready & !ab0aeb;
assign dead61 = hbusreq2_p & deacbf | !hbusreq2_p & v84563c;
assign adaf0a = hbusreq2_p & adaed7 | !hbusreq2_p & adaf00;
assign a5f909 = hbusreq2 & a5f907 | !hbusreq2 & a5f908;
assign b29fcd = hmaster0_p & b29fc7 | !hmaster0_p & b29fcc;
assign ab058a = hlock2_p & ab0588 | !hlock2_p & ab0589;
assign a5f208 = hbusreq2 & c3bcf8 | !hbusreq2 & v84563c;
assign a5eb99 = hmaster1_p & a5eb98 | !hmaster1_p & a5ea4a;
assign a5f7be = hready & a5f9f6 | !hready & v84563c;
assign deae68 = hlock0_p & deae67 | !hlock0_p & v84563c;
assign a5fbe6 = hlock1_p & a5fbe5 | !hlock1_p & v84563c;
assign a5ea51 = hlock1_p & a5fc78 | !hlock1_p & a5ea50;
assign cea1b8 = hbusreq2_p & cea1b7 | !hbusreq2_p & cea85d;
assign af34f0 = hlock3_p & af34ef | !hlock3_p & af3495;
assign a5eec1 = hbusreq1_p & a5fc8f | !hbusreq1_p & !v84563c;
assign adaecb = hmaster1_p & adaec9 | !hmaster1_p & adaeca;
assign a5fb9f = hburst0_p & d5edb8 | !hburst0_p & a5fb9e;
assign b29829 = hbusreq2_p & b29828 | !hbusreq2_p & v84563c;
assign b2995c = hbusreq2_p & b2995b | !hbusreq2_p & !b2994a;
assign b29ac1 = hbusreq2_p & b29ac0 | !hbusreq2_p & b29ab4;
assign c3b6e0 = locked_p & v84563c | !locked_p & !c3b635;
assign c3b62f = hbusreq3 & c3b629 | !hbusreq3 & c3b62e;
assign a5f490 = hgrant1_p & a5f486 | !hgrant1_p & a5f485;
assign a5f944 = hlock0_p & a5f943 | !hlock0_p & v845641;
assign adaef8 = hmaster0_p & adaef4 | !hmaster0_p & adaef7;
assign a5ee93 = hmaster0_p & a5ee82 | !hmaster0_p & a5ee92;
assign ab0b44 = hbusreq0_p & b29d34 | !hbusreq0_p & deacbe;
assign dea701 = jx1_p & dea6f0 | !jx1_p & dea700;
assign ce9d40 = hmaster0_p & ce9d37 | !hmaster0_p & ce9d3f;
assign cea3d9 = stateG10_1_p & deacb4 | !stateG10_1_p & cea3d8;
assign b29f0a = hburst0 & deadb9 | !hburst0 & b29f09;
assign b29a77 = hlock1_p & v84565a | !hlock1_p & !b29a76;
assign cea385 = hlock2_p & cea384 | !hlock2_p & cea383;
assign c3b6f9 = hready & c3b6f8 | !hready & !deae50;
assign adaed2 = hmaster1_p & adaed0 | !hmaster1_p & adaed1;
assign a5fd28 = hbusreq2_p & a5fd27 | !hbusreq2_p & v84563c;
assign cea325 = locked_p & cea324 | !locked_p & !dead0a;
assign ab0cd4 = hbusreq2_p & ab0cd3 | !hbusreq2_p & v845644;
assign a5f420 = hbusreq2 & a5f40d | !hbusreq2 & a5f41f;
assign cea0f4 = hready_p & cea862 | !hready_p & cea0f3;
assign ab0c7d = hgrant2_p & ab0c7b | !hgrant2_p & ab0c7c;
assign c3bd89 = hmaster1_p & c3bd85 | !hmaster1_p & c3bd88;
assign ab06ce = hlock2_p & ab06cd | !hlock2_p & b29a7b;
assign a5ee17 = hlock0_p & a5f36f | !hlock0_p & a5ee14;
assign ab063f = hmaster1_p & ab0ad2 | !hmaster1_p & ab0bee;
assign a5f096 = hbusreq2_p & a5f095 | !hbusreq2_p & v845641;
assign a5e9bc = hbusreq0_p & a5fb30 | !hbusreq0_p & ab0c31;
assign c3b8ab = hlock2_p & c3b7ea | !hlock2_p & !c3b7e6;
assign ab0c2e = hready & b29a5a | !hready & !v84565a;
assign cea289 = hgrant2_p & cea287 | !hgrant2_p & cea288;
assign a5fa21 = hready & a5fa1b | !hready & a5fa20;
assign b29fdd = hready & deadba | !hready & !v84563c;
assign cea464 = hlock2_p & cea463 | !hlock2_p & cea44d;
assign v8c607d = stateG2_p & v84563c | !stateG2_p & v8c6449;
assign a5f438 = hbusreq1 & a5f437 | !hbusreq1 & !v84563c;
assign ce9d36 = hgrant2_p & ce9d34 | !hgrant2_p & ce9d35;
assign a5fa86 = hgrant1_p & v84563c | !hgrant1_p & ab055a;
assign ab0643 = hmaster1_p & v84563c | !hmaster1_p & ab0ade;
assign cea295 = hready & cea292 | !hready & cea294;
assign adaeed = hlock0_p & adaebd | !hlock0_p & adaeec;
assign b29d56 = hbusreq3 & b29d55 | !hbusreq3 & c3bceb;
assign deacbf = hlock0_p & deacbe | !hlock0_p & v84563c;
assign a5f2fa = hgrant2_p & a5fbc4 | !hgrant2_p & a5f2f9;
assign cea159 = hbusreq2_p & cea85e | !hbusreq2_p & v84563c;
assign v845658 = hmaster1_p & v84563c | !hmaster1_p & !v84563c;
assign c3bcce = hgrant2_p & c3bcca | !hgrant2_p & c3bccd;
assign a5e9b3 = hready & a5fa59 | !hready & !c3bc09;
assign a5ee0a = hbusreq2_p & a5ee09 | !hbusreq2_p & a5ee05;
assign c3b830 = decide_p & c3b82f | !decide_p & v845660;
assign deacb3 = start_p & v845652 | !start_p & v84563c;
assign dead14 = hlock0_p & deacfa | !hlock0_p & deace9;
assign ab0593 = hlock0_p & deae51 | !hlock0_p & !ab0591;
assign v845641 = hready & v84563c | !hready & !v84563c;
assign ab0b7d = hlock0_p & v84563c | !hlock0_p & !b29d66;
assign a5fca7 = hready & a5fca1 | !hready & a5fca6;
assign a5fc0f = hlock1_p & a5fbab | !hlock1_p & a5fc0e;
assign ab0653 = hready_p & ab0651 | !hready_p & !ab0652;
assign a5f6f0 = hlock0_p & a5f6ed | !hlock0_p & a5f6ef;
assign c3b768 = hlock2_p & c3b6ab | !hlock2_p & !c3b6a1;
assign ab06ff = hgrant2_p & ab06fc | !hgrant2_p & ab06fe;
assign ab0b17 = hlock0_p & deada8 | !hlock0_p & !deac86;
assign d40d84 = hgrant2_p & d40d60 | !hgrant2_p & d40d83;
assign deadf8 = locked_p & v84563c | !locked_p & !dead8a;
assign cea877 = hbusreq2_p & cea86d | !hbusreq2_p & cea86c;
assign cea39a = hmaster0_p & cea388 | !hmaster0_p & cea399;
assign dea6bb = hlock2_p & dea6ba | !hlock2_p & v84563c;
assign v97045a = decide_p & v97042d | !decide_p & v97044d;
assign ab0670 = hlock0_p & v845660 | !hlock0_p & !dead7f;
assign a5eb4c = hbusreq3 & a5eb4b | !hbusreq3 & v84563c;
assign b29f9f = hready & c3bdbd | !hready & v84563c;
assign dea730 = hbusreq2_p & dead95 | !hbusreq2_p & dead94;
assign a5fa14 = hgrant1_p & a5fa12 | !hgrant1_p & a5fa13;
assign b29fa5 = hgrant2_p & c3bcfb | !hgrant2_p & !b29fa4;
assign a5ee7e = hgrant0_p & a5ee36 | !hgrant0_p & a5ee7d;
assign b8ace2 = hready_p & b8acd9 | !hready_p & b8ace1;
assign cea173 = hbusreq3 & cea172 | !hbusreq3 & cea15c;
assign ab0bc3 = hmaster0_p & ab0bbf | !hmaster0_p & ab0bc2;
assign a5ef73 = hbusreq2_p & a5f593 | !hbusreq2_p & a5ef6d;
assign a5f96e = hlock0_p & a5f96a | !hlock0_p & a5f96d;
assign a5f1a7 = hlock2 & v845641 | !hlock2 & v84563c;
assign b29f7c = hlock2 & b29f7a | !hlock2 & b29f7b;
assign a5ea23 = hbusreq3 & a5ea20 | !hbusreq3 & !a5ea22;
assign a5f380 = hlock0_p & a5f37b | !hlock0_p & !a5f37f;
assign b29fd8 = hlock1_p & v84565a | !hlock1_p & !b29fd7;
assign a5fb2d = hlock2_p & a5fb29 | !hlock2_p & a5fb2c;
assign c3bdd2 = hlock2_p & c3bdd1 | !hlock2_p & !deada8;
assign a5f027 = hbusreq0 & a5f026 | !hbusreq0 & v845644;
assign deacf0 = hbusreq3 & deacef | !hbusreq3 & v84563c;
assign cea2ee = hmaster0_p & cea1c4 | !hmaster0_p & cea2ed;
assign b266ab = hbusreq1_p & b266a0 | !hbusreq1_p & v84563c;
assign ab0acc = hlock2_p & ab0acb | !hlock2_p & cea15a;
assign a5f92c = hbusreq2_p & a5fd27 | !hbusreq2_p & v84564d;
assign cea332 = hgrant1_p & deadb9 | !hgrant1_p & cea271;
assign cea4a9 = hbusreq3 & cea49e | !hbusreq3 & cea422;
assign c3bcd5 = decide_p & c3bcd4 | !decide_p & v845660;
assign c3b7e8 = hlock0_p & c3bdcf | !hlock0_p & !deada8;
assign b29cbf = hbusreq2_p & b29cbc | !hbusreq2_p & v84563c;
assign ab050e = hbusreq3 & ab0d06 | !hbusreq3 & ab050d;
assign a5f29c = hbusreq3 & a5f299 | !hbusreq3 & a5f29b;
assign a5fcd5 = hmastlock_p & a5fcd4 | !hmastlock_p & !v84563c;
assign c3bc9b = hbusreq3 & c3bc9a | !hbusreq3 & c3bc70;
assign b29e52 = hgrant2_p & b29e51 | !hgrant2_p & b29e49;
assign a5fd05 = hbusreq2 & a5fcd2 | !hbusreq2 & !a5fcdf;
assign af34f5 = hmaster1_p & d40d60 | !hmaster1_p & af34f4;
assign a5f4e3 = hlock1_p & a60187 | !hlock1_p & a5f4c9;
assign a81ccb = decide_p & a81cc7 | !decide_p & a81cca;
assign cea425 = hbusreq2_p & cea421 | !hbusreq2_p & cea420;
assign deae4e = hlock1_p & deacf7 | !hlock1_p & !deae4d;
assign a5ec31 = jx1_p & a5ebee | !jx1_p & a5ec30;
assign deaeb1 = hbusreq2_p & deaeb0 | !hbusreq2_p & deaeaf;
assign cea369 = hbusreq2_p & cea367 | !hbusreq2_p & !cea197;
assign a5f95b = hbusreq2_p & a5f95a | !hbusreq2_p & v84563c;
assign af3c66 = hbusreq2_p & af3c65 | !hbusreq2_p & af3c63;
assign d40d6e = hlock1_p & d40d2b | !hlock1_p & d40d6d;
assign a5f9c3 = hlock0_p & a5f9c2 | !hlock0_p & v84563c;
assign deadfa = hlock2_p & deadf9 | !hlock2_p & v84563c;
assign c3b803 = hlock2_p & c3bc94 | !hlock2_p & !c3b7b0;
assign a5eed6 = decide_p & a5eeb5 | !decide_p & a5eed5;
assign deac60 = hbusreq3 & deac5f | !hbusreq3 & v84563c;
assign b2a008 = hmaster1_p & b2a006 | !hmaster1_p & b2a007;
assign ab0c41 = hbusreq2_p & ab0c40 | !hbusreq2_p & v84563c;
assign c3bd50 = hgrant2_p & c3bd4e | !hgrant2_p & c3bd4f;
assign a81ced = hmaster0_p & a81cec | !hmaster0_p & a81cc3;
assign a5f940 = hbusreq1_p & a5f8dd | !hbusreq1_p & a60193;
assign dead1c = hbusreq3 & dead1b | !hbusreq3 & v84563c;
assign ab063b = decide_p & ab063a | !decide_p & !v845662;
assign b29d94 = hlock2 & b29d92 | !hlock2 & b29d93;
assign ab059b = hlock0_p & v84563c | !hlock0_p & !b2997c;
assign af3498 = hmaster1_p & af3497 | !hmaster1_p & d40d60;
assign ab0b6e = hmaster0_p & ab0b5a | !hmaster0_p & ab0b6d;
assign a5ea07 = hlock2 & a5f1a2 | !hlock2 & a5ea06;
assign af3c3f = hready_p & af3c3a | !hready_p & af3c3e;
assign ab0c5d = hbusreq0_p & c3bd5f | !hbusreq0_p & v84565a;
assign d40d79 = hlock3_p & d40d78 | !hlock3_p & d40d5b;
assign b26693 = hmastlock_p & b26692 | !hmastlock_p & !v84563c;
assign a5ebec = hready_p & a5eba3 | !hready_p & a5ebeb;
assign a5fb02 = hbusreq3 & a5fafd | !hbusreq3 & v84563c;
assign a5ea00 = hbusreq2_p & a5e9ff | !hbusreq2_p & a5f199;
assign a5f28d = hgrant3_p & a5f95f | !hgrant3_p & a5f28c;
assign ab0582 = hgrant2_p & ab0580 | !hgrant2_p & ab0581;
assign a5fc6d = locked_p & v84563c | !locked_p & a5fc6c;
assign b29ce5 = hlock0_p & b29ce4 | !hlock0_p & !deadb2;
assign a5ee47 = hbusreq1 & a5ee46 | !hbusreq1 & v84563c;
assign a5efa7 = hlock0_p & a60141 | !hlock0_p & a5ee66;
assign b29998 = hmaster1_p & b29997 | !hmaster1_p & b29981;
assign c3bd4d = hlock2_p & c3bd4c | !hlock2_p & !cea887;
assign af348c = hbusreq2_p & af348b | !hbusreq2_p & d40d51;
assign deacf4 = start_p & deac4a | !start_p & deacf3;
assign ab0cf2 = hgrant2_p & ab0be2 | !hgrant2_p & ab0ca2;
assign b26752 = hmaster0_p & b2674b | !hmaster0_p & !b26751;
assign a5fc23 = hlock0_p & a5fc22 | !hlock0_p & a5fb91;
assign a5ee04 = hready_p & a5f3de | !hready_p & a5ee03;
assign cea271 = hbusreq1_p & deadb9 | !hbusreq1_p & !v84563c;
assign b29e9b = hgrant2_p & b29e99 | !hgrant2_p & b29e9a;
assign cea0c1 = hbusreq3 & cea0be | !hbusreq3 & cea0c0;
assign a5f4c9 = hgrant1_p & a5f4c8 | !hgrant1_p & a5f4c7;
assign a5fbee = hmastlock_p & a5fbed | !hmastlock_p & v84563c;
assign c3bcbe = decide_p & c3bcbd | !decide_p & !v845660;
assign b29b0b = hgrant3_p & b29a9f | !hgrant3_p & b29b0a;
assign adaf15 = hmaster1_p & adaf00 | !hmaster1_p & v84563c;
assign cea37a = hready & cea151 | !hready & cea376;
assign deae26 = hbusreq3 & deae20 | !hbusreq3 & deae25;
assign b266ef = hlock1_p & v84563c | !hlock1_p & b266ee;
assign cea278 = hbusreq3 & cea25b | !hbusreq3 & cea277;
assign c3b64c = hbusreq2_p & c3b64b | !hbusreq2_p & c3b64a;
assign a5f089 = hlock0_p & a5f726 | !hlock0_p & v84563c;
assign a60169 = hlock1_p & a60168 | !hlock1_p & v84563c;
assign ab06be = hlock0_p & ab06bb | !hlock0_p & !ab06bd;
assign deada7 = start_p & v845652 | !start_p & !deada6;
assign b26706 = hmaster0_p & b26702 | !hmaster0_p & b26705;
assign a5fbc5 = hgrant2_p & a5fbc4 | !hgrant2_p & v84563c;
assign b29a55 = hmaster1_p & b29a54 | !hmaster1_p & v84563c;
assign a5ee75 = hlock2 & a5f3ba | !hlock2 & a5ee74;
assign b29e6f = hmaster1_p & b29e6c | !hmaster1_p & !b29e6e;
assign a5f080 = hbusreq2 & a5f07e | !hbusreq2 & a5f07f;
assign c3b7ee = hmaster0_p & c3b7e1 | !hmaster0_p & c3b7ed;
assign a5f937 = hgrant1_p & v84563c | !hgrant1_p & a5f936;
assign a5f3b1 = hbusreq2 & a5f36b | !hbusreq2 & a5f3b0;
assign cea3cc = hlock1_p & v84563c | !hlock1_p & !cea255;
assign ab0539 = hbusreq1_p & v84563c | !hbusreq1_p & ab0538;
assign b299e6 = decide_p & b299e5 | !decide_p & b29e57;
assign af3c5a = hlock2_p & af3c59 | !hlock2_p & af3c58;
assign b29efc = hlock2 & deacb7 | !hlock2 & b29efb;
assign ab0af4 = hlock2 & ab0af2 | !hlock2 & ab0af3;
assign ce9e25 = hmaster0_p & ce9e24 | !hmaster0_p & ce9d2e;
assign af3c20 = hgrant2_p & af3c1a | !hgrant2_p & af3c1f;
assign b26725 = hlock2_p & b266a4 | !hlock2_p & !b266a2;
assign a5f930 = hbusreq1_p & a5fb8b | !hbusreq1_p & a60168;
assign cea2b5 = hlock3_p & cea29c | !hlock3_p & cea2b4;
assign ab0cf0 = hgrant2_p & ab0be2 | !hgrant2_p & ab0cef;
assign dea726 = hlock2_p & dea724 | !hlock2_p & !dea725;
assign af35b0 = hmaster1_p & af352c | !hmaster1_p & af358b;
assign ab067c = hbusreq3 & ab067b | !hbusreq3 & v845660;
assign a5fb33 = hbusreq2 & a5fb31 | !hbusreq2 & a5fb32;
assign deac4f = hburst1 & deac4e | !hburst1 & v84563c;
assign a5fbfa = hlock1_p & adaee9 | !hlock1_p & a5fbf9;
assign dead03 = hmaster0_p & deace8 | !hmaster0_p & dead02;
assign ce9d57 = hmaster1_p & ce9d4e | !hmaster1_p & cea178;
assign a5ea47 = hlock2_p & a5ea41 | !hlock2_p & a5ea46;
assign b29ebf = hlock0_p & dead7f | !hlock0_p & !b29ebe;
assign a5f83b = hlock1_p & a5f837 | !hlock1_p & a5f83a;
assign a5fc7b = stateA1_p & d615cf | !stateA1_p & a5fc75;
assign b2671a = hbusreq2_p & b26719 | !hbusreq2_p & b26717;
assign a5f6f9 = hlock2 & a5fc44 | !hlock2 & a5f6f8;
assign a5f2df = hready_p & a5f29f | !hready_p & a5f2de;
assign c3b799 = hlock2_p & c3b797 | !hlock2_p & !c3b798;
assign ab0692 = hlock0_p & b29f10 | !hlock0_p & !b29f1f;
assign a5f375 = hlock1_p & a5fc84 | !hlock1_p & !a5f374;
assign b29d0d = hlock0_p & deadde | !hlock0_p & !v84563c;
assign b26781 = hmaster1_p & b266ae | !hmaster1_p & b2675f;
assign a5f4f0 = hready & v84563c | !hready & a5f4ef;
assign ab06f5 = hbusreq2_p & ab06f4 | !hbusreq2_p & ab06f3;
assign a5f1f5 = hlock0_p & a5f1f4 | !hlock0_p & a5f9a3;
assign a5ef6f = hbusreq2_p & a5f593 | !hbusreq2_p & a5ef6e;
assign a5f290 = locked_p & v84563c | !locked_p & a5f28f;
assign a5f20f = hbusreq0 & a5f20c | !hbusreq0 & !a5f20e;
assign b29cec = hbusreq2_p & b29ceb | !hbusreq2_p & c3bc21;
assign a5f3cb = hbusreq1 & a5f3ca | !hbusreq1 & !v84563c;
assign ab0ca7 = hbusreq2_p & ab0c83 | !hbusreq2_p & dead2e;
assign ab0bb2 = hbusreq3 & ab0ba2 | !hbusreq3 & cea15a;
assign a5efda = hbusreq3 & a5efd7 | !hbusreq3 & a5efd9;
assign ce9cde = hbusreq3_p & ce9cdd | !hbusreq3_p & cea1a8;
assign a5fcc7 = hready & a5fcc5 | !hready & a5fcc6;
assign a5f787 = hready & a5f783 | !hready & a5f786;
assign c3bd93 = hmaster0_p & c3bd89 | !hmaster0_p & c3bd92;
assign c3b751 = hlock2_p & c3b637 | !hlock2_p & c3b635;
assign b266fc = hlock2_p & b266fa | !hlock2_p & b266fb;
assign c3b814 = hlock0_p & c3be00 | !hlock0_p & v845660;
assign ab06d1 = hlock0_p & b29f79 | !hlock0_p & !ab06bd;
assign c3b61f = hgrant3_p & c3bdf7 | !hgrant3_p & !c3b61e;
assign a5fa28 = hbusreq2_p & a5fa27 | !hbusreq2_p & v84563c;
assign a5ea1f = hbusreq0_p & a5fcd2 | !hbusreq0_p & v84563c;
assign b29966 = hready & c3b6be | !hready & v84563c;
assign b2674f = hbusreq2_p & b266b3 | !hbusreq2_p & !b266bc;
assign af34d6 = hbusreq2_p & af34d5 | !hbusreq2_p & af3c4c;
assign af3561 = hgrant1_p & af352c | !hgrant1_p & af3560;
assign c3bd44 = hbusreq2_p & c3bd24 | !hbusreq2_p & deac1e;
assign adaf17 = decide_p & adaed5 | !decide_p & adaf16;
assign ab0b36 = hmaster1_p & v84563c | !hmaster1_p & ab0b35;
assign ab06f2 = hbusreq2_p & ab0674 | !hbusreq2_p & b29a4d;
assign c3bc7b = locked_p & c3bc7a | !locked_p & dead0c;
assign cea2e9 = locked_p & cea2e8 | !locked_p & b26697;
assign v970454 = hgrant3_p & v970430 | !hgrant3_p & v970453;
assign b29d23 = hgrant2_p & b29d1f | !hgrant2_p & b29d22;
assign a5fc14 = hlock0_p & a5fc11 | !hlock0_p & !a5fc13;
assign af3486 = hbusreq2_p & af3c81 | !hbusreq2_p & af3c80;
assign dead15 = hlock2_p & dead14 | !hlock2_p & deace9;
assign b29ff0 = hmaster1_p & b29e5c | !hmaster1_p & b29edd;
assign c3bc6a = hmaster1_p & c3bc5f | !hmaster1_p & c3bc69;
assign deadf0 = hbusreq2_p & deadef | !hbusreq2_p & !v84563c;
assign cea32a = hmaster1_p & cea31e | !hmaster1_p & cea329;
assign cea44a = locked_p & deae59 | !locked_p & !cea38d;
assign deae63 = hbusreq3 & deae5e | !hbusreq3 & deae62;
assign a5ee2e = hbusreq1 & a5ee2c | !hbusreq1 & a5ee2d;
assign ab05e3 = hlock0_p & b29832 | !hlock0_p & v8c6711;
assign a5ee89 = hbusreq2_p & a5ee88 | !hbusreq2_p & a5ee87;
assign a5fbd8 = hbusreq1 & a5fbd7 | !hbusreq1 & !a5fba2;
assign dead92 = hbusreq1_p & v84563c | !hbusreq1_p & deacdf;
assign b299f1 = hmaster1_p & b29f75 | !hmaster1_p & !b299ed;
assign a5fc97 = hmaster0_p & a5fc6f | !hmaster0_p & a5fc96;
assign a5ea28 = hbusreq0_p & a5fccc | !hbusreq0_p & v84563c;
assign b29a3d = hlock2_p & v84563c | !hlock2_p & !b29a3c;
assign ab0b95 = hlock0_p & v84563c | !hlock0_p & b266a8;
assign a5ef7c = hlock2 & a5ef7b | !hlock2 & a5f36e;
assign a5f13a = hbusreq2_p & a5f123 | !hbusreq2_p & a5f109;
assign a5ee13 = locked_p & a5f3a0 | !locked_p & a5f38f;
assign ab0c8d = hlock2 & ab0c8a | !hlock2 & ab0c8c;
assign a5fd0f = hbusreq0_p & a5fccb | !hbusreq0_p & a5fcce;
assign c3b808 = hbusreq2_p & c3b807 | !hbusreq2_p & !c3b7ad;
assign a5f707 = hbusreq1_p & v970408 | !hbusreq1_p & !a5fbab;
assign a5f037 = hgrant3_p & a5f02d | !hgrant3_p & a5f036;
assign ab0626 = hlock2_p & ab056a | !hlock2_p & ab0563;
assign a5f8d2 = hmastlock_p & a60196 | !hmastlock_p & !v84563c;
assign cea1ae = start_p & cea1aa | !start_p & !cea1ad;
assign b29fad = hbusreq2_p & b29fac | !hbusreq2_p & v84563c;
assign a5f068 = hlock0_p & a5f065 | !hlock0_p & a5f067;
assign a60140 = hready & v84563c | !hready & v845646;
assign ab0c14 = hlock0_p & v84563c | !hlock0_p & ab0c13;
assign dea6d9 = hmaster0_p & dea6d8 | !hmaster0_p & !v84563c;
assign cea433 = hlock1_p & deac52 | !hlock1_p & !cea408;
assign c3b6b0 = hlock0_p & c3b6ae | !hlock0_p & !c3b6af;
assign a5f36e = hready & v84563c | !hready & !v845648;
assign deae6e = hmaster0_p & deae64 | !hmaster0_p & deae6d;
assign b29a89 = hgrant2_p & b29a7e | !hgrant2_p & b29a88;
assign ab0ad0 = decide_p & ab0acf | !decide_p & v84563c;
assign a5f8d3 = hbusreq1_p & a5f8d2 | !hbusreq1_p & !a60177;
assign ab0ad1 = hlock0_p & v84563c | !hlock0_p & v84565a;
assign a5fce1 = hmastlock_p & a5fce0 | !hmastlock_p & !v84563c;
assign ce9dbb = decide_p & ce9dba | !decide_p & v84563c;
assign a5f99c = hlock2_p & a5f99b | !hlock2_p & v84563c;
assign ab05ec = decide_p & ab05eb | !decide_p & v84563c;
assign a5f40a = hlock1_p & deac52 | !hlock1_p & a5f409;
assign b29a96 = hlock2_p & b29d2e | !hlock2_p & !b29a7c;
assign a5efb3 = hbusreq2_p & a5efad | !hbusreq2_p & a5efb2;
assign cea41b = hready & deae90 | !hready & cea29f;
assign a5fce8 = hbusreq0 & a5fcdb | !hbusreq0 & !a5fce7;
assign b29a45 = hbusreq3 & b29d5a | !hbusreq3 & v84563c;
assign b29d25 = hmaster0_p & b29cdb | !hmaster0_p & !b29d24;
assign c3bbf9 = hlock1_p & v84563c | !hlock1_p & !c3bbf8;
assign b29b27 = hmaster0_p & b29b25 | !hmaster0_p & b29b26;
assign deacd5 = hbusreq2_p & deacd2 | !hbusreq2_p & deacbe;
assign c3b723 = hbusreq3 & c3b718 | !hbusreq3 & c3b722;
assign ab05bc = hmaster1_p & ab0589 | !hmaster1_p & dead2e;
assign a81cf4 = hmaster1_p & v84563c | !hmaster1_p & a81cf3;
assign c3bbd5 = hlock2_p & c3bbd4 | !hlock2_p & !c3bbd3;
assign b29d34 = hready & deacbe | !hready & v84563c;
assign a5fa65 = hready & a5fa62 | !hready & a5fa64;
assign cea404 = hlock1_p & v84565a | !hlock1_p & !v845646;
assign a5f02c = decide_p & a5f02b | !decide_p & v84563c;
assign ab0c71 = hbusreq2_p & ab0bd6 | !hbusreq2_p & ab0b3b;
assign b29f98 = hgrant2_p & c3bcfb | !hgrant2_p & !b29f97;
assign a5f8e9 = hlock1_p & v84563c | !hlock1_p & a5f8e8;
assign a5ee62 = hlock2 & a5f3a1 | !hlock2 & a5ee39;
assign af356c = hmaster1_p & af356b | !hmaster1_p & af3566;
assign ce9cd0 = hmaster1_p & cea879 | !hmaster1_p & !cea1a1;
assign a5f534 = hlock1_p & a5fa1c | !hlock1_p & a5f533;
assign a5fabc = hbusreq0 & a5fa9e | !hbusreq0 & !a5fabb;
assign a5fd25 = hlock2 & a5fd24 | !hlock2 & !v84563c;
assign a5f540 = hready & v84563c | !hready & !a5f53f;
assign b29fc6 = hgrant2_p & dead3e | !hgrant2_p & !b29fc5;
assign a5fcff = hready & a5fcfd | !hready & a5fcfe;
assign dead2b = hgrant0_p & dead03 | !hgrant0_p & dead2a;
assign cea29b = hmaster1_p & cea1a3 | !hmaster1_p & cea29a;
assign deae3d = hmaster0_p & deae39 | !hmaster0_p & deae3c;
assign a5f23a = hbusreq2 & a5f238 | !hbusreq2 & a5f239;
assign deae32 = hlock0_p & deae31 | !hlock0_p & !v84563c;
assign ab05df = hlock0_p & b298a4 | !hlock0_p & !ab05de;
assign cea276 = hlock2_p & cea275 | !hlock2_p & v84563c;
assign a5fc5b = locked_p & a5fc5a | !locked_p & v84563c;
assign a5eddb = hlock0_p & a5edda | !hlock0_p & a5f576;
assign cea3ab = hbusreq3 & cea3aa | !hbusreq3 & !cea3a7;
assign b29ffa = decide_p & b29ff9 | !decide_p & v84563c;
assign a5ef9b = hbusreq2_p & a5ef9a | !hbusreq2_p & a5ee0c;
assign a5ea3c = hlock2 & v84563c | !hlock2 & v845641;
assign a5ef8a = hbusreq2_p & a5edd6 | !hbusreq2_p & a5ef89;
assign deae6b = hbusreq2_p & deae66 | !hbusreq2_p & deae65;
assign c06d34 = stateG3_1_p & v845670 | !stateG3_1_p & !v84563c;
assign dea6d2 = hbusreq2_p & dea6d1 | !hbusreq2_p & !deadba;
assign a5edfb = locked_p & v845641 | !locked_p & a5edfa;
assign a5ee82 = hmaster1_p & a5ee81 | !hmaster1_p & v84563c;
assign dea731 = hbusreq3 & dea730 | !hbusreq3 & !v84563c;
assign a5f8b5 = hbusreq1_p & deac52 | !hbusreq1_p & !deaca1;
assign c3b6ae = hready & c3b6a6 | !hready & c3bd5d;
assign a5fb94 = hready & a5fb8a | !hready & !a5fb8c;
assign c3bdfc = hbusreq2_p & c3bdfb | !hbusreq2_p & c3bc5c;
assign a5f45c = hlock0_p & a5f440 | !hlock0_p & !a5f45b;
assign a5fcaa = hready & b2672b | !hready & a5fca9;
assign a5f41c = hlock1_p & v84563c | !hlock1_p & ab055c;
assign b29fb8 = hlock2 & b29fb6 | !hlock2 & b29fb7;
assign c98b95 = hgrant1_p & v84563c | !hgrant1_p & v845646;
assign ce9d21 = hbusreq3 & ce9d1f | !hbusreq3 & ce9d20;
assign ab05b4 = hlock0_p & v84563c | !hlock0_p & !ab05b3;
assign a5ee5a = hlock1_p & a5fbe1 | !hlock1_p & a5ee52;
assign ab06fd = hlock0_p & c3bd8d | !hlock0_p & v845660;
assign a5f8e2 = hbusreq1_p & a5f8dd | !hbusreq1_p & !a5fbab;
assign af34b8 = hlock1_p & d40d33 | !hlock1_p & !af34b7;
assign dea74a = hmaster0_p & dea749 | !hmaster0_p & !v84563c;
assign c3bd9f = hgrant2_p & c3bc6d | !hgrant2_p & c3bd9e;
assign v8567b4 = hmaster0_p & v877992 | !hmaster0_p & v845646;
assign c3bbd1 = hlock1_p & v84563c | !hlock1_p & !deac56;
assign a5ef50 = hgrant1_p & b8acda | !hgrant1_p & v84563c;
assign af3c2e = hlock0_p & af3c2c | !hlock0_p & af3c2d;
assign b29d61 = hbusreq3 & b29d60 | !hbusreq3 & c3bceb;
assign b29f6b = hbusreq2_p & b29f69 | !hbusreq2_p & v84563c;
assign cea42f = hready & cea42e | !hready & cea3bf;
assign cea480 = hgrant1_p & cea47f | !hgrant1_p & deae7f;
assign deac7a = hlock1_p & v84563c | !hlock1_p & !v84565a;
assign c3bd7c = hlock2_p & c3bd7b | !hlock2_p & c3bc3c;
assign a5f045 = hgrant3_p & a5f03d | !hgrant3_p & a5f044;
assign a5fbf7 = hgrant2_p & a5fbd6 | !hgrant2_p & a5fbf6;
assign b29ece = hlock2_p & b29ecd | !hlock2_p & v845660;
assign c3bda9 = hlock0_p & c3bce6 | !hlock0_p & !c3bce5;
assign b29a44 = hmaster1_p & b29a3f | !hmaster1_p & b29a43;
assign a5f332 = hbusreq0 & a5f330 | !hbusreq0 & !a5f331;
assign a5f549 = hlock0_p & a5fa6c | !hlock0_p & a5f36e;
assign cea465 = hbusreq2_p & cea464 | !hbusreq2_p & cea463;
assign a5fb84 = hbusreq2_p & v84563c | !hbusreq2_p & a5fb83;
assign ab0c96 = hlock1_p & b2a020 | !hlock1_p & !v84563c;
assign a5f2eb = hbusreq2_p & a5f2ea | !hbusreq2_p & a60142;
assign deae1b = decide_p & deae1a | !decide_p & v84563c;
assign bdb585 = hlock0_p & bdb584 | !hlock0_p & v84565a;
assign dead66 = hmaster1_p & dead63 | !hmaster1_p & dead65;
assign dea6cb = hlock0_p & dea6ca | !hlock0_p & !deada8;
assign ab0cae = hlock0_p & ab0cad | !hlock0_p & ab0c89;
assign b29f94 = hmaster0_p & b29f8c | !hmaster0_p & b29f93;
assign ab0bfa = hready & dead6e | !hready & !v84563c;
assign a5fc3b = hbusreq3 & a5fc31 | !hbusreq3 & a5fc3a;
assign a5f07c = hbusreq0 & a5f07b | !hbusreq0 & !v84563c;
assign ab0c1c = hlock0_p & v84563c | !hlock0_p & !v845660;
assign a5f325 = hlock2_p & a5f324 | !hlock2_p & v84563c;
assign a5f08c = hbusreq2_p & a5f08a | !hbusreq2_p & a5f08b;
assign a5eb9a = hmaster0_p & a5eb99 | !hmaster0_p & a5ea6d;
assign a5f572 = hgrant1_p & b29928 | !hgrant1_p & b29923;
assign b29a9a = hgrant2_p & b29a97 | !hgrant2_p & b29a99;
assign dead6b = hbusreq3_p & dead52 | !hbusreq3_p & dead6a;
assign adaec4 = hmastlock_p & adaec3 | !hmastlock_p & v84563c;
assign ce9df1 = hbusreq0_p & cea17a | !hbusreq0_p & !cea18d;
assign a5eae5 = hlock0_p & a5f248 | !hlock0_p & !a5eae4;
assign b29976 = hlock3_p & b29958 | !hlock3_p & b29975;
assign b29fa8 = hmaster1_p & b29d64 | !hmaster1_p & b29fa7;
assign a5f35b = hgrant2_p & v84563c | !hgrant2_p & a5f344;
assign b29b35 = hgrant3_p & b29b1b | !hgrant3_p & b29b34;
assign a5f11f = hlock1_p & a5f11b | !hlock1_p & a5f11e;
assign c3bda2 = hgrant2_p & c3bc6d | !hgrant2_p & c3bda1;
assign a5f8de = stateA1_p & v84563c | !stateA1_p & a81ca6;
assign ab05c5 = hlock0_p & v84563c | !hlock0_p & ab0598;
assign adaf0f = decide_p & adaefd | !decide_p & adaf0e;
assign ab0617 = locked_p & deae59 | !locked_p & !ab0610;
assign b29ea5 = hready & deacf7 | !hready & v84563c;
assign adaecf = hbusreq2_p & adaece | !hbusreq2_p & v84563c;
assign ab0ca1 = hmaster1_p & ab0c94 | !hmaster1_p & ab0ca0;
assign a5fd12 = hlock0_p & v845660 | !hlock0_p & a5fd11;
assign c3bdf9 = locked_p & v84563c | !locked_p & c3bdf8;
assign a5fb65 = hmaster1_p & a5fb37 | !hmaster1_p & a5fb64;
assign a5f705 = hbusreq1_p & a5f704 | !hbusreq1_p & !a5fc84;
assign d40d7b = hmastlock_p & d40d7a | !hmastlock_p & v84563c;
assign cea190 = hbusreq2_p & cea15b | !hbusreq2_p & cea18f;
assign b29f03 = start_p & cea1aa | !start_p & !v84563c;
assign ab06ef = hmaster0_p & ab06e5 | !hmaster0_p & ab06ee;
assign c3bdb9 = hburst1 & v84566c | !hburst1 & !v84563c;
assign b29d67 = hlock0_p & b29d66 | !hlock0_p & !v84563c;
assign dea6c5 = hmaster0_p & dea6c1 | !hmaster0_p & dea6c4;
assign cea407 = stateG10_1_p & deaca1 | !stateG10_1_p & cea3bc;
assign c3bc6b = hmaster0_p & c3bc57 | !hmaster0_p & c3bc6a;
assign b298ad = hbusreq2_p & b298ac | !hbusreq2_p & v84563c;
assign a5f543 = hbusreq1 & a5f493 | !hbusreq1 & v84565a;
assign c3b732 = hbusreq2_p & c3b64b | !hbusreq2_p & c3b731;
assign c3b81b = hbusreq2_p & c3b81a | !hbusreq2_p & !c3b7b0;
assign bdb59c = hready_p & bdb583 | !hready_p & bdb59b;
assign a5fb10 = stateG10_1_p & v84563c | !stateG10_1_p & a60167;
assign a5f58a = hmaster1_p & a5f54e | !hmaster1_p & a5f589;
assign ab054c = hlock0_p & ab054b | !hlock0_p & !b2992b;
assign cea181 = decide_p & cea180 | !decide_p & a57859;
assign a5fbde = locked_p & a5fbdb | !locked_p & a5fbdd;
assign a5fc63 = hgrant2_p & a5fc62 | !hgrant2_p & v84563c;
assign a5ead0 = hready & a60168 | !hready & a5f786;
assign a5eef2 = hbusreq2_p & a5eef1 | !hbusreq2_p & !a5eef0;
assign deac54 = stateG10_1_p & v84565a | !stateG10_1_p & deac53;
assign c3bd38 = hmastlock_p & deacb3 | !hmastlock_p & !v84563c;
assign b29b11 = hmaster0_p & b29b0f | !hmaster0_p & b29b10;
assign af352e = hbusreq1_p & v84563c | !hbusreq1_p & af352c;
assign a5f475 = hlock2_p & a5f45c | !hlock2_p & !a5f474;
assign ab0614 = hbusreq2_p & ab060f | !hbusreq2_p & ab0613;
assign b2998e = hlock2 & b298ab | !hlock2 & b2998d;
assign ab074b = hmaster0_p & ab0749 | !hmaster0_p & ab074a;
assign a5f990 = hlock0_p & a5f98f | !hlock0_p & a5fad4;
assign a5eef4 = hbusreq2_p & a5eede | !hbusreq2_p & a5eedb;
assign c3bc90 = hbusreq0_p & b266a8 | !hbusreq0_p & c3bc8b;
assign af3c5c = hmaster1_p & af3c53 | !hmaster1_p & af3c5b;
assign a5f1c4 = hbusreq2_p & a5f1c3 | !hbusreq2_p & v84563c;
assign ce9d59 = hgrant0_p & v84563c | !hgrant0_p & ce9d58;
assign a5ee38 = hready & v84563c | !hready & !deae59;
assign a5fbc0 = locked_p & v84563c | !locked_p & v845641;
assign a5f961 = hlock2_p & a5f960 | !hlock2_p & v84563c;
assign b2678b = decide_p & b2678a | !decide_p & b26783;
assign cea3a3 = hmaster1_p & cea3a2 | !hmaster1_p & v84563c;
assign ab0c85 = hlock0_p & v845660 | !hlock0_p & c3bce5;
assign a5f712 = hmastlock_p & a5f711 | !hmastlock_p & v84563c;
assign a5fa26 = hlock2 & v84563c | !hlock2 & a5fa25;
assign b29f19 = hmastlock_p & b29f18 | !hmastlock_p & !v84563c;
assign ab0ace = hbusreq3 & ab0acd | !hbusreq3 & v84563c;
assign a5eb54 = decide_p & a5eb4e | !decide_p & !a5eb53;
assign deac4d = stateA1_p & v84563c | !stateA1_p & deac4c;
assign a5f291 = hlock0_p & a5f290 | !hlock0_p & v84563c;
assign c3b6fa = locked_p & c3b6f9 | !locked_p & !c3b625;
assign a5f09c = hlock0_p & a5f727 | !hlock0_p & v84563c;
assign c3b825 = locked_p & c3b824 | !locked_p & !c3bcdb;
assign a5fc71 = locked_p & v84563c | !locked_p & !a5fc70;
assign c3bc08 = hgrant1_p & c3bbd2 | !hgrant1_p & c3bbf7;
assign a5f2fc = hmaster0_p & a5f2fb | !hmaster0_p & a5f1bf;
assign cea0b7 = hlock1_p & v84563c | !hlock1_p & !cea0b6;
assign a5f459 = hlock1_p & a5fa1d | !hlock1_p & a5f458;
assign a9b9e1 = hgrant0_p & a9b9d8 | !hgrant0_p & a9b9e0;
assign deae18 = hmaster0_p & deae16 | !hmaster0_p & deae17;
assign c3b892 = hgrant2_p & c3b808 | !hgrant2_p & c3b891;
assign a5f2e6 = hready & v84563c | !hready & !deacec;
assign cea43f = hmaster0_p & cea428 | !hmaster0_p & cea43e;
assign ab0516 = hlock2_p & b298a4 | !hlock2_p & ab0515;
assign ab072f = decide_p & ab072e | !decide_p & !v845662;
assign b2999c = hready & c3b6f8 | !hready & !v84563c;
assign b2a005 = hbusreq2_p & b2a004 | !hbusreq2_p & v84563c;
assign ab0686 = hmaster1_p & ab0685 | !hmaster1_p & v84563c;
assign a5f14d = hlock2_p & a5f145 | !hlock2_p & a5f14c;
assign b299cf = hbusreq3 & b299ce | !hbusreq3 & b2995c;
assign deae05 = locked_p & deae04 | !locked_p & !dead8a;
assign cea148 = hlock0_p & b2669d | !hlock0_p & v84563c;
assign b29e71 = decide_p & b29e70 | !decide_p & v84563c;
assign a5f495 = hready & a5f492 | !hready & a5f494;
assign c3bc17 = hlock2_p & c3bc15 | !hlock2_p & !c3bc16;
assign ab0af5 = hlock2_p & ab0af1 | !hlock2_p & ab0af4;
assign a5f556 = hlock1_p & a60172 | !hlock1_p & a5f555;
assign ce9dc8 = hlock0_p & cea2ae | !hlock0_p & ce9dc7;
assign dead85 = hbusreq3 & v845660 | !hbusreq3 & dead84;
assign b29a58 = decide_p & b29a57 | !decide_p & v84563c;
assign b29a8b = hmaster0_p & b29a6f | !hmaster0_p & !b29a8a;
assign a5f3d2 = locked_p & v84563c | !locked_p & a5f3c8;
assign cea2e7 = hlock1_p & v84563c | !hlock1_p & cea2e6;
assign a5ee43 = hbusreq1 & a5fb89 | !hbusreq1 & v84563c;
assign a5eeb5 = hlock3_p & a5ee7e | !hlock3_p & a5eeb4;
assign b29f45 = hbusreq2_p & b29f43 | !hbusreq2_p & v84563c;
assign a5ea19 = hbusreq0 & a5ea18 | !hbusreq0 & a5ea0f;
assign ab0c70 = hmaster1_p & ab0c6f | !hmaster1_p & ab0c47;
assign ab05a8 = hlock2 & ab0521 | !hlock2 & ab05a7;
assign a5f9a4 = hlock0_p & a5f9a1 | !hlock0_p & a5f9a3;
assign dead41 = locked_p & dead40 | !locked_p & v84563c;
assign a5f470 = hlock1_p & a5f837 | !hlock1_p & a5f458;
assign b29b61 = jx2_p & b2a01d | !jx2_p & b29b60;
assign cea1c6 = hmaster1_p & cea1c3 | !hmaster1_p & cea1c5;
assign a5f52a = hlock1_p & a60177 | !hlock1_p & !a5f4cc;
assign c3b80e = hmaster1_p & c3b806 | !hmaster1_p & c3b80d;
assign a5fb31 = hlock2 & a5fa5b | !hlock2 & a5fb30;
assign dea6dd = hgrant3_p & deaead | !hgrant3_p & !dea6dc;
assign a5ea88 = hbusreq2_p & a5f089 | !hbusreq2_p & a5ea60;
assign b29d58 = hlock0_p & b266a8 | !hlock0_p & v84563c;
assign cea4aa = hbusreq2_p & cea49b | !hbusreq2_p & cea49a;
assign a5ef31 = decide_p & a5eefa | !decide_p & a5ef30;
assign c3bc99 = hlock0_p & b26720 | !hlock0_p & c3bc90;
assign ab0b58 = hbusreq2_p & ab0b57 | !hbusreq2_p & ab0b56;
assign b29b0d = hbusreq2_p & b29b0c | !hbusreq2_p & v84563c;
assign dea748 = hgrant2_p & dea744 | !hgrant2_p & dea747;
assign a5f753 = hbusreq2 & a5fcbc | !hbusreq2 & v84563c;
assign b29984 = locked_p & b29983 | !locked_p & !v84563c;
assign c3b8b4 = hmaster0_p & c3b8b3 | !hmaster0_p & c3b7ed;
assign a5fc07 = hlock2 & a5fbff | !hlock2 & a5fc06;
assign c3b693 = hgrant1_p & c3b692 | !hgrant1_p & deae74;
assign deae24 = hlock2_p & deae23 | !hlock2_p & !deadba;
assign d40d73 = hgrant2_p & d40d72 | !hgrant2_p & v84563c;
assign b29cd9 = hbusreq3 & b29cd7 | !hbusreq3 & b29cd8;
assign af34ea = hmaster1_p & af34e9 | !hmaster1_p & af3c64;
assign a5efe1 = hbusreq2_p & a5f547 | !hbusreq2_p & a5efe0;
assign a5ef7d = hlock0_p & a5edcc | !hlock0_p & a5ef6b;
assign b29a53 = hbusreq2_p & b29a52 | !hbusreq2_p & v84563c;
assign af3c64 = hlock0_p & af3c5e | !hlock0_p & af3c62;
assign c3bd65 = hbusreq2_p & c3bd63 | !hbusreq2_p & c3bc20;
assign dead1a = hlock0_p & dead19 | !hlock0_p & deacfb;
assign a5ee8b = hbusreq1 & a5ee8a | !hbusreq1 & !v84563c;
assign b266f2 = hgrant2_p & b266ed | !hgrant2_p & b266f1;
assign a5ebea = hgrant0_p & v84563c | !hgrant0_p & a5ebe9;
assign c3be06 = hmaster0_p & c3be05 | !hmaster0_p & c3bda3;
assign af3578 = hready_p & af3539 | !hready_p & af3577;
assign ce9d50 = hmaster0_p & ce9d4b | !hmaster0_p & ce9d4f;
assign b29f56 = hlock2 & b29f52 | !hlock2 & b29f55;
assign c3b67c = hready & c3b67b | !hready & c3bd2c;
assign c3b64e = hmaster1_p & c3b64d | !hmaster1_p & v84563c;
assign c3b755 = hmaster0_p & c3b754 | !hmaster0_p & c3b6f2;
assign b29ae5 = hbusreq2_p & b29ae4 | !hbusreq2_p & !b29ae3;
assign deac7c = hbusreq2_p & deac72 | !hbusreq2_p & !deac7b;
assign a5f03e = hbusreq2_p & a5f01c | !hbusreq2_p & v84563c;
assign c3bc63 = locked_p & c3bc62 | !locked_p & b2671f;
assign deaea3 = hlock2_p & deaea2 | !hlock2_p & !v84563c;
assign b29d03 = hlock2_p & b29d02 | !hlock2_p & b29cea;
assign b2990b = hlock2_p & v84563c | !hlock2_p & b2990a;
assign af3535 = hmaster0_p & af3530 | !hmaster0_p & af3534;
assign cea234 = hbusreq3 & cea15e | !hbusreq3 & v84563c;
assign c3bdd3 = hbusreq2_p & c3bdd2 | !hbusreq2_p & v84565a;
assign a5fcf8 = hlock1_p & v84563c | !hlock1_p & a5fcf7;
assign cea197 = hlock0_p & cea196 | !hlock0_p & !v84563c;
assign a5f288 = hmaster1_p & v84563c | !hmaster1_p & a5f287;
assign a5ea06 = hlock0_p & a5f946 | !hlock0_p & a5f1a3;
assign b29eaf = hlock0_p & b29eac | !hlock0_p & !b29eae;
assign a5ebdc = hbusreq2 & a5ea2a | !hbusreq2 & a5eb36;
assign ab0521 = hlock0_p & v84563c | !hlock0_p & !b298aa;
assign a5fc53 = hbusreq1 & a5fbd7 | !hbusreq1 & a5fc52;
assign cea362 = hmaster0_p & cea361 | !hmaster0_p & cea2f7;
assign b299a6 = hmaster0_p & b2999b | !hmaster0_p & b299a5;
assign b299eb = hbusreq3_p & b299ac | !hbusreq3_p & b299ea;
assign a5fb62 = hbusreq2_p & a5fb5f | !hbusreq2_p & a5fb5e;
assign cea85c = locked_p & v84563c | !locked_p & !v845646;
assign af348d = hgrant2_p & af348a | !hgrant2_p & af348c;
assign b29ebc = hlock0_p & b29ebb | !hlock0_p & v845660;
assign a5fbbf = hmaster0_p & a5fb7f | !hmaster0_p & a5fbbe;
assign b29f09 = hburst1 & deadb9 | !hburst1 & b29f08;
assign b29ea8 = hready & deae02 | !hready & !dead33;
assign adaee4 = hbusreq2_p & adaee3 | !hbusreq2_p & v84563c;
assign b29a4d = hlock0_p & c3bce5 | !hlock0_p & !v84563c;
assign v97044a = hgrant2_p & v970449 | !hgrant2_p & v84563c;
assign b298a1 = hlock0_p & b298a0 | !hlock0_p & v84563c;
assign a5ee59 = locked_p & a5ee58 | !locked_p & !v845641;
assign b266d5 = hbusreq2_p & b266d3 | !hbusreq2_p & b266d2;
assign a5e9cd = hgrant2_p & a5e9ae | !hgrant2_p & a5e9cc;
assign a5f409 = hgrant1_p & a5f3f5 | !hgrant1_p & a5f3f4;
assign a5efbd = hgrant2_p & a5efbc | !hgrant2_p & v84563c;
assign c3bcf4 = hbusreq2_p & c3bcf3 | !hbusreq2_p & c3bbbc;
assign ab0532 = hmaster0_p & ab0527 | !hmaster0_p & ab0531;
assign b29d8e = hbusreq2_p & b29d86 | !hbusreq2_p & b29d8d;
assign b29f36 = hbusreq3 & b29efe | !hbusreq3 & b29f35;
assign a5ebc1 = hbusreq2 & a5f198 | !hbusreq2 & a5e9c9;
assign ab0b4b = hbusreq3 & c3bc3c | !hbusreq3 & !ab0b4a;
assign deadd3 = hbusreq1_p & v84563c | !hbusreq1_p & !v84565a;
assign v97043f = locked_p & v97043e | !locked_p & v84563c;
assign b29fb2 = hbusreq1_p & deacf7 | !hbusreq1_p & v84563c;
assign b2678d = hgrant3_p & b26772 | !hgrant3_p & b2678c;
assign ab062c = hbusreq2_p & ab0626 | !hbusreq2_p & ab062b;
assign ce9d2e = hmaster1_p & ce9d2d | !hmaster1_p & cea188;
assign a5fbfd = hready & a5fbf9 | !hready & !deae02;
assign ab0c42 = hbusreq3 & ab0c35 | !hbusreq3 & ab0c41;
assign ab0529 = hlock0_p & v84563c | !hlock0_p & cea38d;
assign d40d4e = hbusreq2_p & d40d36 | !hbusreq2_p & d40d33;
assign c3bd7f = hmaster0_p & c3bd73 | !hmaster0_p & !c3bd7e;
assign c3b714 = hlock1_p & v84563c | !hlock1_p & !c3b713;
assign a5efeb = hgrant2_p & a5efe5 | !hgrant2_p & a5efea;
assign a81cd8 = hmaster0_p & a81cd3 | !hmaster0_p & a81cd7;
assign ab05cd = hbusreq2_p & ab05cc | !hbusreq2_p & ab05ac;
assign a5fc49 = hready & a5fc48 | !hready & v9703fc;
assign deaca2 = hlock1_p & deaca1 | !hlock1_p & v84563c;
assign b29d5e = hlock0_p & b29d5d | !hlock0_p & !v84563c;
assign dea753 = hmaster1_p & dea750 | !hmaster1_p & dea752;
assign b29d97 = hbusreq3 & b29d96 | !hbusreq3 & c3bcfb;
assign dead37 = hmaster1_p & dead2f | !hmaster1_p & !dead36;
assign b2997f = hlock2_p & v845660 | !hlock2_p & b2997e;
assign ab0c02 = hbusreq2_p & ab0c01 | !hbusreq2_p & ab0acb;
assign a5fc61 = hbusreq2_p & a5fc60 | !hbusreq2_p & v84563c;
assign c3b82f = hlock3_p & c3b819 | !hlock3_p & c3b82e;
assign ab0c32 = hlock0_p & v84563c | !hlock0_p & ab0c31;
assign b29826 = locked_p & b29825 | !locked_p & cea37b;
assign a5eb44 = hmaster1_p & a5eb43 | !hmaster1_p & v84563c;
assign af350d = decide_p & af350c | !decide_p & af34f9;
assign a5ee31 = hlock0_p & a5ee30 | !hlock0_p & a5ee28;
assign a5f217 = hgrant2_p & v84563c | !hgrant2_p & a5f754;
assign deacb0 = hbusreq3 & deaca2 | !hbusreq3 & !deacaf;
assign c3bde6 = hbusreq3 & c3bde5 | !hbusreq3 & c3bcfb;
assign cea395 = hlock0_p & cea38a | !hlock0_p & cea393;
assign a5f4f1 = hlock0_p & a5f36e | !hlock0_p & a5f4f0;
assign a5eb97 = hbusreq0 & a5eb96 | !hbusreq0 & a5f084;
assign jx1 = !aa0e0c;
assign ab056b = hlock0_p & ab0adc | !hlock0_p & !b29949;
assign a5f39c = hmaster1_p & a5f393 | !hmaster1_p & a5f39b;
assign c3b74a = hmaster0_p & c3b749 | !hmaster0_p & c3b6d1;
assign v97045c = hgrant3_p & v970459 | !hgrant3_p & v97045b;
assign a5eed1 = hbusreq2 & a5f3db | !hbusreq2 & v845660;
assign a5f00e = hmaster1_p & a5f00d | !hmaster1_p & v84563c;
assign a5f729 = hbusreq0_p & a5f726 | !hbusreq0_p & a5f728;
assign a5fb1c = hgrant1_p & a5fb1b | !hgrant1_p & a60186;
assign b26743 = hlock0_p & b266ae | !hlock0_p & b266a0;
assign c3bd15 = hlock1_p & v84563c | !hlock1_p & !c3bd14;
assign b29cdf = hready & deadb2 | !hready & v84563c;
assign ab06a5 = hbusreq2_p & ab06a4 | !hbusreq2_p & ab06a3;
assign a5fc8f = hmastlock_p & a5fc8e | !hmastlock_p & !v84563c;
assign c3bc0e = hbusreq2_p & c3bc05 | !hbusreq2_p & c3bc0d;
assign a5f440 = hready & a5f438 | !hready & a5f43f;
assign stateG10_3 = !b0d8fd;
assign b299a8 = hlock3_p & b2999a | !hlock3_p & b299a7;
assign b29a62 = stateG10_1_p & c3bd38 | !stateG10_1_p & c3b683;
assign b2993d = hready & b29939 | !hready & c3b694;
assign c3bc75 = hlock0_p & c3bc52 | !hlock0_p & v845660;
assign ab0ae2 = hbusreq2_p & ab0adf | !hbusreq2_p & ab0add;
assign af3588 = hgrant0_p & af357d | !hgrant0_p & af3587;
assign a5ee52 = hbusreq1_p & a5fc51 | !hbusreq1_p & v84563c;
assign ab0674 = hlock0_p & b29ec6 | !hlock0_p & v845660;
assign a5e9dc = hbusreq3 & a5e9d9 | !hbusreq3 & a5e9db;
assign a5fc56 = locked_p & a5fc55 | !locked_p & v84563c;
assign a5fcca = hmaster1_p & v84563c | !hmaster1_p & a5fcc9;
assign a5f367 = locked_p & a5f366 | !locked_p & a60140;
assign ab06e5 = hmaster1_p & ab06dd | !hmaster1_p & ab06e4;
assign c3bd6c = hbusreq2_p & c3bd6b | !hbusreq2_p & v84563c;
assign dea6e1 = hbusreq2_p & dea6e0 | !hbusreq2_p & dea6df;
assign deac10 = hlock3_p & deac0f | !hlock3_p & v84563c;
assign c3bc03 = hready & deac19 | !hready & c3bc02;
assign a5eb90 = hlock2_p & a5eb8e | !hlock2_p & a5eb8f;
assign a5edec = locked_p & a5ede8 | !locked_p & a5edeb;
assign cea8a3 = hgrant2_p & cea89f | !hgrant2_p & cea8a2;
assign a5edcc = hready & v84563c | !hready & c3b6a0;
assign b29f84 = decide_p & b29f83 | !decide_p & v84563c;
assign a5ebc9 = hgrant2_p & a5ebc3 | !hgrant2_p & a5ebc8;
assign af35a6 = hmaster1_p & af3541 | !hmaster1_p & af354c;
assign a5fb6d = hlock2_p & a5fb6c | !hlock2_p & v84563c;
assign cea444 = hlock0_p & cea38a | !hlock0_p & cea37b;
assign cea175 = hmaster1_p & cea171 | !hmaster1_p & cea174;
assign cea2f1 = locked_p & cea15f | !locked_p & !dead0a;
assign cea490 = hgrant3_p & cea442 | !hgrant3_p & cea48f;
assign deac9b = hbusreq2_p & deac89 | !hbusreq2_p & deac87;
assign a81cf8 = locked_p & a81cf7 | !locked_p & v84563c;
assign a5f15e = hbusreq2_p & a5f15d | !hbusreq2_p & a5f15c;
assign b266e1 = hlock0_p & b266dc | !hlock0_p & b266e0;
assign c3bd06 = hmaster1_p & v84563c | !hmaster1_p & c3bd05;
assign c3bca1 = hbusreq3 & c3bca0 | !hbusreq3 & !dead2e;
assign dead7a = start_p & v845652 | !start_p & c07311;
assign af34be = hbusreq2_p & af34bd | !hbusreq2_p & af34bc;
assign deace7 = hbusreq3 & deace6 | !hbusreq3 & v84563c;
assign cea2b3 = hmaster1_p & cea86e | !hmaster1_p & cea29a;
assign a5f711 = start_p & v845654 | !start_p & v84563c;
assign a5fb1f = hlock1_p & v9703fb | !hlock1_p & a5fb1e;
assign ab0cdd = hmaster0_p & ab0cd9 | !hmaster0_p & ab0cdc;
assign a6018d = hlock0_p & a60179 | !hlock0_p & a6018c;
assign a5f3a4 = hlock0_p & a5f3a3 | !hlock0_p & a5f3a1;
assign dead9c = hbusreq3 & dead9b | !hbusreq3 & !v84563c;
assign b29fd7 = hgrant1_p & b29f0b | !hgrant1_p & b29f0d;
assign ab05ae = hgrant2_p & ab05ad | !hgrant2_p & cea15a;
assign a5f516 = hready & a5f515 | !hready & !c3b6a6;
assign c3bc4e = hlock0_p & c3bc4d | !hlock0_p & !deace1;
assign af349a = decide_p & af3496 | !decide_p & af3499;
assign deace3 = locked_p & v84563c | !locked_p & deace1;
assign c3b6c2 = hbusreq2_p & c3b6c1 | !hbusreq2_p & c3b6a1;
assign a5f2d3 = hbusreq2_p & a5f949 | !hbusreq2_p & v84563c;
assign ab0c24 = hmaster1_p & ab0c1f | !hmaster1_p & ab0c23;
assign dea749 = hmaster1_p & dea748 | !hmaster1_p & !v84563c;
assign a5ef3b = hlock0_p & a5ee83 | !hlock0_p & a5ef3a;
assign deade1 = hlock2_p & deade0 | !hlock2_p & !v84563c;
assign dea787 = hbusreq2_p & deae24 | !hbusreq2_p & deae23;
assign cea0e7 = hbusreq3 & cea887 | !hbusreq3 & !deacaa;
assign cea488 = hbusreq2_p & cea484 | !hbusreq2_p & cea483;
assign ab0adf = hlock2_p & ab0add | !hlock2_p & ab0ade;
assign ab0546 = hmastlock_p & b29f0a | !hmastlock_p & c3b676;
assign af3563 = hlock0_p & af3562 | !hlock0_p & af352c;
assign a5f93f = hlock0_p & a5f93e | !hlock0_p & !v84563c;
assign deadbb = stateG10_1_p & deacb4 | !stateG10_1_p & deadba;
assign cea43d = hgrant2_p & cea43b | !hgrant2_p & cea43c;
assign af3c72 = hmaster0_p & af3c6f | !hmaster0_p & af3c71;
assign b29aad = hlock0_p & b29d79 | !hlock0_p & !b29e4d;
assign deac5d = hlock2_p & deac5c | !hlock2_p & deac5b;
assign cea89d = hlock2_p & cea89c | !hlock2_p & deacaa;
assign cea1ba = hburst0 & v84563c | !hburst0 & cea1b9;
assign a5f2f5 = locked_p & v84563c | !locked_p & a5f2f4;
assign dead0e = hlock0_p & dead0b | !hlock0_p & dead0d;
assign a5f326 = hbusreq2_p & a5f325 | !hbusreq2_p & v84563c;
assign b29b1a = decide_p & b29b19 | !decide_p & v84563c;
assign cea161 = locked_p & cea15f | !locked_p & !cea160;
assign a5fd19 = hgrant0_p & a5fceb | !hgrant0_p & a5fd18;
assign ab0d06 = hbusreq2_p & ab0d05 | !hbusreq2_p & ab0d03;
assign b29e4b = hmaster1_p & b29e48 | !hmaster1_p & b29e4a;
assign a5eaef = hbusreq2_p & a5eadd | !hbusreq2_p & a5eadb;
assign ab06af = hlock1_p & deaca0 | !hlock1_p & ab06ae;
assign a5ef5a = hlock2_p & a5ef53 | !hlock2_p & a5ef59;
assign c3bbf4 = hgrant2_p & c3bbf0 | !hgrant2_p & c3bbf3;
assign af3c4e = hlock1_p & d40d33 | !hlock1_p & af3c4d;
assign a5fb78 = hbusreq2_p & a5fb77 | !hbusreq2_p & a5fb74;
assign b29fcb = hgrant2_p & dead3e | !hgrant2_p & !b29fca;
assign cea3aa = hlock0_p & cea37b | !hlock0_p & cea3a9;
assign a5f210 = hmaster1_p & v84563c | !hmaster1_p & a5f20f;
assign a5ea83 = hlock0_p & a5ea82 | !hlock0_p & !a5ea5b;
assign a5ee69 = hbusreq2 & a5ee67 | !hbusreq2 & a5ee68;
assign a5f01f = hbusreq2_p & a5f01c | !hbusreq2_p & a5fa37;
assign a5f953 = hbusreq2_p & a5f952 | !hbusreq2_p & v84563c;
assign cea19e = hbusreq2_p & cea19a | !hbusreq2_p & cea0bf;
assign af34cc = hmaster0_p & af34c0 | !hmaster0_p & af34cb;
assign a5f0a6 = hbusreq0 & a5f0a5 | !hbusreq0 & !v84563c;
assign ab0608 = hbusreq2_p & ab0594 | !hbusreq2_p & ab0607;
assign a5f97f = start_p & a5fba3 | !start_p & a5f97e;
assign ab05d9 = hready_p & ab05d7 | !hready_p & !ab05d8;
assign b266d4 = hbusreq2_p & b266d3 | !hbusreq2_p & b266ca;
assign cea168 = hbusreq2_p & cea154 | !hbusreq2_p & v84563c;
assign a5f6ec = hready & a5fb8a | !hready & a5f6e6;
assign b29d81 = hlock0_p & deace9 | !hlock0_p & !v84563c;
assign cea33a = hgrant2_p & cea338 | !hgrant2_p & cea339;
assign bdb5aa = hgrant0_p & bdb5a4 | !hgrant0_p & bdb5a9;
assign c3bc56 = hbusreq3 & c3bc50 | !hbusreq3 & c3bc55;
assign a5f26d = hbusreq2 & a5fce7 | !hbusreq2 & !v84563c;
assign a5fab1 = hlock0_p & a5fab0 | !hlock0_p & !v84563c;
assign deadee = hlock0_p & deaded | !hlock0_p & !v84563c;
assign ab0cba = hgrant0_p & ab0cb3 | !hgrant0_p & !ab0cb9;
assign cea347 = hmaster0_p & cea346 | !hmaster0_p & cea239;
assign c3b6b9 = hmaster1_p & c3b6b8 | !hmaster1_p & !deacaa;
assign a5f0ae = hbusreq0 & a5f0ad | !hbusreq0 & v84563c;
assign a5eea4 = hbusreq1 & a5eea3 | !hbusreq1 & !v84563c;
assign dea6be = hmaster0_p & deaeb2 | !hmaster0_p & dea6bd;
assign af3c56 = hlock1_p & d40d33 | !hlock1_p & af3c4c;
assign ab0c3c = hlock0_p & v84563c | !hlock0_p & !b29a65;
assign b29f0f = hlock1_p & v84565a | !hlock1_p & !b29f0e;
assign af357d = hmaster0_p & af3536 | !hmaster0_p & af357c;
assign a5f95d = hmaster0_p & a5f959 | !hmaster0_p & a5f95c;
assign cea31d = hbusreq2_p & cea16b | !hbusreq2_p & v845660;
assign a5f46d = hmastlock_p & a5f833 | !hmastlock_p & v84563c;
assign deae43 = hmaster1_p & deae42 | !hmaster1_p & deade4;
assign a5f1f6 = hready & v84563c | !hready & dead0c;
assign ab0578 = hmaster0_p & ab0555 | !hmaster0_p & ab0577;
assign a5f99a = hmaster0_p & a5f968 | !hmaster0_p & a5f999;
assign c3b66e = hlock2_p & c3b66c | !hlock2_p & !c3b66b;
assign af34de = hgrant2_p & af34dd | !hgrant2_p & af3c64;
assign af35c2 = hbusreq3_p & af35a2 | !hbusreq3_p & af35c1;
assign af3c6a = start_p & v84563c | !start_p & !af3c69;
assign a5fcb3 = hbusreq2 & a5fc7f | !hbusreq2 & a5fc91;
assign a5f303 = hmaster1_p & a5f302 | !hmaster1_p & a5f215;
assign ab0be5 = hgrant2_p & ab0be2 | !hgrant2_p & ab0be4;
assign b2676e = decide_p & b2676b | !decide_p & b2676d;
assign c3bd3a = hgrant1_p & c3bd39 | !hgrant1_p & c3bd37;
assign ab0517 = hbusreq2_p & ab0516 | !hbusreq2_p & b298a4;
assign a60179 = hready & a60171 | !hready & a60178;
assign b2992a = hlock1_p & c3b683 | !hlock1_p & !b29929;
assign c3b77e = hgrant3_p & c3b777 | !hgrant3_p & c3b77d;
assign a5f7b4 = hready & v84563c | !hready & a5f9f9;
assign ab0604 = hbusreq2_p & ab0603 | !hbusreq2_p & ab058d;
assign deaead = hready_p & deae70 | !hready_p & deaeac;
assign a5f7cb = hready & v84563c | !hready & !ab06af;
assign a5f01e = hbusreq0 & a5fae2 | !hbusreq0 & a5f01d;
assign bdb5a3 = hmaster1_p & bdb598 | !hmaster1_p & !v84565a;
assign ab061a = hlock2 & ab05dc | !hlock2 & ab0619;
assign a5ef05 = hmaster1_p & a5edf5 | !hmaster1_p & v84563c;
assign b29fe5 = hgrant2_p & b29fe2 | !hgrant2_p & b29fe4;
assign cea453 = hbusreq2_p & cea452 | !hbusreq2_p & cea37b;
assign c3bdca = hmaster0_p & c3bdc4 | !hmaster0_p & c3bdc9;
assign af3c22 = hgrant2_p & af3c21 | !hgrant2_p & af3c1f;
assign af349c = hlock0_p & af3c5d | !hlock0_p & af3c4c;
assign b299dc = hmaster0_p & b299db | !hmaster0_p & b2997a;
assign a5f0ec = hlock2_p & a5f0e6 | !hlock2_p & a5f0eb;
assign a5fbc9 = hlock2 & a5fb74 | !hlock2 & a5fbc8;
assign c3b893 = hmaster1_p & c3b88f | !hmaster1_p & c3b892;
assign cea298 = hbusreq2_p & cea297 | !hbusreq2_p & v84563c;
assign cea420 = hlock0_p & cea41f | !hlock0_p & cea405;
assign b29fd5 = hlock2_p & b29fd1 | !hlock2_p & !b29fd4;
assign a5f744 = hbusreq2 & a5f742 | !hbusreq2 & a5f743;
assign ab0ae6 = hlock0_p & v84563c | !hlock0_p & !b29a5a;
assign a5f9e8 = hready & a5f9e7 | !hready & deadb2;
assign b29cf0 = hready & c3bc02 | !hready & !v84563c;
assign ab0612 = hlock0_p & v84563c | !hlock0_p & ab0611;
assign cea492 = hmaster1_p & cea491 | !hmaster1_p & v84563c;
assign ab0cb6 = hmaster1_p & ab0cb4 | !hmaster1_p & ab0cb5;
assign b29ae2 = hready & c3bd37 | !hready & c3b683;
assign c3b676 = hburst0 & v84563c | !hburst0 & c3b675;
assign ce9d42 = decide_p & ce9d41 | !decide_p & v84563c;
assign cea16d = locked_p & v84563c | !locked_p & !cea16c;
assign c3bbbf = hbusreq3 & c3bbbe | !hbusreq3 & v84563c;
assign c3bce0 = locked_p & dead7b | !locked_p & !v84563c;
assign c3b63e = hbusreq3 & c3b638 | !hbusreq3 & c3b63d;
assign c3b632 = hlock0_p & c3bbbb | !hlock0_p & c3b631;
assign c3bc96 = hbusreq2_p & c3bc95 | !hbusreq2_p & !v84563c;
assign a60170 = hlock1_p & a6016f | !hlock1_p & !v84563c;
assign af34f7 = hmaster1_p & af34f6 | !hmaster1_p & d40d60;
assign b29d84 = hlock0_p & b29d83 | !hlock0_p & !v84563c;
assign b29e98 = decide_p & b29e97 | !decide_p & b29e57;
assign a81d0a = decide_p & a81cc6 | !decide_p & a81cff;
assign af3c70 = hbusreq2_p & af3c5e | !hbusreq2_p & af3c4c;
assign ab0563 = hlock0_p & v84563c | !hlock0_p & !b29947;
assign c3bdf4 = hmaster1_p & c3bd6c | !hmaster1_p & c3bd72;
assign a5f9f5 = hgrant1_p & a5f9f4 | !hgrant1_p & a60168;
assign a5fa12 = stateG10_1_p & v970407 | !stateG10_1_p & v9703fb;
assign a5f145 = hlock0_p & a5f864 | !hlock0_p & a5f144;
assign ab051e = hbusreq3 & ab051d | !hbusreq3 & ab0517;
assign a5f492 = hbusreq1 & a5f491 | !hbusreq1 & v84563c;
assign af34ef = hmaster0_p & af34ee | !hmaster0_p & af348f;
assign a5f947 = hlock0_p & a5f946 | !hlock0_p & a5f8c5;
assign bdb587 = hbusreq2_p & bdb586 | !hbusreq2_p & v84565a;
assign af3531 = hbusreq2_p & v84563c | !hbusreq2_p & af352c;
assign cea440 = hlock3_p & cea41a | !hlock3_p & cea43f;
assign af34aa = hmaster1_p & af34a5 | !hmaster1_p & af34a9;
assign ab0b66 = hlock0_p & ab0b64 | !hlock0_p & ab0b65;
assign a5ea21 = hbusreq0_p & a5fcdf | !hbusreq0_p & !v84563c;
assign deaddc = hgrant2_p & deadd8 | !hgrant2_p & deaddb;
assign a5f8c7 = hbusreq2 & a5f8c1 | !hbusreq2 & a5f8c6;
assign ab0713 = hlock2_p & ab06b8 | !hlock2_p & ab0712;
assign b29a1a = hmaster0_p & b29e48 | !hmaster0_p & b29a19;
assign ab0b3a = hlock2_p & ab0b38 | !hlock2_p & ab0b39;
assign a5f29e = hmaster0_p & a5f29d | !hmaster0_p & !a5f755;
assign cea1b1 = hmastlock_p & cea1b0 | !hmastlock_p & !v84563c;
assign a5fb76 = hlock0_p & a5fb75 | !hlock0_p & a5fb73;
assign a5efd8 = hlock0_p & a5fa6c | !hlock0_p & a5ef6b;
assign c3b642 = hlock2_p & c3b640 | !hlock2_p & c3b641;
assign cea327 = hlock2_p & cea326 | !hlock2_p & !cea17a;
assign c3bd67 = hmaster1_p & c3bcd1 | !hmaster1_p & c3bd66;
assign cea246 = start_p & cea1aa | !start_p & v84563c;
assign dead4c = hmaster0_p & dead44 | !hmaster0_p & !dead4b;
assign dead26 = hbusreq2_p & deacfe | !hbusreq2_p & dead25;
assign cea35b = hlock0_p & dead19 | !hlock0_p & v845660;
assign deacfa = locked_p & deacf9 | !locked_p & !b2671f;
assign c3bcaf = hlock3_p & c3bc9f | !hlock3_p & c3bcae;
assign a5eb4e = hmaster0_p & a5eb4d | !hmaster0_p & a5f0a0;
assign ab0cd6 = hbusreq3 & ab0cd4 | !hbusreq3 & ab0cd5;
assign a5f560 = hready & a5f520 | !hready & a5f40c;
assign d40d91 = hmaster0_p & d40d90 | !hmaster0_p & d40d60;
assign a5f3f0 = stateG10_1_p & v84563c | !stateG10_1_p & a5f3ef;
assign dead3d = hlock2_p & v845660 | !hlock2_p & !v84563c;
assign af3c40 = hgrant3_p & af3c2a | !hgrant3_p & af3c3f;
assign c3bc0c = hbusreq2_p & c3bc0b | !hbusreq2_p & deac7b;
assign a5fbe4 = start_p & v8e1935 | !start_p & !a5fbac;
assign c3b6d8 = hlock2_p & c3b6d6 | !hlock2_p & c3b6d7;
assign a5ead4 = hlock0_p & a5fa5e | !hlock0_p & a5ead1;
assign b26716 = hbusreq0_p & b266b8 | !hbusreq0_p & !b26715;
assign adaec3 = start_p & a81ca6 | !start_p & adaec2;
assign a5f8bb = hlock0_p & a5f8b8 | !hlock0_p & a5f8ba;
assign deae89 = hbusreq3 & deae7b | !hbusreq3 & deae88;
assign dead95 = hlock2_p & dead94 | !hlock2_p & !v84563c;
assign af3510 = hbusreq3_p & af34fc | !hbusreq3_p & af350f;
assign a5f284 = hbusreq2_p & a5f283 | !hbusreq2_p & v84563c;
assign af3c63 = hlock0_p & af3c5d | !hlock0_p & af3c62;
assign a5f040 = hgrant2_p & a5f03f | !hgrant2_p & a5f020;
assign c3b72c = hready_p & c3b711 | !hready_p & c3b72b;
assign ab0ce8 = hbusreq2_p & ab0ce7 | !hbusreq2_p & ab0b5f;
assign c3b638 = hbusreq2_p & c3b633 | !hbusreq2_p & c3b637;
assign a5f251 = hbusreq2 & a5f250 | !hbusreq2 & ab0c31;
assign d40d53 = hgrant2_p & d40d4e | !hgrant2_p & d40d52;
assign dead22 = hbusreq2_p & deacfe | !hbusreq2_p & dead21;
assign ab0cc2 = hlock0_p & v84563c | !hlock0_p & !b29ae2;
assign a5f2c7 = hbusreq2 & ab0c31 | !hbusreq2 & a5f908;
assign a5f094 = hlock0_p & a5f71d | !hlock0_p & v84563c;
assign v9703fe = hmaster1_p & v9703fd | !hmaster1_p & v84563c;
assign deaeab = hlock3_p & deae8f | !hlock3_p & deaeaa;
assign cea3eb = hlock0_p & cea3dc | !hlock0_p & cea3ea;
assign deae7b = hbusreq2_p & deae7a | !hbusreq2_p & !deadb2;
assign a5f199 = hbusreq2 & a5f198 | !hbusreq2 & a5fa6b;
assign dea765 = hbusreq2_p & deae07 | !hbusreq2_p & v84563c;
assign a5ea26 = hmaster1_p & a5ea23 | !hmaster1_p & a5ea25;
assign a5ea7d = hready & a5f6e4 | !hready & v84563c;
assign c3bdc4 = hmaster1_p & c3bdb8 | !hmaster1_p & c3bdc3;
assign a5fbac = stateA1_p & a81ca7 | !stateA1_p & !v84563c;
assign c3b62d = hlock2_p & c3b62c | !hlock2_p & !c3b62b;
assign ab0672 = hbusreq2_p & ab0671 | !hbusreq2_p & ab066f;
assign b2995a = hbusreq2_p & b29959 | !hbusreq2_p & !b29943;
assign c3b6fc = hlock2_p & c3b6fb | !hlock2_p & !c3b6e3;
assign a5efc1 = hbusreq2 & a5efc0 | !hbusreq2 & a5ee77;
assign cea32e = hlock3_p & cea2f9 | !hlock3_p & cea32d;
assign a5f8cb = hbusreq2 & a5f8c9 | !hbusreq2 & a5f8ca;
assign c3b649 = locked_p & v84563c | !locked_p & !v845648;
assign ab0b5a = hmaster1_p & ab0b54 | !hmaster1_p & ab0b59;
assign d40d94 = hlock2_p & d40d51 | !hlock2_p & d40d33;
assign a5f20d = hbusreq2 & a5fc93 | !hbusreq2 & !v84563c;
assign a5fa58 = hbusreq3 & a5fa28 | !hbusreq3 & a5fa57;
assign a5f751 = hbusreq2_p & a5f750 | !hbusreq2_p & v84563c;
assign ab0b38 = hlock2 & ab0ad1 | !hlock2 & ab0b37;
assign ab0b87 = hmaster1_p & ab0b71 | !hmaster1_p & ab0b86;
assign a60185 = stateA1_p & a60184 | !stateA1_p & c06d34;
assign cea26e = hgrant1_p & cea26c | !hgrant1_p & cea26d;
assign c3bd42 = hbusreq2_p & c3bd41 | !hbusreq2_p & v84563c;
assign a5f153 = hready & v84563c | !hready & v845648;
assign deac6b = hgrant1_p & deac52 | !hgrant1_p & deac6a;
assign a5f569 = hbusreq2_p & a5f568 | !hbusreq2_p & a5f567;
assign a81cfe = hmaster0_p & a81cfa | !hmaster0_p & a81cfd;
assign b29e5a = hready_p & b29e58 | !hready_p & b29e59;
assign a5f47a = hbusreq3 & a5f478 | !hbusreq3 & !a5f479;
assign b29d37 = hbusreq2_p & b29d35 | !hbusreq2_p & b29d36;
assign a5fbcd = hlock2_p & a5fbca | !hlock2_p & a5fbcc;
assign deaea5 = hbusreq2_p & deaea3 | !hbusreq2_p & deae95;
assign c3b643 = hbusreq2_p & c3b642 | !hbusreq2_p & c3b640;
assign a5f394 = hbusreq0_p & a5f385 | !hbusreq0_p & a5f390;
assign a9b9db = hmaster1_p & v84563c | !hmaster1_p & a9b9da;
assign a5f836 = hlock1_p & a5f833 | !hlock1_p & a5f835;
assign c98b9f = hready_p & v8c6711 | !hready_p & c98b9e;
assign cea1a5 = hmaster0_p & cea1a2 | !hmaster0_p & !cea1a4;
assign ab0cfb = hgrant2_p & ab0cfa | !hgrant2_p & ab0c62;
assign deac89 = hlock2_p & deac87 | !hlock2_p & deac88;
assign c3b6d1 = hmaster1_p & c3b6ca | !hmaster1_p & c3b6d0;
assign c3b6c6 = hready & c3b6c4 | !hready & c3b6c5;
assign ab0bd9 = hlock0_p & v84565a | !hlock0_p & ab0bd8;
assign c3b6f0 = hbusreq2_p & c3b6ef | !hbusreq2_p & !c3b656;
assign af3509 = hgrant0_p & af3506 | !hgrant0_p & af3508;
assign a5f1b7 = hbusreq2_p & a5f1b6 | !hbusreq2_p & v84563c;
assign ce9d15 = hlock3_p & ce9cfd | !hlock3_p & ce9d14;
assign a5f5a3 = hlock0_p & a5f5a2 | !hlock0_p & a5f495;
assign dea75a = hmaster0_p & dea753 | !hmaster0_p & dea759;
assign cea2a1 = hlock0_p & cea2a0 | !hlock0_p & v84563c;
assign c3bcfe = hbusreq2_p & c3bcfd | !hbusreq2_p & v84563c;
assign b2996c = hbusreq2_p & b2996b | !hbusreq2_p & !b2994b;
assign a5f3f5 = stateG10_1_p & v84563c | !stateG10_1_p & a5f3f4;
assign a5ea70 = hgrant2_p & a5ea35 | !hgrant2_p & a5f089;
assign c3bcb5 = hmaster1_p & v84563c | !hmaster1_p & c3bcb4;
assign a5f988 = hmastlock_p & a5f987 | !hmastlock_p & !v84563c;
assign a5f38d = hlock1_p & b266a0 | !hlock1_p & !v84563c;
assign a5f592 = hbusreq2 & a5f4f0 | !hbusreq2 & a5f4f1;
assign b29960 = hbusreq3 & b2995e | !hbusreq3 & b2995f;
assign a5f48a = hready & a5f489 | !hready & !c3b694;
assign ce9d32 = hbusreq3 & ce9d30 | !hbusreq3 & ce9d31;
assign b26730 = hgrant2_p & b26726 | !hgrant2_p & !b2672f;
assign a5fbf6 = hbusreq3 & a5fbf5 | !hbusreq3 & v84563c;
assign b29d3c = hbusreq2_p & b29d35 | !hbusreq2_p & !v84563c;
assign af34e2 = hlock3_p & af34cd | !hlock3_p & af34e1;
assign b26783 = hgrant0_p & b26780 | !hgrant0_p & b26782;
assign b29f4f = hgrant2_p & b29cfb | !hgrant2_p & b29d05;
assign dea762 = hbusreq2_p & deae13 | !hbusreq2_p & deae12;
assign deaca0 = start_p & v845652 | !start_p & !v8c607d;
assign c3bd77 = hbusreq1_p & c3bd11 | !hbusreq1_p & c3bbd2;
assign b29919 = hgrant1_p & b29918 | !hgrant1_p & deacbc;
assign af34d4 = hgrant2_p & af34d3 | !hgrant2_p & af3c5e;
assign ab06b9 = hgrant1_p & b29ee9 | !hgrant1_p & ab06a9;
assign cea85e = hlock2_p & cea85d | !hlock2_p & v84563c;
assign c3bda6 = hlock0_p & c3bcee | !hlock0_p & !c3bcdb;
assign a5eedc = hlock0_p & a5f565 | !hlock0_p & a5f560;
assign ab05b0 = hbusreq0_p & ab0598 | !hbusreq0_p & ab05af;
assign ce9dfe = hgrant2_p & cea15e | !hgrant2_p & !ce9dfd;
assign b29972 = hbusreq2_p & b29971 | !hbusreq2_p & v84563c;
assign b26737 = hbusreq2_p & b26722 | !hbusreq2_p & b26736;
assign ab0735 = hmaster0_p & ab0733 | !hmaster0_p & ab0734;
assign b29d83 = locked_p & v84563c | !locked_p & b29d82;
assign adaef2 = locked_p & adaef1 | !locked_p & v84563c;
assign af358f = hmaster0_p & af358c | !hmaster0_p & af358e;
assign a5f22f = hready & a60168 | !hready & a5f797;
assign c3b639 = locked_p & v84563c | !locked_p & deae59;
assign b29ab1 = hlock2_p & b29ab0 | !hlock2_p & b29d81;
assign cea15f = hready & dead08 | !hready & v84563c;
assign c3b6b3 = hbusreq2_p & c3b6b2 | !hbusreq2_p & !c3b6b1;
assign a5fcfc = hready & a5fcf6 | !hready & a5fcfb;
assign c3bc47 = hready & b2671f | !hready & !v84563c;
assign a5eb8f = hbusreq2 & a5f09c | !hbusreq2 & a5fc1a;
assign b266b4 = hlock2_p & b266b2 | !hlock2_p & b266b3;
assign c3bc39 = hbusreq2_p & c3bc38 | !hbusreq2_p & v84563c;
assign v84566e = stateG2_p & v84563c | !stateG2_p & !v84563c;
assign ab0ba2 = hlock0_p & v84563c | !hlock0_p & ab0ba1;
assign ab06c8 = hgrant1_p & b29eea | !hgrant1_p & b29f76;
assign a5fae6 = hbusreq0 & a5fae4 | !hbusreq0 & !a5fae5;
assign a5f6e5 = hbusreq1_p & a5fb8c | !hbusreq1_p & !a5fb8b;
assign cea374 = hbusreq1_p & dead33 | !hbusreq1_p & !v84563c;
assign ab06d7 = hmaster0_p & ab06c7 | !hmaster0_p & ab06d6;
assign b26774 = hbusreq2_p & b26773 | !hbusreq2_p & b26713;
assign c3bbfc = hlock0_p & c3bbf9 | !hlock0_p & !c3bbfb;
assign dea7a1 = hmaster1_p & dea7a0 | !hmaster1_p & dea731;
assign a5f4ef = hbusreq1 & c3b6a0 | !hbusreq1 & v84563c;
assign cea0d2 = hbusreq3 & cea0ca | !hbusreq3 & cea86e;
assign cea447 = hmaster1_p & cea446 | !hmaster1_p & cea85f;
assign c3bdbc = hlock1_p & deae02 | !hlock1_p & !c3bdbb;
assign af34c5 = hlock2_p & af3c63 | !hlock2_p & af3c4c;
assign af348a = hbusreq2_p & af3489 | !hbusreq2_p & d40d33;
assign a5fc81 = hlock0_p & a5fc7a | !hlock0_p & a5fc80;
assign af3c16 = hmaster0_p & af3c15 | !hmaster0_p & af3c14;
assign dead8f = hlock2_p & dead2e | !hlock2_p & !v84563c;
assign ab0c0f = hlock2_p & ab0c0e | !hlock2_p & v84563c;
assign ce9ccd = hready_p & ce9cbe | !hready_p & !ce9ccc;
assign a5fd37 = hbusreq2_p & a5fd36 | !hbusreq2_p & v84563c;
assign a5ea9b = hbusreq0_p & a5fc7f | !hbusreq0_p & !v84563c;
assign b8aced = hgrant0_p & b8acd9 | !hgrant0_p & b8acec;
assign a5ef8d = hbusreq0 & a5ef8a | !hbusreq0 & a5ef8c;
assign ab06c1 = hlock0_p & b2a00e | !hlock0_p & v84563c;
assign ab0551 = hbusreq2_p & ab0540 | !hbusreq2_p & ab053e;
assign ab066e = hbusreq2_p & ab066d | !hbusreq2_p & ab066b;
assign b29fc5 = hbusreq2_p & b29fc4 | !hbusreq2_p & v84563c;
assign af3c2a = hready_p & af3c18 | !hready_p & af3c29;
assign ab0703 = hlock3_p & ab06f0 | !hlock3_p & ab0702;
assign ce9d71 = hgrant2_p & cea338 | !hgrant2_p & ce9d70;
assign cea37b = hready & deae5a | !hready & deae59;
assign a5f3c8 = hready & a5f3c7 | !hready & v84563c;
assign a5eb48 = hready_p & a5eaa4 | !hready_p & a5eb47;
assign a5f378 = hlock1_p & a5fbab | !hlock1_p & !a5f377;
assign c3bd22 = hlock0_p & c3bd17 | !hlock0_p & !c3bd21;
assign a5f842 = hlock1_p & a5f83f | !hlock1_p & a5f841;
assign a5ef17 = hmaster1_p & a5edfe | !hmaster1_p & a5ef16;
assign a5f979 = hbusreq2 & a5f978 | !hbusreq2 & a5f6fa;
assign a81cfa = hmaster1_p & v84563c | !hmaster1_p & a81cf9;
assign c3b6ce = hbusreq2_p & c3b6cd | !hbusreq2_p & c3b6b1;
assign b29d99 = hmaster1_p & b29d91 | !hmaster1_p & b29d98;
assign b29eb7 = hmastlock_p & b29eb6 | !hmastlock_p & !v84563c;
assign af354d = hlock0_p & af3548 | !hlock0_p & af354c;
assign a5ee24 = locked_p & v845646 | !locked_p & v845641;
assign b29fda = hready & b29f19 | !hready & v84563c;
assign c3b7b6 = hlock3_p & c3b7aa | !hlock3_p & !c3b7b5;
assign ab0c1f = hbusreq3 & ab0c1b | !hbusreq3 & ab0c1e;
assign a6016d = stateA1_p & a81ca7 | !stateA1_p & a6016c;
assign ab0c5b = hlock1_p & v84565a | !hlock1_p & !ab0c5a;
assign b2670b = hlock0_p & b266a8 | !hlock0_p & !b26695;
assign ce9d26 = hbusreq2_p & cea286 | !hbusreq2_p & !cea887;
assign a5fa1d = hmastlock_p & v970407 | !hmastlock_p & !v84563c;
assign b26761 = hbusreq2_p & b26699 | !hbusreq2_p & !b26757;
assign a5eb93 = hlock0_p & a5fc1c | !hlock0_p & v84563c;
assign b29d78 = hready & b29d77 | !hready & !v84563c;
assign af3565 = hgrant2_p & af355e | !hgrant2_p & af3564;
assign a81ca9 = hmastlock_p & a81ca8 | !hmastlock_p & v84563c;
assign cea24d = start_p & cea1aa | !start_p & !cea24c;
assign a5fc9c = hbusreq3 & a5fc9b | !hbusreq3 & v84563c;
assign ab0b71 = hgrant2_p & ab0b70 | !hgrant2_p & cea15a;
assign ab0ba9 = hlock0_p & v84563c | !hlock0_p & !ab0ba8;
assign a5eea2 = hbusreq1 & a5eea1 | !hbusreq1 & !v84563c;
assign ab06b2 = hlock0_p & ab06ac | !hlock0_p & !ab06b1;
assign cea367 = hlock2_p & cea366 | !hlock2_p & v84563c;
assign dead75 = start_p & v845652 | !start_p & !dead74;
assign c3b726 = hbusreq3 & c3b724 | !hbusreq3 & c3b725;
assign bdb5b6 = hmaster0_p & bdb5b5 | !hmaster0_p & !bdb595;
assign b2673d = hbusreq2_p & b2673c | !hbusreq2_p & b2673b;
assign a5ee7c = hmaster1_p & a5ee6b | !hmaster1_p & a5ee7b;
assign a5f7cf = hlock2_p & a5f7bc | !hlock2_p & a5f7ce;
assign a81ce7 = hgrant2_p & a81ce6 | !hgrant2_p & v84563c;
assign c3b70f = hgrant0_p & c3b6ff | !hgrant0_p & c3b70e;
assign b26740 = hmaster0_p & b26731 | !hmaster0_p & !b2673f;
assign b29a66 = hlock0_p & b29a65 | !hlock0_p & !v84563c;
assign a5f389 = hbusreq2 & a5f385 | !hbusreq2 & a5f388;
assign a81ce2 = hlock1_p & a81ca9 | !hlock1_p & a81ce1;
assign ab0ccf = decide_p & ab0cce | !decide_p & !v845662;
assign b29feb = hgrant3_p & b29f85 | !hgrant3_p & b29fea;
assign a5edf3 = hbusreq3 & a5edec | !hbusreq3 & !a5edf2;
assign af3501 = hmaster0_p & af3500 | !hmaster0_p & af34aa;
assign bdb5b1 = hlock2_p & bdb58b | !hlock2_p & !v84565a;
assign a5fbec = hbusreq1 & a5fbeb | !hbusreq1 & a5fbb6;
assign a5f804 = hgrant1_p & a5f7f6 | !hgrant1_p & a5f7f5;
assign cea44e = hlock2_p & cea44c | !hlock2_p & cea44d;
assign a5f14c = hbusreq2 & a5f146 | !hbusreq2 & a5f14b;
assign c3bdac = hmaster1_p & c3bda8 | !hmaster1_p & c3bdab;
assign a5f863 = hbusreq1 & a5f861 | !hbusreq1 & !a5f862;
assign cea31f = hburst1 & v84563c | !hburst1 & !v84566c;
assign a5fa1f = hgrant1_p & a5fa1e | !hgrant1_p & a5fa1c;
assign ab0be2 = hbusreq2_p & ab0b6f | !hbusreq2_p & v845644;
assign ab0af2 = hlock0_p & v84563c | !hlock0_p & !deac52;
assign dead08 = hlock1_p & deacf7 | !hlock1_p & v84563c;
assign dead01 = hbusreq3 & dead00 | !hbusreq3 & v84563c;
assign a5f98e = hlock2 & a5f985 | !hlock2 & a5f98d;
assign ab0b93 = hbusreq2_p & ab0b8f | !hbusreq2_p & ab0b92;
assign af35b5 = hbusreq2_p & af35b4 | !hbusreq2_p & af352c;
assign c3bbd3 = hlock1_p & c3bbd2 | !hlock1_p & deac5a;
assign a5f9db = stateA1_p & v84563c | !stateA1_p & !a5f9da;
assign dead50 = decide_p & deacda | !decide_p & !v84563c;
assign d40d70 = hgrant2_p & v84563c | !hgrant2_p & d40d6f;
assign b29e6d = hbusreq2_p & b29d17 | !hbusreq2_p & b29cbb;
assign a5fcc2 = hmaster0_p & a5fcae | !hmaster0_p & a5fcc1;
assign b299db = hmaster1_p & b299da | !hmaster1_p & c3bceb;
assign a5ee4d = locked_p & a5ee4c | !locked_p & a60140;
assign a5efad = hlock2_p & a5efaa | !hlock2_p & a5efac;
assign a5f32c = hbusreq2_p & a5f325 | !hbusreq2_p & a5fa6d;
assign b29eed = hready & b29eec | !hready & v84563c;
assign ab06bc = hready & deaca1 | !hready & deaca0;
assign deadc8 = hbusreq3 & deadb5 | !hbusreq3 & deadc7;
assign af359b = hmaster1_p & v84563c | !hmaster1_p & af359a;
assign cea280 = hready & deac57 | !hready & c98b96;
assign b29d9b = hgrant0_p & b29d63 | !hgrant0_p & !b29d9a;
assign cea272 = hgrant1_p & cea270 | !hgrant1_p & cea271;
assign dea6cf = hlock1_p & v84565a | !hlock1_p & !dea6ce;
assign a81ceb = decide_p & a81cd9 | !decide_p & a81cea;
assign a5ea1d = hmaster0_p & a5e9eb | !hmaster0_p & a5ea1c;
assign dead06 = hbusreq2_p & dead05 | !hbusreq2_p & deace1;
assign a5f1ff = hlock0_p & a5f726 | !hlock0_p & a5f729;
assign deac3f = hgrant2_p & deac2a | !hgrant2_p & deac3e;
assign a5f6f7 = hbusreq2 & a5f6f1 | !hbusreq2 & a5f6f6;
assign b29ec4 = hbusreq3 & b29eb2 | !hbusreq3 & b29ec3;
assign b29abd = locked_p & deae02 | !locked_p & !v84563c;
assign dea79b = hlock3_p & dea78b | !hlock3_p & dea75a;
assign a81d01 = hready_p & a81ceb | !hready_p & a81d00;
assign c3bd72 = hbusreq2_p & c3bd71 | !hbusreq2_p & !deacaa;
assign a5f1e5 = locked_p & a5f1d6 | !locked_p & v845641;
assign a5eb9f = hgrant2_p & a5eb9d | !hgrant2_p & a5eb9e;
assign c3bc50 = hbusreq2_p & c3bc4f | !hbusreq2_p & c3bc4c;
assign dea6fd = decide_p & dea6f7 | !decide_p & !v84563c;
assign b26754 = hlock3_p & b26741 | !hlock3_p & b26753;
assign ab0cbd = hready & deadde | !hready & !v84565a;
assign a5fb79 = hready & v84563c | !hready & !b26697;
assign a5f926 = hbusreq2_p & a5f925 | !hbusreq2_p & v84563c;
assign ab0d00 = hgrant3_p & ab0ce5 | !hgrant3_p & !ab0cff;
assign b29efa = hready & deacb7 | !hready & !v84563c;
assign b2674d = hbusreq2_p & b2674c | !hbusreq2_p & !b26715;
assign d40d31 = hmastlock_p & d40d30 | !hmastlock_p & v84563c;
assign a5f1a8 = hbusreq2 & a5f1a7 | !hbusreq2 & v84563c;
assign b299cd = hlock2_p & v84563c | !hlock2_p & !b29948;
assign deacd7 = hgrant2_p & deacd4 | !hgrant2_p & deacd6;
assign a5f6e3 = hbusreq3_p & a5fd1c | !hbusreq3_p & a5f6e2;
assign deae61 = hlock2_p & deae60 | !hlock2_p & !v84563c;
assign a5f3b8 = hbusreq0_p & a5f36b | !hbusreq0_p & a5f38f;
assign a5f26a = hmaster1_p & a5f269 | !hmaster1_p & a5f958;
assign a5fcd2 = locked_p & a5fcd1 | !locked_p & c3bd5f;
assign ab0689 = decide_p & ab0688 | !decide_p & v84563c;
assign c3bc69 = hbusreq3 & c3bc68 | !hbusreq3 & c3bc5e;
assign ab06f7 = hmaster1_p & ab06f1 | !hmaster1_p & ab06f6;
assign a5f3bb = hlock0_p & a5f36e | !hlock0_p & a5f3b8;
assign a5efaa = hbusreq2 & a5efa8 | !hbusreq2 & a5efa9;
assign a5fb92 = hbusreq0_p & v84563c | !hbusreq0_p & a5fb91;
assign b26723 = hbusreq2_p & b26722 | !hbusreq2_p & b26721;
assign a5fbb8 = locked_p & a5fbb7 | !locked_p & v84563c;
assign cea165 = hbusreq3 & cea164 | !hbusreq3 & cea15c;
assign deadab = hgrant1_p & deada9 | !hgrant1_p & deadaa;
assign a60193 = hmastlock_p & a60192 | !hmastlock_p & v84563c;
assign ab0690 = hbusreq2_p & ab068f | !hbusreq2_p & ab068e;
assign a5fb22 = hlock2_p & a5fb21 | !hlock2_p & v84563c;
assign ab0c8f = hbusreq2_p & ab0c8e | !hbusreq2_p & ab0b5f;
assign b0c0fe = hready_p & b29e57 | !hready_p & !v845658;
assign ab0699 = hlock0_p & b29f1d | !hlock0_p & !b29f1f;
assign a5f24e = hready & a5f833 | !hready & !a5f83f;
assign c3bd08 = hlock3_p & c3bcf7 | !hlock3_p & !c3bd07;
assign b29d6b = hbusreq3 & b29d6a | !hbusreq3 & c3bcfb;
assign ab0ca5 = hmaster0_p & ab0ca1 | !hmaster0_p & ab0ca4;
assign adaf19 = decide_p & adaed5 | !decide_p & adaf0e;
assign a5f039 = hbusreq0 & a5fd37 | !hbusreq0 & a5f038;
assign af3590 = hgrant0_p & af358a | !hgrant0_p & af358f;
assign a5ee91 = hbusreq0 & a5ee89 | !hbusreq0 & !a5ee90;
assign ab05e1 = hbusreq3 & ab05dd | !hbusreq3 & ab05e0;
assign ce9d4d = hbusreq2_p & cea16b | !hbusreq2_p & cea35b;
assign deacd3 = hbusreq2_p & deacd2 | !hbusreq2_p & v84563c;
assign ab057b = hbusreq2_p & ab0560 | !hbusreq2_p & ab0565;
assign b29f31 = hready & deadc4 | !hready & !v84563c;
assign v84564b = hbusreq2 & v84563c | !hbusreq2 & !v84563c;
assign a5f4c7 = hbusreq1_p & a60186 | !hbusreq1_p & v84563c;
assign ab0bcb = hmaster1_p & dead53 | !hmaster1_p & ab0bca;
assign cea86c = hlock0_p & deac19 | !hlock0_p & v84563c;
assign a5fb29 = hbusreq2 & a5fb28 | !hbusreq2 & ab0c32;
assign ce9ddb = hmaster0_p & ce9dda | !hmaster0_p & ce9d3f;
assign cea3ad = hmaster0_p & cea3a3 | !hmaster0_p & cea3ac;
assign d40d82 = hlock1_p & d40d33 | !hlock1_p & !d40d3b;
assign c3bc85 = locked_p & cea151 | !locked_p & b2671f;
assign a5fb36 = hbusreq3 & a5fb35 | !hbusreq3 & a5fb2d;
assign ab0c48 = hbusreq2_p & ab0c46 | !hbusreq2_p & ab0add;
assign b29ead = hready & deae02 | !hready & v84563c;
assign a5f3de = decide_p & a5f3c2 | !decide_p & a5f3dd;
assign b266ff = hgrant2_p & b266fd | !hgrant2_p & b266fe;
assign ab0533 = hlock3_p & ab0520 | !hlock3_p & ab0532;
assign cea44c = hlock0_p & cea379 | !hlock0_p & cea44b;
assign c3b625 = hready & c3b624 | !hready & v84563c;
assign b29ff6 = hbusreq2_p & b29f7d | !hbusreq2_p & b29cbb;
assign ab0b0c = hlock2 & ab0b09 | !hlock2 & ab0b0b;
assign a5fc05 = locked_p & a5fc04 | !locked_p & v845641;
assign a5f709 = hready & a5f706 | !hready & a5f708;
assign ab0655 = hbusreq3_p & ab0654 | !hbusreq3_p & ab0bf8;
assign c3bd87 = hlock2_p & c3bd86 | !hlock2_p & dead2e;
assign c3bcc7 = hbusreq2_p & c3bcc6 | !hbusreq2_p & !v84563c;
assign v970433 = hmaster0_p & v84563c | !hmaster0_p & v970432;
assign a5edc2 = hlock2 & a5edbf | !hlock2 & a5edc1;
assign a5ee49 = locked_p & a5ee48 | !locked_p & a5f36b;
assign c3bbea = hlock2_p & c3bbe8 | !hlock2_p & deacaa;
assign c3bc6f = hlock2_p & c3bc6e | !hlock2_p & v845660;
assign c3bce9 = hbusreq2_p & c3bce8 | !hbusreq2_p & c3bbbc;
assign cea33c = hmaster0_p & cea33b | !hmaster0_p & cea29b;
assign ab0b56 = hlock0_p & c3bc52 | !hlock0_p & v84563c;
assign b8acda = stateG10_1_p & v84563c | !stateG10_1_p & v845646;
assign b840b2 = hready_p & b840b1 | !hready_p & b840ae;
assign c3bc59 = hlock2_p & c3bc58 | !hlock2_p & b2670b;
assign a5fba5 = start_p & a5fba3 | !start_p & a5fba4;
assign c3b6aa = hlock2_p & c3b6a9 | !hlock2_p & !c3b698;
assign a5edd5 = hlock0_p & a5edd4 | !hlock0_p & a5f55b;
assign v845643 = hbusreq0 & v84563c | !hbusreq0 & !v84563c;
assign ab0c2c = hlock3_p & ab0c19 | !hlock3_p & ab0c2b;
assign cea462 = locked_p & cea376 | !locked_p & cea37b;
assign dead80 = hlock0_p & dead7e | !hlock0_p & !dead7f;
assign deacab = hlock0_p & deacaa | !hlock0_p & v84563c;
assign b29eab = hready & dead33 | !hready & !v84563c;
assign af3c27 = hmaster0_p & v877992 | !hmaster0_p & af3c26;
assign a5f8b7 = hlock1_p & a60172 | !hlock1_p & a5f8b6;
assign ce9cba = hgrant2_p & ce9cb9 | !hgrant2_p & !cea15c;
assign b29d21 = hbusreq2_p & b29d17 | !hbusreq2_p & v84563c;
assign a5fd16 = hgrant2_p & a5fd14 | !hgrant2_p & a5fd15;
assign a5fcc5 = hlock1_p & deac52 | !hlock1_p & deac53;
assign b29950 = hready & b2994d | !hready & c3b6a6;
assign deacb1 = hgrant2_p & deacae | !hgrant2_p & deacb0;
assign dead94 = hlock0_p & dead93 | !hlock0_p & !v84563c;
assign ab0580 = hbusreq2_p & ab057f | !hbusreq2_p & ab0572;
assign a5fc0d = hmastlock_p & a5fc0c | !hmastlock_p & !v84563c;
assign a5ee80 = hlock2_p & a5ee7f | !hlock2_p & a5ee08;
assign b2a015 = hbusreq2_p & b29f5a | !hbusreq2_p & b29cbb;
assign a5ee1b = hbusreq1_p & a5fc48 | !hbusreq1_p & v84563c;
assign ab055c = hgrant1_p & ab055b | !hgrant1_p & ab055a;
assign deadc7 = hbusreq2_p & deadc6 | !hbusreq2_p & v84563c;
assign a5f03c = decide_p & a5f03b | !decide_p & v84563c;
assign c3b871 = decide_p & c3b870 | !decide_p & v845660;
assign b29d30 = hbusreq2_p & b29d2f | !hbusreq2_p & v84563c;
assign ce9cb7 = hmaster0_p & ce9cb6 | !hmaster0_p & cea450;
assign a5f29a = hbusreq2 & a5fc91 | !hbusreq2 & !v84563c;
assign cea0f2 = hlock3_p & cea0d7 | !hlock3_p & cea0f1;
assign deacdd = locked_p & v84563c | !locked_p & !b26697;
assign a5f7f9 = hlock1_p & a5fbab | !hlock1_p & !a5f7f8;
assign ce9d54 = hbusreq2_p & ce9d53 | !hbusreq2_p & ce9d52;
assign b26729 = hlock1_p & v84563c | !hlock1_p & !b266da;
assign stateG3_1 = !a81d0d;
assign v845656 = hmaster0_p & v84563c | !hmaster0_p & !v84563c;
assign cea355 = hmaster0_p & cea354 | !hmaster0_p & cea2b3;
assign v970452 = decide_p & v970451 | !decide_p & v97044d;
assign b29ec9 = hbusreq2_p & b29ec8 | !hbusreq2_p & v84563c;
assign b29f1c = hlock1_p & b29f19 | !hlock1_p & b29f1b;
assign dea6f6 = hmaster0_p & dea6f3 | !hmaster0_p & !dea6f5;
assign cea3da = hgrant1_p & cea3d9 | !hgrant1_p & deae7f;
assign a5eecb = hgrant2_p & a5eeca | !hgrant2_p & v84563c;
assign deacf9 = hlock1_p & deacf7 | !hlock1_p & deacf8;
assign b8ace4 = locked_p & v84563c | !locked_p & b8ace3;
assign c3b801 = decide_p & c3b800 | !decide_p & v845660;
assign a5fc90 = hready & a5fc8c | !hready & a5fc8f;
assign deacf2 = hburst0_p & c07311 | !hburst0_p & deacf1;
assign ab0af9 = hlock1_p & v84563c | !hlock1_p & deacbd;
assign b29ed0 = hbusreq3 & b29ecf | !hbusreq3 & dead84;
assign b2672f = hbusreq2_p & b2672e | !hbusreq2_p & b2672d;
assign a5fc6f = hmaster1_p & v84563c | !hmaster1_p & a5fc6e;
assign b29d05 = hbusreq2_p & b29cf8 | !hbusreq2_p & !v84563c;
assign b29f6d = hmaster1_p & b29f68 | !hmaster1_p & b29f6c;
assign c3b77c = decide_p & c3b77b | !decide_p & v845660;
assign b2a019 = decide_p & b2a018 | !decide_p & !b29e57;
assign a5ea6e = hmaster0_p & a5ea4b | !hmaster0_p & a5ea6d;
assign c3bdda = hbusreq3 & c3bdd3 | !hbusreq3 & c3bdd9;
assign b29981 = hgrant2_p & b29980 | !hgrant2_p & !b29c3c;
assign b2a001 = hmaster0_p & b2a000 | !hmaster0_p & b29f93;
assign ab0637 = hbusreq2_p & ab0573 | !hbusreq2_p & ab0636;
assign b29f38 = hbusreq3 & b29f37 | !hbusreq3 & b29f35;
assign deaeb4 = hlock0_p & deaeb3 | !hlock0_p & v84563c;
assign deae56 = hbusreq3 & deae54 | !hbusreq3 & deae55;
assign c3bd4b = hready & c3bbd3 | !hready & cea887;
assign a5fa9e = hbusreq2_p & a5fa8c | !hbusreq2_p & a5fa8b;
assign a5f4e5 = hbusreq1_p & v9703fb | !hbusreq1_p & v84565a;
assign b29fca = hbusreq2_p & b29fc9 | !hbusreq2_p & v84563c;
assign a5fad2 = hbusreq0_p & a5fa2d | !hbusreq0_p & v84563c;
assign ab071c = hbusreq3 & ab071a | !hbusreq3 & ab071b;
assign a5f082 = hbusreq2_p & a5f081 | !hbusreq2_p & a5fb7b;
assign a5f582 = hlock0_p & a5f581 | !hlock0_p & a5f576;
assign deadf6 = decide_p & deadf5 | !decide_p & v84563c;
assign a5f511 = hbusreq2_p & a5f4f3 | !hbusreq2_p & a5f510;
assign a5ea92 = hbusreq0 & a5f0ab | !hbusreq0 & v84563c;
assign a5fa0e = stateG10_1_p & v970408 | !stateG10_1_p & a60187;
assign d40d3b = stateG10_1_p & d40d3a | !stateG10_1_p & !d40d33;
assign a5fa5f = hlock0_p & a5fa5d | !hlock0_p & a5fa5e;
assign b29d0f = hbusreq2_p & b29d0e | !hbusreq2_p & !b29d0d;
assign a5f56b = hlock1_p & a6016f | !hlock1_p & !a5f56a;
assign a5f211 = hmaster0_p & a5f20a | !hmaster0_p & a5f210;
assign a5f7ba = hready & v84563c | !hready & !ab0aee;
assign a5f23c = hbusreq2_p & a5f23b | !hbusreq2_p & v84563c;
assign c3bcd7 = hgrant3_p & c3bcbf | !hgrant3_p & !c3bcd6;
assign a5f72f = hbusreq3 & a5f72e | !hbusreq3 & v84563c;
assign af3493 = hgrant2_p & af348a | !hgrant2_p & af3492;
assign a5ef38 = hbusreq2 & a5ee13 | !hbusreq2 & a5ef37;
assign c3bccc = hbusreq2_p & c3bcc8 | !hbusreq2_p & c3bc0d;
assign b29e50 = hbusreq2_p & b29e4f | !hbusreq2_p & v84563c;
assign a5f942 = hlock1_p & a60193 | !hlock1_p & a5f941;
assign b29959 = hlock2_p & v84563c | !hlock2_p & !b29943;
assign a5f51b = hready & a5f515 | !hready & a5f51a;
assign c3bc72 = hlock0_p & b26697 | !hlock0_p & c3bc4d;
assign a5f9c6 = hbusreq3 & a601a6 | !hbusreq3 & a5f9c5;
assign a5eefa = hlock3_p & a5eef9 | !hlock3_p & a5ede4;
assign b29fb5 = locked_p & b29fb4 | !locked_p & c3bcdb;
assign cea411 = hgrant2_p & cea406 | !hgrant2_p & cea410;
assign d40d77 = hmaster1_p & d40d31 | !hmaster1_p & d40d47;
assign b2982e = hlock1_p & dead7b | !hlock1_p & b2982d;
assign ce9d6e = hbusreq2_p & cea297 | !hbusreq2_p & cea296;
assign a5f28b = decide_p & a5f25a | !decide_p & a5f28a;
assign a5ee19 = hlock2_p & a5ee15 | !hlock2_p & a5ee18;
assign a5f020 = hbusreq0 & a5fae7 | !hbusreq0 & a5f01f;
assign a5f43b = hbusreq1_p & a5fa1d | !hbusreq1_p & v84563c;
assign b29ff9 = hmaster0_p & b29ff5 | !hmaster0_p & !b29ff8;
assign c3b6a0 = hlock1_p & v84565a | !hlock1_p & v84563c;
assign deac4b = hburst1_p & v8c6449 | !hburst1_p & v84563c;
assign b29f86 = hlock0_p & b29ecc | !hlock0_p & c3bcdb;
assign a5edce = hlock2 & a5edcd | !hlock2 & a5f36e;
assign dea75e = hbusreq2_p & deadfa | !hbusreq2_p & v84563c;
assign cea2f3 = hlock2_p & cea2f2 | !hlock2_p & !cea17a;
assign v97042f = decide_p & v97042e | !decide_p & v9703ff;
assign ce9e23 = hgrant2_p & ce9d26 | !hgrant2_p & ce9e22;
assign ab0c22 = hbusreq2_p & ab0c21 | !hbusreq2_p & v84563c;
assign a5f968 = hmaster1_p & a5f962 | !hmaster1_p & a5f967;
assign ab0bff = locked_p & ab0bfe | !locked_p & !v84563c;
assign ab0649 = hlock3_p & ab0642 | !hlock3_p & ab0648;
assign b299ad = hlock2_p & v84563c | !hlock2_p & !b29991;
assign cea3a9 = hbusreq0_p & cea37b | !hbusreq0_p & !cea38d;
assign a5f3c6 = hbusreq1_p & b26695 | !hbusreq1_p & v84563c;
assign b26747 = hbusreq2_p & b266a8 | !hbusreq2_p & !b26695;
assign b8ace6 = hmaster1_p & b8ace5 | !hmaster1_p & !v84563c;
assign a5fc65 = hmaster0_p & a5fc59 | !hmaster0_p & a5fc64;
assign dea758 = hgrant2_p & deadf0 | !hgrant2_p & dea757;
assign deae2d = decide_p & deae2c | !decide_p & !v84563c;
assign ab0b60 = hlock2_p & ab0b5f | !hlock2_p & dead2e;
assign a5eef6 = hbusreq3 & a5eef4 | !hbusreq3 & !a5eef5;
assign cea8a1 = hbusreq2_p & cea89d | !hbusreq2_p & cea89c;
assign ab0ca0 = hgrant2_p & ab0b70 | !hgrant2_p & ab0c9f;
assign a5f727 = hready & a5fb71 | !hready & !b266a0;
assign a5faaf = hlock1_p & a60177 | !hlock1_p & !a5faae;
assign cea861 = hlock3_p & cea860 | !hlock3_p & v84563c;
assign a5e9c1 = hlock1_p & a5fbab | !hlock1_p & !a5e9c0;
assign b26779 = hlock2_p & b26736 | !hlock2_p & b266ae;
assign c3b7d1 = hlock2_p & c3b7cc | !hlock2_p & !c3b7d0;
assign cea387 = hbusreq3 & cea37f | !hbusreq3 & cea386;
assign a5fb6f = stateA1_p & v8e1935 | !stateA1_p & v84563c;
assign c3b84c = hbusreq2_p & c3b84b | !hbusreq2_p & !c3b84a;
assign a5f293 = hlock2_p & a5f292 | !hlock2_p & v84563c;
assign cea183 = hready_p & cea181 | !hready_p & cea182;
assign deac56 = hgrant1_p & deac54 | !hgrant1_p & deac55;
assign deae0f = hbusreq2_p & deae0e | !hbusreq2_p & dead39;
assign b29f77 = hgrant1_p & b29ee9 | !hgrant1_p & b29f76;
assign c3bdcf = hready & c3bd5c | !hready & c3bdce;
assign adaecd = hbusreq2_p & adaecc | !hbusreq2_p & v84563c;
assign v970444 = hbusreq1_p & v9703fc | !hbusreq1_p & v97043e;
assign c3b718 = hbusreq2_p & c3b717 | !hbusreq2_p & !c3b6a8;
assign a5fb6b = locked_p & v84563c | !locked_p & a5fb6a;
assign a5fc08 = start_p & a6016a | !start_p & a5fbdf;
assign dea6e4 = hmaster0_p & dea6e3 | !hmaster0_p & deae6d;
assign c3bdf7 = hready_p & c3bdea | !hready_p & c3bdf6;
assign cea192 = hmaster1_p & cea15d | !hmaster1_p & cea191;
assign b266da = stateG10_1_p & b26693 | !stateG10_1_p & b266a1;
assign c3bc83 = hgrant2_p & c3bc78 | !hgrant2_p & c3bc82;
assign d40d47 = hgrant2_p & d40d45 | !hgrant2_p & d40d46;
assign b29ab0 = hlock2 & b29aad | !hlock2 & b29aaf;
assign deac61 = hbusreq2_p & deac5d | !hbusreq2_p & deac5c;
assign b29fa3 = hlock2_p & b29f9b | !hlock2_p & !b29fa2;
assign a5efa9 = hlock0_p & a5fbc0 | !hlock0_p & a5ee68;
assign c3b68e = hbusreq3 & c3b68c | !hbusreq3 & c3b68d;
assign cea409 = hlock1_p & deac51 | !hlock1_p & !cea408;
assign a5f734 = hbusreq2_p & a5f733 | !hbusreq2_p & v84563c;
assign cea8ad = hlock2_p & cea8ac | !hlock2_p & v84563c;
assign v970431 = hlock0_p & v9703fd | !hlock0_p & v84563c;
assign ab0746 = hlock0_p & b29f99 | !hlock0_p & !ab0745;
assign a5f6df = hmaster0_p & a5f6da | !hmaster0_p & a5f6de;
assign cea0f0 = hmaster1_p & cea0e9 | !hmaster1_p & cea0ef;
assign c3bd36 = start_p & v845652 | !start_p & !c3bd35;
assign a5fbc3 = hlock2_p & a5fbc2 | !hlock2_p & v84563c;
assign deacc4 = hgrant2_p & deacc0 | !hgrant2_p & deacc3;
assign cea0b5 = hbusreq3 & cea8ae | !hbusreq3 & cea86e;
assign a5f924 = hbusreq2 & a5f91a | !hbusreq2 & a5f923;
assign b8acf0 = hready_p & b8acee | !hready_p & b8acef;
assign ab0640 = hgrant2_p & ab0b2d | !hgrant2_p & ab0b30;
assign bdb59a = hmaster0_p & bdb599 | !hmaster0_p & !bdb598;
assign ab05a6 = hlock2 & ab0d03 | !hlock2 & ab05a5;
assign b29923 = hbusreq1_p & v84563c | !hbusreq1_p & !deadba;
assign b29cea = hlock2 & b29ce7 | !hlock2 & b29ce9;
assign b2a007 = hgrant2_p & b29e95 | !hgrant2_p & !b29fa4;
assign a5f472 = hready & a5f46f | !hready & a5f471;
assign b26756 = hmastlock_p & b2669e | !hmastlock_p & v84563c;
assign deae03 = hbusreq1_p & v84563c | !hbusreq1_p & deae02;
assign a5efd5 = hbusreq3 & a5efd2 | !hbusreq3 & a5efd4;
assign a5f2fe = hbusreq2 & a5fc71 | !hbusreq2 & v84563c;
assign cea460 = hlock0_p & cea38e | !hlock0_p & !cea38d;
assign b29a4b = hbusreq2_p & b29a4a | !hbusreq2_p & v84563c;
assign c3b8b6 = hready_p & c3b896 | !hready_p & c3b8b5;
assign b298a3 = hbusreq2_p & b298a2 | !hbusreq2_p & v84563c;
assign c3b77a = hgrant0_p & dead2e | !hgrant0_p & c3b779;
assign ab074d = decide_p & ab074c | !decide_p & v845662;
assign b29d65 = hlock0_p & b29d51 | !hlock0_p & !v84563c;
assign c3b70b = hbusreq2_p & c3b70a | !hbusreq2_p & !c3b656;
assign a5f0a4 = hbusreq0 & a5f0a3 | !hbusreq0 & v84563c;
assign deae8a = hbusreq2_p & deae7a | !hbusreq2_p & deae79;
assign a5efca = hgrant2_p & a5efc9 | !hgrant2_p & v84563c;
assign a5eb6f = hbusreq2_p & a5f198 | !hbusreq2_p & a5f199;
assign b2999e = hlock0_p & b2999d | !hlock0_p & !b29986;
assign a9b9ed = decide_p & bdb581 | !decide_p & a9b9d2;
assign a5fb99 = hlock0_p & a5fb98 | !hlock0_p & a5fb92;
assign a5f6d1 = hbusreq2_p & a5f6d0 | !hbusreq2_p & v84563c;
assign c3b7bd = hlock0_p & c3bd17 | !hlock0_p & !deadb2;
assign dead83 = hbusreq3 & dead79 | !hbusreq3 & dead82;
assign a5ef51 = hlock1_p & v84565a | !hlock1_p & a5ef50;
assign b29952 = hlock2 & b2994f | !hlock2 & b29951;
assign c3bdfb = hlock2_p & c3bdfa | !hlock2_p & dead2e;
assign c3b6a8 = hready & c3b6a7 | !hready & deada8;
assign a5ee5f = locked_p & a5ee5e | !locked_p & v845641;
assign a60147 = decide_p & a60146 | !decide_p & v84563c;
assign a5f1ce = hmaster1_p & a5f1c4 | !hmaster1_p & a5f1cd;
assign a5ede1 = hbusreq0 & a5eddf | !hbusreq0 & a5ede0;
assign af34ce = hmaster1_p & af349d | !hmaster1_p & af34a1;
assign ab054e = hlock2_p & ab054c | !hlock2_p & ab054d;
assign af3c5d = locked_p & d40d33 | !locked_p & af3c4e;
assign deae08 = hbusreq2_p & deae07 | !hbusreq2_p & v845660;
assign a5ea90 = hbusreq2 & a5f0ab | !hbusreq2 & a5ea8f;
assign b2a00e = hready & deac7a | !hready & !v84563c;
assign c3b6cf = hbusreq2_p & c3b6cd | !hbusreq2_p & c3b6cc;
assign a5f9a2 = hready & a5fbdd | !hready & b2672b;
assign a9b9e4 = hgrant2_p & v84563c | !hgrant2_p & !a9b9d0;
assign a5fc95 = hbusreq3 & a5fc94 | !hbusreq3 & v84563c;
assign a5f8dc = start_p & a5f8d8 | !start_p & !a5f8db;
assign ab0c61 = hbusreq2_p & ab0c60 | !hbusreq2_p & ab0b23;
assign af3c7f = hlock1_p & af3c49 | !hlock1_p & !d40d41;
assign a5f108 = hbusreq0_p & a5f82c | !hbusreq0_p & ab0c31;
assign dea6df = hlock0_p & dea6de | !hlock0_p & !v84563c;
assign b29f05 = hburst0 & deacb3 | !hburst0 & b29f04;
assign a5f8d7 = hlock0_p & a5f8d6 | !hlock0_p & v84563c;
assign deadd6 = hlock0_p & deadd5 | !hlock0_p & !v84563c;
assign b29f87 = hlock2_p & b29f86 | !hlock2_p & dead2e;
assign a5f1e7 = hbusreq2 & a5f1e4 | !hbusreq2 & !a5f1e6;
assign ab0c73 = hgrant2_p & ab0c71 | !hgrant2_p & ab0c72;
assign a5ef46 = hmaster1_p & a5ef45 | !hmaster1_p & !v84563c;
assign a5ef8c = hbusreq2_p & a5eddc | !hbusreq2_p & a5ef8b;
assign a5fb5d = hbusreq0_p & a5fb2a | !hbusreq0_p & v84563c;
assign b29cba = decide_p & b29cb9 | !decide_p & v84563c;
assign deae79 = hlock0_p & deae76 | !hlock0_p & !deadb2;
assign ab0c12 = hmaster1_p & ab0c0d | !hmaster1_p & ab0c11;
assign ab05cf = hlock0_p & v84563c | !hlock0_p & ab05b0;
assign b29d7c = hlock0_p & b29d79 | !hlock0_p & !b29d7b;
assign adaedd = hmaster1_p & v84563c | !hmaster1_p & adaedc;
assign ab0c8b = locked_p & c3bd8b | !locked_p & !v84563c;
assign c3b852 = hmaster1_p & c3b851 | !hmaster1_p & c3b7e0;
assign deac72 = hlock2_p & deac71 | !hlock2_p & deac52;
assign ab0bdf = hready_p & ab0bcd | !hready_p & ab0bde;
assign c3bdc7 = hbusreq2_p & c3bdc6 | !hbusreq2_p & v845660;
assign ab05ee = hlock0_p & v84563c | !hlock0_p & !ab05ed;
assign a5f268 = hbusreq2 & a5fccb | !hbusreq2 & v84563c;
assign af3503 = hmaster0_p & af3502 | !hmaster0_p & af34cb;
assign a5ea5b = hbusreq0_p & a5fc5e | !hbusreq0_p & v84563c;
assign cea467 = hmaster0_p & cea45f | !hmaster0_p & cea466;
assign d40d72 = hbusreq2_p & d40d2c | !hbusreq2_p & d40d68;
assign b29978 = hready_p & b29910 | !hready_p & b29977;
assign stateA1 = b2678e;
assign ab0cb4 = hgrant2_p & ab0bba | !hgrant2_p & ab0c93;
assign dea6d5 = hbusreq2_p & dea6d1 | !hbusreq2_p & dea6d0;
assign a6019b = hlock2_p & a6018d | !hlock2_p & a6019a;
assign b26758 = hbusreq0_p & b26699 | !hbusreq0_p & !b26757;
assign a5f547 = hlock2_p & a5f538 | !hlock2_p & a5f546;
assign a5fcfd = hlock1_p & deac52 | !hlock1_p & deac54;
assign a5f3b6 = hbusreq2_p & a5f3b2 | !hbusreq2_p & a5f3b5;
assign b29abb = locked_p & b29aba | !locked_p & !v84563c;
assign ab0639 = hmaster1_p & ab0634 | !hmaster1_p & !ab0638;
assign deadcb = hgrant2_p & deadc8 | !hgrant2_p & deadca;
assign c3be00 = locked_p & v84563c | !locked_p & c3bdff;
assign a5fc76 = stateA1_p & v84563c | !stateA1_p & !a5fc75;
assign adaef7 = hmaster1_p & adaef6 | !hmaster1_p & v84563c;
assign b29e4d = locked_p & b29e4c | !locked_p & v84563c;
assign b29914 = hbusreq1_p & v84563c | !hbusreq1_p & !deaca1;
assign c07311 = stateG3_1_p & v845670 | !stateG3_1_p & !v845670;
assign b299a4 = hgrant2_p & b299a3 | !hgrant2_p & !b29c3c;
assign a5eed3 = hmaster1_p & a5eed0 | !hmaster1_p & a5eed2;
assign cea29d = hgrant1_p & deac52 | !hgrant1_p & deac55;
assign a5f536 = hready & a5f531 | !hready & a5f535;
assign b29d54 = hlock2_p & v84563c | !hlock2_p & b29d53;
assign a5ee4b = hbusreq1 & a5fbd9 | !hbusreq1 & v84563c;
assign a5fce3 = hmastlock_p & a5fce2 | !hmastlock_p & v84563c;
assign c3b7f5 = hlock1_p & c3bbd2 | !hlock1_p & c3b7f4;
assign ab0c88 = hmaster1_p & ab0c84 | !hmaster1_p & ab0c87;
assign dea733 = hlock0_p & deae30 | !hlock0_p & v84563c;
assign b266cb = hbusreq1_p & b266ca | !hbusreq1_p & b26693;
assign af356a = hbusreq2_p & af355f | !hbusreq2_p & af352c;
assign ce9d2c = hbusreq2_p & cea297 | !hbusreq2_p & cea366;
assign c3bdb2 = hlock2_p & c3bdb1 | !hlock2_p & !c3bca0;
assign ce9cd2 = hlock3_p & ce9cd1 | !hlock3_p & cea18a;
assign a5f300 = hmaster1_p & a5f2ff | !hmaster1_p & a5f751;
assign b29ffc = locked_p & v84563c | !locked_p & !c3bdf8;
assign dea6f4 = hgrant2_p & deacd3 | !hgrant2_p & deacd5;
assign af34e9 = hgrant2_p & af3c50 | !hgrant2_p & af3c70;
assign a5f1db = hbusreq2_p & a5f1da | !hbusreq2_p & v84563c;
assign dea74c = hbusreq3 & dea74b | !hbusreq3 & deae40;
assign cea38e = locked_p & v84563c | !locked_p & !cea38d;
assign ab0628 = hlock2_p & ab056b | !hlock2_p & ab0564;
assign c3bd7a = hready & c3bd79 | !hready & deada8;
assign b29b5f = jx1_p & b29b36 | !jx1_p & b29a21;
assign deae5d = hlock2_p & deae5c | !hlock2_p & !v84563c;
assign a5faeb = hmaster0_p & a5f9cb | !hmaster0_p & a5faea;
assign ab05ff = hmaster1_p & ab05f8 | !hmaster1_p & ab05fe;
assign cea150 = hbusreq1_p & deae02 | !hbusreq1_p & v84563c;
assign c3bd2d = hready & cea26f | !hready & c3bd2c;
assign b29cdd = hready & deadac | !hready & !v84563c;
assign c3b888 = decide_p & c3b887 | !decide_p & !v845660;
assign a5edc6 = hlock1_p & a5fa1c | !hlock1_p & a5f4cc;
assign b29f5f = hmaster0_p & b29f47 | !hmaster0_p & !b29f5e;
assign deae94 = hlock1_p & v84565a | !hlock1_p & !c98b95;
assign a5f70e = hbusreq2 & a5f70d | !hbusreq2 & !v84563c;
assign ab05d4 = hmaster0_p & ab05c9 | !hmaster0_p & ab05d3;
assign a5f0ac = hbusreq0_p & a5fc71 | !hbusreq0_p & v84563c;
assign c3bc18 = hbusreq2_p & c3bc17 | !hbusreq2_p & !c3bc16;
assign a5fcac = hbusreq3 & a5fcab | !hbusreq3 & v84563c;
assign b266c1 = hbusreq2_p & b266a8 | !hbusreq2_p & b266ae;
assign b29d63 = hmaster0_p & b29d57 | !hmaster0_p & b29d62;
assign dea6f8 = decide_p & dea6f7 | !decide_p & v84563c;
assign v8c6711 = hlock1_p & v84563c | !hlock1_p & v845646;
assign a5ea45 = hlock0_p & a5ea44 | !hlock0_p & a5ea40;
assign a5eae7 = hready & a5f11b | !hready & a5f837;
assign a5f084 = hbusreq2_p & a5f083 | !hbusreq2_p & a5fbc1;
assign a5f334 = hmaster1_p & a5f6db | !hmaster1_p & a5f333;
assign ab0b51 = hready_p & ab0ad0 | !hready_p & ab0b50;
assign deae35 = hbusreq2_p & dead8f | !hbusreq2_p & v845644;
assign cea340 = hgrant3_p & cea2b7 | !hgrant3_p & cea33f;
assign cea238 = hbusreq3 & cea237 | !hbusreq3 & v84563c;
assign af34b6 = hmastlock_p & af3c4a | !hmastlock_p & !v84563c;
assign c3b6e9 = hbusreq2_p & c3b6e8 | !hbusreq2_p & !c3b625;
assign c3b721 = hlock2_p & c3b720 | !hlock2_p & !c3b71f;
assign b29f96 = hlock2_p & b29f95 | !hlock2_p & v845660;
assign c3bdb7 = hbusreq2_p & c3bdb6 | !hbusreq2_p & v845660;
assign ab0b32 = hgrant2_p & ab0b2e | !hgrant2_p & ab0b31;
assign a5f4a5 = hlock1_p & a60168 | !hlock1_p & a5f4a4;
assign a5f4fb = hbusreq1 & a5f4fa | !hbusreq1 & !v84563c;
assign c3bc44 = hlock3_p & c3bc2f | !hlock3_p & !c3bc43;
assign ab0c98 = locked_p & ab0c97 | !locked_p & !v84563c;
assign dea76e = hlock3_p & v84563c | !hlock3_p & dea76d;
assign d40d5a = hmaster1_p & d40d59 | !hmaster1_p & d40d54;
assign ab05da = hgrant3_p & ab0587 | !hgrant3_p & !ab05d9;
assign c3bdd5 = hready & cea331 | !hready & c3bdd4;
assign ab05f7 = hbusreq2_p & ab0560 | !hbusreq2_p & ab05f5;
assign cea3f9 = hlock0_p & cea3f8 | !hlock0_p & cea3cd;
assign a5f1cb = hbusreq2 & a5f1c8 | !hbusreq2 & a5f1ca;
assign a5f07e = hlock0_p & a5f71e | !hlock0_p & v84563c;
assign c3b7ea = hlock0_p & c3b613 | !hlock0_p & !v84563c;
assign ab0b69 = hbusreq2_p & ab0b68 | !hbusreq2_p & ab0b66;
assign a5eaf5 = hmaster1_p & a5eaf4 | !hmaster1_p & a5f163;
assign a5f047 = jx1_p & a5f014 | !jx1_p & a5f046;
assign cea334 = hready & cea331 | !hready & cea333;
assign a5f4ea = hready & a5f4e4 | !hready & a5f4e9;
assign a5fc2b = hbusreq2 & a5fc2a | !hbusreq2 & a5fc29;
assign af3533 = hlock0_p & v84563c | !hlock0_p & af3532;
assign a5f90a = hlock2_p & a5f909 | !hlock2_p & v84563c;
assign a5edca = hbusreq2 & a5edc2 | !hbusreq2 & a5edc9;
assign a5fcc0 = hgrant2_p & a5fcbe | !hgrant2_p & a5fcbf;
assign a5ea2e = hmaster0_p & a5ea26 | !hmaster0_p & a5ea2d;
assign a5f08e = hbusreq3 & a5f08d | !hbusreq3 & v84563c;
assign a5edd1 = hbusreq2_p & a5edcb | !hbusreq2_p & a5edd0;
assign ab05ba = hmaster0_p & ab05a0 | !hmaster0_p & ab05b9;
assign ab073d = hmaster0_p & ab073b | !hmaster0_p & ab073c;
assign a5fc4e = hmaster0_p & v84563c | !hmaster0_p & a5fc4d;
assign c3b774 = hmaster0_p & c3b773 | !hmaster0_p & c3bcd3;
assign deac2a = hbusreq3 & deac20 | !hbusreq3 & v84563c;
assign ab0c1e = hbusreq2_p & ab0c1d | !hbusreq2_p & v84563c;
assign d40d6c = hmaster0_p & v84563c | !hmaster0_p & d40d6b;
assign c3b7a4 = hmaster1_p & c3b79f | !hmaster1_p & c3b7a3;
assign c3bdaf = hready & c3bdae | !hready & !dead6e;
assign a5ea30 = hready_p & a5f0b1 | !hready_p & a5ea2f;
assign ab0bae = hlock0_p & b29ecc | !hlock0_p & v845660;
assign a5f958 = hbusreq2_p & a5f957 | !hbusreq2_p & v84563c;
assign a5edba = hbusreq2 & a5edac | !hbusreq2 & a5edb9;
assign ab0cdf = hbusreq2_p & ab0c6d | !hbusreq2_p & v845644;
assign a5efdd = hbusreq2_p & a5f4f3 | !hbusreq2_p & a5ef79;
assign a81caf = stateG2_p & v84563c | !stateG2_p & !v845672;
assign a5eb83 = hmaster0_p & a5eb76 | !hmaster0_p & a5eb82;
assign a5f83f = hmastlock_p & a5f83e | !hmastlock_p & v84563c;
assign a5fbc2 = hbusreq2 & a60142 | !hbusreq2 & a5fbc1;
assign a5f718 = hbusreq2 & a5f717 | !hbusreq2 & v84563c;
assign c3bc21 = hlock0_p & v84565a | !hlock0_p & !v84563c;
assign ab0bf6 = decide_p & ab0bf5 | !decide_p & !v845662;
assign a81ce4 = hgrant2_p & v84563c | !hgrant2_p & a81ce3;
assign af357f = hlock1_p & af352c | !hlock1_p & af357e;
assign c3bcc5 = hlock0_p & cea29f | !hlock0_p & !v84563c;
assign c3bc8d = hbusreq2_p & b266a8 | !hbusreq2_p & c3bc8c;
assign a5f55b = hbusreq0_p & a5f4ee | !hbusreq0_p & a5f4fc;
assign a5fa5d = hready & a60168 | !hready & a5f9f9;
assign deae8f = hmaster0_p & deae8e | !hmaster0_p & !v84563c;
assign b29aaf = hlock0_p & b29aae | !hlock0_p & !dead77;
assign ab0cd7 = hbusreq2_p & ab0c21 | !hbusreq2_p & v845644;
assign ab05ac = hlock2 & ab05aa | !hlock2 & ab05ab;
assign c3bc29 = hbusreq3 & c3bc18 | !hbusreq3 & c3bc28;
assign b29926 = hlock1_p & c3b683 | !hlock1_p & !b29925;
assign ab0bc8 = hready_p & ab0bc6 | !hready_p & !ab0bc7;
assign a5f13b = hbusreq0 & a5f13a | !hbusreq0 & !ab0c31;
assign c3b873 = hgrant3_p & c3b802 | !hgrant3_p & c3b872;
assign a5ee77 = hlock0_p & v845641 | !hlock0_p & a5ee76;
assign a9b9d9 = locked_p & c3b6a0 | !locked_p & !v84563c;
assign ab0b8b = hlock2 & ab0b88 | !hlock2 & ab0b8a;
assign a5fa67 = hlock0_p & a5fa65 | !hlock0_p & !a5fa66;
assign cea2b1 = hbusreq2_p & cea2b0 | !hbusreq2_p & !deacaa;
assign b29ae8 = hbusreq3 & b29d20 | !hbusreq3 & b29ae7;
assign a5fbeb = hlock1_p & a5f9dd | !hlock1_p & v84563c;
assign dead6e = hmastlock_p & dead6d | !hmastlock_p & !v84563c;
assign ab0b3f = hbusreq3 & v84563c | !hbusreq3 & ab0b3e;
assign b2676b = hmaster0_p & b2676a | !hmaster0_p & !b266bd;
assign a81cc8 = locked_p & a81cb1 | !locked_p & v84563c;
assign cea163 = hlock2_p & cea162 | !hlock2_p & !dead72;
assign a5f457 = hbusreq1 & a5f456 | !hbusreq1 & v84563c;
assign a5f6fa = hready & v84563c | !hready & !dead33;
assign a5f373 = hbusreq2_p & a5f372 | !hbusreq2_p & a5f36d;
assign ab05c7 = hbusreq2_p & ab05c6 | !hbusreq2_p & ab059c;
assign a5f590 = hlock2_p & a5f58d | !hlock2_p & a5f58f;
assign dead97 = hbusreq3 & dead96 | !hbusreq3 & !v84563c;
assign b29ecc = locked_p & v84563c | !locked_p & !c3bc47;
assign dea789 = hgrant2_p & dea785 | !hgrant2_p & dea788;
assign dead5f = hgrant2_p & deacad | !hgrant2_p & deacaf;
assign b26698 = locked_p & b26693 | !locked_p & !b26697;
assign ab059f = hgrant2_p & ab059e | !hgrant2_p & cea15a;
assign a5f8f5 = hbusreq0 & a5f8f3 | !hbusreq0 & !a5f8f4;
assign c3bd81 = decide_p & c3bd80 | !decide_p & v845660;
assign b29ccb = hbusreq2_p & b29cca | !hbusreq2_p & !b29cc9;
assign a5ee67 = hlock2 & a5ee13 | !hlock2 & a5ee66;
assign ce9cc8 = hbusreq3 & ce9cc6 | !hbusreq3 & ce9cc7;
assign af3c54 = hbusreq1_p & d40d33 | !hbusreq1_p & af3c4c;
assign a5ee6e = hlock0_p & a60141 | !hlock0_p & a5ee6d;
assign a5eb2a = hbusreq2 & a5ea27 | !hbusreq2 & a5ea8f;
assign af3c2c = locked_p & v84563c | !locked_p & v8c6711;
assign a5f328 = hbusreq2 & a5f321 | !hbusreq2 & v845641;
assign a5fb82 = locked_p & v84563c | !locked_p & a5fb81;
assign dea6c7 = hlock3_p & v84563c | !hlock3_p & dea6c6;
assign a5fcf7 = hbusreq1_p & v84563c | !hbusreq1_p & !a5fcd7;
assign b29943 = hlock0_p & b29942 | !hlock0_p & !v84563c;
assign ab0b10 = hbusreq3 & ab0b0d | !hbusreq3 & ab0b0f;
assign af3494 = hmaster1_p & af3493 | !hmaster1_p & af348e;
assign a5eeda = hready & a5f520 | !hready & a5f3f7;
assign c3bc5a = hlock0_p & cea341 | !hlock0_p & deacdf;
assign a5f78e = hlock0_p & a5f787 | !hlock0_p & a5f78d;
assign c3bc4c = hlock0_p & b2669d | !hlock0_p & !deace1;
assign a81cce = hmaster1_p & v84563c | !hmaster1_p & a81ccd;
assign c3bce2 = hlock2_p & c3bce1 | !hlock2_p & !dead7f;
assign b266b9 = hmaster1_p & b266b8 | !hmaster1_p & b266a2;
assign a5f171 = hbusreq0_p & a5f9e8 | !hbusreq0_p & a5fa2d;
assign cea449 = hbusreq2_p & cea445 | !hbusreq2_p & cea448;
assign c3bbf2 = hbusreq2_p & c3bbea | !hbusreq2_p & c3bbe8;
assign a5ea81 = hready & a5fc09 | !hready & a5fc0d;
assign cea1a8 = hgrant3_p & cea18c | !hgrant3_p & cea1a7;
assign b2675e = locked_p & b2675d | !locked_p & b2672b;
assign a5ee87 = hlock0_p & a5ee86 | !hlock0_p & a5ee14;
assign deadb3 = hlock0_p & deadac | !hlock0_p & !deadb2;
assign af3489 = hlock2_p & af3c7b | !hlock2_p & d40d33;
assign cea48d = hlock3_p & cea48c | !hlock3_p & cea43f;
assign a81cde = hlock0_p & a81caa | !hlock0_p & a81cdd;
assign cea46b = hmaster1_p & cea46a | !hmaster1_p & cea178;
assign a5ea3f = hbusreq0 & a5ea3b | !hbusreq0 & a5ea3e;
assign c3bc97 = hbusreq3 & c3bc93 | !hbusreq3 & c3bc96;
assign c3b827 = hlock2_p & c3b826 | !hlock2_p & !c3b7ab;
assign ab0586 = decide_p & ab0585 | !decide_p & v84563c;
assign deae48 = decide_p & deae47 | !decide_p & v84563c;
assign a5fcef = locked_p & v845641 | !locked_p & !v84563c;
assign a5f1eb = hmaster1_p & v84563c | !hmaster1_p & a5f1ea;
assign a5ea3a = hlock2_p & a5fbd3 | !hlock2_p & a5ea39;
assign cea45f = hmaster1_p & cea444 | !hmaster1_p & v84563c;
assign ab0606 = hbusreq0_p & b298aa | !hbusreq0_p & cea44a;
assign a5f3d9 = hbusreq2_p & a5f3d2 | !hbusreq2_p & a5f3d8;
assign a5f73e = hbusreq3 & a5f73d | !hbusreq3 & v84563c;
assign ab0519 = hbusreq0_p & b298a0 | !hbusreq0_p & b299d7;
assign deae21 = hgrant1_p & deadba | !hgrant1_p & deadbc;
assign a5ea17 = hlock2_p & a5ea16 | !hlock2_p & a5f196;
assign ce9ddc = decide_p & ce9ddb | !decide_p & v84563c;
assign af3546 = stateG10_1_p & v84563c | !stateG10_1_p & af352e;
assign a5f880 = hready & a5f87c | !hready & !a5f87f;
assign a5f9a0 = hready & a5fbdd | !hready & !b26729;
assign b29f68 = hgrant2_p & b29f64 | !hgrant2_p & b29f67;
assign a5f295 = hbusreq3 & a5f294 | !hbusreq3 & v84563c;
assign b2673f = hmaster1_p & b26738 | !hmaster1_p & !b2673e;
assign ab0bd4 = hlock0_p & v84563c | !hlock0_p & b29e67;
assign b29b1c = hlock0_p & c3bcef | !hlock0_p & v84563c;
assign a5f955 = hbusreq2_p & a5f954 | !hbusreq2_p & !v84563c;
assign a5fab3 = hlock0_p & a5fab2 | !hlock0_p & v84563c;
assign a5f2f3 = hlock0_p & a5f2f2 | !hlock0_p & a5f728;
assign c3b778 = hmaster1_p & c3bca4 | !hmaster1_p & c3b703;
assign a60176 = start_p & a81ca6 | !start_p & a60175;
assign a5f965 = hbusreq2 & a5f964 | !hbusreq2 & a5fb7b;
assign a5f2ca = hmaster1_p & a5f2c9 | !hmaster1_p & a5f926;
assign deace2 = hlock0_p & deacdd | !hlock0_p & deace1;
assign af34dc = hlock2_p & af3c64 | !hlock2_p & af3c4c;
assign ab0715 = hlock0_p & b29fd9 | !hlock0_p & !b29fdc;
assign a5fc47 = start_p & v845654 | !start_p & !a5fc46;
assign a5ee2c = hlock1_p & a5fbae | !hlock1_p & !a5ee1e;
assign a5f74e = hbusreq2_p & a5f74d | !hbusreq2_p & !v84563c;
assign a5edf1 = hready & a5edee | !hready & a5edf0;
assign af3c37 = hmaster0_p & af3c36 | !hmaster0_p & af3c35;
assign af3c6c = hmaster1_p & af3c6b | !hmaster1_p & af3c4c;
assign a5fd39 = hmaster0_p & v84563c | !hmaster0_p & a5fd38;
assign c3b7aa = hmaster0_p & c3b7a4 | !hmaster0_p & c3b7a9;
assign b29ab7 = hmaster1_p & b29ab6 | !hmaster1_p & b29d64;
assign deadbd = hgrant1_p & deadbb | !hgrant1_p & deadbc;
assign ab0b2d = hbusreq2_p & ab0b24 | !hbusreq2_p & ab0b23;
assign b29faa = hgrant0_p & b29f94 | !hgrant0_p & !b29fa9;
assign af34c3 = hbusreq2_p & af34b0 | !hbusreq2_p & af3c4c;
assign c3b844 = hlock0_p & c3bdd0 | !hlock0_p & deada8;
assign a5f8d5 = hlock1_p & a60177 | !hlock1_p & !a5f8d4;
assign cea474 = hmaster0_p & cea46b | !hmaster0_p & cea473;
assign a5f3d0 = hbusreq3 & a5f3c9 | !hbusreq3 & !a5f3cf;
assign ab0cdb = hbusreq3 & ab0cda | !hbusreq3 & v84564a;
assign ce9d5a = hlock3_p & ce9d51 | !hlock3_p & ce9d59;
assign cea24f = hburst0 & cea24d | !hburst0 & cea24e;
assign a5f577 = hlock0_p & a5f575 | !hlock0_p & !a5f576;
assign a5f6ce = hgrant0_p & a60144 | !hgrant0_p & a5fbc5;
assign a5eeb3 = hmaster0_p & a5ee9a | !hmaster0_p & a5eeb2;
assign c3b6ed = hbusreq2_p & c3b6ec | !hbusreq2_p & !c3b6e0;
assign cea89f = hbusreq3 & cea88d | !hbusreq3 & cea89e;
assign b29fab = hlock0_p & c3bcf8 | !hlock0_p & c3bcdb;
assign a5f4cf = hlock1_p & a60177 | !hlock1_p & !a5f4ce;
assign a5f7fa = hbusreq1_p & a5fa1d | !hbusreq1_p & !a60177;
assign a5ee1d = hbusreq1 & a5ee1c | !hbusreq1 & !v84563c;
assign ab0bef = hmaster1_p & ab0bed | !hmaster1_p & ab0bee;
assign ab0c01 = hlock2_p & ab0bfd | !hlock2_p & ab0c00;
assign deac9d = hgrant2_p & deac9a | !hgrant2_p & deac9c;
assign deadb4 = hlock2_p & deadb3 | !hlock2_p & !deadb2;
assign c3b656 = hlock0_p & c3b625 | !hlock0_p & c3b655;
assign deae41 = hbusreq2_p & deadd7 | !hbusreq2_p & v845644;
assign ab0602 = hready_p & ab05ec | !hready_p & ab0601;
assign a5f2d5 = hmaster1_p & a5fd28 | !hmaster1_p & a5f2d4;
assign a5f321 = hlock0_p & a5f320 | !hlock0_p & ab0c31;
assign deae46 = hmaster1_p & dead63 | !hmaster1_p & !deae45;
assign a5ee70 = hbusreq0_p & a5fbc0 | !hbusreq0_p & a5ee68;
assign ab062e = hbusreq2_p & ab0628 | !hbusreq2_p & ab062d;
assign a5eee1 = hlock1_p & a5fbab | !hlock1_p & !a5f434;
assign dead35 = hlock0_p & dead34 | !hlock0_p & v84563c;
assign b29edf = hmaster0_p & b29eda | !hmaster0_p & b29ede;
assign a5e9da = hbusreq2_p & a5e9d5 | !hbusreq2_p & a5e9d4;
assign b29eb0 = hlock2 & b29eaa | !hlock2 & b29eaf;
assign cea199 = hbusreq2_p & cea198 | !hbusreq2_p & !v84563c;
assign cea889 = hlock2_p & cea888 | !hlock2_p & !cea887;
assign b29f61 = hbusreq2_p & b29f60 | !hbusreq2_p & !v84563c;
assign ab0599 = hlock0_p & b298a4 | !hlock0_p & ab0598;
assign a5eea0 = hlock2 & a5ee9d | !hlock2 & a5ee9f;
assign ce9cc1 = hlock2_p & ce9cc0 | !hlock2_p & !cea405;
assign c3b7b7 = decide_p & c3b7b6 | !decide_p & v845660;
assign af35aa = hmaster1_p & af352c | !hmaster1_p & af352f;
assign b2994b = hlock2 & b29948 | !hlock2 & b2994a;
assign a5ea8b = hmaster1_p & a5ea8a | !hmaster1_p & v84563c;
assign af3586 = hmaster1_p & af3585 | !hmaster1_p & af3533;
assign af35a8 = decide_p & af35a7 | !decide_p & af3576;
assign cea442 = hready_p & cea3af | !hready_p & cea441;
assign cea286 = hlock2_p & cea283 | !hlock2_p & !cea887;
assign ab0527 = hmaster1_p & ab0526 | !hmaster1_p & v84563c;
assign a5e9e6 = hbusreq0 & a5e9e1 | !hbusreq0 & a5f15c;
assign d40d2a = start_p & v84563c | !start_p & d40d29;
assign b29d6d = hlock1_p & dead6e | !hlock1_p & b29d6c;
assign a5fb7e = hbusreq3 & a5fb78 | !hbusreq3 & a5fb7d;
assign a5edee = hbusreq1 & a5eded | !hbusreq1 & !v84563c;
assign a5eec3 = hready & a5eec0 | !hready & a5eec2;
assign ab06e7 = hlock0_p & ab06e6 | !hlock0_p & !dead34;
assign a5f3ef = hbusreq1_p & a60168 | !hbusreq1_p & v84563c;
assign a5ebc3 = hbusreq0 & a5ebc2 | !hbusreq0 & v845641;
assign b29f3c = hready & deac57 | !hready & v84563c;
assign a5fb7d = hbusreq2_p & a5fb7c | !hbusreq2_p & a5fb7b;
assign ab0c58 = hgrant2_p & ab0b03 | !hgrant2_p & ab0b0f;
assign dead47 = hbusreq3 & dead46 | !hbusreq3 & !dead39;
assign d40d64 = hready_p & d40d2e | !hready_p & d40d63;
assign deacbd = hgrant1_p & v84563c | !hgrant1_p & deacbc;
assign ab056d = hbusreq2_p & ab0560 | !hbusreq2_p & ab056c;
assign b26770 = hmaster0_p & b2676f | !hmaster0_p & !b26705;
assign a5f7bc = hbusreq2 & a5f7a4 | !hbusreq2 & a5f7bb;
assign a5f82b = hlock1_p & a5f828 | !hlock1_p & a5f82a;
assign a5ea0d = hbusreq2 & a5ea07 | !hbusreq2 & a5ea06;
assign a5f973 = hlock1_p & v84563c | !hlock1_p & !a5fb8d;
assign a5e9eb = hmaster1_p & a5e9dd | !hmaster1_p & a5e9ea;
assign a5f39a = hbusreq2_p & a5f399 | !hbusreq2_p & a5f395;
assign a5fa6f = hbusreq2_p & a5fa56 | !hbusreq2_p & a5fa6e;
assign b29f8e = hlock2 & b29f8d | !hlock2 & b29ecd;
assign bdb5a1 = hgrant0_p & bdb59e | !hgrant0_p & bdb5a0;
assign a5ee60 = hlock0_p & a5ee59 | !hlock0_p & !a5ee5f;
assign a5f071 = hlock0_p & a5f06f | !hlock0_p & a5f070;
assign a5f099 = hmaster1_p & a5f092 | !hmaster1_p & a5f098;
assign cea265 = start_p & deac4a | !start_p & !v84563c;
assign c3bcf6 = hmaster1_p & c3bbbf | !hmaster1_p & c3bcf5;
assign a5ee26 = hready & a5ee25 | !hready & !v84563c;
assign b29d5c = hready & dead6e | !hready & !deae02;
assign a5efbf = hlock0_p & a5ee38 | !hlock0_p & a5efbe;
assign af34a4 = hmaster1_p & af349f | !hmaster1_p & af34a3;
assign hgrant0 = !ab076c;
assign deadfe = hlock2_p & deadfd | !hlock2_p & v84563c;
assign b29f54 = hready & b29f53 | !hready & v84563c;
assign a9b9d1 = hmaster1_p & a9b9d0 | !hmaster1_p & !v84563c;
assign deac5a = hgrant1_p & deac54 | !hgrant1_p & deac53;
assign a5fc8d = stateA1_p & v845652 | !stateA1_p & !v845654;
assign ab0676 = hbusreq2_p & ab0675 | !hbusreq2_p & ab0b80;
assign dea6fb = hlock3_p & v84563c | !hlock3_p & dea6fa;
assign ab0bb4 = hmaster1_p & ab0b9a | !hmaster1_p & ab0bb3;
assign a5efb5 = hmaster1_p & a5efb4 | !hmaster1_p & a5fbc5;
assign a81cd6 = hgrant2_p & a81cd5 | !hgrant2_p & v84563c;
assign b29fa6 = hmaster1_p & b29f98 | !hmaster1_p & b29fa5;
assign af358d = hgrant2_p & af352d | !hgrant2_p & af3531;
assign c3b807 = hlock2_p & c3bc75 | !hlock2_p & !c3b7ad;
assign ab0684 = hbusreq2_p & ab0683 | !hbusreq2_p & !b29b1c;
assign b2997d = hlock0_p & b2997c | !hlock0_p & !v84563c;
assign ab06ad = stateG10_1_p & deacb3 | !stateG10_1_p & deaca0;
assign ab0738 = hlock0_p & b29f3d | !hlock0_p & !ab0737;
assign a5fa60 = hlock2 & a5fa5c | !hlock2 & a5fa5f;
assign c3b80b = hlock2_p & c3b809 | !hlock2_p & !c3b80a;
assign ab0c9a = hready & ab0c96 | !hready & dead40;
assign cea486 = hbusreq3 & cea47e | !hbusreq3 & cea485;
assign cea418 = hgrant2_p & cea416 | !hgrant2_p & cea417;
assign a5edd8 = hlock1_p & v84565a | !hlock1_p & b29929;
assign c3bdbe = hready & c3bdbc | !hready & c3bdbd;
assign c3b813 = hbusreq2_p & c3b811 | !hbusreq2_p & !c3b812;
assign deadd5 = hlock1_p & v84565a | !hlock1_p & !deadd4;
assign bdb5a8 = hmaster1_p & bdb5a7 | !hmaster1_p & !bdb598;
assign b29ee6 = hburst1 & b29ee5 | !hburst1 & v84563c;
assign be34df = hgrant2_p & v84563c | !hgrant2_p & v84564a;
assign a5f93d = hbusreq2_p & a5f93c | !hbusreq2_p & a5fad6;
assign a5f188 = hgrant1_p & a5fa0e | !hgrant1_p & a5f187;
assign a5ea39 = hbusreq2 & a5f094 | !hbusreq2 & a5fbc6;
assign a5f369 = hready & a5f365 | !hready & !a5f368;
assign b26745 = hmaster1_p & b26744 | !hmaster1_p & !b26718;
assign a5f197 = hlock2_p & a5f194 | !hlock2_p & a5f196;
assign a5f570 = hgrant1_p & a5f56e | !hgrant1_p & a5f56f;
assign a5eb3b = hgrant2_p & a5eb38 | !hgrant2_p & a5eb3a;
assign b29ea1 = decide_p & b29ea0 | !decide_p & b29e57;
assign ab0c7e = hmaster1_p & ab0c73 | !hmaster1_p & ab0c7d;
assign c3bcbc = hmaster1_p & c3bc36 | !hmaster1_p & c3bc21;
assign b29aa3 = hlock0_p & deace1 | !hlock0_p & !v84563c;
assign a5ef07 = hbusreq1 & a5ef06 | !hbusreq1 & !v84563c;
assign ce9db8 = hbusreq3 & ce9db7 | !hbusreq3 & v84563c;
assign b2993f = hlock2 & b2993b | !hlock2 & b2993e;
assign b29830 = hlock1_p & dead7b | !hlock1_p & !b2982f;
assign a5f521 = hready & a5f520 | !hready & a5f4a7;
assign a5f305 = hgrant0_p & a5f301 | !hgrant0_p & a5f304;
assign ce9d34 = hbusreq2_p & cea2b0 | !hbusreq2_p & cea887;
assign af350f = hgrant3_p & af34ff | !hgrant3_p & af350e;
assign a5ef86 = hlock0_p & a5f581 | !hlock0_p & a5f36e;
assign a5fc58 = hgrant2_p & v84563c | !hgrant2_p & a5fc57;
assign a5f599 = hgrant2_p & a5f595 | !hgrant2_p & a5f598;
assign c3b67a = hgrant1_p & c3b679 | !hgrant1_p & deae7f;
assign c3bca8 = hlock2_p & dead77 | !hlock2_p & v84563c;
assign a5fca1 = hbusreq1 & a5fc9e | !hbusreq1 & !a5fca0;
assign a5f01c = hlock2_p & a5fa37 | !hlock2_p & v845644;
assign a5f1d4 = hlock0_p & a5f1d3 | !hlock0_p & a5fc2c;
assign cea357 = hready_p & cea348 | !hready_p & cea356;
assign a5f526 = hlock0_p & a5f521 | !hlock0_p & a5f525;
assign ab0571 = hlock0_p & ab056f | !hlock0_p & ab0570;
assign ab06a3 = hlock0_p & b29f3d | !hlock0_p & !deaca2;
assign a5ea64 = hlock2 & a5f1a2 | !hlock2 & a5fbc1;
assign ab0ae0 = hbusreq2_p & ab0adf | !hbusreq2_p & ab0ade;
assign a5f09f = hbusreq3 & a5f09e | !hbusreq3 & v84563c;
assign c3b661 = hbusreq1_p & deada8 | !hbusreq1_p & c3b660;
assign a5f3a6 = hlock2_p & a5f3a2 | !hlock2_p & a5f3a5;
assign a5ef33 = hgrant3_p & a5ee04 | !hgrant3_p & a5ef32;
assign b29a42 = hbusreq2_p & b29a41 | !hbusreq2_p & v84563c;
assign ab06ca = hready & ab06c9 | !hready & v84563c;
assign a5fc46 = stateA1_p & v84566e | !stateA1_p & a5f9da;
assign a5eb46 = hgrant0_p & v84563c | !hgrant0_p & a5eb45;
assign c3b7ff = hmaster0_p & c3b7f0 | !hmaster0_p & c3b7fe;
assign cea177 = hgrant0_p & cea158 | !hgrant0_p & cea176;
assign a5f45a = hbusreq1 & a5f459 | !hbusreq1 & v84565a;
assign a5f066 = locked_p & a5f6fa | !locked_p & v84563c;
assign dea7b4 = jx0_p & dea701 | !jx0_p & dea7b3;
assign c3b6ab = hlock0_p & c3bbe2 | !hlock0_p & !c3b6a1;
assign v970421 = hbusreq2_p & v970420 | !hbusreq2_p & v84563c;
assign a5fb8d = hbusreq1_p & a5fb8c | !hbusreq1_p & dead6e;
assign a5f3cf = locked_p & a5f3ce | !locked_p & v84563c;
assign ab06bb = hready & ab06ba | !hready & v84563c;
assign d40d80 = hbusreq1_p & d40d31 | !hbusreq1_p & d40d7b;
assign a5f434 = hbusreq1_p & a5f828 | !hbusreq1_p & v84563c;
assign b29994 = hlock0_p & b29993 | !hlock0_p & !v84563c;
assign a5f1a3 = hbusreq0_p & v84563c | !hbusreq0_p & ab0c31;
assign b29fe6 = hmaster1_p & b29fe5 | !hmaster1_p & b29f46;
assign ce9cbc = hmaster0_p & ce9cbb | !hmaster0_p & cea45c;
assign af34b4 = hbusreq2_p & af34b3 | !hbusreq2_p & af3c4c;
assign a5fc7e = hready & a5fc7d | !hready & b2982c;
assign a5eecd = hbusreq2 & a5f3c9 | !hbusreq2 & !a5f3cf;
assign dea6ce = hgrant1_p & deadba | !hgrant1_p & deae7f;
assign a5fa1a = hgrant1_p & a5fa0e | !hgrant1_p & a60187;
assign deacf8 = hbusreq1_p & v84563c | !hbusreq1_p & deacf7;
assign cea3fa = hlock1_p & deac52 | !hlock1_p & !v845646;
assign a5ef93 = hmaster0_p & a5ef92 | !hmaster0_p & !a5ee01;
assign deac20 = hbusreq2_p & deac1f | !hbusreq2_p & v84565a;
assign c3b79c = hlock0_p & c3bce0 | !hlock0_p & dead7f;
assign a5e9d7 = hbusreq0 & a5e9d6 | !hbusreq0 & v845641;
assign a60146 = hlock3_p & a60145 | !hlock3_p & v84563c;
assign ce9cc9 = hgrant2_p & ce9cc5 | !hgrant2_p & ce9cc8;
assign a5ee55 = hbusreq1_p & v9703fc | !hbusreq1_p & v84563c;
assign deaea7 = hbusreq2_p & deaea3 | !hbusreq2_p & deaea2;
assign v8e1935 = hburst0_p & v84563c | !hburst0_p & v845654;
assign a5ea7c = hlock0_p & a5ea7b | !hlock0_p & a5ea4e;
assign cea267 = hburst0 & v84563c | !hburst0 & cea266;
assign a5fd3a = decide_p & a5fd39 | !decide_p & v84563c;
assign ab05e0 = hbusreq2_p & ab0524 | !hbusreq2_p & ab05df;
assign a5f53e = hlock0_p & a5f4ee | !hlock0_p & a5f53d;
assign c3bd86 = hlock0_p & c3bc52 | !hlock0_p & !c3bce5;
assign b2a013 = hgrant2_p & b2a011 | !hgrant2_p & b2a012;
assign c3be02 = hlock2_p & c3be01 | !hlock2_p & v845660;
assign b8acdc = hlock1_p & v84563c | !hlock1_p & b8acdb;
assign deadc5 = hlock0_p & deadbe | !hlock0_p & !deadc4;
assign ab0b0e = hlock0_p & ab0adc | !hlock0_p & !v84563c;
assign b26735 = locked_p & v84563c | !locked_p & b26734;
assign ab0bde = decide_p & ab0bdd | !decide_p & v84563c;
assign a5fc0b = hlock1_p & a5fba2 | !hlock1_p & a5fc0a;
assign a5f248 = hready & a5f247 | !hready & a5f7fc;
assign a5ee99 = hgrant2_p & a5ee98 | !hgrant2_p & v84563c;
assign a5fd09 = hbusreq2_p & a5fd05 | !hbusreq2_p & !a5fd08;
assign c3bd9d = hlock2_p & c3bd9c | !hlock2_p & !cea17a;
assign a5ea3d = hlock2_p & a5fbc1 | !hlock2_p & a5ea3c;
assign ab058d = hlock0_p & ab0b5e | !hlock0_p & !cea38d;
assign ab0c8a = hlock0_p & ab0b64 | !hlock0_p & ab0c89;
assign cea19a = hlock2_p & cea0bf | !hlock2_p & !v84563c;
assign ab06cb = hlock0_p & ab06ca | !hlock0_p & !ab068c;
assign af3c61 = hbusreq2_p & af3c60 | !hbusreq2_p & af3c4c;
assign b840ac = hmaster1_p & v84564f | !hmaster1_p & v845647;
assign dea76f = decide_p & dea76e | !decide_p & v84563c;
assign b29f1e = hlock0_p & b29f10 | !hlock0_p & b29f1d;
assign be34e7 = hgrant0_p & v84564a | !hgrant0_p & be34df;
assign a5f8be = hlock1_p & a60172 | !hlock1_p & a5f8bd;
assign a81cb0 = start_p & v84563c | !start_p & a81caf;
assign a5ee73 = hbusreq0_p & a5ee38 | !hbusreq0_p & a5ee65;
assign b2a017 = hmaster1_p & b29e9e | !hmaster1_p & !b2a016;
assign b8acdf = hmaster1_p & b8acdc | !hmaster1_p & !v84563c;
assign a5ea54 = hbusreq0_p & a5fc5c | !hbusreq0_p & v84563c;
assign af3c23 = hmaster1_p & af3c20 | !hmaster1_p & af3c22;
assign a5fc18 = hlock2 & v84563c | !hlock2 & a5fc17;
assign a81d06 = hmaster1_p & a81cf1 | !hmaster1_p & v84563c;
assign ce9cc2 = hbusreq2_p & ce9cc1 | !hbusreq2_p & !cea405;
assign dea79e = hgrant3_p & dea75d | !hgrant3_p & !dea79d;
assign b299ac = hgrant3_p & b29978 | !hgrant3_p & b299ab;
assign a5fb9c = hbusreq2_p & a5fb9b | !hbusreq2_p & a5fb93;
assign b29f34 = hlock2_p & b29f1e | !hlock2_p & !b29f33;
assign b2677d = hmaster0_p & b2677c | !hmaster0_p & !b2673f;
assign a5f56d = hbusreq1_p & v9703fb | !hbusreq1_p & !deadb9;
assign cea249 = hmastlock_p & cea248 | !hmastlock_p & v84566c;
assign deadfb = hbusreq2_p & deadfa | !hbusreq2_p & v845660;
assign ab0b4a = hbusreq2_p & ab0b46 | !hbusreq2_p & ab0b45;
assign a5ee7a = hbusreq2_p & a5ee79 | !hbusreq2_p & a5ee78;
assign b29fba = hbusreq2_p & b29fb9 | !hbusreq2_p & v84563c;
assign a5fc8c = hmastlock_p & a5fc8b | !hmastlock_p & !v84563c;
assign dead7c = hbusreq1_p & dead7b | !hbusreq1_p & !v84563c;
assign dea6c3 = hgrant2_p & dea6c2 | !hgrant2_p & dead3b;
assign a5f1d2 = hready & a5f1d1 | !hready & !a5fb8c;
assign c3b6cc = hlock0_p & c3b6cb | !hlock0_p & c3b6af;
assign dead89 = hbusreq1_p & v84563c | !hbusreq1_p & !b26695;
assign ab0cad = locked_p & c3bdaf | !locked_p & !v84563c;
assign cea41c = hlock0_p & cea41b | !hlock0_p & cea3fb;
assign ab053e = hlock0_p & ab053d | !hlock0_p & !b2991b;
assign cea29e = hlock1_p & v84563c | !hlock1_p & !cea29d;
assign bfbd19 = stateG3_1_p & v84563c | !stateG3_1_p & bfbd18;
assign a5fd00 = locked_p & a5fcfc | !locked_p & a5fcff;
assign b29999 = hmaster0_p & b29982 | !hmaster0_p & b29998;
assign b29d07 = hgrant2_p & b29cfc | !hgrant2_p & b29d06;
assign a5ef88 = hbusreq0 & a5ef85 | !hbusreq0 & a5ef87;
assign c3b749 = hmaster1_p & c3b6a1 | !hmaster1_p & !deacaa;
assign a5ef6c = hlock0_p & a5f4f0 | !hlock0_p & a5ef6b;
assign b29aa5 = hlock2_p & v845660 | !hlock2_p & b29aa4;
assign ab0cec = hlock2_p & ab0ceb | !hlock2_p & v84563c;
assign c3bde2 = hready_p & c3bdcd | !hready_p & c3bde1;
assign c3bc70 = hbusreq2_p & c3bc6f | !hbusreq2_p & c3bc6e;
assign a5f828 = start_p & v8e1935 | !start_p & !c06d34;
assign a5f976 = hlock0_p & a5f975 | !hlock0_p & a5f72b;
assign d40d3c = hbusreq1_p & d40d33 | !hbusreq1_p & v84563c;
assign a5f085 = hbusreq0 & a5f082 | !hbusreq0 & a5f084;
assign a5f936 = hbusreq1_p & v84563c | !hbusreq1_p & deac52;
assign ab06b0 = hready & deacb7 | !hready & ab06af;
assign b299a3 = hbusreq2_p & b299a2 | !hbusreq2_p & b29995;
assign b299e2 = hgrant2_p & b299e1 | !hgrant2_p & !b29c3c;
assign a5f861 = hlock1_p & a60172 | !hlock1_p & deac56;
assign b2677b = hgrant2_p & b26778 | !hgrant2_p & b2677a;
assign dea6fa = hgrant0_p & dead2d | !hgrant0_p & dead3c;
assign v970457 = decide_p & v84563c | !decide_p & v970456;
assign ab071e = hmaster1_p & ab071d | !hmaster1_p & ab06a7;
assign cea422 = hbusreq2_p & cea421 | !hbusreq2_p & cea405;
assign b2998c = locked_p & deae59 | !locked_p & b2997c;
assign ab0510 = hlock0_p & b298a4 | !hlock0_p & b298a0;
assign b29eb5 = hburst1 & dead7a | !hburst1 & b29eb4;
assign af3c29 = decide_p & af3c28 | !decide_p & v8567b4;
assign b299de = hlock0_p & b29992 | !hlock0_p & v84563c;
assign ab0be4 = hbusreq2_p & cea15a | !hbusreq2_p & cea18f;
assign b299e7 = hmaster0_p & b299d3 | !hmaster0_p & !b29957;
assign ab0bc6 = decide_p & ab0bc5 | !decide_p & v845662;
assign a5f122 = hbusreq2 & a5f110 | !hbusreq2 & a5f121;
assign ab0cb9 = hmaster0_p & ab0cb6 | !hmaster0_p & ab0cb8;
assign a5fc13 = locked_p & a5fc12 | !locked_p & v845641;
assign ab0c64 = hmaster1_p & ab0c58 | !hmaster1_p & !ab0c63;
assign a5f20a = hmaster1_p & a5f209 | !hmaster1_p & a5f751;
assign b29f50 = hlock1_p & deac51 | !hlock1_p & b29ee9;
assign ab0552 = hbusreq2_p & ab054e | !hbusreq2_p & ab054c;
assign a5fad4 = hbusreq0_p & v845641 | !hbusreq0_p & v84563c;
assign ab0c9c = hlock0_p & v84563c | !hlock0_p & !ab0c9b;
assign b29f46 = hgrant2_p & b29f44 | !hgrant2_p & b29f45;
assign a5f844 = hlock0_p & a5f83c | !hlock0_p & a5f843;
assign a5f213 = hbusreq2 & a5fcab | !hbusreq2 & v84563c;
assign b29eb4 = start_p & cea1aa | !start_p & b29eb3;
assign b29953 = hlock2_p & b29952 | !hlock2_p & b29943;
assign c3b7f4 = hgrant1_p & c3bd12 | !hgrant1_p & c3bd77;
assign af3c3a = decide_p & af3c39 | !decide_p & v8567b4;
assign cea39d = locked_p & deae59 | !locked_p & !cea39c;
assign a5ea76 = hlock2_p & a5ea75 | !hlock2_p & a5ea46;
assign a5fba7 = hbusreq1_p & a5fba6 | !hbusreq1_p & a5fba2;
assign a5f1f8 = hlock0_p & a5f1f7 | !hlock0_p & v84563c;
assign a5eb70 = hbusreq0 & a5eb6f | !hbusreq0 & v845641;
assign deadaa = hbusreq1_p & deada8 | !hbusreq1_p & !deac51;
assign deadde = hmastlock_p & deaca0 | !hmastlock_p & v84566c;
assign af3c5e = locked_p & d40d33 | !locked_p & af3c4c;
assign ab06f6 = hgrant2_p & ab06f2 | !hgrant2_p & ab06f5;
assign a5f3bc = hbusreq2 & a5f3ba | !hbusreq2 & a5f3bb;
assign c3bd02 = hlock0_p & c3bcdb | !hlock0_p & c3bd01;
assign cea376 = hlock1_p & v84563c | !hlock1_p & !cea374;
assign a5f2dc = hmaster1_p & a5f2db | !hmaster1_p & !a5f958;
assign a5ee0d = hbusreq2_p & a5ee09 | !hbusreq2_p & a5ee0c;
assign a9b9de = hgrant2_p & a9b9dd | !hgrant2_p & !v84563c;
assign dea6dc = hready_p & dea6c8 | !hready_p & !dea6db;
assign ab0d02 = jx0_p & ab0bf9 | !jx0_p & ab0d01;
assign a60175 = stateA1_p & a60174 | !stateA1_p & !v8c6449;
assign ab0b8c = hlock0_p & v84563c | !hlock0_p & !deace9;
assign a5f4ce = hgrant1_p & a5f4cd | !hgrant1_p & a5f4cc;
assign cea436 = hlock2_p & cea435 | !hlock2_p & cea3fb;
assign c3bcd9 = hready & cea1b3 | !hready & c3bc61;
assign ab05e7 = hlock0_p & b29832 | !hlock0_p & ab05e6;
assign a5f6d6 = hbusreq2_p & a5f6d2 | !hbusreq2_p & a5fa6d;
assign af349e = hlock2_p & af349c | !hlock2_p & af349d;
assign v970450 = hmaster0_p & v97044f | !hmaster0_p & v97042a;
assign ab076c = jx2_p & ab0d02 | !jx2_p & ab076b;
assign ab0c44 = hlock0_p & v84563c | !hlock0_p & ab0c43;
assign ab0b90 = hlock0_p & v84563c | !hlock0_p & !b29d88;
assign b299d6 = hready_p & b299cc | !hready_p & b299d5;
assign af3c49 = hmastlock_p & af3c48 | !hmastlock_p & v84563c;
assign a5eadd = hlock2_p & a5eadb | !hlock2_p & a5eadc;
assign c3bd8d = locked_p & v84563c | !locked_p & !c3bcef;
assign af34ac = hlock2_p & af3c5f | !hlock2_p & af3c4c;
assign b29cfe = hready & deada8 | !hready & v84563c;
assign cea47b = hready & cea47a | !hready & cea40a;
assign b29ed1 = hmaster1_p & b29c3d | !hmaster1_p & b29ed0;
assign af34c2 = hbusreq2_p & af34c1 | !hbusreq2_p & af3c6b;
assign af359d = hmaster1_p & af359c | !hmaster1_p & af3574;
assign b29b0f = hmaster1_p & b29b0e | !hmaster1_p & b29a50;
assign dea6ed = decide_p & dea6ec | !decide_p & v84563c;
assign d40d87 = hgrant2_p & d40d86 | !hgrant2_p & d40d60;
assign a5eb35 = hgrant2_p & a5eb2b | !hgrant2_p & a5eb34;
assign a81ce3 = locked_p & a81ce2 | !locked_p & v84563c;
assign a5f555 = hgrant1_p & a5f3f5 | !hgrant1_p & b29914;
assign a5eb37 = hbusreq2 & a5ea24 | !hbusreq2 & a5eb36;
assign c3b805 = hbusreq2_p & c3b7a5 | !hbusreq2_p & c3bc94;
assign v845660 = locked_p & v84563c | !locked_p & !v84563c;
assign b8ace0 = hmaster0_p & b8acdf | !hmaster0_p & b8acdc;
assign a5fbff = hlock0_p & a5fbfc | !hlock0_p & a5fbfe;
assign a5f58f = hbusreq2 & a5f4ee | !hbusreq2 & a5f58e;
assign deac71 = hlock0_p & deac6c | !hlock0_p & deac52;
assign a5f073 = hlock2_p & a5f071 | !hlock2_p & a5f072;
assign a5fcdf = locked_p & a5fcde | !locked_p & v84563c;
assign a5f3f2 = hlock1_p & a60168 | !hlock1_p & a5f3f1;
assign a5ee02 = hmaster0_p & a5edf4 | !hmaster0_p & a5ee01;
assign adaf1b = hgrant3_p & adaf18 | !hgrant3_p & adaf1a;
assign bdb5ba = hbusreq3_p & bdb5ad | !hbusreq3_p & bdb5b9;
assign b266af = hlock0_p & b266ad | !hlock0_p & b266ae;
assign c3b717 = hlock2_p & c3b716 | !hlock2_p & !c3b6a8;
assign ab075b = hmaster0_p & ab0759 | !hmaster0_p & ab075a;
assign bdb5b8 = hready_p & bdb5a2 | !hready_p & !bdb5b7;
assign b26721 = hlock0_p & b26720 | !hlock0_p & b266a8;
assign cea0bc = hlock1_p & v84563c | !hlock1_p & !cea0bb;
assign dea6bf = hbusreq2_p & deaeb0 | !hbusreq2_p & v84563c;
assign c3b876 = hmaster1_p & c3b7b3 | !hmaster1_p & c3bcb4;
assign c3bd98 = hready & dead0a | !hready & !v84563c;
assign cea0be = hbusreq2_p & cea0b9 | !hbusreq2_p & cea0bd;
assign a5ef34 = hlock0_p & a5ee83 | !hlock0_p & a5ee13;
assign dead04 = hlock0_p & deacdd | !hlock0_p & deace3;
assign adaf11 = hgrant3_p & adaedb | !hgrant3_p & adaf10;
assign b29cbb = hlock0_p & v84565a | !hlock0_p & v84563c;
assign a5efde = hlock0_p & a5fa6c | !hlock0_p & a5ef5e;
assign a5ea1c = hmaster1_p & a5ea1a | !hmaster1_p & a5ea1b;
assign c3b7d6 = hbusreq3 & c3b7d4 | !hbusreq3 & c3b7d5;
assign a5f8c0 = hlock0_p & a5f8bf | !hlock0_p & v845641;
assign deae59 = hlock1_p & v84563c | !hlock1_p & !v845646;
assign a5f98c = locked_p & a5f98b | !locked_p & !v845641;
assign af354f = hbusreq2_p & af354e | !hbusreq2_p & af354c;
assign a5e9ae = hbusreq0 & a5f19a | !hbusreq0 & a5e9ad;
assign b2671e = hbusreq2_p & b2671d | !hbusreq2_p & !b26695;
assign c3bd71 = hlock2_p & c3bd4b | !hlock2_p & cea887;
assign deadf4 = hmaster0_p & deade5 | !hmaster0_p & !deadf3;
assign dead19 = locked_p & v84563c | !locked_p & !dead18;
assign a5efc6 = hgrant0_p & a5efa5 | !hgrant0_p & a5efc5;
assign af35be = hgrant0_p & af35bb | !hgrant0_p & af35bd;
assign ab0b0a = hready & deadde | !hready & ab0aeb;
assign a5eea8 = hbusreq2 & a5eea0 | !hbusreq2 & !a5eea7;
assign a5eb51 = hbusreq3 & a5eb4f | !hbusreq3 & a5eb50;
assign a5f56f = hbusreq1_p & v9703fb | !hbusreq1_p & !deadba;
assign a81cf0 = hmastlock_p & a81cef | !hmastlock_p & v84563c;
assign a5ef76 = hmaster1_p & a5ef75 | !hmaster1_p & v84563c;
assign dead51 = hready_p & dead4f | !hready_p & !dead50;
assign ab0c5a = hgrant1_p & c3b660 | !hgrant1_p & ab0c59;
assign ab0cc4 = hlock0_p & v84563c | !hlock0_p & ab0cc3;
assign deae66 = hlock2_p & deae65 | !hlock2_p & !v84563c;
assign a5f092 = hbusreq3 & a5f089 | !hbusreq3 & v84563c;
assign a5eaec = hbusreq0 & a5eaeb | !hbusreq0 & !ab0c31;
assign adaece = hlock2_p & adaec4 | !hlock2_p & v84563c;
assign bdb599 = hmaster1_p & v84565a | !hmaster1_p & !bdb598;
assign c3b88b = hlock2_p & c3b7a6 | !hlock2_p & c3b7b1;
assign b8ace5 = hgrant2_p & v8c6711 | !hgrant2_p & b8ace4;
assign a5fbd4 = hlock2_p & a5fbd3 | !hlock2_p & v84563c;
assign cea17e = hmaster0_p & cea17d | !hmaster0_p & cea178;
assign ab066c = hlock0_p & c3bcf8 | !hlock0_p & !ab066a;
assign a5f232 = hlock2 & a5f22e | !hlock2 & a5f231;
assign a5eb3f = hbusreq0_p & a5fce5 | !hbusreq0_p & !v84563c;
assign b266a3 = locked_p & v84563c | !locked_p & !b266a2;
assign b29cc8 = hlock1_p & deadde | !hlock1_p & deac5a;
assign ab0b01 = hlock2 & ab0afb | !hlock2 & ab0b00;
assign cea1aa = stateA1_p & v845652 | !stateA1_p & !v84563c;
assign c3bdba = hburst0 & v84566c | !hburst0 & c3bdb9;
assign ab0aef = hready & b29a5a | !hready & ab0aee;
assign a5f38b = hlock1_p & a5fb71 | !hlock1_p & v84563c;
assign a5f4ed = hbusreq1 & c3b697 | !hbusreq1 & v84563c;
assign b29f5d = hgrant2_p & b29f5b | !hgrant2_p & b29f5c;
assign cea328 = hbusreq2_p & cea327 | !hbusreq2_p & v845660;
assign a5fd0a = hbusreq3 & a5fd09 | !hbusreq3 & v84563c;
assign b2997a = hmaster1_p & b298a3 | !hmaster1_p & b29829;
assign c3b6c5 = hlock1_p & deada8 | !hlock1_p & c3b6c3;
assign a5ead2 = hlock0_p & a5ead0 | !hlock0_p & a5ead1;
assign v845646 = hbusreq1_p & v84563c | !hbusreq1_p & !v84563c;
assign ce9d72 = hmaster1_p & ce9d71 | !hmaster1_p & !ce9d28;
assign ab05f0 = hbusreq0_p & b29949 | !hbusreq0_p & b29946;
assign ab055e = hready & b29917 | !hready & ab055d;
assign a5f73d = hbusreq2_p & a5f73c | !hbusreq2_p & v84563c;
assign c3b71d = hlock1_p & c3b683 | !hlock1_p & deadba;
assign a5ef44 = hmaster0_p & a5ef43 | !hmaster0_p & a5f3c0;
assign a5fbf2 = hlock0_p & a5fbf1 | !hlock0_p & a5fbe9;
assign a5fca0 = hlock1_p & a5fc84 | !hlock1_p & a5fc9f;
assign c3b616 = hbusreq2_p & c3b615 | !hbusreq2_p & !v84563c;
assign a5f1bd = hbusreq2_p & a5f72d | !hbusreq2_p & v84563c;
assign b29d71 = hlock2_p & v84563c | !hlock2_p & !b29d70;
assign dea768 = hlock0_p & dea767 | !hlock0_p & v84563c;
assign cea37d = hlock0_p & cea379 | !hlock0_p & cea37c;
assign dead8c = hlock0_p & dead8b | !hlock0_p & !v84563c;
assign a5fcab = locked_p & a5fca7 | !locked_p & a5fcaa;
assign deaced = locked_p & v84563c | !locked_p & !deacec;
assign ab0cc5 = hlock2 & v84563c | !hlock2 & ab0cc4;
assign a5f54d = hbusreq2_p & a5f547 | !hbusreq2_p & a5f54c;
assign a5ea9c = hbusreq0_p & a5fc91 | !hbusreq0_p & !v84563c;
assign a5eb49 = hgrant3_p & a5ea30 | !hgrant3_p & a5eb48;
assign a5fbe1 = hmastlock_p & a5fbe0 | !hmastlock_p & v84563c;
assign c3b812 = hlock0_p & c3bd8d | !hlock0_p & v84563c;
assign dea7ab = decide_p & dea7aa | !decide_p & v84563c;
assign deae9c = hgrant2_p & deae98 | !hgrant2_p & deae9b;
assign b266b2 = hlock0_p & b2669d | !hlock0_p & b266b1;
assign b29962 = hmaster1_p & b29961 | !hmaster1_p & b29e65;
assign a5eff9 = hmaster0_p & a5eff8 | !hmaster0_p & a5ef17;
assign c3b685 = hlock1_p & deadb9 | !hlock1_p & deadc3;
assign b2992e = hbusreq2_p & b2992d | !hbusreq2_p & !b2992c;
assign a5f37f = locked_p & a5f37e | !locked_p & v845641;
assign b29988 = hready & deae4e | !hready & c3b622;
assign a5ef62 = hbusreq2_p & a5ef5a | !hbusreq2_p & a5ef61;
assign b29b20 = hbusreq2_p & b29b1f | !hbusreq2_p & !b29b1e;
assign b29ab8 = hmaster0_p & b29aac | !hmaster0_p & b29ab7;
assign c3bbfa = hgrant1_p & c3bbf6 | !hgrant1_p & c3bbd2;
assign cea336 = hlock2_p & cea335 | !hlock2_p & v84563c;
assign a5f395 = hlock0_p & a60141 | !hlock0_p & a5f394;
assign c3b74f = hmaster1_p & c3b74e | !hmaster1_p & c3bc5e;
assign b29a41 = hlock2_p & v84563c | !hlock2_p & b29a40;
assign c3b645 = hmaster1_p & c3b63e | !hmaster1_p & c3b644;
assign c3b734 = hmaster1_p & c3b733 | !hmaster1_p & c3bcb4;
assign a81cc4 = hmaster0_p & a81cb6 | !hmaster0_p & a81cc3;
assign ab0700 = hmaster1_p & ab06ff | !hmaster1_p & ab0bbb;
assign b29fd3 = hlock0_p & b29f57 | !hlock0_p & b29fd2;
assign a5f1ae = hbusreq1 & v84563c | !hbusreq1 & a5f1ad;
assign a5eee7 = hbusreq1_p & a5f455 | !hbusreq1_p & v84563c;
assign locked = c3b8cc;
assign cea493 = hmaster0_p & cea492 | !hmaster0_p & cea3ac;
assign af3585 = hgrant2_p & af3584 | !hgrant2_p & af3531;
assign ab050f = hmaster1_p & ab050e | !hmaster1_p & ab0ace;
assign a5fa00 = hready & a5f9f6 | !hready & v84565a;
assign v970413 = hlock1_p & v9703fc | !hlock1_p & v84563c;
assign a5f589 = hgrant2_p & a5f585 | !hgrant2_p & a5f588;
assign a5f7ce = hbusreq2 & a5f7c4 | !hbusreq2 & a5f7cd;
assign a5f422 = hbusreq2_p & a5f421 | !hbusreq2_p & a5f420;
assign c3b690 = hmaster1_p & c3b68f | !hmaster1_p & c3bccf;
assign a5f289 = hmaster0_p & a5f286 | !hmaster0_p & a5f288;
assign a5fb54 = hbusreq0 & a5fa8b | !hbusreq0 & a5fb4d;
assign a5fb88 = stateA1_p & v84563c | !stateA1_p & a5fb87;
assign a5f7f6 = stateG10_1_p & v970408 | !stateG10_1_p & a5f7f5;
assign c3b6e4 = hlock2_p & c3b6e2 | !hlock2_p & !c3b6e3;
assign b298b1 = hbusreq2_p & b298b0 | !hbusreq2_p & v84563c;
assign c3bcc2 = hmaster0_p & c3bcc1 | !hmaster0_p & c3bc71;
assign a5f11b = hmastlock_p & a5f11a | !hmastlock_p & v84563c;
assign c3bce3 = hbusreq2_p & c3bce2 | !hbusreq2_p & v84563c;
assign dead73 = hlock0_p & dead71 | !hlock0_p & !dead72;
assign a5fb74 = hlock0_p & v84563c | !hlock0_p & a5fb73;
assign adaedf = hlock1_p & adaebc | !hlock1_p & v84563c;
assign ab0cc0 = hlock2_p & ab0cbf | !hlock2_p & ab0c33;
assign ab0cf4 = hmaster0_p & ab0cf1 | !hmaster0_p & ab0cf3;
assign a5fd1a = decide_p & a5fb67 | !decide_p & a5fd19;
assign b26763 = hmaster1_p & b26762 | !hmaster1_p & !b266b3;
assign b29d72 = hbusreq2_p & b29d71 | !hbusreq2_p & v84563c;
assign a5f2da = hbusreq2_p & a5f2d9 | !hbusreq2_p & !v84563c;
assign ab0b04 = hbusreq3 & ab0af7 | !hbusreq3 & ab0b03;
assign ab06df = hbusreq2_p & ab06de | !hbusreq2_p & b29a4d;
assign b29a65 = hready & c3bd3b | !hready & b29a64;
assign c3bd8a = hlock1_p & v84563c | !hlock1_p & !dead6e;
assign a5f591 = hbusreq2_p & a5f590 | !hbusreq2_p & a5f58f;
assign ab06c6 = hbusreq3 & b29a7b | !hbusreq3 & ab06b5;
assign a5fbdd = hlock1_p & v84563c | !hlock1_p & a5fbdc;
assign a60186 = start_p & v8e1935 | !start_p & !a60185;
assign a5f22d = hready & a5f8b4 | !hready & a5f786;
assign c3bc60 = hbusreq1_p & dead6e | !hbusreq1_p & !v84563c;
assign a81cae = decide_p & a81cad | !decide_p & a81cac;
assign a5f1d1 = hlock1_p & a5f9dd | !hlock1_p & a5f1d0;
assign a5f0d5 = hlock0_p & a5f78d | !hlock0_p & a5f0d0;
assign c3bdb0 = locked_p & c3bdaf | !locked_p & !c3bcdb;
assign b26709 = hready_p & b266c4 | !hready_p & b26708;
assign b266e0 = hlock1_p & b266ca | !hlock1_p & b266df;
assign a5fab0 = hready & a5faac | !hready & a5faaf;
assign c3bdc6 = hlock2_p & c3bdc5 | !hlock2_p & v845660;
assign af3567 = hmaster1_p & af3565 | !hmaster1_p & af3566;
assign a81cc0 = hlock2_p & a81cb1 | !hlock2_p & v84563c;
assign c3bda3 = hmaster1_p & c3bc71 | !hmaster1_p & c3bda2;
assign c3bc9e = hmaster0_p & c3bc84 | !hmaster0_p & c3bc9d;
assign a5fc5e = hready & a5fc51 | !hready & v9703fc;
assign a5f3f7 = hlock1_p & a60172 | !hlock1_p & a5f3f6;
assign b29a7e = hbusreq2_p & b29a7d | !hbusreq2_p & c3bc21;
assign a5efd4 = hbusreq2_p & a5efd3 | !hbusreq2_p & a5ef6e;
assign b29b29 = decide_p & b29b28 | !decide_p & b29e57;
assign ab0bd8 = hbusreq0_p & b29e67 | !hbusreq0_p & deacbe;
assign a5fbda = hbusreq1 & a5fbd9 | !hbusreq1 & !a5fbab;
assign c3b6e7 = hmaster0_p & c3b6da | !hmaster0_p & c3b6e6;
assign a5f9df = hgrant1_p & a5f9de | !hgrant1_p & a5f9dd;
assign v970435 = hgrant2_p & v84563c | !hgrant2_p & v970434;
assign cea1a9 = hbusreq3_p & cea184 | !hbusreq3_p & cea1a8;
assign a5f36c = locked_p & a5f369 | !locked_p & a5f36b;
assign a5f8ed = hready & a60192 | !hready & !a60176;
assign a5f991 = hbusreq2 & a5f98e | !hbusreq2 & !a5f990;
assign a5ef7f = hbusreq2_p & a5edcb | !hbusreq2_p & a5ef7e;
assign a5f0a0 = hmaster1_p & a5f09f | !hmaster1_p & v84563c;
assign ce9e5e = jx1_p & ce9e29 | !jx1_p & ce9cde;
assign af34fc = hgrant3_p & af349b | !hgrant3_p & af34fb;
assign a5efb6 = hlock0_p & a5ee13 | !hlock0_p & a5ef3a;
assign b29a5b = hlock0_p & b29a5a | !hlock0_p & !v84563c;
assign a81d0c = hgrant3_p & a81d09 | !hgrant3_p & a81d0b;
assign cea16f = hbusreq2_p & cea16b | !hbusreq2_p & cea16e;
assign af35b4 = hlock2_p & af3563 | !hlock2_p & af352c;
assign a5f06f = locked_p & a5f6f2 | !locked_p & v845641;
assign b29ecd = hlock0_p & b29ecc | !hlock0_p & c3bd8e;
assign deaea2 = hlock0_p & deaea1 | !hlock0_p & !v84563c;
assign ab073b = hmaster1_p & ab06b5 | !hmaster1_p & ab073a;
assign c3b8cc = jx2_p & c3b621 | !jx2_p & c3b8cb;
assign a5f17c = hbusreq0_p & a5fb13 | !hbusreq0_p & ab0c31;
assign af3599 = hmaster0_p & af3597 | !hmaster0_p & af3598;
assign a5f9c4 = hlock2_p & a5f9c3 | !hlock2_p & v84563c;
assign a5eba2 = hgrant0_p & v84563c | !hgrant0_p & a5eba1;
assign c98ba3 = hready_p & c98ba1 | !hready_p & c98ba2;
assign a5f256 = hmaster0_p & a5f255 | !hmaster0_p & a5f8f7;
assign ab06ac = hready & ab06ab | !hready & v84563c;
assign c3b66b = hready & c3b66a | !hready & deadb2;
assign b29ae3 = hlock0_p & b29ae2 | !hlock0_p & !v84563c;
assign a5fb89 = start_p & v84563c | !start_p & a5fb88;
assign a5f520 = hbusreq1 & a5f3ef | !hbusreq1 & v84563c;
assign b29833 = locked_p & b29831 | !locked_p & !b29832;
assign b29907 = hlock0_p & cea37b | !hlock0_p & !v84563c;
assign c3b7ae = hbusreq3 & c3b7ad | !hbusreq3 & !v845644;
assign b26711 = hbusreq2_p & b26710 | !hbusreq2_p & b2670e;
assign c3b845 = hlock2_p & c3b7e8 | !hlock2_p & !c3b844;
assign c3b701 = hbusreq2_p & c3b700 | !hbusreq2_p & !c3b625;
assign b29a87 = hlock2_p & b29a86 | !hlock2_p & b29a7c;
assign c3b772 = hbusreq3_p & c3b72d | !hbusreq3_p & !c3b771;
assign cea18b = decide_p & cea18a | !decide_p & v84563c;
assign af3571 = locked_p & v84563c | !locked_p & af352c;
assign c3bdaa = hlock2_p & c3bda9 | !hlock2_p & dead2e;
assign c3b6b6 = hmaster1_p & c3b6ad | !hmaster1_p & c3b6b5;
assign dead82 = hbusreq2_p & dead81 | !hbusreq2_p & v84563c;
assign ab0c6c = hbusreq2_p & ab0c6b | !hbusreq2_p & v84563c;
assign b29a1d = decide_p & b29a1c | !decide_p & b29e57;
assign a5efe9 = hbusreq2_p & a5f583 | !hbusreq2_p & a5efe8;
assign a5efaf = hbusreq0_p & a5ee65 | !hbusreq0_p & a5efae;
assign a5fa70 = hbusreq3 & a5fa6a | !hbusreq3 & a5fa6f;
assign a5edf2 = locked_p & a5edf1 | !locked_p & v84563c;
assign cea2e4 = hburst0 & cea2e2 | !hburst0 & cea2e3;
assign ab0adc = hready & c98b96 | !hready & v84563c;
assign b26714 = hbusreq2_p & b2670c | !hbusreq2_p & b26713;
assign c3b699 = hlock2_p & c3b696 | !hlock2_p & !c3b698;
assign b29a8f = hbusreq2_p & b29a8e | !hbusreq2_p & !c3bc21;
assign b29a6d = hgrant2_p & b29a69 | !hgrant2_p & b29a6c;
assign cea26b = hmastlock_p & cea26a | !hmastlock_p & v84563c;
assign deae7f = hbusreq1_p & deadba | !hbusreq1_p & !v84563c;
assign d40d96 = hbusreq2_p & d40d94 | !hbusreq2_p & d40d51;
assign c3bcd1 = hgrant2_p & c3bc06 | !hgrant2_p & c3bc0e;
assign cea3d8 = hbusreq1_p & deadba | !hbusreq1_p & !cea26a;
assign v868347 = jx1_p & v84563c | !jx1_p & !v84563c;
assign a5fb8e = hlock1_p & a5fb8b | !hlock1_p & !a5fb8d;
assign v9703fc = hmastlock_p & v9703fb | !hmastlock_p & v84563c;
assign ab05f5 = hlock2 & ab05ee | !hlock2 & ab05f1;
assign a5f383 = hbusreq3 & a5f373 | !hbusreq3 & !a5f382;
assign a5f945 = hlock2 & a5f93f | !hlock2 & a5f944;
assign cea253 = hgrant1_p & cea251 | !hgrant1_p & cea252;
assign a5eea1 = hlock1_p & a5fc09 | !hlock1_p & !a5ee52;
assign c3b636 = locked_p & v84563c | !locked_p & c3b635;
assign af35bd = hmaster0_p & af35bc | !hmaster0_p & af359d;
assign c3b72a = hlock3_p & c3b729 | !hlock3_p & !c3b6d2;
assign ab0b24 = hlock2_p & ab0b21 | !hlock2_p & ab0b23;
assign ab0511 = hlock0_p & v84563c | !hlock0_p & b298a0;
assign a5f749 = hmaster0_p & a5f73f | !hmaster0_p & a5f748;
assign a5f742 = hlock0_p & a5f6e9 | !hlock0_p & a5f741;
assign a9b9ef = hgrant3_p & a9b9ee | !hgrant3_p & !a9b9eb;
assign ab0ba4 = locked_p & v84563c | !locked_p & b29d8a;
assign a5fa11 = hlock1_p & a6016f | !hlock1_p & !a5fa10;
assign a5f3b2 = hlock2_p & a5f3af | !hlock2_p & a5f3b1;
assign ab0b5c = hlock0_p & v845660 | !hlock0_p & !b29d87;
assign cea2f4 = hbusreq2_p & cea2f3 | !hbusreq2_p & cea15a;
assign ab0c0a = hlock2 & ab0c06 | !hlock2 & ab0c09;
assign a5f15f = hbusreq0 & a5f14e | !hbusreq0 & a5f15e;
assign cea1b4 = hready & cea1b3 | !hready & cea151;
assign deae96 = hlock2_p & deae95 | !hlock2_p & !v84563c;
assign a5f6e7 = hready & a5f6e4 | !hready & a5f6e6;
assign a5edf9 = hbusreq2 & a5edf5 | !hbusreq2 & a5edf8;
assign dead3b = hbusreq2_p & dead3a | !hbusreq2_p & dead39;
assign af34a6 = hlock0_p & af3c4f | !hlock0_p & af3c6b;
assign a5f24c = hready & a5f828 | !hready & a5fa1d;
assign b29e97 = hgrant0_p & c3bceb | !hgrant0_p & !b29e96;
assign cea1a0 = hgrant2_p & cea19c | !hgrant2_p & cea19f;
assign c3b62b = locked_p & dead7b | !locked_p & !v845648;
assign a81d03 = hmaster1_p & a81cdc | !hmaster1_p & v84563c;
assign a5fcb4 = hbusreq2_p & a5fcb0 | !hbusreq2_p & !a5fcb3;
assign b29aab = hgrant2_p & b29aa6 | !hgrant2_p & !b29aaa;
assign b2a00f = hlock0_p & b2a00e | !hlock0_p & !c3bd60;
assign a5f529 = hbusreq1 & a5f528 | !hbusreq1 & !v84563c;
assign a5f3c5 = hready & a5f3c4 | !hready & v84563c;
assign a5f78d = hready & a5f9f6 | !hready & deac52;
assign ab0b49 = hbusreq3 & c3bc3c | !hbusreq3 & !ab0b48;
assign c3b68b = hbusreq3 & c3b66f | !hbusreq3 & c3b68a;
assign a5fa6d = hlock0_p & a5fa6c | !hlock0_p & v84563c;
assign af34ec = hgrant0_p & af34e5 | !hgrant0_p & af34eb;
assign adaf0e = hgrant0_p & adaf04 | !hgrant0_p & adaf0d;
assign c3b70c = hgrant2_p & c3b70b | !hgrant2_p & v845660;
assign ab0ce2 = hmaster1_p & ab0bd7 | !hmaster1_p & ab0ce1;
assign b29a6a = hbusreq2_p & b29a5c | !hbusreq2_p & v84563c;
assign c3b64a = hlock0_p & c3b648 | !hlock0_p & c3b649;
assign ab0610 = hready & deae67 | !hready & v845646;
assign a5f6fb = hbusreq2 & a5f6f9 | !hbusreq2 & a5f6fa;
assign c3bc67 = hlock2_p & c3bc64 | !hlock2_p & !c3bc66;
assign cea389 = locked_p & v84563c | !locked_p & !cea378;
assign a5ea79 = hgrant2_p & a5ea74 | !hgrant2_p & a5ea78;
assign a5ef18 = hmaster0_p & a5ef05 | !hmaster0_p & a5ef17;
assign v84564a = hbusreq2_p & v84563c | !hbusreq2_p & !v84563c;
assign b29f0e = hgrant1_p & b29f0c | !hgrant1_p & b29f0d;
assign c3bc43 = hmaster0_p & cea0e8 | !hmaster0_p & c3bc42;
assign dea79f = hbusreq2_p & deae33 | !hbusreq2_p & deae32;
assign cea269 = hburst1 & v84563c | !hburst1 & deac4e;
assign ab057d = hready & c3b6c5 | !hready & deada8;
assign deaea9 = hmaster1_p & deaea6 | !hmaster1_p & deaea8;
assign ab0bb5 = hmaster0_p & ab0b87 | !hmaster0_p & ab0bb4;
assign a5fb69 = hready_p & a60147 | !hready_p & a5fb68;
assign c3b651 = hlock0_p & deae59 | !hlock0_p & v845648;
assign af34f1 = hmaster1_p & d40d60 | !hmaster1_p & af3497;
assign c3b6f5 = hmaster1_p & c3b6d7 | !hmaster1_p & dead2e;
assign a5f71d = hready & a5fb73 | !hready & b266a2;
assign af34bb = locked_p & af34b5 | !locked_p & af34ba;
assign a5ef9e = hlock0_p & a5ee12 | !hlock0_p & a5ef9d;
assign ab0687 = hmaster0_p & ab0682 | !hmaster0_p & ab0686;
assign a5f029 = hmaster1_p & a5f92d | !hmaster1_p & a5f028;
assign a5fc24 = hbusreq2_p & v84563c | !hbusreq2_p & a5fc23;
assign v97040b = hlock1_p & v9703fc | !hlock1_p & v97040a;
assign ab064a = decide_p & ab0649 | !decide_p & v84563c;
assign af3596 = hlock3_p & af3595 | !hlock3_p & af356d;
assign af3c13 = hlock2_p & af3c12 | !hlock2_p & v845646;
assign a5f57e = hlock1_p & a5f8d2 | !hlock1_p & a5f57d;
assign c3b798 = hlock0_p & c3bcdc | !hlock0_p & dead77;
assign adaee0 = locked_p & adaedf | !locked_p & v84563c;
assign dead4e = hlock3_p & dead2b | !hlock3_p & dead4d;
assign d40d66 = start_p & v84563c | !start_p & !c06d34;
assign a5f239 = hlock0_p & a5f8ca | !hlock0_p & a5f233;
assign b2995f = hbusreq2_p & b2995b | !hbusreq2_p & v84563c;
assign bdb59f = hmaster1_p & v845660 | !hmaster1_p & c3bca4;
assign a5fa8c = hlock2_p & a5fa89 | !hlock2_p & a5fa8b;
assign b29f63 = hbusreq2_p & b29f62 | !hbusreq2_p & !v84563c;
assign cea391 = locked_p & v84563c | !locked_p & !cea380;
assign af35ac = hmaster1_p & af352c | !hmaster1_p & af3581;
assign a5f1f2 = hbusreq1 & v84563c | !hbusreq1 & !a5f1f1;
assign a5f204 = hmaster1_p & v84563c | !hmaster1_p & a5f203;
assign c3b8ae = hbusreq2_p & c3b8ab | !hbusreq2_p & c3b7ea;
assign b29d5a = hbusreq2_p & b29d59 | !hbusreq2_p & v84563c;
assign a5fae9 = hgrant2_p & a5fae3 | !hgrant2_p & a5fae8;
assign a5ee25 = hbusreq1 & a5fb71 | !hbusreq1 & v84563c;
assign b29a94 = hgrant2_p & b29a90 | !hgrant2_p & b29a93;
assign ab056f = hready & b2994d | !hready & c3bd5d;
assign d40d8d = hgrant3_p & d40d64 | !hgrant3_p & d40d8c;
assign b29aa8 = hlock0_p & b29aa7 | !hlock0_p & !v84563c;
assign d40d5c = hlock3_p & d40d56 | !hlock3_p & d40d5b;
assign a5f385 = locked_p & v84563c | !locked_p & a5f36b;
assign a5eec5 = hbusreq0_p & a5f3cf | !hbusreq0_p & a5eec4;
assign c3b820 = hlock2_p & c3b81f | !hlock2_p & !c3b80a;
assign cea2f6 = hmaster1_p & cea2f0 | !hmaster1_p & cea2f5;
assign cea2b7 = hready_p & cea23c | !hready_p & cea2b6;
assign ab0bed = hgrant2_p & ab0beb | !hgrant2_p & ab0bec;
assign c3b663 = hgrant1_p & c3b662 | !hgrant1_p & deae74;
assign d40d9c = hgrant3_p & d40d93 | !hgrant3_p & d40d9b;
assign b29ea9 = locked_p & b29ea8 | !locked_p & !v84563c;
assign a5f757 = decide_p & a5f74a | !decide_p & a5f756;
assign cea414 = hlock0_p & cea3cd | !hlock0_p & cea412;
assign c3bc86 = hlock0_p & c3bc85 | !hlock0_p & !c3bc65;
assign b8ace9 = locked_p & v8c6711 | !locked_p & b8ace3;
assign a5f750 = hbusreq2 & a5fc6d | !hbusreq2 & v84563c;
assign b266bd = hmaster1_p & b266ba | !hmaster1_p & b266bc;
assign b29f39 = hgrant2_p & b29f36 | !hgrant2_p & b29f38;
assign cea2b0 = hlock2_p & cea2af | !hlock2_p & cea887;
assign deac87 = hlock0_p & deac6c | !hlock0_p & deac86;
assign ab0c47 = hbusreq2_p & ab0c46 | !hbusreq2_p & ab0ade;
assign a5f3dc = hmaster1_p & a5f3d9 | !hmaster1_p & a5f3db;
assign af35a2 = hgrant3_p & af3578 | !hgrant3_p & af35a1;
assign a5f1b2 = hready & a5f1ac | !hready & !a5f1b1;
assign a5fc9d = hbusreq1_p & a5fc78 | !hbusreq1_p & !a5fc7d;
assign dead33 = hmastlock_p & dead32 | !hmastlock_p & !v84563c;
assign ce9d33 = hgrant2_p & cea2a8 | !hgrant2_p & ce9d32;
assign dea782 = hbusreq2_p & deae1f | !hbusreq2_p & !deada8;
assign ab0678 = hmaster1_p & ab0673 | !hmaster1_p & ab0677;
assign a5f363 = jx0_p & a5f6e3 | !jx0_p & a5f362;
assign c3bca3 = hmaster0_p & dead2e | !hmaster0_p & c3bca2;
assign af3518 = hlock0_p & v84563c | !hlock0_p & v845642;
assign a5f887 = hgrant2_p & a5f885 | !hgrant2_p & a5f886;
assign a5f721 = hlock2_p & a5f720 | !hlock2_p & v84563c;
assign deae70 = decide_p & deae6f | !decide_p & v84563c;
assign c3bcc0 = hgrant2_p & c3bc6d | !hgrant2_p & c3bc81;
assign cea40d = hlock2_p & cea40c | !hlock2_p & cea3fb;
assign ab0589 = hlock0_p & v845660 | !hlock0_p & cea37b;
assign ab06c0 = hlock2_p & ab06bf | !hlock2_p & b29a7b;
assign a5fd36 = hlock2_p & a5fd35 | !hlock2_p & a5fad6;
assign adaebf = hmaster0_p & adaebe | !hmaster0_p & v84563c;
assign a5e9cf = hmaster1_p & a5e9cd | !hmaster1_p & a5e9ce;
assign cea427 = hgrant2_p & cea423 | !hgrant2_p & cea426;
assign a5eb40 = hbusreq2 & a5eb3e | !hbusreq2 & a5eb3f;
assign cea32f = decide_p & cea32e | !decide_p & a57859;
assign c3bd3f = hlock0_p & c3bd2d | !hlock0_p & !c3bd3e;
assign cea879 = hgrant2_p & cea86f | !hgrant2_p & cea878;
assign a6018c = hready & a60189 | !hready & a6018b;
assign b29d36 = hlock2 & deacbe | !hlock2 & b29d34;
assign c3b6ff = hmaster0_p & c3b6f5 | !hmaster0_p & c3b6fe;
assign b29990 = locked_p & c3bbba | !locked_p & !cea38d;
assign cea0d5 = hgrant2_p & cea0d2 | !hgrant2_p & cea0d4;
assign a5ef3a = hbusreq0_p & a5ee13 | !hbusreq0_p & a5f390;
assign ab0bb7 = hbusreq3 & c3bca0 | !hbusreq3 & !v845660;
assign cea35c = hlock2_p & cea35b | !hlock2_p & v845660;
assign ab052c = hlock2_p & b29832 | !hlock2_p & ab052b;
assign a5ef0c = hbusreq0_p & a5edec | !hbusreq0_p & !a5ef0b;
assign a9b9da = hgrant2_p & v84563c | !hgrant2_p & !a9b9d9;
assign cea179 = hlock1_p & dead76 | !hlock1_p & v84563c;
assign a5f03a = hmaster1_p & a5fd28 | !hmaster1_p & a5f039;
assign a5fc52 = hlock1_p & a5fc51 | !hlock1_p & v84563c;
assign c3bd11 = hmastlock_p & c3bd10 | !hmastlock_p & v84566c;
assign ab0740 = hlock2_p & ab067a | !hlock2_p & !b29b1c;
assign a5f3a1 = locked_p & a5f3a0 | !locked_p & a5f36b;
assign b29f9b = hlock0_p & b29f99 | !hlock0_p & b29f9a;
assign a5fcd1 = hready & a5fb8b | !hready & v84563c;
assign c3bdbd = hlock1_p & deae02 | !hlock1_p & !v84563c;
assign ab067e = hmaster0_p & ab0678 | !hmaster0_p & ab067d;
assign a5f0d0 = hbusreq0_p & a5f7be | !hbusreq0_p & a5f7ba;
assign c3b7e1 = hmaster1_p & c3b7d7 | !hmaster1_p & c3b7e0;
assign b299ef = hmaster0_p & b299ec | !hmaster0_p & !b299ee;
assign ab06a8 = hmaster1_p & ab06a0 | !hmaster1_p & ab06a7;
assign a5efa3 = hbusreq0 & a5ef9f | !hbusreq0 & !a5efa2;
assign cea342 = hlock0_p & cea341 | !hlock0_p & v84563c;
assign a5f596 = hbusreq2_p & a5f590 | !hbusreq2_p & a5f58d;
assign ab06e1 = hlock0_p & b29f9a | !hlock0_p & !dead41;
assign af3492 = hbusreq2_p & af348b | !hbusreq2_p & d40d33;
assign cea45d = hmaster0_p & cea455 | !hmaster0_p & cea45c;
assign c3b73c = hmaster1_p & c3b737 | !hmaster1_p & c3b73b;
assign a5f09d = hbusreq2_p & a5f09b | !hbusreq2_p & a5f09c;
assign c3b710 = hlock3_p & c3b6f4 | !hlock3_p & c3b70f;
assign a5eb87 = hmaster1_p & a5eb86 | !hmaster1_p & !a5ea25;
assign a5ea2a = hbusreq0_p & a5fcce | !hbusreq0_p & v84563c;
assign d40d7f = hmaster0_p & d40d60 | !hmaster0_p & d40d7e;
assign a5fc59 = hmaster1_p & v84563c | !hmaster1_p & a5fc58;
assign b29f8b = hbusreq2_p & b29f8a | !hbusreq2_p & v84563c;
assign af34ee = hmaster1_p & af3c49 | !hmaster1_p & af3487;
assign b29cfb = hbusreq2_p & b29cf8 | !hbusreq2_p & v84563c;
assign a5f3d5 = hbusreq1_p & a5fc69 | !hbusreq1_p & !v84563c;
assign cea8a7 = hmastlock_p & deacb3 | !hmastlock_p & v84566c;
assign deac63 = hgrant2_p & deac60 | !hgrant2_p & deac62;
assign ab05fd = hbusreq2_p & ab057f | !hbusreq2_p & ab05fc;
assign a5fc60 = hlock2_p & a5fc5f | !hlock2_p & v84563c;
assign c3b878 = decide_p & c3b877 | !decide_p & !v845660;
assign cea354 = hmaster1_p & cea2a7 | !hmaster1_p & cea2b1;
assign v97043a = hmaster1_p & v970439 | !hmaster1_p & v84563c;
assign af3c1a = hbusreq2_p & af3c19 | !hbusreq2_p & v845646;
assign b2997c = hready & deae5a | !hready & !v84563c;
assign a5eb3d = hbusreq2 & a5ea1f | !hbusreq2 & !a5ea21;
assign ab0722 = hmaster0_p & ab071e | !hmaster0_p & ab06c4;
assign b29837 = hbusreq3 & b29829 | !hbusreq3 & b29836;
assign a5f4a2 = hbusreq1_p & a60167 | !hbusreq1_p & v84563c;
assign ab06cc = hlock0_p & ab06ca | !hlock0_p & !ab06b1;
assign b29f32 = hlock0_p & b29f1f | !hlock0_p & b29f31;
assign deadce = hbusreq1_p & v84563c | !hbusreq1_p & !deac52;
assign af34e6 = locked_p & af3c49 | !locked_p & af34ba;
assign cea170 = hbusreq3 & cea16f | !hbusreq3 & cea15c;
assign v97042a = hmaster1_p & v970421 | !hmaster1_p & v970429;
assign a5f022 = hmaster1_p & a5f6db | !hmaster1_p & a5f021;
assign v97042d = hmaster0_p & v97042c | !hmaster0_p & v97042a;
assign a5f35f = decide_p & a5f335 | !decide_p & a5f35e;
assign b2675c = hbusreq1_p & b26693 | !hbusreq1_p & !b26756;
assign dead8e = hbusreq2_p & dead8d | !hbusreq2_p & v84563c;
assign af3c52 = hlock2_p & af3c51 | !hlock2_p & af3c50;
assign v845670 = stateG3_0_p & v84563c | !stateG3_0_p & !v84563c;
assign a5f74c = hbusreq2_p & a5f74b | !hbusreq2_p & v84563c;
assign cea14e = hbusreq2_p & cea149 | !hbusreq2_p & cea14d;
assign ab0bbc = hbusreq3 & v84563c | !hbusreq3 & ab0bba;
assign a5f2d7 = hbusreq2 & a5fcd9 | !hbusreq2 & !v84563c;
assign b29ee9 = hmastlock_p & deac50 | !hmastlock_p & v84566c;
assign adaf09 = hmaster1_p & v84563c | !hmaster1_p & adaf08;
assign dead7e = locked_p & dead7d | !locked_p & !v84563c;
assign af35c5 = jx2_p & af3c10 | !jx2_p & !af35c4;
assign cea338 = hbusreq3 & cea298 | !hbusreq3 & cea337;
assign ce9db6 = hbusreq3 & ce9db5 | !hbusreq3 & v84563c;
assign cea8ab = hlock1_p & v84563c | !hlock1_p & !cea8aa;
assign a5fc67 = hlock3_p & a5fc42 | !hlock3_p & a5fc66;
assign ab059d = hlock2_p & ab059a | !hlock2_p & ab059c;
assign b2676d = hmaster0_p & b2676c | !hmaster0_p & b266c2;
assign ab0717 = hlock2_p & ab0715 | !hlock2_p & ab0716;
assign c3bd9b = locked_p & c3bc7a | !locked_p & c3bd9a;
assign dea766 = hlock1_p & deacdf | !hlock1_p & v84563c;
assign a5eb47 = decide_p & a5eb1c | !decide_p & a5eb46;
assign cea884 = hready & deac57 | !hready & cea883;
assign a5f8f3 = hbusreq2_p & a5f8cc | !hbusreq2_p & a5fad1;
assign a5f1b1 = hbusreq1 & dead40 | !hbusreq1 & a5f1b0;
assign a5ee85 = hbusreq2_p & a5ee80 | !hbusreq2_p & a5ee84;
assign a5f297 = hmaster0_p & a5f296 | !hmaster0_p & a5f748;
assign b29d52 = locked_p & v84563c | !locked_p & !b29d51;
assign a5f0da = hbusreq2 & a5f0d5 | !hbusreq2 & a5f0d9;
assign b29d6a = hbusreq2_p & b29d69 | !hbusreq2_p & b29d68;
assign deae3a = hbusreq2_p & dead9a | !hbusreq2_p & v845644;
assign cea491 = hbusreq3 & cea44a | !hbusreq3 & cea3a1;
assign cea187 = hmaster1_p & v84563c | !hmaster1_p & !deacaa;
assign af35a9 = hready_p & af35a5 | !hready_p & af35a8;
assign a5eb94 = hbusreq2 & a5ea60 | !hbusreq2 & a5eb93;
assign a5f7f4 = start_p & v8e1935 | !start_p & a5f7f3;
assign b29a8a = hmaster1_p & b29a89 | !hmaster1_p & !b299ed;
assign b29d4c = hmaster1_p & b29d3e | !hmaster1_p & b29d4b;
assign af357a = hbusreq0_p & v84563c | !hbusreq0_p & af3579;
assign cea479 = hgrant1_p & cea478 | !hgrant1_p & cea255;
assign a5fbf3 = hbusreq2 & a5fbe9 | !hbusreq2 & a5fbf2;
assign cea3e8 = hlock1_p & v84565a | !hlock1_p & !deae7f;
assign adaed5 = hmaster0_p & adaed4 | !hmaster0_p & adaed2;
assign a5ea63 = hbusreq2_p & a5ea5f | !hbusreq2_p & a5ea62;
assign b29ff5 = hmaster1_p & b29ff4 | !hmaster1_p & b29f6c;
assign adaf00 = locked_p & adaeff | !locked_p & v84563c;
assign cea396 = hlock2_p & cea394 | !hlock2_p & cea395;
assign cea33d = hlock3_p & cea33c | !hlock3_p & cea2b4;
assign deae9a = hbusreq2_p & deae96 | !hbusreq2_p & deae95;
assign ab0633 = hbusreq2_p & ab0560 | !hbusreq2_p & ab0632;
assign b29a7a = hlock2 & b29ce0 | !hlock2 & b29a79;
assign c3b810 = hlock0_p & c3b80f | !hlock0_p & !dead77;
assign ab0b7b = hlock2 & ab0b78 | !hlock2 & ab0b7a;
assign a5ebca = hmaster1_p & a5ebc9 | !hmaster1_p & a5f163;
assign b26789 = hmaster1_p & b26788 | !hmaster1_p & !b266e5;
assign deada0 = decide_p & dead9f | !decide_p & v84563c;
assign a5f013 = hgrant3_p & a5ef95 | !hgrant3_p & a5f012;
assign a5fbe8 = hready & a5fbe3 | !hready & a5fbe7;
assign a5e9d5 = hlock2_p & a5e9d4 | !hlock2_p & a5f199;
assign a5eaa2 = hmaster0_p & a5ea99 | !hmaster0_p & a5eaa1;
assign a9b9d7 = hmaster1_p & v84563c | !hmaster1_p & !a9b9d6;
assign a5f9de = stateG10_1_p & v84563c | !stateG10_1_p & a5f9dd;
assign b29e99 = hbusreq2_p & v84564c | !hbusreq2_p & !v845644;
assign a5ef06 = hbusreq1_p & a5fcd5 | !hbusreq1_p & !v84563c;
assign a5fca5 = hlock1_p & a5fc87 | !hlock1_p & a5fca4;
assign a5ea86 = hbusreq2_p & a5ea85 | !hbusreq2_p & a5ea62;
assign c3b6af = hbusreq0_p & c3b698 | !hbusreq0_p & c3b6a1;
assign deade5 = hmaster1_p & deaddc | !hmaster1_p & deade4;
assign a5f21a = hgrant0_p & a5f211 | !hgrant0_p & a5f219;
assign cea472 = hgrant2_p & cea471 | !hgrant2_p & !v845660;
assign a5fc29 = hlock0_p & v84563c | !hlock0_p & a5fc28;
assign cea2e2 = start_p & v84563c | !start_p & cea1ad;
assign a81cac = hmaster0_p & a81cab | !hmaster0_p & v84563c;
assign ce9cda = decide_p & ce9cd9 | !decide_p & a57859;
assign b29a20 = hgrant3_p & b299f5 | !hgrant3_p & b29a1f;
assign af3c59 = hlock0_p & af3c57 | !hlock0_p & af3c58;
assign cea48b = hmaster1_p & cea48a | !hmaster1_p & !cea1a1;
assign a5ec23 = hready_p & a5f035 | !hready_p & a5ec21;
assign deae8c = hbusreq3 & deae8a | !hbusreq3 & deae8b;
assign af3c31 = hgrant2_p & af3c2b | !hgrant2_p & af3c30;
assign c3b677 = hmastlock_p & cea26a | !hmastlock_p & c3b676;
assign a5e9c3 = hlock1_p & a60177 | !hlock1_p & !a5e9c2;
assign b29f7e = hbusreq2_p & b29f7d | !hbusreq2_p & v84565a;
assign a5fbcc = hbusreq2 & a5fbcb | !hbusreq2 & a5fbc6;
assign b2990f = hlock3_p & b298a9 | !hlock3_p & b2990e;
assign deadea = hgrant2_p & deacbf | !hgrant2_p & deacc2;
assign ce9e0a = hmaster0_p & ce9e09 | !hmaster0_p & ce9d4f;
assign a5ee0c = hlock0_p & a60141 | !hlock0_p & a5f38f;
assign a5ef53 = hlock0_p & a5ef52 | !hlock0_p & a5f4fc;
assign c3bcf9 = hlock2_p & c3bcf8 | !hlock2_p & v84563c;
assign af34fa = decide_p & af34f0 | !decide_p & af34f9;
assign a5f4cb = hbusreq1 & a5f4ca | !hbusreq1 & !v84563c;
assign a5ee6c = hlock0_p & a60140 | !hlock0_p & a5f3b8;
assign dead56 = hmaster0_p & dead55 | !hmaster0_p & dead54;
assign deae0c = locked_p & v84563c | !locked_p & !deae0b;
assign dea76b = hmaster1_p & dea76a | !hmaster1_p & dead3c;
assign af3c4a = stateA1_p & v84563c | !stateA1_p & v845674;
assign a5f883 = hbusreq2 & a5f882 | !hbusreq2 & v84563c;
assign a5ee66 = locked_p & v84563c | !locked_p & a5ee65;
assign a5f783 = hlock1_p & a60167 | !hlock1_p & a5f9f5;
assign a81cdc = locked_p & a81cdb | !locked_p & v84563c;
assign c3bc4a = hlock2_p & c3bc49 | !hlock2_p & dead2e;
assign a5fc8a = stateA1_p & v845652 | !stateA1_p & a81ca6;
assign a5f0a2 = hlock3_p & a5f090 | !hlock3_p & a5f0a1;
assign b29f3d = hready & deac5b | !hready & v84563c;
assign c3bc52 = locked_p & v84563c | !locked_p & c3bc51;
assign c3bce5 = hready & deace1 | !hready & v84563c;
assign c3bbf8 = hgrant1_p & c3bbf6 | !hgrant1_p & c3bbf7;
assign a9b9eb = hready_p & a9b9ea | !hready_p & !v84563c;
assign b29f79 = hready & b29f78 | !hready & v84563c;
assign ce9cc4 = hbusreq2_p & ce9cc3 | !hbusreq2_p & !cea405;
assign dead0a = hlock1_p & v84563c | !hlock1_p & !dead09;
assign deae2f = hgrant3_p & deadf7 | !hgrant3_p & !deae2e;
assign b29a50 = hbusreq3 & b29a4f | !hbusreq3 & v84563c;
assign a5fc41 = hmaster0_p & a5fbf8 | !hmaster0_p & a5fc40;
assign a5fcf2 = hbusreq1_p & a5fb8b | !hbusreq1_p & !a5fcd5;
assign a5e9c5 = hbusreq0_p & a5fb32 | !hbusreq0_p & ab0c31;
assign deae23 = hlock0_p & deae22 | !hlock0_p & !deadba;
assign c3bccf = hgrant2_p & c3bbef | !hgrant2_p & c3bbf2;
assign ab0574 = hbusreq2_p & ab0573 | !hbusreq2_p & !ab0572;
assign bdb5a7 = hgrant2_p & v84565a | !hgrant2_p & !bdb598;
assign c3b82a = hbusreq2_p & c3b7a5 | !hbusreq2_p & c3b829;
assign a5ef11 = hbusreq1 & a5ef10 | !hbusreq1 & !v84563c;
assign b29954 = hbusreq2_p & b29953 | !hbusreq2_p & !v84563c;
assign deac9f = hmaster0_p & deac64 | !hmaster0_p & !deac9e;
assign a5fbc7 = locked_p & v84563c | !locked_p & a5fbc6;
assign a5ea12 = hlock0_p & a5ea11 | !hlock0_p & a5e9b4;
assign b29cbd = hbusreq2_p & b29cbc | !hbusreq2_p & b29cbb;
assign b2993a = hready & b29939 | !hready & !v84563c;
assign a5f998 = hbusreq0 & a5f97b | !hbusreq0 & !a5f997;
assign ab06ab = hlock1_p & v84565a | !hlock1_p & ab06aa;
assign a5ef8e = hgrant2_p & a5ef88 | !hgrant2_p & a5ef8d;
assign a5ee8f = hlock2_p & a5ee8e | !hlock2_p & !a5ee31;
assign b29f52 = hlock0_p & b29f51 | !hlock0_p & c3bd61;
assign b26741 = hgrant0_p & b2671c | !hgrant0_p & b26740;
assign b29a9d = hlock3_p & b29a8b | !hlock3_p & b29a9c;
assign b266e6 = hmaster1_p & b266d6 | !hmaster1_p & b266e5;
assign deacaf = hbusreq2_p & deacac | !hbusreq2_p & deacab;
assign a5fc93 = hlock0_p & a5fc89 | !hlock0_p & a5fc92;
assign cea484 = hlock2_p & cea483 | !hlock2_p & cea3ea;
assign a9b9e0 = hmaster0_p & a9b9db | !hmaster0_p & !a9b9df;
assign ab0c19 = hmaster0_p & ab0c12 | !hmaster0_p & ab0c18;
assign cea3af = decide_p & cea3ae | !decide_p & v84563c;
assign a5f8d9 = hburst1_p & c07311 | !hburst1_p & c06d34;
assign af3c6d = hmaster0_p & af3c6c | !hmaster0_p & af3c4c;
assign a5ef27 = hmaster1_p & a5ef26 | !hmaster1_p & v84563c;
assign deadd8 = hbusreq3 & deadd2 | !hbusreq3 & deadd7;
assign deae6a = hbusreq3 & deae69 | !hbusreq3 & !v84563c;
assign deae4f = locked_p & deae4e | !locked_p & !v84563c;
assign a5f96d = hbusreq0_p & a5f726 | !hbusreq0_p & a5f96c;
assign b299cb = hmaster0_p & b299b0 | !hmaster0_p & b2990d;
assign c3b61d = decide_p & c3b61c | !decide_p & v845660;
assign c3b6de = hready & c3b622 | !hready & c3b6dd;
assign a5f986 = stateA1_p & a5fb9d | !stateA1_p & a5fc75;
assign ce9cd1 = hmaster0_p & ce9cd0 | !hmaster0_p & cea1a4;
assign a5f838 = hmastlock_p & v845654 | !hmastlock_p & !v84563c;
assign c3bd8f = hlock0_p & c3bd8c | !hlock0_p & !c3bd8e;
assign deae2a = hmaster1_p & deae29 | !hmaster1_p & !v84563c;
assign a5ee78 = hbusreq2 & a5ee75 | !hbusreq2 & a5ee77;
assign b266b8 = locked_p & b26694 | !locked_p & b26695;
assign a5f042 = hmaster0_p & a5f6da | !hmaster0_p & a5f041;
assign a5fc4b = hbusreq0 & a5fc45 | !hbusreq0 & a5fc4a;
assign cea36e = hmaster0_p & cea36d | !hmaster0_p & cea29b;
assign cea1c2 = hbusreq2_p & cea1c1 | !hbusreq2_p & v84563c;
assign adaef0 = hbusreq1_p & adaebc | !hbusreq1_p & adaeea;
assign b29d7e = locked_p & b29d7d | !locked_p & !v84563c;
assign ab06d5 = hgrant2_p & ab06cf | !hgrant2_p & ab06d4;
assign dea6f3 = hmaster1_p & v84563c | !hmaster1_p & !dead5f;
assign a5f94f = hmaster1_p & a5f92d | !hmaster1_p & a5f94e;
assign a5fc6a = hbusreq1_p & v84563c | !hbusreq1_p & !a5fc69;
assign ab05aa = hlock0_p & v84563c | !hlock0_p & !b29990;
assign ab0c28 = hbusreq2_p & ab0c27 | !hbusreq2_p & v84563c;
assign a5ea49 = hbusreq0 & a5ea48 | !hbusreq0 & a5f084;
assign a5f0a7 = hbusreq3 & a5f0a4 | !hbusreq3 & !a5f0a6;
assign adaf0c = hmaster1_p & adaf0b | !hmaster1_p & v84563c;
assign c3b6d7 = hlock0_p & c3b631 | !hlock0_p & !c3b625;
assign deacfc = hbusreq0_p & deace9 | !hbusreq0_p & deacfb;
assign af358a = hmaster0_p & af3536 | !hmaster0_p & af3589;
assign c98b96 = hlock1_p & v84563c | !hlock1_p & c98b95;
assign a5ea24 = hbusreq0_p & a5fcc8 | !hbusreq0_p & v84563c;
assign dea75c = decide_p & dea75b | !decide_p & v84563c;
assign deae92 = hlock2_p & deae91 | !hlock2_p & !v84563c;
assign a5f1e3 = hlock0_p & a5f1e2 | !hlock0_p & !a5fc2c;
assign b29e55 = hgrant0_p & b29e47 | !hgrant0_p & !b29e54;
assign a5f52b = hbusreq1 & a5f52a | !hbusreq1 & !v84563c;
assign c3b850 = hbusreq3 & c3b84e | !hbusreq3 & c3b84f;
assign a5fb03 = hmaster1_p & v84563c | !hmaster1_p & a5fb02;
assign a5f970 = locked_p & a5f96f | !locked_p & v845641;
assign a5fc1f = hbusreq2_p & a5fc19 | !hbusreq2_p & a5fc1e;
assign a5fb11 = hgrant1_p & a5fb10 | !hgrant1_p & a60167;
assign ab05db = hbusreq0_p & b29990 | !hbusreq0_p & cea44a;
assign dea6c8 = decide_p & dea6c7 | !decide_p & v84563c;
assign a5f08d = hbusreq0 & a5f08c | !hbusreq0 & a5fbc1;
assign ab0c30 = hlock2 & ab0ae6 | !hlock2 & ab0c2f;
assign a5f6d4 = hbusreq3 & a5f6d1 | !hbusreq3 & a5f6d3;
assign a5f539 = stateG10_1_p & v84563c | !stateG10_1_p & deadd3;
assign c3bd5c = hlock1_p & v84563c | !hlock1_p & !c3bd5b;
assign dead45 = hlock2_p & dead34 | !hlock2_p & v84563c;
assign a5e9e8 = hbusreq2_p & a5e9e0 | !hbusreq2_p & a5e9df;
assign b29ffe = hlock2_p & b29ffd | !hlock2_p & dead2e;
assign af34d2 = hlock2_p & af3c5e | !hlock2_p & af3c4c;
assign b29fed = hbusreq2_p & b29fec | !hbusreq2_p & v84563c;
assign ab0bbf = hmaster1_p & ab0bbb | !hmaster1_p & ab0bbe;
assign dead90 = hbusreq2_p & dead8f | !hbusreq2_p & v84563c;
assign dea74e = hbusreq2_p & deadd7 | !hbusreq2_p & deadd6;
assign b29fc3 = hlock0_p & b29fc2 | !hlock0_p & b29f9a;
assign b26773 = hlock2_p & b26713 | !hlock2_p & b26743;
assign a5fbb4 = hlock0_p & a5fbb2 | !hlock0_p & !a5fbb3;
assign v970409 = stateG10_1_p & v970408 | !stateG10_1_p & v9703fc;
assign a5fc44 = locked_p & a5fc43 | !locked_p & v84563c;
assign b29b17 = hmaster1_p & b29b16 | !hmaster1_p & b29a6e;
assign ab0c76 = hlock1_p & deada8 | !hlock1_p & ab0c75;
assign ab05c2 = hbusreq2_p & ab05c1 | !hbusreq2_p & ab05c0;
assign a5f96b = hready & v84566c | !hready & b266a0;
assign deae10 = hgrant2_p & dead39 | !hgrant2_p & deae0f;
assign a5ee5e = hready & a5ee5b | !hready & a5ee5d;
assign a5edc8 = hready & a5f531 | !hready & a5edc7;
assign a5fb2a = hready & v84563c | !hready & !cea29f;
assign ce9cf8 = hbusreq3 & cea14a | !hbusreq3 & v84563c;
assign d40d44 = hlock2_p & d40d43 | !hlock2_p & d40d42;
assign ab0736 = decide_p & ab0735 | !decide_p & v84563c;
assign a5f1da = hlock2_p & a5f1d9 | !hlock2_p & a5f979;
assign a5edff = hbusreq0_p & a5edf5 | !hbusreq0_p & a5edfb;
assign ab0621 = hgrant2_p & ab0620 | !hgrant2_p & cea15a;
assign a5fcd8 = hready & a5fcd5 | !hready & a5fcd7;
assign a5fcad = hgrant2_p & a5fc9c | !hgrant2_p & a5fcac;
assign cea2a4 = hready & cea0bc | !hready & cea29f;
assign ab05a0 = hmaster1_p & ab059f | !hmaster1_p & ab0b71;
assign a5f195 = hlock0_p & a5f8b9 | !hlock0_p & v84563c;
assign c3b7a6 = hlock0_p & c3bdf9 | !hlock0_p & v845660;
assign b29979 = hmaster1_p & b298a3 | !hmaster1_p & c3bceb;
assign ab0bfe = hready & b2a020 | !hready & !v84563c;
assign v970436 = hmaster1_p & v84563c | !hmaster1_p & v970435;
assign b29b23 = hbusreq2_p & b29b22 | !hbusreq2_p & v84563c;
assign a5f485 = hbusreq1_p & a5f9dd | !hbusreq1_p & v84563c;
assign cea3b9 = stateG10_1_p & deacb4 | !stateG10_1_p & cea3b8;
assign af34da = hbusreq2_p & af34d9 | !hbusreq2_p & af3c6b;
assign a5f544 = hready & v84563c | !hready & a5f543;
assign c3b885 = hgrant2_p & c3b7dc | !hgrant2_p & c3b884;
assign ab0c89 = hbusreq0_p & deace9 | !hbusreq0_p & c3bd8d;
assign b266be = hmaster0_p & b266b9 | !hmaster0_p & b266bd;
assign a5f9a7 = hlock0_p & a5f9a6 | !hlock0_p & v84563c;
assign b29827 = hlock0_p & b29826 | !hlock0_p & !v84563c;
assign a5fae5 = hbusreq2_p & a5fab4 | !hbusreq2_p & a5fab1;
assign cea8a0 = hbusreq2_p & cea889 | !hbusreq2_p & cea888;
assign a5fcdd = start_p & a5fba3 | !start_p & a5fcdc;
assign b2991c = hlock0_p & b2991b | !hlock0_p & !v84563c;
assign a5f8b8 = hready & a5f8b4 | !hready & a5f8b7;
assign ab056a = hlock0_p & ab0adc | !hlock0_p & !b29947;
assign cea236 = hlock2_p & cea235 | !hlock2_p & v84563c;
assign ce9d55 = hgrant2_p & cea15e | !hgrant2_p & !ce9d54;
assign ab0755 = hgrant2_p & ab06b5 | !hgrant2_p & ab0754;
assign c3b687 = hlock0_p & c3b67c | !hlock0_p & !c3b686;
assign a5fb98 = locked_p & a5fb97 | !locked_p & v84563c;
assign a5fc80 = hbusreq0_p & a5fc7a | !hbusreq0_p & !a5fc7f;
assign b29934 = hmaster1_p & b29933 | !hmaster1_p & b29e65;
assign ce9e29 = hbusreq3_p & ce9db0 | !hbusreq3_p & ce9e28;
assign v97044d = hgrant0_p & v970443 | !hgrant0_p & v97044c;
assign ab05d2 = hgrant2_p & ab05d1 | !hgrant2_p & cea15a;
assign ab06fa = hlock2 & ab06f8 | !hlock2 & ab06f9;
assign dea735 = hbusreq3 & dea734 | !hbusreq3 & !v84563c;
assign a5eaf2 = hbusreq0 & a5eaf1 | !hbusreq0 & !ab0c31;
assign ab0c0b = hlock2_p & ab0c03 | !hlock2_p & ab0c0a;
assign a5f0aa = hmaster1_p & a5f0a7 | !hmaster1_p & a5f0a9;
assign af3c80 = hlock0_p & af3c7d | !hlock0_p & af3c7f;
assign ce9cfd = hmaster0_p & ce9cf9 | !hmaster0_p & ce9cfc;
assign adaefc = hmaster0_p & adaefb | !hmaster0_p & adaed2;
assign a5f86d = hlock0_p & a5f864 | !hlock0_p & a5f86c;
assign dead63 = hgrant2_p & dead61 | !hgrant2_p & dead62;
assign dea73d = hbusreq2_p & deadb4 | !hbusreq2_p & !deadb2;
assign c3b715 = hready & c3b714 | !hready & c3bdce;
assign ab0c80 = hlock3_p & ab0c65 | !hlock3_p & ab0c7f;
assign a5eeb8 = hbusreq1 & a5eeb7 | !hbusreq1 & !v84563c;
assign ab052f = hlock0_p & v84563c | !hlock0_p & !cea3a9;
assign a5ee35 = hmaster1_p & a5ee0d | !hmaster1_p & a5ee34;
assign a5eb8e = hbusreq2 & a5f08b | !hbusreq2 & a5eb8d;
assign b2669b = hlock2_p & b2669a | !hlock2_p & b26699;
assign a5f1c8 = hlock0_p & a5f71e | !hlock0_p & a5f71d;
assign dead9e = hmaster0_p & dead98 | !hmaster0_p & dead9d;
assign a5f8e6 = hlock0_p & a5f8e5 | !hlock0_p & !v845641;
assign c3b613 = hready & deac7a | !hready & v845648;
assign ab05b8 = hgrant2_p & ab05b7 | !hgrant2_p & cea15a;
assign af3552 = hmaster1_p & af3541 | !hmaster1_p & af3551;
assign a5f9fa = hready & a5f9f6 | !hready & a5f9f9;
assign b2998a = hlock0_p & b29989 | !hlock0_p & !deae51;
assign ab05b1 = hlock0_p & b298a4 | !hlock0_p & ab05b0;
assign a5f455 = hmastlock_p & a5f828 | !hmastlock_p & v84563c;
assign a60144 = hbusreq2_p & a60143 | !hbusreq2_p & a60142;
assign a5fc79 = hready & a5fc78 | !hready & v84563c;
assign ab0b67 = hlock0_p & dead72 | !hlock0_p & !ab0b65;
assign a5f8cd = hbusreq2_p & a5f8cc | !hbusreq2_p & a5fad6;
assign ab069a = hlock2_p & ab0692 | !hlock2_p & ab0699;
assign a5f1e4 = hlock2 & a5f1de | !hlock2 & a5f1e3;
assign a5f3b9 = hlock0_p & a5f39e | !hlock0_p & a5f3b8;
assign ab058f = hready & deae4e | !hready & c3b6dd;
assign c3bcec = hbusreq3 & c3bce9 | !hbusreq3 & c3bceb;
assign b29abc = hlock0_p & b29abb | !hlock0_p & !b29e4d;
assign b29d4e = hlock3_p & b29d25 | !hlock3_p & b29d4d;
assign c3b7df = hbusreq2_p & c3b7dd | !hbusreq2_p & c3b7db;
assign cea3db = hlock1_p & v84565a | !hlock1_p & !cea3da;
assign b29f90 = hlock2 & dead35 | !hlock2 & b29f8f;
assign ab0c08 = locked_p & ab0c07 | !locked_p & !v84563c;
assign b298ae = locked_p & deae59 | !locked_p & !b29832;
assign a5ead5 = hbusreq2 & a5ead3 | !hbusreq2 & a5ead4;
assign a5f580 = hbusreq1 & a5f57e | !hbusreq1 & a5f57f;
assign b299a1 = hlock2 & b2999e | !hlock2 & b299a0;
assign a5e9b9 = hgrant1_p & a60168 | !hgrant1_p & a5f174;
assign a5f530 = hbusreq1_p & a60187 | !hbusreq1_p & v84563c;
assign b29ed6 = hbusreq3 & b29ed4 | !hbusreq3 & b29ed5;
assign cea446 = hbusreq2_p & cea445 | !hbusreq2_p & cea443;
assign c3b706 = hlock0_p & c3b705 | !hlock0_p & !c3b626;
assign ab0564 = hlock0_p & v84563c | !hlock0_p & !b29949;
assign ab0c92 = hlock2_p & ab0b95 | !hlock2_p & v84563c;
assign ab0671 = hlock2_p & ab066f | !hlock2_p & ab0670;
assign deadf2 = hgrant2_p & deadf0 | !hgrant2_p & deadf1;
assign c3bd61 = hbusreq0_p & c3bd5f | !hbusreq0_p & c3bd60;
assign b29f10 = hready & b29f0f | !hready & v84563c;
assign a5edb6 = hlock1_p & a5fa1c | !hlock1_p & a5f4ce;
assign a5f6f4 = hready & v84563c | !hready & !dead6e;
assign c3bdc1 = hlock2_p & c3bdc0 | !hlock2_p & !cea17a;
assign ab0525 = hbusreq2_p & ab0524 | !hbusreq2_p & ab0522;
assign cea14c = locked_p & v84563c | !locked_p & cea14b;
assign d40d56 = hmaster0_p & d40d48 | !hmaster0_p & d40d55;
assign a5f254 = hbusreq3 & a5f23c | !hbusreq3 & !a5f253;
assign deadb1 = hgrant1_p & deada9 | !hgrant1_p & deada8;
assign a5fd15 = hbusreq3 & a5fd10 | !hbusreq3 & v84563c;
assign a5e9d9 = hbusreq0 & a5f195 | !hbusreq0 & v845641;
assign b298a6 = hlock2_p & v84563c | !hlock2_p & b298a5;
assign cea451 = hmaster0_p & cea447 | !hmaster0_p & cea450;
assign a5fcf5 = hlock1_p & a5fbab | !hlock1_p & a5fcf4;
assign a5f8c9 = hlock2 & a5fa8b | !hlock2 & a5f8c8;
assign ab064f = hgrant0_p & bdb59e | !hgrant0_p & !ab064e;
assign a601a6 = hbusreq2_p & a6019b | !hbusreq2_p & a6019a;
assign cea3bc = hbusreq1_p & deaca1 | !hbusreq1_p & !v84565a;
assign c3bdd8 = hlock2_p & c3bdd7 | !hlock2_p & !deadba;
assign a5ee9c = locked_p & a5ee9b | !locked_p & a5f39e;
assign deae64 = hmaster1_p & deae63 | !hmaster1_p & v84563c;
assign a5f900 = hready & v84563c | !hready & a5f8ff;
assign b29fa1 = hlock0_p & dead41 | !hlock0_p & !b29fa0;
assign a9b9e6 = hgrant2_p & a9b9d0 | !hgrant2_p & !v84563c;
assign adaec9 = hlock1_p & adaec4 | !hlock1_p & adaec8;
assign af3c42 = hready_p & v8567b4 | !hready_p & af3c41;
assign ab05a4 = locked_p & ab05a3 | !locked_p & b2997c;
assign deae5a = hlock1_p & b26695 | !hlock1_p & !v845646;
assign ab05c9 = hmaster1_p & ab05c8 | !hmaster1_p & ab0bbb;
assign a5f907 = hlock0_p & a5f906 | !hlock0_p & ab0c31;
assign deae09 = hmaster1_p & dead2d | !hmaster1_p & deae08;
assign cea41e = hbusreq2_p & cea41d | !hbusreq2_p & cea3fb;
assign ab0541 = hbusreq2_p & ab0540 | !hbusreq2_p & ab053f;
assign cea193 = hmaster0_p & cea192 | !hmaster0_p & cea15d;
assign cea1b3 = hlock1_p & v84563c | !hlock1_p & !cea1b2;
assign dea72f = hbusreq3 & dea72d | !hbusreq3 & dea72e;
assign b29aea = hmaster1_p & b29ae9 | !hmaster1_p & b29a6e;
assign af3538 = hlock3_p & af3535 | !hlock3_p & af3537;
assign a5fb35 = hbusreq2_p & a5fb34 | !hbusreq2_p & v84563c;
assign af352d = locked_p & af352c | !locked_p & v84563c;
assign a5f3d7 = hready & a5f3d4 | !hready & a5f3d6;
assign c3b8b3 = hmaster1_p & c3b8af | !hmaster1_p & c3b8b2;
assign a5fc03 = locked_p & a5fc02 | !locked_p & v84563c;
assign a5efcc = hmaster0_p & a5efcb | !hmaster0_p & a5eed3;
assign a5ea96 = hbusreq0_p & a5fcab | !hbusreq0_p & v84563c;
assign cea38b = hlock0_p & cea389 | !hlock0_p & cea38a;
assign a5eef7 = hgrant2_p & a5eef3 | !hgrant2_p & a5eef6;
assign a5f6ee = hready & a5f9dd | !hready & !dead6e;
assign cea406 = hbusreq2_p & cea3fc | !hbusreq2_p & cea405;
assign deae14 = hbusreq2_p & deae13 | !hbusreq2_p & dead39;
assign deac1e = hlock0_p & deac19 | !hlock0_p & v84565a;
assign dea6c1 = hmaster1_p & dea6c0 | !hmaster1_p & dead3c;
assign a5efe3 = hbusreq2_p & a5f568 | !hbusreq2_p & a5ef84;
assign a5ea0f = hbusreq2_p & a5ea0e | !hbusreq2_p & v845641;
assign cea273 = hlock1_p & v84563c | !hlock1_p & !cea272;
assign a5f994 = hready & v84563c | !hready & !dead7b;
assign a5efb2 = hbusreq2 & a5efb1 | !hbusreq2 & a5ee26;
assign deae28 = hbusreq3 & deae27 | !hbusreq3 & deae25;
assign cea3a8 = hbusreq3 & cea3a4 | !hbusreq3 & !cea3a7;
assign dea727 = hbusreq2_p & dea726 | !hbusreq2_p & dea724;
assign b299ae = hbusreq2_p & b299ad | !hbusreq2_p & v84563c;
assign a5ede6 = hbusreq1_p & a5fb8b | !hbusreq1_p & v84563c;
assign dea6da = hlock3_p & dea6d9 | !hlock3_p & deaeaa;
assign b29d87 = hready & deacdf | !hready & b266a0;
assign c3b776 = decide_p & c3b775 | !decide_p & v845660;
assign ab0cea = hmaster0_p & ab0ce9 | !hmaster0_p & ab0c90;
assign c3b7ed = hmaster1_p & c3b7ec | !hmaster1_p & c3bcd2;
assign v970446 = locked_p & v970445 | !locked_p & v84563c;
assign a5f8db = stateA1_p & a60184 | !stateA1_p & a5f8da;
assign c3bcdb = hready & b26695 | !hready & v84563c;
assign ce9cd8 = hgrant0_p & v84563c | !hgrant0_p & cea178;
assign ab0590 = locked_p & ab058f | !locked_p & !b29832;
assign ab0597 = hmaster0_p & ab058c | !hmaster0_p & ab0596;
assign ab0c62 = hbusreq2_p & ab0c60 | !hbusreq2_p & ab0b21;
assign a5efc7 = hmaster1_p & a5f3d8 | !hmaster1_p & v84563c;
assign c3b697 = hlock1_p & deac52 | !hlock1_p & v84563c;
assign a5fb5f = hlock2_p & a5fb5e | !hlock2_p & a5fad6;
assign a5f160 = hbusreq2_p & a5f14d | !hbusreq2_p & a5f145;
assign v970434 = locked_p & v970413 | !locked_p & v84563c;
assign b29cd5 = hbusreq2_p & b29cd4 | !hbusreq2_p & deacab;
assign a5eeb1 = hgrant2_p & a5eeb0 | !hgrant2_p & v84563c;
assign af3c7d = hlock1_p & af3c49 | !hlock1_p & !d40d3d;
assign a5ea40 = hbusreq0_p & a5fc56 | !hbusreq0_p & v84563c;
assign b29a84 = hready & b29a83 | !hready & c3bdce;
assign bdb589 = hgrant2_p & bdb587 | !hgrant2_p & bdb588;
assign ab0bdc = hmaster1_p & ab0bd7 | !hmaster1_p & !ab0bdb;
assign a5f882 = hlock2 & a5fafd | !hlock2 & a5f881;
assign c3bd00 = hmaster1_p & c3bcfc | !hmaster1_p & c3bcff;
assign v970451 = hlock3_p & v970450 | !hlock3_p & v97042d;
assign cea3a1 = hbusreq2_p & cea3a0 | !hbusreq2_p & cea39f;
assign a5eee3 = hready & a5eee2 | !hready & a5f43f;
assign a5fbb1 = hready & a5fba8 | !hready & a5fbb0;
assign a5f2e3 = hready & a5fb81 | !hready & !b26734;
assign c3bbc0 = hlock3_p & c3bbbf | !hlock3_p & !v84563c;
assign a5fa02 = hlock2 & a5f9e9 | !hlock2 & a5fa01;
assign b2a000 = hmaster1_p & b29fff | !hmaster1_p & b29f8b;
assign ab0ae5 = hmaster1_p & ab0ad2 | !hmaster1_p & ab0ae4;
assign a60195 = hbusreq1 & a60169 | !hbusreq1 & a60194;
assign ab06eb = hlock0_p & b2a002 | !hlock0_p & v845660;
assign c3bc07 = hbusreq3 & c3bbfe | !hbusreq3 & c3bc06;
assign a5f567 = hbusreq2 & a5f561 | !hbusreq2 & a5f566;
assign cea155 = hbusreq2_p & cea154 | !hbusreq2_p & cea153;
assign a5f471 = hbusreq1 & a5f470 | !hbusreq1 & v84565a;
assign b29eb2 = hbusreq2_p & b29eb1 | !hbusreq2_p & v84563c;
assign c3bd4f = hbusreq2_p & c3bd4d | !hbusreq2_p & c3bbe8;
assign a5fbd6 = hbusreq3 & a5fbce | !hbusreq3 & a5fbd5;
assign ab0685 = hbusreq3 & ab0684 | !hbusreq3 & !v84563c;
assign c3b79a = hbusreq2_p & c3b799 | !hbusreq2_p & c3b797;
assign ab0c06 = hlock0_p & v84563c | !hlock0_p & !ab0c05;
assign cea378 = hready & v8c6711 | !hready & v845646;
assign adaf13 = hmaster0_p & adaf12 | !hmaster0_p & v84563c;
assign af3c3c = hmaster0_p & af3c3b | !hmaster0_p & af3c23;
assign ab0b3b = hlock0_p & v84563c | !hlock0_p & deacbe;
assign b29d50 = hready_p & b29cba | !hready_p & b29d4f;
assign c3b889 = hready_p & c3b878 | !hready_p & c3b888;
assign a5f98a = hlock1_p & a5fc84 | !hlock1_p & a5f989;
assign a5edf0 = hbusreq1 & a5edef | !hbusreq1 & !v84563c;
assign ab0acf = hlock3_p & ab0ace | !hlock3_p & v84563c;
assign a5eadf = hbusreq0 & a5ead7 | !hbusreq0 & a5eade;
assign af35b9 = hmaster0_p & af35b8 | !hmaster0_p & af3567;
assign c3bc2e = hmaster1_p & c3bc10 | !hmaster1_p & c3bc2d;
assign b29d9a = hmaster0_p & b29d75 | !hmaster0_p & b29d99;
assign af3558 = hlock2_p & af3541 | !hlock2_p & v84563c;
assign a5f09b = hlock0_p & a5f6e9 | !hlock0_p & v84563c;
assign deae50 = hlock1_p & dead6e | !hlock1_p & dead76;
assign af3550 = hbusreq2_p & af354e | !hbusreq2_p & af354d;
assign b29ec8 = hlock2_p & b29ec7 | !hlock2_p & v845660;
assign a5f41f = hlock0_p & a5f41e | !hlock0_p & a5f40d;
assign b29ce7 = hlock0_p & deac52 | !hlock0_p & !v84563c;
assign a5fba9 = stateA1_p & a81ca7 | !stateA1_p & c07311;
assign a5f0d1 = hlock0_p & a5f0c3 | !hlock0_p & a5f0d0;
assign af359f = hgrant0_p & af3599 | !hgrant0_p & af359e;
assign b29d6f = locked_p & b29d6d | !locked_p & b29d6e;
assign a5f6eb = hlock0_p & a5f6e8 | !hlock0_p & a5f6ea;
assign ab06f0 = hgrant0_p & ab0be1 | !hgrant0_p & !ab06ef;
assign ab0cb7 = hgrant2_p & ab0bba | !hgrant2_p & ab0ca2;
assign ab052e = hbusreq3 & ab052a | !hbusreq3 & ab052d;
assign cea887 = hlock1_p & deada8 | !hlock1_p & v84563c;
assign b29a7c = hlock2 & b29ce7 | !hlock2 & b29a7b;
assign b299d4 = hmaster0_p & b299d3 | !hmaster0_p & b29974;
assign b29985 = hready & deae50 | !hready & v84563c;
assign ab0554 = hgrant2_p & ab0550 | !hgrant2_p & ab0553;
assign a5f515 = hbusreq1 & a5f485 | !hbusreq1 & v84563c;
assign b29fc0 = hlock1_p & v84563c | !hlock1_p & c3bdbb;
assign deade3 = hbusreq2_p & deade1 | !hbusreq2_p & !deacab;
assign cea0c0 = hbusreq2_p & cea86d | !hbusreq2_p & !cea0bf;
assign ab0c0d = hbusreq3 & ab0c02 | !hbusreq3 & ab0c0c;
assign af35af = hmaster0_p & af35aa | !hmaster0_p & af3589;
assign a5ebee = hbusreq3_p & a5eb49 | !hbusreq3_p & a5ebed;
assign c3b628 = hlock2_p & c3b627 | !hlock2_p & !c3b626;
assign a5f3be = hbusreq2_p & a5f3bd | !hbusreq2_p & a5f3b9;
assign b29f8c = hmaster1_p & b29f88 | !hmaster1_p & b29f8b;
assign a5fa5a = hready & a5fa59 | !hready & !c3bdce;
assign b29d59 = hlock2_p & v84563c | !hlock2_p & b29d58;
assign b299e4 = hmaster0_p & b299e3 | !hmaster0_p & b29998;
assign a5fc11 = locked_p & a5fc10 | !locked_p & !v84563c;
assign b29ed8 = hbusreq2_p & b29ed7 | !hbusreq2_p & v84563c;
assign a5f11d = stateG10_1_p & a5f11c | !stateG10_1_p & a5f11b;
assign d40d2c = locked_p & d40d2b | !locked_p & v84563c;
assign a5fba1 = start_p & a6016a | !start_p & a5fba0;
assign a5ee0f = hlock1_p & v84563c | !hlock1_p & ab05a1;
assign a5f18c = hlock1_p & a60177 | !hlock1_p & !a5f18b;
assign cea47d = hlock2_p & cea47c | !hlock2_p & cea3cd;
assign ab0b55 = hlock0_p & v845660 | !hlock0_p & b29d51;
assign a81cef = start_p & v84563c | !start_p & !v845672;
assign c3bcd3 = hmaster1_p & c3bcd1 | !hmaster1_p & c3bcd2;
assign cea0ee = hbusreq3 & v84563c | !hbusreq3 & cea877;
assign cea18d = locked_p & v845648 | !locked_p & !v84563c;
assign a5f377 = hbusreq1_p & v970408 | !hbusreq1_p & v84563c;
assign a5f138 = hbusreq2_p & a5f0ec | !hbusreq2_p & a5f0e6;
assign ab060d = hlock0_p & v84563c | !hlock0_p & b29992;
assign a5f0a5 = hbusreq0_p & a5fc89 | !hbusreq0_p & !v84563c;
assign b29a3e = hbusreq2_p & b29a3d | !hbusreq2_p & v84563c;
assign dea750 = hgrant2_p & dea74c | !hgrant2_p & dea74f;
assign stateG3_2 = !d40d9d;
assign a5fbdf = stateA1_p & a5fb9d | !stateA1_p & !a5fb87;
assign a5f8c2 = hgrant1_p & v84563c | !hgrant1_p & b29914;
assign c3b82d = hmaster0_p & c3b823 | !hmaster0_p & c3b82c;
assign ce9dd3 = hbusreq2_p & cea2b0 | !hbusreq2_p & ce9dc8;
assign ab06dd = hgrant2_p & ab06db | !hgrant2_p & ab06dc;
assign c3bd91 = hbusreq2_p & c3bd90 | !hbusreq2_p & c3bc5c;
assign b266e2 = hlock2_p & b266e1 | !hlock2_p & b266e0;
assign ab0b8a = hlock0_p & v84563c | !hlock0_p & !ab0b89;
assign a5f587 = hbusreq2_p & a5f583 | !hbusreq2_p & a5f577;
assign dea6e2 = hbusreq3 & dea6e1 | !hbusreq3 & deae62;
assign af3580 = locked_p & af357f | !locked_p & v84563c;
assign b29c3c = hbusreq2_p & b29c3b | !hbusreq2_p & v84563c;
assign a5f8f2 = hbusreq0 & a5f8cd | !hbusreq0 & !a5f8f1;
assign deae25 = hbusreq2_p & deae24 | !hbusreq2_p & v84563c;
assign b840b1 = hgrant0_p & v845643 | !hgrant0_p & b840b0;
assign c3bc79 = locked_p & v845648 | !locked_p & dead0a;
assign dea6c4 = hmaster1_p & dea6c3 | !hmaster1_p & dea6c0;
assign d40d85 = hmaster1_p & d40d60 | !hmaster1_p & d40d84;
assign a5fc9f = hbusreq1_p & a5fc84 | !hbusreq1_p & a5fc8c;
assign a5f162 = hbusreq0 & a5f160 | !hbusreq0 & a5f161;
assign cea36c = hgrant2_p & cea368 | !hgrant2_p & cea36b;
assign af34bd = hlock2_p & af34bc | !hlock2_p & af34bb;
assign a5fb66 = hmaster0_p & a5fb03 | !hmaster0_p & a5fb65;
assign c3bd73 = hmaster1_p & c3bd6d | !hmaster1_p & c3bd72;
assign a5ef78 = hlock2 & a5ef5f | !hlock2 & a5f36e;
assign a5eb39 = hbusreq0_p & a5fd00 | !hbusreq0_p & v84563c;
assign b29e53 = hmaster1_p & b29e52 | !hmaster1_p & !b29e4a;
assign d40d7a = start_p & v84563c | !start_p & bfbd19;
assign c3b71b = hlock1_p & v84563c | !hlock1_p & !c3b71a;
assign a5ec33 = jx2_p & a5f363 | !jx2_p & a5ec32;
assign a5ee11 = hready & a5f365 | !hready & a5ee10;
assign ab0cf7 = hbusreq2_p & ab0c6d | !hbusreq2_p & ab0b0e;
assign a5f012 = hready_p & a5efce | !hready_p & a5f011;
assign ab0b7a = hlock0_p & v84563c | !hlock0_p & ab0b79;
assign dea6bd = hmaster1_p & deaeb5 | !hmaster1_p & dea6bc;
assign ab0b46 = hlock2_p & ab0b45 | !hlock2_p & ab0b23;
assign c3b81c = hgrant2_p & c3b81b | !hgrant2_p & c3b7a5;
assign b2992d = hlock2_p & v84563c | !hlock2_p & !b2992c;
assign ab05be = hbusreq2_p & ab0589 | !hbusreq2_p & ab05bd;
assign c3b6b8 = hbusreq3 & c3b698 | !hbusreq3 & c3b6a1;
assign a5ef36 = locked_p & a60140 | !locked_p & a5ef35;
assign a5f1a4 = hlock0_p & v84563c | !hlock0_p & a5f1a3;
assign b299d8 = hlock0_p & b299d7 | !hlock0_p & v84563c;
assign a5efc4 = hmaster1_p & a5efbd | !hmaster1_p & a5efc3;
assign a5f2de = decide_p & a5f2d6 | !decide_p & !a5f2dd;
assign a5f95f = hready_p & a5f757 | !hready_p & a5f95e;
assign a81ccc = hready_p & a81cae | !hready_p & a81ccb;
assign a5ea74 = hbusreq0 & a5ea73 | !hbusreq0 & a5ea3e;
assign b2671c = hmaster0_p & b26712 | !hmaster0_p & b2671b;
assign dead17 = hbusreq3 & dead16 | !hbusreq3 & v84563c;
assign b26704 = hbusreq2_p & b26703 | !hbusreq2_p & !b266a0;
assign b2674b = hmaster1_p & b26748 | !hmaster1_p & b2674a;
assign dead02 = hmaster1_p & deacf0 | !hmaster1_p & dead01;
assign a5fce9 = hbusreq3 & a5fce8 | !hbusreq3 & v84563c;
assign b2998d = hlock0_p & b2998c | !hlock0_p & !v84563c;
assign ab05e5 = hbusreq3 & ab052a | !hbusreq3 & ab05e4;
assign dead53 = hbusreq2_p & v84563c | !hbusreq2_p & v845644;
assign af3c79 = stateG10_1_p & d40d33 | !stateG10_1_p & af3c49;
assign a5eed5 = hgrant0_p & a5eec9 | !hgrant0_p & a5eed4;
assign a5eb8a = hready_p & a5eb54 | !hready_p & a5eb89;
assign cea0ba = hbusreq1_p & v84565a | !hbusreq1_p & !v84563c;
assign b299f4 = decide_p & b299f3 | !decide_p & v84563c;
assign ab064c = hgrant0_p & ab0be1 | !hgrant0_p & !ab0b71;
assign ab0af6 = hlock0_p & v84563c | !hlock0_p & !v84565a;
assign deacc5 = hlock0_p & deaca1 | !hlock0_p & v84563c;
assign a5ea1a = hgrant2_p & a5ea10 | !hgrant2_p & a5ea19;
assign b266ad = locked_p & v84563c | !locked_p & b266ac;
assign cea169 = hbusreq3 & cea168 | !hbusreq3 & cea159;
assign a5f3b4 = hready & a5f38c | !hready & !a5f3b3;
assign af359a = hgrant2_p & af356f | !hgrant2_p & af352d;
assign a5fa22 = hlock0_p & a5fa16 | !hlock0_p & !a5fa21;
assign af3c11 = locked_p & v845646 | !locked_p & v8c6711;
assign ab0c3e = hlock0_p & v84563c | !hlock0_p & ab0c3d;
assign dea6ef = hgrant3_p & dea6ee | !hgrant3_p & !v84563c;
assign a5f3ae = hmaster1_p & a5f3ad | !hmaster1_p & v84563c;
assign v84564f = hbusreq3 & v84563c | !hbusreq3 & !v84563c;
assign a5ee45 = locked_p & a5ee44 | !locked_p & a60140;
assign af3536 = hmaster1_p & v84563c | !hmaster1_p & af352f;
assign b29fb9 = hlock2_p & b29fb8 | !hlock2_p & !b29f90;
assign c3bde8 = hmaster1_p & c3bcb4 | !hmaster1_p & c3bd05;
assign a5f436 = hgrant1_p & a5f435 | !hgrant1_p & a5f434;
assign ab0c05 = locked_p & ab0c04 | !locked_p & !v84563c;
assign d40d68 = locked_p & d40d67 | !locked_p & v84563c;
assign ab0b99 = hbusreq3 & ab0b98 | !hbusreq3 & cea15a;
assign a5fc4d = hmaster1_p & v84563c | !hmaster1_p & a5fc4c;
assign a5f5a9 = hlock0_p & a5f5a8 | !hlock0_p & a5f4b8;
assign cea2a6 = hlock2_p & cea2a5 | !hlock2_p & v84563c;
assign ab052b = hlock0_p & v84563c | !hlock0_p & b29832;
assign deacb8 = hbusreq2_p & deacb7 | !hbusreq2_p & v84563c;
assign a5eeee = hready & a5eee8 | !hready & a5f471;
assign ab063d = hgrant3_p & ab0602 | !hgrant3_p & !ab063c;
assign ab071a = hbusreq2_p & ab0713 | !hbusreq2_p & ab06b8;
assign ab0acb = hlock0_p & b298a4 | !hlock0_p & v845660;
assign ab0bf3 = hgrant2_p & ab0bf2 | !hgrant2_p & ab0b30;
assign af3496 = hlock3_p & af3490 | !hlock3_p & af3495;
assign a5ef82 = hlock0_p & a5f560 | !hlock0_p & a5ef81;
assign cea359 = hmaster1_p & cea358 | !hmaster1_p & cea1c4;
assign d40d6b = hmaster1_p & v84563c | !hmaster1_p & d40d6a;
assign ce9d31 = hbusreq2_p & cea2a6 | !hbusreq2_p & cea2a5;
assign a5f1d8 = hlock0_p & a5f1d7 | !hlock0_p & a5f72b;
assign cea1bb = hmastlock_p & cea1ba | !hmastlock_p & v84563c;
assign a5ea58 = hlock1_p & a5fc84 | !hlock1_p & a5ea57;
assign a5f87b = hbusreq2 & a5f86d | !hbusreq2 & a5f87a;
assign ab0b15 = hready & deae1d | !hready & c3bd5d;
assign c3b6ad = hgrant2_p & c3b6a3 | !hgrant2_p & c3b6ac;
assign v970455 = hmaster1_p & v97043f | !hmaster1_p & v84563c;
assign a5eecf = hbusreq2_p & a5eecd | !hbusreq2_p & !a5eece;
assign ab0b19 = hbusreq2_p & ab0b18 | !hbusreq2_p & !ab0b17;
assign a5ea7a = hmaster1_p & a5ea70 | !hmaster1_p & a5ea79;
assign ce9e0c = decide_p & ce9e0b | !decide_p & a57859;
assign c3b692 = stateG10_1_p & deacb4 | !stateG10_1_p & c3b691;
assign c3bd84 = hlock2_p & c3bd83 | !hlock2_p & dead2e;
assign cea33f = hready_p & cea32f | !hready_p & cea33e;
assign ab075d = hready_p & ab074d | !hready_p & !ab075c;
assign v970459 = hready_p & v970457 | !hready_p & v970458;
assign a5ee09 = hlock2_p & a5ee05 | !hlock2_p & a5ee08;
assign a5eebe = hlock0_p & a5f3c9 | !hlock0_p & a5eebd;
assign b266c4 = decide_p & b266bf | !decide_p & b266c3;
assign a5fb8b = hmastlock_p & deacf4 | !hmastlock_p & v84563c;
assign a5f94d = hbusreq0 & a5f94c | !hbusreq0 & a5f94a;
assign a5fa88 = hready & a60168 | !hready & a5fa87;
assign a5f287 = hgrant2_p & v84563c | !hgrant2_p & a5f95b;
assign ab05e9 = hbusreq3 & ab052f | !hbusreq3 & ab05e8;
assign d615cf = stateG3_1_p & v84563c | !stateG3_1_p & !v845670;
assign a5fca9 = hlock1_p & v84563c | !hlock1_p & a5fca8;
assign ab0651 = decide_p & ab0650 | !decide_p & v845662;
assign v845662 = hgrant0_p & v84563c | !hgrant0_p & !v84563c;
assign ab06f9 = hlock0_p & b29fb5 | !hlock0_p & !dead34;
assign cea27b = hgrant2_p & cea278 | !hgrant2_p & cea27a;
assign b29f40 = hready & deaca2 | !hready & !v84563c;
assign deaddf = hlock1_p & deadde | !hlock1_p & !deadd4;
assign dea78a = hmaster1_p & dea789 | !hmaster1_p & !v84563c;
assign ab0c21 = hlock2_p & ab0c20 | !hlock2_p & v84563c;
assign a5f8f7 = hmaster1_p & a5f6db | !hmaster1_p & a5f8f6;
assign deadb9 = start_p & v845652 | !start_p & !v8c6449;
assign a5f360 = hready_p & a5f306 | !hready_p & a5f35f;
assign a5ebe7 = hgrant2_p & a5ebdd | !hgrant2_p & a5ebe6;
assign af3c38 = hgrant0_p & v8567b4 | !hgrant0_p & af3c37;
assign a5f1f1 = hlock1_p & a5fc0d | !hlock1_p & !v84563c;
assign ab0618 = hbusreq0_p & b29993 | !hbusreq0_p & ab0617;
assign a5fad5 = hlock0_p & v84563c | !hlock0_p & a5fad4;
assign adaeeb = locked_p & adaeea | !locked_p & v84563c;
assign c3b7ac = hbusreq3 & c3b7ab | !hbusreq3 & dead39;
assign d40d3e = hlock1_p & d40d31 | !hlock1_p & !d40d3d;
assign a5fc17 = hlock0_p & v845641 | !hlock0_p & a5fbc0;
assign c3b6eb = hmaster1_p & c3b6ea | !hmaster1_p & c3bcc0;
assign b2994e = hready & b2994d | !hready & !v84563c;
assign cea29f = hlock1_p & v84563c | !hlock1_p & !c98b95;
assign ab0623 = hmaster0_p & ab0616 | !hmaster0_p & ab0622;
assign a5f932 = hlock1_p & a60168 | !hlock1_p & a5f931;
assign v97045d = hbusreq3_p & v970454 | !hbusreq3_p & v97045c;
assign b29e68 = hlock2 & b29e67 | !hlock2 & b29d34;
assign c3b7fd = hgrant2_p & c3b7f9 | !hgrant2_p & c3b7fc;
assign a5f934 = hlock0_p & a5f933 | !hlock0_p & v845641;
assign a81d08 = decide_p & a81cc6 | !decide_p & a81d07;
assign b29d24 = hmaster1_p & b29d07 | !hmaster1_p & !b29d23;
assign cea424 = hbusreq2_p & cea41d | !hbusreq2_p & cea41c;
assign c3bc6e = hlock0_p & v845648 | !hlock0_p & v845660;
assign b298b3 = hmaster1_p & b298b2 | !hmaster1_p & v84563c;
assign a5e9b5 = hlock0_p & a5e9b3 | !hlock0_p & a5e9b4;
assign a5fd02 = hgrant2_p & a5fcf1 | !hgrant2_p & a5fd01;
assign cea3b7 = hmastlock_p & cea24f | !hmastlock_p & v84563c;
assign cea2eb = hlock2_p & cea2ea | !hlock2_p & v84563c;
assign a5f4cc = hbusreq1_p & v9703fb | !hbusreq1_p & v84563c;
assign ce9cbe = decide_p & ce9cbd | !decide_p & a57859;
assign af3c25 = hgrant2_p & af3c1a | !hgrant2_p & v845646;
assign ce9d4a = hgrant2_p & cea15e | !hgrant2_p & !ce9d49;
assign a5f06d = hlock2_p & a5f068 | !hlock2_p & a5f06c;
assign a5ee15 = hlock0_p & a5ee12 | !hlock0_p & a5ee14;
assign a5fa0f = hbusreq1_p & a60187 | !hbusreq1_p & !a6016f;
assign b26728 = hlock1_p & b26693 | !hlock1_p & b26727;
assign ab0642 = hmaster0_p & ab063f | !hmaster0_p & ab0641;
assign a5f9e1 = hready & a5f9e0 | !hready & !c3bd16;
assign b29e72 = hready_p & b29e5f | !hready_p & b29e71;
assign deacf6 = hburst0 & deacf4 | !hburst0 & deacf5;
assign adaee6 = hmaster1_p & adaee5 | !hmaster1_p & v84563c;
assign a5f17e = hlock2 & a5f172 | !hlock2 & a5f17d;
assign c3b712 = stateG10_1_p & deada8 | !stateG10_1_p & c3b661;
assign a5ef97 = locked_p & v84563c | !locked_p & a5ef35;
assign c3bcee = locked_p & v84563c | !locked_p & !c3bcdb;
assign a5f70b = hready & a5f704 | !hready & v970408;
assign a5f9c2 = hready & v84563c | !hready & c98b96;
assign cea40e = hready & c98b96 | !hready & c98b95;
assign ab0c10 = hbusreq2_p & ab0c0f | !hbusreq2_p & ab0acb;
assign a5fd1c = hgrant3_p & a5fb69 | !hgrant3_p & a5fd1b;
assign deae4b = hbusreq3_p & deae2f | !hbusreq3_p & deae4a;
assign a5efe7 = hbusreq2_p & a5f568 | !hbusreq2_p & a5efe6;
assign ab055f = hlock0_p & v84563c | !hlock0_p & !ab055e;
assign cea46e = hbusreq2_p & cea46d | !hbusreq2_p & cea44a;
assign c3bdc0 = hlock0_p & c3bdbf | !hlock0_p & !c3bd9b;
assign a5f494 = hbusreq1 & c3b6bd | !hbusreq1 & !a5f493;
assign af3505 = hmaster1_p & af3c4c | !hmaster1_p & af3c58;
assign a5eeb6 = hmaster1_p & a5f3d2 | !hmaster1_p & v84563c;
assign b8acee = decide_p & b8ace8 | !decide_p & b8aced;
assign a5f57c = hbusreq1 & a5f57b | !hbusreq1 & v84563c;
assign d40d90 = hmaster1_p & d40d7b | !hmaster1_p & d40d60;
assign ce9d10 = hlock0_p & deacec | !hlock0_p & v84563c;
assign c3b77f = hbusreq3_p & c3b77e | !hbusreq3_p & !c3bcd7;
assign af3573 = hbusreq0_p & v84563c | !hbusreq0_p & af3571;
assign c98ba1 = hgrant0_p & v8c6711 | !hgrant0_p & c98ba0;
assign ab0757 = hbusreq2_p & ab06a4 | !hbusreq2_p & ab0756;
assign cea39b = locked_p & deae59 | !locked_p & cea37b;
assign c3bc0f = hbusreq3 & c3bc0c | !hbusreq3 & c3bc0e;
assign af35bb = hmaster0_p & af35ba | !hmaster0_p & af3598;
assign v970447 = hgrant2_p & v84563c | !hgrant2_p & v970446;
assign a5ef2b = hgrant2_p & a5ef2a | !hgrant2_p & v84563c;
assign a5ef89 = hlock0_p & a5edd4 | !hlock0_p & a5ef81;
assign cea255 = hbusreq1_p & deaca1 | !hbusreq1_p & !v84563c;
assign ab0ca4 = hmaster1_p & ab0b71 | !hmaster1_p & ab0ca3;
assign a5fcdc = stateA1_p & a60174 | !stateA1_p & !cea24b;
assign b29a40 = hlock0_p & c3bce6 | !hlock0_p & v84563c;
assign a5f00f = hmaster0_p & a5f00e | !hmaster0_p & a5ef2e;
assign adaef5 = hbusreq2_p & adaebd | !hbusreq2_p & adaeeb;
assign a5ef09 = hbusreq1 & a5ef08 | !hbusreq1 & !v84563c;
assign ce9cfb = hbusreq3 & ce9cfa | !hbusreq3 & v84563c;
assign b26718 = hlock0_p & b26699 | !hlock0_p & b26716;
assign ce9d46 = hlock0_p & cea2f1 | !hlock0_p & !cea17a;
assign cea438 = hgrant2_p & cea432 | !hgrant2_p & cea437;
assign af34c9 = hbusreq2_p & af34c8 | !hbusreq2_p & af34c7;
assign c3b683 = hmastlock_p & deadb9 | !hmastlock_p & !v84563c;
assign cea31a = hbusreq2_p & cea2eb | !hbusreq2_p & v84563c;
assign a5efe2 = hgrant2_p & a5efdd | !hgrant2_p & a5efe1;
assign v9703fa = stateA1_p & v84566e | !stateA1_p & !v84563c;
assign b29fe1 = hbusreq2_p & b29fe0 | !hbusreq2_p & v84563c;
assign b26733 = hbusreq2_p & b26732 | !hbusreq2_p & !b26715;
assign a5fcc9 = hbusreq3 & a5fcc8 | !hbusreq3 & v84563c;
assign a5f9f9 = hlock1_p & a60172 | !hlock1_p & a5f9f8;
assign a5f939 = hready & v84563c | !hready & a5f938;
assign b29825 = hready & b29824 | !hready & !deaeb6;
assign a5fbf9 = start_p & v84563c | !start_p & a5fb87;
assign cea8a9 = hbusreq1_p & deadde | !hbusreq1_p & !v84563c;
assign ab0b82 = hbusreq2_p & ab0b81 | !hbusreq2_p & v84563c;
assign a5f087 = hmaster1_p & a5f07d | !hmaster1_p & a5f086;
assign dead68 = decide_p & dead67 | !decide_p & v84563c;
assign a5f943 = hready & a5f942 | !hready & a5f8d2;
assign cea2e6 = hbusreq1_p & cea2e5 | !hbusreq1_p & v84563c;
assign cea256 = hgrant1_p & deacb5 | !hgrant1_p & cea255;
assign b29a56 = hmaster0_p & b29a51 | !hmaster0_p & b29a55;
assign c3b6bc = hgrant1_p & c3b692 | !hgrant1_p & c3b691;
assign a5fa2d = hready & v84563c | !hready & !v84565a;
assign ab0744 = hgrant2_p & ab0741 | !hgrant2_p & ab0743;
assign a5fb9d = stateG2_p & v84563c | !stateG2_p & d615cf;
assign deaeaf = hlock0_p & deaeae | !hlock0_p & v84563c;
assign ab0bb0 = hbusreq2_p & ab0baf | !hbusreq2_p & v84563c;
assign af34f3 = locked_p & af3c49 | !locked_p & d40d82;
assign a5fc39 = hlock2_p & a5fc38 | !hlock2_p & v84563c;
assign b29ed3 = hlock2_p & c3bcf8 | !hlock2_p & !v84563c;
assign ab06e8 = hlock2 & ab066b | !hlock2 & ab06e7;
assign a5f71b = hbusreq3 & a5f6fd | !hbusreq3 & !a5f71a;
assign ab0560 = hlock2 & ab053f | !hlock2 & ab055f;
assign cea380 = hready & v8c6711 | !hready & !v84563c;
assign b29a1f = hready_p & b29a1d | !hready_p & b29a1e;
assign af34a8 = hlock2_p & af34a6 | !hlock2_p & af34a7;
assign b299ff = hgrant0_p & c3bceb | !hgrant0_p & !b29d64;
assign ab06b6 = hbusreq2_p & ab06b4 | !hbusreq2_p & ab06b5;
assign dead87 = hmaster1_p & deac0f | !hmaster1_p & dead85;
assign a81cc6 = hmaster0_p & a81cc5 | !hmaster0_p & a81cc3;
assign dead12 = hgrant2_p & dead07 | !hgrant2_p & dead11;
assign b8ace7 = hmaster0_p & b8ace6 | !hmaster0_p & b8ace5;
assign cea1b6 = hlock0_p & cea1b5 | !hlock0_p & v84563c;
assign ab0ce4 = decide_p & ab0ce3 | !decide_p & v84563c;
assign ce9d12 = hbusreq3 & ce9d11 | !hbusreq3 & v84563c;
assign af35b2 = hgrant0_p & af35af | !hgrant0_p & af35b1;
assign b29a8e = hlock2_p & v84563c | !hlock2_p & !c3bc21;
assign a5f3cd = hbusreq1 & a5f3cc | !hbusreq1 & !v84563c;
assign a5ef13 = locked_p & a5ef12 | !locked_p & v84563c;
assign cea3ef = hbusreq2_p & cea3cf | !hbusreq2_p & cea3ce;
assign a5fc3e = hbusreq3 & a5fc3d | !hbusreq3 & v84563c;
assign b29f0c = stateG10_1_p & b29f06 | !stateG10_1_p & b29f0b;
assign ab0b34 = hmaster0_p & ab0ae5 | !hmaster0_p & ab0b33;
assign af34fe = decide_p & af3495 | !decide_p & af3499;
assign a5e9f1 = hready & a5f9e7 | !hready & c3bbfb;
assign b29cdb = hmaster1_p & b29cc1 | !hmaster1_p & b29cda;
assign deae7a = hlock2_p & deae79 | !hlock2_p & !deadb2;
assign a5f785 = hgrant1_p & deac52 | !hgrant1_p & a5f784;
assign a5f3c3 = hbusreq1_p & a5fc78 | !hbusreq1_p & v84563c;
assign c3b653 = hbusreq2_p & c3b652 | !hbusreq2_p & c3b651;
assign cea321 = hbusreq1_p & v84566c | !hbusreq1_p & !cea320;
assign ab0ba6 = hlock0_p & v84563c | !hlock0_p & ab0ba5;
assign a5f8cf = hbusreq1_p & a60192 | !hbusreq1_p & !a5f8ce;
assign dead8a = hlock1_p & b26695 | !hlock1_p & !dead89;
assign c3bd63 = hlock2_p & c3bd62 | !hlock2_p & !c3bc3c;
assign a5f398 = hbusreq2 & a5f396 | !hbusreq2 & a5f397;
assign hgrant2 = !b29b61;
assign cea1a2 = hmaster1_p & cea1a0 | !hmaster1_p & cea1a1;
assign a81ce5 = hmaster1_p & v84563c | !hmaster1_p & a81ce4;
assign a5fd22 = hbusreq2 & a5fd21 | !hbusreq2 & ab0c32;
assign b29a92 = hbusreq2_p & b29a8e | !hbusreq2_p & v84563c;
assign cea0b8 = hlock0_p & cea0b7 | !hlock0_p & v84563c;
assign a5f903 = hlock2_p & a5f902 | !hlock2_p & v84563c;
assign a5fa6b = hlock0_p & v845641 | !hlock0_p & v84563c;
assign a5efb7 = locked_p & v84563c | !locked_p & a5efae;
assign a5ea53 = locked_p & a5ea52 | !locked_p & v845641;
assign dea746 = hbusreq2_p & deadc6 | !hbusreq2_p & deadc5;
assign c3b703 = hgrant2_p & dead3e | !hgrant2_p & cea18d;
assign deadd0 = hlock1_p & deac52 | !hlock1_p & !deadcf;
assign ab0b62 = hbusreq3 & ab0b5d | !hbusreq3 & ab0b61;
assign b29946 = hlock1_p & v84565a | !hlock1_p & !b8acdb;
assign a5ea37 = hbusreq2_p & a5f08a | !hbusreq2_p & a5fb6c;
assign ab0b5e = locked_p & v84563c | !locked_p & !b29832;
assign a5ee21 = hbusreq1 & a5ee1f | !hbusreq1 & !a5ee20;
assign b29e4a = hgrant2_p & dead3e | !hgrant2_p & !b29e49;
assign cea3f2 = hgrant2_p & cea3ee | !hgrant2_p & cea3f1;
assign a5fcf0 = hbusreq2 & a5fcc8 | !hbusreq2 & a5fcef;
assign c3bcde = hlock2_p & c3bcdd | !hlock2_p & !dead77;
assign a5f8ff = hlock1_p & v84566c | !hlock1_p & a5f8fe;
assign cea323 = hlock1_p & deae02 | !hlock1_p & v84566c;
assign a5ea9e = hbusreq2_p & a5ea9a | !hbusreq2_p & !a5ea9d;
assign adaee9 = start_p & v84563c | !start_p & d5edb8;
assign ab0cd0 = hready_p & ab0cbc | !hready_p & !ab0ccf;
assign a81cd4 = hlock2_p & a81caa | !hlock2_p & v84563c;
assign b29fdf = hlock2 & b29fdc | !hlock2 & b29fde;
assign a5f238 = hlock2 & a5fa8a | !hlock2 & a5f237;
assign b26777 = hlock2_p & b266af | !hlock2_p & b266a0;
assign a5f206 = hgrant0_p & a5f1ec | !hgrant0_p & a5f205;
assign a5f218 = hmaster1_p & v84563c | !hmaster1_p & a5f217;
assign c3bcab = hgrant2_p & c3bcaa | !hgrant2_p & !v845660;
assign ab053b = hgrant1_p & ab053a | !hgrant1_p & v84563c;
assign af3583 = hlock2_p & af352d | !hlock2_p & v84563c;
assign a5fa63 = hgrant1_p & v9703fb | !hgrant1_p & a5fa13;
assign af3c68 = hmaster0_p & af3c5c | !hmaster0_p & af3c67;
assign c3b7a7 = hbusreq2_p & c3b7a5 | !hbusreq2_p & c3b7a6;
assign dead71 = locked_p & dead70 | !locked_p & !v84563c;
assign a5f6f2 = hready & v84563c | !hready & a5f6e6;
assign v845648 = hlock1_p & v84563c | !hlock1_p & !v84563c;
assign start = !a9b9f0;
assign cea431 = hlock2_p & cea430 | !hlock2_p & cea3fb;
assign ab066a = hbusreq0_p & dead34 | !hbusreq0_p & b29eac;
assign deac79 = hbusreq3 & deac78 | !hbusreq3 & v84563c;
assign b29b18 = hmaster1_p & b29a9a | !hmaster1_p & b29e6e;
assign a5f331 = hbusreq2_p & a5f8f0 | !hbusreq2_p & !v84563c;
assign a5f9da = hburst0_p & v845672 | !hburst0_p & a5f9d9;
assign a5fbf0 = hready & a5fbec | !hready & a5fbef;
assign b266a9 = hlock0_p & b2669d | !hlock0_p & b266a8;
assign ce9d20 = hbusreq2_p & cea276 | !hbusreq2_p & cea275;
assign c3b816 = hgrant2_p & c3b813 | !hgrant2_p & c3b815;
assign ab0b22 = hbusreq0_p & b29cf2 | !hbusreq0_p & v84565a;
assign v970439 = hgrant2_p & v970438 | !hgrant2_p & v84563c;
assign a5e9ba = hlock1_p & a5fb8b | !hlock1_p & a5e9b9;
assign c3bc9c = hgrant2_p & c3bc97 | !hgrant2_p & c3bc9b;
assign a5f73b = hbusreq2 & a5f71d | !hbusreq2 & a5f73a;
assign a5f97a = hlock2_p & a5f977 | !hlock2_p & a5f979;
assign b840ae = hmaster0_p & b840ac | !hmaster0_p & b840ad;
assign a5ef91 = hbusreq3 & a5ef0b | !hbusreq3 & a5ef13;
assign c3b76e = hmaster0_p & c3b76d | !hmaster0_p & c3b6b6;
assign cea370 = hready_p & cea364 | !hready_p & cea36f;
assign bdb58b = hlock0_p & cea0bc | !hlock0_p & !v84565a;
assign ab0cfd = hmaster0_p & ab0cf9 | !hmaster0_p & ab0cfc;
assign a5f58d = hlock0_p & a5f58c | !hlock0_p & a5f4ee;
assign b29ac3 = hmaster1_p & b29ac2 | !hmaster1_p & b29e48;
assign c3bda1 = hbusreq2_p & c3bcf3 | !hbusreq2_p & c3bc6e;
assign cea17c = hgrant2_p & v84563c | !hgrant2_p & cea17b;
assign cea293 = hgrant1_p & deaca1 | !hgrant1_p & cea255;
assign c3b7a0 = hlock0_p & c3bce6 | !hlock0_p & v845660;
assign a5f393 = hbusreq3 & a5f392 | !hbusreq3 & a5fbc0;
assign b29d49 = hbusreq3 & v84563c | !hbusreq3 & b29d1e;
assign af3540 = hgrant1_p & af353f | !hgrant1_p & af352c;
assign b29975 = hmaster0_p & b29962 | !hmaster0_p & b29974;
assign ab0b09 = hlock0_p & v84563c | !hlock0_p & !deadde;
assign af3569 = hmaster1_p & v84563c | !hmaster1_p & af354c;
assign af356e = hlock3_p & af3568 | !hlock3_p & af356d;
assign a5fca2 = hbusreq1_p & v84563c | !hbusreq1_p & !b2982c;
assign d40d36 = hlock1_p & d40d31 | !hlock1_p & d40d35;
assign b29ab6 = hgrant2_p & b29ab5 | !hgrant2_p & !b29d5a;
assign ab068f = hlock2_p & ab068d | !hlock2_p & ab068e;
assign a5f1b4 = hlock2 & a5fc56 | !hlock2 & a5f1b3;
assign a5f43e = hlock1_p & v84565a | !hlock1_p & deac18;
assign c3b84f = hbusreq2_p & c3b84b | !hbusreq2_p & c3b849;
assign ab0cc7 = hbusreq2_p & ab0cc6 | !hbusreq2_p & v84563c;
assign b29fd1 = hlock0_p & b29f51 | !hlock0_p & c3bd5f;
assign a5f7c3 = hlock0_p & a5f7c0 | !hlock0_p & a5f7c2;
assign a5edf7 = hready & a5edf6 | !hready & v84563c;
assign ab06ee = hmaster1_p & ab06ed | !hmaster1_p & ab0b71;
assign a5ef9d = hbusreq0_p & a5f3a1 | !hbusreq0_p & a5f390;
assign adaed8 = hmaster1_p & adaed7 | !hmaster1_p & v84563c;
assign b29a63 = hgrant1_p & b29a62 | !hgrant1_p & c3b683;
assign a5ef43 = hmaster1_p & a5ef42 | !hmaster1_p & v84563c;
assign b266a2 = hlock1_p & b26695 | !hlock1_p & b266a1;
assign a5f37d = hbusreq1 & a5f377 | !hbusreq1 & v84563c;
assign ab06c4 = hmaster1_p & ab06c3 | !hmaster1_p & !ab0640;
assign b29abe = hlock0_p & b29abd | !hlock0_p & !dead77;
assign b2677f = hmaster1_p & b266ae | !hmaster1_p & b266a3;
assign a5fb72 = hbusreq1_p & v84563c | !hbusreq1_p & a5fb71;
assign cea4ab = hbusreq3 & cea4aa | !hbusreq3 & cea425;
assign af34c0 = hmaster1_p & af34b2 | !hmaster1_p & af34bf;
assign c3b8ca = jx1_p & c3b8b8 | !jx1_p & c3b77f;
assign a5f124 = hbusreq2_p & a5f123 | !hbusreq2_p & !a5f122;
assign a5ee00 = hlock0_p & a5edf5 | !hlock0_p & a5edff;
assign c3b7b1 = hlock0_p & c3bcef | !hlock0_p & !v84563c;
assign a5ea8e = hlock3_p & a5ea6f | !hlock3_p & a5ea8d;
assign a5f984 = locked_p & a5f983 | !locked_p & v84563c;
assign a60188 = hlock1_p & a60187 | !hlock1_p & v84563c;
assign cea35f = hbusreq2_p & cea2f3 | !hbusreq2_p & cea18f;
assign ab05fb = hbusreq2_p & ab057f | !hbusreq2_p & ab05fa;
assign d40d76 = hgrant0_p & d40d6c | !hgrant0_p & d40d75;
assign v85f3c3 = stateG3_0_p & v84563c | !stateG3_0_p & v845674;
assign a5f4a8 = hready & a5f4a6 | !hready & a5f4a7;
assign c3b6c3 = hgrant1_p & c3b6a4 | !hgrant1_p & c3b691;
assign a5eada = hbusreq0_p & v84563c | !hbusreq0_p & a5f8ca;
assign cea330 = hgrant1_p & cea26b | !hgrant1_p & cea26d;
assign a5f02b = hlock3_p & a5f023 | !hlock3_p & a5f02a;
assign a5e9e1 = hbusreq2_p & a5e9e0 | !hbusreq2_p & a5f14c;
assign cea363 = hgrant0_p & cea35a | !hgrant0_p & cea362;
assign a5ef28 = hbusreq2 & a5edec | !hbusreq2 & !a5edf2;
assign b26787 = hbusreq2_p & b26785 | !hbusreq2_p & b266f0;
assign af348e = hlock0_p & af3c49 | !hlock0_p & d40d33;
assign b29e5e = hmaster0_p & b29e5d | !hmaster0_p & b29e5c;
assign ab0b6a = hlock2_p & ab0b5f | !hlock2_p & v845660;
assign a5f94b = hbusreq0 & a5f93d | !hbusreq0 & a5f94a;
assign a5e9d3 = hbusreq0 & a5e9d2 | !hbusreq0 & v845641;
assign a81cc2 = hlock0_p & a81cb1 | !hlock0_p & v84563c;
assign ab0b89 = locked_p & dead6e | !locked_p & b29d82;
assign a5ee28 = hbusreq0_p & a5ee24 | !hbusreq0_p & a5ee27;
assign a5eee9 = hready & a5eee8 | !hready & a5f45a;
assign a5efea = hbusreq0 & a5efe7 | !hbusreq0 & !a5efe9;
assign b29918 = stateG10_1_p & v84563c | !stateG10_1_p & deacbc;
assign b29d92 = hlock0_p & b26695 | !hlock0_p & !v84563c;
assign a5f24b = hbusreq2 & a5f24a | !hbusreq2 & !ab0c31;
assign a5ef5f = hlock0_p & a5f4fc | !hlock0_p & a5ef5e;
assign ab0730 = hready_p & ab0704 | !hready_p & !ab072f;
assign c3bddd = hgrant2_p & c3bdda | !hgrant2_p & c3bddc;
assign c3bcb2 = hgrant3_p & c3bc46 | !hgrant3_p & c3bcb1;
assign bdb5b2 = hbusreq2_p & bdb5b1 | !hbusreq2_p & !v84565a;
assign deae86 = hlock0_p & deae81 | !hlock0_p & !deadc4;
assign b29f7a = hlock0_p & b29f79 | !hlock0_p & c3bd61;
assign b266e7 = hlock2_p & b266d2 | !hlock2_p & b26695;
assign c3b7fa = hlock0_p & c3bd7a | !hlock0_p & deada8;
assign b26695 = hmastlock_p & b26694 | !hmastlock_p & v84566c;
assign a5f500 = hlock2 & a5f4fc | !hlock2 & a5f36e;
assign ab0bd6 = hlock2_p & ab0b38 | !hlock2_p & ab0bd5;
assign a5fc5c = locked_p & a5fc04 | !locked_p & v84563c;
assign ab0ce9 = hmaster1_p & ab0ce8 | !hmaster1_p & ab0c87;
assign c3b6a6 = hlock1_p & v84563c | !hlock1_p & !c3b6a5;
assign deacef = hbusreq2_p & deacea | !hbusreq2_p & deacee;
assign af3c3d = hlock3_p & af3c3c | !hlock3_p & af3c27;
assign a5f201 = hlock2_p & a5f200 | !hlock2_p & v84563c;
assign ce9d3e = hgrant2_p & cea25b | !hgrant2_p & ce9d3d;
assign b29e9c = hmaster1_p & b29e9b | !hmaster1_p & b29e65;
assign b29d74 = hgrant2_p & b29d6b | !hgrant2_p & !b29d73;
assign bdb5ae = decide_p & bdb581 | !decide_p & v845660;
assign b29a5d = hbusreq2_p & b29a5c | !hbusreq2_p & !b29a5b;
assign b2990a = hlock0_p & b29832 | !hlock0_p & v84563c;
assign b29fe8 = hlock3_p & b29fe7 | !hlock3_p & b29f82;
assign b29cf8 = hlock2_p & b29cf7 | !hlock2_p & v84563c;
assign ab0b03 = hbusreq2_p & ab0b02 | !hbusreq2_p & v84563c;
assign a5f344 = hbusreq2_p & a5f343 | !hbusreq2_p & v84563c;
assign v845672 = stateG3_1_p & v84563c | !stateG3_1_p & !v84563c;
assign a5f120 = hready & a5f11f | !hready & a5f83b;
assign ab069c = hbusreq3 & ab0690 | !hbusreq3 & ab069b;
assign dea700 = hbusreq3_p & dea6ff | !hbusreq3_p & dead6a;
assign b29edd = hbusreq3 & b29edc | !hbusreq3 & !v84564a;
assign a5eaa0 = hgrant2_p & a5ea9f | !hgrant2_p & a5f0ae;
assign a5fc1b = hlock2 & a5fb91 | !hlock2 & a5fc1a;
assign a5f32d = hbusreq3 & a5f32a | !hbusreq3 & a5f32c;
assign c3b754 = hmaster1_p & c3b753 | !hmaster1_p & c3bcc0;
assign a5f74a = hlock3_p & a5f731 | !hlock3_p & a5f749;
assign ab0c6e = hbusreq2_p & ab0c6d | !hbusreq2_p & v84563c;
assign b29ea3 = hgrant3_p & b29e72 | !hgrant3_p & b29ea2;
assign c3b779 = hmaster0_p & c3b778 | !hmaster0_p & c3bca4;
assign af3c50 = locked_p & af3c49 | !locked_p & af3c4c;
assign b266fa = hlock0_p & b266cd | !hlock0_p & b266bb;
assign a81cf6 = hbusreq1_p & a81cb1 | !hbusreq1_p & a81cf0;
assign c3bde9 = hmaster0_p & c3bde7 | !hmaster0_p & c3bde8;
assign a5fba3 = stateA1_p & a81ca6 | !stateA1_p & !v845654;
assign a81cd2 = hgrant2_p & v84563c | !hgrant2_p & a81cd1;
assign a60167 = start_p & v84563c | !start_p & a60166;
assign adaf02 = hlock0_p & adaed7 | !hlock0_p & adaf01;
assign a5f46f = hbusreq1 & a5f46e | !hbusreq1 & v84563c;
assign a5f024 = hbusreq2_p & a5fd36 | !hbusreq2_p & a5fad6;
assign c3bd80 = hlock3_p & c3bd68 | !hlock3_p & !c3bd7f;
assign deac0f = hbusreq3 & v845660 | !hbusreq3 & v84563c;
assign deace5 = hlock2_p & deace2 | !hlock2_p & deace4;
assign dea751 = hbusreq2_p & deade1 | !hbusreq2_p & deade0;
assign cea477 = decide_p & cea476 | !decide_p & a57859;
assign adaf04 = hmaster0_p & v84563c | !hmaster0_p & adaf03;
assign c3bcc9 = hbusreq2_p & c3bcc8 | !hbusreq2_p & !v84563c;
assign deae5c = hlock0_p & deae5b | !hlock0_p & !v84563c;
assign deae3c = hmaster1_p & dead54 | !hmaster1_p & deae3b;
assign bdb5a5 = hgrant2_p & bdb598 | !hgrant2_p & !v84565a;
assign cea86e = hbusreq2_p & cea86d | !hbusreq2_p & v84563c;
assign a60198 = hready & a60195 | !hready & a60197;
assign ab05f3 = hbusreq3 & ab05ef | !hbusreq3 & ab05f2;
assign c3b6ea = hgrant2_p & c3b6e9 | !hgrant2_p & c3bc70;
assign c3bcad = hmaster0_p & c3bca7 | !hmaster0_p & !c3bcac;
assign ab0ae3 = hbusreq3 & ab0ad6 | !hbusreq3 & ab0ae2;
assign a5ea68 = hbusreq0 & a5ea63 | !hbusreq0 & a5ea67;
assign b29ec1 = hlock2 & b29ebf | !hlock2 & b29ec0;
assign ce9e20 = hgrant2_p & cea368 | !hgrant2_p & ce9e1f;
assign a5fceb = hmaster0_p & a5fcca | !hmaster0_p & a5fcea;
assign ce9d5b = decide_p & ce9d5a | !decide_p & a57859;
assign adaed7 = locked_p & adaec4 | !locked_p & v84563c;
assign ce9cb9 = hbusreq2_p & ce9cb8 | !hbusreq2_p & !cea38d;
assign stateG10_1 = !c98ba4;
assign a5eaed = hbusreq3 & a5eadf | !hbusreq3 & !a5eaec;
assign c3bc5e = hbusreq2_p & c3bc5d | !hbusreq2_p & c3bc5c;
assign a5ea61 = hlock0_p & a5fc1a | !hlock0_p & v84563c;
assign b2676f = hmaster1_p & b266a0 | !hmaster1_p & !b266e0;
assign a5ef7b = hlock0_p & a5edcc | !hlock0_p & a5ef5e;
assign cea365 = hready & cea0bc | !hready & !c98b95;
assign a5fcd7 = hmastlock_p & a5fcd6 | !hmastlock_p & v84563c;
assign ab0719 = hbusreq3 & ab0714 | !hbusreq3 & ab0718;
assign ab0cf6 = decide_p & ab0cf5 | !decide_p & v845662;
assign b2673b = hlock0_p & b26720 | !hlock0_p & b266b1;
assign a5eb96 = hbusreq2_p & a5eb95 | !hbusreq2_p & a5ea69;
assign a5fa42 = hlock2 & a5fa2e | !hlock2 & a5fa41;
assign c3bc93 = hbusreq2_p & c3bc92 | !hbusreq2_p & !dead21;
assign a81cb5 = hlock1_p & a81cb1 | !hlock1_p & v84563c;
assign ab0be8 = hgrant0_p & ab0be1 | !hgrant0_p & !ab0be7;
assign ab0b94 = hbusreq3 & ab0b93 | !hbusreq3 & ab0b70;
assign ab0cb1 = hbusreq2_p & ab0cb0 | !hbusreq2_p & v845660;
assign a5fcb6 = hgrant2_p & a5fcb5 | !hgrant2_p & a5fc73;
assign deae30 = hlock1_p & deacdf | !hlock1_p & dead92;
assign ab061f = hlock2 & ab052f | !hlock2 & ab061e;
assign ab05a9 = hlock2_p & ab05a6 | !hlock2_p & ab05a8;
assign c3b6da = hmaster1_p & c3b6d9 | !hmaster1_p & c3bc5e;
assign c3bca0 = hlock0_p & dead77 | !hlock0_p & v84563c;
assign a5ea10 = hbusreq0 & a5ea00 | !hbusreq0 & a5ea0f;
assign a5ede8 = hready & a5ede7 | !hready & v84563c;
assign a5fc01 = hlock1_p & a5fb8b | !hlock1_p & a5fc00;
assign ce9d22 = hgrant2_p & cea278 | !hgrant2_p & ce9d21;
assign dea76d = hgrant0_p & dead2d | !hgrant0_p & dea76c;
assign a5f93a = hlock0_p & a5f939 | !hlock0_p & a5f8c5;
assign a5ee07 = hlock0_p & a5f387 | !hlock0_p & a5f36b;
assign a5ef3c = hbusreq2_p & a5ef39 | !hbusreq2_p & a5ef3b;
assign a5fb7a = locked_p & v84563c | !locked_p & a5fb79;
assign ab060e = hlock2 & ab0529 | !hlock2 & ab060d;
assign a5f959 = hmaster1_p & a5f956 | !hmaster1_p & a5f958;
assign c3b618 = hbusreq2_p & c3b615 | !hbusreq2_p & c3bc0d;
assign a5fcce = locked_p & v845641 | !locked_p & v84565a;
assign af3c4c = hmastlock_p & af3c4b | !hmastlock_p & v84563c;
assign b299f2 = hmaster0_p & b299f0 | !hmaster0_p & !b299f1;
assign a81cda = start_p & a81ca6 | !start_p & c07311;
assign deace9 = locked_p & v84563c | !locked_p & b26695;
assign cea470 = hlock2_p & cea395 | !hlock2_p & cea3aa;
assign c3bc80 = hlock2_p & c3bc7f | !hlock2_p & cea18d;
assign v970449 = hbusreq2_p & v9703fd | !hbusreq2_p & v97043f;
assign c3b679 = stateG10_1_p & deacb4 | !stateG10_1_p & c3b678;
assign a5f26e = hbusreq2_p & a5f26d | !hbusreq2_p & !v84563c;
assign ab0cbf = hlock2 & ab0b09 | !hlock2 & ab0cbe;
assign b29e9e = hgrant2_p & b29e9d | !hgrant2_p & b29d05;
assign a5ea84 = hbusreq2 & a5ea80 | !hbusreq2 & !a5ea83;
assign a5f035 = decide_p & a5f034 | !decide_p & v84563c;
assign ab062b = hlock0_p & ab0adc | !hlock0_p & !ab05ed;
assign af3c33 = hmaster0_p & af3c32 | !hmaster0_p & af3c31;
assign a5f922 = hready & v84563c | !hready & a5f921;
assign c3bbf6 = stateG10_1_p & cea8a7 | !stateG10_1_p & c3bbd2;
assign deadec = hgrant1_p & v84563c | !hgrant1_p & deadeb;
assign a5f216 = hmaster1_p & a5f212 | !hmaster1_p & a5f215;
assign a5fb4c = hready & a60192 | !hready & v9703fb;
assign a5ee8d = locked_p & a5ee8c | !locked_p & !v845641;
assign a9b9d5 = hready_p & a9b9d4 | !hready_p & v84563c;
assign a5f2d9 = hbusreq2 & a5fce5 | !hbusreq2 & !v84563c;
assign c3bd04 = hbusreq2_p & c3bd03 | !hbusreq2_p & v84563c;
assign b29cd7 = hbusreq2_p & b29cca | !hbusreq2_p & v84563c;
assign c3bcf1 = hbusreq0_p & c3bcee | !hbusreq0_p & c3bcf0;
assign c3b63d = hbusreq2_p & c3b63c | !hbusreq2_p & c3b63b;
assign dead0c = hlock1_p & b26695 | !hlock1_p & dead09;
assign ab0576 = hgrant2_p & ab0574 | !hgrant2_p & ab0575;
assign b29fce = hgrant0_p & b29fbc | !hgrant0_p & !b29fcd;
assign deacc1 = hbusreq2_p & deaca1 | !hbusreq2_p & v84563c;
assign a60197 = hbusreq1 & v84563c | !hbusreq1 & a60196;
assign c3b884 = hbusreq2_p & c3b7dc | !hbusreq2_p & c3b883;
assign a5f6d8 = hgrant2_p & a5f6d4 | !hgrant2_p & a5f6d7;
assign c3b7ef = hbusreq3 & c3b7e4 | !hbusreq3 & c3b7e6;
assign a5ebc8 = hbusreq0 & a5ebc7 | !hbusreq0 & v845641;
assign a5eb75 = hgrant2_p & a5eb70 | !hgrant2_p & a5eb74;
assign a5f805 = hlock1_p & a5f7f5 | !hlock1_p & a5f804;
assign af357c = hmaster1_p & af3531 | !hmaster1_p & af357b;
assign b29ce8 = hready & deac52 | !hready & v84565a;
assign a5f11a = start_p & v845654 | !start_p & a5f7f3;
assign d40d2e = hmaster0_p & d40d2d | !hmaster0_p & v84563c;
assign deae0a = hmaster0_p & deae00 | !hmaster0_p & deae09;
assign a5f885 = hbusreq2_p & a5f884 | !hbusreq2_p & v84563c;
assign b29ff2 = decide_p & b29ff1 | !decide_p & v84563c;
assign b29eba = hready & b29eb9 | !hready & v84563c;
assign b2672b = hlock1_p & b26695 | !hlock1_p & b266da;
assign dea6eb = hmaster1_p & dea6ea | !hmaster1_p & !dead5f;
assign a81cd9 = hgrant0_p & a81ccf | !hgrant0_p & a81cd8;
assign cea15b = hlock2_p & cea15a | !hlock2_p & v845660;
assign a5eea6 = locked_p & a5eea5 | !locked_p & !v845641;
assign d40d9a = decide_p & d40d99 | !decide_p & d40d8a;
assign a5ee3b = hlock2 & a5ee37 | !hlock2 & a5ee3a;
assign ab0aed = hgrant1_p & ab0aec | !hgrant1_p & ab0aeb;
assign cea2f8 = hmaster0_p & cea2f6 | !hmaster0_p & cea2f7;
assign c3bd46 = hgrant2_p & c3bd43 | !hgrant2_p & c3bd45;
assign b29f67 = hbusreq3 & b29f65 | !hbusreq3 & b29f66;
assign a5fce4 = hready & a5fce1 | !hready & a5fce3;
assign a5fbba = hlock2_p & a5fbb4 | !hlock2_p & !a5fbb9;
assign a5fcc6 = hlock1_p & v84563c | !hlock1_p & deacbc;
assign a5ec21 = decide_p & a5ec20 | !decide_p & v84563c;
assign c3bc5b = hbusreq2_p & c3bc59 | !hbusreq2_p & c3bc5a;
assign ab0bfc = hlock0_p & v84563c | !hlock0_p & !ab0bfb;
assign a5eec7 = hbusreq0 & a5eebe | !hbusreq0 & !a5eec6;
assign deae45 = hgrant2_p & deadf0 | !hgrant2_p & deae44;
assign b299b0 = hmaster1_p & b299af | !hmaster1_p & b29e5c;
assign cea35a = hmaster0_p & cea359 | !hmaster0_p & cea2ed;
assign ce9d53 = hlock2_p & ce9d52 | !hlock2_p & !ce9d47;
assign c3b73e = decide_p & c3b73d | !decide_p & !v845660;
assign a5edde = hbusreq0 & a5edd7 | !hbusreq0 & a5eddd;
assign ab050b = hlock0_p & v84563c | !hlock0_p & !b29833;
assign b29a4f = hbusreq2_p & b29a4e | !hbusreq2_p & v84563c;
assign b26765 = hgrant0_p & b2675b | !hgrant0_p & b26764;
assign af3c1c = hlock0_p & v8c6711 | !hlock0_p & v845646;
assign b29f07 = stateA1_p & v8c6449 | !stateA1_p & cea24b;
assign c3b822 = hgrant2_p & c3b81e | !hgrant2_p & c3b821;
assign b2a010 = hlock2_p & b2a00f | !hlock2_p & v84563c;
assign cea2ae = hready & cea2ac | !hready & cea2ad;
assign b2995d = hbusreq3 & b2995a | !hbusreq3 & b2995c;
assign b266b6 = hmaster1_p & b266b0 | !hmaster1_p & b266b5;
assign dea6ff = hgrant3_p & dea6f9 | !hgrant3_p & !dea6fe;
assign dead2d = hbusreq2_p & dead2c | !hbusreq2_p & v845660;
assign dea72c = hmaster0_p & dea729 | !hmaster0_p & dea72b;
assign b29f65 = hbusreq2_p & b29f60 | !hbusreq2_p & v84563c;
assign af3c7a = hgrant1_p & af3c79 | !hgrant1_p & af3c49;
assign c3b61b = hmaster1_p & c3b61a | !hmaster1_p & c3bd50;
assign af35a0 = decide_p & af3596 | !decide_p & af359f;
assign c3b60b = decide_p & c3b60a | !decide_p & v845660;
assign a5f0e5 = hbusreq0_p & v84563c | !hbusreq0_p & a5f7cb;
assign ab0587 = hready_p & ab0534 | !hready_p & ab0586;
assign cea275 = hlock0_p & cea274 | !hlock0_p & v84563c;
assign adaebd = locked_p & adaebc | !locked_p & v84563c;
assign deac51 = hmastlock_p & deac50 | !hmastlock_p & !v84563c;
assign a5fd34 = hbusreq0_p & a5fd23 | !hbusreq0_p & v84563c;
assign af3c6f = hmaster1_p & af3c50 | !hmaster1_p & af3c58;
assign a5fb37 = hgrant2_p & a5fb2f | !hgrant2_p & a5fb36;
assign a5ee97 = hlock2_p & a5ee96 | !hlock2_p & a5ee3e;
assign af3c34 = hgrant0_p & af3c16 | !hgrant0_p & af3c33;
assign a5f365 = hbusreq1 & a5f364 | !hbusreq1 & v84563c;
assign a5f7f3 = stateA1_p & d40d29 | !stateA1_p & !c06d34;
assign cea198 = hlock2_p & cea197 | !hlock2_p & !v84563c;
assign c3b665 = hready & c3b664 | !hready & c3bd16;
assign b266d2 = hlock0_p & b266cd | !hlock0_p & b266ca;
assign ab0530 = hbusreq3 & ab052f | !hbusreq3 & ab052d;
assign b298a8 = hbusreq3 & b298a3 | !hbusreq3 & b298a7;
assign a5ee64 = hlock2_p & a5ee61 | !hlock2_p & a5ee63;
assign cea45b = hgrant2_p & cea45a | !hgrant2_p & !cea15c;
assign ab06e3 = hbusreq2_p & ab06e2 | !hbusreq2_p & ab06e0;
assign b29d2b = hgrant2_p & b29d29 | !hgrant2_p & b29d2a;
assign cea167 = hmaster1_p & cea15d | !hmaster1_p & cea166;
assign a5f14a = hready & a60195 | !hready & a5f149;
assign b29ac5 = hgrant0_p & c3bceb | !hgrant0_p & !b29ac4;
assign ab0523 = hlock0_p & v84563c | !hlock0_p & !b298ae;
assign a5ee92 = hmaster1_p & a5ee85 | !hmaster1_p & a5ee91;
assign deadff = hbusreq2_p & deadfe | !hbusreq2_p & v845660;
assign deacfe = hlock0_p & deace9 | !hlock0_p & deacfc;
assign ab0680 = hbusreq3 & ab067f | !hbusreq3 & dead2e;
assign a5f176 = hlock1_p & a5fb8b | !hlock1_p & a5f175;
assign dead31 = stateG2_p & v84563c | !stateG2_p & !c07311;
assign a5edeb = hready & a5edea | !hready & v84563c;
assign b29823 = hbusreq1_p & b2a020 | !hbusreq1_p & dead33;
assign a5ea67 = hbusreq2_p & a5ea66 | !hbusreq2_p & a5ea3c;
assign cea0d7 = hmaster0_p & cea8a4 | !hmaster0_p & cea0d6;
assign ab0c34 = hlock2_p & ab0c30 | !hlock2_p & ab0c33;
assign c3b6e2 = hlock0_p & c3b6df | !hlock0_p & !c3b6e1;
assign a5fb86 = hburst1_p & d5edb8 | !hburst1_p & v84563c;
assign b8acd7 = jx0_p & v8565cf | !jx0_p & !v84563c;
assign a5fc26 = hgrant2_p & a5fc20 | !hgrant2_p & a5fc25;
assign a5f82c = hready & a5f82b | !hready & a5fa1d;
assign a5eb8c = locked_p & v84563c | !locked_p & a5eb8b;
assign c98b9e = decide_p & c98b96 | !decide_p & v8c6711;
assign ce9d6f = hbusreq2_p & cea336 | !hbusreq2_p & cea335;
assign b29927 = hbusreq1_p & v84563c | !hbusreq1_p & !deadb9;
assign a5efb9 = hlock0_p & a5ee66 | !hlock0_p & a5efb8;
assign a5f39e = hready & v84563c | !hready & c3b624;
assign b26731 = hmaster1_p & b26724 | !hmaster1_p & b26730;
assign adaec6 = hmastlock_p & adaec5 | !hmastlock_p & v84563c;
assign cea1be = hready & cea1bd | !hready & dead7d;
assign a5f755 = hmaster1_p & v84563c | !hmaster1_p & a5f754;
assign a5ea2c = hbusreq0 & a5ea2b | !hbusreq0 & v84563c;
assign deac5f = hbusreq2_p & deac5d | !hbusreq2_p & deac5b;
assign dea6f1 = hmaster1_p & deac3f | !hmaster1_p & !v84563c;
assign a5f594 = hbusreq2_p & a5f593 | !hbusreq2_p & a5f592;
assign b299ed = hgrant2_p & b29d1e | !hgrant2_p & b29d21;
assign a5785a = hready_p & a57859 | !hready_p & !v845656;
assign a5f487 = hgrant1_p & a5f486 | !hgrant1_p & a5f9dd;
assign c3bd3d = hlock1_p & deadb9 | !hlock1_p & c3bd3c;
assign a5eeae = hbusreq2 & a5eead | !hbusreq2 & a5ee71;
assign c3bca5 = hbusreq3 & cea17a | !hbusreq3 & !cea18d;
assign a5f2f8 = hlock2_p & a5f2f7 | !hlock2_p & v84563c;
assign a5f193 = hlock0_p & a5f18d | !hlock0_p & !a5f192;
assign b266bb = hbusreq0_p & b26695 | !hbusreq0_p & !b266a0;
assign af35c4 = jx0_p & af3511 | !jx0_p & !af35c3;
assign cea27a = hbusreq3 & cea279 | !hbusreq3 & cea277;
assign v97043c = hgrant0_p & v970433 | !hgrant0_p & v97043b;
assign a5ee50 = hlock0_p & a5ee4d | !hlock0_p & a5ee4f;
assign b29fb0 = hbusreq2_p & b29faf | !hbusreq2_p & v84563c;
assign a5eb42 = hbusreq0 & a5eb41 | !hbusreq0 & v84563c;
assign cea398 = hbusreq3 & cea397 | !hbusreq3 & cea391;
assign a5f323 = hlock0_p & a5fa6c | !hlock0_p & ab0c31;
assign a5f574 = hbusreq1 & a5f571 | !hbusreq1 & !a5f573;
assign a5f075 = hbusreq0 & a5f06e | !hbusreq0 & a5f074;
assign b29835 = hlock2_p & v84563c | !hlock2_p & !b29834;
assign a5f92f = hlock0_p & a5f92e | !hlock0_p & a5f8ba;
assign c3bd13 = hbusreq1_p & c3bd11 | !hbusreq1_p & !v84563c;
assign ab0c9f = hbusreq2_p & ab0c9e | !hbusreq2_p & cea15a;
assign c3bd6a = hbusreq2_p & c3bd69 | !hbusreq2_p & v84563c;
assign b29996 = hbusreq2_p & b2998f | !hbusreq2_p & b29995;
assign c3b8ac = hbusreq2_p & c3b8ab | !hbusreq2_p & !c3b7e6;
assign b29831 = hready & b2982e | !hready & b29830;
assign a5f54b = hlock0_p & a5fa6c | !hlock0_p & a5f4f0;
assign v84564d = hlock2 & v84563c | !hlock2 & !v84563c;
assign a5fd10 = hlock0_p & a5fccb | !hlock0_p & a5fd0f;
assign a5f723 = hbusreq3 & a5f722 | !hbusreq3 & v84563c;
assign a5f3d3 = hbusreq1_p & b266a0 | !hbusreq1_p & !v84563c;
assign b29ee7 = hburst0 & b29ee5 | !hburst0 & b29ee6;
assign cea24b = hburst0_p & v84563c | !hburst0_p & cea24a;
assign a5ea35 = hbusreq2_p & a5ea33 | !hbusreq2_p & a5ea34;
assign a81cb2 = stateG10_1_p & v84563c | !stateG10_1_p & a81cb1;
assign ce9cc6 = hbusreq2_p & ce9cc1 | !hbusreq2_p & ce9cc0;
assign a5f3a3 = locked_p & a60140 | !locked_p & a5f36e;
assign b29d4a = hbusreq3 & v84563c | !hbusreq3 & b29d21;
assign cea14a = hbusreq2_p & cea149 | !hbusreq2_p & cea148;
assign deae98 = hbusreq3 & deae93 | !hbusreq3 & deae97;
assign ab068d = hlock0_p & b29eed | !hlock0_p & !ab068c;
assign a5ee33 = hbusreq2_p & a5ee32 | !hbusreq2_p & a5ee29;
assign a5faab = hgrant1_p & a60193 | !hgrant1_p & a5faaa;
assign a5fafb = hlock1_p & a60186 | !hlock1_p & v84563c;
assign a5f532 = stateG10_1_p & v9703fb | !stateG10_1_p & a5f4e5;
assign a5fc77 = start_p & deac4a | !start_p & a5fc76;
assign a5f6fd = hbusreq2_p & a5f6fc | !hbusreq2_p & a60142;
assign a5fb68 = decide_p & a5fb67 | !decide_p & v84563c;
assign ce9e27 = hready_p & ce9e0c | !hready_p & ce9e26;
assign a5ea5e = hbusreq2 & a5f089 | !hbusreq2 & a5fa6b;
assign cea172 = hbusreq2_p & cea16b | !hbusreq2_p & cea16a;
assign a5eafc = hmaster0_p & a5eaf5 | !hmaster0_p & a5e9cf;
assign dead44 = hmaster1_p & dead3c | !hmaster1_p & dead43;
assign ab0b65 = hbusreq0_p & deace9 | !hbusreq0_p & b29d88;
assign a5f473 = hlock0_p & a5f472 | !hlock0_p & a5f45b;
assign a5eef0 = hbusreq2 & a5eee9 | !hbusreq2 & a5eeef;
assign cea283 = hlock0_p & cea280 | !hlock0_p & !cea887;
assign a5f858 = hbusreq3 & a5f7d0 | !hbusreq3 & !a5f857;
assign ce9d49 = hbusreq2_p & ce9d48 | !hbusreq2_p & ce9d46;
assign ab0cab = locked_p & ab0caa | !locked_p & !v84563c;
assign a5edb7 = hbusreq1 & a5edb6 | !hbusreq1 & c3b6a0;
assign a5ea98 = hgrant2_p & a5ea95 | !hgrant2_p & a5ea97;
assign cea3a5 = hlock0_p & cea39c | !hlock0_p & cea380;
assign c3bdff = hready & dead18 | !hready & !v84563c;
assign a5efd1 = hlock2_p & a5efd0 | !hlock2_p & a5ef59;
assign ab0afa = hready & ab0af9 | !hready & v84563c;
assign c3b73a = hbusreq2_p & c3b652 | !hbusreq2_p & c3b739;
assign a5f86a = hlock1_p & a5fa1c | !hlock1_p & v84565a;
assign af352f = hlock1_p & v84563c | !hlock1_p & af352e;
assign c3b6b5 = hgrant2_p & c3b6b3 | !hgrant2_p & c3b6b4;
assign a5f6db = hgrant2_p & a5fa57 | !hgrant2_p & a5fa6f;
assign b2a002 = locked_p & v84563c | !locked_p & !c3bdff;
assign b29d3e = hgrant2_p & b29d38 | !hgrant2_p & b29d3d;
assign af34ae = locked_p & d40d33 | !locked_p & af3c56;
assign a60142 = hlock0_p & a60141 | !hlock0_p & v84563c;
assign cea860 = hbusreq3 & cea85f | !hbusreq3 & v84563c;
assign cea3be = hgrant1_p & cea3bd | !hgrant1_p & cea255;
assign deae62 = hbusreq2_p & deae61 | !hbusreq2_p & deae60;
assign a5ee5c = hlock1_p & a5fbe5 | !hlock1_p & a5ee55;
assign a5ee9a = hmaster1_p & a5ee99 | !hmaster1_p & v84563c;
assign ab05eb = hmaster0_p & ab05e2 | !hmaster0_p & ab05ea;
assign c3b81f = hlock0_p & c3bdbf | !hlock0_p & !cea17a;
assign a5f4f3 = hlock2_p & a5f4ec | !hlock2_p & a5f4f2;
assign c3bc92 = hlock2_p & c3bc91 | !hlock2_p & !dead21;
assign b29a3c = hlock0_p & c3bce0 | !hlock0_p & !v84563c;
assign a5ee9e = locked_p & a5ee4e | !locked_p & a5f36e;
assign a5efa5 = hmaster0_p & a5ef9c | !hmaster0_p & a5efa4;
assign b298aa = locked_p & c3bbba | !locked_p & cea37b;
assign af35a4 = hmaster0_p & af35a3 | !hmaster0_p & af3534;
assign b29e4e = hlock2 & b29e4d | !hlock2 & dead77;
assign c3bc05 = hlock2_p & c3bc04 | !hlock2_p & !v84563c;
assign cea195 = decide_p & cea194 | !decide_p & a57859;
assign b2999a = hgrant0_p & b2997b | !hgrant0_p & !b29999;
assign a5fcfa = hlock1_p & a5fcdd | !hlock1_p & a5fcf9;
assign a5f010 = hgrant0_p & a5eff9 | !hgrant0_p & a5f00f;
assign d40d58 = hbusreq2_p & d40d31 | !hbusreq2_p & d40d33;
assign b8acf3 = jx0_p & b8acf2 | !jx0_p & v84563c;
assign b29d5f = hlock2_p & v84563c | !hlock2_p & !b29d5e;
assign deae07 = hlock2_p & deae06 | !hlock2_p & v84563c;
assign cea29a = hgrant2_p & cea298 | !hgrant2_p & cea299;
assign a5eef9 = hmaster0_p & a5eef8 | !hmaster0_p & a5f58a;
assign a5f2e8 = hlock0_p & a5f2e7 | !hlock0_p & v84563c;
assign b29909 = hbusreq2_p & b29908 | !hbusreq2_p & v84563c;
assign b29a79 = hlock0_p & b29a78 | !hlock0_p & !deadb2;
assign a9b9e7 = hmaster1_p & a9b9e6 | !hmaster1_p & !v84563c;
assign ab0644 = hbusreq2_p & ab0bda | !hbusreq2_p & ab0b23;
assign a5fb30 = hready & a60167 | !hready & v84563c;
assign a5f917 = hlock1_p & a5fa1c | !hlock1_p & !deadd4;
assign ab05a2 = hlock1_p & dead6e | !hlock1_p & !ab05a1;
assign a5efce = decide_p & a5efc6 | !decide_p & a5efcd;
assign cea157 = hmaster1_p & cea14f | !hmaster1_p & cea156;
assign a5f090 = hmaster0_p & a5f087 | !hmaster0_p & a5f08f;
assign cea408 = hgrant1_p & cea407 | !hgrant1_p & cea255;
assign a5f714 = hmastlock_p & a81cda | !hmastlock_p & !v84563c;
assign af34ca = hgrant2_p & af34c6 | !hgrant2_p & af34c9;
assign c3bd25 = hbusreq2_p & c3bd24 | !hbusreq2_p & v84565a;
assign c3bd39 = stateG10_1_p & c3bd38 | !stateG10_1_p & c3bd37;
assign cea40b = hready & cea409 | !hready & cea40a;
assign a5fcbb = hbusreq0_p & c3bcf8 | !hbusreq0_p & a5fc71;
assign a5f840 = stateG10_1_p & adaec6 | !stateG10_1_p & a5f83f;
assign a5ea94 = hbusreq2 & a5f0a8 | !hbusreq2 & a5ea8f;
assign a5f4ba = hlock2 & a5f496 | !hlock2 & a5f4b9;
assign ab0beb = hbusreq2_p & ab0bea | !hbusreq2_p & v845644;
assign a5f2f1 = hready & a5fc21 | !hready & !b26734;
assign a5efa1 = hlock0_p & a5ee23 | !hlock0_p & !a5efa0;
assign c3b65b = decide_p & c3b65a | !decide_p & v845660;
assign dea6d0 = hlock0_p & dea6cf | !hlock0_p & !deadba;
assign aa0e0c = jx2_p & v84563c | !jx2_p & !aa0e0b;
assign a5ee41 = hgrant2_p & a5ee40 | !hgrant2_p & v84563c;
assign b29a82 = hgrant1_p & deada8 | !hgrant1_p & c3b691;
assign bdb580 = hmaster1_p & v845660 | !hmaster1_p & !v84563c;
assign cea3bf = hlock1_p & v84563c | !hlock1_p & !cea3be;
assign deac34 = hbusreq2_p & deac1f | !hbusreq2_p & deac1e;
assign ab0b4e = hmaster0_p & ab0b36 | !hmaster0_p & ab0b4d;
assign c3bbbb = locked_p & v84563c | !locked_p & c3bbba;
assign a5eb9d = hbusreq0 & a5eb9c | !hbusreq0 & v84563c;
assign b29a47 = hmaster0_p & b29a44 | !hmaster0_p & b29a46;
assign a5eec9 = hmaster0_p & a5eeb6 | !hmaster0_p & a5eec8;
assign a5ea4d = locked_p & v845641 | !locked_p & v84563c;
assign c3b708 = hbusreq2_p & c3b707 | !hbusreq2_p & !c3b6e0;
assign c3b88d = hlock2_p & c3b814 | !hlock2_p & c3b829;
assign b29f81 = hmaster1_p & b29f75 | !hmaster1_p & !b29f80;
assign b29f59 = hlock2 & deacc5 | !hlock2 & b29f58;
assign c3b738 = hbusreq0_p & v845648 | !hbusreq0_p & c3b72f;
assign deae16 = hmaster1_p & deae10 | !hmaster1_p & deae15;
assign ab0592 = hlock0_p & ab0590 | !hlock0_p & ab0591;
assign dea725 = hlock0_p & dead72 | !hlock0_p & dead77;
assign a5f927 = hmaster1_p & a5f90c | !hmaster1_p & a5f926;
assign a5f99e = hgrant2_p & a5fbc4 | !hgrant2_p & a5f99d;
assign ab0bda = hlock2_p & ab0bd9 | !hlock2_p & ab0b23;
assign c3b71e = hlock1_p & deadb9 | !hlock1_p & deadba;
assign a5fa20 = hlock1_p & a5fa1c | !hlock1_p & a5fa1f;
assign ab0514 = hbusreq2_p & ab0512 | !hbusreq2_p & ab0513;
assign c3b6f7 = hbusreq2_p & c3b6d7 | !hbusreq2_p & c3b6f6;
assign c3be04 = hgrant2_p & c3bc6d | !hgrant2_p & c3be03;
assign b29d69 = hlock2_p & v845660 | !hlock2_p & b29d68;
assign a5ea6b = hbusreq0 & a5ea6a | !hbusreq0 & a5fbc1;
assign c3bc35 = hlock2_p & v84565a | !hlock2_p & !v84563c;
assign c3b6a4 = stateG10_1_p & deada8 | !stateG10_1_p & c3b691;
assign deae36 = hbusreq3 & deae34 | !hbusreq3 & deae35;
assign cea47e = hbusreq2_p & cea47d | !hbusreq2_p & cea3cd;
assign c3b621 = jx0_p & c3bcd8 | !jx0_p & c3b620;
assign jx0 = !af35c5;
assign c3b8b1 = hbusreq2_p & c3b7dd | !hbusreq2_p & c3b8b0;
assign bdb59d = hmaster1_p & dead2e | !hmaster1_p & v845660;
assign b29a98 = hlock2_p & b29d39 | !hlock2_p & !b29a7c;
assign c3bd5e = hready & c3bd5c | !hready & c3bd5d;
assign b29b25 = hmaster1_p & b29b24 | !hmaster1_p & b29aab;
assign a5f1f4 = locked_p & a5f1f3 | !locked_p & a5f9a2;
assign ce9cd3 = decide_p & ce9cd2 | !decide_p & v84563c;
assign a5f53a = hgrant1_p & a5f539 | !hgrant1_p & deadd3;
assign cea43b = hbusreq2_p & cea43a | !hbusreq2_p & cea414;
assign b26767 = decide_p & b26707 | !decide_p & !b26765;
assign a5fc91 = locked_p & a5fc90 | !locked_p & v84563c;
assign a5eedf = hbusreq2_p & a5eede | !hbusreq2_p & a5eedd;
assign a5fb2c = hbusreq2 & a5fb2b | !hbusreq2 & !v84563c;
assign a81cf2 = hbusreq0_p & a81cc8 | !hbusreq0_p & a81cf1;
assign b2991a = hlock1_p & deaca1 | !hlock1_p & !b29919;
assign ab0631 = hmaster1_p & ab0630 | !hmaster1_p & ab0bee;
assign cea458 = hgrant2_p & cea457 | !hgrant2_p & !cea15c;
assign ab0c82 = hready_p & ab0c2d | !hready_p & ab0c81;
assign c3b895 = hgrant0_p & c3bc5e | !hgrant0_p & c3b894;
assign a5f1e1 = hready & a5f1e0 | !hready & a5fbae;
assign a5f6e9 = hready & v84563c | !hready & b26695;
assign c3bdd1 = hlock0_p & c3bdcf | !hlock0_p & !c3bdd0;
assign cea3a6 = hlock2_p & cea3a5 | !hlock2_p & cea380;
assign a5eeac = hlock0_p & a5f387 | !hlock0_p & a5ee6d;
assign c3b6dc = hbusreq2_p & c3b6d8 | !hbusreq2_p & c3b6db;
assign b29956 = hgrant2_p & b2991e | !hgrant2_p & b29930;
assign b29a21 = hbusreq3_p & b29a20 | !hbusreq3_p & b29ea3;
assign a5f07b = hbusreq2_p & a5f07a | !hbusreq2_p & a5f077;
assign af34b2 = hgrant2_p & af34ad | !hgrant2_p & af34b1;
assign b29a9b = hmaster1_p & b29a9a | !hmaster1_p & b299ed;
assign cea0ca = hbusreq2_p & cea0b9 | !hbusreq2_p & v84563c;
assign ab0c17 = hbusreq3 & ab0c16 | !hbusreq3 & v84563c;
assign ab0635 = hbusreq2_p & ab0573 | !hbusreq2_p & !ab05fa;
assign a5f40d = hready & a5f3f3 | !hready & a5f40c;
assign adaeba = stateG2_p & v84563c | !stateG2_p & d5edb8;
assign a5f972 = hlock2 & a5f96e | !hlock2 & a5f971;
assign b29f5b = hbusreq2_p & b29f5a | !hbusreq2_p & v84565a;
assign a5eaf0 = hbusreq0 & a5eaee | !hbusreq0 & a5eaef;
assign a5f1cf = hlock0_p & a5f6ea | !hlock0_p & a5f96d;
assign cea1c0 = hlock0_p & cea1bf | !hlock0_p & v84563c;
assign ce9cdd = hgrant3_p & ce9cd4 | !hgrant3_p & ce9cdc;
assign adaefa = decide_p & adaee8 | !decide_p & adaef9;
assign v970407 = start_p & v8e1935 | !start_p & v84563c;
assign ab059a = hlock2 & ab0510 | !hlock2 & ab0599;
assign a5f3da = hbusreq0_p & a5f3d2 | !hbusreq0_p & a5f3d8;
assign ab0c94 = hgrant2_p & ab0b70 | !hgrant2_p & ab0c93;
assign a5f1c1 = hgrant0_p & a5f99a | !hgrant0_p & a5f1c0;
assign a5fbce = hbusreq2_p & a5fbcd | !hbusreq2_p & a5fbcc;
assign a5f8ee = hlock2 & a5fb4d | !hlock2 & a5f8ed;
assign b29b1e = hlock2 & b29b1c | !hlock2 & b29b1d;
assign deacad = hbusreq2_p & deacac | !hbusreq2_p & v84563c;
assign a5fc1d = hlock0_p & a5fc1a | !hlock0_p & a5fc1c;
assign a5ee57 = hbusreq1 & a5ee56 | !hbusreq1 & !v84563c;
assign ab0c26 = hlock0_p & v84563c | !hlock0_p & !ab0c25;
assign a5f08f = hmaster1_p & a5f08e | !hmaster1_p & a60145;
assign deac19 = hlock1_p & v84563c | !hlock1_p & deac18;
assign cea482 = hready & cea481 | !hready & cea333;
assign d40d8f = hmaster0_p & d40d8e | !hmaster0_p & v84563c;
assign deae2c = hlock3_p & deae2b | !hlock3_p & deadf4;
assign cea393 = hbusreq0_p & cea38a | !hbusreq0_p & cea38e;
assign af3c67 = hmaster1_p & af3c61 | !hmaster1_p & af3c66;
assign deae39 = hmaster1_p & deae36 | !hmaster1_p & deae38;
assign adaec1 = decide_p & adaec0 | !decide_p & adaebf;
assign ab05dd = hbusreq2_p & ab05aa | !hbusreq2_p & ab05dc;
assign ab0c78 = hlock0_p & ab0c77 | !hlock0_p & !ab0c5d;
assign a5f2ed = hmaster0_p & a5f2ec | !hmaster0_p & a5f999;
assign dead91 = hbusreq3 & dead8e | !hbusreq3 & dead90;
assign b266cc = hgrant1_p & b266ca | !hgrant1_p & b266cb;
assign a5f08a = hbusreq2 & a5f089 | !hbusreq2 & a5fb6c;
assign af3490 = hmaster0_p & af3488 | !hmaster0_p & af348f;
assign a5fb96 = hlock0_p & a5fb95 | !hlock0_p & a5fb92;
assign b29d88 = locked_p & v84563c | !locked_p & !b29d87;
assign dea769 = hbusreq2_p & deae0e | !hbusreq2_p & dea768;
assign ab06bf = hlock2 & ab06b8 | !hlock2 & ab06be;
assign ab06fc = hbusreq2_p & ab06fb | !hbusreq2_p & b29ab2;
assign b26775 = hmaster1_p & b26774 | !hmaster1_p & b26711;
assign ab053c = hlock1_p & v84563c | !hlock1_p & ab053b;
assign d40d7d = hlock0_p & d40d31 | !hlock0_p & d40d7c;
assign ab0b37 = hlock0_p & v84563c | !hlock0_p & c3bd60;
assign a5fbb6 = hmastlock_p & a5fbb5 | !hmastlock_p & v84563c;
assign b29974 = hmaster1_p & b29973 | !hmaster1_p & b29956;
assign af34d9 = hlock2_p & af3c50 | !hlock2_p & af3c6b;
assign b29939 = hlock1_p & deac51 | !hlock1_p & !c3b693;
assign a5f8e8 = hgrant1_p & v84563c | !hgrant1_p & b29923;
assign af3575 = hmaster1_p & af3572 | !hmaster1_p & af3574;
assign b29ecb = hmaster1_p & b29ec4 | !hmaster1_p & b29eca;
assign a5eae9 = hbusreq2 & a5eae6 | !hbusreq2 & a5eae8;
assign a5fd27 = hlock2_p & a5fd22 | !hlock2_p & a5fd26;
assign ab0742 = hlock2_p & ab06eb | !hlock2_p & ab06fd;
assign a5fc74 = hburst1_p & d615cf | !hburst1_p & !v84563c;
assign c3bbe2 = hready & cea29f | !hready & v845648;
assign a5fc85 = stateA1_p & a81ca7 | !stateA1_p & !cea1ac;
assign a5f35d = hmaster0_p & a5f35c | !hmaster0_p & a5f288;
assign a5ef0a = hready & a5ef07 | !hready & a5ef09;
assign ab05c4 = hmaster0_p & ab05bc | !hmaster0_p & ab05c3;
assign a5f110 = hlock0_p & a5f806 | !hlock0_p & a5f108;
assign v97044f = hmaster1_p & v9703fc | !hmaster1_p & v970413;
assign deae6c = hbusreq3 & deae6b | !hbusreq3 & !v84563c;
assign b29f97 = hbusreq2_p & b29f96 | !hbusreq2_p & v84563c;
assign a5f2fb = hmaster1_p & a5f2fa | !hmaster1_p & a5f1b8;
assign af34d0 = hmaster1_p & af34cf | !hmaster1_p & af34a7;
assign a5f6e0 = decide_p & a5f6df | !decide_p & v84563c;
assign deae1e = hlock0_p & deae1d | !hlock0_p & !deada8;
assign ab0c83 = hlock2_p & ab0b5b | !hlock2_p & dead2e;
assign v970416 = hmaster1_p & v97040b | !hmaster1_p & v970413;
assign b29987 = hlock0_p & b29984 | !hlock0_p & !b29986;
assign ce9cce = hgrant3_p & ce9cb3 | !hgrant3_p & ce9ccd;
assign ab067a = hlock0_p & b29ffc | !hlock0_p & v845660;
assign af34e4 = hmaster1_p & af3c70 | !hmaster1_p & af3c50;
assign c3bc4f = hlock2_p & c3bc4c | !hlock2_p & c3bc4e;
assign a5faac = hlock1_p & a6016f | !hlock1_p & !a5faab;
assign a9b9dc = hlock2_p & a9b9d0 | !hlock2_p & v845660;
assign a5f1df = hbusreq1_p & a5f988 | !hbusreq1_p & a5fba6;
assign dead6d = start_p & v845652 | !start_p & !dead6c;
assign ab05b6 = hlock2_p & ab05b2 | !hlock2_p & ab05b5;
assign c3bc7c = hlock0_p & c3bc79 | !hlock0_p & !c3bc7b;
assign deae12 = hlock0_p & deae11 | !hlock0_p & v84563c;
assign c3b6d4 = decide_p & c3b6d3 | !decide_p & v845660;
assign a5f381 = hlock2_p & a5f380 | !hlock2_p & !a5f37f;
assign b2996f = hlock0_p & c3b6c5 | !hlock0_p & deada8;
assign d40d42 = hlock1_p & d40d31 | !hlock1_p & !d40d41;
assign c3bdb5 = hmaster0_p & c3bdac | !hmaster0_p & c3bdb4;
assign b29a91 = hbusreq2_p & b29a8c | !hbusreq2_p & v84563c;
assign a5edac = hlock2 & a5f5a3 | !hlock2 & a5f5a9;
assign a81cdf = hmaster1_p & v84563c | !hmaster1_p & a81cde;
assign v970438 = hbusreq2_p & v970437 | !hbusreq2_p & v84563c;
assign dea737 = hmaster0_p & dea732 | !hmaster0_p & dea736;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hbusreq2_p = 0;
  hlock2_p = 0;
  hbusreq3_p = 0;
  hlock3_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmaster1_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  hgrant2_p = 0;
  hgrant3_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  stateG10_2_p = 0;
  stateG10_3_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hbusreq2_p = hbusreq2;
  hlock2_p = hlock2;
  hbusreq3_p = hbusreq3;
  hlock3_p = hlock3;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmaster1_p = hmaster1;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  hgrant2_p = hgrant2;
  hgrant3_p = hgrant3;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  stateG10_2_p = stateG10_2;
  stateG10_3_p = stateG10_3;
  jx0_p = jx0;
  jx1_p = jx1;
  jx2_p = jx2;
    end
endmodule

