module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, StoB_REQ4_n, StoB_REQ5_n, StoB_REQ6_n, StoB_REQ7_n, StoB_REQ8_n, StoB_REQ9_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoS_ACK4_n, BtoS_ACK5_n, BtoS_ACK6_n, BtoS_ACK7_n, BtoS_ACK8_n, BtoS_ACK9_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, SLC2_n, SLC3_n, jx0_n, jx1_n, jx2_n, jx3_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844fbd;
  wire v90612e;
  wire v9093a9;
  wire v8a1fe3;
  wire v844fa1;
  wire v93f8f0;
  wire v90dd2f;
  wire v905764;
  wire v911fc7;
  wire v911946;
  wire v9091c6;
  wire v9078da;
  wire v903d1e;
  wire v908429;
  wire v9093ec;
  wire v90adcb;
  wire v906046;
  wire v844f9f;
  wire v91058e;
  wire v9076a8;
  wire v93dffe;
  wire v93fc02;
  wire v93e681;
  wire v903e85;
  wire v844f9d;
  wire v87a21f;
  wire v93e2de;
  wire v9134df;
  wire v863a78;
  wire v9132b0;
  wire v911509;
  wire v9122e7;
  wire v9097c3;
  wire v844f9b;
  wire v9052de;
  wire v910f6e;
  wire v910243;
  wire v90962d;
  wire v93faf8;
  wire v90776b;
  wire v8b98d4;
  wire v910710;
  wire v93f744;
  wire v90da41;
  wire v87a1d0;
  wire v911ebf;
  wire v93f838;
  wire v93e47b;
  wire v93e8f6;
  wire v9057cb;
  wire v90a850;
  wire v844fbb;
  wire v904182;
  wire v9300af;
  wire v863444;
  wire v93f79a;
  wire v910b33;
  wire v906c71;
  wire v93fd50;
  wire v90f8f5;
  wire v90a27c;
  wire v89f9d7;
  wire v90767a;
  wire v905702;
  wire v90a3e0;
  wire v905978;
  wire v93e8d3;
  wire v93f81b;
  wire v90f500;
  wire v93ec83;
  wire v93f41e;
  wire v909dd6;
  wire v89f7e7;
  wire v93e86c;
  wire v9049a9;
  wire v87a1f0;
  wire v90fe49;
  wire v90611f;
  wire v93fc8e;
  wire v909174;
  wire v90a134;
  wire v93f69d;
  wire v93db03;
  wire v93fddd;
  wire v9080a0;
  wire v93e13e;
  wire v910644;
  wire v9098e3;
  wire v90adef;
  wire v93fc81;
  wire v90f994;
  wire v93fa2e;
  wire v93fb85;
  wire v86341e;
  wire v93fde5;
  wire v906a80;
  wire v90e9e1;
  wire v93fbb6;
  wire v93fb5d;
  wire v93fcd0;
  wire v907a33;
  wire v908fb5;
  wire v912190;
  wire v91086f;
  wire v93f698;
  wire v93fcdd;
  wire v90a1c6;
  wire v90a61d;
  wire v909ba1;
  wire v910b96;
  wire v903da9;
  wire v91104c;
  wire v90804e;
  wire v907aa0;
  wire v93fafd;
  wire v8a924b;
  wire v91195c;
  wire v9082d3;
  wire v910820;
  wire v87a1f2;
  wire v9113de;
  wire v90ff24;
  wire v907d33;
  wire v90811c;
  wire v87c9bf;
  wire v906acc;
  wire v93fb5c;
  wire v905d28;
  wire v910f3a;
  wire v93fb13;
  wire v93fa40;
  wire v93fe04;
  wire v90d00f;
  wire v93f864;
  wire v93fdbd;
  wire v90a233;
  wire v9041e4;
  wire v93f8ee;
  wire v906414;
  wire v90569e;
  wire v90999b;
  wire v93f362;
  wire v90932c;
  wire v90e79a;
  wire v91229f;
  wire v8d3791;
  wire v909845;
  wire v90f83e;
  wire v93f07c;
  wire v90cbf3;
  wire v904d51;
  wire v907bd1;
  wire v8a8fa3;
  wire v90469d;
  wire v93e8cc;
  wire v911498;
  wire v91a9a2;
  wire v93fa58;
  wire v93f6db;
  wire v910242;
  wire v9077f7;
  wire v90a241;
  wire v9047b1;
  wire v93fa5e;
  wire v90e774;
  wire v91229e;
  wire v9074a6;
  wire v93f5c0;
  wire v907122;
  wire v8b99b4;
  wire v93f69c;
  wire v87e087;
  wire v905e84;
  wire v9045c0;
  wire v908357;
  wire v909df9;
  wire v93fde4;
  wire v9085b3;
  wire v90631b;
  wire v93fe01;
  wire v93f67b;
  wire v903c5b;
  wire v88b9b7;
  wire v90d6ca;
  wire v93fb03;
  wire v90888d;
  wire v909222;
  wire v908a03;
  wire v93e90d;
  wire v93e948;
  wire v90df02;
  wire v9043a5;
  wire v89e0d7;
  wire v9079ac;
  wire v93fc32;
  wire v93f916;
  wire v90567d;
  wire v9074f5;
  wire v9053ed;
  wire v913a94;
  wire v90927b;
  wire v90cf52;
  wire v85ea96;
  wire v904926;
  wire v910ee7;
  wire v887bb8;
  wire v910d81;
  wire v9042fa;
  wire v907d8f;
  wire v8b9d25;
  wire v907ef2;
  wire v93fa03;
  wire v8b9b9b;
  wire v90809e;
  wire v90aaa8;
  wire v93e731;
  wire v904d7e;
  wire v907d9d;
  wire v90f6b5;
  wire v93fb34;
  wire v9056e2;
  wire v93e037;
  wire v92ffd6;
  wire v93e94e;
  wire v906275;
  wire v9091a2;
  wire v911328;
  wire v8a928a;
  wire v844fcd;
  wire v9081c2;
  wire v844fa9;
  wire v86e7cf;
  wire v90cfd5;
  wire v93fe1a;
  wire v844fcf;
  wire v85eb14;
  wire v93fd98;
  wire v909546;
  wire v8c8823;
  wire v87f17d;
  wire v869aeb;
  wire v87c51f;
  wire v910f82;
  wire v907e86;
  wire v9074fa;
  wire v93fda8;
  wire v93faf2;
  wire v911680;
  wire v93db4a;
  wire v90ea74;
  wire v90ad47;
  wire v906201;
  wire v911090;
  wire v90df44;
  wire v90dfbc;
  wire v91086c;
  wire v93f818;
  wire v93eda4;
  wire v93fdd2;
  wire v909691;
  wire v8d37f5;
  wire v90ad39;
  wire v9079bf;
  wire v908aa8;
  wire v90fb0e;
  wire v93fd0f;
  wire v90db9e;
  wire v90927a;
  wire v863428;
  wire v907417;
  wire v863a3f;
  wire v93e7ac;
  wire v90987f;
  wire v93f793;
  wire v8b9c07;
  wire v904b4f;
  wire v863b2f;
  wire v908e92;
  wire v9052f0;
  wire v93f7f4;
  wire v872e5f;
  wire v93fa96;
  wire v910fcd;
  wire v87c9b3;
  wire v93f9d2;
  wire v908836;
  wire v93f87f;
  wire v9070e2;
  wire v93fd51;
  wire v909337;
  wire v903e7a;
  wire v93f6aa;
  wire v863ad6;
  wire v8b9f15;
  wire v90e3bf;
  wire v905292;
  wire v90738b;
  wire v93e9c8;
  wire v93f74a;
  wire v93fd5f;
  wire v93e648;
  wire v909043;
  wire v9043ec;
  wire v93fbb0;
  wire v93f755;
  wire v90e144;
  wire v9300a5;
  wire v93f6cf;
  wire v8d37d6;
  wire v93fc48;
  wire v93e80c;
  wire v93fc2d;
  wire v9051ae;
  wire v903d68;
  wire v93fbce;
  wire v8ebd2a;
  wire v844fab;
  wire v93fd76;
  wire v907e3f;
  wire v89e10d;
  wire v87f17f;
  wire v93f776;
  wire v93e701;
  wire v903c0d;
  wire v90d8f3;
  wire v93fd59;
  wire v93fc68;
  wire v93fc94;
  wire v90d22b;
  wire v906c8b;
  wire v844f99;
  wire v884481;
  wire v844f97;
  wire v844f95;
  wire v9047e4;
  wire v9060ea;
  wire v8b5f61;
  wire v904234;
  wire v9104ad;
  wire v93fbe5;
  wire v91ae94;
  wire v908127;
  wire v90e611;
  wire v908fba;
  wire v909e2c;
  wire v93fbba;
  wire v9093db;
  wire v93f6a4;
  wire v93f7f5;
  wire v906d08;
  wire v906642;
  wire v9056ad;
  wire v91023b;
  wire v9055bd;
  wire v93f70c;
  wire v93f6fc;
  wire v90fb2b;
  wire v908107;
  wire v909661;
  wire v90cf49;
  wire v8bbc51;
  wire v93f734;
  wire v93fb2a;
  wire v93fbcd;
  wire v909bff;
  wire v910c0f;
  wire v90fe92;
  wire v911311;
  wire v87b4fc;
  wire v93e48f;
  wire v905da3;
  wire v910bf8;
  wire v9054c6;
  wire v93fb29;
  wire v93f216;
  wire v90479a;
  wire v9071c7;
  wire v93f689;
  wire v85eabe;
  wire v906a79;
  wire v911d8e;
  wire v93fe14;
  wire v93f714;
  wire v93f722;
  wire v93f7fb;
  wire v93faf7;
  wire v93e8ab;
  wire v91ddca;
  wire v91053d;
  wire v93faca;
  wire v85f28b;
  wire v93fd1b;
  wire v908e7f;
  wire v904cc8;
  wire v90a18c;
  wire v90f2f8;
  wire v93fbdc;
  wire v90d651;
  wire v93eef4;
  wire v91aa04;
  wire v911bcf;
  wire v9052ba;
  wire v909722;
  wire v911951;
  wire v8ee1a9;
  wire v907ccf;
  wire v904f76;
  wire v8a9267;
  wire v90893a;
  wire v903d0c;
  wire v904e2f;
  wire v93f8bb;
  wire v90606d;
  wire v93fc3e;
  wire v90d972;
  wire v904bcb;
  wire v872442;
  wire v89e08c;
  wire v93fa3a;
  wire v90722c;
  wire v9095bf;
  wire v86f4a3;
  wire v93f9a9;
  wire v93f85e;
  wire v93ea50;
  wire v90ed41;
  wire v863a37;
  wire v913348;
  wire v90a5ef;
  wire v93fa55;
  wire v8bb868;
  wire v90a6f4;
  wire v93fa90;
  wire v90a9e4;
  wire v86313d;
  wire v911451;
  wire v93fb09;
  wire v93e77b;
  wire v93fc9b;
  wire v904e70;
  wire v912687;
  wire v93f9c6;
  wire v93f7f1;
  wire v905718;
  wire v910b7a;
  wire v903b7c;
  wire v93f7d9;
  wire v904cb5;
  wire v90ddf9;
  wire v93fdc9;
  wire v93fe2d;
  wire v93fc09;
  wire v907ce3;
  wire v93fc75;
  wire v8b4990;
  wire v93efbb;
  wire v93f6ce;
  wire v905434;
  wire v90f864;
  wire v93ec07;
  wire v904fc8;
  wire v903f21;
  wire v89e0da;
  wire v93fc65;
  wire v93fe2b;
  wire v8f382c;
  wire v907048;
  wire v872746;
  wire v93fe34;
  wire v89f840;
  wire v93f765;
  wire v90ad2f;
  wire v9300c0;
  wire v908c12;
  wire v93eaa8;
  wire v93f6d3;
  wire v90a29a;
  wire v90815c;
  wire v93faec;
  wire v88d074;
  wire v93e898;
  wire v903d90;
  wire v90e93c;
  wire v90f810;
  wire v90474e;
  wire v90f2de;
  wire v93ef1d;
  wire v905eaa;
  wire v9102bf;
  wire v90add3;
  wire v93fbf0;
  wire v87a1f9;
  wire v909927;
  wire v910f51;
  wire v903e7f;
  wire v8633b7;
  wire v9083d0;
  wire v8b9dbd;
  wire v90f7a1;
  wire v9054b5;
  wire v90664a;
  wire v93fc2b;
  wire v904dd8;
  wire v93f3a8;
  wire v910c50;
  wire v93fa5b;
  wire v93fc10;
  wire v93f78a;
  wire v8b9ba5;
  wire v909a70;
  wire v93f2a2;
  wire v93daf2;
  wire v904b99;
  wire v910230;
  wire v930036;
  wire v90caf3;
  wire v903d5e;
  wire v9132dc;
  wire v9083f0;
  wire v912f4e;
  wire v907fc6;
  wire v93fd3a;
  wire v909ecc;
  wire v90817e;
  wire v906195;
  wire v9059a0;
  wire v93f75c;
  wire v93f8d1;
  wire v907e6b;
  wire v8ee188;
  wire v908743;
  wire v8b9f38;
  wire v9121b6;
  wire v93f682;
  wire v908e8e;
  wire v90dcfd;
  wire v912291;
  wire v86dc4b;
  wire v904afe;
  wire v906c3f;
  wire v93fb33;
  wire v885188;
  wire v909be8;
  wire v9048c6;
  wire v93f770;
  wire v93e150;
  wire v85f240;
  wire v912265;
  wire v93f9f6;
  wire v93e816;
  wire v93f9e7;
  wire v910461;
  wire v93e105;
  wire v9080c5;
  wire v93f955;
  wire v904628;
  wire v909dde;
  wire v85cd12;
  wire v93fb92;
  wire v93e85e;
  wire v93ee3b;
  wire v93fa1f;
  wire v93ecb9;
  wire v93f769;
  wire v909e8a;
  wire v93fd75;
  wire v906ec1;
  wire v93fb41;
  wire v911b50;
  wire v93e9ea;
  wire v88d7c9;
  wire v913662;
  wire v90e8da;
  wire v93fb81;
  wire v910f4e;
  wire v89f920;
  wire v93e713;
  wire v907f31;
  wire v90e02c;
  wire v910d99;
  wire v91355f;
  wire v89e086;
  wire v93f6ad;
  wire v93fb26;
  wire v9051ba;
  wire v904c80;
  wire v904345;
  wire v9057f8;
  wire v905d68;
  wire v9042a0;
  wire v93fe73;
  wire v907b84;
  wire v87f181;
  wire v87d990;
  wire v907301;
  wire v93e203;
  wire v9114cf;
  wire v93e281;
  wire v863abb;
  wire v91a6ea;
  wire v93f694;
  wire v93fb19;
  wire v909e99;
  wire v93fe0a;
  wire v8d371f;
  wire v91315c;
  wire v9091b4;
  wire v904ff8;
  wire v93e288;
  wire v90ad75;
  wire v905ba8;
  wire v93f71d;
  wire v908d14;
  wire v909c74;
  wire v90dcf6;
  wire v93fa74;
  wire v91334f;
  wire v8b9c3a;
  wire v904a8a;
  wire v863359;
  wire v8f37fc;
  wire v93fd42;
  wire v9056a0;
  wire v93fbf4;
  wire v93fc89;
  wire v89e05b;
  wire v90cf68;
  wire v90d443;
  wire v90a4bb;
  wire v910c29;
  wire v90859f;
  wire v9117b1;
  wire v90ea51;
  wire v93fe36;
  wire v93f824;
  wire v93df06;
  wire v93f0b0;
  wire v904432;
  wire v90df4b;
  wire v93f1c4;
  wire v93fdb2;
  wire v93f9bc;
  wire v883cbe;
  wire v93fe46;
  wire v90a348;
  wire v90a525;
  wire v93f82b;
  wire v906f55;
  wire v8b4976;
  wire v93faa1;
  wire v9087b1;
  wire v9087d1;
  wire v858fc9;
  wire v910bb8;
  wire v90d5a3;
  wire v906a6b;
  wire v93fc40;
  wire v8b4a08;
  wire v90636b;
  wire v93fbcf;
  wire v911853;
  wire v93fddc;
  wire v93f883;
  wire v93e882;
  wire v90a7b2;
  wire v93f7ea;
  wire v904200;
  wire v9060d2;
  wire v93f9f3;
  wire v93fa84;
  wire v93f5b9;
  wire v8b9bb4;
  wire v8b98b7;
  wire v904013;
  wire v89e06e;
  wire v904d81;
  wire v90f8ce;
  wire v904632;
  wire v909197;
  wire v88bb45;
  wire v90831e;
  wire v90467c;
  wire v93f9bf;
  wire v908cff;
  wire v905146;
  wire v9085f5;
  wire v90d7d2;
  wire v9131cb;
  wire v910f41;
  wire v87cb21;
  wire v844fb3;
  wire v909082;
  wire v8b49f1;
  wire v911c0f;
  wire v93f87b;
  wire v90adc4;
  wire v93fcbe;
  wire v93fce5;
  wire v9099e1;
  wire v907607;
  wire v93e577;
  wire v93f685;
  wire v90f2ff;
  wire v93fcdb;
  wire v907be9;
  wire v9121bb;
  wire v93f9ac;
  wire v93fd9c;
  wire v908d55;
  wire v93e7af;
  wire v93e89f;
  wire v911c6f;
  wire v93fc04;
  wire v90980d;
  wire v93fd9e;
  wire v9123a2;
  wire v906627;
  wire v93fdfe;
  wire v910cf1;
  wire v90873f;
  wire v90e6e5;
  wire v90db9f;
  wire v93fcd4;
  wire v904779;
  wire v910825;
  wire v871033;
  wire v9047b7;
  wire v90937e;
  wire v9072c8;
  wire v909f4c;
  wire v9075d4;
  wire v93fb68;
  wire v93f66f;
  wire v8a8fed;
  wire v91879a;
  wire v93f148;
  wire v905810;
  wire v87c525;
  wire v90a784;
  wire v93e76f;
  wire v93e8cb;
  wire v93fb08;
  wire v905d04;
  wire v93fca0;
  wire v905adf;
  wire v9080f5;
  wire v93fe1b;
  wire v90a89f;
  wire v85ea99;
  wire v90fc5e;
  wire v87a97c;
  wire v93fbd6;
  wire v93fd11;
  wire v90eed2;
  wire v90acaa;
  wire v93fb64;
  wire v93fbe6;
  wire v93ee22;
  wire v90a102;
  wire v93f9f4;
  wire v90a8c3;
  wire v90e7d7;
  wire v90decc;
  wire v93f9dd;
  wire v93e602;
  wire v90603e;
  wire v8b9e12;
  wire v8f229e;
  wire v913522;
  wire v93f709;
  wire v93f941;
  wire v8839a7;
  wire v910383;
  wire v93fdd5;
  wire v907017;
  wire v90d22a;
  wire v907e91;
  wire v903c81;
  wire v93fa3d;
  wire v905a21;
  wire v904e00;
  wire v90851b;
  wire v90ff7e;
  wire v910e44;
  wire v93f6a0;
  wire v905d97;
  wire v93f8d3;
  wire v93fcc8;
  wire v9117e5;
  wire v93fd60;
  wire v90e019;
  wire v905b55;
  wire v863b26;
  wire v90dc0d;
  wire v90664c;
  wire v93f69a;
  wire v93f107;
  wire v85eaff;
  wire v909cea;
  wire v90da8b;
  wire v93fb93;
  wire v9043fc;
  wire v9121a7;
  wire v90d7a0;
  wire v89f8bc;
  wire v91a992;
  wire v93e296;
  wire v90dd77;
  wire v93fb38;
  wire v93e896;
  wire v908d05;
  wire v870fb9;
  wire v93def0;
  wire v93fbb9;
  wire v90526b;
  wire v8a9209;
  wire v9103b5;
  wire v90f309;
  wire v9056f9;
  wire v91231a;
  wire v911b4d;
  wire v90ada1;
  wire v90936b;
  wire v93e2fa;
  wire v93f51d;
  wire v908f29;
  wire v93fb45;
  wire v9098bb;
  wire v881ec0;
  wire v90a002;
  wire v913a60;
  wire v93fb1d;
  wire v907f0e;
  wire v910dda;
  wire v910c4e;
  wire v90931a;
  wire v8f381e;
  wire v93fe69;
  wire v909fd6;
  wire v93f1a6;
  wire v904c53;
  wire v910525;
  wire v90e073;
  wire v90a541;
  wire v93f389;
  wire v89e07c;
  wire v8b9bd8;
  wire v93005b;
  wire v930037;
  wire v93f70d;
  wire v909224;
  wire v911a1e;
  wire v91071f;
  wire v90e159;
  wire v93f871;
  wire v90a62c;
  wire v93e259;
  wire v90a926;
  wire v93f69b;
  wire v90a6d8;
  wire v93f766;
  wire v912ef3;
  wire v90f1b9;
  wire v90d634;
  wire v93fc0f;
  wire v909f4b;
  wire v907b86;
  wire v93fb39;
  wire v90fbfd;
  wire v905d2c;
  wire v93f6a6;
  wire v93f9a7;
  wire v905a88;
  wire v90add9;
  wire v93fafc;
  wire v8b9ecf;
  wire v9056b0;
  wire v93fc77;
  wire v93fe3f;
  wire v93e3a1;
  wire v904da8;
  wire v911bb8;
  wire v93f87c;
  wire v93e440;
  wire v93f0a7;
  wire v9097bf;
  wire v859639;
  wire v8a921d;
  wire v9101d0;
  wire v9085e8;
  wire v905dc1;
  wire v87c4e7;
  wire v89f7c7;
  wire v903b0f;
  wire v9132f8;
  wire v93fd64;
  wire v90de74;
  wire v8b9972;
  wire v90fa88;
  wire v90f629;
  wire v90cc4a;
  wire v911933;
  wire v90e361;
  wire v93fe5d;
  wire v906769;
  wire v93fa06;
  wire v911a92;
  wire v90767c;
  wire v90d6e8;
  wire v93f754;
  wire v904f32;
  wire v93f696;
  wire v89b107;
  wire v86345d;
  wire v90e8f5;
  wire v908eea;
  wire v93fbd2;
  wire v912ec8;
  wire v908553;
  wire v907468;
  wire v93e1dc;
  wire v93f853;
  wire v93f7fa;
  wire v908805;
  wire v91043e;
  wire v9104ca;
  wire v93fac1;
  wire v93f290;
  wire v907cc6;
  wire v93fabf;
  wire v9051e9;
  wire v87bf17;
  wire v908d1f;
  wire v90aa64;
  wire v913a54;
  wire v8f37f3;
  wire v906d3f;
  wire v93fca7;
  wire v910d5a;
  wire v90e1dd;
  wire v93fa66;
  wire v904f85;
  wire v906e08;
  wire v90a3f5;
  wire v90e612;
  wire v91247e;
  wire v93ecf7;
  wire v8b4a10;
  wire v90523b;
  wire v9135e7;
  wire v9049ac;
  wire v9080a7;
  wire v90813f;
  wire v887a80;
  wire v93fa4d;
  wire v9100b7;
  wire v909f00;
  wire v908acd;
  wire v93fda4;
  wire v89f95b;
  wire v93f75f;
  wire v93f7d5;
  wire v90ea98;
  wire v93eb1d;
  wire v93f0b8;
  wire v910d2f;
  wire v93f9fe;
  wire v903b68;
  wire v90d59e;
  wire v93fb74;
  wire v90799d;
  wire v906f72;
  wire v93e0c9;
  wire v8b9c01;
  wire v93f746;
  wire v91a733;
  wire v904d40;
  wire v9064cc;
  wire v904e3e;
  wire v909efe;
  wire v90f7a9;
  wire v91db5b;
  wire v910d62;
  wire v85ea72;
  wire v9102bb;
  wire v91a6dc;
  wire v93fb80;
  wire v93f6b6;
  wire v8b6034;
  wire v844fc1;
  wire v93f753;
  wire v844fa5;
  wire v93fde7;
  wire v9063d8;
  wire v911452;
  wire v93fdcc;
  wire v93ed00;
  wire v93fd3d;
  wire v90df7f;
  wire v93e310;
  wire v93f63b;
  wire v904adb;
  wire v9099ee;
  wire v93f860;
  wire v93fc15;
  wire v904c52;
  wire v93fa16;
  wire v912cf4;
  wire v93fc71;
  wire v8bbc68;
  wire v91104b;
  wire v93fc64;
  wire v93facb;
  wire v905824;
  wire v909eab;
  wire v9078b3;
  wire v9104d5;
  wire v903fee;
  wire v907102;
  wire v93f70b;
  wire v910f62;
  wire v93fd94;
  wire v93ef57;
  wire v872067;
  wire v9044b1;
  wire v89fe58;
  wire v930005;
  wire v910515;
  wire v93fdbc;
  wire v91a747;
  wire v93faf5;
  wire v9063b2;
  wire v93fd2e;
  wire v91343f;
  wire v93e262;
  wire v93fa54;
  wire v93f827;
  wire v93fad2;
  wire v90470d;
  wire v93f7e6;
  wire v93ec1d;
  wire v91a6d3;
  wire v910289;
  wire v90711a;
  wire v93f1ad;
  wire v93f2a4;
  wire v908237;
  wire v93fcc4;
  wire v908073;
  wire v93f6dd;
  wire v909dcc;
  wire v90549c;
  wire v90a196;
  wire v911428;
  wire v93fa9c;
  wire v904f64;
  wire v9124b8;
  wire v90a2fc;
  wire v93fdd4;
  wire v93f8bf;
  wire v9051d8;
  wire v90531e;
  wire v93f91a;
  wire v90e433;
  wire v93fdfd;
  wire v909e28;
  wire v90897e;
  wire v93e800;
  wire v93fa52;
  wire v9057d4;
  wire v93f1cb;
  wire v93ed15;
  wire v909bdf;
  wire v9082be;
  wire v90e9a1;
  wire v93e751;
  wire v93fdda;
  wire v90e261;
  wire v906338;
  wire v93e115;
  wire v906491;
  wire v93f39f;
  wire v9061f2;
  wire v93faa8;
  wire v907679;
  wire v93e9d8;
  wire v89f8b8;
  wire v93f85b;
  wire v93fa69;
  wire v90930e;
  wire v93ef40;
  wire v92fffd;
  wire v8633ec;
  wire v906b4a;
  wire v93f634;
  wire v863a00;
  wire v90775f;
  wire v93fc24;
  wire v93f751;
  wire v907c69;
  wire v89c5bd;
  wire v90606c;
  wire v905199;
  wire v85ea93;
  wire v904f5e;
  wire v9051cd;
  wire v903cef;
  wire v905246;
  wire v90e5b4;
  wire v93e3f1;
  wire v9042d2;
  wire v93e189;
  wire v93f19b;
  wire v908df3;
  wire v90926e;
  wire v90575e;
  wire v90e140;
  wire v93fb1c;
  wire v904074;
  wire v90fcd2;
  wire v93e589;
  wire v904f2e;
  wire v8b9e17;
  wire v93e9d1;
  wire v908e52;
  wire v93fd8f;
  wire v8b4a13;
  wire v93ebb5;
  wire v93e0a0;
  wire v905636;
  wire v90901d;
  wire v9084ef;
  wire v93fb24;
  wire v93f7be;
  wire v93f785;
  wire v93f06e;
  wire v93f825;
  wire v90968f;
  wire v90fa80;
  wire v90490e;
  wire v93f784;
  wire v9103e5;
  wire v93e548;
  wire v93e838;
  wire v93fd19;
  wire v905ba4;
  wire v903bf8;
  wire v93f918;
  wire v93f856;
  wire v90ef1a;
  wire v90ba31;
  wire v93f917;
  wire v903b56;
  wire v93f830;
  wire v906d83;
  wire v911586;
  wire v93f9f5;
  wire v904253;
  wire v863a64;
  wire v91047b;
  wire v904b1b;
  wire v93ea7f;
  wire v90fb00;
  wire v903cd1;
  wire v909a08;
  wire v909dc9;
  wire v8b99c6;
  wire v844fc3;
  wire v9046a7;
  wire v93f937;
  wire v906b64;
  wire v912fc9;
  wire v90a23c;
  wire v93f3f2;
  wire v91209b;
  wire v907200;
  wire v90f4dd;
  wire v93fdc0;
  wire v90834a;
  wire v93e671;
  wire v90dc57;
  wire v93efb8;
  wire v904677;
  wire v904b94;
  wire v904c4f;
  wire v93f8a3;
  wire v90583b;
  wire v9050ba;
  wire v93fbcc;
  wire v87c541;
  wire v907b07;
  wire v93ea9e;
  wire v93ef38;
  wire v90ed7e;
  wire v90712d;
  wire v93f897;
  wire v911826;
  wire v93e682;
  wire v93f6d0;
  wire v8a9250;
  wire v905291;
  wire v93f7a1;
  wire v90a774;
  wire v90748c;
  wire v90fa03;
  wire v91a70f;
  wire v93fd4a;
  wire v912d1a;
  wire v904e3a;
  wire v93f90f;
  wire v904fee;
  wire v904d56;
  wire v90542e;
  wire v93f729;
  wire v93f6c4;
  wire v8b9bbf;
  wire v90620e;
  wire v93f7fc;
  wire v90536f;
  wire v90ed80;
  wire v907bb9;
  wire v90505e;
  wire v87261e;
  wire v9082e6;
  wire v91007f;
  wire v9078eb;
  wire v9094f2;
  wire v90de0e;
  wire v905b6a;
  wire v9096ca;
  wire v93f56e;
  wire v913399;
  wire v904fd6;
  wire v910b22;
  wire v90a1c0;
  wire v88c2af;
  wire v908ffc;
  wire v911435;
  wire v90f0c5;
  wire v906034;
  wire v90f4fb;
  wire v93e0e6;
  wire v90ef0d;
  wire v89b1a4;
  wire v90e978;
  wire v906255;
  wire v90855a;
  wire v93fc0a;
  wire v93f119;
  wire v93f1b4;
  wire v93e228;
  wire v907e7e;
  wire v93fd12;
  wire v93fa7e;
  wire v910527;
  wire v93e3cf;
  wire v89f983;
  wire v93f9af;
  wire v90fb76;
  wire v908a34;
  wire v904f52;
  wire v93f1c8;
  wire v9131c9;
  wire v904e16;
  wire v9062b5;
  wire v909637;
  wire v906623;
  wire v9045f4;
  wire v9076a7;
  wire v908f27;
  wire v87c21e;
  wire v9049d0;
  wire v93fdeb;
  wire v90a6d6;
  wire v93fdc4;
  wire v93fce8;
  wire v93fd48;
  wire v9096f0;
  wire v911f1f;
  wire v90d52b;
  wire v90ee51;
  wire v93003e;
  wire v90a63a;
  wire v90a2b5;
  wire v93f927;
  wire v913332;
  wire v93dfc0;
  wire v8b9e82;
  wire v90fc92;
  wire v906ae9;
  wire v93fcc9;
  wire v863a47;
  wire v93f910;
  wire v93f6ea;
  wire v90f83a;
  wire v90534f;
  wire v90810f;
  wire v8d37c1;
  wire v904725;
  wire v93f111;
  wire v9051bb;
  wire v9058f3;
  wire v86c2d0;
  wire v93e295;
  wire v93e8de;
  wire v913619;
  wire v86e433;
  wire v9132e5;
  wire v89c5e3;
  wire v908eba;
  wire v9085fc;
  wire v906c66;
  wire v90ae9a;
  wire v9046a6;
  wire v93f738;
  wire v8a8b0a;
  wire v90f624;
  wire v8a8fb1;
  wire v93fce7;
  wire v911102;
  wire v886f59;
  wire v93e402;
  wire v90deff;
  wire v8b98be;
  wire v93f7ad;
  wire v93fc7d;
  wire v90ee6d;
  wire v93ec50;
  wire v9082a3;
  wire v93fdfb;
  wire v912679;
  wire v93fdde;
  wire v93f762;
  wire v908e01;
  wire v93e933;
  wire v859635;
  wire v93ee4b;
  wire v8a8fdd;
  wire v905461;
  wire v93e9b9;
  wire v93fa17;
  wire v9096ae;
  wire v93fd25;
  wire v90db6b;
  wire v93fc5d;
  wire v88c601;
  wire v93f908;
  wire v93fb31;
  wire v93fe20;
  wire v9082e4;
  wire v905396;
  wire v904b58;
  wire v9098ba;
  wire v904663;
  wire v93fce2;
  wire v889a9e;
  wire v903fe9;
  wire v93fd23;
  wire v90e945;
  wire v85ea5f;
  wire v93e404;
  wire v93f7b7;
  wire v93e14f;
  wire v93f0a3;
  wire v905c01;
  wire v90d2b7;
  wire v906256;
  wire v93f68a;
  wire v93f541;
  wire v93f690;
  wire v9046f9;
  wire v90dc9c;
  wire v9133ba;
  wire v8f2234;
  wire v905df9;
  wire v89f844;
  wire v93ee84;
  wire v906c6e;
  wire v909078;
  wire v93db3f;
  wire v872e32;
  wire v908834;
  wire v909ca5;
  wire v90932e;
  wire v93e650;
  wire v909080;
  wire v93fbd8;
  wire v908797;
  wire v90e6f1;
  wire v93fa44;
  wire v906cc5;
  wire v90d662;
  wire v90eece;
  wire v90a149;
  wire v8633c3;
  wire v8ee17f;
  wire v906cd3;
  wire v906913;
  wire v90748b;
  wire v9126bb;
  wire v90798e;
  wire v9132ed;
  wire v90729a;
  wire v93ef46;
  wire v93fb0f;
  wire v93fc19;
  wire v909297;
  wire v90d7e7;
  wire v91218a;
  wire v85f258;
  wire v90460c;
  wire v93f796;
  wire v90ae72;
  wire v93ee1b;
  wire v908636;
  wire v912d1c;
  wire v904430;
  wire v90eda0;
  wire v93f6df;
  wire v93e9e3;
  wire v90decf;
  wire v93f652;
  wire v93f9d5;
  wire v93fbc2;
  wire v90fe5c;
  wire v88c832;
  wire v91071e;
  wire v93f922;
  wire v904520;
  wire v90ad02;
  wire v90a181;
  wire v90441c;
  wire v8b9d27;
  wire v90e526;
  wire v93e37e;
  wire v93f805;
  wire v93e97c;
  wire v90d1ca;
  wire v90759b;
  wire v93f155;
  wire v93fb83;
  wire v87a1b7;
  wire v93fd6f;
  wire v90ed3d;
  wire v908df7;
  wire v93f32b;
  wire v910d10;
  wire v904296;
  wire v9120f4;
  wire v93f821;
  wire v89f93b;
  wire v85eaf1;
  wire v93f5e9;
  wire v9098ab;
  wire v9086b7;
  wire v90a216;
  wire v90e4ec;
  wire v93f61e;
  wire v9089bf;
  wire v9097b1;
  wire v87c55f;
  wire v90598f;
  wire v91a6e7;
  wire v87bf0e;
  wire v93fcb9;
  wire v908e73;
  wire v9099e8;
  wire v85f243;
  wire v93f80d;
  wire v8f3874;
  wire v93f282;
  wire v87c558;
  wire v9052f2;
  wire v9097db;
  wire v904025;
  wire v9096a3;
  wire v909823;
  wire v9090d6;
  wire v93e269;
  wire v93fa72;
  wire v909cb1;
  wire v89f90b;
  wire v904ba7;
  wire v93fe48;
  wire v8a8f89;
  wire v93fb27;
  wire v8b9c2c;
  wire v91016c;
  wire v90ff47;
  wire v90432c;
  wire v93debb;
  wire v85eac9;
  wire v903d0b;
  wire v908f85;
  wire v909c72;
  wire v93fcf9;
  wire v93e6fe;
  wire v90e546;
  wire v905136;
  wire v93f1cf;
  wire v90ec05;
  wire v8ee1cd;
  wire v93f727;
  wire v90cfda;
  wire v910d56;
  wire v93e168;
  wire v93fd5c;
  wire v91162e;
  wire v90e251;
  wire v9096fd;
  wire v9124c5;
  wire v90f7d3;
  wire v93fb61;
  wire v910d70;
  wire v93ec4d;
  wire v904ae0;
  wire v91305d;
  wire v93fcc5;
  wire v90ae5a;
  wire v93f7b8;
  wire v93f7f0;
  wire v93e9e5;
  wire v93fd77;
  wire v909928;
  wire v90ee37;
  wire v9043f4;
  wire v91a757;
  wire v9043c7;
  wire v912673;
  wire v90fbfe;
  wire v911185;
  wire v93f928;
  wire v90604e;
  wire v906bf5;
  wire v910117;
  wire v93daaf;
  wire v907a13;
  wire v903e62;
  wire v89b100;
  wire v93f535;
  wire v93f6a7;
  wire v93f906;
  wire v93ed96;
  wire v910056;
  wire v90d217;
  wire v90f07f;
  wire v9097c6;
  wire v90a1db;
  wire v8ee1a7;
  wire v93f2a8;
  wire v93f8c1;
  wire v90cbf6;
  wire v8d37bd;
  wire v9090d1;
  wire v8b9c2b;
  wire v907c8c;
  wire v93fd21;
  wire v9044b8;
  wire v909705;
  wire v905537;
  wire v904995;
  wire v93e684;
  wire v904654;
  wire v908f32;
  wire v904313;
  wire v93fdc6;
  wire v90f8c9;
  wire v90ea8a;
  wire v911c50;
  wire v93fc9a;
  wire v93f88f;
  wire v912124;
  wire v908816;
  wire v8b9d49;
  wire v90a2b8;
  wire v93f82e;
  wire v93e385;
  wire v904df8;
  wire v93f74f;
  wire v8f22a5;
  wire v93f8a0;
  wire v91003a;
  wire v93ecb6;
  wire v8ee181;
  wire v93fb37;
  wire v87cb9e;
  wire v90d4ff;
  wire v909e7f;
  wire v93fa81;
  wire v93ec26;
  wire v909d18;
  wire v93fb2e;
  wire v93f731;
  wire v8b9e6b;
  wire v93fc06;
  wire v93fad7;
  wire v93f936;
  wire v85eacb;
  wire v904757;
  wire v9054c9;
  wire v93fb1a;
  wire v904765;
  wire v93f6b8;
  wire v87a979;
  wire v90a798;
  wire v912643;
  wire v90cbf7;
  wire v910cda;
  wire v93f28b;
  wire v93f811;
  wire v904221;
  wire v911815;
  wire v913342;
  wire v8810ad;
  wire v93fb6e;
  wire v93e0fb;
  wire v92fff5;
  wire v90744a;
  wire v909366;
  wire v90d78b;
  wire v93f588;
  wire v93fa08;
  wire v93ebf5;
  wire v906d77;
  wire v93f646;
  wire v863450;
  wire v9109e6;
  wire v9045b2;
  wire v905838;
  wire v90e2e7;
  wire v8b9c52;
  wire v9051da;
  wire v90656f;
  wire v904590;
  wire v93fc7e;
  wire v93fcd9;
  wire v93e535;
  wire v9043e5;
  wire v93f76e;
  wire v8a8f6f;
  wire v90cc57;
  wire v93fcda;
  wire v906315;
  wire v9082ba;
  wire v9114c0;
  wire v93f7fd;
  wire v91a99a;
  wire v93fd1e;
  wire v86d7d1;
  wire v90f1cb;
  wire v90e38d;
  wire v93ef01;
  wire v91026f;
  wire v907383;
  wire v90a8ac;
  wire v93fd78;
  wire v9135b9;
  wire v93dab8;
  wire v90d718;
  wire v8f22ee;
  wire v93f8c6;
  wire v93ee38;
  wire v93f989;
  wire v863346;
  wire v90481b;
  wire v93fa73;
  wire v90d5bd;
  wire v910cee;
  wire v93fd55;
  wire v9118f0;
  wire v93fcf2;
  wire v8728ef;
  wire v93fc07;
  wire v93f86a;
  wire v93ece6;
  wire v85cca5;
  wire v91a6f1;
  wire v87e0d8;
  wire v92ffd3;
  wire v93fd3e;
  wire v93f29c;
  wire v93fc26;
  wire v9070f7;
  wire v911db6;
  wire v93fe29;
  wire v90a2b9;
  wire v93f7b1;
  wire v93fd1f;
  wire v905dd8;
  wire v91146e;
  wire v912481;
  wire v90eed7;
  wire v93de80;
  wire v90a314;
  wire v90a07e;
  wire v89f852;
  wire v909ab9;
  wire v9126b6;
  wire v8f3849;
  wire v904434;
  wire v93eb9e;
  wire v93fd33;
  wire v85f2b9;
  wire v90a0b5;
  wire v93f77c;
  wire v93fbaa;
  wire v89b116;
  wire v93e2c2;
  wire v90faaf;
  wire v9067c1;
  wire v906c48;
  wire v8b9c3f;
  wire v90df22;
  wire v93e549;
  wire v93fcea;
  wire v90809d;
  wire v90496b;
  wire v93f9ad;
  wire v88b848;
  wire v910b21;
  wire v93fba3;
  wire v89fe24;
  wire v8b989a;
  wire v8880f2;
  wire v90d731;
  wire v907a1b;
  wire v93fdbe;
  wire v93f9ff;
  wire v873a26;
  wire v913079;
  wire v8b98bd;
  wire v911760;
  wire v904e53;
  wire v93fcf4;
  wire v9133ad;
  wire v93fa56;
  wire v908083;
  wire v905252;
  wire v93f687;
  wire v89f984;
  wire v93f665;
  wire v910bd7;
  wire v8f3853;
  wire v89e0b4;
  wire v905425;
  wire v93fdf0;
  wire v906534;
  wire v90789d;
  wire v930106;
  wire v93fded;
  wire v9090c9;
  wire v93fdba;
  wire v908a98;
  wire v93db10;
  wire v93fd40;
  wire v93f92e;
  wire v8848d6;
  wire v93fda7;
  wire v908096;
  wire v909666;
  wire v90a0e8;
  wire v905d73;
  wire v906461;
  wire v93e68f;
  wire v9045df;
  wire v89f905;
  wire v93fc28;
  wire v93fc1a;
  wire v90690e;
  wire v93f681;
  wire v93f9a4;
  wire v905381;
  wire v906ad1;
  wire v903aff;
  wire v90f79b;
  wire v910495;
  wire v911ec2;
  wire v905285;
  wire v909ea8;
  wire v88036c;
  wire v85f268;
  wire v90a098;
  wire v908a2f;
  wire v9134c0;
  wire v9088de;
  wire v8f22e0;
  wire v93e7c2;
  wire v93fb0a;
  wire v93f005;
  wire v9077be;
  wire v90f8e7;
  wire v93fbff;
  wire v909cee;
  wire v90a1f7;
  wire v93f8e4;
  wire v904e47;
  wire v90d442;
  wire v909cf3;
  wire v93f64f;
  wire v93fbbe;
  wire v93fdaf;
  wire v93e9ce;
  wire v93faeb;
  wire v93fae6;
  wire v8b4977;
  wire v907898;
  wire v93e78b;
  wire v906c8c;
  wire v93e337;
  wire v907add;
  wire v906717;
  wire v93edc8;
  wire v89f82d;
  wire v93fa99;
  wire v93fe00;
  wire v8b9efa;
  wire v8633ef;
  wire v906cf5;
  wire v906495;
  wire v911bc2;
  wire v90cc41;
  wire v903c09;
  wire v93f92f;
  wire v903d01;
  wire v9064b4;
  wire v87c503;
  wire v93f6e2;
  wire v87c4c5;
  wire v903c80;
  wire v8b9d28;
  wire v93ec24;
  wire v93f699;
  wire v90f304;
  wire v8b9d84;
  wire v90f62b;
  wire v906038;
  wire v85eaa2;
  wire v9041a7;
  wire v93fd49;
  wire v93f9da;
  wire v909001;
  wire v903b4e;
  wire v90517f;
  wire v93f781;
  wire v912fb2;
  wire v93f8b2;
  wire v907664;
  wire v863478;
  wire v844fb5;
  wire v905972;
  wire v903c65;
  wire v93faa4;
  wire v905ed9;
  wire v90eea7;
  wire v93eed6;
  wire v93fe07;
  wire v8b49ad;
  wire v90515d;
  wire v93e819;
  wire v93f8e0;
  wire v93e6af;
  wire v903fef;
  wire v871b18;
  wire v911c73;
  wire v93f739;
  wire v93e024;
  wire v90d880;
  wire v90443a;
  wire v93e2e6;
  wire v910e17;
  wire v90d21a;
  wire v8a927b;
  wire v90aa8a;
  wire v907c59;
  wire v870d72;
  wire v903b9c;
  wire v93f98c;
  wire v90ba1a;
  wire v93f6ca;
  wire v93fa1b;
  wire v90fc7f;
  wire v904809;
  wire v904b45;
  wire v8a8f74;
  wire v89e11b;
  wire v906416;
  wire v90a7f2;
  wire v90f787;
  wire v87575e;
  wire v90a9fc;
  wire v8c737b;
  wire v90414b;
  wire v91a9b9;
  wire v90a175;
  wire v904575;
  wire v9050a5;
  wire v9130c9;
  wire v93ed2a;
  wire v87c54e;
  wire v906dea;
  wire v912378;
  wire v907069;
  wire v93eaf0;
  wire v90653d;
  wire v908250;
  wire v90fe91;
  wire v93ee82;
  wire v8a8fac;
  wire v91100a;
  wire v93f8c3;
  wire v93df55;
  wire v90a30e;
  wire v9082fc;
  wire v906042;
  wire v90e36f;
  wire v90a451;
  wire v93fe1e;
  wire v93fca3;
  wire v93f0a9;
  wire v93fa91;
  wire v9124ae;
  wire v93f4e9;
  wire v905487;
  wire v907995;
  wire v9113fb;
  wire v906c2f;
  wire v904aae;
  wire v93f345;
  wire v90a334;
  wire v93006d;
  wire v910e2d;
  wire v93f994;
  wire v93f771;
  wire v90a876;
  wire v93dc15;
  wire v93e68d;
  wire v907e88;
  wire v93f627;
  wire v93fe0d;
  wire v93f745;
  wire v93f2b9;
  wire v9115cb;
  wire v9077c7;
  wire v93fb66;
  wire v90dec9;
  wire v90628f;
  wire v8ee1bc;
  wire v906c20;
  wire v93dbf1;
  wire v91dc98;
  wire v905a9e;
  wire v93f78f;
  wire v90efef;
  wire v909c3b;
  wire v90f391;
  wire v9072b7;
  wire v93f893;
  wire v93fdb3;
  wire v90567a;
  wire v910226;
  wire v87a98d;
  wire v904b7f;
  wire v91038c;
  wire v90512d;
  wire v93e162;
  wire v9075db;
  wire v90dd1f;
  wire v90ad6c;
  wire v905d8b;
  wire v90e133;
  wire v90919c;
  wire v9133ea;
  wire v85ea79;
  wire v904aac;
  wire v93e5bf;
  wire v9044a5;
  wire v87ca8a;
  wire v89f9c3;
  wire v90f38b;
  wire v93e9c7;
  wire v93fade;
  wire v93f92c;
  wire v93eb22;
  wire v906541;
  wire v93f8fa;
  wire v91364c;
  wire v904141;
  wire v90a214;
  wire v93e371;
  wire v908fb8;
  wire v911c82;
  wire v93f6cb;
  wire v909b02;
  wire v90a4bf;
  wire v93fdaa;
  wire v9091dd;
  wire v90f5f8;
  wire v90444f;
  wire v8b9c4f;
  wire v90ad6f;
  wire v91a71d;
  wire v93fdee;
  wire v90787b;
  wire v93fe75;
  wire v90529c;
  wire v904fbf;
  wire v85e94c;
  wire v907da6;
  wire v908546;
  wire v8ee1d1;
  wire v93f875;
  wire v912ec5;
  wire v907edc;
  wire v90f5ff;
  wire v93fd35;
  wire v93fce9;
  wire v90728a;
  wire v93ee39;
  wire v910e84;
  wire v910e66;
  wire v910910;
  wire v90d59c;
  wire v93fc46;
  wire v93f28c;
  wire v9109e5;
  wire v93f743;
  wire v9070d5;
  wire v90515a;
  wire v93ea3e;
  wire v90f7d1;
  wire v93ed29;
  wire v91336c;
  wire v90cee9;
  wire v93f896;
  wire v90fbc8;
  wire v904bdb;
  wire v90d64c;
  wire v93e335;
  wire v93ca43;
  wire v90aa42;
  wire v93fd90;
  wire v906ac6;
  wire v93fa27;
  wire v911013;
  wire v93fd67;
  wire v909458;
  wire v90d9b3;
  wire v93fe39;
  wire v9093d9;
  wire v93fa28;
  wire v8639e7;
  wire v903fa3;
  wire v90ebe8;
  wire v93f444;
  wire v93fd96;
  wire v90991f;
  wire v86d767;
  wire v90d704;
  wire v910db7;
  wire v93fced;
  wire v90dc09;
  wire v91a9b6;
  wire v93fcbd;
  wire v90567c;
  wire v93f899;
  wire v90d81c;
  wire v93efa3;
  wire v93faa6;
  wire v93fd8a;
  wire v93f764;
  wire v908ff3;
  wire v906d80;
  wire v90a2f1;
  wire v90e437;
  wire v93fbc1;
  wire v93e3a5;
  wire v85eadc;
  wire v93fab8;
  wire v93fcf0;
  wire v904af3;
  wire v89e119;
  wire v93f280;
  wire v907840;
  wire v90d4cc;
  wire v906d41;
  wire v906b3d;
  wire v93fb6f;
  wire v905803;
  wire v89f9bc;
  wire v93e86e;
  wire v9096f3;
  wire v93f7f6;
  wire v93fdfa;
  wire v90a3f6;
  wire v9091e3;
  wire v9087d2;
  wire v904d89;
  wire v903c2a;
  wire v93e875;
  wire v90a4f9;
  wire v9042ba;
  wire v909f68;
  wire v909b10;
  wire v93f813;
  wire v93fb7d;
  wire v93e723;
  wire v93fd97;
  wire v93fb4a;
  wire v910543;
  wire v93f284;
  wire v8633bd;
  wire v906f62;
  wire v93f77b;
  wire v90df61;
  wire v93fa5d;
  wire v905dc0;
  wire v93fae3;
  wire v907c85;
  wire v90824e;
  wire v93f050;
  wire v93fbea;
  wire v905d0a;
  wire v909347;
  wire v89f966;
  wire v91093d;
  wire v93fa36;
  wire v9135e9;
  wire v93fc42;
  wire v9100a9;
  wire v93f6ae;
  wire v93f728;
  wire v9111d3;
  wire v90dc2c;
  wire v90e5b9;
  wire v91007d;
  wire v93fc5a;
  wire v90f4f7;
  wire v91aa7d;
  wire v90d8d5;
  wire v8a8faa;
  wire v90f33b;
  wire v93f6de;
  wire v904436;
  wire v909b55;
  wire v90aeb7;
  wire v90d84e;
  wire v90e339;
  wire v908209;
  wire v93f787;
  wire v90e4f2;
  wire v93fa15;
  wire v93e519;
  wire v911b74;
  wire v907e33;
  wire v87ba4e;
  wire v8bbc54;
  wire v90459f;
  wire v91a9de;
  wire v907eaa;
  wire v93f7d7;
  wire v93f979;
  wire v90d370;
  wire v93fd84;
  wire v91267e;
  wire v908867;
  wire v867045;
  wire v93fac5;
  wire v904f1a;
  wire v90efe2;
  wire v910be8;
  wire v905556;
  wire v90df5b;
  wire v9051e8;
  wire v93f792;
  wire v904ec6;
  wire v90e8fd;
  wire v93f6ed;
  wire v908b06;
  wire v903f5a;
  wire v93fb69;
  wire v90ad0b;
  wire v90a629;
  wire v8ee1c7;
  wire v9060c1;
  wire v9101cc;
  wire v9052ef;
  wire v93f293;
  wire v90eaab;
  wire v93f6c6;
  wire v89b1a0;
  wire v909d71;
  wire v93f58c;
  wire v908515;
  wire v913632;
  wire v911944;
  wire v91164f;
  wire v9099ef;
  wire v93dc30;
  wire v911b78;
  wire v8b9dfa;
  wire v908681;
  wire v90484c;
  wire v909c0e;
  wire v8b9f3e;
  wire v93f9c5;
  wire v90a8cd;
  wire v92ffd9;
  wire v93fc3d;
  wire v90fb54;
  wire v93fb8d;
  wire v93f7b3;
  wire v89f9cd;
  wire v8b70a3;
  wire v904fbb;
  wire v93fbfc;
  wire v93fe30;
  wire v908a76;
  wire v904f93;
  wire v93f82a;
  wire v8b99a1;
  wire v9130c5;
  wire v906570;
  wire v905322;
  wire v906d92;
  wire v909eb5;
  wire v8b7122;
  wire v90e9e2;
  wire v9072b4;
  wire v8f3879;
  wire v93f6bc;
  wire v90cc30;
  wire v90eef9;
  wire v93e7d1;
  wire v910c51;
  wire v9050e0;
  wire v93f926;
  wire v905325;
  wire v910919;
  wire v913072;
  wire v90891d;
  wire v9088ff;
  wire v910e69;
  wire v93e5da;
  wire v906a51;
  wire v90f88e;
  wire v93f895;
  wire v93dac8;
  wire v905841;
  wire v93fa86;
  wire v93eaca;
  wire v90a1bc;
  wire v911b48;
  wire v9056bd;
  wire v910469;
  wire v90d0fd;
  wire v90f5fc;
  wire v907684;
  wire v90e856;
  wire v8b9eca;
  wire v905467;
  wire v93efae;
  wire v909a7c;
  wire v89b1a2;
  wire v93f749;
  wire v86ccf1;
  wire v90ad77;
  wire v91aa51;
  wire v9057c1;
  wire v90ef1b;
  wire v93e126;
  wire v93f75b;
  wire v93fb43;
  wire v93db85;
  wire v90854b;
  wire v90da97;
  wire v876439;
  wire v93e77a;
  wire v93f29e;
  wire v913561;
  wire v90f9be;
  wire v9062d9;
  wire v903df5;
  wire v93ec44;
  wire v90805e;
  wire v93f88a;
  wire v905a20;
  wire v85dee0;
  wire v93eece;
  wire v9130af;
  wire v8b9c5f;
  wire v9051c9;
  wire v93f6d5;
  wire v906df6;
  wire v863477;
  wire v93fe68;
  wire v9090dd;
  wire v93fada;
  wire v910f2e;
  wire v9101ae;
  wire v9043b9;
  wire v93f4cd;
  wire v93e10c;
  wire v9045f3;
  wire v89fdce;
  wire v9096f7;
  wire v93fc63;
  wire v93e7d4;
  wire v904088;
  wire v90a5b8;
  wire v93eceb;
  wire v880d7e;
  wire v93fca2;
  wire v93f970;
  wire v8ee1f5;
  wire v90856f;
  wire v91a6d5;
  wire v93e77d;
  wire v93f1aa;
  wire v93f9f0;
  wire v9050e7;
  wire v903ddc;
  wire v8706e4;
  wire v89e042;
  wire v93f9ab;
  wire v9100ff;
  wire v93fc4c;
  wire v8f22ad;
  wire v908000;
  wire v93f7e3;
  wire v910e72;
  wire v90fa41;
  wire v8b98fe;
  wire v86345c;
  wire v93ec81;
  wire v93fcd5;
  wire v93f8b9;
  wire v9054e2;
  wire v93e835;
  wire v9133f0;
  wire v93fd57;
  wire v90548c;
  wire v93ec6f;
  wire v912383;
  wire v909434;
  wire v906c6f;
  wire v93fd5b;
  wire v93f8f7;
  wire v9300cb;
  wire v8b9e3d;
  wire v93e0c5;
  wire v93fd16;
  wire v93fd0e;
  wire v908af7;
  wire v911fe3;
  wire v8857fd;
  wire v93fe56;
  wire v90a91e;
  wire v9070e3;
  wire v91cfc7;
  wire v93f977;
  wire v906d58;
  wire v906f44;
  wire v9083d3;
  wire v93f6c3;
  wire v93dee2;
  wire v89f803;
  wire v90479c;
  wire v90e1d0;
  wire v910c37;
  wire v9059b7;
  wire v907da3;
  wire v93fbe2;
  wire v910473;
  wire v905597;
  wire v90a430;
  wire v93ef13;
  wire v905329;
  wire v9065d3;
  wire v90e44c;
  wire v93fa0d;
  wire v90e88f;
  wire v90a588;
  wire v93da97;
  wire v909bd3;
  wire v93df0a;
  wire v93f85d;
  wire v8b497a;
  wire v90f8d6;
  wire v93fcc1;
  wire v90a604;
  wire v93fe49;
  wire v90ad0a;
  wire v9067d4;
  wire v907c01;
  wire v93fb57;
  wire v863add;
  wire v93effa;
  wire v91091b;
  wire v87010f;
  wire v93fa51;
  wire v90f2f6;
  wire v903c46;
  wire v8b9b9f;
  wire v90ded0;
  wire v93fdd9;
  wire v87283f;
  wire v905194;
  wire v9091fe;
  wire v911973;
  wire v8d3799;
  wire v8a9289;
  wire v93fb95;
  wire v8b9d0f;
  wire v93fa53;
  wire v911941;
  wire v9132eb;
  wire v8f3825;
  wire v9107aa;
  wire v9050d2;
  wire v90fb89;
  wire v906b66;
  wire v90a47f;
  wire v904931;
  wire v93f093;
  wire v9071f0;
  wire v93f6d2;
  wire v907bee;
  wire v910f1b;
  wire v904258;
  wire v91026d;
  wire v90a9c5;
  wire v912d04;
  wire v9070cb;
  wire v90ae53;
  wire v93f9b4;
  wire v90db49;
  wire v93fc0e;
  wire v93fbf9;
  wire v906665;
  wire v8b9c46;
  wire v90ac9e;
  wire v90a4bd;
  wire v93faef;
  wire v93ea75;
  wire v907524;
  wire v90dec8;
  wire v90ae6a;
  wire v93e655;
  wire v93e14a;
  wire v911d61;
  wire v905d37;
  wire v90d698;
  wire v89f92f;
  wire v93f7f9;
  wire v8b5f55;
  wire v93f29d;
  wire v9115e3;
  wire v906492;
  wire v910b91;
  wire v93fab0;
  wire v9058f1;
  wire v93e138;
  wire v93f97f;
  wire v9102cc;
  wire v93f324;
  wire v93f76d;
  wire v93fc4d;
  wire v911005;
  wire v9073c3;
  wire v90aaca;
  wire v90e32f;
  wire v9102f4;
  wire v85eaa5;
  wire v903e8d;
  wire v93fd14;
  wire v93fc8d;
  wire v93e9de;
  wire v870489;
  wire v910d6d;
  wire v907bbb;
  wire v8b9cd2;
  wire v9132d3;
  wire v91097b;
  wire v93fc1f;
  wire v8739eb;
  wire v90a1fa;
  wire v905a5b;
  wire v93f7d6;
  wire v90fae7;
  wire v93fb78;
  wire v87bae8;
  wire v8b9f37;
  wire v913169;
  wire v93f6fb;
  wire v90aa3b;
  wire v904a61;
  wire v90d93b;
  wire v90a75f;
  wire v93fc7b;
  wire v908e8b;
  wire v93eda5;
  wire v93de99;
  wire v93f6eb;
  wire v93f7a9;
  wire v89e121;
  wire v93f223;
  wire v90e3ed;
  wire v904bd4;
  wire v9102aa;
  wire v91143a;
  wire v93fd38;
  wire v907517;
  wire v93f7ca;
  wire v903bfc;
  wire v90d629;
  wire v905397;
  wire v93f680;
  wire v90ecfa;
  wire v910e55;
  wire v93f91c;
  wire v87a203;
  wire v863a97;
  wire v90a5a4;
  wire v907120;
  wire v908fb4;
  wire v908ad9;
  wire v93f986;
  wire v90ede1;
  wire v908ed6;
  wire v9134bc;
  wire v90ef16;
  wire v93e596;
  wire v93e097;
  wire v90d3ff;
  wire v93f89e;
  wire v93fd4e;
  wire v93f6d8;
  wire v91aa3f;
  wire v90dcb3;
  wire v90e2d7;
  wire v93f8f4;
  wire v911f15;
  wire v85de34;
  wire v911ed7;
  wire v93fa4e;
  wire v93f7e8;
  wire v93fbac;
  wire v85ea42;
  wire v90f0a8;
  wire v93f779;
  wire v905de8;
  wire v86f5de;
  wire v906983;
  wire v93fdd1;
  wire v908f73;
  wire v91a73f;
  wire v93f314;
  wire v90cf0e;
  wire v93f202;
  wire v906226;
  wire v93fdae;
  wire v93e048;
  wire v909e90;
  wire v89e108;
  wire v90844d;
  wire v910101;
  wire v907299;
  wire v908edf;
  wire v93fb91;
  wire v93f80a;
  wire v93fe47;
  wire v903d12;
  wire v90e76a;
  wire v87b42f;
  wire v90e8bf;
  wire v91137e;
  wire v908138;
  wire v90468d;
  wire v90f1b8;
  wire v908bf7;
  wire v93fcad;
  wire v90d5a9;
  wire v93faff;
  wire v90fd1c;
  wire v908a4f;
  wire v907c71;
  wire v87c534;
  wire v90441e;
  wire v93fad5;
  wire v93f6fa;
  wire v90e893;
  wire v906e3d;
  wire v93f852;
  wire v906131;
  wire v93f6b2;
  wire v906e3b;
  wire v90a1fe;
  wire v86ce19;
  wire v907a32;
  wire v9112d1;
  wire v912f3d;
  wire v904671;
  wire v904dcf;
  wire v93fcc0;
  wire v906c10;
  wire v8a8fda;
  wire v90ba2c;
  wire v90a97c;
  wire v87a2ad;
  wire v93fe6a;
  wire v9068b6;
  wire v90827d;
  wire v907472;
  wire v90d0b6;
  wire v90575f;
  wire v9133d2;
  wire v93fe37;
  wire v93e70c;
  wire v8b830b;
  wire v89fdcf;
  wire v8b99bb;
  wire v90501e;
  wire v90a86b;
  wire v93fbb2;
  wire v93fbdd;
  wire v93f80e;
  wire v903e70;
  wire v904d39;
  wire v86fef2;
  wire v9078a1;
  wire v90a20d;
  wire v909cc1;
  wire v93fa4f;
  wire v93fb14;
  wire v8821a1;
  wire v85ea62;
  wire v93f27f;
  wire v93f840;
  wire v910380;
  wire v9094ed;
  wire v90a20e;
  wire v93fcd8;
  wire v93f87e;
  wire v8f37ef;
  wire v90d27b;
  wire v9107ca;
  wire v91137c;
  wire v93f7c4;
  wire v93f6f5;
  wire v93f9b0;
  wire v911edd;
  wire v907e7a;
  wire v93f518;
  wire v8f22ea;
  wire v90a8e9;
  wire v90f9b6;
  wire v911937;
  wire v90d054;
  wire v906fc1;
  wire v90a4e6;
  wire v93fb48;
  wire v91141d;
  wire v9054bc;
  wire v909649;
  wire v90684c;
  wire v93fd7f;
  wire v93fdb4;
  wire v9040a9;
  wire v90eed3;
  wire v906adf;
  wire v909a12;
  wire v907bca;
  wire v9117db;
  wire v905aaa;
  wire v93eba3;
  wire v89c580;
  wire v89fd94;
  wire v90aa3c;
  wire v93fd1c;
  wire v90ff07;
  wire v93fad0;
  wire v886fce;
  wire v93f8ff;
  wire v93fa46;
  wire v90e25e;
  wire v90824f;
  wire v93f6c9;
  wire v905b62;
  wire v93fc18;
  wire v93fc0b;
  wire v9119f8;
  wire v9081aa;
  wire v907e8f;
  wire v86d690;
  wire v93df15;
  wire v9099f2;
  wire v9061b3;
  wire v90acfe;
  wire v904603;
  wire v905170;
  wire v93f8a9;
  wire v90ad3d;
  wire v9087b7;
  wire v909d1c;
  wire v93f73a;
  wire v8b9f34;
  wire v87de8d;
  wire v87c547;
  wire v93fa8d;
  wire v93fa75;
  wire v905540;
  wire v912173;
  wire v93fa47;
  wire v93db04;
  wire v89f9e4;
  wire v844fbf;
  wire v906ce1;
  wire v911a33;
  wire v844fa3;
  wire v912fad;
  wire v93f037;
  wire v93f894;
  wire v93f720;
  wire v93f66b;
  wire v8807b1;
  wire v910b4b;
  wire v904fd2;
  wire v908106;
  wire v93f8b4;
  wire v93e137;
  wire v93fb3f;
  wire v90f947;
  wire v90879a;
  wire v910b05;
  wire v905618;
  wire v93f31f;
  wire v93fa4c;
  wire v91a76f;
  wire v906b5f;
  wire v8d195d;
  wire v9071ed;
  wire v8d37d4;
  wire v8f22d1;
  wire v88e67b;
  wire v93f701;
  wire v9115a7;
  wire v88b606;
  wire v85e142;
  wire v93fb58;
  wire v93001e;
  wire v90425a;
  wire v910cbf;
  wire v93eade;
  wire v908ae5;
  wire v9049b2;
  wire v93e853;
  wire v909367;
  wire v93fc6d;
  wire v90f5bd;
  wire v93f098;
  wire v91051a;
  wire v907683;
  wire v93f5ff;
  wire v8b49cc;
  wire v93fa29;
  wire v907abc;
  wire v93f92a;
  wire v9112e1;
  wire v907e73;
  wire v908436;
  wire v910fe2;
  wire v93fdf1;
  wire v93f6a2;
  wire v93dc08;
  wire v904847;
  wire v90736f;
  wire v93e4c1;
  wire v9086d9;
  wire v90fb82;
  wire v93fce3;
  wire v93e975;
  wire v93f490;
  wire v90a96f;
  wire v90ed6e;
  wire v93fe5a;
  wire v90e988;
  wire v905f24;
  wire v89fd8d;
  wire v93fad3;
  wire v93e301;
  wire v93f8b8;
  wire v905aa1;
  wire v906d4c;
  wire v905e43;
  wire v93e136;
  wire v93e60f;
  wire v93dee0;
  wire v93f6fe;
  wire v9045bb;
  wire v93fbf3;
  wire v93eb43;
  wire v93e886;
  wire v9110a7;
  wire v93fa05;
  wire v90aca4;
  wire v90f9ed;
  wire v911a89;
  wire v87c566;
  wire v91aa43;
  wire v93fde9;
  wire v8f2274;
  wire v93fd1a;
  wire v911880;
  wire v910403;
  wire v8ee172;
  wire v90980a;
  wire v93fae2;
  wire v93e6c2;
  wire v909365;
  wire v89f894;
  wire v93fc97;
  wire v91359a;
  wire v89f796;
  wire v904b9e;
  wire v904ba3;
  wire v90e333;
  wire v90539a;
  wire v93faf4;
  wire v90d5c3;
  wire v93fe61;
  wire v93fe72;
  wire v93fe1f;
  wire v90456e;
  wire v903b7b;
  wire v93fac6;
  wire v9113b2;
  wire v903c6e;
  wire v907633;
  wire v93fc98;
  wire v90a36a;
  wire v9117de;
  wire v906209;
  wire v9105f4;
  wire v93f73c;
  wire v93fd00;
  wire v93f6f4;
  wire v9076cf;
  wire v93e2a0;
  wire v93e4b4;
  wire v91214b;
  wire v904da6;
  wire v904abd;
  wire v93fd01;
  wire v93f8ec;
  wire v93f73e;
  wire v90a49d;
  wire v908ed2;
  wire v93e193;
  wire v91aa2a;
  wire v904b09;
  wire v93f9d7;
  wire v87ca3a;
  wire v85f2b0;
  wire v93fe21;
  wire v90edd1;
  wire v93fd44;
  wire v90a074;
  wire v93e852;
  wire v8b6009;
  wire v8660c5;
  wire v8b4a3a;
  wire v844fb1;
  wire v909c45;
  wire v93fd32;
  wire v908f48;
  wire v93f15e;
  wire v863b25;
  wire v93ecc4;
  wire v93fd7a;
  wire v903cf9;
  wire v9056d9;
  wire v93fd8d;
  wire v93fcf3;
  wire v9124cb;
  wire v906b57;
  wire v909187;
  wire v904de5;
  wire v908e7c;
  wire v911383;
  wire v93f72f;
  wire v90ecba;
  wire v906c91;
  wire v911b4e;
  wire v8b9b94;
  wire v93fb36;
  wire v93fe3d;
  wire v93f21c;
  wire v93fd79;
  wire v87c4fa;
  wire v93f085;
  wire v903b70;
  wire v910958;
  wire v93fba8;
  wire v91a9b7;
  wire v905511;
  wire v93fa95;
  wire v906d53;
  wire v93f91d;
  wire v9097da;
  wire v90aa5e;
  wire v90df59;
  wire v93f90a;
  wire v8f60f9;
  wire v93fbe4;
  wire v93f136;
  wire v904ee9;
  wire v8b9b71;
  wire v93faab;
  wire v909a7b;
  wire v93e03a;
  wire v93fc4a;
  wire v89f79e;
  wire v904f14;
  wire v93fe64;
  wire v93fbb7;
  wire v908cf4;
  wire v912f40;
  wire v90d8d8;
  wire v93fc27;
  wire v904ecc;
  wire v93f990;
  wire v93fbb8;
  wire v880314;
  wire v93f6e9;
  wire v93f960;
  wire v9107e7;
  wire v93ec72;
  wire v9114c9;
  wire v90671f;
  wire v910ff7;
  wire v90e6f5;
  wire v93fc9d;
  wire v870dd6;
  wire v90edca;
  wire v908e75;
  wire v93fdf3;
  wire v9083c5;
  wire v93f5db;
  wire v93f912;
  wire v910237;
  wire v904b8c;
  wire v93ec47;
  wire v93f074;
  wire v904abe;
  wire v90ea47;
  wire v903fc8;
  wire v93f9e3;
  wire v90fa18;
  wire v910d28;
  wire v93fc67;
  wire v90e373;
  wire v90e1c3;
  wire v904ebe;
  wire v93fbaf;
  wire v87e7f5;
  wire v93fd63;
  wire v904753;
  wire v913449;
  wire v90d727;
  wire v8b9e71;
  wire v90f9fc;
  wire v909a21;
  wire v93db12;
  wire v93fb2b;
  wire v93fe17;
  wire v93fc4e;
  wire v8b9d1b;
  wire v93fbb3;
  wire v93fa9d;
  wire v910cf2;
  wire v86f729;
  wire v93f854;
  wire v904c38;
  wire v90f88a;
  wire v93f782;
  wire v90cc7a;
  wire v910ca7;
  wire v93df10;
  wire v93ec28;
  wire v90ee4b;
  wire v909d9c;
  wire v906638;
  wire v93edbf;
  wire v93dc87;
  wire v903c1f;
  wire v913a64;
  wire v9104bd;
  wire v93e31b;
  wire v9117e2;
  wire v90d057;
  wire v89e0d5;
  wire v93f9ef;
  wire v93fb1b;
  wire v88932d;
  wire v908d10;
  wire v93dbe9;
  wire v88dbe7;
  wire v90a4da;
  wire v90cbfd;
  wire v93fcf1;
  wire v9045e6;
  wire v8b9ebe;
  wire v9132d2;
  wire v8f22ce;
  wire v9119f9;
  wire v90edf6;
  wire v93fd86;
  wire v93f291;
  wire v905d9c;
  wire v903afe;
  wire v93f5f6;
  wire v90a563;
  wire v9096f1;
  wire v87a28e;
  wire v91143f;
  wire v93fcc2;
  wire v90ae1b;
  wire v904878;
  wire v93fd18;
  wire v90e925;
  wire v8b9d4b;
  wire v9104f8;
  wire v90f0bd;
  wire v9057c9;
  wire v904a80;
  wire v90a2bd;
  wire v9133dc;
  wire v93fccd;
  wire v907559;
  wire v910915;
  wire v904dc1;
  wire v90dedf;
  wire v90faf6;
  wire v91a796;
  wire v93f95a;
  wire v93fb11;
  wire v90e841;
  wire v93f855;
  wire v93f735;
  wire v9043c2;
  wire v85acd3;
  wire v905460;
  wire v93fc53;
  wire v90dd67;
  wire v9133ec;
  wire v9075e7;
  wire v90d5d1;
  wire v904f22;
  wire v91268b;
  wire v910c3a;
  wire v9107c7;
  wire v93e156;
  wire v910f4d;
  wire v93fb0b;
  wire v863363;
  wire v93f533;
  wire v93f965;
  wire v906af3;
  wire v93e33e;
  wire v93f6e5;
  wire v85ea76;
  wire v911724;
  wire v90966d;
  wire v904b04;
  wire v90944f;
  wire v909995;
  wire v93edf1;
  wire v90e1cf;
  wire v91107f;
  wire v90477e;
  wire v904eea;
  wire v8b9ce2;
  wire v93fd4f;
  wire v90eea6;
  wire v9054a8;
  wire v93f7b9;
  wire v93f736;
  wire v8f22ca;
  wire v90e027;
  wire v93fba0;
  wire v9049bf;
  wire v8f22e3;
  wire v903cda;
  wire v904bbf;
  wire v884fc2;
  wire v90f478;
  wire v93faae;
  wire v8b9b56;
  wire v90e958;
  wire v93fc76;
  wire v93fd74;
  wire v93fcc6;
  wire v93f65b;
  wire v93f919;
  wire v93f9b8;
  wire v93f8d4;
  wire v907494;
  wire v93fa64;
  wire v90e7e2;
  wire v908ef9;
  wire v8b9ec2;
  wire v89e12f;
  wire v844fb9;
  wire v93f878;
  wire v93f2da;
  wire v8b496d;
  wire v906b43;
  wire v9046de;
  wire v93fb86;
  wire v905847;
  wire v90fbad;
  wire v90a59e;
  wire v93e391;
  wire v93fa7c;
  wire v90d879;
  wire v8b9dff;
  wire v9114a0;
  wire v904bf3;
  wire v93f7bf;
  wire v91042d;
  wire v93ee87;
  wire v910bf9;
  wire v908410;
  wire v930032;
  wire v93ef30;
  wire v93fe5b;
  wire v9058f4;
  wire v92ffb9;
  wire v906ff5;
  wire v93f7af;
  wire v90762a;
  wire v93fd3c;
  wire v9062b3;
  wire v90765f;
  wire v90ad9a;
  wire v90683e;
  wire v863b34;
  wire v909a26;
  wire v93fa87;
  wire v908533;
  wire v90f78a;
  wire v91003b;
  wire v93ef4c;
  wire v906dd6;
  wire v90729e;
  wire v91080f;
  wire v85f278;
  wire v93fe45;
  wire v90d7e8;
  wire v93f558;
  wire v904b00;
  wire v90d59a;
  wire v9105ed;
  wire v93fe6e;
  wire v93fd2b;
  wire v91305b;
  wire v93e356;
  wire v8c7343;
  wire v9091be;
  wire v909f04;
  wire v93fdf8;
  wire v90d7ce;
  wire v90a2aa;
  wire v93f898;
  wire v93fe66;
  wire v904ede;
  wire v93eb39;
  wire v93fc35;
  wire v9054a2;
  wire v909f63;
  wire v905971;
  wire v93e652;
  wire v9101b8;
  wire v9088a3;
  wire v905186;
  wire v909430;
  wire v93fc22;
  wire v905ffe;
  wire v93fd9a;
  wire v87179f;
  wire v93f7c8;
  wire v90f547;
  wire v93e00f;
  wire v93fb9c;
  wire v93fa35;
  wire v903cd2;
  wire v905cd2;
  wire v85ea9a;
  wire v90657d;
  wire v90e19c;
  wire v930028;
  wire v93fc78;
  wire v85eacf;
  wire v90e6b0;
  wire v90e000;
  wire v8f22a2;
  wire v91071c;
  wire v93fac3;
  wire v904ed4;
  wire v93f3db;
  wire v91aa06;
  wire v90fc6d;
  wire v904b51;
  wire v93fbf8;
  wire v93ec0d;
  wire v904f1b;
  wire v91024c;
  wire v93fdb6;
  wire v93fc69;
  wire v93fe4c;
  wire v911312;
  wire v911318;
  wire v903ec3;
  wire v90d543;
  wire v910b0e;
  wire v93fdcb;
  wire v907f05;
  wire v911417;
  wire v93faa7;
  wire v91247f;
  wire v905835;
  wire v86cda0;
  wire v93f9fa;
  wire v873bc3;
  wire v910d4a;
  wire v90e315;
  wire v8b49bf;
  wire v90fe87;
  wire v90fe55;
  wire v93f092;
  wire v8b9ef8;
  wire v909492;
  wire v93ea4f;
  wire v9068ce;
  wire v911023;
  wire v90962e;
  wire v90a300;
  wire v90d9a0;
  wire v907d03;
  wire v89e0ce;
  wire v90a6ae;
  wire v93f8d0;
  wire v93e77c;
  wire v93f7bd;
  wire v908693;
  wire v88c1f9;
  wire v93f7ec;
  wire v90ed77;
  wire v93fad4;
  wire v93f59b;
  wire v904886;
  wire v93f7a8;
  wire v9080b4;
  wire v93f90d;
  wire v910840;
  wire v910e32;
  wire v908a2c;
  wire v93fc31;
  wire v908f4b;
  wire v93f5cb;
  wire v93fae1;
  wire v913433;
  wire v8b9bd9;
  wire v90a733;
  wire v8b9e96;
  wire v93fbd0;
  wire v9095ec;
  wire v90638b;
  wire v93f045;
  wire v863b37;
  wire v903db9;
  wire v90ea4c;
  wire v93ebe6;
  wire v93e065;
  wire v93fbd3;
  wire v903e08;
  wire v93f8a2;
  wire v93fc01;
  wire v90e083;
  wire v9132d4;
  wire v90521f;
  wire v8a9231;
  wire v93fbd4;
  wire v8b9f21;
  wire v906e15;
  wire v93e450;
  wire v909f36;
  wire v90949f;
  wire v904b41;
  wire v906d63;
  wire v910fd2;
  wire v93f2dc;
  wire v8f382e;
  wire v93fd22;
  wire v9049fd;
  wire v90809b;
  wire v90faf1;
  wire v904c72;
  wire v91a762;
  wire v911365;
  wire v907d8a;
  wire v89b0e5;
  wire v93df9f;
  wire v93dfb4;
  wire v93e72a;
  wire v9092a8;
  wire v9134c4;
  wire v93e855;
  wire v89f97d;
  wire v93e369;
  wire v904ef2;
  wire v907717;
  wire v93fa3f;
  wire v93fdce;
  wire v9041e6;
  wire v904c99;
  wire v9040fb;
  wire v86f60a;
  wire v93f2c6;
  wire v93f7c7;
  wire v909b54;
  wire v9084ae;
  wire v89f84e;
  wire v909119;
  wire v8633ac;
  wire v909918;
  wire v90965e;
  wire v93faf1;
  wire v93fcba;
  wire v93fdbf;
  wire v86dd54;
  wire v90417d;
  wire v93f584;
  wire v93e996;
  wire v903db7;
  wire v9110fe;
  wire v93fa0a;
  wire v909805;
  wire v911a72;
  wire v90f2f4;
  wire v93dbaa;
  wire v905ff9;
  wire v90a08d;
  wire v884dd3;
  wire v909c08;
  wire v93e148;
  wire v9134fe;
  wire v91a9b4;
  wire v90539f;
  wire v93f51c;
  wire v93f8b1;
  wire v8f3826;
  wire v911c11;
  wire v93f12b;
  wire v905f25;
  wire v90dd28;
  wire v9082a5;
  wire v9058d5;
  wire v90546e;
  wire v93fbc7;
  wire v910416;
  wire v93fbee;
  wire v93f4ac;
  wire v907722;
  wire v904303;
  wire v90aeb8;
  wire v93fa2b;
  wire v93f85a;
  wire v93eb70;
  wire v87a20b;
  wire v90ee83;
  wire v93f84d;
  wire v904988;
  wire v8b9c31;
  wire v907a2f;
  wire v86ce77;
  wire v90f161;
  wire v87a242;
  wire v93f5d9;
  wire v93e70e;
  wire v905d92;
  wire v93fb72;
  wire v93fe35;
  wire v908751;
  wire v90828a;
  wire v90f6b4;
  wire v8b9e73;
  wire v93fcb2;
  wire v8f383a;
  wire v8a8f5e;
  wire v905775;
  wire v903c4d;
  wire v93f7ab;
  wire v903d4f;
  wire v93e45c;
  wire v909c15;
  wire v9084f4;
  wire v910d41;
  wire v907b6c;
  wire v907710;
  wire v90ccbd;
  wire v908aae;
  wire v909312;
  wire v93f492;
  wire v93fde2;
  wire v880d77;
  wire v907b01;
  wire v89f927;
  wire v910ffd;
  wire v9086f1;
  wire v93f10b;
  wire v93f02f;
  wire v91262e;
  wire v90edb9;
  wire v93dc2c;
  wire v908176;
  wire v90a9cc;
  wire v906f1e;
  wire v910c20;
  wire v90e62f;
  wire v90d42a;
  wire v90dcfa;
  wire v93e4f9;
  wire v8b9c00;
  wire v90fe7e;
  wire v863418;
  wire v88a51e;
  wire v93f8de;
  wire v904794;
  wire v93dffa;
  wire v90561f;
  wire v93fdb1;
  wire v903b98;
  wire v90fa02;
  wire v90d9b7;
  wire v90a419;
  wire v909dd5;
  wire v93f767;
  wire v910704;
  wire v87a2ae;
  wire v904a90;
  wire v91db5a;
  wire v93fc29;
  wire v930097;
  wire v93fb3a;
  wire v903b7d;
  wire v87a253;
  wire v93f89f;
  wire v9074ce;
  wire v93f768;
  wire v9050cc;
  wire v90a620;
  wire v89f98c;
  wire v93fda1;
  wire v93fe2e;
  wire v9106a7;
  wire v9187aa;
  wire v905038;
  wire v911b43;
  wire v93f8a1;
  wire v913a6f;
  wire v93e773;
  wire v90749b;
  wire v93fbde;
  wire v93f69e;
  wire v904fcd;
  wire v904f5c;
  wire v909415;
  wire v907897;
  wire v93fc5f;
  wire v93e23c;
  wire v90d5c7;
  wire v93e370;
  wire v93fd47;
  wire v93fb5e;
  wire v93f9db;
  wire v906538;
  wire v90408b;
  wire v9071f8;
  wire v85ead8;
  wire v93fa7b;
  wire v93fde6;
  wire v90667f;
  wire v93ebbb;
  wire v93f334;
  wire v903e94;
  wire v863a38;
  wire v93e27a;
  wire v903c83;
  wire v93f7b0;
  wire v93f702;
  wire v8b8638;
  wire v908e7e;
  wire v93fe31;
  wire v89f916;
  wire v93f30c;
  wire v93db1d;
  wire v91aa45;
  wire v9044c6;
  wire v93f8a6;
  wire v90a5ee;
  wire v93e5b8;
  wire v904ab4;
  wire v911cba;
  wire v86333d;
  wire v93f8c5;
  wire v908d2a;
  wire v9095e0;
  wire v906024;
  wire v903d21;
  wire v888002;
  wire v86e831;
  wire v9051f4;
  wire v90dca4;
  wire v93fa6d;
  wire v93f57d;
  wire v904ab2;
  wire v93fd8b;
  wire v89f8bd;
  wire v93fd0d;
  wire v93db7f;
  wire v93fbe1;
  wire v904cde;
  wire v90719c;
  wire v93fb44;
  wire v91232c;
  wire v93e643;
  wire v909be7;
  wire v8b5f5d;
  wire v87a671;
  wire v8b98f4;
  wire v90acc5;
  wire v93efb0;
  wire v93f70a;
  wire v909941;
  wire v9079a8;
  wire v90f0a1;
  wire v93fc49;
  wire v93fab9;
  wire v93f881;
  wire v93e439;
  wire v93e1ed;
  wire v93fdb0;
  wire v904775;
  wire v93fe27;
  wire v87a991;
  wire v93f9d4;
  wire v8b9d35;
  wire v93e4b9;
  wire v930099;
  wire v93f6c1;
  wire v86e625;
  wire v89e0fb;
  wire v87c4ee;
  wire v90ace9;
  wire v93f29a;
  wire v93fcbf;
  wire v9068fc;
  wire v93ea16;
  wire v909c39;
  wire v906d2a;
  wire v90deaa;
  wire v90f36b;
  wire v93ea28;
  wire v8b9c3e;
  wire v93fd4c;
  wire v85ea4f;
  wire v87a25e;
  wire v90faf9;
  wire v912405;
  wire v93f058;
  wire v93e0b5;
  wire v90caed;
  wire v8f223b;
  wire v93fe57;
  wire v91a6f0;
  wire v93fb7a;
  wire v904fb4;
  wire v87ec92;
  wire v93df31;
  wire v93fc17;
  wire v93dc29;
  wire v89f8ef;
  wire v9050ae;
  wire v8b9b88;
  wire v93f7c9;
  wire v93eaa1;
  wire v907799;
  wire v93faed;
  wire v93fcb1;
  wire v93fac4;
  wire v908e4b;
  wire v9112d5;
  wire v93f7de;
  wire v89f8fd;
  wire v904bc1;
  wire v907bfd;
  wire v9043fa;
  wire v93f6bd;
  wire v93eb13;
  wire v910e82;
  wire v90860a;
  wire v909353;
  wire v907634;
  wire v93f203;
  wire v91aa52;
  wire v93fdb7;
  wire v93f7ff;
  wire v904ae4;
  wire v89f948;
  wire v910cc4;
  wire v93fbc0;
  wire v93f7a5;
  wire v93fdc1;
  wire v93f68f;
  wire v93fd93;
  wire v93ec8c;
  wire v89f7e3;
  wire v90d4c9;
  wire v93f82f;
  wire v93fc1d;
  wire v93f959;
  wire v909dec;
  wire v93f75e;
  wire v90e906;
  wire v89e0a6;
  wire v91a799;
  wire v911909;
  wire v9068b7;
  wire v93fa04;
  wire v8f381b;
  wire v904fe6;
  wire v91134b;
  wire v86fe09;
  wire v905dcf;
  wire v90a1fd;
  wire v93fb73;
  wire v93f97e;
  wire v9047eb;
  wire v9079f4;
  wire v90878b;
  wire v90e926;
  wire v90866d;
  wire v9056ac;
  wire v93f870;
  wire v93f8e2;
  wire v9095b9;
  wire v9044c3;
  wire v93fb53;
  wire v907f25;
  wire v910f78;
  wire v90a799;
  wire v90557c;
  wire v8f37f1;
  wire v9068c8;
  wire v93fb9a;
  wire v90dc0a;
  wire v909b01;
  wire v85ea51;
  wire v93f812;
  wire v93fd43;
  wire v93f307;
  wire v904f88;
  wire v93faad;
  wire v90921e;
  wire v93f7bc;
  wire v912178;
  wire v85eb17;
  wire v93e5d4;
  wire v9081ef;
  wire v90ec4b;
  wire v863a7b;
  wire v905355;
  wire v93fda9;
  wire v93fcfe;
  wire v904f0d;
  wire v93f68b;
  wire v9041fc;
  wire v87c52b;
  wire v909b56;
  wire v9086f8;
  wire v93fd52;
  wire v909746;
  wire v9093f3;
  wire v93f97c;
  wire v93f708;
  wire v906c0f;
  wire v9115ae;
  wire v907b54;
  wire v905d7a;
  wire v906fd0;
  wire v90dcca;
  wire v8b9e97;
  wire v91306c;
  wire v90513b;
  wire v9113ea;
  wire v93fbec;
  wire v93fe0e;
  wire v866af4;
  wire v907751;
  wire v93e672;
  wire v906915;
  wire v93f86b;
  wire v8b9eb0;
  wire v92ffc9;
  wire v93f7ce;
  wire v912f42;
  wire v909f7e;
  wire v93e781;
  wire v90d789;
  wire v904b91;
  wire v93dade;
  wire v9095d0;
  wire v8850b3;
  wire v905405;
  wire v87c9f1;
  wire v93e95e;
  wire v90decb;
  wire v8f22bd;
  wire v9061b0;
  wire v93fd0c;
  wire v93fabb;
  wire v911008;
  wire v93f16d;
  wire v93fd07;
  wire v93f795;
  wire v863a2d;
  wire v93fa57;
  wire v93f7e2;
  wire v90f0c4;
  wire v906e30;
  wire v906c0c;
  wire v93fd9b;
  wire v908346;
  wire v903bb1;
  wire v910f5a;
  wire v9067d3;
  wire v903cc5;
  wire v906320;
  wire v910260;
  wire v90dcf0;
  wire v93fb71;
  wire v93f3b9;
  wire v8714f5;
  wire v93fa76;
  wire v8893bb;
  wire v9103bc;
  wire v89f9da;
  wire v93f589;
  wire v906321;
  wire v8ebcf9;
  wire v93fa3c;
  wire v90aa76;
  wire v903c1c;
  wire v90d46a;
  wire v93fbeb;
  wire v93f760;
  wire v93e6f6;
  wire v911b47;
  wire v93fbfa;
  wire v93fce6;
  wire v91066d;
  wire v85eb28;
  wire v904ef7;
  wire v93f9e0;
  wire v8ebd0e;
  wire v8b9d37;
  wire v90e8fa;
  wire v911833;
  wire v93f6f3;
  wire v906b71;
  wire v93fbe8;
  wire v908a3d;
  wire v9057fa;
  wire v90e95b;
  wire v93e903;
  wire v90fa8a;
  wire v904f4d;
  wire v93e41f;
  wire v9134e2;
  wire v8cec7e;
  wire v93e915;
  wire v910dfa;
  wire v908006;
  wire v93fe44;
  wire v905b81;
  wire v93f999;
  wire v93eadd;
  wire v90738c;
  wire v889d4b;
  wire v93f0c0;
  wire v90d1c9;
  wire v93f93c;
  wire v9117e1;
  wire v913067;
  wire v905d63;
  wire v90fc26;
  wire v93f0a6;
  wire v9064e9;
  wire v90d86f;
  wire v9054b6;
  wire v90871b;
  wire v8b9d0e;
  wire v87c517;
  wire v90d5b3;
  wire v904dea;
  wire v904bda;
  wire v93f2fd;
  wire v93fe11;
  wire v909d4d;
  wire v90da38;
  wire v90839e;
  wire v93f70f;
  wire v912172;
  wire v93f844;
  wire v90f164;
  wire v93e9dd;
  wire v930114;
  wire v93fd95;
  wire v910490;
  wire v93ed1c;
  wire v9084d0;
  wire v88d5cd;
  wire v90fb5d;
  wire v90a3da;
  wire v86344b;
  wire v90630d;
  wire v93fa1e;
  wire v90a6ac;
  wire v93e8a1;
  wire v909bbd;
  wire v93fd1d;
  wire v93f83a;
  wire v8b714e;
  wire v930083;
  wire v9044b4;
  wire v884261;
  wire v903cb1;
  wire v93f889;
  wire v93fd89;
  wire v9044c9;
  wire v90d866;
  wire v908fe9;
  wire v910545;
  wire v93e704;
  wire v93f088;
  wire v904ba4;
  wire v906df1;
  wire v93fa7d;
  wire v905408;
  wire v907815;
  wire v93ef5c;
  wire v905a80;
  wire v911edb;
  wire v93ed70;
  wire v93e926;
  wire v909525;
  wire v9081b9;
  wire v907168;
  wire v90a0cb;
  wire v93f3ea;
  wire v93f888;
  wire v905d66;
  wire v90d87f;
  wire v9104aa;
  wire v8f3869;
  wire v9055c0;
  wire v903d60;
  wire v93fabd;
  wire v91a771;
  wire v93f707;
  wire v93dfc7;
  wire v9052ce;
  wire v93fb20;
  wire v93fcb4;
  wire v911a00;
  wire v91a7a3;
  wire v89f7e2;
  wire v90e2dc;
  wire v90f8c2;
  wire v904808;
  wire v91086d;
  wire v93fae4;
  wire v8fe223;
  wire v905ca1;
  wire v90d3cc;
  wire v93f8f8;
  wire v9109ee;
  wire v93fe06;
  wire v93f865;
  wire v911c01;
  wire v91062b;
  wire v93fbd7;
  wire v910081;
  wire v93f8b7;
  wire v90d6fa;
  wire v930016;
  wire v93e829;
  wire v90a557;
  wire v8b9e60;
  wire v904115;
  wire v93ef76;
  wire v90add6;
  wire v93fc6f;
  wire v90f819;
  wire v911b68;
  wire v93fd8e;
  wire v93fdf7;
  wire v905660;
  wire v93fd87;
  wire v909107;
  wire v93fc2a;
  wire v90636e;
  wire v91216e;
  wire v909adc;
  wire v90468f;
  wire v903f58;
  wire v93fd6d;
  wire v93ecd6;
  wire v93f6f0;
  wire v906fec;
  wire v912fa9;
  wire v90d364;
  wire v9085c8;
  wire v93fdd0;
  wire v90cb3d;
  wire v9100bd;
  wire v9088bc;
  wire v90e9f7;
  wire v907091;
  wire v906cc7;
  wire v9079f7;
  wire v9121a6;
  wire v905791;
  wire v90f0a2;
  wire v93f7f7;
  wire v8b9c50;
  wire v91aa44;
  wire v93f7bb;
  wire v907b58;
  wire v90d71a;
  wire v91093c;
  wire v908574;
  wire v909357;
  wire v904da2;
  wire v8b9e40;
  wire v904736;
  wire v93f521;
  wire v9095df;
  wire v93f7e5;
  wire v93fac8;
  wire v88e55e;
  wire v9059ef;
  wire v90a0d7;
  wire v90419d;
  wire v903c40;
  wire v93f790;
  wire v90a602;
  wire v93f7ae;
  wire v93fc86;
  wire v93fc66;
  wire v906fcc;
  wire v904614;
  wire v93fb8a;
  wire v89c59e;
  wire v89f8e5;
  wire v93fa49;
  wire v9106af;
  wire v907b21;
  wire v93fc38;
  wire v9124a6;
  wire v89e0c5;
  wire v909180;
  wire v8f22d0;
  wire v90894d;
  wire v9051ea;
  wire v93e610;
  wire v906e04;
  wire v904132;
  wire v9119fd;
  wire v93fc4f;
  wire v90d250;
  wire v90e772;
  wire v9083cf;
  wire v87c533;
  wire v93fd09;
  wire v93e9cc;
  wire v909058;
  wire v90f5b6;
  wire v9099e3;
  wire v93f9e8;
  wire v87052e;
  wire v90a485;
  wire v90946a;
  wire v903fb2;
  wire v93f96e;
  wire v91cc2d;
  wire v93fdac;
  wire v90fa5e;
  wire v93ec9d;
  wire v93f723;
  wire v93000b;
  wire v9132d6;
  wire v8b4983;
  wire v8b9c55;
  wire v907e36;
  wire v91109f;
  wire v912672;
  wire v9056c5;
  wire v90caeb;
  wire v93f462;
  wire v9115b6;
  wire v93f945;
  wire v872187;
  wire v93fa3b;
  wire v90a44f;
  wire v9097f3;
  wire v8858ac;
  wire v90dc28;
  wire v93eb41;
  wire v93f064;
  wire v86deed;
  wire v930109;
  wire v85e7ba;
  wire v93fa8f;
  wire v905d7e;
  wire v91148d;
  wire v9300c6;
  wire v93f5ae;
  wire v911b9a;
  wire v904901;
  wire v906327;
  wire v93fbb1;
  wire v905312;
  wire v90dc08;
  wire v863ac4;
  wire v907292;
  wire v904d75;
  wire v93fb05;
  wire v908ee8;
  wire v93fafe;
  wire v93ecb0;
  wire v90a884;
  wire v93fdb8;
  wire v918724;
  wire v90eab9;
  wire v8b9e9f;
  wire v93fe38;
  wire v93fd85;
  wire v871483;
  wire v9060e9;
  wire v9077f6;
  wire v909d2b;
  wire v90ad48;
  wire v905b5d;
  wire v93fb00;
  wire v9091c7;
  wire v90ee74;
  wire v93ea5d;
  wire v93fac9;
  wire v93f83f;
  wire v8a8fa0;
  wire v93f33e;
  wire v909b74;
  wire v93e1c0;
  wire v91230c;
  wire v9045f0;
  wire v863aee;
  wire v93fa93;
  wire v910937;
  wire v93f82d;
  wire v93fd73;
  wire v91a6e9;
  wire v910642;
  wire v90fc5f;
  wire v85eaed;
  wire v91aa76;
  wire v93fb8f;
  wire v93fb8c;
  wire v9115ab;
  wire v907ad8;
  wire v93fb6c;
  wire v91150c;
  wire v8b9d5d;
  wire v90a7ea;
  wire v8d37d8;
  wire v93ec67;
  wire v9098a3;
  wire v913265;
  wire v906b07;
  wire v904e13;
  wire v90cbea;
  wire v93f892;
  wire v8d37be;
  wire v90ea21;
  wire v8633df;
  wire v910221;
  wire v93f0bf;
  wire v9048d7;
  wire v87c537;
  wire v90712c;
  wire v93fc34;
  wire v93f511;
  wire v90d9fd;
  wire v92ffda;
  wire v90a902;
  wire v91194f;
  wire v907b65;
  wire v90f3e4;
  wire v93f87a;
  wire v903fb0;
  wire v905665;
  wire v870615;
  wire v87a21e;
  wire v93fda0;
  wire v903c43;
  wire v93fd2c;
  wire v908322;
  wire v90ad69;
  wire v863aa0;
  wire v8b9e6e;
  wire v9080a8;
  wire v93e5e5;
  wire v912f16;
  wire v910062;
  wire v93fccc;
  wire v91071b;
  wire v88946f;
  wire v93f7dc;
  wire v90cfa8;
  wire v91082c;
  wire v93fce0;
  wire v93ef2e;
  wire v93f68c;
  wire v93f02c;
  wire v90a20a;
  wire v93f52d;
  wire v905619;
  wire v8a9205;
  wire v90e172;
  wire v90a207;
  wire v93fcf7;
  wire v906657;
  wire v903b1a;
  wire v93fa22;
  wire v88403f;
  wire v93e32d;
  wire v911150;
  wire v9078f8;
  wire v90494f;
  wire v93f5d7;
  wire v93fc6c;
  wire v904852;
  wire v904bc0;
  wire v909d90;
  wire v9089ef;
  wire v906ce5;
  wire v89f830;
  wire v8d373a;
  wire v93f26c;
  wire v93fb4f;
  wire v8f383c;
  wire v907a4d;
  wire v93faac;
  wire v90a5c0;
  wire v905ac3;
  wire v93e69c;
  wire v93f9f7;
  wire v908545;
  wire v91336b;
  wire v85eb2b;
  wire v87ca35;
  wire v93dfc2;
  wire v871df8;
  wire v90e94e;
  wire v90cbec;
  wire v93f73d;
  wire v9118a3;
  wire v93f04f;
  wire v93f8a5;
  wire v90441d;
  wire v93fe55;
  wire v90752a;
  wire v9045fa;
  wire v90f1ab;
  wire v93fbfe;
  wire v909289;
  wire v910ea0;
  wire v9099a1;
  wire v912477;
  wire v93f78c;
  wire v90f66c;
  wire v93fe0c;
  wire v90d999;
  wire v93f9a1;
  wire v89e122;
  wire v93e05f;
  wire v906c67;
  wire v910fda;
  wire v907d8b;
  wire v90998d;
  wire v863a03;
  wire v90fb4b;
  wire v91192b;
  wire v93e919;
  wire v8b9f23;
  wire v93fe4b;
  wire v93f801;
  wire v8b9c87;
  wire v9054bd;
  wire v91132f;
  wire v89fe59;
  wire v93eff8;
  wire v87a993;
  wire v905f54;
  wire v908ae0;
  wire v93fac0;
  wire v90d0b8;
  wire v93fb82;
  wire v90f7d6;
  wire v93fe52;
  wire v90a33b;
  wire v90e341;
  wire v904a0b;
  wire v93fcbc;
  wire v93fd04;
  wire v9062ae;
  wire v85ef3a;
  wire v903db4;
  wire v93fd6c;
  wire v91e95f;
  wire v904357;
  wire v90950c;
  wire v8b98f1;
  wire v905539;
  wire v93f110;
  wire v906cc8;
  wire v93deab;
  wire v93fb3b;
  wire v89e097;
  wire v91a6d1;
  wire v93f6cc;
  wire v90efea;
  wire v90423b;
  wire v90451f;
  wire v9073c5;
  wire v93fa4b;
  wire v90667d;
  wire v863afc;
  wire v9109f4;
  wire v911552;
  wire v913362;
  wire v8b9ee1;
  wire v90f575;
  wire v9099fa;
  wire v90eef5;
  wire v93eec4;
  wire v93f6fd;
  wire v90ebcd;
  wire v91aa12;
  wire v93006b;
  wire v911b83;
  wire v93f8d2;
  wire v93f7d2;
  wire v90648f;
  wire v910fd8;
  wire v93f678;
  wire v90738d;
  wire v903fac;
  wire v90d6ef;
  wire v91267b;
  wire v88aff7;
  wire v9059b8;
  wire v904a70;
  wire v86e277;
  wire v93f8af;
  wire v90ec5d;
  wire v90fca6;
  wire v90808b;
  wire v913428;
  wire v907c76;
  wire v90d32d;
  wire v93fc93;
  wire v8b9cc5;
  wire v93fc45;
  wire v90e770;
  wire v93ed6a;
  wire v93f869;
  wire v87c4d9;
  wire v90ee63;
  wire v87c9b1;
  wire v9063de;
  wire v913a2b;
  wire v91a6f7;
  wire v90508f;
  wire v93f470;
  wire v93f8ae;
  wire v90cbcc;
  wire v93e470;
  wire v93fa25;
  wire v89f97f;
  wire v93fb2f;
  wire v90723b;
  wire v8b9ce5;
  wire v90f7e4;
  wire v903b83;
  wire v93fdf6;
  wire v93fe5c;
  wire v90ebde;
  wire v863b1a;
  wire v93f664;
  wire v87b2ea;
  wire v90986f;
  wire v8b4981;
  wire v90dab9;
  wire v903eef;
  wire v93fe71;
  wire v93e188;
  wire v91325d;
  wire v93f7a2;
  wire v90914c;
  wire v9133d9;
  wire v906d2b;
  wire v91325f;
  wire v93f962;
  wire v93e6e0;
  wire v90861d;
  wire v9040cd;
  wire v8b49dc;
  wire v90f2f9;
  wire v911167;
  wire v90f0aa;
  wire v907ff8;
  wire v9118ff;
  wire v9041e0;
  wire v909dc5;
  wire v93fc6a;
  wire v93f783;
  wire v904f23;
  wire v904d08;
  wire v9058e9;
  wire v93f6ec;
  wire v903fa0;
  wire v903ba1;
  wire v91359e;
  wire v9051c3;
  wire v85eaab;
  wire v93f28a;
  wire v93f747;
  wire v93f763;
  wire v8b9c53;
  wire v90f383;
  wire v93fb7f;
  wire v90666d;
  wire v93f815;
  wire v86eecd;
  wire v90819e;
  wire v8baf9a;
  wire v90444d;
  wire v90ad03;
  wire v93ed09;
  wire v909924;
  wire v9077a9;
  wire v904c75;
  wire v909016;
  wire v93fb5a;
  wire v93f797;
  wire v90f320;
  wire v91dd4f;
  wire v910e6e;
  wire v93f6dc;
  wire v91a75e;
  wire v912384;
  wire v87a261;
  wire v904008;
  wire v93faf9;
  wire v9115a9;
  wire v93fcdc;
  wire v913068;
  wire v906b22;
  wire v89f9dc;
  wire v905da0;
  wire v909878;
  wire v93fda6;
  wire v93df39;
  wire v9098f2;
  wire v90466e;
  wire v90cfc7;
  wire v93fadc;
  wire v90ed2f;
  wire v8b9de1;
  wire v9100f8;
  wire v88de63;
  wire v88e6c4;
  wire v8d1873;
  wire v93f76b;
  wire v906a5c;
  wire v93f91f;
  wire v90e6f8;
  wire v904610;
  wire v93f822;
  wire v906fba;
  wire v90a4b7;
  wire v86345f;
  wire v905697;
  wire v87c51e;
  wire v90500e;
  wire v93f6a9;
  wire v93fc16;
  wire v9098b1;
  wire v904ccb;
  wire v90eaad;
  wire v905168;
  wire v8b9dcb;
  wire v9110a9;
  wire v90dcc6;
  wire v90944d;
  wire v90f4f8;
  wire v93f7dd;
  wire v93f7d3;
  wire v9101c0;
  wire v93facc;
  wire v907b60;
  wire v8b9996;
  wire v8b495a;
  wire v93f204;
  wire v93f6c7;
  wire v90fc42;
  wire v8b9960;
  wire v903e2f;
  wire v904a3b;
  wire v918886;
  wire v93f2bd;
  wire v912334;
  wire v93f6f9;
  wire v91090e;
  wire v907061;
  wire v90ff49;
  wire v93f882;
  wire v8b9e1d;
  wire v904e93;
  wire v9083b1;
  wire v93e3dd;
  wire v90600b;
  wire v90d933;
  wire v90de9c;
  wire v8ee1f9;
  wire v93f9bb;
  wire v90541b;
  wire v87c4d2;
  wire v9067ab;
  wire v93fe54;
  wire v93f8ad;
  wire v906663;
  wire v870bc2;
  wire v90a097;
  wire v90ee7e;
  wire v91132a;
  wire v93e5f1;
  wire v905077;
  wire v909dc3;
  wire v9384b0;
  wire v844fb7;
  wire v908068;
  wire v93fc84;
  wire v93f901;
  wire v93e51c;
  wire v93f9b9;
  wire v87ca92;
  wire v908325;
  wire v93f5d1;
  wire v93fb3e;
  wire v913435;
  wire v9062f7;
  wire v904e48;
  wire v90e3e1;
  wire v90468e;
  wire v9110ab;
  wire v912fed;
  wire v93f2d9;
  wire v90e40b;
  wire v906fbf;
  wire v9063e0;
  wire v90fcbf;
  wire v906d38;
  wire v93fe41;
  wire v9091b2;
  wire v904a04;
  wire v90a112;
  wire v93fd17;
  wire v93fda3;
  wire v9059d6;
  wire v89f988;
  wire v93f8cf;
  wire v904ae8;
  wire v9053de;
  wire v93f7ac;
  wire v91080c;
  wire v9124bc;
  wire v90accf;
  wire v9133b0;
  wire v90f7ce;
  wire v93f77a;
  wire v9049e4;
  wire v9073b6;
  wire v93fccb;
  wire v93ed91;
  wire v90a786;
  wire v93fb7b;
  wire v904755;
  wire v907adb;
  wire v9047cd;
  wire v91a9cd;
  wire v93f2a0;
  wire v93f6e1;
  wire v90460e;
  wire v93f826;
  wire v905d36;
  wire v93fcfc;
  wire v8b9c1e;
  wire v910bea;
  wire v90ec84;
  wire v909fb2;
  wire v93fcd6;
  wire v907206;
  wire v91006b;
  wire v90995e;
  wire v90ea1f;
  wire v909157;
  wire v90917f;
  wire v90edb8;
  wire v93fc9f;
  wire v93fa70;
  wire v9109dc;
  wire v93fc85;
  wire v93f6b7;
  wire v90a5c1;
  wire v903f97;
  wire v93f23c;
  wire v93fa89;
  wire v93f9be;
  wire v93eb20;
  wire v8a9222;
  wire v93fdd7;
  wire v906037;
  wire v8ebd28;
  wire v9077b1;
  wire v9108ff;
  wire v93f81c;
  wire v90491c;
  wire v93fce1;
  wire v9046d6;
  wire v93fd2f;
  wire v90a53b;
  wire v90d877;
  wire v90f16d;
  wire v93f32a;
  wire v90acc4;
  wire v85ea7f;
  wire v93dfe2;
  wire v91a9e1;
  wire v90d0f9;
  wire v93fb3c;
  wire v86346f;
  wire v904d38;
  wire v93f8ca;
  wire v909e9d;
  wire v93f8ab;
  wire v91268a;
  wire v86337d;
  wire v93fb88;
  wire v8b4a12;
  wire v9101be;
  wire v93fda2;
  wire v93fd54;
  wire v93fe5f;
  wire v9131d1;
  wire v91155d;
  wire v93f83c;
  wire v904714;
  wire v930076;
  wire v9134cc;
  wire v9085ac;
  wire v910c5b;
  wire v9103e4;
  wire v907580;
  wire v9089e7;
  wire v905748;
  wire v90d7cb;
  wire v879731;
  wire v908fd6;
  wire v93ebab;
  wire v905a12;
  wire v90a4d4;
  wire v89f881;
  wire v93fd06;
  wire v91035c;
  wire v9075fd;
  wire v9113c0;
  wire v873ad7;
  wire v93f7f8;
  wire v904e38;
  wire v863476;
  wire v93f7e9;
  wire v93e007;
  wire v89f7dd;
  wire v904b77;
  wire v90446a;
  wire v93fcb7;
  wire v8b99b9;
  wire v93ebd1;
  wire v89f930;
  wire v8ee1a3;
  wire v90cbfc;
  wire v93f6bf;
  wire v907f0b;
  wire v93eabc;
  wire v93f8b5;
  wire v90fc87;
  wire v90a2df;
  wire v907965;
  wire v904568;
  wire v90d9b2;
  wire v904eba;
  wire v93fb96;
  wire v9124a9;
  wire v93e791;
  wire v90d546;
  wire v93f97d;
  wire v89f8a9;
  wire v9058c2;
  wire v93fbb4;
  wire v93e8f1;
  wire v90752d;
  wire v93fb21;
  wire v93fd3b;
  wire v904ba1;
  wire v907e81;
  wire v90fa0b;
  wire v85eaf3;
  wire v93f7c3;
  wire v90a4c6;
  wire v93fda5;
  wire v909383;
  wire v904d1a;
  wire v93fa85;
  wire v8ebce4;
  wire v93fdea;
  wire v93fdc8;
  wire v90e028;
  wire v907469;
  wire v90f9f3;
  wire v93e54b;
  wire v8b9ee2;
  wire v906c35;
  wire v905204;
  wire v8ee186;
  wire v93defa;
  wire v93fd20;
  wire v9066e0;
  wire v907018;
  wire v904b63;
  wire v905366;
  wire v90479e;
  wire v93fe33;
  wire v9047f0;
  wire v90985e;
  wire v90e304;
  wire v882135;
  wire v93fb9d;
  wire v93f320;
  wire v93f972;
  wire v9111a4;
  wire v8b5ff8;
  wire v93fd68;
  wire v93ed58;
  wire v90dff3;
  wire v93ecad;
  wire v913592;
  wire v93f279;
  wire v9056a4;
  wire v8b5f4d;
  wire v9135db;
  wire v93fd8c;
  wire v8b9884;
  wire v93f88d;
  wire v90a59b;
  wire v903b91;
  wire v93faf0;
  wire v904091;
  wire v93e2b8;
  wire v906eb2;
  wire v93eaa6;
  wire v93f6da;
  wire v93fb51;
  wire v906c94;
  wire v930047;
  wire v93fd9f;
  wire v93e1dd;
  wire v904838;
  wire v9135d1;
  wire v90cecd;
  wire v907110;
  wire v93e810;
  wire v910ebb;
  wire v93f6f8;
  wire v93f77e;
  wire v910867;
  wire v90f2da;
  wire v90a07b;
  wire v93f9cb;
  wire v913a39;
  wire v93f9c7;
  wire v93fc47;
  wire v861331;
  wire v93fb77;
  wire v93f833;
  wire v9135f1;
  wire v907bd4;
  wire v93f6ff;
  wire v904dfc;
  wire v93fe15;
  wire v90ef07;
  wire v878dab;
  wire v93fb5f;
  wire v90fc9a;
  wire v90a229;
  wire v8824ac;
  wire v91063d;
  wire v9104e0;
  wire v86335a;
  wire v8ee173;
  wire v904340;
  wire v93f90e;
  wire v90da92;
  wire v93eeda;
  wire v93f81e;
  wire v93fa82;
  wire v93f7b4;
  wire v86dde6;
  wire v8f3865;
  wire v9042b8;
  wire v90a2c8;
  wire v93f692;
  wire v89f80d;
  wire v904521;
  wire v9300da;
  wire v87a20d;
  wire v93e5fc;
  wire v8b9e6c;
  wire v93fac2;
  wire v9111cf;
  wire v90f52f;
  wire v93f94a;
  wire v89f938;
  wire v93f6ac;
  wire v8b9ec9;
  wire v90d47d;
  wire v90a90b;
  wire v8b9e4f;
  wire v93f913;
  wire v905653;
  wire v93fa2a;
  wire v90a4a1;
  wire v88b191;
  wire v90a33f;
  wire v93f98d;
  wire v93fb07;
  wire v907d70;
  wire v93fa80;
  wire v8f3868;
  wire v908a35;
  wire v90da35;
  wire v90f3f8;
  wire v93f6ab;
  wire v87c4c4;
  wire v906a84;
  wire v93f7e1;
  wire v88b26d;
  wire v905486;
  wire v93f695;
  wire v9043bd;
  wire v91335a;
  wire v913225;
  wire v905b92;
  wire v93eec9;
  wire v90710d;
  wire v93e230;
  wire v907f74;
  wire v907321;
  wire v93f7ef;
  wire v907685;
  wire v93fd13;
  wire v93f94b;
  wire v907916;
  wire v9050ad;
  wire v91a7a5;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg StoB_REQ4_p;
  input StoB_REQ4_n;
  reg StoB_REQ5_p;
  input StoB_REQ5_n;
  reg StoB_REQ6_p;
  input StoB_REQ6_n;
  reg StoB_REQ7_p;
  input StoB_REQ7_n;
  reg StoB_REQ8_p;
  input StoB_REQ8_n;
  reg StoB_REQ9_p;
  input StoB_REQ9_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoS_ACK4_p;
  output BtoS_ACK4_n;
  reg BtoS_ACK5_p;
  output BtoS_ACK5_n;
  reg BtoS_ACK6_p;
  output BtoS_ACK6_n;
  reg BtoS_ACK7_p;
  output BtoS_ACK7_n;
  reg BtoS_ACK8_p;
  output BtoS_ACK8_n;
  reg BtoS_ACK9_p;
  output BtoS_ACK9_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg SLC2_p;
  output SLC2_n;
  reg SLC3_p;
  output SLC3_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  reg jx3_p;
  output jx3_n;
  wire ENQ_n;
  wire SLC3_n;

assign v88b191 = BtoS_ACK9_p & v8824ac | !BtoS_ACK9_p & v90a4a1;
assign v909187 = jx0_p & v844f95 | !jx0_p & !v863b25;
assign v91359e = StoB_REQ0_p & v909058 | !StoB_REQ0_p & v903ba1;
assign v906cc5 = jx2_p & v93fbd8 | !jx2_p & v93fa44;
assign v93e7af = BtoS_ACK9_p & v907607 | !BtoS_ACK9_p & v908d55;
assign v90932e = BtoS_ACK0_p & v90fc92 | !BtoS_ACK0_p & v909ca5;
assign v89e0ce = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v907d03;
assign v93f665 = BtoS_ACK0_p & v9046a6 | !BtoS_ACK0_p & v89f984;
assign v90417d = StoB_REQ8_p & v86f60a | !StoB_REQ8_p & v86dd54;
assign v93f793 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v90987f;
assign v903cd2 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93fa35;
assign v93fdb8 = StoB_REQ8_p & v907e36 | !StoB_REQ8_p & v90a884;
assign v93fb6c = StoB_REQ6_p & v909107 | !StoB_REQ6_p & v907ad8;
assign v89f796 = ENQ_p & v911a33 | !ENQ_p & v93fc97;
assign v93f827 = BtoS_ACK8_p & v87f17f | !BtoS_ACK8_p & v844f91;
assign v93fa74 = StoB_REQ8_p & v93f769 | !StoB_REQ8_p & v90dcf6;
assign v9041e0 = BtoS_ACK9_p & v93e05f | !BtoS_ACK9_p & v9118ff;
assign v8b4977 = StoB_REQ1_p & v904ae0 | !StoB_REQ1_p & !v93fae6;
assign v908e8e = BtoS_ACK6_p & v93f9c6 | !BtoS_ACK6_p & v93f682;
assign v90d6fa = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v93f8b7;
assign v908a2f = StoB_REQ6_p & v90f79b | !StoB_REQ6_p & v90a098;
assign v90ee37 = jx0_p & v909928 | !jx0_p & v93f6fc;
assign v93efb8 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v90dc57;
assign v9300cb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f8f7;
assign v9300a5 = BtoS_ACK8_p & v9074fa | !BtoS_ACK8_p & v90e144;
assign v93f815 = BtoS_ACK8_p & v90451f | !BtoS_ACK8_p & v90666d;
assign v93fa73 = jx1_p & v93ee38 | !jx1_p & v90481b;
assign v903c65 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v905972;
assign v908cf4 = jx1_p & v844f91 | !jx1_p & v93fbb7;
assign v90723b = StoB_REQ8_p & v909289 | !StoB_REQ8_p & v93fb2f;
assign v93fad3 = ENQ_p & v93f92a | !ENQ_p & v89fd8d;
assign v93fa15 = BtoS_ACK8_p & v8b5f61 | !BtoS_ACK8_p & !v90e4f2;
assign v90a0cb = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v907168;
assign v93f922 = StoB_REQ6_p & v93e9e3 | !StoB_REQ6_p & v91071e;
assign v90a33f = jx3_p & v9113c0 | !jx3_p & v88b191;
assign v93fac9 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v93ea5d;
assign v93f5ae = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v9300c6;
assign v93f7b0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v903c83;
assign v90515d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b49ad;
assign v909cc1 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v90a20d;
assign v9056e2 = DEQ_p & v9074f5 | !DEQ_p & v93fb34;
assign v93f720 = BtoS_ACK7_p & v93f894 | !BtoS_ACK7_p & v844fa3;
assign v909c74 = jx2_p & v9091b4 | !jx2_p & !v908d14;
assign v90468f = jx0_p & v909107 | !jx0_p & !v909adc;
assign v93dfc0 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v9123a2;
assign v9046f9 = BtoS_ACK8_p & v93fc5d | !BtoS_ACK8_p & v93f690;
assign v93fbc0 = BtoS_ACK6_p & v90860a | !BtoS_ACK6_p & v910cc4;
assign v910cbf = BtoS_ACK8_p & v906b5f | !BtoS_ACK8_p & !v90425a;
assign v93f77e = StoB_REQ9_p & v9135d1 | !StoB_REQ9_p & v93f6f8;
assign v908693 = StoB_REQ8_p & v8b9ef8 | !StoB_REQ8_p & v93f7bd;
assign v905791 = StoB_REQ1_p & v905660 | !StoB_REQ1_p & v9121a6;
assign v91ae94 = StoB_REQ7_p & v93fbe5 | !StoB_REQ7_p & !v910710;
assign v906adf = StoB_REQ6_p & v90664a | !StoB_REQ6_p & v90eed3;
assign v90a1f7 = BtoS_ACK0_p & v913619 | !BtoS_ACK0_p & v909cee;
assign v904d1a = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v909383;
assign v910ca7 = jx1_p & v90cc7a | !jx1_p & v9043f4;
assign v93fcd8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90a20e;
assign v93f29c = RtoB_ACK0_p & v87e0d8 | !RtoB_ACK0_p & v93fd3e;
assign v909ca5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v908834;
assign v844fb3 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v903cf9 = jx0_p & v844f91 | !jx0_p & v863b25;
assign v93e6f6 = BtoS_ACK7_p & v907f25 | !BtoS_ACK7_p & v93f760;
assign v90fcd2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v904074;
assign v93dfb4 = ENQ_p & v90fbad | !ENQ_p & v844f91;
assign v90da97 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v90854b;
assign v90aa5e = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v844f91;
assign v93fcb2 = EMPTY_p & v907722 | !EMPTY_p & v8b9e73;
assign v9047cd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v906fbf;
assign v93dffe = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v9076a8;
assign v93f2da = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v93f878;
assign v93f8e0 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93e819;
assign v93f69c = BtoS_ACK2_p & v9076a8 | !BtoS_ACK2_p & v8b99b4;
assign v91134b = BtoS_ACK6_p & v89f8bd | !BtoS_ACK6_p & v9044c6;
assign v90459f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93e681;
assign v90804e = StoB_REQ7_p & v910710 | !StoB_REQ7_p & v905764;
assign v908545 = BtoR_REQ0_p & v93f9f7 | !BtoR_REQ0_p & v93fb4f;
assign v9059ef = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v88e55e;
assign v93f6dd = BtoS_ACK1_p & v906627 | !BtoS_ACK1_p & v93def0;
assign v8b9d35 = jx2_p & v8b98f4 | !jx2_p & v93f9d4;
assign v909347 = jx3_p & v905d0a | !jx3_p & v844f91;
assign v905ba8 = BtoS_ACK6_p & v90ad75 | !BtoS_ACK6_p & v844f91;
assign v90a08d = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v93e2c2;
assign v90787b = jx0_p & v844f91 | !jx0_p & !v844f99;
assign v89e0a6 = jx1_p & v93f7b0 | !jx1_p & !v903e94;
assign v93f5cb = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v908f4b;
assign v93fa25 = jx1_p & v869aeb | !jx1_p & !v93e470;
assign v90f88a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v904c38;
assign v93fe33 = BtoS_ACK6_p & v90479e | !BtoS_ACK6_p & v8ebce4;
assign v93ecd6 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v8f3869;
assign v8b9e71 = BtoS_ACK9_p & v93fd7a | !BtoS_ACK9_p & v90d727;
assign v93f29a = jx1_p & v93f768 | !jx1_p & v844f91;
assign v909df9 = StoB_REQ6_p & v908357 | !StoB_REQ6_p & v844f91;
assign v912481 = jx2_p & v90e38d | !jx2_p & v91146e;
assign v93f888 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v93f3ea;
assign v913362 = BtoS_ACK8_p & v93f73d | !BtoS_ACK8_p & v911552;
assign v93fc2a = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v907168;
assign v904e16 = BtoS_ACK1_p & v906255 | !BtoS_ACK1_p & !v9131c9;
assign v90748b = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v906913;
assign v93f9f3 = jx1_p & v9060d2 | !jx1_p & v910c50;
assign v93eda4 = jx3_p & v844f91 | !jx3_p & !v93f818;
assign v91086c = BtoS_ACK8_p & v9074fa | !BtoS_ACK8_p & !v90dfbc;
assign v93e1dd = jx2_p & v93fda5 | !jx2_p & !v93fd9f;
assign v911b83 = BtoS_ACK0_p & v93fb3b | !BtoS_ACK0_p & v93006b;
assign v93e9cc = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v93fd09;
assign v93fa4f = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v909cc1;
assign v89e0d5 = ENQ_p & v93f15e | !ENQ_p & v844f91;
assign v90fc92 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v863a37;
assign v93e643 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91232c;
assign v93faff = jx2_p & v904bd4 | !jx2_p & v90d5a9;
assign v93fdd1 = BtoS_ACK7_p & v911f15 | !BtoS_ACK7_p & v906983;
assign v91062b = StoB_REQ0_p & v93f3ea | !StoB_REQ0_p & v911c01;
assign v9135e9 = DEQ_p & v93fa36 | !DEQ_p & v90a2f1;
assign v93fb82 = BtoS_ACK0_p & v93ea50 | !BtoS_ACK0_p & v90d0b8;
assign v93f8c6 = BtoS_ACK6_p & v90d718 | !BtoS_ACK6_p & v8f22ee;
assign v90e8fa = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8b9d37;
assign v90496b = BtoS_ACK6_p & v90d718 | !BtoS_ACK6_p & v90809d;
assign v90893a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v910243;
assign v86346f = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & v90d877;
assign v906c6e = BtoS_ACK0_p & v93dfc0 | !BtoS_ACK0_p & v93ee84;
assign v93eed6 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v90eea7;
assign v90606c = jx1_p & v89c5bd | !jx1_p & v905ba8;
assign v87f181 = jx2_p & v844f91 | !jx2_p & !v844f91;
assign v91aa43 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v93f098;
assign v8706e4 = jx1_p & v9088ff | !jx1_p & v90805e;
assign v93f085 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v87c4fa;
assign v912173 = EMPTY_p & v844f91 | !EMPTY_p & v905540;
assign v93fc40 = jx0_p & v93db03 | !jx0_p & v906a6b;
assign v90a89f = BtoS_ACK2_p & v9123a2 | !BtoS_ACK2_p & v93fe1b;
assign v9079a8 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v909941;
assign v93f9ab = jx2_p & v8706e4 | !jx2_p & !v89e042;
assign v904234 = jx1_p & v9093ec | !jx1_p & !v90d22b;
assign v93fce7 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v90e978;
assign v8b9bb4 = StoB_REQ8_p & v93f9bc | !StoB_REQ8_p & v93f5b9;
assign v90d27b = StoB_REQ1_p & v907472 | !StoB_REQ1_p & v93fc28;
assign v90d999 = StoB_REQ7_p & v871df8 | !StoB_REQ7_p & v93fe0c;
assign v85eaf1 = StoB_REQ6_p & v904296 | !StoB_REQ6_p & v89f93b;
assign v8b9eca = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v90e856;
assign v93f9be = BtoS_ACK6_p & v93fa89 | !BtoS_ACK6_p & v9091b2;
assign v93f78a = BtoS_ACK7_p & v93fc09 | !BtoS_ACK7_p & !v93fc10;
assign v93f699 = BtoS_ACK9_p & v93e168 | !BtoS_ACK9_p & v93ec24;
assign v910b0e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v906ff5;
assign v909525 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93e926;
assign v9121a6 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v9079f7;
assign v93fb44 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90719c;
assign v9050cc = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93f768;
assign v93fe1a = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v90cfd5;
assign v906f72 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v90799d;
assign v93f83a = jx0_p & v90aeb7 | !jx0_p & !v90690e;
assign v9121a7 = jx0_p & v93f714 | !jx0_p & !v844f91;
assign v906b43 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b496d;
assign v905619 = StoB_REQ6_p & v91194f | !StoB_REQ6_p & v93f52d;
assign v8858ac = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v9097f3;
assign v93f290 = BtoS_ACK0_p & v90873f | !BtoS_ACK0_p & v93fac1;
assign v908ef9 = BtoR_REQ0_p & v93f8d4 | !BtoR_REQ0_p & v90e7e2;
assign v911328 = RtoB_ACK1_p & v90f6b5 | !RtoB_ACK1_p & v9091a2;
assign v90f8c9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93fdc6;
assign v93fde9 = stateG12_p & v911a33 | !stateG12_p & v91aa43;
assign v93faa6 = jx2_p & v844f91 | !jx2_p & v93efa3;
assign v93fcb7 = BtoS_ACK1_p & v93fccb | !BtoS_ACK1_p & v90446a;
assign v88c1f9 = BtoS_ACK8_p & v90fe87 | !BtoS_ACK8_p & v908693;
assign BtoS_ACK7_n = !v8b4a3a;
assign v910825 = StoB_REQ1_p & v9052de | !StoB_REQ1_p & v844f91;
assign v9100f8 = BtoS_ACK0_p & v93fb3b | !BtoS_ACK0_p & v8b9de1;
assign v93f7a5 = StoB_REQ7_p & v93f8a6 | !StoB_REQ7_p & v93fbc0;
assign v91a992 = jx2_p & v844f91 | !jx2_p & v89f8bc;
assign v909c45 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844fb1;
assign BtoS_ACK0_n = !v89e12f;
assign v93fd95 = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & v87f17f;
assign v863b26 = StoB_REQ8_p & v93fcc8 | !StoB_REQ8_p & v905b55;
assign v89f7e7 = jx0_p & v90767a | !jx0_p & v909dd6;
assign v86333d = jx1_p & v903c83 | !jx1_p & !v93fe31;
assign v93fbbe = StoB_REQ1_p & v904ae0 | !StoB_REQ1_p & !v911680;
assign v8b9b56 = ENQ_p & v87e7f5 | !ENQ_p & v93faae;
assign v905a80 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v93fc68;
assign v93f9d4 = jx1_p & v93e1ed | !jx1_p & v87a991;
assign v9052ba = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v911bcf;
assign v907469 = BtoS_ACK7_p & v907e81 | !BtoS_ACK7_p & v90e028;
assign v909649 = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & !v9054bc;
assign v93fd52 = BtoS_ACK7_p & v907f25 | !BtoS_ACK7_p & v9086f8;
assign v87c547 = DEQ_p & v90acfe | !DEQ_p & v87de8d;
assign v903c43 = jx0_p & v93fda0 | !jx0_p & v93f707;
assign v93dc30 = BtoS_ACK4_p & v844f9f | !BtoS_ACK4_p & v9099ef;
assign v9058d5 = StoB_REQ8_p & v86f60a | !StoB_REQ8_p & v9082a5;
assign v912ec5 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v93f875;
assign v906538 = StoB_REQ7_p & v93fe2e | !StoB_REQ7_p & v93f9db;
assign v93f6fe = StoB_REQ7_p & v904ff8 | !StoB_REQ7_p & v844f91;
assign v8b497a = StoB_REQ8_p & v87f17f | !StoB_REQ8_p & !v93f85d;
assign v93fbb3 = jx0_p & v93fe17 | !jx0_p & v8b9d1b;
assign v90a62c = jx1_p & v93f871 | !jx1_p & v844f91;
assign v9060ea = jx1_p & v884481 | !jx1_p & v9047e4;
assign v9105ed = jx0_p & v93fa7c | !jx0_p & v90d59a;
assign v93f90a = jx0_p & v90aa5e | !jx0_p & v90df59;
assign v9096ca = ENQ_p & v90834a | !ENQ_p & !v905b6a;
assign v93fc07 = BtoS_ACK7_p & v93dab8 | !BtoS_ACK7_p & v8728ef;
assign v91247e = StoB_REQ8_p & v86345d | !StoB_REQ8_p & v90e612;
assign v93fdbe = stateG7_1_p & v89b116 | !stateG7_1_p & v907a1b;
assign v8b9eb0 = StoB_REQ3_p & v908eea | !StoB_REQ3_p & !v844f9f;
assign v93fe2d = jx1_p & v9095bf | !jx1_p & !v86313d;
assign v90e38d = jx1_p & v87f17d | !jx1_p & v90f1cb;
assign v90fb2b = jx0_p & v93f70c | !jx0_p & v93f6fc;
assign v93f692 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v90a2c8;
assign v93f8ca = StoB_REQ6_p & v904d38 | !StoB_REQ6_p & v906d38;
assign v93fccb = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93f9a9;
assign v91a6e7 = BtoS_ACK0_p & v90810f | !BtoS_ACK0_p & !v90598f;
assign v93f852 = jx1_p & v844f91 | !jx1_p & !v906e3d;
assign v905653 = StoB_REQ8_p & v93f7b4 | !StoB_REQ8_p & v93f913;
assign v89f905 = BtoS_ACK7_p & v911185 | !BtoS_ACK7_p & !v9045df;
assign v91a6f1 = BtoS_ACK9_p & v93f76e | !BtoS_ACK9_p & v85cca5;
assign v90de74 = BtoS_ACK9_p & v93e3a1 | !BtoS_ACK9_p & v93fd64;
assign v93ee39 = BtoS_ACK8_p & v90529c | !BtoS_ACK8_p & v90728a;
assign v90a602 = jx3_p & v93fa7d | !jx3_p & !v93f790;
assign v8b9f21 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v91305b;
assign v907da3 = BtoS_ACK6_p & v93f9c6 | !BtoS_ACK6_p & v9059b7;
assign v89e05b = BtoS_ACK9_p & v93e85e | !BtoS_ACK9_p & v93fc89;
assign v863428 = BtoS_ACK9_p & v9074fa | !BtoS_ACK9_p & v90927a;
assign v93f707 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v844f95;
assign v93f82d = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v910937;
assign v904bda = jx3_p & v844f91 | !jx3_p & v93e27a;
assign v909c39 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93ea16;
assign v9078da = BtoS_ACK8_p & v93f8f0 | !BtoS_ACK8_p & v9091c6;
assign v90e93c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90611f;
assign v863a38 = jx1_p & v844f91 | !jx1_p & !v903e94;
assign v904ab2 = BtoS_ACK6_p & v908d2a | !BtoS_ACK6_p & v93f57d;
assign v91a9a2 = ENQ_p & v8a1fe3 | !ENQ_p & v911498;
assign v90f624 = StoB_REQ1_p & v9046a6 | !StoB_REQ1_p & v844f9b;
assign v9102cc = BtoS_ACK6_p & v91aa51 | !BtoS_ACK6_p & v93f97f;
assign v93e671 = BtoS_ACK8_p & v908237 | !BtoS_ACK8_p & !v90897e;
assign v911a1e = jx2_p & v844f91 | !jx2_p & v909224;
assign v93f8a5 = jx0_p & v90aeb7 | !jx0_p & v844f91;
assign v910c3a = StoB_REQ0_p & v909cc1 | !StoB_REQ0_p & v844f91;
assign v93fd79 = jx1_p & v863b25 | !jx1_p & v93f21c;
assign v90ee74 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v9091c7;
assign v89f881 = BtoS_ACK7_p & v913435 | !BtoS_ACK7_p & v90accf;
assign v93fd0e = BtoS_ACK6_p & v910e72 | !BtoS_ACK6_p & v93fd16;
assign v93fbc7 = StoB_REQ9_p & v93f2c6 | !StoB_REQ9_p & v90546e;
assign v9063b2 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93faf5;
assign v871483 = ENQ_p & v93e704 | !ENQ_p & v93fe38;
assign v904ab4 = BtoS_ACK7_p & v93e27a | !BtoS_ACK7_p & v93e5b8;
assign v90567d = RtoB_ACK0_p & v93f916 | !RtoB_ACK0_p & v91a9a2;
assign v863b2f = jx1_p & v904b4f | !jx1_p & v844f91;
assign v906d63 = BtoS_ACK0_p & v8c7343 | !BtoS_ACK0_p & v904b41;
assign v913433 = stateG12_p & v910840 | !stateG12_p & v93fae1;
assign v93fb20 = jx1_p & v93fabd | !jx1_p & v9052ce;
assign v93f870 = ENQ_p & v93f89f | !ENQ_p & v9056ac;
assign v90cbec = jx1_p & v910f82 | !jx1_p & !v90ede1;
assign v9066e0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fd20;
assign v91071f = BtoS_ACK7_p & v93fc04 | !BtoS_ACK7_p & v911a1e;
assign v93fc71 = BtoS_ACK1_p & v906627 | !BtoS_ACK1_p & v90a89f;
assign v904fd2 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v910b4b;
assign v904b00 = jx2_p & v93f558 | !jx2_p & v844f91;
assign v91a9de = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90459f;
assign v86eecd = StoB_REQ9_p & v903eef | !StoB_REQ9_p & v93f815;
assign v90d9fd = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v907168;
assign v93fcbd = jx3_p & v844f91 | !jx3_p & v91a9b6;
assign v91cc2d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8f3869;
assign v913a94 = EMPTY_p & v90567d | !EMPTY_p & v9053ed;
assign v93f26c = ENQ_p & v93e704 | !ENQ_p & v8d373a;
assign v909058 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93e9cc;
assign v8b9d1b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93fc4e;
assign v90481b = StoB_REQ7_p & v93f989 | !StoB_REQ7_p & v863346;
assign v909d2b = StoB_REQ3_p & v93fd8e | !StoB_REQ3_p & v87c533;
assign v93f881 = jx0_p & v9079a8 | !jx0_p & v93fab9;
assign v907799 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93eaa1;
assign v904628 = jx0_p & v844f91 | !jx0_p & v90893a;
assign v90d054 = jx0_p & v90a8e9 | !jx0_p & v911937;
assign v90a214 = jx1_p & v89e11b | !jx1_p & v904141;
assign v904430 = StoB_REQ1_p & v904b58 | !StoB_REQ1_p & v872e32;
assign v93fc5d = jx2_p & v93fd25 | !jx2_p & v90db6b;
assign v93fa89 = jx0_p & v9091b2 | !jx0_p & v93fb3e;
assign v9113fb = jx1_p & v9050a5 | !jx1_p & v8b49ad;
assign v904901 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v911b9a;
assign v9300c0 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v90ad2f;
assign v9048c6 = jx3_p & v93fa3a | !jx3_p & !v909be8;
assign v904ba1 = EMPTY_p & v904714 | !EMPTY_p & v93fd3b;
assign v906f55 = StoB_REQ0_p & v93df06 | !StoB_REQ0_p & v93f82b;
assign v93f2b9 = BtoS_ACK9_p & v908250 | !BtoS_ACK9_p & v93f745;
assign v90a300 = BtoS_ACK1_p & v90a59e | !BtoS_ACK1_p & v90962e;
assign v8b9ebe = BtoS_ACK6_p & v93f90a | !BtoS_ACK6_p & v844f91;
assign v93fcc6 = EMPTY_p & v89e0d5 | !EMPTY_p & v93fd74;
assign v909adc = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v91216e;
assign v90744a = jx3_p & v90e546 | !jx3_p & !v92fff5;
assign v9110a9 = BtoS_ACK8_p & v93f73d | !BtoS_ACK8_p & v8b9dcb;
assign v906042 = BtoS_ACK6_p & v91a9b9 | !BtoS_ACK6_p & v9082fc;
assign v90f7e4 = StoB_REQ9_p & v910ea0 | !StoB_REQ9_p & v8b9ce5;
assign v90edf6 = jx2_p & v9045e6 | !jx2_p & v9119f9;
assign v93ebe6 = BtoS_ACK6_p & v90ea4c | !BtoS_ACK6_p & v90762a;
assign v93f8ad = jx3_p & v87f17f | !jx3_p & v93fe54;
assign v93fb57 = stateG12_p & v844f91 | !stateG12_p & !v907c01;
assign v89e086 = BtoS_ACK8_p & v93fb92 | !BtoS_ACK8_p & v91355f;
assign v90a097 = BtoS_ACK9_p & v93f9bb | !BtoS_ACK9_p & v870bc2;
assign v90cee9 = BtoS_ACK8_p & v85e94c | !BtoS_ACK8_p & v91336c;
assign v8f383c = BtoR_REQ0_p & v906ce5 | !BtoR_REQ0_p & v93fb4f;
assign v904808 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v90f8c2;
assign v8848d6 = BtoS_ACK6_p & v93fcc9 | !BtoS_ACK6_p & v93f92e;
assign v913348 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v863a37;
assign v87bf17 = jx1_p & v907be9 | !jx1_p & v9051e9;
assign v93f7f7 = StoB_REQ0_p & v93fd87 | !StoB_REQ0_p & v90f0a2;
assign v86cda0 = StoB_REQ8_p & v93eb39 | !StoB_REQ8_p & v905835;
assign v93fd32 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v909c45;
assign v93e54b = jx1_p & v90e3e1 | !jx1_p & v844f91;
assign v93f92e = jx0_p & v93fd40 | !jx0_p & !v907a13;
assign v90690e = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v93fc1a;
assign v907e7a = StoB_REQ7_p & v8821a1 | !StoB_REQ7_p & v911edd;
assign v904755 = jx1_p & v93f910 | !jx1_p & !v844f91;
assign v93fe4b = BtoS_ACK7_p & v910fda | !BtoS_ACK7_p & v8b9f23;
assign v904a04 = jx0_p & v9091b2 | !jx0_p & v913435;
assign v90736f = StoB_REQ8_p & v90f947 | !StoB_REQ8_p & v904847;
assign v89f983 = jx1_p & v93f1b4 | !jx1_p & !v93e3cf;
assign v93f6cf = BtoS_ACK9_p & v9074fa | !BtoS_ACK9_p & v9300a5;
assign v93e3cf = StoB_REQ7_p & v910527 | !StoB_REQ7_p & v93f119;
assign v9047b7 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v93ecb9 = jx2_p & v93fa1f | !jx2_p & !v844f91;
assign v93f7d2 = jx0_p & v93f8d2 | !jx0_p & v844f91;
assign v93fb5a = BtoS_ACK2_p & v906cc8 | !BtoS_ACK2_p & v909016;
assign v90425a = StoB_REQ8_p & v9071ed | !StoB_REQ8_p & v93001e;
assign v93f959 = ENQ_p & v93df31 | !ENQ_p & v93fc1d;
assign v9051c3 = BtoS_ACK0_p & v93fb3b | !BtoS_ACK0_p & v91359e;
assign v93fae6 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v90d1ca;
assign v911826 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v93f897;
assign v9132e5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86e433;
assign v93e835 = BtoS_ACK0_p & v876439 | !BtoS_ACK0_p & v9054e2;
assign v8b9d0f = jx0_p & v8b9c5f | !jx0_p & v93fb95;
assign v8b495a = jx3_p & v93f78c | !jx3_p & !v89f9dc;
assign v907aa0 = BtoS_ACK4_p & v844f9f | !BtoS_ACK4_p & !v9300af;
assign v9074ce = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v863a78;
assign v93e138 = StoB_REQ6_p & v9058f1 | !StoB_REQ6_p & v91026d;
assign v908ae0 = StoB_REQ1_p & v93e926 | !StoB_REQ1_p & v905f54;
assign v93f7ec = StoB_REQ9_p & v909492 | !StoB_REQ9_p & v88c1f9;
assign v93f970 = jx1_p & v91ae94 | !jx1_p & !v93fca2;
assign v9133ad = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fcf4;
assign v909dd6 = StoB_REQ6_p & v93f41e | !StoB_REQ6_p & v844f91;
assign v93fdce = jx0_p & v844f91 | !jx0_p & !v93fa3f;
assign v93fb41 = jx0_p & v844f91 | !jx0_p & !v910243;
assign v90acc5 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v913a6f;
assign v9074f5 = RtoB_ACK0_p & v904d51 | !RtoB_ACK0_p & v9077f7;
assign v9124a9 = jx1_p & v90f07f | !jx1_p & !v93fb96;
assign v906fd0 = jx3_p & v844f91 | !jx3_p & v905d7a;
assign v93fcf0 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v908eea;
assign v93fc46 = BtoS_ACK6_p & v910910 | !BtoS_ACK6_p & v90d59c;
assign v91192b = BtoS_ACK6_p & v90ede1 | !BtoS_ACK6_p & v90fb4b;
assign v906ae9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90fc92;
assign v844fc3 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & !v844f91;
assign v909691 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9b;
assign v93fe38 = jx3_p & v93fa7d | !jx3_p & !v8b9e9f;
assign v93fe00 = BtoS_ACK0_p & v93f7ad | !BtoS_ACK0_p & v93fa99;
assign v90ddf9 = BtoS_ACK7_p & v93f7d9 | !BtoS_ACK7_p & !v904cb5;
assign v90e44c = BtoS_ACK7_p & v93f9ab | !BtoS_ACK7_p & !v9065d3;
assign v93f1cb = BtoS_ACK9_p & v93fcc4 | !BtoS_ACK9_p & v9057d4;
assign v905ca1 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fe223;
assign v89fe58 = BtoS_ACK6_p & v90ad75 | !BtoS_ACK6_p & v9044b1;
assign v9104f8 = jx3_p & v844f91 | !jx3_p & v8b9d4b;
assign v86f5de = jx1_p & v85ea42 | !jx1_p & !v905de8;
assign v909b56 = jx1_p & v87c52b | !jx1_p & !v904f88;
assign v90a7b2 = StoB_REQ6_p & v911853 | !StoB_REQ6_p & v93e882;
assign v93f1ad = BtoS_ACK9_p & v844fa5 | !BtoS_ACK9_p & !v90711a;
assign v90811c = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v90a3e0;
assign v906b66 = StoB_REQ2_p & v87b4fc | !StoB_REQ2_p & v90fb89;
assign v907b86 = StoB_REQ7_p & v93f70d | !StoB_REQ7_p & v909f4b;
assign v93f805 = StoB_REQ0_p & v93f7f5 | !StoB_REQ0_p & v93e37e;
assign v9051cd = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v904f5e;
assign v906275 = EMPTY_p & v907bd1 | !EMPTY_p & v93e94e;
assign v93fbd3 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v93e00f;
assign v93fe0a = BtoS_ACK8_p & v91a6ea | !BtoS_ACK8_p & v93f769;
assign v90512d = jx2_p & v91038c | !jx2_p & v93eaf0;
assign v909924 = stateG7_1_p & v904f23 | !stateG7_1_p & v93ed09;
assign v909222 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90888d;
assign v93faf5 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v91a747;
assign v90d5a9 = jx1_p & v85ea42 | !jx1_p & !v93fcad;
assign v89f984 = StoB_REQ0_p & v93db4a | !StoB_REQ0_p & v91305d;
assign v93f895 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v90f88e;
assign v93fda3 = jx1_p & v9062f7 | !jx1_p & v93fd17;
assign v93fd94 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v910f62;
assign v93fcf7 = jx1_p & v911edb | !jx1_p & v90a207;
assign v93fb11 = ENQ_p & v93f95a | !ENQ_p & v910915;
assign v90712c = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v87c537;
assign v93fb72 = ENQ_p & v90fbad | !ENQ_p & v93e70e;
assign v89b1a2 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v909a7c;
assign v90a5ef = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v913348;
assign v93f723 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v91a771;
assign v93f7f8 = jx2_p & v93fb7b | !jx2_p & !v873ad7;
assign v906a51 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v93e5da;
assign v93fe11 = FULL_p & v909dec | !FULL_p & v93f2fd;
assign v90d22b = jx0_p & v844f9f | !jx0_p & v844f9d;
assign v908ee8 = StoB_REQ7_p & v903fb2 | !StoB_REQ7_p & v93fb05;
assign v93f7e2 = StoB_REQ9_p & v93f86b | !StoB_REQ9_p & v93fa57;
assign v91164f = StoB_REQ8_p & v87f17f | !StoB_REQ8_p & v907eaa;
assign v90efea = StoB_REQ7_p & v871df8 | !StoB_REQ7_p & v93f6cc;
assign v93fda9 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v909c39;
assign v93fd77 = BtoS_ACK6_p & v8a8b0a | !BtoS_ACK6_p & v93e9e5;
assign v90f819 = jx3_p & v93fa7d | !jx3_p & !v93fc6f;
assign v90cf49 = jx2_p & v93f6a4 | !jx2_p & v909661;
assign v93f79a = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & v863444;
assign v90ea4c = jx0_p & v93fa7c | !jx0_p & v910243;
assign v913522 = BtoS_ACK6_p & v9072c8 | !BtoS_ACK6_p & v8f229e;
assign v90d718 = jx0_p & v844f91 | !jx0_p & !v93fc0a;
assign v93f291 = BtoS_ACK8_p & v93dbe9 | !BtoS_ACK8_p & v93fd86;
assign v906cc8 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v93fd2b;
assign v93f771 = BtoS_ACK6_p & v8b49ad | !BtoS_ACK6_p & v93f994;
assign v8b4a12 = jx1_p & v93fb3c | !jx1_p & !v93fb88;
assign v93f818 = BtoS_ACK9_p & v9074fa | !BtoS_ACK9_p & v91086c;
assign v904ccb = BtoS_ACK6_p & v90ede1 | !BtoS_ACK6_p & !v9098b1;
assign v93fcea = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v93e549;
assign v90a4bd = BtoS_ACK7_p & v9107aa | !BtoS_ACK7_p & !v90ac9e;
assign v911b4d = BtoS_ACK0_p & v90873f | !BtoS_ACK0_p & v91231a;
assign v93fa96 = jx3_p & v844f91 | !jx3_p & !v872e5f;
assign v93fc0f = BtoS_ACK6_p & v871033 | !BtoS_ACK6_p & v844f91;
assign v90494f = ENQ_p & v9083cf | !ENQ_p & v9078f8;
assign v93fd47 = jx0_p & v9074ce | !jx0_p & v863a78;
assign v93fdc4 = jx0_p & v93f119 | !jx0_p & v906623;
assign v91a7a3 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v911a00;
assign v90ea8a = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v90f8c9;
assign v90ee7e = jx3_p & v87f17f | !jx3_p & v90a097;
assign v909be7 = jx0_p & v909e2c | !jx0_p & !v93e643;
assign v85ead8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9071f8;
assign v93fc31 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v908a2c;
assign v93e8a1 = jx1_p & v93fc68 | !jx1_p & !v90fb5d;
assign v8b9e17 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v904f2e;
assign v863478 = BtoR_REQ1_p & v913079 | !BtoR_REQ1_p & v907664;
assign v93f894 = jx1_p & v844fa3 | !jx1_p & !v93f037;
assign v93f936 = BtoS_ACK6_p & v8b9d27 | !BtoS_ACK6_p & v93fad7;
assign v90873f = StoB_REQ1_p & v93e2de | !StoB_REQ1_p & v844f91;
assign v93fe44 = jx3_p & v844f91 | !jx3_p & v908006;
assign v9051e9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fabf;
assign v93fbb6 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v90e9e1;
assign v9043a5 = BtoS_ACK8_p & v903da9 | !BtoS_ACK8_p & v90df02;
assign v904714 = ENQ_p & v908325 | !ENQ_p & v93f83c;
assign v93f2c6 = BtoS_ACK8_p & v904b00 | !BtoS_ACK8_p & v86f60a;
assign v93edbf = jx2_p & v906638 | !jx2_p & v910ca7;
assign v93fdf8 = StoB_REQ7_p & v9058f3 | !StoB_REQ7_p & v909f04;
assign v93f7ca = StoB_REQ9_p & v908e8b | !StoB_REQ9_p & v907517;
assign v90aa42 = StoB_REQ8_p & v90529c | !StoB_REQ8_p & v93ca43;
assign v90a134 = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & v909174;
assign v9119fd = StoB_REQ8_p & v90d866 | !StoB_REQ8_p & v904132;
assign v93f977 = BtoS_ACK6_p & v9130af | !BtoS_ACK6_p & v91cfc7;
assign v93f9fa = BtoS_ACK8_p & v90a2aa | !BtoS_ACK8_p & v86cda0;
assign v9042d2 = ENQ_p & v93f753 | !ENQ_p & v90e5b4;
assign v903c83 = jx0_p & v863a78 | !jx0_p & v844f91;
assign v93fb39 = jx1_p & v93fc0f | !jx1_p & !v907b86;
assign v8b9d28 = BtoS_ACK8_p & v910d56 | !BtoS_ACK8_p & !v903c80;
assign v91194f = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v90a902;
assign v93fab0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910b91;
assign v93fc63 = StoB_REQ2_p & v905702 | !StoB_REQ2_p & v909078;
assign v907e86 = jx1_p & v910f82 | !jx1_p & v844f91;
assign v93f926 = StoB_REQ7_p & v87f17d | !StoB_REQ7_p & v9050e0;
assign v863346 = BtoS_ACK6_p & v905537 | !BtoS_ACK6_p & v87f17d;
assign v8a921d = stateG12_p & v90adc4 | !stateG12_p & v859639;
assign v8ebcf9 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v906321;
assign v90548c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v93fd57;
assign v93f6d3 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v93eaa8;
assign v93fac0 = BtoS_ACK1_p & v93f85e | !BtoS_ACK1_p & v908ae0;
assign v93e6af = jx0_p & v844f91 | !jx0_p & v90515d;
assign v91229f = BtoS_ACK7_p & v93e47b | !BtoS_ACK7_p & v90e79a;
assign v90cfa8 = StoB_REQ6_p & v93f511 | !StoB_REQ6_p & v93f7dc;
assign v93f9db = BtoS_ACK6_p & v93fd47 | !BtoS_ACK6_p & v93fb5e;
assign v863363 = BtoS_ACK6_p & v93f91d | !BtoS_ACK6_p & v93fb0b;
assign v93f81b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93e8d3;
assign v89e10d = jx1_p & v844f91 | !jx1_p & !v87f17d;
assign v9124cb = StoB_REQ7_p & v93fcf3 | !StoB_REQ7_p & v863b25;
assign v903c6e = jx2_p & v90456e | !jx2_p & !v9113b2;
assign v93f87e = BtoS_ACK0_p & v876439 | !BtoS_ACK0_p & v93fcd8;
assign v909434 = StoB_REQ2_p & v905702 | !StoB_REQ2_p & !v93f765;
assign v909492 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8b9ef8;
assign v93ef1d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v906642;
assign v90e133 = BtoS_ACK0_p & v86c2d0 | !BtoS_ACK0_p & v905d8b;
assign v93e2e6 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v90443a;
assign v90808b = jx2_p & v90fca6 | !jx2_p & v863afc;
assign v93f9c6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v844f97;
assign v90a525 = StoB_REQ1_p & v93f824 | !StoB_REQ1_p & v90a348;
assign v908ae5 = BtoS_ACK9_p & v8d195d | !BtoS_ACK9_p & v93eade;
assign v91a70f = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v90fa03;
assign v904575 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9046a6;
assign v90a002 = BtoS_ACK6_p & v871033 | !BtoS_ACK6_p & v881ec0;
assign v911365 = StoB_REQ9_p & v93f045 | !StoB_REQ9_p & v91a762;
assign v904da2 = StoB_REQ0_p & v91216e | !StoB_REQ0_p & v909357;
assign v907bca = BtoS_ACK6_p & v90cc30 | !BtoS_ACK6_p & !v909a12;
assign v90f33b = EMPTY_p & v90d8d5 | !EMPTY_p & !v8a8faa;
assign v93f76e = StoB_REQ8_p & v87f17d | !StoB_REQ8_p & v9043e5;
assign v906d08 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v93f7f5;
assign v8b9e6c = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v93e5fc;
assign v93f280 = BtoS_ACK1_p & v86c2d0 | !BtoS_ACK1_p & v89e119;
assign v9133b0 = BtoS_ACK7_p & v91080c | !BtoS_ACK7_p & v90accf;
assign v90ac9e = jx2_p & v9070cb | !jx2_p & v8b9c46;
assign v904aae = jx0_p & v8a927b | !jx0_p & v8b49ad;
assign v93fa56 = BtoS_ACK0_p & v913619 | !BtoS_ACK0_p & v9133ad;
assign v878dab = RtoB_ACK1_p & v904ba1 | !RtoB_ACK1_p & v90ef07;
assign v93e816 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v93f9f6;
assign v904aac = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85ea79;
assign v90542e = RtoB_ACK0_p & v904e3a | !RtoB_ACK0_p & v904d56;
assign v93eb39 = BtoS_ACK7_p & v904b00 | !BtoS_ACK7_p & v904ede;
assign v906a6b = BtoS_ACK0_p & v93e77b | !BtoS_ACK0_p & v90d5a3;
assign v93f8c5 = jx2_p & v86333d | !jx2_p & v9074ce;
assign v90ae53 = StoB_REQ0_p & v9071c7 | !StoB_REQ0_p & v93fdd4;
assign v8b5f4d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a4c6;
assign v8b98d4 = StoB_REQ8_p & v906046 | !StoB_REQ8_p & v90776b;
assign v903cc5 = jx0_p & v9067d3 | !jx0_p & !v844f91;
assign v8824ac = StoB_REQ8_p & v93f7f8 | !StoB_REQ8_p & v90a229;
assign v93f588 = jx1_p & v93f119 | !jx1_p & !v87f17d;
assign v907898 = BtoS_ACK1_p & v93fce7 | !BtoS_ACK1_p & v8b4977;
assign v90937e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9047b7;
assign v93fbdd = jx0_p & v8b99bb | !jx0_p & v93fbb2;
assign v905d7a = BtoS_ACK9_p & v93e27a | !BtoS_ACK9_p & v911cba;
assign v93e402 = StoB_REQ6_p & v8a8fb1 | !StoB_REQ6_p & v886f59;
assign v93ea50 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v93f85e;
assign v863359 = jx3_p & v93e105 | !jx3_p & !v904a8a;
assign v93e105 = BtoS_ACK9_p & v93e150 | !BtoS_ACK9_p & v910461;
assign v906cf5 = BtoS_ACK6_p & v8b9d27 | !BtoS_ACK6_p & v8633ef;
assign v9089bf = StoB_REQ0_p & v93f70c | !StoB_REQ0_p & v93f61e;
assign v93fb6f = BtoS_ACK1_p & v8bb868 | !BtoS_ACK1_p & v906b3d;
assign v90e925 = StoB_REQ9_p & v93f291 | !StoB_REQ9_p & v93fd18;
assign v907edc = jx0_p & v844f91 | !jx0_p & !v912ec5;
assign v90cecd = jx1_p & v930047 | !jx1_p & !v882135;
assign v8f37fc = jx2_p & v93fb81 | !jx2_p & !v908d14;
assign v9093db = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v93fbba;
assign v90e32f = jx0_p & v911005 | !jx0_p & v90aaca;
assign v9070f7 = EMPTY_p & v904025 | !EMPTY_p & v93fc26;
assign v880314 = jx1_p & v93fbb8 | !jx1_p & v906256;
assign v910b05 = StoB_REQ7_p & v90d22b | !StoB_REQ7_p & v844f91;
assign v910525 = ENQ_p & v90adc4 | !ENQ_p & v844f91;
assign v93fd68 = StoB_REQ9_p & v90f9f3 | !StoB_REQ9_p & v8b5ff8;
assign v8a9289 = jx0_p & v85dee0 | !jx0_p & v8d3799;
assign v93fd07 = jx2_p & v93f16d | !jx2_p & v85ead8;
assign v904a90 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844fb9;
assign v93f746 = ENQ_p & v85eaff | !ENQ_p & v8b9c01;
assign v93f4ac = ENQ_p & v90fbad | !ENQ_p & v93fbee;
assign v89c59e = StoB_REQ3_p & v905702 | !StoB_REQ3_p & v844fb9;
assign v903ddc = BtoS_ACK8_p & v93fb43 | !BtoS_ACK8_p & !v9050e7;
assign v9096a3 = BtoS_ACK7_p & v93f119 | !BtoS_ACK7_p & !v90d52b;
assign v903d4f = jx0_p & v910fd2 | !jx0_p & !v90690e;
assign v93e8ab = jx2_p & v93f216 | !jx2_p & v93faf7;
assign v905291 = BtoS_ACK9_p & v87f17f | !BtoS_ACK9_p & v844f91;
assign v9045c0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v905e84;
assign v90a59e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v90e978;
assign v9042a0 = StoB_REQ9_p & v909e8a | !StoB_REQ9_p & v905d68;
assign v8a8fa3 = DEQ_p & v904d51 | !DEQ_p & v907bd1;
assign v87a21e = BtoS_ACK6_p & v86344b | !BtoS_ACK6_p & v870615;
assign v911586 = DEQ_p & v906d83 | !DEQ_p & v93f19b;
assign v904cde = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93fbe1;
assign v9070e2 = jx0_p & v93f87f | !jx0_p & v844f91;
assign v93fd1f = StoB_REQ8_p & v93fe29 | !StoB_REQ8_p & v93f7b1;
assign v90a629 = stateG12_p & v90ad0b | !stateG12_p & !v93fd59;
assign v9060d2 = StoB_REQ7_p & v8b4a08 | !StoB_REQ7_p & v904200;
assign v887bb8 = jx1_p & v844f91 | !jx1_p & v93f864;
assign v9134c4 = jx1_p & v93fe6e | !jx1_p & v9058f3;
assign v93f107 = stateG12_p & v90adc4 | !stateG12_p & v93f69a;
assign v905b92 = ENQ_p & v93fb51 | !ENQ_p & v844f91;
assign v9054bd = jx2_p & v8b9c87 | !jx2_p & v90cbec;
assign v85ea62 = StoB_REQ3_p & v908eea | !StoB_REQ3_p & v9074a6;
assign v907b07 = StoB_REQ9_p & v87c541 | !StoB_REQ9_p & v844f91;
assign v93fd60 = jx1_p & v93fce5 | !jx1_p & v844f91;
assign v93fb3f = jx1_p & v913332 | !jx1_p & !v844f91;
assign v90d32d = BtoS_ACK9_p & v93f73d | !BtoS_ACK9_p & v907c76;
assign v8b9e60 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v90a557;
assign v909845 = BtoS_ACK8_p & v903da9 | !BtoS_ACK8_p & v8d3791;
assign v90e1cf = jx1_p & v93f085 | !jx1_p & v93edf1;
assign v90ccbd = BtoS_ACK8_p & v90a733 | !BtoS_ACK8_p & v907710;
assign v909353 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v93fd0d;
assign v909a26 = jx0_p & v90d879 | !jx0_p & v93fa7c;
assign v93eb9e = jx2_p & v904434 | !jx2_p & v93fcf2;
assign v91137e = jx2_p & v90d93b | !jx2_p & v90e8bf;
assign v907d03 = BtoS_ACK0_p & v93e391 | !BtoS_ACK0_p & v90d9a0;
assign v905702 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9d;
assign v870dd6 = jx1_p & v90e6f5 | !jx1_p & v93fc9d;
assign v91104b = BtoS_ACK0_p & v906627 | !BtoS_ACK0_p & v8bbc68;
assign v9097f3 = StoB_REQ2_p & v9099e3 | !StoB_REQ2_p & v90a44f;
assign v9074a6 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v9300af;
assign v90dfbc = BtoS_ACK7_p & v93faf2 | !BtoS_ACK7_p & !v90df44;
assign v86d7d1 = BtoS_ACK8_p & v90cc57 | !BtoS_ACK8_p & v93fd1e;
assign v90dc57 = StoB_REQ9_p & v93e671 | !StoB_REQ9_p & v844f91;
assign v93f864 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90d00f;
assign v93fac4 = BtoS_ACK9_p & v9050cc | !BtoS_ACK9_p & v93fcb1;
assign v90a784 = BtoS_ACK8_p & v93fc04 | !BtoS_ACK8_p & v87c525;
assign v9134bc = jx2_p & v93f986 | !jx2_p & v908ed6;
assign v9045f3 = BtoS_ACK1_p & v93f85e | !BtoS_ACK1_p & v93ec07;
assign v905e84 = BtoS_ACK1_p & v93dffe | !BtoS_ACK1_p & v87e087;
assign v93f960 = BtoS_ACK7_p & v93fbe4 | !BtoS_ACK7_p & v93f6e9;
assign v93ea9e = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v907b07;
assign v91097b = StoB_REQ8_p & v90a4bd | !StoB_REQ8_p & v9132d3;
assign v9047e4 = jx0_p & v844f97 | !jx0_p & v844f95;
assign v90e9a1 = DEQ_p & v909bdf | !DEQ_p & v9082be;
assign v909c0e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90484c;
assign v93fc4a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93e03a;
assign v85ea9a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v905cd2;
assign v90eda0 = BtoS_ACK1_p & v90fc92 | !BtoS_ACK1_p & v904430;
assign v93fd00 = RtoB_ACK0_p & v93f73c | !RtoB_ACK0_p & v87c566;
assign v90a112 = BtoS_ACK6_p & v906fbf | !BtoS_ACK6_p & v904a04;
assign v93fd09 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v87c533;
assign v909c08 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v884dd3;
assign v90f2da = jx3_p & v844f91 | !jx3_p & v910867;
assign v904bc1 = jx2_p & v89f8fd | !jx2_p & v93f768;
assign v85ea99 = StoB_REQ1_p & v90a89f | !StoB_REQ1_p & v844f91;
assign v905366 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v904b63;
assign v910ea0 = BtoS_ACK8_p & v93f73d | !BtoS_ACK8_p & !v909289;
assign v8f37ef = StoB_REQ6_p & v93f87e | !StoB_REQ6_p & v9068b6;
assign v911167 = BtoS_ACK7_p & v9054bd | !BtoS_ACK7_p & v90f2f9;
assign v90e159 = BtoS_ACK8_p & v93fc04 | !BtoS_ACK8_p & v91071f;
assign v8bbc54 = stateG7_1_p & v907e33 | !stateG7_1_p & v87ba4e;
assign v93f739 = StoB_REQ7_p & v911c73 | !StoB_REQ7_p & v90515d;
assign v903e70 = jx1_p & v93f80e | !jx1_p & !v844f91;
assign v907c71 = BtoS_ACK8_p & v93fdae | !BtoS_ACK8_p & v908a4f;
assign v904e3e = EMPTY_p & v910525 | !EMPTY_p & v9064cc;
assign v90ff47 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v91016c;
assign v903b0f = StoB_REQ8_p & v93e296 | !StoB_REQ8_p & v89f7c7;
assign v90a207 = StoB_REQ7_p & v90f3e4 | !StoB_REQ7_p & v90e172;
assign v85ef3a = BtoS_ACK8_p & v89e122 | !BtoS_ACK8_p & v9062ae;
assign v93f3ea = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v90a0cb;
assign v905d63 = BtoS_ACK8_p & v93f29a | !BtoS_ACK8_p & v913067;
assign v9071f0 = BtoS_ACK0_p & v93f85e | !BtoS_ACK0_p & v93f093;
assign v9067c1 = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & !v90faaf;
assign v9085e8 = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & v9121a7;
assign v93f6aa = BtoS_ACK7_p & v93fdd2 | !BtoS_ACK7_p & v903e7a;
assign v93ecad = ENQ_p & v908325 | !ENQ_p & v90dff3;
assign v904926 = jx1_p & v844f91 | !jx1_p & v911509;
assign v909082 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fb3;
assign v905718 = jx1_p & v912687 | !jx1_p & v93f7f1;
assign v90eed3 = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & !v906a51;
assign v9109f4 = jx2_p & v863a03 | !jx2_p & v863afc;
assign v93f744 = jx1_p & v910710 | !jx1_p & v844f91;
assign v93f7f4 = BtoS_ACK8_p & v9074fa | !BtoS_ACK8_p & v9052f0;
assign v904d39 = jx2_p & v8b830b | !jx2_p & v903e70;
assign v9077be = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v93f005;
assign v909bbd = jx2_p & v93e8a1 | !jx2_p & !v93fa1e;
assign BtoS_ACK4_n = !v87a2ae;
assign v90a0d7 = StoB_REQ8_p & v9088bc | !StoB_REQ8_p & v9059ef;
assign v90636e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v93fc2a;
assign v866af4 = BtoS_ACK6_p & v903e94 | !BtoS_ACK6_p & v93fe0e;
assign v93fb81 = jx1_p & v88d7c9 | !jx1_p & v90e8da;
assign v93f8a6 = BtoS_ACK6_p & v903e94 | !BtoS_ACK6_p & v9044c6;
assign v93f889 = BtoS_ACK6_p & v90630d | !BtoS_ACK6_p & !v903cb1;
assign v907bbb = jx1_p & v93e9de | !jx1_p & !v910d6d;
assign v8ee1f9 = BtoR_REQ1_p & v93fc16 | !BtoR_REQ1_p & v90de9c;
assign v8b9c55 = jx2_p & v93f96e | !jx2_p & v8b4983;
assign v93f8ff = BtoS_ACK6_p & v9130af | !BtoS_ACK6_p & v844f91;
assign v90faf1 = BtoS_ACK7_p & v903db9 | !BtoS_ACK7_p & v90809b;
assign v90a49d = jx3_p & v93f73e | !jx3_p & v844f91;
assign v910b7a = jx2_p & v93fb09 | !jx2_p & !v905718;
assign v8ee1a3 = BtoS_ACK6_p & v90a786 | !BtoS_ACK6_p & v89f930;
assign v911a33 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v906ce1;
assign v93fa8d = EMPTY_p & v9061b3 | !EMPTY_p & v87c547;
assign v9121bb = BtoS_ACK7_p & v93fce5 | !BtoS_ACK7_p & v907be9;
assign v93fb69 = StoB_REQ9_p & v90d370 | !StoB_REQ9_p & v903f5a;
assign v906fcc = ENQ_p & v93e704 | !ENQ_p & v93fc66;
assign v906321 = StoB_REQ0_p & v910f5a | !StoB_REQ0_p & v93f589;
assign v93f0a3 = BtoS_ACK6_p & v8a8b0a | !BtoS_ACK6_p & v93e14f;
assign v908546 = BtoS_ACK6_p & v91a9b9 | !BtoS_ACK6_p & v844f91;
assign v903d60 = jx0_p & v90ad39 | !jx0_p & !v9055c0;
assign v905665 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v903fb0;
assign v93fdee = EMPTY_p & v9077c7 | !EMPTY_p & v91a71d;
assign v90991f = jx1_p & v8639e7 | !jx1_p & v90515a;
assign v93fc2b = BtoS_ACK6_p & v93f9c6 | !BtoS_ACK6_p & !v90664a;
assign v93f882 = RtoB_ACK0_p & v90ff49 | !RtoB_ACK0_p & v90ad03;
assign v904dcf = EMPTY_p & v903d12 | !EMPTY_p & v904671;
assign v93f66b = StoB_REQ8_p & v93f894 | !StoB_REQ8_p & v93f720;
assign v9113de = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87a1f2;
assign v8ee188 = BtoS_ACK6_p & v910230 | !BtoS_ACK6_p & v907e6b;
assign v903c09 = StoB_REQ6_p & v911bc2 | !StoB_REQ6_p & v90cc41;
assign v93fcc0 = RtoB_ACK1_p & v907120 | !RtoB_ACK1_p & v904dcf;
assign v93006b = StoB_REQ0_p & v909525 | !StoB_REQ0_p & v91aa12;
assign v904340 = BtoS_ACK0_p & v93fccb | !BtoS_ACK0_p & v8ee173;
assign v90da8b = jx1_p & v871033 | !jx1_p & !v909f4c;
assign v93f29d = BtoS_ACK0_p & v876439 | !BtoS_ACK0_p & v8b5f55;
assign v93e650 = jx0_p & v906c6e | !jx0_p & !v90932e;
assign v93f7b1 = jx2_p & v90a2b9 | !jx2_p & v87f17d;
assign v90987f = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v93e7ac;
assign v907524 = jx1_p & v8b9d0f | !jx1_p & !v9090dd;
assign v910230 = jx0_p & v90ed41 | !jx0_p & v93fa55;
assign v904bf3 = jx0_p & v844f91 | !jx0_p & v90d879;
assign v903b98 = DEQ_p & v910ffd | !DEQ_p & v93fdb1;
assign v87a98d = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v910226;
assign v904654 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93e684;
assign v93f763 = StoB_REQ7_p & v90ebde | !StoB_REQ7_p & v93f747;
assign v912477 = jx3_p & v93dfc2 | !jx3_p & !v9099a1;
assign v903c81 = BtoS_ACK7_p & v93e8cb | !BtoS_ACK7_p & v907e91;
assign v908a34 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v90fb76;
assign v9091be = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c7343;
assign v93ed15 = jx3_p & v93f1ad | !jx3_p & !v93f1cb;
assign v9115a7 = StoB_REQ7_p & v93fbf0 | !StoB_REQ7_p & v844f91;
assign v93fbeb = jx1_p & v93fd43 | !jx1_p & !v90d46a;
assign v93f9bb = jx2_p & v87c51f | !jx2_p & v844f91;
assign v910062 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v912f16;
assign v8b9d0e = RtoB_ACK0_p & v9054b6 | !RtoB_ACK0_p & v90871b;
assign v910c29 = EMPTY_p & v90d443 | !EMPTY_p & v90a4bb;
assign v90e073 = DEQ_p & v904c53 | !DEQ_p & v910525;
assign v93f58c = BtoS_ACK7_p & v9104ad | !BtoS_ACK7_p & !v909d71;
assign v905b55 = BtoS_ACK7_p & v93fd60 | !BtoS_ACK7_p & v90e019;
assign v93e32d = StoB_REQ9_p & v8b9e6e | !StoB_REQ9_p & v88403f;
assign v90a563 = BtoS_ACK6_p & v88932d | !BtoS_ACK6_p & v93f5f6;
assign v90e6f1 = BtoS_ACK6_p & v93f910 | !BtoS_ACK6_p & v908797;
assign v90de9c = RtoB_ACK1_p & v907061 | !RtoB_ACK1_p & v90d933;
assign v90f810 = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & v90e93c;
assign v887a80 = jx2_p & v90d634 | !jx2_p & v90813f;
assign v90d879 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fa7c;
assign v905618 = jx1_p & v90879a | !jx1_p & !v910b05;
assign v90e3ed = StoB_REQ7_p & v93ee3b | !StoB_REQ7_p & v904a61;
assign v93e5bf = BtoS_ACK0_p & v8bb868 | !BtoS_ACK0_p & v904aac;
assign v9133ba = jx2_p & v90dc9c | !jx2_p & !v93f6ea;
assign v93fca0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v905d04;
assign v93ec67 = jx2_p & v8d37d8 | !jx2_p & v90cb3d;
assign v93f92a = jx3_p & v907abc | !jx3_p & v911a33;
assign v93f5d1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90534f;
assign v90ae72 = StoB_REQ1_p & v93f908 | !StoB_REQ1_p & v905df9;
assign v93f8af = jx0_p & v909107 | !jx0_p & v844f91;
assign v93001e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v93fb58;
assign v93fad4 = stateG12_p & v90fbad | !stateG12_p & v90ed77;
assign v93f728 = DEQ_p & v90df61 | !DEQ_p & v93f6ae;
assign v85eac9 = jx1_p & v93debb | !jx1_p & v90d52b;
assign v872e5f = BtoS_ACK9_p & v9074fa | !BtoS_ACK9_p & v93f7f4;
assign v904ba3 = jx3_p & v844f91 | !jx3_p & !v904b9e;
assign v906e30 = jx3_p & v8b9b88 | !jx3_p & v90f0c4;
assign v89f9cd = StoB_REQ8_p & v87f17f | !StoB_REQ8_p & v93f7b3;
assign v91051a = BtoS_ACK7_p & v87f17f | !BtoS_ACK7_p & !v909367;
assign v9113c0 = BtoS_ACK9_p & v904e48 | !BtoS_ACK9_p & v9075fd;
assign v93eb20 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f9be;
assign v9070d5 = BtoS_ACK6_p & v8b49ad | !BtoS_ACK6_p & v844f91;
assign v903da9 = jx2_p & v910b96 | !jx2_p & v93faf8;
assign v9077a9 = StoB_REQ3_p & v93fd8e | !StoB_REQ3_p & v93fbd3;
assign v93fcd9 = StoB_REQ7_p & v9093ec | !StoB_REQ7_p & v93fc7e;
assign v93fbd4 = BtoS_ACK0_p & v8c7343 | !BtoS_ACK0_p & v8a9231;
assign v904e38 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a786;
assign v93fa9c = BtoS_ACK0_p & v93e2de | !BtoS_ACK0_p & v911428;
assign v911090 = jx1_p & v906201 | !jx1_p & v844f91;
assign v93fad0 = jx3_p & v90f2f6 | !jx3_p & !v90ff07;
assign v87c541 = BtoS_ACK8_p & v90e261 | !BtoS_ACK8_p & v93e9d8;
assign v93f9a1 = jx1_p & v869aeb | !jx1_p & !v90d999;
assign v912643 = BtoS_ACK0_p & v90810f | !BtoS_ACK0_p & !v90a798;
assign v93fdbf = jx2_p & v90965e | !jx2_p & v93fcba;
assign v91024c = BtoS_ACK0_p & v93e391 | !BtoS_ACK0_p & v904f1b;
assign v93f02c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v93f68c;
assign v90d704 = BtoS_ACK7_p & v910e66 | !BtoS_ACK7_p & v86d767;
assign v93f6de = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v844f91;
assign v93f792 = BtoS_ACK6_p & v93e681 | !BtoS_ACK6_p & v9051e8;
assign v87a993 = StoB_REQ2_p & v93ed70 | !StoB_REQ2_p & v93eff8;
assign v90e772 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v90d250;
assign v93e310 = jx1_p & v93fc94 | !jx1_p & v90df7f;
assign v904436 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v93f6de;
assign v93f5db = StoB_REQ9_p & v9107e7 | !StoB_REQ9_p & v9083c5;
assign v93fc6a = ENQ_p & v93fdf6 | !ENQ_p & v909dc5;
assign v93fba8 = BtoS_ACK8_p & v911b4e | !BtoS_ACK8_p & v910958;
assign v93ec8c = StoB_REQ8_p & v904ab4 | !StoB_REQ8_p & v93fd93;
assign v90a0b5 = BtoS_ACK8_p & v93f7b1 | !BtoS_ACK8_p & v85f2b9;
assign v911fc7 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v905764;
assign v9090c9 = StoB_REQ2_p & v908127 | !StoB_REQ2_p & v912ec8;
assign v8b4976 = BtoS_ACK0_p & v90a5ef | !BtoS_ACK0_p & v906f55;
assign v8633b7 = StoB_REQ6_p & v909927 | !StoB_REQ6_p & v903e7f;
assign v911933 = jx3_p & v844f91 | !jx3_p & v90cc4a;
assign v93ef4c = BtoS_ACK6_p & v93fa7c | !BtoS_ACK6_p & v90762a;
assign v90aaa8 = ENQ_p & v910242 | !ENQ_p & v844f91;
assign v90919c = StoB_REQ2_p & v93fd5c | !StoB_REQ2_p & v844f91;
assign v8b9b94 = jx0_p & v863b25 | !jx0_p & !v844f95;
assign v90631b = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v9085b3;
assign v8d195d = StoB_REQ8_p & v90f947 | !StoB_REQ8_p & v906b5f;
assign v93e0e6 = BtoR_REQ0_p & v911435 | !BtoR_REQ0_p & v90f4fb;
assign v93fde6 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fa7b;
assign v863a78 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9134df;
assign v90e6e5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90873f;
assign v89f9c3 = jx1_p & v844f91 | !jx1_p & v87ca8a;
assign v93e78b = StoB_REQ0_p & v93db4a | !StoB_REQ0_p & v907898;
assign v87d990 = jx3_p & v93e105 | !jx3_p & !v87f181;
assign v904b41 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90949f;
assign v93e0b5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f058;
assign v905c01 = StoB_REQ0_p & v93f70c | !StoB_REQ0_p & !v844f91;
assign v90f4fb = EMPTY_p & v904c4f | !EMPTY_p & v906034;
assign v93f69d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90a134;
assign v93fd21 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v907c8c;
assign v93f63b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9052de;
assign v9044b4 = jx0_p & v90ea74 | !jx0_p & !v93fdfa;
assign v90f864 = StoB_REQ2_p & v908127 | !StoB_REQ2_p & v905434;
assign v9117e1 = BtoS_ACK7_p & v906d2a | !BtoS_ACK7_p & v93f93c;
assign v905381 = StoB_REQ1_p & v93f908 | !StoB_REQ1_p & v93fdba;
assign v905835 = BtoS_ACK7_p & v909f63 | !BtoS_ACK7_p & v91247f;
assign v904dea = BtoR_REQ0_p & v90d1c9 | !BtoR_REQ0_p & v90d5b3;
assign v909a12 = jx0_p & v906adf | !jx0_p & !v910473;
assign v9059b8 = BtoS_ACK9_p & v9073c5 | !BtoS_ACK9_p & v88aff7;
assign v9118a3 = jx1_p & v87f17d | !jx1_p & v871df8;
assign v9088bc = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v9100bd;
assign v93e9e5 = jx0_p & v90ae5a | !jx0_p & !v93f7f0;
assign v93fd8a = BtoS_ACK7_p & v90529c | !BtoS_ACK7_p & v93faa6;
assign v90ec5d = BtoS_ACK6_p & v871df8 | !BtoS_ACK6_p & v93f8af;
assign v910f41 = RtoB_ACK1_p & v905146 | !RtoB_ACK1_p & v9131cb;
assign v93fd9e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90980d;
assign v908f27 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v9076a7;
assign v93fa1e = jx1_p & v86344b | !jx1_p & v90630d;
assign v907018 = jx1_p & v93defa | !jx1_p & v9066e0;
assign v93faae = jx3_p & v90f478 | !jx3_p & v844f91;
assign v913067 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9117e1;
assign v90d59c = jx0_p & v844f91 | !jx0_p & v8a927b;
assign v93f72f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v911383;
assign v93fb3c = StoB_REQ7_p & v90e6f1 | !StoB_REQ7_p & v90d0f9;
assign v907a4d = ENQ_p & v93e704 | !ENQ_p & v9078f8;
assign v90a876 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f771;
assign v93f85b = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v89f8b8;
assign v93e450 = BtoS_ACK2_p & v91305b | !BtoS_ACK2_p & v906e15;
assign v8b9c2b = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v93fd5c;
assign v93ee38 = StoB_REQ7_p & v910710 | !StoB_REQ7_p & v93f8c6;
assign v9057d4 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93fa52;
assign v90722c = jx2_p & v906c8b | !jx2_p & !v844f91;
assign v9112e1 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844fa3;
assign v93fdc6 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v904313;
assign v90f0c4 = BtoS_ACK9_p & v907bfd | !BtoS_ACK9_p & v93f7e2;
assign v904d08 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v93fe71;
assign v909b54 = jx1_p & v93f7c7 | !jx1_p & v9058f3;
assign v910fe2 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v908436;
assign v904e53 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v911760;
assign v908006 = BtoS_ACK9_p & v9044c3 | !BtoS_ACK9_p & v910dfa;
assign v904ef7 = ENQ_p & v93f89f | !ENQ_p & v85eb28;
assign v93fa72 = BtoS_ACK9_p & v93e228 | !BtoS_ACK9_p & !v93e269;
assign v93f736 = RtoB_ACK0_p & v93f7b9 | !RtoB_ACK0_p & v904dc1;
assign v8b5f55 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f7f9;
assign v90a098 = BtoS_ACK0_p & v93e295 | !BtoS_ACK0_p & v85f268;
assign v93edf1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v863363;
assign v8b99bb = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v89fdcf;
assign v9094f2 = EMPTY_p & v9082e6 | !EMPTY_p & v9078eb;
assign v907be9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fcdb;
assign v93f521 = jx0_p & v91aa44 | !jx0_p & !v904736;
assign v90a102 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93ee22;
assign v910cc4 = jx0_p & v909e2c | !jx0_p & !v89f948;
assign v93fd5c = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v905702;
assign v903afe = jx2_p & v905d9c | !jx2_p & v908d10;
assign v911a89 = jx3_p & v844f91 | !jx3_p & !v90f9ed;
assign v93fce2 = BtoS_ACK0_p & v913619 | !BtoS_ACK0_p & v904663;
assign v93e2de = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v87a21f;
assign v903b1a = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v906657;
assign v93fb0f = jx0_p & v906623 | !jx0_p & v93ef46;
assign v93dfc7 = jx0_p & v91a771 | !jx0_p & !v93f707;
assign v904f22 = EMPTY_p & v90dedf | !EMPTY_p & v90d5d1;
assign v93fd42 = BtoS_ACK7_p & v906ec1 | !BtoS_ACK7_p & v8f37fc;
assign v910c20 = BtoS_ACK7_p & v93ea4f | !BtoS_ACK7_p & v906f1e;
assign v904bdb = jx3_p & v844f91 | !jx3_p & v90fbc8;
assign v9079f7 = StoB_REQ2_p & v93fdf7 | !StoB_REQ2_p & v906cc7;
assign v861331 = BtoS_ACK7_p & v907e81 | !BtoS_ACK7_p & v93fc47;
assign v93fabb = BtoS_ACK6_p & v90860a | !BtoS_ACK6_p & v93fd0c;
assign v8b9c46 = jx1_p & v906665 | !jx1_p & !v844f91;
assign v904fbf = jx1_p & v87c54e | !jx1_p & v844f91;
assign v93fda1 = jx1_p & v93f768 | !jx1_p & v89f98c;
assign v90a63a = BtoS_ACK8_p & v93fdeb | !BtoS_ACK8_p & !v93003e;
assign v90729a = BtoS_ACK0_p & v90810f | !BtoS_ACK0_p & !v9132ed;
assign v909f04 = jx0_p & v9091be | !jx0_p & !v844f9d;
assign v92ffd6 = RtoB_ACK0_p & v91a9a2 | !RtoB_ACK0_p & v907bd1;
assign v86d690 = ENQ_p & v844f91 | !ENQ_p & v907e8f;
assign v8f22e3 = BtoS_ACK7_p & v93f9e3 | !BtoS_ACK7_p & v9049bf;
assign v9087b7 = RtoB_ACK0_p & v90ad3d | !RtoB_ACK0_p & v844f91;
assign v93fd78 = BtoS_ACK7_p & v87f17d | !BtoS_ACK7_p & v90a8ac;
assign v93fa3b = StoB_REQ6_p & v90f5b6 | !StoB_REQ6_p & v872187;
assign v93e672 = jx2_p & v907751 | !jx2_p & v844f91;
assign v9096f3 = BtoS_ACK6_p & v91a9b9 | !BtoS_ACK6_p & v93e86e;
assign v93fd0f = jx2_p & v87c51f | !jx2_p & !v90fb0e;
assign v93eff8 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v89fe59;
assign v93fbb2 = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & !v90a86b;
assign v91143f = jx1_p & v9096f1 | !jx1_p & v87a28e;
assign v93fc89 = StoB_REQ9_p & v909e8a | !StoB_REQ9_p & v93fbf4;
assign v930028 = BtoS_ACK0_p & v8c7343 | !BtoS_ACK0_p & v90e19c;
assign v90f994 = StoB_REQ9_p & v911ebf | !StoB_REQ9_p & v93fc81;
assign v906226 = ENQ_p & v844f91 | !ENQ_p & v93f202;
assign v90a3e0 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v905702;
assign v93fccc = StoB_REQ1_p & v90712c | !StoB_REQ1_p & v910062;
assign v913435 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fb3e;
assign v907bd1 = ENQ_p & v8a1fe3 | !ENQ_p & v844f91;
assign BtoR_REQ0_n = !v8f3879;
assign v90a926 = jx0_p & v844f91 | !jx0_p & v93fcbe;
assign v9072b4 = RtoB_ACK1_p & v905322 | !RtoB_ACK1_p & !v90e9e2;
assign v904d81 = jx3_p & v93fa3a | !jx3_p & !v89e06e;
assign v9115e3 = StoB_REQ6_p & v93f29d | !StoB_REQ6_p & v9071f0;
assign v90d9b3 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v906c20;
assign v93f7dd = BtoS_ACK8_p & v90451f | !BtoS_ACK8_p & v90f4f8;
assign v93e70c = BtoS_ACK6_p & v91aa51 | !BtoS_ACK6_p & v93fe37;
assign v93db03 = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v93f69d;
assign v905325 = jx1_p & v93e7d1 | !jx1_p & !v93f926;
assign v907f05 = BtoS_ACK6_p & v93fa7c | !BtoS_ACK6_p & v93fdcb;
assign v910fda = jx2_p & v906c67 | !jx2_p & v90cbec;
assign v904253 = BtoR_REQ0_p & v93f918 | !BtoR_REQ0_p & v93f9f5;
assign v905408 = jx1_p & v9093ec | !jx1_p & v90fb5d;
assign v93f203 = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v907634;
assign v93fe2e = jx0_p & v9074ce | !jx0_p & v844f91;
assign v9046de = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v906b43;
assign v93e535 = jx1_p & v93fcd9 | !jx1_p & v87f17d;
assign v910f82 = jx0_p & v844f9b | !jx0_p & v844f91;
assign v90a4b7 = BtoS_ACK9_p & v9073c5 | !BtoS_ACK9_p & v906fba;
assign v903ec3 = BtoS_ACK6_p & v93fa7c | !BtoS_ACK6_p & v911318;
assign v906638 = jx1_p & v93f085 | !jx1_p & v909d9c;
assign v93fdc8 = jx1_p & v93fdea | !jx1_p & !v844f91;
assign v90567c = ENQ_p & v9093d9 | !ENQ_p & v93fcbd;
assign v844f9f = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & !v844f91;
assign v8b9e6b = BtoS_ACK0_p & v93f7ad | !BtoS_ACK0_p & v93f731;
assign v93fb7f = BtoS_ACK7_p & v90f575 | !BtoS_ACK7_p & v90f383;
assign v863b25 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f95;
assign v9060e9 = RtoB_ACK0_p & v93fd85 | !RtoB_ACK0_p & v871483;
assign v907e88 = BtoS_ACK7_p & v906c2f | !BtoS_ACK7_p & v93e68d;
assign v90f4f8 = StoB_REQ8_p & v8b9dcb | !StoB_REQ8_p & v90944d;
assign v93f9ac = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9121bb;
assign v93ea5d = StoB_REQ0_p & v93fd87 | !StoB_REQ0_p & v90ee74;
assign v906e15 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b9f21;
assign v93dbe9 = jx2_p & v844f91 | !jx2_p & v908d10;
assign v9076cf = stateG7_1_p & v93fd00 | !stateG7_1_p & v93f6f4;
assign v91080f = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v90729e;
assign v9061b0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8f22bd;
assign v8633bd = RtoB_ACK0_p & v93f284 | !RtoB_ACK0_p & v93fd67;
assign v905dc1 = jx1_p & v93fc0f | !jx1_p & !v9085e8;
assign v93fd76 = jx1_p & v844f91 | !jx1_p & v87f17d;
assign v9080c5 = jx1_p & v93fc68 | !jx1_p & v844f91;
assign v88d5cd = StoB_REQ7_p & v9093ec | !StoB_REQ7_p & !v93fc68;
assign v90fb76 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v89f840;
assign v93fb0a = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v904313;
assign v86ce19 = jx3_p & v908ad9 | !jx3_p & v90a1fe;
assign v908acd = StoB_REQ9_p & v90e159 | !StoB_REQ9_p & v909f00;
assign v93eb70 = BtoS_ACK6_p & v89f84e | !BtoS_ACK6_p & v93f85a;
assign v90628f = jx1_p & v844f91 | !jx1_p & v93faa4;
assign v93f490 = jx2_p & v9086d9 | !jx2_p & !v93e975;
assign v9078eb = DEQ_p & v91007f | !DEQ_p & v904e3a;
assign v90477e = BtoS_ACK7_p & v9114c9 | !BtoS_ACK7_p & !v91107f;
assign v86deed = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v93f064;
assign v8b9e40 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v904da2;
assign v8f3869 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f99;
assign v9086f8 = jx2_p & v909b56 | !jx2_p & v93fb73;
assign v93fa28 = jx0_p & v844f91 | !jx0_p & !v906a79;
assign v88036c = BtoS_ACK1_p & v93dfc0 | !BtoS_ACK1_p & v909ea8;
assign v93fbaa = BtoS_ACK9_p & v93fd1f | !BtoS_ACK9_p & v93f77c;
assign v908aa8 = BtoS_ACK6_p & v910f82 | !BtoS_ACK6_p & v9079bf;
assign v930032 = jx0_p & v93fa7c | !jx0_p & v90d879;
assign v93fa22 = StoB_REQ8_p & v863aa0 | !StoB_REQ8_p & v903b1a;
assign v9081c2 = RtoB_ACK0_p & v844fcd | !RtoB_ACK0_p & !v844f91;
assign v8b4981 = jx2_p & v863b1a | !jx2_p & v90986f;
assign v904091 = jx3_p & v844f91 | !jx3_p & v93faf0;
assign v89f82d = BtoS_ACK1_p & v90e978 | !BtoS_ACK1_p & v9120f4;
assign v93fc28 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8b98bd;
assign v93fd97 = StoB_REQ9_p & v93e875 | !StoB_REQ9_p & v93e723;
assign v93fbe8 = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v906b71;
assign v93e781 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v909f7e;
assign v909995 = BtoS_ACK8_p & v93fbe4 | !BtoS_ACK8_p & v90944f;
assign v903b70 = BtoS_ACK7_p & v93fd79 | !BtoS_ACK7_p & v93f085;
assign v93ef5c = BtoS_ACK6_p & v87f17d | !BtoS_ACK6_p & v9093ec;
assign v90d546 = BtoS_ACK7_p & v907965 | !BtoS_ACK7_p & v93e791;
assign v93e4b4 = DEQ_p & v93e2a0 | !DEQ_p & v89f796;
assign v8b4a13 = jx1_p & v91ae94 | !jx1_p & v93fd8f;
assign v93f69e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fbde;
assign v905537 = jx0_p & v93e8de | !jx0_p & !v89c5e3;
assign v93fa08 = jx1_p & v90d52b | !jx1_p & v87f17d;
assign v904995 = StoB_REQ1_p & v90e251 | !StoB_REQ1_p & v906bf5;
assign v93fd48 = StoB_REQ7_p & v910527 | !StoB_REQ7_p & v93fce8;
assign v90844d = BtoS_ACK7_p & v911f15 | !BtoS_ACK7_p & v89e108;
assign v9090d1 = StoB_REQ7_p & v910710 | !StoB_REQ7_p & !v8d37bd;
assign v9055c0 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8f3869;
assign v91cfc7 = jx0_p & v93fe56 | !jx0_p & v9070e3;
assign v90da38 = DEQ_p & v889d4b | !DEQ_p & v909d4d;
assign v90523b = BtoS_ACK9_p & v9043fc | !BtoS_ACK9_p & v8b4a10;
assign v91db5a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v904a90;
assign v93fc32 = jx3_p & v908429 | !jx3_p & v9079ac;
assign v910f2e = jx1_p & v93fe68 | !jx1_p & !v93fada;
assign v91db5b = DEQ_p & v93f0b8 | !DEQ_p & v90f7a9;
assign v9078b3 = BtoS_ACK6_p & v90df7f | !BtoS_ACK6_p & v909eab;
assign v906657 = jx2_p & v93fcf7 | !jx2_p & v908322;
assign v908e7c = jx0_p & v904de5 | !jx0_p & v863b25;
assign v908af7 = StoB_REQ7_p & v93f7e3 | !StoB_REQ7_p & v93fd0e;
assign v93f223 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v89e121;
assign v9097bf = stateG7_1_p & v8b9ecf | !stateG7_1_p & v93f0a7;
assign v90a9c5 = jx0_p & v9071f0 | !jx0_p & v91026d;
assign v911880 = StoB_REQ7_p & v89f920 | !StoB_REQ7_p & v844f91;
assign v90d47d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b9ec9;
assign v93fbac = BtoS_ACK6_p & v8b9b9f | !BtoS_ACK6_p & v844f91;
assign v906f44 = StoB_REQ6_p & v93fe56 | !StoB_REQ6_p & v90856f;
assign v93f2a2 = StoB_REQ9_p & v93fdc9 | !StoB_REQ9_p & v909a70;
assign v93f8b5 = BtoS_ACK8_p & v93f7f8 | !BtoS_ACK8_p & v93eabc;
assign v907017 = StoB_REQ7_p & v8839a7 | !StoB_REQ7_p & v93fdd5;
assign v911815 = jx2_p & v93e385 | !jx2_p & v904221;
assign v93fc64 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v93e8d3;
assign v863a37 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v844f91;
assign v93f770 = jx1_p & v903d0c | !jx1_p & !v844f91;
assign v9075e7 = RtoB_ACK0_p & v904dc1 | !RtoB_ACK0_p & v9133ec;
assign v911944 = jx3_p & v90a629 | !jx3_p & v913632;
assign v91100a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8a8fac;
assign v904b1b = EMPTY_p & v93fd19 | !EMPTY_p & v91047b;
assign v8d37c1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v90810f;
assign v91146e = jx1_p & v905dd8 | !jx1_p & v91026f;
assign v93f6d5 = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v9051c9;
assign v911bc2 = BtoS_ACK0_p & v90534f | !BtoS_ACK0_p & v9089bf;
assign v90468e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90e3e1;
assign v90e019 = jx1_p & v907be9 | !jx1_p & v8b49f1;
assign v8d37d4 = BtoS_ACK8_p & v90f947 | !BtoS_ACK8_p & !v9071ed;
assign v93003e = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v90ee51;
assign v8f381b = BtoS_ACK6_p & v9068b7 | !BtoS_ACK6_p & v93fa04;
assign v93fe64 = jx0_p & v93fc4a | !jx0_p & v904f14;
assign v909d90 = RtoB_ACK0_p & v93f7ae | !RtoB_ACK0_p & v91a6e9;
assign v907206 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v905434;
assign v904bd4 = jx1_p & v93f223 | !jx1_p & !v90e3ed;
assign v93ec72 = jx1_p & v909187 | !jx1_p & !v93f91d;
assign v8b9d27 = jx0_p & v886f59 | !jx0_p & !v93fc7d;
assign v93f781 = DEQ_p & v9041a7 | !DEQ_p & v93fd3e;
assign v93f092 = jx1_p & v844f91 | !jx1_p & v9046de;
assign v90e926 = StoB_REQ9_p & v911cba | !StoB_REQ9_p & v90878b;
assign v913a6f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93f8a1;
assign v93df0a = ENQ_p & v844f91 | !ENQ_p & !v909bd3;
assign v90da41 = jx2_p & v93f744 | !jx2_p & v844f91;
assign v91107f = jx2_p & v90e1cf | !jx2_p & v90966d;
assign v93f9d5 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v93f652;
assign v89f894 = BtoS_ACK9_p & v93e136 | !BtoS_ACK9_p & v909365;
assign v905597 = jx0_p & v93fbe2 | !jx0_p & v910473;
assign v93fcda = BtoS_ACK6_p & v9096ae | !BtoS_ACK6_p & v87f17d;
assign v90e304 = BtoS_ACK6_p & v93fb3e | !BtoS_ACK6_p & v844f91;
assign v93f694 = jx1_p & v86f4a3 | !jx1_p & v844f91;
assign v844fbd = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844f91;
assign v93f6f9 = ENQ_p & v912477 | !ENQ_p & v912334;
assign v88bb45 = RtoB_ACK0_p & v9048c6 | !RtoB_ACK0_p & v9051ba;
assign v910d99 = BtoS_ACK7_p & v906ec1 | !BtoS_ACK7_p & v90e02c;
assign v903e7a = jx2_p & v87c51f | !jx2_p & !v909337;
assign v90f6b4 = RtoB_ACK0_p & v93fb72 | !RtoB_ACK0_p & v90828a;
assign v93f32b = StoB_REQ1_p & v906642 | !StoB_REQ1_p & !v908df7;
assign v90f0a8 = BtoS_ACK6_p & v90ad75 | !BtoS_ACK6_p & v93fd4e;
assign v93f896 = StoB_REQ9_p & v93ee39 | !StoB_REQ9_p & v90cee9;
assign v93f989 = BtoS_ACK6_p & v9058f3 | !BtoS_ACK6_p & v87f17d;
assign v93defa = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ee186;
assign v88c601 = StoB_REQ2_p & v908127 | !StoB_REQ2_p & v844f91;
assign v8ebd0e = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & !v904182;
assign jx1_n = !v8ee1f9;
assign v90eece = jx1_p & v93f111 | !jx1_p & !v9085fc;
assign v9300c6 = jx2_p & v91148d | !jx2_p & v8b4983;
assign v9093a9 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v90612e;
assign v9133d2 = BtoS_ACK0_p & v913348 | !BtoS_ACK0_p & v90575f;
assign v93e228 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v93f1b4;
assign v913a2b = BtoS_ACK1_p & v93deab | !BtoS_ACK1_p & v9063de;
assign v93f937 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & !v9046a7;
assign v93fdf0 = BtoS_ACK6_p & v8a8b0a | !BtoS_ACK6_p & v905425;
assign v90a5b8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v904088;
assign v93f1c4 = jx1_p & v91ae94 | !jx1_p & v90df4b;
assign v93fbde = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v90749b;
assign v93f6eb = jx0_p & v844f91 | !jx0_p & !v90cc30;
assign v93f6db = stateG12_p & v8a1fe3 | !stateG12_p & v93fa58;
assign v93fc45 = DEQ_p & v86e277 | !DEQ_p & v8b9cc5;
assign v90ad2f = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v93f765;
assign v8d37f5 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v909691;
assign v93f98d = ENQ_p & v908325 | !ENQ_p & v90a33f;
assign v903d01 = BtoS_ACK6_p & v90a216 | !BtoS_ACK6_p & !v93f92f;
assign v93f7bd = BtoS_ACK7_p & v93ea4f | !BtoS_ACK7_p & v93e77c;
assign v906a79 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v85eabe;
assign v90e261 = jx2_p & v863abb | !jx2_p & v844f91;
assign v9043f4 = BtoS_ACK6_p & v912679 | !BtoS_ACK6_p & v90ee37;
assign v8b98f4 = jx1_p & v93fd8b | !jx1_p & !v87a671;
assign v906315 = jx1_p & v910710 | !jx1_p & v93fcda;
assign v909dde = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v904628;
assign v9091dd = StoB_REQ9_p & v91364c | !StoB_REQ9_p & v93fdaa;
assign v8b9f38 = jx1_p & v93fc3e | !jx1_p & v908743;
assign v93f853 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v93e1dc;
assign v906cc7 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v907091;
assign v9058f3 = jx0_p & v844f91 | !jx0_p & !v844f9d;
assign v93f97c = StoB_REQ9_p & v911cba | !StoB_REQ9_p & v9093f3;
assign v90f7d1 = jx2_p & v93f743 | !jx2_p & v93ea3e;
assign v903cb1 = jx0_p & v90d6e8 | !jx0_p & !v93f6fc;
assign v909918 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8633ac;
assign v90460c = jx0_p & v844f91 | !jx0_p & !v85f258;
assign v90d59e = BtoS_ACK7_p & v93fd60 | !BtoS_ACK7_p & v903b68;
assign v911013 = jx3_p & v844f91 | !jx3_p & v93fa27;
assign v93fdbc = BtoS_ACK7_p & v912cf4 | !BtoS_ACK7_p & !v910515;
assign v93f6e5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v93e33e;
assign v908fb4 = StoB_REQ9_p & v87f17f | !StoB_REQ9_p & v93fd76;
assign v93fd89 = jx1_p & v884261 | !jx1_p & v93f889;
assign v93f045 = BtoS_ACK8_p & v904b00 | !BtoS_ACK8_p & v90638b;
assign v909b55 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v904436;
assign v93fd6d = jx1_p & v911edb | !jx1_p & v903f58;
assign v9053ed = DEQ_p & v9074f5 | !DEQ_p & v91a9a2;
assign v9067ab = BtoS_ACK8_p & v93f9bb | !BtoS_ACK8_p & !v87c4d2;
assign v90caf3 = jx1_p & v903d0c | !jx1_p & v930036;
assign v93fda4 = BtoS_ACK9_p & v93e3a1 | !BtoS_ACK9_p & v908acd;
assign v93f6bd = jx2_p & v9043fa | !jx2_p & v9074ce;
assign v910d10 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v93f32b;
assign v90d370 = BtoS_ACK8_p & v93fd76 | !BtoS_ACK8_p & v93f979;
assign v91a75e = jx0_p & v93f6dc | !jx0_p & v844f91;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v93f999 = RtoB_ACK0_p & v906c0c | !RtoB_ACK0_p & v905b81;
assign v93fc4d = StoB_REQ0_p & v9071c7 | !StoB_REQ0_p & v93fb45;
assign v90606d = BtoS_ACK6_p & v910243 | !BtoS_ACK6_p & !v93f8bb;
assign v90e8bf = jx1_p & v93fbac | !jx1_p & !v87b42f;
assign v907120 = EMPTY_p & v93df0a | !EMPTY_p & v90a5a4;
assign v905748 = BtoS_ACK7_p & v907580 | !BtoS_ACK7_p & v9089e7;
assign v93e00f = StoB_REQ4_p & v90f547 | !StoB_REQ4_p & v844f91;
assign v85eacb = StoB_REQ7_p & v93fd77 | !StoB_REQ7_p & v93f936;
assign v905b6a = jx3_p & v90de0e | !jx3_p & v844f91;
assign v91104c = StoB_REQ8_p & v906046 | !StoB_REQ8_p & v903da9;
assign v90cbfc = jx1_p & v844f91 | !jx1_p & v8ee1a3;
assign v93fac3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v91071c;
assign v93f80e = BtoS_ACK6_p & v8b9b9f | !BtoS_ACK6_p & v93fbdd;
assign v8b9b88 = BtoS_ACK9_p & v9050cc | !BtoS_ACK9_p & v9050ae;
assign v93f284 = ENQ_p & v93eed6 | !ENQ_p & v910543;
assign v93fa57 = BtoS_ACK8_p & v904bc1 | !BtoS_ACK8_p & v863a2d;
assign v913072 = StoB_REQ7_p & v910919 | !StoB_REQ7_p & v90eef9;
assign v89f830 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v91a7a3;
assign v9095e0 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v87a21f;
assign v90408b = jx1_p & v9074ce | !jx1_p & v906538;
assign v907168 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9d;
assign v8ebce4 = jx0_p & v93fa85 | !jx0_p & !v844f91;
assign v90ecfa = jx2_p & v87f17f | !jx2_p & v844f91;
assign v90fb82 = StoB_REQ7_p & v9121b6 | !StoB_REQ7_p & v844f91;
assign v87e7f5 = jx3_p & v93fbaf | !jx3_p & v93f15e;
assign v909dc5 = jx3_p & v93f78c | !jx3_p & !v9041e0;
assign v905a5b = jx3_p & v90f2f6 | !jx3_p & !v90a1fa;
assign v93fdac = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v91cc2d;
assign v93f64f = jx1_p & v9090d1 | !jx1_p & v909cf3;
assign v8b99b4 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v907122;
assign v85eadc = EMPTY_p & v909458 | !EMPTY_p & v93e3a5;
assign v909cf3 = StoB_REQ7_p & v93f9a4 | !StoB_REQ7_p & v90d442;
assign v905a12 = stateG12_p & v908325 | !stateG12_p & v93ebab;
assign v93f9a9 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v844f91;
assign v89fe59 = StoB_REQ3_p & v90f547 | !StoB_REQ3_p & v93fd2b;
assign v90a1c6 = stateG12_p & v8a1fe3 | !stateG12_p & v93fcdd;
assign v911428 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90a196;
assign v90f83e = StoB_REQ9_p & v911ebf | !StoB_REQ9_p & v909845;
assign v903db7 = BtoS_ACK9_p & v89f97d | !BtoS_ACK9_p & v93e996;
assign v90e361 = ENQ_p & v90adc4 | !ENQ_p & v911933;
assign v9045f0 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v91230c;
assign v93f833 = BtoS_ACK9_p & v907e81 | !BtoS_ACK9_p & v93fb77;
assign v93fb24 = BtoS_ACK6_p & v90ad75 | !BtoS_ACK6_p & !v9084ef;
assign v90921e = jx2_p & v93faad | !jx2_p & v93fb73;
assign v90d8d8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v912f40;
assign SLC1_n = v89f9e4;
assign v9085fc = jx0_p & v93e8de | !jx0_p & !v908eba;
assign v90a90b = jx1_p & v93f6ac | !jx1_p & !v90d47d;
assign v8b4990 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fc75;
assign v93f685 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v93e577;
assign v91a9b7 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93fba8;
assign v908cff = EMPTY_p & v909197 | !EMPTY_p & v93f9bf;
assign v859639 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v9117e5;
assign v904765 = BtoS_ACK0_p & v90810f | !BtoS_ACK0_p & !v93fb1a;
assign v85ea93 = BtoS_ACK7_p & v93e115 | !BtoS_ACK7_p & v905199;
assign v90f320 = BtoS_ACK1_p & v93deab | !BtoS_ACK1_p & v93f797;
assign v93fd57 = StoB_REQ1_p & v93e7d4 | !StoB_REQ1_p & v90d7e7;
assign v9118f0 = StoB_REQ7_p & v9114c0 | !StoB_REQ7_p & v93fd55;
assign v9099ef = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v904182;
assign v90ea21 = RtoB_ACK0_p & v8d37be | !RtoB_ACK0_p & v906fcc;
assign v93f9e7 = BtoS_ACK8_p & v93f770 | !BtoS_ACK8_p & !v93e816;
assign v90d1c9 = EMPTY_p & v93eadd | !EMPTY_p & v93f0c0;
assign v93fd01 = BtoS_ACK8_p & v909367 | !BtoS_ACK8_p & !v904abd;
assign v903cef = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v9051cd;
assign v93f8ec = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v93fd01;
assign v904590 = stateG12_p & v9109e6 | !stateG12_p & v90656f;
assign v908138 = BtoS_ACK7_p & v90d3ff | !BtoS_ACK7_p & v91137e;
assign v93f646 = BtoS_ACK8_p & v909366 | !BtoS_ACK8_p & !v906d77;
assign v913449 = BtoS_ACK8_p & v93ecc4 | !BtoS_ACK8_p & v904753;
assign v90a2bd = StoB_REQ8_p & v93dbe9 | !StoB_REQ8_p & v904a80;
assign v93fde5 = jx1_p & v93f8f0 | !jx1_p & v844f91;
assign v8f382e = BtoS_ACK6_p & v909f04 | !BtoS_ACK6_p & v93f2dc;
assign v903ba1 = BtoS_ACK1_p & v93deab | !BtoS_ACK1_p & v903fa0;
assign v90432c = BtoS_ACK6_p & v93fc0a | !BtoS_ACK6_p & v90ff47;
assign v9063d8 = BtoS_ACK8_p & v93fde7 | !BtoS_ACK8_p & !v844fa5;
assign v93f753 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & !v844fc1;
assign v906541 = jx2_p & v89f9c3 | !jx2_p & v93eb22;
assign v908834 = BtoS_ACK1_p & v90fc92 | !BtoS_ACK1_p & v872e32;
assign v90a36a = BtoS_ACK8_p & v906b5f | !BtoS_ACK8_p & !v93fc98;
assign v93fa64 = DEQ_p & v93fc76 | !DEQ_p & v907494;
assign v90a9cc = BtoS_ACK9_p & v90fe55 | !BtoS_ACK9_p & v908176;
assign v90ee51 = BtoS_ACK7_p & v9096f0 | !BtoS_ACK7_p & !v90d52b;
assign v93f216 = jx1_p & v91ae94 | !jx1_p & v93fb29;
assign v85eb17 = BtoS_ACK8_p & v9095b9 | !BtoS_ACK8_p & v912178;
assign v8714f5 = StoB_REQ3_p & v93fd9b | !StoB_REQ3_p & !v904182;
assign v90dd28 = jx2_p & v905f25 | !jx2_p & v93fcba;
assign v93f6f0 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v93ecd6;
assign v9063de = StoB_REQ1_p & v904436 | !StoB_REQ1_p & v87c9b1;
assign v90caed = jx1_p & v93e0b5 | !jx1_p & v93fb3a;
assign v90dca4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9051f4;
assign v930106 = BtoS_ACK7_p & v93fc5d | !BtoS_ACK7_p & v90789d;
assign v907f25 = jx2_p & v93fb53 | !jx2_p & v844f91;
assign v93f908 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v88c601;
assign v93e27a = jx2_p & v863a38 | !jx2_p & v844f91;
assign v93fcc1 = jx1_p & v8b9eca | !jx1_p & v844f91;
assign v844fb5 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v93f320 = jx2_p & v907018 | !jx2_p & !v93fb9d;
assign v880d7e = jx0_p & v9096f7 | !jx0_p & v93eceb;
assign v93f7b7 = BtoS_ACK0_p & v9046a6 | !BtoS_ACK0_p & v93e404;
assign v93f747 = BtoS_ACK6_p & v9099fa | !BtoS_ACK6_p & v93f28a;
assign v90d7cb = StoB_REQ8_p & v910c5b | !StoB_REQ8_p & v905748;
assign v9135f1 = jx3_p & v844f91 | !jx3_p & v93f833;
assign v90f8c2 = StoB_REQ2_p & v93ed70 | !StoB_REQ2_p & v90e2dc;
assign v9070e3 = BtoS_ACK0_p & v9047b7 | !BtoS_ACK0_p & !v90a91e;
assign v9109e5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v908546;
assign v90dc28 = StoB_REQ1_p & v93f9e8 | !StoB_REQ1_p & v8858ac;
assign v911b78 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v93dc30;
assign v908797 = jx0_p & v906d08 | !jx0_p & !v844f91;
assign v93f8bb = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v90569e;
assign v911ed7 = StoB_REQ7_p & v93ee3b | !StoB_REQ7_p & v85de34;
assign v91a6d1 = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v89e097;
assign v93fdb6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91024c;
assign v90549c = BtoS_ACK0_p & v906627 | !BtoS_ACK0_p & v909dcc;
assign v9114c0 = BtoS_ACK6_p & v912679 | !BtoS_ACK6_p & v87f17d;
assign v93f6a9 = EMPTY_p & v909924 | !EMPTY_p & !v90500e;
assign v912f4e = jx1_p & v9095bf | !jx1_p & !v910230;
assign v9121b6 = BtoS_ACK6_p & v910243 | !BtoS_ACK6_p & v90569e;
assign v9099fa = jx0_p & v89e097 | !jx0_p & v844f91;
assign v93fdda = BtoS_ACK9_p & v907e3f | !BtoS_ACK9_p & v903c0d;
assign v93fafe = jx1_p & v911edb | !jx1_p & v908ee8;
assign v91a6f7 = StoB_REQ0_p & v909b55 | !StoB_REQ0_p & v913a2b;
assign v90856f = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v8ee1f5;
assign v910f5a = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v903bb1;
assign v8728ef = jx2_p & v93fa73 | !jx2_p & v93fcf2;
assign v91155d = BtoS_ACK9_p & v93fcd6 | !BtoS_ACK9_p & v9131d1;
assign v90541b = jx2_p & v93fda8 | !jx2_p & !v844f91;
assign v92ffd9 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v90a8cd;
assign v90d93b = jx1_p & v93fbe5 | !jx1_p & !v904a61;
assign v93fa3a = BtoS_ACK9_p & v904e2f | !BtoS_ACK9_p & v89e08c;
assign v910f1b = BtoS_ACK1_p & v913348 | !BtoS_ACK1_p & v907bee;
assign v90944d = BtoS_ACK7_p & v90f575 | !BtoS_ACK7_p & v90dcc6;
assign v9052ef = jx0_p & v90ea74 | !jx0_p & v93fdfa;
assign v906d80 = jx3_p & v844f91 | !jx3_p & v908ff3;
assign v8a9250 = stateG7_1_p & v90ed7e | !stateG7_1_p & v93f6d0;
assign v90f547 = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & v844fbb;
assign v90810f = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v90534f;
assign v90444d = ENQ_p & v93fdf6 | !ENQ_p & v8baf9a;
assign v8b9e3d = BtoS_ACK0_p & v9062d9 | !BtoS_ACK0_p & v9300cb;
assign v93fd17 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a112;
assign v93dbaa = jx1_p & v904bf3 | !jx1_p & v9058f3;
assign v9051f4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86e831;
assign v90557c = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v90a799;
assign v93000b = jx0_p & v93f723 | !jx0_p & !v93f707;
assign v9114c9 = jx2_p & v93ec72 | !jx2_p & !v8f60f9;
assign v90a1fa = BtoS_ACK9_p & v8f3825 | !BtoS_ACK9_p & v8739eb;
assign v904adb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v844f99;
assign v93fa82 = jx2_p & v93eeda | !jx2_p & !v93f81e;
assign v909d4d = RtoB_ACK0_p & v909dec | !RtoB_ACK0_p & v93fe11;
assign v90fbfe = BtoS_ACK8_p & v93fc5d | !BtoS_ACK8_p & v912673;
assign v93daaf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910117;
assign v9082e6 = stateG7_1_p & v90505e | !stateG7_1_p & v87261e;
assign v90d442 = BtoS_ACK6_p & v905537 | !BtoS_ACK6_p & v904e47;
assign v93fbb1 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v906327;
assign v8a9209 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90526b;
assign v904313 = StoB_REQ3_p & v905702 | !StoB_REQ3_p & v90decf;
assign v93f77c = StoB_REQ9_p & v86d7d1 | !StoB_REQ9_p & v90a0b5;
assign v93f2a8 = jx1_p & v93f9af | !jx1_p & !v9085fc;
assign v89f966 = ENQ_p & v93f893 | !ENQ_p & v909347;
assign v90776b = jx2_p & v9097c3 | !jx2_p & v93faf8;
assign v90531e = BtoS_ACK6_p & v93f63b | !BtoS_ACK6_p & v9051d8;
assign v93e189 = jx3_p & v93fdda | !jx3_p & v844f91;
assign v85f28b = jx3_p & v93fd59 | !jx3_p & !v93faca;
assign v86ce77 = StoB_REQ8_p & v904b00 | !StoB_REQ8_p & v907a2f;
assign v8f22a2 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v90e000;
assign v9093d9 = jx3_p & v93fe39 | !jx3_p & v93eed6;
assign v93f82f = BtoS_ACK9_p & v907bfd | !BtoS_ACK9_p & v90d4c9;
assign v911bcf = jx3_p & v91aa04 | !jx3_p & v844f91;
assign v93f119 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fc0a;
assign v906c8c = BtoS_ACK0_p & v911102 | !BtoS_ACK0_p & v93e78b;
assign v89b1a4 = BtoR_REQ1_p & v8b9bbf | !BtoR_REQ1_p & v90ef0d;
assign v858fc9 = jx1_p & v93fc3e | !jx1_p & v9087d1;
assign v8f22ad = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fc4c;
assign v909180 = StoB_REQ6_p & v90690e | !StoB_REQ6_p & v89e0c5;
assign v91195c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a924b;
assign v93e9ea = BtoS_ACK6_p & v93fb41 | !BtoS_ACK6_p & v911b50;
assign v93fc9a = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v911c50;
assign v93fdcb = jx0_p & v910b0e | !jx0_p & v90762a;
assign v904753 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fd63;
assign v93f709 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93e577;
assign v906e04 = jx2_p & v93e610 | !jx2_p & v93fd89;
assign v93db85 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v9088ff;
assign v910b96 = jx1_p & v909ba1 | !jx1_p & v9122e7;
assign v93e2c2 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v90e978;
assign v91a799 = jx2_p & v89e0a6 | !jx2_p & v844f91;
assign v9085ac = jx1_p & v844f91 | !jx1_p & v93e51c;
assign v910545 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v908fe9;
assign v93f6f3 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v911833;
assign v93f8cf = jx0_p & v913435 | !jx0_p & v93fb3e;
assign v903c1c = BtoS_ACK6_p & v90860a | !BtoS_ACK6_p & v90aa76;
assign v910e55 = jx3_p & v844f91 | !jx3_p & v90ecfa;
assign v93df9f = ENQ_p & v93f59b | !ENQ_p & v89b0e5;
assign v90d9b2 = jx1_p & v90accf | !jx1_p & v904568;
assign v903aff = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v906ad1;
assign v90d5a3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v910bb8;
assign v93e602 = StoB_REQ1_p & v906642 | !StoB_REQ1_p & !v844f91;
assign v93f826 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90460e;
assign v93f8ae = jx0_p & v93f470 | !jx0_p & v844f91;
assign v93eb13 = BtoS_ACK6_p & v903c83 | !BtoS_ACK6_p & v904f5c;
assign v8b5ff8 = BtoS_ACK8_p & v85eaf3 | !BtoS_ACK8_p & v9111a4;
assign v9041fc = BtoS_ACK6_p & v9068b7 | !BtoS_ACK6_p & v93f68b;
assign v93f69b = jx0_p & v844f91 | !jx0_p & v90f2ff;
assign v9057fa = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v908a3d;
assign v907a33 = jx1_p & v911fc7 | !jx1_p & !v844fbd;
assign v90a86b = StoB_REQ0_p & v910bd7 | !StoB_REQ0_p & !v90501e;
assign v93f88f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fc9a;
assign v89f8a9 = BtoS_ACK8_p & v93e007 | !BtoS_ACK8_p & v93f97d;
assign v90efe2 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v904f1a;
assign v91a762 = BtoS_ACK8_p & v90a733 | !BtoS_ACK8_p & v904c72;
assign v8807b1 = jx1_p & v844f91 | !jx1_p & v93f037;
assign v90767c = RtoB_ACK1_p & v90a541 | !RtoB_ACK1_p & v911a92;
assign v90443a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v906642;
assign v89e0c5 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v9124a6;
assign v93fd75 = jx1_p & v904628 | !jx1_p & v844f91;
assign v85eaff = jx3_p & v93f107 | !jx3_p & v90adc4;
assign v905aaa = jx1_p & v9040a9 | !jx1_p & !v9117db;
assign v93fb96 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v904eba;
assign v93e77b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v844f99;
assign v844f91 = 1;
assign v844fbb = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & !v844f91;
assign v93db4a = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v911680;
assign v909d18 = BtoS_ACK0_p & v90deff | !BtoS_ACK0_p & v93ec26;
assign v905d37 = StoB_REQ2_p & v87b4fc | !StoB_REQ2_p & v911d61;
assign v93f844 = EMPTY_p & v909dec | !EMPTY_p & v912172;
assign v85f278 = BtoS_ACK8_p & v863b34 | !BtoS_ACK8_p & v91080f;
assign v904757 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93f6a7;
assign v906046 = jx2_p & v90adcb | !jx2_p & v844f91;
assign v91080c = jx1_p & v913435 | !jx1_p & v93f7ac;
assign v93ecb0 = jx2_p & v93fafe | !jx2_p & v8b4983;
assign v93f6c1 = BtoS_ACK8_p & v93db1d | !BtoS_ACK8_p & v930099;
assign v90ae5a = BtoS_ACK0_p & v9046a6 | !BtoS_ACK0_p & v93fcc5;
assign v90e841 = BtoS_ACK6_p & v88932d | !BtoS_ACK6_p & v9132d2;
assign v930097 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93fc29;
assign v90d84e = jx0_p & v90aeb7 | !jx0_p & v85f258;
assign v905312 = jx3_p & v93fa7d | !jx3_p & !v93fbb1;
assign v907634 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v909353;
assign v905a9e = BtoS_ACK7_p & v93dbf1 | !BtoS_ACK7_p & v91dc98;
assign v91325f = BtoS_ACK0_p & v93ea50 | !BtoS_ACK0_p & v906d2b;
assign v9097c6 = jx1_p & v90f07f | !jx1_p & v90d7a0;
assign v9115cb = jx3_p & v90a9fc | !jx3_p & v93f2b9;
assign v9047b1 = RtoB_ACK0_p & v91a9a2 | !RtoB_ACK0_p & v90a241;
assign v93fc49 = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v90f0a1;
assign v9134fe = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93e148;
assign v9117e2 = jx3_p & v8b9e71 | !jx3_p & v93e31b;
assign v8f223b = BtoS_ACK7_p & v906d2a | !BtoS_ACK7_p & v90caed;
assign v9043c2 = BtoS_ACK7_p & v93dbe9 | !BtoS_ACK7_p & v93f735;
assign v908e73 = BtoS_ACK6_p & v90a216 | !BtoS_ACK6_p & !v93fcb9;
assign v8ee186 = BtoS_ACK6_p & v906c35 | !BtoS_ACK6_p & v905204;
assign v8f22ce = BtoS_ACK6_p & v912679 | !BtoS_ACK6_p & v9132d2;
assign v93f9d2 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v909691;
assign v90789d = jx2_p & v93f687 | !jx2_p & v906534;
assign v93fd8b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v904ab2;
assign v90a216 = jx0_p & v93f762 | !jx0_p & !v93fc0a;
assign v910919 = jx0_p & v90eef9 | !jx0_p & v844f91;
assign v93f86a = StoB_REQ8_p & v93fd78 | !StoB_REQ8_p & v93fc07;
assign v90d7e7 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v905702;
assign v93f7e6 = BtoS_ACK9_p & v93fa54 | !BtoS_ACK9_p & !v90470d;
assign v90fa5e = jx0_p & v93f87f | !jx0_p & !v93fdac;
assign v911d8e = jx0_p & v93f689 | !jx0_p & v906a79;
assign v93fda7 = jx1_p & v913332 | !jx1_p & v8848d6;
assign v905146 = BtoR_REQ0_p & v90467c | !BtoR_REQ0_p & v908cff;
assign v93fa1f = jx1_p & v93fbe5 | !jx1_p & v93ee3b;
assign v90d217 = jx0_p & v93f689 | !jx0_p & !v910056;
assign v93fa69 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93f85b;
assign v93f690 = BtoS_ACK7_p & v93fc5d | !BtoS_ACK7_p & v93f541;
assign v863aee = StoB_REQ8_p & v9088bc | !StoB_REQ8_p & v9045f0;
assign v90ed77 = BtoS_ACK9_p & v90fe55 | !BtoS_ACK9_p & v93f7ec;
assign v90e9f7 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v9088bc;
assign v909289 = BtoS_ACK7_p & v93f04f | !BtoS_ACK7_p & !v93fbfe;
assign v93e975 = jx1_p & v90fb82 | !jx1_p & v93fce3;
assign v93e723 = BtoS_ACK8_p & v90512d | !BtoS_ACK8_p & v93fb7d;
assign v93fccd = StoB_REQ9_p & v93f291 | !StoB_REQ9_p & v9133dc;
assign v93fd87 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v905660;
assign v93f12b = StoB_REQ7_p & v9041e6 | !StoB_REQ7_p & v911c11;
assign v908eea = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v904182;
assign v93f52d = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v90a20a;
assign v93fa93 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v863aee;
assign v93fe0c = jx0_p & v90f66c | !jx0_p & v844f91;
assign v93fa95 = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v844f91;
assign v90e7e2 = EMPTY_p & v89e0d5 | !EMPTY_p & v93fa64;
assign v90729e = BtoS_ACK7_p & v91003b | !BtoS_ACK7_p & v906dd6;
assign v93e440 = jx3_p & v844f91 | !jx3_p & v93f87c;
assign v93f6fc = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v909297 = StoB_REQ7_p & v910710 | !StoB_REQ7_p & !v93fc19;
assign v93f0b8 = RtoB_ACK0_p & v904c53 | !RtoB_ACK0_p & v90fa88;
assign v93e933 = StoB_REQ6_p & v8d37c1 | !StoB_REQ6_p & v93fc0a;
assign v90738c = ENQ_p & v904f0d | !ENQ_p & v93fe44;
assign v90d972 = BtoS_ACK7_p & v90893a | !BtoS_ACK7_p & v93fc3e;
assign v93e68d = jx2_p & v910e2d | !jx2_p & v93dc15;
assign v93f8f0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844fa1;
assign v87c4ee = jx3_p & v93f334 | !jx3_p & v89e0fb;
assign v93e9e3 = BtoS_ACK0_p & v86e433 | !BtoS_ACK0_p & v93f6df;
assign v91026d = BtoS_ACK0_p & v913348 | !BtoS_ACK0_p & v904258;
assign v93e262 = ENQ_p & v93f753 | !ENQ_p & !v91343f;
assign v9083b1 = stateG7_1_p & v93f882 | !stateG7_1_p & v904e93;
assign v909dec = ENQ_p & v93f89f | !ENQ_p & v844f91;
assign v8b9c3a = StoB_REQ9_p & v93fe0a | !StoB_REQ9_p & v91334f;
assign v9098ba = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v904b58;
assign v90d789 = StoB_REQ0_p & v909cc1 | !StoB_REQ0_p & v93e781;
assign v93fa53 = StoB_REQ7_p & v8a9289 | !StoB_REQ7_p & v8b9d0f;
assign v90e315 = jx3_p & v90d7e8 | !jx3_p & v910d4a;
assign v90854b = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v91058e;
assign v909ea8 = StoB_REQ1_p & v93f908 | !StoB_REQ1_p & v905285;
assign v904886 = BtoS_ACK7_p & v90d879 | !BtoS_ACK7_p & v906dd6;
assign v904abe = jx1_p & v844f91 | !jx1_p & v909c45;
assign v86e7cf = DEQ_p & v844f91 | !DEQ_p & !v844fa9;
assign v9050ad = RtoB_ACK1_p & v93e230 | !RtoB_ACK1_p & v907916;
assign v909823 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9096a3;
assign v90a5ee = jx1_p & v844f91 | !jx1_p & !v93f8a6;
assign v93fc6d = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v909367;
assign v93ec24 = StoB_REQ9_p & v93fded | !StoB_REQ9_p & v8b9d28;
assign v93e136 = StoB_REQ8_p & v90f947 | !StoB_REQ8_p & v905e43;
assign v904ebe = BtoS_ACK9_p & v93f074 | !BtoS_ACK9_p & v90e1c3;
assign v90f2de = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v90474e;
assign v9095b9 = jx2_p & v93f8e2 | !jx2_p & v844f91;
assign v909c72 = BtoS_ACK8_p & v93f1b4 | !BtoS_ACK8_p & !v908f85;
assign v93f769 = BtoS_ACK7_p & v93f955 | !BtoS_ACK7_p & v93ecb9;
assign v93f779 = BtoS_ACK6_p & v90cc30 | !BtoS_ACK6_p & v93fd4e;
assign v904d89 = jx2_p & v93f7f6 | !jx2_p & v9087d2;
assign v930036 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v910230;
assign v93fcd4 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90db9f;
assign v93f7c4 = BtoS_ACK0_p & v913561 | !BtoS_ACK0_p & v91137c;
assign v90df5b = BtoS_ACK0_p & v93fc02 | !BtoS_ACK0_p & v905556;
assign v93fa3f = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v907717;
assign v91043e = StoB_REQ1_p & v90631b | !StoB_REQ1_p & v844f91;
assign v90a8e9 = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v8f22ea;
assign v906495 = StoB_REQ7_p & v93fdf0 | !StoB_REQ7_p & v906cf5;
assign v90e437 = FULL_p & v90ad6f | !FULL_p & v90a2f1;
assign v93f78c = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v87ca35;
assign v93f795 = BtoS_ACK7_p & v93f6bd | !BtoS_ACK7_p & v93fd07;
assign v93dfc2 = BtoS_ACK9_p & v89e10d | !BtoS_ACK9_p & v87ca35;
assign v9050e7 = BtoS_ACK7_p & v93e10c | !BtoS_ACK7_p & !v93f9f0;
assign v90962d = StoB_REQ6_p & v910243 | !StoB_REQ6_p & v844f91;
assign v8b6034 = BtoR_REQ1_p & v90767c | !BtoR_REQ1_p & v93f6b6;
assign v90ba1a = StoB_REQ8_p & v871b18 | !StoB_REQ8_p & v93f98c;
assign v8fe223 = StoB_REQ0_p & v909525 | !StoB_REQ0_p & v93fae4;
assign v911b48 = StoB_REQ8_p & v905325 | !StoB_REQ8_p & v90a1bc;
assign v90eef9 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v90cc30;
assign v90e02c = jx2_p & v93fb81 | !jx2_p & !v907f31;
assign v93fb78 = jx2_p & v90fae7 | !jx2_p & v844f91;
assign v90ad6c = BtoS_ACK1_p & v86c2d0 | !BtoS_ACK1_p & v90dd1f;
assign v9048d7 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v90f547;
assign v93fac6 = StoB_REQ7_p & v93fc2b | !StoB_REQ7_p & v844f91;
assign v9058f4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93fe5b;
assign v87cb21 = BtoR_REQ1_p & v90859f | !BtoR_REQ1_p & v910f41;
assign v905ff9 = jx2_p & v93dbaa | !jx2_p & v844f91;
assign v9079bf = jx0_p & v90ad39 | !jx0_p & v844f91;
assign v93fe5f = BtoS_ACK8_p & v909fb2 | !BtoS_ACK8_p & v93fd54;
assign v906983 = jx2_p & v93fa4e | !jx2_p & v86f5de;
assign v90cc41 = BtoS_ACK0_p & v906255 | !BtoS_ACK0_p & v9097b1;
assign v912679 = jx0_p & v93fdfb | !jx0_p & !v844f95;
assign v90a541 = EMPTY_p & v910e44 | !EMPTY_p & v90e073;
assign v904ae8 = jx0_p & v913435 | !jx0_p & v9091b2;
assign v9126b6 = StoB_REQ7_p & v910710 | !StoB_REQ7_p & v909ab9;
assign v906bf5 = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & v90604e;
assign v87ca92 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93f9b9;
assign v9077c7 = ENQ_p & v93eed6 | !ENQ_p & v9115cb;
assign v90828a = FULL_p & v93dfb4 | !FULL_p & v908751;
assign v90469d = EMPTY_p & v86341e | !EMPTY_p & v8a8fa3;
assign v9123a2 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9f;
assign v909cb1 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844fbb;
assign v90fb0e = jx1_p & v908aa8 | !jx1_p & v844f91;
assign v910c0f = stateG7_1_p & v844f91 | !stateG7_1_p & v909bff;
assign v93fbf0 = BtoS_ACK6_p & v904e70 | !BtoS_ACK6_p & v90add3;
assign v90aeb8 = stateG12_p & v90fbad | !stateG12_p & v904303;
assign v93fa06 = DEQ_p & v90fa88 | !DEQ_p & v906769;
assign v907b65 = jx0_p & v93f511 | !jx0_p & !v91194f;
assign v909661 = jx1_p & v9055bd | !jx1_p & v908107;
assign v8a8fdd = jx1_p & v9082a3 | !jx1_p & v93ee4b;
assign v8b9e73 = DEQ_p & v905d92 | !DEQ_p & v90f6b4;
assign v93fe31 = jx0_p & v844f9f | !jx0_p & !v908e7e;
assign v90484c = BtoS_ACK2_p & v9076a8 | !BtoS_ACK2_p & v908681;
assign v904c80 = jx2_p & v93fb81 | !jx2_p & !v844f91;
assign v904d38 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86346f;
assign v91336c = StoB_REQ8_p & v90728a | !StoB_REQ8_p & v93ed29;
assign v90ae6a = jx0_p & v910bf8 | !jx0_p & v93fd21;
assign v87ca8a = BtoS_ACK6_p & v91a9b9 | !BtoS_ACK6_p & v9044a5;
assign v909dcc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f6dd;
assign v913265 = StoB_REQ8_p & v9088bc | !StoB_REQ8_p & v9098a3;
assign v912405 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v90faf9;
assign v93f7a8 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v904886;
assign v93fafd = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v907aa0;
assign v908127 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v904182;
assign v90d6ef = StoB_REQ8_p & v911552 | !StoB_REQ8_p & v903fac;
assign v91aa51 = jx0_p & v86ccf1 | !jx0_p & v90ad77;
assign v904663 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9098ba;
assign v93fa4d = BtoS_ACK7_p & v93e259 | !BtoS_ACK7_p & v887a80;
assign v93f8f7 = BtoS_ACK1_p & v8bb868 | !BtoS_ACK1_p & v93fd5b;
assign v90539f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91a9b4;
assign v93f0c0 = DEQ_p & v889d4b | !DEQ_p & v905b81;
assign v90deaa = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844fbb;
assign v93fd5b = StoB_REQ1_p & v93e7d4 | !StoB_REQ1_p & v906c6f;
assign v85ea76 = jx0_p & v906af3 | !jx0_p & v93f6e5;
assign v9045b2 = jx1_p & v93debb | !jx1_p & v87f17d;
assign v910e69 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v90a233;
assign v89e0d7 = StoB_REQ9_p & v911ebf | !StoB_REQ9_p & v9043a5;
assign v93fb80 = BtoR_REQ0_p & v910d62 | !BtoR_REQ0_p & v91a6dc;
assign v93e548 = RtoB_ACK0_p & v9103e5 | !RtoB_ACK0_p & v863a00;
assign v85eabe = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v906642;
assign v93f722 = jx0_p & v93f714 | !jx0_p & !v93f6fc;
assign v903f21 = BtoS_ACK1_p & v93f85e | !BtoS_ACK1_p & v904fc8;
assign v93dee0 = jx1_p & v8f22d1 | !jx1_p & !v93e60f;
assign v909224 = jx1_p & v844f91 | !jx1_p & !v93f70d;
assign v93fcc5 = StoB_REQ0_p & v9071c7 | !StoB_REQ0_p & v91305d;
assign v91aa45 = StoB_REQ8_p & v93e27a | !StoB_REQ8_p & v93db1d;
assign v881ec0 = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v9098bb;
assign v90897e = BtoS_ACK7_p & v908073 | !BtoS_ACK7_p & !v909e28;
assign v89f9bc = BtoS_ACK0_p & v8bb868 | !BtoS_ACK0_p & v905803;
assign v903c80 = StoB_REQ8_p & v89f905 | !StoB_REQ8_p & v87c4c5;
assign v90cbcc = BtoS_ACK6_p & v9099fa | !BtoS_ACK6_p & v93f8ae;
assign v90ff49 = ENQ_p & v912477 | !ENQ_p & v93facc;
assign v90e000 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90e6b0;
assign v903d1e = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v9078da;
assign v90eaad = jx1_p & v9043ec | !jx1_p & !v904ccb;
assign v903b68 = jx1_p & v907be9 | !jx1_p & v844f91;
assign v880d77 = RtoB_ACK0_p & v93fde2 | !RtoB_ACK0_p & v93f4ac;
assign v93fc42 = EMPTY_p & v90ad6f | !EMPTY_p & v9135e9;
assign v90fb54 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fc3d;
assign v90ec4b = jx3_p & v844f91 | !jx3_p & v9081ef;
assign v90ef16 = jx1_p & v93db85 | !jx1_p & !v844f91;
assign v87ec92 = stateG12_p & v93f89f | !stateG12_p & v904fb4;
assign v90ecba = jx1_p & v93ecc4 | !jx1_p & v93f72f;
assign v93e94e = DEQ_p & v93e731 | !DEQ_p & v92ffd6;
assign v93fde7 = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & v844f91;
assign v93f6ca = jx0_p & v90515d | !jx0_p & v8b49ad;
assign v90831e = DEQ_p & v88bb45 | !DEQ_p & v9051ba;
assign v93e1dc = StoB_REQ1_p & v907468 | !StoB_REQ1_p & v844f91;
assign v910527 = jx0_p & v93f119 | !jx0_p & !v844f91;
assign v90ebde = BtoS_ACK6_p & v871df8 | !BtoS_ACK6_p & v93fe5c;
assign v871b18 = jx1_p & v93e819 | !jx1_p & v903fef;
assign v93f9f5 = EMPTY_p & v9082be | !EMPTY_p & v911586;
assign v909f36 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93e450;
assign v93e269 = StoB_REQ9_p & v903c0d | !StoB_REQ9_p & v9090d6;
assign v910e84 = jx1_p & v93e6af | !jx1_p & v844f91;
assign v93f093 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v904931;
assign v93fce1 = jx0_p & v909157 | !jx0_p & v90491c;
assign v93fcb4 = jx2_p & v9104aa | !jx2_p & v93fb20;
assign v93f362 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v90999b;
assign v8b9bbf = RtoB_ACK1_p & v90583b | !RtoB_ACK1_p & v93f6c4;
assign v906ce1 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v844fbf;
assign v904736 = StoB_REQ6_p & v909adc | !StoB_REQ6_p & v8b9e40;
assign v905d2c = BtoS_ACK7_p & v93e259 | !BtoS_ACK7_p & v90fbfd;
assign v93fb05 = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v904d75;
assign v93f90f = jx3_p & v93fbcc | !jx3_p & v844f91;
assign v9086b7 = StoB_REQ7_p & v93f0a3 | !StoB_REQ7_p & v9098ab;
assign v90a1bc = BtoS_ACK7_p & v90891d | !BtoS_ACK7_p & v93eaca;
assign v90adcb = jx1_p & v9093ec | !jx1_p & v844f91;
assign v9056a4 = StoB_REQ8_p & v907e81 | !StoB_REQ8_p & v93f279;
assign v906b4a = BtoS_ACK9_p & v8633ec | !BtoS_ACK9_p & v93fa69;
assign v90d21a = BtoS_ACK0_p & v93fe07 | !BtoS_ACK0_p & v910e17;
assign v93fb9c = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v93e00f;
assign v90d7a0 = BtoS_ACK6_p & v93e89f | !BtoS_ACK6_p & v9121a7;
assign v89f84e = jx0_p & v844f91 | !jx0_p & v93fa7c;
assign v9078a1 = BtoS_ACK8_p & v93fdd9 | !BtoS_ACK8_p & !v86fef2;
assign v90467c = EMPTY_p & v909197 | !EMPTY_p & v90831e;
assign v93e9ce = StoB_REQ0_p & v93db4a | !StoB_REQ0_p & v93fdaf;
assign v93fc1d = jx3_p & v908e4b | !jx3_p & v93f82f;
assign v90fc87 = jx1_p & v906fbf | !jx1_p & v90a786;
assign v8b9c01 = jx3_p & v93e0c9 | !jx3_p & v844f91;
assign v90da35 = StoB_REQ8_p & v907469 | !StoB_REQ8_p & v908a35;
assign v90fc7f = BtoS_ACK6_p & v93f6ca | !BtoS_ACK6_p & v93fa1b;
assign v93fe71 = StoB_REQ3_p & v87c533 | !StoB_REQ3_p & v93fbd3;
assign v909dc9 = RtoB_ACK1_p & v904253 | !RtoB_ACK1_p & v909a08;
assign v93fcb9 = jx0_p & v87c55f | !jx0_p & !v87bf0e;
assign v85e142 = jx1_p & v9115a7 | !jx1_p & v88b606;
assign v88b26d = RtoB_ACK0_p & v93f98d | !RtoB_ACK0_p & v93f7e1;
assign v90e62f = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v910c20;
assign v904610 = StoB_REQ8_p & v913428 | !StoB_REQ8_p & v90e6f8;
assign v93fbcf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90636b;
assign v90ea51 = StoB_REQ8_p & v90722c | !StoB_REQ8_p & v9117b1;
assign v93fc8d = BtoS_ACK6_p & v8b9b9f | !BtoS_ACK6_p & v93fd14;
assign DEQ_n = !v8c8823;
assign v9078f8 = jx3_p & v93fa7d | !jx3_p & !v911150;
assign v93ed91 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fccb;
assign v93fde4 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v90a3e0;
assign v93fdfd = jx1_p & v90531e | !jx1_p & v90e433;
assign v90e76a = jx0_p & v93f714 | !jx0_p & v844f91;
assign v9042b8 = jx1_p & v90accf | !jx1_p & v8f3865;
assign v91137c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9107ca;
assign v912190 = StoB_REQ8_p & v93fbb6 | !StoB_REQ8_p & !v908fb5;
assign v910dfa = StoB_REQ9_p & v93e27a | !StoB_REQ9_p & v93e915;
assign v89e0b4 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8f3853;
assign v93f6a6 = StoB_REQ8_p & v91071f | !StoB_REQ8_p & v905d2c;
assign v93fe29 = jx2_p & v911db6 | !jx2_p & v87f17d;
assign v93e4f9 = BtoS_ACK9_p & v90fe55 | !BtoS_ACK9_p & v90dcfa;
assign v90ea1f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90995e;
assign v89c5e3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v913619;
assign v8ee1a7 = BtoS_ACK7_p & v911185 | !BtoS_ACK7_p & !v90a1db;
assign v908681 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b9dfa;
assign v90e774 = EMPTY_p & v91a9a2 | !EMPTY_p & v93fa5e;
assign v91007d = EMPTY_p & v90ad6f | !EMPTY_p & v90e5b9;
assign v93fbce = BtoR_REQ0_p & v903d68 | !BtoR_REQ0_p & v87c9b3;
assign v89fe24 = StoB_REQ8_p & v90eed7 | !StoB_REQ8_p & v93fba3;
assign v8f37f3 = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v913a54;
assign v906ad1 = BtoS_ACK1_p & v93dfc0 | !BtoS_ACK1_p & v905381;
assign v93fa54 = StoB_REQ8_p & v87f17f | !StoB_REQ8_p & !v844f91;
assign v93fdf6 = jx3_p & v93dfc2 | !jx3_p & !v903b83;
assign v90dec8 = jx2_p & v93ea75 | !jx2_p & !v907524;
assign v90f164 = BtoR_REQ0_p & v90839e | !BtoR_REQ0_p & v93f844;
assign v908d1f = StoB_REQ1_p & v93fc8e | !StoB_REQ1_p & !v844f91;
assign v93fb58 = jx2_p & v93f701 | !jx2_p & !v85e142;
assign v93f136 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v909187;
assign v904013 = StoB_REQ9_p & v883cbe | !StoB_REQ9_p & v8b98b7;
assign v8633ac = BtoS_ACK6_p & v89f84e | !BtoS_ACK6_p & v909119;
assign v87a97c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90fc5e;
assign v93e855 = jx2_p & v9134c4 | !jx2_p & v844f91;
assign v90809e = ENQ_p & v90a61d | !ENQ_p & v8b9b9b;
assign v9063e0 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v93f6a7;
assign v93df15 = RtoB_ACK0_p & v886fce | !RtoB_ACK0_p & v86d690;
assign v89e097 = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v93fb3b;
assign v8ee1cd = jx2_p & v863a47 | !jx2_p & v90ec05;
assign v91343f = jx3_p & v93fdcc | !jx3_p & !v93fd2e;
assign v909cee = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fbff;
assign v87a21f = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9d;
assign v87de8d = RtoB_ACK0_p & v87a203 | !RtoB_ACK0_p & v9112d1;
assign v91a747 = StoB_REQ8_p & v93fdbc | !StoB_REQ8_p & !v844f91;
assign v9044c3 = StoB_REQ8_p & v93e27a | !StoB_REQ8_p & v9095b9;
assign v93eeda = jx1_p & v844f91 | !jx1_p & v90da92;
assign v87e0d8 = jx3_p & v904590 | !jx3_p & !v91a6f1;
assign v93fe20 = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v93fb31;
assign v93fe4c = BtoS_ACK0_p & v93e391 | !BtoS_ACK0_p & v93fc69;
assign v910958 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v903b70;
assign v8893bb = StoB_REQ2_p & v908346 | !StoB_REQ2_p & v93fa76;
assign v907ff8 = BtoS_ACK8_p & v89e122 | !BtoS_ACK8_p & v90f0aa;
assign v90891d = jx1_p & v93e7d1 | !jx1_p & v913072;
assign v90e25e = StoB_REQ7_p & v93f8ff | !StoB_REQ7_p & v93fa46;
assign v90ebe8 = jx2_p & v8ee1d1 | !jx2_p & v903fa3;
assign v93fe72 = RtoB_ACK1_p & v905aa1 | !RtoB_ACK1_p & v93fe61;
assign v90f8e7 = StoB_REQ1_p & v904e53 | !StoB_REQ1_p & v9077be;
assign v90f309 = StoB_REQ1_p & v906acc | !StoB_REQ1_p & v844f91;
assign v93f005 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v93fb0a;
assign v90e9e2 = BtoR_REQ0_p & v844fa9 | !BtoR_REQ0_p & v8b7122;
assign v90fa02 = EMPTY_p & v89f927 | !EMPTY_p & v903b98;
assign v90dc0d = BtoS_ACK8_p & v93f6a0 | !BtoS_ACK8_p & v863b26;
assign v93fdaf = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v93fbbe;
assign v93fb77 = BtoS_ACK8_p & v907e81 | !BtoS_ACK8_p & v861331;
assign v907916 = BtoR_REQ0_p & v93f7ef | !BtoR_REQ0_p & v93f94b;
assign v910867 = BtoS_ACK9_p & v9056a4 | !BtoS_ACK9_p & v93f77e;
assign v89e0fb = BtoS_ACK9_p & v91aa45 | !BtoS_ACK9_p & v86e625;
assign v90f5bd = BtoS_ACK7_p & v87f17f | !BtoS_ACK7_p & v844f91;
assign v909080 = BtoS_ACK6_p & v93fcc9 | !BtoS_ACK6_p & v93e650;
assign v93deab = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v906cc8;
assign v93fd7f = jx0_p & v90a4e6 | !jx0_p & v90684c;
assign v90cbf7 = StoB_REQ6_p & v912643 | !StoB_REQ6_p & v909637;
assign v910b21 = jx2_p & v88b848 | !jx2_p & v93fcf2;
assign v90ff24 = BtoS_ACK0_p & v93fc02 | !BtoS_ACK0_p & v9113de;
assign v90a9e4 = StoB_REQ6_p & v93fa55 | !StoB_REQ6_p & v93fa90;
assign v93f854 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86f729;
assign v90a3f6 = jx0_p & v93e9c7 | !jx0_p & !v93fdfa;
assign v87c537 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v9048d7;
assign v904847 = jx2_p & v905618 | !jx2_p & !v93dc08;
assign v93fdb3 = BtoS_ACK7_p & v90515d | !BtoS_ACK7_p & v89e11b;
assign v93f7bf = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v904bf3;
assign v9051e8 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v90df5b;
assign v907091 = StoB_REQ3_p & v93fd8e | !StoB_REQ3_p & v844f9f;
assign v93fcd5 = StoB_REQ1_p & v93ec07 | !StoB_REQ1_p & v93ec81;
assign v9132d4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90e083;
assign v89e0da = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v903f21;
assign v93f68f = jx2_p & v93fdc1 | !jx2_p & v85ead8;
assign v85ea96 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v90cf52;
assign v93fd25 = jx1_p & v9093ec | !jx1_p & v9096ae;
assign v908df7 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v90ed3d;
assign v93f768 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9074ce;
assign v93f73e = BtoS_ACK9_p & v93fc6d | !BtoS_ACK9_p & v93f8ec;
assign v93f7f9 = BtoS_ACK1_p & v90da97 | !BtoS_ACK1_p & v89f92f;
assign v93fdc1 = jx1_p & v910e82 | !jx1_p & !v93f7a5;
assign v903fa3 = jx1_p & v8639e7 | !jx1_p & v844f91;
assign v906d2b = StoB_REQ0_p & v909058 | !StoB_REQ0_p & v9133d9;
assign v93f15e = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v908f48;
assign v905d28 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v93fb5c;
assign v90f9fc = jx1_p & v93ecc4 | !jx1_p & v904ee9;
assign v93fd23 = jx1_p & v910710 | !jx1_p & v903fe9;
assign v90a850 = StoB_REQ7_p & v910710 | !StoB_REQ7_p & !v9057cb;
assign v87c4c5 = BtoS_ACK7_p & v93f8c1 | !BtoS_ACK7_p & !v93f6e2;
assign v910bea = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fb3e;
assign v905978 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v90a3e0;
assign v93f23c = jx2_p & v90a5c1 | !jx2_p & !v903f97;
assign v93fad5 = jx3_p & v908ad9 | !jx3_p & v90441e;
assign v904af3 = StoB_REQ2_p & v93fcf0 | !StoB_REQ2_p & v844f91;
assign v910056 = BtoS_ACK0_p & v90534f | !BtoS_ACK0_p & v93ed96;
assign v93f85a = jx0_p & v844f91 | !jx0_p & v90762a;
assign v90fe55 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v90fe87;
assign v844fc1 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v844f91;
assign v908533 = BtoS_ACK6_p & v909a26 | !BtoS_ACK6_p & v93fa87;
assign v9054c6 = jx0_p & v910bf8 | !jx0_p & v844f9d;
assign v9047eb = BtoS_ACK7_p & v93e27a | !BtoS_ACK7_p & v93f97e;
assign v90468d = BtoS_ACK8_p & v90d3ff | !BtoS_ACK8_p & v908138;
assign v906663 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v93f9bb;
assign v9113b2 = jx1_p & v903b7b | !jx1_p & v93fac6;
assign v93fb8f = StoB_REQ1_p & v905660 | !StoB_REQ1_p & v91aa76;
assign v909ecc = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v93fd3a;
assign v90d933 = BtoR_REQ0_p & v90600b | !BtoR_REQ0_p & v91090e;
assign v90a430 = BtoS_ACK6_p & v90cc30 | !BtoS_ACK6_p & v905597;
assign v905a20 = jx1_p & v93db85 | !jx1_p & !v93f88a;
assign v90d71a = StoB_REQ2_p & v93fc2a | !StoB_REQ2_p & v907b58;
assign v9071c7 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v90479a;
assign v93e810 = BtoS_ACK7_p & v8b9ee2 | !BtoS_ACK7_p & v907110;
assign v905f54 = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v87a993;
assign v93f962 = StoB_REQ6_p & v90f5b6 | !StoB_REQ6_p & v91325f;
assign v8b830b = jx1_p & v91ae94 | !jx1_p & !v93e70c;
assign v93fd04 = BtoS_ACK7_p & v9054bd | !BtoS_ACK7_p & v93fcbc;
assign v90fc9a = jx1_p & v93fb5f | !jx1_p & !v910bea;
assign v93f754 = jx0_p & v90d6e8 | !jx0_p & v844f91;
assign v910bf9 = StoB_REQ7_p & v93ee87 | !StoB_REQ7_p & v90d879;
assign v93e13e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9080a0;
assign v93fdd0 = BtoS_ACK6_p & v90630d | !BtoS_ACK6_p & v9085c8;
assign v93fd9b = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9f;
assign v93fbc2 = StoB_REQ1_p & v904b58 | !StoB_REQ1_p & v93f9d5;
assign v911db6 = jx1_p & v913332 | !jx1_p & v87f17d;
assign v908325 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v87ca92;
assign v93fd11 = StoB_REQ1_p & v93e8d3 | !StoB_REQ1_p & v844f91;
assign v90aeb7 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v909b55;
assign v91a9b6 = BtoS_ACK9_p & v90aa42 | !BtoS_ACK9_p & v90dc09;
assign v904d7e = DEQ_p & v93e731 | !DEQ_p & v91a9a2;
assign v930076 = jx1_p & v9062f7 | !jx1_p & v844f91;
assign v91a99a = jx2_p & v906315 | !jx2_p & v93f7fd;
assign v907722 = stateG7_1_p & v93fa0a | !stateG7_1_p & v93f4ac;
assign v93e882 = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v93f883;
assign v90dab9 = BtoS_ACK7_p & v910fda | !BtoS_ACK7_p & v8b4981;
assign v93fc65 = BtoS_ACK0_p & v93ea50 | !BtoS_ACK0_p & v89e0da;
assign v93fadc = StoB_REQ1_p & v905660 | !StoB_REQ1_p & v90cfc7;
assign v90441c = jx1_p & v909297 | !jx1_p & v90a181;
assign v93fe49 = StoB_REQ8_p & v87f17f | !StoB_REQ8_p & !v90a604;
assign v93e5b8 = jx2_p & v90a5ee | !jx2_p & v844f91;
assign v89f844 = BtoS_ACK1_p & v93dfc0 | !BtoS_ACK1_p & v905df9;
assign v93fb13 = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v910f3a;
assign v90567a = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fdb3;
assign v90fc42 = stateG7_1_p & v8b9996 | !stateG7_1_p & v93f6c7;
assign v93f07c = BtoS_ACK9_p & v91104c | !BtoS_ACK9_p & v90f83e;
assign v93fab9 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fc49;
assign v912fad = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v844fa3;
assign v906913 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v906cd3;
assign v93e14a = StoB_REQ3_p & v911311 | !StoB_REQ3_p & v907aa0;
assign v90f6b5 = BtoR_REQ0_p & v913a94 | !BtoR_REQ0_p & v907d9d;
assign v9105f4 = jx3_p & v93fdf1 | !jx3_p & !v906209;
assign v9134cc = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v930076;
assign v93f897 = StoB_REQ9_p & v90712d | !StoB_REQ9_p & v844f91;
assign v910f78 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v87a21f;
assign v911185 = jx2_p & v90dc9c | !jx2_p & !v90ec05;
assign v93fa8f = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v85e7ba;
assign v913a60 = jx0_p & v93f714 | !jx0_p & v93f685;
assign v88e67b = StoB_REQ7_p & v93f7e3 | !StoB_REQ7_p & v844f91;
assign v8b9f37 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v87bae8;
assign v910461 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v93f9e7;
assign v908250 = StoB_REQ8_p & v93ed2a | !StoB_REQ8_p & v90653d;
assign v904f4d = jx1_p & v87c52b | !jx1_p & !v90fa8a;
assign v93fc48 = ENQ_p & v93eda4 | !ENQ_p & v8d37d6;
assign v90d7e8 = BtoS_ACK9_p & v9114a0 | !BtoS_ACK9_p & v93fe45;
assign v93f7c9 = jx1_p & v93e0b5 | !jx1_p & v85ead8;
assign v93f990 = jx0_p & v90d8d8 | !jx0_p & v904ecc;
assign v93e875 = BtoS_ACK8_p & v93ed2a | !BtoS_ACK8_p & v903c2a;
assign v910cf1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fdfe;
assign v93e391 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90a59e;
assign v93f8b8 = DEQ_p & v93fad3 | !DEQ_p & v93e301;
assign v90cf68 = jx3_p & v93e105 | !jx3_p & !v89e05b;
assign v88b848 = jx1_p & v93f9ad | !jx1_p & v90481b;
assign v93ee4b = StoB_REQ7_p & v912679 | !StoB_REQ7_p & v859635;
assign v90986f = jx1_p & v93fd51 | !jx1_p & !v87b2ea;
assign v91879a = BtoS_ACK6_p & v93e89f | !BtoS_ACK6_p & !v8a8fed;
assign v93f97d = StoB_REQ8_p & v93eabc | !StoB_REQ8_p & v90d546;
assign v90d1ca = StoB_REQ2_p & v90fe49 | !StoB_REQ2_p & v908a34;
assign v909458 = stateG7_1_p & v90d64c | !stateG7_1_p & v93fd67;
assign v93fe17 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93fb2b;
assign v91132f = jx0_p & v90ed41 | !jx0_p & v844f91;
assign v93f749 = BtoS_ACK9_p & v910c51 | !BtoS_ACK9_p & v89b1a2;
assign v93fd6c = BtoS_ACK9_p & v93e05f | !BtoS_ACK9_p & v903db4;
assign v93e5da = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & !v910e69;
assign v90a53b = jx1_p & v93eb20 | !jx1_p & v93fd2f;
assign v863450 = StoB_REQ9_p & v93fd76 | !StoB_REQ9_p & v93f646;
assign v91aa04 = stateG12_p & v844f91 | !stateG12_p & !v87f17f;
assign v93e2a0 = RtoB_ACK0_p & v93fad3 | !RtoB_ACK0_p & v91359a;
assign v90decf = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v89f840;
assign v90ad03 = ENQ_p & v912477 | !ENQ_p & v8baf9a;
assign v90cb3d = jx1_p & v912fa9 | !jx1_p & v93fdd0;
assign v93fc5f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v907897;
assign v8b9e4f = jx2_p & v9042b8 | !jx2_p & !v90a90b;
assign v93f9bf = DEQ_p & v88bb45 | !DEQ_p & v87d990;
assign v907a1b = jx3_p & v9109e6 | !jx3_p & !v90d731;
assign v93e371 = BtoS_ACK6_p & v8b49ad | !BtoS_ACK6_p & v90d21a;
assign v906769 = RtoB_ACK0_p & v90f629 | !RtoB_ACK0_p & v93fe5d;
assign v93f776 = StoB_REQ8_p & v87f17f | !StoB_REQ8_p & v89e10d;
assign v9135d1 = BtoS_ACK8_p & v907e81 | !BtoS_ACK8_p & v904838;
assign v9097db = BtoS_ACK9_p & v93e9b9 | !BtoS_ACK9_p & v9052f2;
assign v9051ba = jx3_p & v93e105 | !jx3_p & !v93fb26;
assign v8b9ef8 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v93f092;
assign v93fe46 = StoB_REQ2_p & v93fe36 | !StoB_REQ2_p & !v93fd3a;
assign v85eaab = StoB_REQ6_p & v90f5b6 | !StoB_REQ6_p & v9051c3;
assign v93f979 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fd76;
assign v9117de = StoB_REQ9_p & v8d37d4 | !StoB_REQ9_p & v90a36a;
assign v90e88f = BtoS_ACK8_p & v9101ae | !BtoS_ACK8_p & !v93fa0d;
assign v93f39f = jx1_p & v93fbe5 | !jx1_p & v906491;
assign v9082ba = BtoS_ACK6_p & v8a8b0a | !BtoS_ACK6_p & v87f17d;
assign v93e188 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v93fe71;
assign v93f65b = BtoR_REQ0_p & v93fba0 | !BtoR_REQ0_p & v93fcc6;
assign v93e007 = jx2_p & v863476 | !jx2_p & !v93f7e9;
assign v93fbba = jx0_p & v909e2c | !jx0_p & v844f9d;
assign v90cbfd = StoB_REQ8_p & v93dbe9 | !StoB_REQ8_p & v90a4da;
assign v906c35 = jx0_p & v844f91 | !jx0_p & v93fb3e;
assign v93e89f = jx0_p & v844f97 | !jx0_p & !v844f91;
assign v90a4a1 = StoB_REQ9_p & v86dde6 | !StoB_REQ9_p & v93fa2a;
assign v8f381e = BtoS_ACK8_p & v93fb93 | !BtoS_ACK8_p & v90931a;
assign v93e77d = BtoS_ACK6_p & v93e126 | !BtoS_ACK6_p & v91a6d5;
assign v90f2ff = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v93f685;
assign v89f7e2 = StoB_REQ3_p & v90f547 | !StoB_REQ3_p & v844f9f;
assign v9102bf = BtoS_ACK0_p & v93e77b | !BtoS_ACK0_p & v905eaa;
assign v906c10 = StoB_REQ3_p & v908eea | !StoB_REQ3_p & !v844f91;
assign v93fbb4 = BtoS_ACK9_p & v89f7dd | !BtoS_ACK9_p & v9058c2;
assign v90799d = BtoS_ACK8_p & v93f6a0 | !BtoS_ACK8_p & v93fb74;
assign v9112d1 = FULL_p & v844f91 | !FULL_p & v907a32;
assign v93f928 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v909078;
assign v910101 = StoB_REQ8_p & v90e2d7 | !StoB_REQ8_p & v90844d;
assign v8f3865 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90da92;
assign v9049fd = jx1_p & v93e065 | !jx1_p & v93fd22;
assign v93f762 = StoB_REQ0_p & v844f97 | !StoB_REQ0_p & v90855a;
assign v93f51c = jx0_p & v844f91 | !jx0_p & v90539f;
assign v904c52 = StoB_REQ8_p & v93fc15 | !StoB_REQ8_p & v844f91;
assign v90e7d7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v90a8c3;
assign v908ed2 = ENQ_p & v93f92a | !ENQ_p & v90a49d;
assign v904521 = BtoS_ACK0_p & v904b63 | !BtoS_ACK0_p & v89f80d;
assign v90a4bb = DEQ_p & v9051ba | !DEQ_p & v93e203;
assign v93f9b8 = DEQ_p & v8f22ca | !DEQ_p & v93f919;
assign v907517 = BtoS_ACK8_p & v93f6fb | !BtoS_ACK8_p & v93fd38;
assign v8b9d4b = BtoS_ACK9_p & v90cbfd | !BtoS_ACK9_p & v90e925;
assign v9071ed = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v90f947;
assign v907da6 = StoB_REQ8_p & v90529c | !StoB_REQ8_p & v85e94c;
assign v908e7f = DEQ_p & v93fd1b | !DEQ_p & v844f91;
assign v85f240 = jx1_p & v90893a | !jx1_p & !v844f91;
assign v93f6ea = jx1_p & v93f910 | !jx1_p & v93e89f;
assign v93f10b = EMPTY_p & v89f927 | !EMPTY_p & v9086f1;
assign v90e1d0 = BtoS_ACK6_p & v906d58 | !BtoS_ACK6_p & v90479c;
assign v9041a7 = RtoB_ACK0_p & v90744a | !RtoB_ACK0_p & v87e0d8;
assign v93f9f7 = EMPTY_p & v905ac3 | !EMPTY_p & v93e69c;
assign v91a733 = ENQ_p & v9101d0 | !ENQ_p & v844f91;
assign v90ad75 = jx0_p & v93f9c6 | !jx0_p & v844f95;
assign v9088de = BtoS_ACK1_p & v90fc92 | !BtoS_ACK1_p & v9134c0;
assign v90f8f5 = BtoS_ACK1_p & v93dffe | !BtoS_ACK1_p & v93fd50;
assign v9044b8 = jx0_p & v844f91 | !jx0_p & !v93fd21;
assign v9079f4 = StoB_REQ8_p & v904ab4 | !StoB_REQ8_p & v9047eb;
assign v909d1c = DEQ_p & v9087b7 | !DEQ_p & v907a32;
assign v90932c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f362;
assign v93fc94 = StoB_REQ7_p & v93fc68 | !StoB_REQ7_p & !v9093ec;
assign v8d37d6 = jx3_p & v844f91 | !jx3_p & !v93f6cf;
assign v90f78a = StoB_REQ7_p & v93ee87 | !StoB_REQ7_p & v908533;
assign v91a7a5 = BtoR_REQ1_p & v878dab | !BtoR_REQ1_p & v9050ad;
assign v93f5e9 = jx0_p & v93fd6f | !jx0_p & !v85eaf1;
assign v9079ac = BtoS_ACK9_p & v91104c | !BtoS_ACK9_p & v89e0d7;
assign v906c48 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v9067c1;
assign v93fc69 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9058f4;
assign v93f6b7 = BtoS_ACK8_p & v907adb | !BtoS_ACK8_p & v93fc85;
assign v9099a1 = BtoS_ACK9_p & v93f73d | !BtoS_ACK9_p & v910ea0;
assign v90479a = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v90fe49;
assign v93e7c2 = BtoS_ACK0_p & v86e433 | !BtoS_ACK0_p & v8f22e0;
assign v93fa47 = BtoR_REQ0_p & v93fa8d | !BtoR_REQ0_p & v912173;
assign v906a80 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fde5;
assign v93fb37 = StoB_REQ0_p & v9071c7 | !StoB_REQ0_p & v8ee181;
assign v8b49cc = StoB_REQ9_p & v93f098 | !StoB_REQ9_p & !v93f5ff;
assign v90851b = BtoS_ACK9_p & v93f66f | !BtoS_ACK9_p & v904e00;
assign v93f6d8 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v93fd4e;
assign v90e40b = jx1_p & v9062f7 | !jx1_p & v93f2d9;
assign v93fd8c = jx2_p & v9135db | !jx2_p & !v93fb9d;
assign v90fc26 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v905d63;
assign v905df9 = BtoS_ACK2_p & v9123a2 | !BtoS_ACK2_p & v8f2234;
assign v90ef1a = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93f856;
assign v93fb3e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f5d1;
assign v93fd8d = jx1_p & v93ecc4 | !jx1_p & v9056d9;
assign v90d78b = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & !v909366;
assign v85f2b9 = StoB_REQ8_p & v90eed7 | !StoB_REQ8_p & v93fd33;
assign v90ad6f = ENQ_p & v93eed6 | !ENQ_p & v844f91;
assign v904ec6 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f792;
assign v908e4b = stateG12_p & v8b9b88 | !stateG12_p & v93fac4;
assign v909dc3 = ENQ_p & v93e5f1 | !ENQ_p & v905077;
assign v93f6c7 = RtoB_ACK0_p & v907b60 | !RtoB_ACK0_p & v93f204;
assign v909722 = DEQ_p & v93fd1b | !DEQ_p & v9052ba;
assign v93f7ce = StoB_REQ2_p & v93fcf0 | !StoB_REQ2_p & v92ffc9;
assign v93fb0b = jx0_p & v9107c7 | !jx0_p & v910f4d;
assign v908096 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v908df7;
assign v90f4dd = BtoS_ACK9_p & v87f17f | !BtoS_ACK9_p & !v907200;
assign v913068 = BtoS_ACK8_p & v90451f | !BtoS_ACK8_p & v93fcdc;
assign v93f941 = jx0_p & v93f70c | !jx0_p & v93f709;
assign v906195 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v90817e;
assign v909eab = jx0_p & v91104b | !jx0_p & v905824;
assign v90f5ff = BtoS_ACK6_p & v9050a5 | !BtoS_ACK6_p & v907edc;
assign v90f3e4 = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v907b65;
assign v90a96f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v93f490;
assign v905556 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910be8;
assign v90a2fc = jx1_p & v91ae94 | !jx1_p & v9124b8;
assign v93f910 = jx0_p & v844f9b | !jx0_p & !v844f91;
assign v904434 = jx1_p & v9126b6 | !jx1_p & v8f3849;
assign v93fd44 = RtoB_ACK0_p & v90e333 | !RtoB_ACK0_p & v93e301;
assign v93f830 = ENQ_p & v907c69 | !ENQ_p & v844f91;
assign v904931 = BtoS_ACK1_p & v93f85e | !BtoS_ACK1_p & v90a47f;
assign v9090dd = StoB_REQ6_p & v93f9c6 | !StoB_REQ6_p & v90cc30;
assign v90a30e = BtoS_ACK0_p & v8bb868 | !BtoS_ACK0_p & v93df55;
assign v909157 = BtoS_ACK0_p & v93fccb | !BtoS_ACK0_p & v90ea1f;
assign v90dcc6 = jx2_p & v93f678 | !jx2_p & v90eaad;
assign v903cd1 = EMPTY_p & v9082be | !EMPTY_p & v90fb00;
assign v912ef3 = BtoS_ACK6_p & v90db9f | !BtoS_ACK6_p & v844f91;
assign v93fb7d = StoB_REQ8_p & v903c2a | !StoB_REQ8_p & v93f813;
assign v93fc9d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fbb7;
assign v904abd = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v904da6;
assign v93f70b = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v907102;
assign v90914c = StoB_REQ1_p & v93e9cc | !StoB_REQ1_p & v93f7a2;
assign v904182 = StoB_REQ5_p & v844fbb | !StoB_REQ5_p & v844f91;
assign v93e8de = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v93e295;
assign v90f9f3 = BtoS_ACK8_p & v907e81 | !BtoS_ACK8_p & v907469;
assign v93fade = jx0_p & v93e9c7 | !jx0_p & !v906a79;
assign v93f92f = jx0_p & v903c09 | !jx0_p & !v87bf0e;
assign v90a7f2 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v906416;
assign v912f40 = StoB_REQ0_p & v93f7f5 | !StoB_REQ0_p & v844f91;
assign v93f75f = ENQ_p & v90adc4 | !ENQ_p & v89f95b;
assign v93ef38 = jx3_p & v93fbcc | !jx3_p & v93ea9e;
assign v8b49ad = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fe07;
assign v90a557 = jx2_p & v93e829 | !jx2_p & v93fb20;
assign v93e115 = jx2_p & v9080c5 | !jx2_p & v844f91;
assign v93fd49 = DEQ_p & v9041a7 | !DEQ_p & v87e0d8;
assign v93dc2c = BtoS_ACK8_p & v90fe87 | !BtoS_ACK8_p & v90edb9;
assign v907add = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v93f32b;
assign v911311 = BtoS_ACK4_p & v844f9f | !BtoS_ACK4_p & !v904182;
assign v88aff7 = StoB_REQ9_p & v913362 | !StoB_REQ9_p & v91267b;
assign v911973 = jx1_p & v93e7d1 | !jx1_p & !v9091fe;
assign v90a798 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9054c9;
assign v903bfc = BtoS_ACK9_p & v90aa3b | !BtoS_ACK9_p & v93f7ca;
assign v93faa7 = jx1_p & v90d543 | !jx1_p & v911417;
assign v8b99c6 = BtoR_REQ1_p & v93fb1c | !BtoR_REQ1_p & v909dc9;
assign v93f7d6 = ENQ_p & v863add | !ENQ_p & !v905a5b;
assign v90f2f8 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v90a18c;
assign v93fbb0 = jx1_p & v9043ec | !jx1_p & v844f91;
assign v93fd50 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v906c71;
assign v93fcdd = BtoS_ACK9_p & v906a80 | !BtoS_ACK9_p & v93f698;
assign v93fd1e = BtoS_ACK7_p & v90cc57 | !BtoS_ACK7_p & v91a99a;
assign v93eade = StoB_REQ9_p & v8d37d4 | !StoB_REQ9_p & v910cbf;
assign v90acc4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9063e0;
assign v93e919 = jx1_p & v908aa8 | !jx1_p & !v91192b;
assign v90e611 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v908127;
assign v907580 = jx1_p & v913435 | !jx1_p & v844f91;
assign v90ad48 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v909d2b;
assign v903fb2 = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v90946a;
assign v906256 = BtoS_ACK6_p & v912679 | !BtoS_ACK6_p & !v90d2b7;
assign v905136 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90534f;
assign v903d68 = EMPTY_p & v9051ae | !EMPTY_p & v910fcd;
assign v90f787 = BtoS_ACK8_p & v90ba1a | !BtoS_ACK8_p & v90a7f2;
assign v91dc98 = jx1_p & v89e11b | !jx1_p & v93faa4;
assign v90a27c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90f8f5;
assign v93f906 = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & !v93f6a7;
assign v93fd74 = DEQ_p & v93fc76 | !DEQ_p & v90dd67;
assign v9091c6 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v911946;
assign v905cd2 = BtoS_ACK2_p & v91305b | !BtoS_ACK2_p & v903cd2;
assign v909107 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v93fd87;
assign v8633ef = jx0_p & v93e337 | !jx0_p & !v8b9efa;
assign v9133dc = BtoS_ACK8_p & v904a80 | !BtoS_ACK8_p & v904878;
assign v93f708 = BtoS_ACK9_p & v9044c3 | !BtoS_ACK9_p & v93f97c;
assign v910e32 = jx1_p & v93f8d0 | !jx1_p & v906dd6;
assign v93f33e = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v8a8fa0;
assign v93fa81 = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & !v909e7f;
assign v90fbfd = jx2_p & v90d634 | !jx2_p & v93fb39;
assign v93f82e = StoB_REQ7_p & v909705 | !StoB_REQ7_p & v90a2b8;
assign v903e08 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v93fbd3;
assign v93f73a = EMPTY_p & v844f91 | !EMPTY_p & v909d1c;
assign v904671 = DEQ_p & v93f6fa | !DEQ_p & v912f3d;
assign v93f825 = StoB_REQ8_p & v93f06e | !StoB_REQ8_p & !v844f91;
assign v93f0a6 = BtoS_ACK9_p & v93fcbf | !BtoS_ACK9_p & v90fc26;
assign v93eaa6 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v9103e4;
assign v9111d3 = EMPTY_p & v93f77b | !EMPTY_p & v93f728;
assign v9056c5 = StoB_REQ2_p & v93fd09 | !StoB_REQ2_p & v912672;
assign v89fdcf = StoB_REQ0_p & v93db4a | !StoB_REQ0_p & v93ebb5;
assign v93fb95 = StoB_REQ6_p & v8d3799 | !StoB_REQ6_p & v903c46;
assign v9101ae = jx2_p & v905a20 | !jx2_p & v910f2e;
assign v906416 = BtoS_ACK7_p & v904b45 | !BtoS_ACK7_p & v89e11b;
assign v93fc53 = jx3_p & v844f91 | !jx3_p & v905460;
assign v912ec8 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v93fbd2;
assign v911509 = jx0_p & v903e85 | !jx0_p & v9132b0;
assign v9130af = jx0_p & v85dee0 | !jx0_p & v93eece;
assign v90728a = BtoS_ACK7_p & v90529c | !BtoS_ACK7_p & v93fce9;
assign v884261 = BtoS_ACK6_p & v86344b | !BtoS_ACK6_p & v9044b4;
assign v93f898 = StoB_REQ8_p & v904b00 | !StoB_REQ8_p & v90a2aa;
assign v90866d = BtoS_ACK9_p & v911909 | !BtoS_ACK9_p & v90e926;
assign v904c72 = StoB_REQ8_p & v90638b | !StoB_REQ8_p & v90faf1;
assign v90ec84 = jx1_p & v8b9c1e | !jx1_p & !v910bea;
assign v863ac4 = ENQ_p & v93e704 | !ENQ_p & v905312;
assign v905847 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93fb86;
assign v8cec7e = StoB_REQ8_p & v93e27a | !StoB_REQ8_p & v9134e2;
assign v90962e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v911023;
assign v905da0 = jx3_p & v93f110 | !jx3_p & v89f9dc;
assign v93fdd2 = jx2_p & v844f91 | !jx2_p & !v907e86;
assign v93fa49 = StoB_REQ2_p & v8b98bd | !StoB_REQ2_p & v89f8e5;
assign v90d057 = ENQ_p & v87e7f5 | !ENQ_p & v9117e2;
assign v906ec1 = jx2_p & v93fd75 | !jx2_p & !v844f91;
assign v93f96e = jx1_p & v911edb | !jx1_p & v903fb2;
assign v93fd0c = jx0_p & v93dade | !jx0_p & !v9061b0;
assign v90cbea = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v904e13;
assign v9088a3 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v9101b8;
assign v909430 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v905186;
assign v93e301 = ENQ_p & v911a33 | !ENQ_p & v844f91;
assign v9049e4 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93f77a;
assign v93fafc = jx3_p & v844f91 | !jx3_p & v90add9;
assign v93fbf4 = BtoS_ACK8_p & v93fb92 | !BtoS_ACK8_p & v9056a0;
assign v93f91f = jx2_p & v906a5c | !jx2_p & v863afc;
assign v908a3d = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v93fbe8;
assign v906414 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f8ee;
assign v93f6f4 = RtoB_ACK0_p & v93f73c | !RtoB_ACK0_p & v89f796;
assign v904d51 = ENQ_p & v90a61d | !ENQ_p & v90cbf3;
assign v9049a9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93e86c;
assign v90fe49 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9b;
assign v93f7a9 = jx0_p & v844f91 | !jx0_p & v93f895;
assign v903c46 = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v9052de;
assign v8b9efa = StoB_REQ6_p & v93edc8 | !StoB_REQ6_p & v93fe00;
assign v90d9a0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90a300;
assign v93fe5a = BtoS_ACK8_p & v904847 | !BtoS_ACK8_p & !v90ed6e;
assign v91aa3f = jx1_p & v93f89e | !jx1_p & !v93f6d8;
assign v93f878 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844fb9;
assign v907840 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f280;
assign v93faac = RtoB_ACK0_p & v907a4d | !RtoB_ACK0_p & v871483;
assign v93e652 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v906cd3;
assign v908357 = BtoS_ACK0_p & v93fc02 | !BtoS_ACK0_p & v9045c0;
assign v910d4a = BtoS_ACK9_p & v93f898 | !BtoS_ACK9_p & v873bc3;
assign v93fe1b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v9080f5;
assign v9052f2 = StoB_REQ9_p & v9046f9 | !StoB_REQ9_p & v87c558;
assign v909ab9 = BtoS_ACK6_p & v90d718 | !BtoS_ACK6_p & v89f852;
assign v908e01 = StoB_REQ6_p & v93fdde | !StoB_REQ6_p & v93f762;
assign v87b4fc = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v911311;
assign v93e337 = StoB_REQ6_p & v93faeb | !StoB_REQ6_p & v906c8c;
assign v93fcc4 = StoB_REQ8_p & v908237 | !StoB_REQ8_p & v844f91;
assign v904088 = BtoS_ACK1_p & v913348 | !BtoS_ACK1_p & v93e7d4;
assign v90f7a1 = StoB_REQ7_p & v93fbf0 | !StoB_REQ7_p & v8b9dbd;
assign v9076a8 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v91058e;
assign v90e5b4 = jx3_p & v93fdda | !jx3_p & v905246;
assign v911b47 = StoB_REQ8_p & v93fb71 | !StoB_REQ8_p & v93e6f6;
assign v908176 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93dc2c;
assign v93fa2e = BtoS_ACK9_p & v8b98d4 | !BtoS_ACK9_p & v90f994;
assign v93ed58 = BtoS_ACK9_p & v93f7c3 | !BtoS_ACK9_p & v93fd68;
assign v9131c9 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93f1c8;
assign v911005 = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v93fc4d;
assign v93fa87 = jx0_p & v90d879 | !jx0_p & v90762a;
assign v88946f = StoB_REQ0_p & v93fc34 | !StoB_REQ0_p & v91071b;
assign v93f701 = jx1_p & v8f22d1 | !jx1_p & !v88e67b;
assign v912124 = BtoS_ACK0_p & v913619 | !BtoS_ACK0_p & v93f88f;
assign v8a8f74 = BtoS_ACK6_p & v8b49ad | !BtoS_ACK6_p & v8a927b;
assign v918886 = EMPTY_p & v90fc42 | !EMPTY_p & !v904a3b;
assign v90f5b6 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v909058;
assign v9050d2 = StoB_REQ3_p & v911311 | !StoB_REQ3_p & v844f91;
assign v8b9c5f = StoB_REQ6_p & v85dee0 | !StoB_REQ6_p & v90ef1b;
assign v90db9e = BtoS_ACK7_p & v93fdd2 | !BtoS_ACK7_p & v93fd0f;
assign v93e2b8 = ENQ_p & v908325 | !ENQ_p & v904091;
assign v912fed = jx0_p & v913435 | !jx0_p & v844f91;
assign v906f62 = RtoB_ACK0_p & v93f284 | !RtoB_ACK0_p & v93f899;
assign v93f9a7 = BtoS_ACK8_p & v89e07c | !BtoS_ACK8_p & v93f6a6;
assign v91aa44 = StoB_REQ6_p & v909107 | !StoB_REQ6_p & v8b9c50;
assign v93fd33 = BtoS_ACK7_p & v90a07e | !BtoS_ACK7_p & v93eb9e;
assign v90636b = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v909174;
assign v87c9f1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v905405;
assign v906c6f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v909434;
assign v93f0b0 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v93df06;
assign v8a9267 = BtoR_REQ1_p & v844fab | !BtoR_REQ1_p & v904f76;
assign v93fc2d = RtoB_ACK0_p & v93fc48 | !RtoB_ACK0_p & v910fcd;
assign v906cd3 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v90e978;
assign v90446a = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v904b77;
assign v93e150 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v93f770;
assign v90caeb = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v9056c5;
assign v93fddd = StoB_REQ6_p & v93db03 | !StoB_REQ6_p & v844f91;
assign v90d5c3 = DEQ_p & v91359a | !DEQ_p & v93faf4;
assign v89f8fd = jx1_p & v93f768 | !jx1_p & !v93f7de;
assign v93fb2b = StoB_REQ0_p & v905da3 | !StoB_REQ0_p & v844f91;
assign v863418 = ENQ_p & v93f59b | !ENQ_p & v90fe7e;
assign v93fce9 = jx2_p & v8ee1d1 | !jx2_p & v93fd35;
assign v93fc0e = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v90db49;
assign v910d2f = DEQ_p & v93f0b8 | !DEQ_p & v90f629;
assign v904ae0 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v90e945;
assign v93fb9d = jx1_p & v90985e | !jx1_p & !v882135;
assign v93df10 = jx2_p & v910cf2 | !jx2_p & v910ca7;
assign v93f9f4 = jx1_p & v93fca0 | !jx1_p & v90a102;
assign v90a3da = jx1_p & v88d5cd | !jx1_p & v90fb5d;
assign v90fe87 = jx1_p & v8b9dff | !jx1_p & v844f91;
assign v9133ec = FULL_p & v89e0d5 | !FULL_p & v90dd67;
assign v86e277 = ENQ_p & v8b98f1 | !ENQ_p & v904a70;
assign v93f2a0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v91a9cd;
assign v90fe5c = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v93fbc2;
assign v9075fd = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v91035c;
assign v9115a9 = BtoS_ACK7_p & v90f575 | !BtoS_ACK7_p & v93faf9;
assign v909e2c = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v908fba;
assign v93fd86 = BtoS_ACK7_p & v93dbe9 | !BtoS_ACK7_p & v90edf6;
assign v90db49 = StoB_REQ0_p & v85eabe | !StoB_REQ0_p & v93fdd4;
assign v9098bb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fb45;
assign v911a00 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v93fcb4;
assign v93f307 = BtoS_ACK6_p & v90860a | !BtoS_ACK6_p & v9044c6;
assign v9050ae = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v89f8ef;
assign v90a2b5 = StoB_REQ9_p & v903c0d | !StoB_REQ9_p & v90a63a;
assign v9050a5 = jx0_p & v904575 | !jx0_p & !v844f99;
assign v904775 = jx0_p & v93fdb0 | !jx0_p & v904f5c;
assign v89f9dc = BtoS_ACK9_p & v9073c5 | !BtoS_ACK9_p & v906b22;
assign v93fc6c = ENQ_p & v9083cf | !ENQ_p & v93fd73;
assign v8b99a1 = DEQ_p & v844f91 | !DEQ_p & !v904f93;
assign v8b98bd = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v905702;
assign v930037 = jx0_p & v93005b | !jx0_p & !v844f91;
assign v90e893 = jx2_p & v87f17f | !jx2_p & v908ed6;
assign v907e3f = StoB_REQ8_p & v93fd76 | !StoB_REQ8_p & v844f91;
assign v904345 = BtoS_ACK7_p & v906ec1 | !BtoS_ACK7_p & v904c80;
assign v906320 = BtoS_ACK6_p & v903e94 | !BtoS_ACK6_p & v903cc5;
assign v90d7ce = jx1_p & v93fe6e | !jx1_p & v93fdf8;
assign v90cfc7 = BtoS_ACK2_p & v906cc8 | !BtoS_ACK2_p & v90466e;
assign v90936b = BtoS_ACK6_p & v90db9f | !BtoS_ACK6_p & v90ada1;
assign v93f7e5 = StoB_REQ7_p & v903f58 | !StoB_REQ7_p & v9095df;
assign v90d86f = jx3_p & v9064e9 | !jx3_p & v844f91;
assign v93fa29 = BtoS_ACK9_p & v93fc6d | !BtoS_ACK9_p & v8b49cc;
assign v909927 = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v87a1f9;
assign v93e7ac = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v909691;
assign v93f6ff = FULL_p & v93fb21 | !FULL_p & v907bd4;
assign v89f98c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a620;
assign v93fa70 = jx1_p & v90e6f1 | !jx1_p & !v844f91;
assign v93f7ef = EMPTY_p & v93f695 | !EMPTY_p & v907321;
assign v93fdbd = jx1_p & v90804e | !jx1_p & v93f864;
assign v8b9f15 = BtoS_ACK9_p & v9074fa | !BtoS_ACK9_p & v863ad6;
assign v91047b = DEQ_p & v905ba4 | !DEQ_p & v863a64;
assign v912fc9 = StoB_REQ9_p & v906b64 | !StoB_REQ9_p & v844f91;
assign v93eb22 = jx1_p & v93f92c | !jx1_p & v844f91;
assign v904e93 = RtoB_ACK0_p & v90ff49 | !RtoB_ACK0_p & v8b9e1d;
assign v9109e6 = BtoS_ACK9_p & v90d78b | !BtoS_ACK9_p & !v863450;
assign v90d3ff = jx2_p & v90fae7 | !jx2_p & v908ed6;
assign v9096f0 = jx1_p & v93f119 | !jx1_p & v93fd48;
assign v9096ae = jx0_p & v93fa17 | !jx0_p & !v89c5e3;
assign v86fe09 = StoB_REQ7_p & v93f8a6 | !StoB_REQ7_p & v91134b;
assign v93ed2a = jx2_p & v90a175 | !jx2_p & v9130c9;
assign v906df6 = StoB_REQ6_p & v93eece | !StoB_REQ6_p & v93f6d5;
assign v8f2234 = StoB_REQ2_p & v908127 | !StoB_REQ2_p & v9080f5;
assign v90ad39 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8d37f5;
assign v90dc0a = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v93fb9a;
assign v89e121 = BtoS_ACK6_p & v93f6eb | !BtoS_ACK6_p & v93f7a9;
assign v93f92c = BtoS_ACK6_p & v9050a5 | !BtoS_ACK6_p & v93fade;
assign v93e0c9 = BtoS_ACK9_p & v905d97 | !BtoS_ACK9_p & v906f72;
assign v93f6dc = StoB_REQ6_p & v909107 | !StoB_REQ6_p & v910e6e;
assign v908237 = jx2_p & v93e310 | !jx2_p & v93f2a4;
assign v912fb2 = EMPTY_p & v85eaa2 | !EMPTY_p & v93f781;
assign v8b9b9b = jx3_p & v908429 | !jx3_p & v93fa03;
assign v93fa5b = jx1_p & v90f7a1 | !jx1_p & v910c50;
assign v907468 = BtoS_ACK2_p & v9123a2 | !BtoS_ACK2_p & v908553;
assign v91aa52 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93f203;
assign v906665 = BtoS_ACK6_p & v8b9b9f | !BtoS_ACK6_p & v93fbf9;
assign v93f77b = stateG7_1_p & v8633bd | !stateG7_1_p & v906f62;
assign v911941 = jx1_p & v93fa53 | !jx1_p & !v93fada;
assign v89f9d7 = BtoS_ACK0_p & v93fc02 | !BtoS_ACK0_p & v90a27c;
assign v93fbd6 = BtoS_ACK0_p & v93fdfe | !BtoS_ACK0_p & v87a97c;
assign v93fa4e = jx1_p & v93f223 | !jx1_p & !v911ed7;
assign v93f7e1 = ENQ_p & v908325 | !ENQ_p & v906a84;
assign v908867 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v91267e;
assign v87a1f2 = BtoS_ACK1_p & v93dffe | !BtoS_ACK1_p & v910820;
assign v90517f = BtoR_REQ0_p & v93f9da | !BtoR_REQ0_p & v903b4e;
assign v93fdba = BtoS_ACK2_p & v9123a2 | !BtoS_ACK2_p & v9090c9;
assign v9068b6 = BtoS_ACK0_p & v93f85e | !BtoS_ACK0_p & v93fe6a;
assign v93fad2 = BtoS_ACK8_p & v87f17f | !BtoS_ACK8_p & !v93fa54;
assign v9073c3 = StoB_REQ0_p & v85eabe | !StoB_REQ0_p & v93fb45;
assign v93fd2b = StoB_REQ4_p & v844f9f | !StoB_REQ4_p & v844f91;
assign v907048 = BtoS_ACK1_p & v913348 | !BtoS_ACK1_p & v8f382c;
assign v911edd = BtoS_ACK6_p & v91aa51 | !BtoS_ACK6_p & v93f9b0;
assign v93e852 = EMPTY_p & v93e301 | !EMPTY_p & v90a074;
assign v908ff3 = BtoS_ACK9_p & v90529c | !BtoS_ACK9_p & v93f764;
assign v93f8f8 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v89f840;
assign v90a233 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v90611f;
assign v904cb5 = jx2_p & v93f6a4 | !jx2_p & !v844f91;
assign v93f8a0 = BtoS_ACK0_p & v90f624 | !BtoS_ACK0_p & v8f22a5;
assign v93fda2 = BtoS_ACK7_p & v93f23c | !BtoS_ACK7_p & v9101be;
assign v93f855 = jx1_p & v844f91 | !jx1_p & v90e841;
assign v910b22 = EMPTY_p & v904c4f | !EMPTY_p & v904fd6;
assign v89e042 = jx1_p & v863477 | !jx1_p & !v9090dd;
assign v89f79e = StoB_REQ0_p & v91218a | !StoB_REQ0_p & v844f91;
assign v93f767 = BtoR_REQ0_p & v90fa02 | !BtoR_REQ0_p & v909dd5;
assign v93fcbe = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f97;
assign v93fd9c = BtoS_ACK8_p & v9099e1 | !BtoS_ACK8_p & v93f9ac;
assign v93f8de = RtoB_ACK0_p & v863418 | !RtoB_ACK0_p & v88a51e;
assign v9096f1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a563;
assign v93f3b9 = BtoS_ACK8_p & v93e27a | !BtoS_ACK8_p & v93fb71;
assign v90a3f5 = jx2_p & v87bf17 | !jx2_p & v906e08;
assign v93f87f = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v908836;
assign v91305d = BtoS_ACK1_p & v9046a6 | !BtoS_ACK1_p & v904ae0;
assign v8b70a3 = BtoS_ACK8_p & v907eaa | !BtoS_ACK8_p & v89f9cd;
assign v904008 = jx1_p & v869aeb | !jx1_p & !v87a261;
assign v90db9f = jx0_p & v910cf1 | !jx0_p & v90e6e5;
assign v905636 = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v93e0a0;
assign v88e6c4 = jx0_p & v88de63 | !jx0_p & v844f91;
assign v93f21c = StoB_REQ7_p & v93fcf3 | !StoB_REQ7_p & v93fe3d;
assign v93fdae = jx2_p & v913169 | !jx2_p & v908ed6;
assign v910d41 = jx2_p & v9084f4 | !jx2_p & v906dd6;
assign v9090d6 = BtoS_ACK8_p & v93f1b4 | !BtoS_ACK8_p & !v909823;
assign v90d59a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v910243;
assign v90adef = StoB_REQ8_p & v87a1d0 | !StoB_REQ8_p & v9098e3;
assign v93f84d = StoB_REQ7_p & v9058f3 | !StoB_REQ7_p & v90ee83;
assign v886f59 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v911102;
assign v90d81c = BtoS_ACK6_p & v90787b | !BtoS_ACK6_p & v93fa28;
assign v93f202 = jx3_p & v908ad9 | !jx3_p & v90cf0e;
assign v93dade = StoB_REQ6_p & v93fa4f | !StoB_REQ6_p & v904b91;
assign v9061f2 = BtoS_ACK6_p & v9099ee | !BtoS_ACK6_p & v844f91;
assign v90e945 = StoB_REQ2_p & v90fe49 | !StoB_REQ2_p & !v844f91;
assign v910cf2 = jx1_p & v844f91 | !jx1_p & v93fa9d;
assign v908751 = ENQ_p & v90fbad | !ENQ_p & v93fe35;
assign v93e684 = BtoS_ACK1_p & v90fc92 | !BtoS_ACK1_p & v904995;
assign v8ee181 = BtoS_ACK1_p & v93fce7 | !BtoS_ACK1_p & v93ecb6;
assign v93e0a0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93ebb5;
assign v93f8ee = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & v9041e4;
assign v9083d0 = jx0_p & v90f2de | !jx0_p & v8633b7;
assign v85f258 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v91218a;
assign v87a1b7 = BtoS_ACK0_p & v911102 | !BtoS_ACK0_p & v93fb83;
assign v93fabd = BtoS_ACK6_p & v86344b | !BtoS_ACK6_p & v903d60;
assign v93fca7 = jx0_p & v90d6e8 | !jx0_p & v93f709;
assign v93ee1b = BtoS_ACK1_p & v93dfc0 | !BtoS_ACK1_p & v90ae72;
assign v93f7d7 = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & v907eaa;
assign v85dee0 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v910825;
assign v905d8b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90ad6c;
assign v90684c = StoB_REQ6_p & v911937 | !StoB_REQ6_p & v909649;
assign v93f927 = BtoS_ACK9_p & v93e228 | !BtoS_ACK9_p & !v90a2b5;
assign v90dc08 = ENQ_p & v9083cf | !ENQ_p & v905312;
assign v93e701 = BtoS_ACK8_p & v89e10d | !BtoS_ACK8_p & v93f776;
assign v93fe52 = jx0_p & v90f7d6 | !jx0_p & v844f91;
assign v906024 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v9095e0;
assign v93f4cd = jx1_p & v9093ec | !jx1_p & v91aa51;
assign v905ba4 = RtoB_ACK0_p & v909bdf | !RtoB_ACK0_p & v93e3f1;
assign v93fd55 = BtoS_ACK6_p & v90a216 | !BtoS_ACK6_p & v87f17d;
assign v904794 = DEQ_p & v93f8de | !DEQ_p & v908751;
assign v905a21 = BtoS_ACK8_p & v93fb68 | !BtoS_ACK8_p & v93fa3d;
assign v903db9 = jx2_p & v863b37 | !jx2_p & v90d879;
assign v87c4c4 = BtoS_ACK9_p & v9056a4 | !BtoS_ACK9_p & v93f6ab;
assign v91232c = BtoS_ACK0_p & v93f702 | !BtoS_ACK0_p & v93fb44;
assign v93f06e = BtoS_ACK7_p & v908073 | !BtoS_ACK7_p & !v93f785;
assign v90fb4b = jx0_p & v91a771 | !jx0_p & v844f91;
assign v863ad6 = BtoS_ACK8_p & v9074fa | !BtoS_ACK8_p & v93f6aa;
assign v93ea16 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9068fc;
assign v908836 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v93f9d2;
assign v870489 = BtoS_ACK6_p & v90cc30 | !BtoS_ACK6_p & v910473;
assign v8d3799 = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v910825;
assign v87010f = BtoS_ACK8_p & v93e7d1 | !BtoS_ACK8_p & !v91091b;
assign v91141d = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v93fb48;
assign BtoS_ACK1_n = !v8b6034;
assign v912265 = jx1_p & v93fc3e | !jx1_p & !v844f91;
assign v90f62b = jx3_p & v9109e6 | !jx3_p & !v91a6f1;
assign v93fced = BtoS_ACK8_p & v93ca43 | !BtoS_ACK8_p & v910db7;
assign v93f6a7 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v90ed3d;
assign v8b5f5d = BtoS_ACK6_p & v89f8bd | !BtoS_ACK6_p & v909be7;
assign v907bee = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & v93f6d2;
assign v93e589 = BtoS_ACK0_p & v906627 | !BtoS_ACK0_p & v90fcd2;
assign v907664 = RtoB_ACK1_p & v90517f | !RtoB_ACK1_p & v93f8b2;
assign v93f755 = jx2_p & v87c51f | !jx2_p & !v93fbb0;
assign v93fd19 = stateG7_1_p & v93e548 | !stateG7_1_p & v93e838;
assign v93e898 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88d074;
assign v93fd12 = StoB_REQ7_p & v87f17d | !StoB_REQ7_p & v907e7e;
assign v93f51d = jx1_p & v907be9 | !jx1_p & v93e2fa;
assign v8f229e = jx0_p & v93f9dd | !jx0_p & v8b9e12;
assign v90444f = jx3_p & v904b7f | !jx3_p & v90f5f8;
assign v93ee82 = BtoS_ACK0_p & v86c2d0 | !BtoS_ACK0_p & v90fe91;
assign v90965e = jx1_p & v909918 | !jx1_p & v9041e6;
assign v93fa55 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v90a5ef;
assign v93dffa = EMPTY_p & v93dfb4 | !EMPTY_p & v904794;
assign v87a261 = StoB_REQ7_p & v90ec5d | !StoB_REQ7_p & v912384;
assign v905540 = DEQ_p & v9087b7 | !DEQ_p & v93fa75;
assign v93fb21 = ENQ_p & v908325 | !ENQ_p & v844f91;
assign v913561 = StoB_REQ1_p & v913348 | !StoB_REQ1_p & v844f9d;
assign v90a2df = jx1_p & v93f1cf | !jx1_p & !v93fb3e;
assign v93ef40 = jx3_p & v93fdda | !jx3_p & v90930e;
assign v863a64 = RtoB_ACK0_p & v9082be | !RtoB_ACK0_p & v908df3;
assign v90604e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93f928;
assign v90e083 = BtoS_ACK2_p & v91305b | !BtoS_ACK2_p & v93fc01;
assign v93fc7e = jx0_p & v844f91 | !jx0_p & !v93f119;
assign v9101c0 = BtoS_ACK9_p & v9073c5 | !BtoS_ACK9_p & v93f7d3;
assign v90e3bf = jx3_p & v844f91 | !jx3_p & !v8b9f15;
assign v85ea51 = jx0_p & v844f91 | !jx0_p & v909b01;
assign v9107c7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v910c3a;
assign v93e9dd = RtoB_ACK1_p & v904dea | !RtoB_ACK1_p & v90f164;
assign v93f7c3 = StoB_REQ8_p & v907e81 | !StoB_REQ8_p & v85eaf3;
assign v904b94 = ENQ_p & v90834a | !ENQ_p & !v904677;
assign v90dec9 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fb66;
assign v89f8bd = jx0_p & v844f9f | !jx0_p & !v8b8638;
assign v907cc6 = jx0_p & v908805 | !jx0_p & v93f290;
assign v93f3f2 = jx3_p & v93f937 | !jx3_p & v90a23c;
assign v903b4e = EMPTY_p & v85eaa2 | !EMPTY_p & v909001;
assign v93f865 = StoB_REQ1_p & v90a0cb | !StoB_REQ1_p & v93fe06;
assign v90f575 = jx2_p & v8b9ee1 | !jx2_p & v90cbec;
assign v90a196 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v906acc;
assign v90d3cc = StoB_REQ6_p & v9081b9 | !StoB_REQ6_p & v905ca1;
assign v908d55 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93fd9c;
assign v93fb68 = jx2_p & v904779 | !jx2_p & v9075d4;
assign v93dc08 = jx1_p & v93f6a2 | !jx1_p & v93fa4c;
assign v905355 = stateG7_1_p & v93f870 | !stateG7_1_p & v863a7b;
assign v904c4f = ENQ_p & v844fc3 | !ENQ_p & !v844f91;
assign v88d074 = BtoS_ACK6_p & v93efbb | !BtoS_ACK6_p & v93faec;
assign v92ffb9 = BtoS_ACK1_p & v90a59e | !BtoS_ACK1_p & v9058f4;
assign v90e526 = StoB_REQ1_p & v90e945 | !StoB_REQ1_p & v90fe49;
assign v9384b0 = EMPTY_p & v91132a | !EMPTY_p & !v909dc3;
assign v913332 = StoB_REQ7_p & v87f17d | !StoB_REQ7_p & !v844f91;
assign v90e144 = BtoS_ACK7_p & v93fdd2 | !BtoS_ACK7_p & v93f755;
assign v90e2dc = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v89f7e2;
assign v89b107 = jx2_p & v844f91 | !jx2_p & v93f696;
assign v93fabf = BtoS_ACK6_p & v90db9f | !BtoS_ACK6_p & v907cc6;
assign v908a76 = jx3_p & v93fe30 | !jx3_p & !v844f91;
assign v910ff7 = BtoS_ACK6_p & v90671f | !BtoS_ACK6_p & v904de5;
assign v93fe30 = stateG12_p & v93fbfc | !stateG12_p & !v844f91;
assign v904ff8 = BtoS_ACK6_p & v904e70 | !BtoS_ACK6_p & v844f91;
assign v93fa0a = ENQ_p & v90fbad | !ENQ_p & v9110fe;
assign v90f161 = BtoS_ACK8_p & v911a72 | !BtoS_ACK8_p & v86ce77;
assign v9056b0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f871;
assign v90683e = BtoS_ACK7_p & v908410 | !BtoS_ACK7_p & v90ad9a;
assign v90a902 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v92ffda;
assign v908fb5 = BtoS_ACK7_p & v93fcd0 | !BtoS_ACK7_p & !v907a33;
assign v90667f = BtoS_ACK8_p & v93e370 | !BtoS_ACK8_p & v93fde6;
assign v907b01 = RtoB_ACK0_p & v93fde2 | !RtoB_ACK0_p & v93fb72;
assign v905204 = jx0_p & v844f91 | !jx0_p & v9091b2;
assign v93fc38 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v907b21;
assign v93f85d = jx1_p & v93e7d1 | !jx1_p & v844f91;
assign v90e9e1 = jx1_p & v844f91 | !jx1_p & !v844fbd;
assign v906038 = RtoB_ACK0_p & v90f304 | !RtoB_ACK0_p & v90f62b;
assign v90546e = BtoS_ACK8_p & v911a72 | !BtoS_ACK8_p & v9058d5;
assign v93fdb4 = BtoS_ACK6_p & v8b9b9f | !BtoS_ACK6_p & v93fd7f;
assign v8d37bd = BtoS_ACK6_p & v90cbf6 | !BtoS_ACK6_p & v906623;
assign v884fc2 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v904bbf;
assign v8b9c53 = jx1_p & v869aeb | !jx1_p & !v93f763;
assign v9132eb = jx2_p & v911973 | !jx2_p & v911941;
assign v90d866 = BtoS_ACK7_p & v909bbd | !BtoS_ACK7_p & !v9044c9;
assign v908ffc = DEQ_p & v91007f | !DEQ_p & v88c2af;
assign v93e168 = StoB_REQ8_p & v8ee1cd | !StoB_REQ8_p & v910d56;
assign v906d41 = StoB_REQ2_p & v8b98bd | !StoB_REQ2_p & !v844f91;
assign v93f7bb = StoB_REQ3_p & v907168 | !StoB_REQ3_p & v93f8f8;
assign v93e9d8 = BtoS_ACK7_p & v93e115 | !BtoS_ACK7_p & v907679;
assign v90748c = BtoS_ACK8_p & v93e115 | !BtoS_ACK8_p & v85ea93;
assign v86e625 = StoB_REQ9_p & v911cba | !StoB_REQ9_p & v93f6c1;
assign v911680 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v90fe49;
assign v909c3b = StoB_REQ9_p & v906c20 | !StoB_REQ9_p & v90efef;
assign v905697 = ENQ_p & v93fda6 | !ENQ_p & v86345f;
assign v903fa0 = StoB_REQ1_p & v93e9cc | !StoB_REQ1_p & v93f6ec;
assign v93f6b8 = BtoS_ACK0_p & v90855a | !BtoS_ACK0_p & !v9097b1;
assign v90539a = FULL_p & v93e301 | !FULL_p & v90e333;
assign v90d0b6 = BtoS_ACK1_p & v913348 | !BtoS_ACK1_p & v907472;
assign v912673 = BtoS_ACK7_p & v93fc5d | !BtoS_ACK7_p & v9043c7;
assign v93fc86 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v90e9f7;
assign v910383 = jx0_p & v93f70c | !jx0_p & !v93f685;
assign v93ec4d = jx1_p & v910710 | !jx1_p & v910d70;
assign v90e8da = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v913662;
assign v9096fd = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v90e251;
assign v93e370 = StoB_REQ8_p & v93fda1 | !StoB_REQ8_p & v90d5c7;
assign v8c737b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86c2d0;
assign v911ec2 = StoB_REQ2_p & v908127 | !StoB_REQ2_p & v910495;
assign v93f90e = jx0_p & v904340 | !jx0_p & v907a13;
assign v86ccf1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f85e;
assign v93fda8 = jx1_p & v87f17d | !jx1_p & !v844f91;
assign v93e70e = jx3_p & v844f91 | !jx3_p & v93f5d9;
assign v93fd4a = jx3_p & v93fbcc | !jx3_p & v91a70f;
assign v93efae = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v905467;
assign v93f9b9 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v93e51c;
assign v93f7be = jx1_p & v90901d | !jx1_p & v93fb24;
assign v9043bd = RtoB_ACK0_p & v90752d | !RtoB_ACK0_p & v90a07b;
assign v906492 = StoB_REQ1_p & v907bee | !StoB_REQ1_p & v8b9c2b;
assign v93f9da = EMPTY_p & v85eaa2 | !EMPTY_p & v93fd49;
assign v93fc93 = jx3_p & v93f110 | !jx3_p & v90d32d;
assign v93f282 = StoB_REQ8_p & v90d662 | !StoB_REQ8_p & v8f3874;
assign v90f7d3 = BtoS_ACK0_p & v913619 | !BtoS_ACK0_p & v9124c5;
assign v9082d3 = BtoS_ACK2_p & v9076a8 | !BtoS_ACK2_p & v91195c;
assign v93efb0 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v90acc5;
assign v93eba3 = jx2_p & v93f518 | !jx2_p & v905aaa;
assign v904c53 = ENQ_p & v85eaff | !ENQ_p & v93f1a6;
assign v907292 = RtoB_ACK0_p & v90dc08 | !RtoB_ACK0_p & v863ac4;
assign v93e713 = StoB_REQ7_p & v89f920 | !StoB_REQ7_p & v910f4e;
assign v9115ab = StoB_REQ0_p & v93fd87 | !StoB_REQ0_p & v93fb8c;
assign v93fc06 = StoB_REQ6_p & v909d18 | !StoB_REQ6_p & v8b9e6b;
assign v93f6d0 = ENQ_p & v844fc3 | !ENQ_p & !v93e682;
assign v93fe66 = jx1_p & v844f91 | !jx1_p & v93f796;
assign v93fa46 = BtoS_ACK6_p & v906d58 | !BtoS_ACK6_p & v844f91;
assign v8660c5 = RtoB_ACK1_p & v87ca3a | !RtoB_ACK1_p & v8b6009;
assign v907eaa = jx1_p & v91a9de | !jx1_p & !v844f91;
assign v9099ee = jx0_p & v93f63b | !jx0_p & v904adb;
assign v87a1f0 = jx1_p & v90a850 | !jx1_p & v9049a9;
assign v8b4983 = jx1_p & v93ec9d | !jx1_p & v9132d6;
assign v93e95e = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v87c9f1;
assign v9095bf = jx0_p & v910243 | !jx0_p & !v90893a;
assign v8f3879 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v9072b4;
assign v90eed2 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v93fd11;
assign v93f293 = BtoS_ACK6_p & v884481 | !BtoS_ACK6_p & v9052ef;
assign v90767a = StoB_REQ6_p & v89f9d7 | !StoB_REQ6_p & v844f91;
assign v93fb38 = jx2_p & v93e76f | !jx2_p & v90da8b;
assign v93dc29 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93fc17;
assign v910910 = jx0_p & v844f91 | !jx0_p & v8b49ad;
assign v911552 = BtoS_ACK7_p & v910fda | !BtoS_ACK7_p & v9109f4;
assign v93df55 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f8c3;
assign v93f9fe = EMPTY_p & v93eb1d | !EMPTY_p & v910d2f;
assign v90752a = jx0_p & v90d6e8 | !jx0_p & !v844f91;
assign v909e28 = jx2_p & v90a2fc | !jx2_p & v93fdfd;
assign v913632 = BtoS_ACK9_p & v8b5f61 | !BtoS_ACK9_p & v908515;
assign v903c4d = BtoS_ACK7_p & v904b00 | !BtoS_ACK7_p & v905775;
assign v8b99b9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fcb7;
assign v93f9f6 = BtoS_ACK7_p & v85f240 | !BtoS_ACK7_p & v912265;
assign v907ad8 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v9115ab;
assign v93fc3d = BtoS_ACK6_p & v93e681 | !BtoS_ACK6_p & v92ffd9;
assign v93fc29 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91db5a;
assign v906627 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v9123a2;
assign v8b9e82 = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v93dfc0;
assign v8f22ee = jx0_p & v844f91 | !jx0_p & !v906623;
assign v93e5e5 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v9080a8;
assign v88dbe7 = jx1_p & v93f136 | !jx1_p & v844f91;
assign v93f6ab = StoB_REQ9_p & v90f9f3 | !StoB_REQ9_p & v90f3f8;
assign v93f9e3 = jx1_p & v863b25 | !jx1_p & v844f91;
assign v907e7e = jx0_p & v844f91 | !jx0_p & v93f119;
assign v910117 = BtoS_ACK1_p & v90fc92 | !BtoS_ACK1_p & v906bf5;
assign v93fc22 = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v909430;
assign v910289 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v844fa5;
assign v907f31 = jx1_p & v910f4e | !jx1_p & v93e713;
assign v9095d0 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v93fd0d;
assign v93f7e8 = BtoS_ACK6_p & v8a9289 | !BtoS_ACK6_p & v844f91;
assign v90a588 = StoB_REQ9_p & v903ddc | !StoB_REQ9_p & v90e88f;
assign v904fee = ENQ_p & v844fc3 | !ENQ_p & !v93f90f;
assign v903e85 = StoB_REQ6_p & v93e681 | !StoB_REQ6_p & v844f91;
assign v90666d = StoB_REQ8_p & v90dab9 | !StoB_REQ8_p & v93fb7f;
assign v93f511 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v93fc34;
assign v8b49dc = jx1_p & v869aeb | !jx1_p & !v9040cd;
assign v90441d = BtoS_ACK6_p & v871df8 | !BtoS_ACK6_p & v93f8a5;
assign v90d22a = jx1_p & v913522 | !jx1_p & !v907017;
assign v93e577 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f70c;
assign v93f972 = BtoS_ACK7_p & v8b9ee2 | !BtoS_ACK7_p & v93f320;
assign v93fc66 = jx3_p & v93fa7d | !jx3_p & !v93fc86;
assign v93f70a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93efb0;
assign v87a2ad = BtoS_ACK1_p & v93f85e | !BtoS_ACK1_p & v90a97c;
assign v93f8b7 = jx0_p & v90d3cc | !jx0_p & !v910081;
assign v91143a = BtoS_ACK7_p & v93de99 | !BtoS_ACK7_p & v9102aa;
assign v8b9c07 = jx0_p & v93f793 | !jx0_p & v844f91;
assign v93fe39 = stateG12_p & v93eed6 | !stateG12_p & v90d9b3;
assign v90a9fc = BtoS_ACK9_p & v93f8e0 | !BtoS_ACK9_p & v87575e;
assign v93f57d = jx0_p & v904f5c | !jx0_p & v93fa6d;
assign v93faa8 = jx1_p & v9061f2 | !jx1_p & v905ba8;
assign v90e1c3 = StoB_REQ9_p & v903fc8 | !StoB_REQ9_p & v90e373;
assign v905838 = BtoS_ACK7_p & v93f588 | !BtoS_ACK7_p & !v9045b2;
assign v9085c8 = jx0_p & v90d364 | !jx0_p & !v93f707;
assign v907d8f = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9042fa;
assign v844fbf = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844f91;
assign v93f680 = FULL_p & v844f91 | !FULL_p & v905397;
assign v90accf = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9124bc;
assign v9102bb = DEQ_p & v904d40 | !DEQ_p & v85ea72;
assign v93fe47 = ENQ_p & v844f91 | !ENQ_p & v93f80a;
assign v9100b7 = StoB_REQ8_p & v91071f | !StoB_REQ8_p & v93fa4d;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v93f4e9 = BtoS_ACK7_p & v93ed2a | !BtoS_ACK7_p & v9124ae;
assign v863476 = jx1_p & v9062f7 | !jx1_p & v904e38;
assign v88d7c9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93e9ea;
assign v90809d = jx0_p & v844f91 | !jx0_p & !v93fcea;
assign v911417 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v907f05;
assign v909941 = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v93f70a;
assign v9051c9 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v9052de;
assign v93faf4 = RtoB_ACK0_p & v89f796 | !RtoB_ACK0_p & v90539a;
assign v90d727 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v913449;
assign v93fe14 = BtoS_ACK6_p & v884481 | !BtoS_ACK6_p & v911d8e;
assign v93e791 = jx2_p & v90d9b2 | !jx2_p & !v9124a9;
assign v93f97e = jx2_p & v905dcf | !jx2_p & v93fb73;
assign v91e95f = jx3_p & v93f78c | !jx3_p & !v93fd6c;
assign v90a91e = StoB_REQ0_p & v906642 | !StoB_REQ0_p & v93e602;
assign v872067 = BtoS_ACK6_p & v9099ee | !BtoS_ACK6_p & v93ef57;
assign v913169 = jx1_p & v8b9f37 | !jx1_p & !v844f91;
assign v910f51 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9041e4;
assign v93fc47 = jx2_p & v844f91 | !jx2_p & !v93f9c7;
assign v93f86b = BtoS_ACK8_p & v93e27a | !BtoS_ACK8_p & v906915;
assign v87a991 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fe27;
assign v93ecf7 = BtoS_ACK8_p & v93fb93 | !BtoS_ACK8_p & v91247e;
assign v9114a0 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8b9dff;
assign v90ad47 = jx0_p & v90ea74 | !jx0_p & v844f91;
assign v910469 = jx0_p & v90eef9 | !jx0_p & v93f895;
assign v8b9d49 = jx0_p & v912d1c | !jx0_p & !v908816;
assign v93fe41 = BtoS_ACK0_p & v93f5d1 | !BtoS_ACK0_p & v906d38;
assign v89f97d = StoB_REQ8_p & v904b00 | !StoB_REQ8_p & v93e855;
assign v90e988 = StoB_REQ9_p & v8d37d4 | !StoB_REQ9_p & v93fe5a;
assign v92ffda = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v90d9fd;
assign v93fc15 = jx2_p & v93e310 | !jx2_p & v93f860;
assign v93f73d = jx2_p & v90e94e | !jx2_p & v90cbec;
assign v86337d = BtoS_ACK6_p & v93fb3e | !BtoS_ACK6_p & v91268a;
assign v906c0c = ENQ_p & v93f89f | !ENQ_p & v906e30;
assign v93f901 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93fc84;
assign v93f27f = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & !v85ea62;
assign v903c5b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f67b;
assign v8bb868 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v844f91;
assign v90f79b = BtoS_ACK0_p & v93e295 | !BtoS_ACK0_p & v903aff;
assign v93f6a0 = jx1_p & v9099e1 | !jx1_p & v844f91;
assign v90f383 = jx2_p & v8b9c53 | !jx2_p & v90986f;
assign v93fcfe = stateG12_p & v93f89f | !stateG12_p & v93fda9;
assign v9054e2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f8b9;
assign v9098b1 = jx0_p & v93fda0 | !jx0_p & !v844f91;
assign v90ad02 = BtoS_ACK6_p & v9096ae | !BtoS_ACK6_p & v904520;
assign v903e62 = jx0_p & v906c6e | !jx0_p & !v907a13;
assign v90441e = BtoS_ACK9_p & v93e048 | !BtoS_ACK9_p & v87c534;
assign v91a9e1 = jx0_p & v906d08 | !jx0_p & !v93dfe2;
assign v93faf1 = BtoS_ACK6_p & v93fa7c | !BtoS_ACK6_p & v844f91;
assign v886fce = ENQ_p & v844f91 | !ENQ_p & !v93fad0;
assign v93ecb6 = StoB_REQ1_p & v904ae0 | !StoB_REQ1_p & v91003a;
assign v90f1ab = jx1_p & v906201 | !jx1_p & !v9045fa;
assign v9104bd = StoB_REQ9_p & v90ee4b | !StoB_REQ9_p & v913a64;
assign v90878b = BtoS_ACK8_p & v91a799 | !BtoS_ACK8_p & v9079f4;
assign v904520 = jx0_p & v912d1c | !jx0_p & !v93f922;
assign v90819e = BtoS_ACK9_p & v9073c5 | !BtoS_ACK9_p & v86eecd;
assign v912d1c = BtoS_ACK0_p & v93e295 | !BtoS_ACK0_p & v908636;
assign v90855a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v906255;
assign v9082a3 = StoB_REQ7_p & v8a8b0a | !StoB_REQ7_p & v93ec50;
assign v93fa51 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v87010f;
assign v93fd90 = BtoS_ACK8_p & v93ca43 | !BtoS_ACK8_p & v91336c;
assign v90664a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v9054b5;
assign v90eef5 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v89fe59;
assign v912fa9 = BtoS_ACK6_p & v86344b | !BtoS_ACK6_p & v906fec;
assign v93fbe2 = StoB_REQ6_p & v9054b5 | !StoB_REQ6_p & v906a51;
assign BtoS_ACK8_n = !v8b99c6;
assign v93fe15 = DEQ_p & v90a07b | !DEQ_p & v904dfc;
assign v8d37be = ENQ_p & v9083cf | !ENQ_p & v93f892;
assign v904b4f = BtoS_ACK6_p & v910f82 | !BtoS_ACK6_p & v8b9c07;
assign v93fd6f = StoB_REQ6_p & v93e97c | !StoB_REQ6_p & v87a1b7;
assign v903fac = BtoS_ACK7_p & v90f575 | !BtoS_ACK7_p & v90738d;
assign v89fdce = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9045f3;
assign v930099 = StoB_REQ8_p & v904ab4 | !StoB_REQ8_p & v93e4b9;
assign v9118ff = StoB_REQ9_p & v903eef | !StoB_REQ9_p & v907ff8;
assign v90e3e1 = jx0_p & v844f91 | !jx0_p & v913435;
assign v93f8d0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a6ae;
assign v90ae1b = BtoS_ACK7_p & v903afe | !BtoS_ACK7_p & v93fcc2;
assign v8b9c3f = BtoS_ACK1_p & v906255 | !BtoS_ACK1_p & !v906c48;
assign v93fc67 = StoB_REQ8_p & v90ea47 | !StoB_REQ8_p & v910d28;
assign v93f95a = jx3_p & v91a796 | !jx3_p & v93f15e;
assign v903e8d = StoB_REQ6_p & v90aaca | !StoB_REQ6_p & v93fc0e;
assign v93f110 = stateG12_p & v905539 | !stateG12_p & !v93f78c;
assign v93ec44 = StoB_REQ6_p & v90f9be | !StoB_REQ6_p & v903df5;
assign v93fb1a = StoB_REQ0_p & v93f70c | !StoB_REQ0_p & v9054c9;
assign v90a8cd = BtoS_ACK0_p & v93fc02 | !BtoS_ACK0_p & v93f9c5;
assign v909337 = jx1_p & v93fd51 | !jx1_p & v844f91;
assign v906c94 = jx0_p & v93f689 | !jx0_p & !v844f91;
assign v89e122 = jx2_p & v93f9a1 | !jx2_p & v90cbec;
assign v9132d3 = BtoS_ACK7_p & v90dec8 | !BtoS_ACK7_p & !v8b9cd2;
assign v90fe91 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fb31;
assign v93f90d = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v9080b4;
assign v93f9e0 = RtoB_ACK0_p & v906c0c | !RtoB_ACK0_p & v904ef7;
assign v93fca3 = jx0_p & v93fe1e | !jx0_p & !v9056ad;
assign v93e203 = RtoB_ACK0_p & v9051ba | !RtoB_ACK0_p & v907301;
assign v9075d4 = jx1_p & v9072c8 | !jx1_p & !v909f4c;
assign v911451 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v86313d;
assign v91132a = ENQ_p & v93f8ad | !ENQ_p & v90ee7e;
assign v90d731 = BtoS_ACK9_p & v93f76e | !BtoS_ACK9_p & v8880f2;
assign v93fbd7 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v91062b;
assign v905810 = jx2_p & v844f91 | !jx2_p & v93f148;
assign v904ba4 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93f979;
assign v8b9c87 = jx1_p & v844f91 | !jx1_p & !v93fe0c;
assign v9104ad = jx2_p & v904234 | !jx2_p & !v9060ea;
assign v87c52b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9041fc;
assign v93fd8e = BtoS_ACK4_p & v844f9f | !BtoS_ACK4_p & v90f547;
assign v90a4d4 = jx3_p & v905a12 | !jx3_p & v908325;
assign v8739eb = StoB_REQ9_p & v93faef | !StoB_REQ9_p & v93fc1f;
assign v90aca4 = StoB_REQ9_p & v8d37d4 | !StoB_REQ9_p & v93fa05;
assign v908743 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ee188;
assign v93f681 = jx0_p & v844f91 | !jx0_p & !v90690e;
assign v908068 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844fb7;
assign v93fa86 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v905841;
assign v91058e = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v844f9f;
assign v93fc16 = RtoB_ACK1_p & v90e770 | !RtoB_ACK1_p & v93f6a9;
assign v93fcf4 = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v904e53;
assign v93f87b = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v911c0f;
assign v91a6d3 = jx3_p & v93ec1d | !jx3_p & v93f753;
assign v89e11b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8a8f74;
assign v93fdf3 = StoB_REQ8_p & v93f960 | !StoB_REQ8_p & !v908e75;
assign v91268b = RtoB_ACK1_p & v93fb1b | !RtoB_ACK1_p & v904f22;
assign v8b5f61 = jx2_p & v906c8b | !jx2_p & v9060ea;
assign v93fdfa = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v910bd7;
assign v93fc17 = BtoS_ACK7_p & v9074ce | !BtoS_ACK7_p & v85ead8;
assign v92fffd = ENQ_p & v93f753 | !ENQ_p & v93ef40;
assign v9044a5 = jx0_p & v90e133 | !jx0_p & v93e5bf;
assign v87a671 = StoB_REQ7_p & v93f8a6 | !StoB_REQ7_p & v8b5f5d;
assign v9068fc = jx1_p & v844f91 | !jx1_p & v93fb3a;
assign v907061 = BtoR_REQ0_p & v918886 | !BtoR_REQ0_p & v91090e;
assign v910bf8 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v905da3;
assign v872442 = BtoS_ACK8_p & v903d0c | !BtoS_ACK8_p & !v904bcb;
assign v9043b9 = StoB_REQ8_p & v93fb43 | !StoB_REQ8_p & v9101ae;
assign v91dd4f = StoB_REQ0_p & v93fd87 | !StoB_REQ0_p & v90f320;
assign v9080a0 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v93fddd;
assign v93fc0b = BtoS_ACK8_p & v93fdae | !BtoS_ACK8_p & v93fc18;
assign v91148d = jx1_p & v911edb | !jx1_p & v905d7e;
assign v907683 = StoB_REQ8_p & v90f5bd | !StoB_REQ8_p & v91051a;
assign v93fd20 = BtoS_ACK6_p & v8a9222 | !BtoS_ACK6_p & v844f91;
assign v912f16 = StoB_REQ2_p & v87c537 | !StoB_REQ2_p & v93e5e5;
assign v93eaa1 = BtoS_ACK7_p & v9074ce | !BtoS_ACK7_p & v93f7c9;
assign v907b6c = BtoS_ACK7_p & v903db9 | !BtoS_ACK7_p & v910d41;
assign v911c11 = BtoS_ACK6_p & v909f04 | !BtoS_ACK6_p & v93fdce;
assign v93f81c = BtoS_ACK0_p & v91a9cd | !BtoS_ACK0_p & v9108ff;
assign v93e295 = StoB_REQ1_p & v86c2d0 | !StoB_REQ1_p & v93dfc0;
assign v907e81 = jx2_p & v844f91 | !jx2_p & !v904755;
assign v89f7c7 = BtoS_ACK7_p & v93e259 | !BtoS_ACK7_p & v87c4e7;
assign v90521f = BtoS_ACK1_p & v93e356 | !BtoS_ACK1_p & v9132d4;
assign v85eaf3 = jx2_p & v90fa0b | !jx2_p & !v904755;
assign v91aa12 = BtoS_ACK1_p & v93deab | !BtoS_ACK1_p & v90ebcd;
assign v90e958 = ENQ_p & v93f95a | !ENQ_p & v844f91;
assign v90aa3b = StoB_REQ8_p & v93fb78 | !StoB_REQ8_p & v93f6fb;
assign v93f6d2 = StoB_REQ2_p & v93fd5c | !StoB_REQ2_p & v93f928;
assign v90719c = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v904cde;
assign v90a884 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v93ecb0;
assign v93e8f1 = jx3_p & v9113c0 | !jx3_p & v93fbb4;
assign v93f6cc = jx0_p & v91a6d1 | !jx0_p & v844f91;
assign v8ee1a9 = EMPTY_p & v93eef4 | !EMPTY_p & v911951;
assign v873ad7 = jx1_p & v93f1cf | !jx1_p & !v844f91;
assign v8d37d8 = jx1_p & v911edb | !jx1_p & v90a7ea;
assign v9114cf = DEQ_p & v9048c6 | !DEQ_p & v93e203;
assign v908bf7 = BtoS_ACK6_p & v90cc30 | !BtoS_ACK6_p & v90e76a;
assign v90f83a = jx2_p & v863a47 | !jx2_p & v93f6ea;
assign v90944f = BtoS_ACK7_p & v93fbe4 | !BtoS_ACK7_p & v904b04;
assign v91003b = jx1_p & v90d879 | !jx1_p & v90f78a;
assign v90efef = BtoS_ACK8_p & v93fb66 | !BtoS_ACK8_p & v93f78f;
assign v9043e5 = jx2_p & v93e535 | !jx2_p & v87f17d;
assign v9095df = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v93f521;
assign v93fc35 = BtoS_ACK8_p & v904b00 | !BtoS_ACK8_p & v93eb39;
assign v863a03 = jx1_p & v869aeb | !jx1_p & !v90998d;
assign v907301 = FULL_p & v907b84 | !FULL_p & v87d990;
assign v870bc2 = BtoS_ACK8_p & v93f9bb | !BtoS_ACK8_p & v906663;
assign v905803 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fb6f;
assign v93ef30 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v908a34;
assign v93e230 = BtoR_REQ0_p & v913225 | !BtoR_REQ0_p & v90710d;
assign v93fb00 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v905b5d;
assign v93fe2b = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & v913348;
assign v93fc85 = BtoS_ACK7_p & v907adb | !BtoS_ACK7_p & v9109dc;
assign v904a0b = jx1_p & v869aeb | !jx1_p & !v90e341;
assign v93ed00 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v906627;
assign v93f70c = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v90600b = EMPTY_p & v9083b1 | !EMPTY_p & !v93e3dd;
assign v870615 = jx0_p & v93e648 | !jx0_p & !v905665;
assign v90a2f1 = ENQ_p & v93eed6 | !ENQ_p & v906d80;
assign v90ad77 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v913348;
assign v904838 = BtoS_ACK7_p & v907e81 | !BtoS_ACK7_p & v93e1dd;
assign v90a29a = BtoS_ACK0_p & v90a6f4 | !BtoS_ACK0_p & v93f6d3;
assign v93ec1d = stateG12_p & v93f753 | !stateG12_p & !v93f7e6;
assign v9100ff = jx0_p & v93f895 | !jx0_p & !v90cc30;
assign v9089ef = DEQ_p & v909d90 | !DEQ_p & v93fc6c;
assign v93fde2 = ENQ_p & v90fbad | !ENQ_p & v93f492;
assign v9047f0 = BtoS_ACK6_p & v93f1cf | !BtoS_ACK6_p & v8ebce4;
assign v907607 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9099e1;
assign v904725 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8d37c1;
assign v911150 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v93e32d;
assign v93f785 = jx2_p & v8b4a13 | !jx2_p & v93f7be;
assign v93fb85 = jx3_p & v908429 | !jx3_p & v93fa2e;
assign v86dc4b = jx2_p & v8b9f38 | !jx2_p & !v912291;
assign v93f783 = ENQ_p & v912477 | !ENQ_p & v909dc5;
assign v93fcad = StoB_REQ7_p & v90f1b8 | !StoB_REQ7_p & v908bf7;
assign v93e704 = jx3_p & v9084d0 | !jx3_p & !v910545;
assign v910dda = jx2_p & v93f51d | !jx2_p & v907f0e;
assign v93fb8c = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93fb8f;
assign v93e8cb = jx2_p & v93e76f | !jx2_p & v9075d4;
assign v90648f = BtoS_ACK6_p & v9099fa | !BtoS_ACK6_p & v93f7d2;
assign v9080a7 = BtoS_ACK6_p & v9072c8 | !BtoS_ACK6_p & v844f91;
assign v93f89f = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v87a253;
assign v93eec9 = DEQ_p & v905b92 | !DEQ_p & v907bd4;
assign v90eea6 = BtoS_ACK9_p & v93db12 | !BtoS_ACK9_p & v93fd4f;
assign v907710 = StoB_REQ8_p & v903c4d | !StoB_REQ8_p & v907b6c;
assign v9072c8 = jx0_p & v871033 | !jx0_p & v90937e;
assign v910ee7 = jx2_p & v904926 | !jx2_p & v90962d;
assign v906af3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93f965;
assign v93e838 = RtoB_ACK0_p & v9103e5 | !RtoB_ACK0_p & v9042d2;
assign v9135b9 = jx1_p & v93fc7e | !jx1_p & v87f17d;
assign v908eba = StoB_REQ6_p & v9132e5 | !StoB_REQ6_p & v89c5e3;
assign v87c9b1 = BtoS_ACK2_p & v906cc8 | !BtoS_ACK2_p & v90ee63;
assign v930005 = jx1_p & v872067 | !jx1_p & v89fe58;
assign v9064cc = DEQ_p & v904d40 | !DEQ_p & v90e361;
assign v904f93 = ENQ_p & v911944 | !ENQ_p & v908a76;
assign v93fe37 = jx0_p & v9068b6 | !jx0_p & v9133d2;
assign v904f85 = StoB_REQ7_p & v910d5a | !StoB_REQ7_p & v93fa66;
assign v909efe = BtoR_REQ0_p & v93f9fe | !BtoR_REQ0_p & v904e3e;
assign v8bbc68 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fc71;
assign v909928 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v905c01;
assign v93df39 = StoB_REQ3_p & v93fd8e | !StoB_REQ3_p & v93e00f;
assign v93f80d = jx2_p & v90441c | !jx2_p & v85f243;
assign v93fdb1 = RtoB_ACK0_p & v93dfb4 | !RtoB_ACK0_p & v90828a;
assign v93da97 = BtoS_ACK9_p & v9043b9 | !BtoS_ACK9_p & v90a588;
assign v909119 = jx0_p & v844f91 | !jx0_p & v905ffe;
assign v909f4c = jx0_p & v844f97 | !jx0_p & !v93fcbe;
assign v8b9996 = RtoB_ACK0_p & v907b60 | !RtoB_ACK0_p & v90444d;
assign v907417 = jx3_p & v844f91 | !jx3_p & !v863428;
assign v8b98fe = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & !v90fa41;
assign v9131d1 = StoB_REQ9_p & v93f6b7 | !StoB_REQ9_p & v93fe5f;
assign v93f796 = BtoS_ACK6_p & v9058f3 | !BtoS_ACK6_p & v90460c;
assign v86341e = ENQ_p & v8a1fe3 | !ENQ_p & v93fb85;
assign v93f6a4 = jx1_p & v91ae94 | !jx1_p & v9093db;
assign v9059d6 = BtoS_ACK7_p & v90e40b | !BtoS_ACK7_p & v93fda3;
assign v8a9222 = jx0_p & v93ed91 | !jx0_p & v93f2a0;
assign v8b9c52 = BtoS_ACK8_p & v909366 | !BtoS_ACK8_p & !v90e2e7;
assign v93faad = jx1_p & v93fd43 | !jx1_p & !v904f88;
assign v89f920 = BtoS_ACK6_p & v93f9c6 | !BtoS_ACK6_p & v844f91;
assign v909078 = StoB_REQ3_p & v905702 | !StoB_REQ3_p & !v844f91;
assign v8f22e0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9088de;
assign v907717 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v904ef2;
assign v93fa80 = jx1_p & v907d70 | !jx1_p & !v882135;
assign v90879a = StoB_REQ7_p & v9093ec | !StoB_REQ7_p & !v844f91;
assign v90faf9 = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v87a25e;
assign v93fb4f = EMPTY_p & v93f26c | !EMPTY_p & v906fcc;
assign v93fb36 = jx0_p & v863b25 | !jx0_p & v904de5;
assign v879731 = BtoS_ACK8_p & v930076 | !BtoS_ACK8_p & v90d7cb;
assign v904f1a = BtoS_ACK2_p & v9076a8 | !BtoS_ACK2_p & v93fac5;
assign v93f5ff = BtoS_ACK8_p & v909367 | !BtoS_ACK8_p & !v907683;
assign v8b9c2c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fb27;
assign v89f9e4 = BtoR_REQ1_p & v93fcc0 | !BtoR_REQ1_p & v93db04;
assign v909a70 = BtoS_ACK8_p & v910b7a | !BtoS_ACK8_p & !v8b9ba5;
assign v89e12f = BtoR_REQ1_p & v91268b | !BtoR_REQ1_p & v8b9ec2;
assign v907ce3 = jx0_p & v93f8bb | !jx0_p & !v910243;
assign v906d3f = BtoS_ACK6_p & v871033 | !BtoS_ACK6_p & v8f37f3;
assign v93fd0d = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v90decf;
assign v8b9d25 = BtoS_ACK8_p & v90cf52 | !BtoS_ACK8_p & v907d8f;
assign v90a1fe = BtoS_ACK9_p & v90e893 | !BtoS_ACK9_p & v906e3b;
assign v907d9d = EMPTY_p & v907bd1 | !EMPTY_p & v904d7e;
assign v90ada1 = jx0_p & v9103b5 | !jx0_p & v911b4d;
assign v906ac6 = StoB_REQ9_p & v93ee39 | !StoB_REQ9_p & v93fd90;
assign v93fb5e = jx0_p & v9074ce | !jx0_p & v904f5c;
assign v905971 = jx0_p & v90762a | !jx0_p & v910243;
assign v90752d = ENQ_p & v90a4d4 | !ENQ_p & v93e8f1;
assign v8b9cd2 = jx2_p & v93f76d | !jx2_p & v907bbb;
assign v907472 = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & !v90827d;
assign v903e7f = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v910f51;
assign v93f1b4 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v93f119;
assign v93f584 = BtoS_ACK8_p & v93e855 | !BtoS_ACK8_p & v90417d;
assign v93ea75 = jx1_p & v9088ff | !jx1_p & v905194;
assign v90775f = stateG7_1_p & v92fffd | !stateG7_1_p & v863a00;
assign v908f29 = StoB_REQ1_p & v90a233 | !StoB_REQ1_p & v844f91;
assign v93fc01 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93f8a2;
assign v904fe6 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8f381b;
assign v907321 = DEQ_p & v9043bd | !DEQ_p & v907f74;
assign v93f883 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fddc;
assign v904e3a = ENQ_p & v844fc3 | !ENQ_p & !v93fd4a;
assign v9043fa = jx1_p & v905038 | !jx1_p & !v9112d5;
assign v93f1aa = jx1_p & v93e77d | !jx1_p & !v844f91;
assign v90414b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8bb868;
assign v8633c3 = jx2_p & v90eece | !jx2_p & !v90a149;
assign v93fba3 = BtoS_ACK7_p & v93dab8 | !BtoS_ACK7_p & v910b21;
assign v907c8c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b9c2b;
assign v90deff = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v90534f;
assign v906dea = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91a9b9;
assign v93de80 = jx0_p & v844f91 | !jx0_p & !v904725;
assign v9133f0 = StoB_REQ6_p & v93e835 | !StoB_REQ6_p & v9096f7;
assign v93f9ef = DEQ_p & v90d057 | !DEQ_p & v89e0d5;
assign v93f66f = StoB_REQ8_p & v93fc04 | !StoB_REQ8_p & v93fb68;
assign v90a6ae = BtoS_ACK6_p & v93fa7c | !BtoS_ACK6_p & v89e0ce;
assign v905396 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v905702;
assign v910e17 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v93e2e6;
assign v909f63 = jx2_p & v9054a2 | !jx2_p & v90d879;
assign v87c51f = jx1_p & v869aeb | !jx1_p & v844f91;
assign v90e8fd = jx1_p & v904ec6 | !jx1_p & !v844f91;
assign v89f95b = jx3_p & v844f91 | !jx3_p & v93fda4;
assign v93f6ed = BtoS_ACK7_p & v93fd84 | !BtoS_ACK7_p & v90e8fd;
assign v93f8a1 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v911b43;
assign v930109 = StoB_REQ6_p & v90a485 | !StoB_REQ6_p & v86deed;
assign v9081b9 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v909525;
assign v89f92f = StoB_REQ1_p & v90a47f | !StoB_REQ1_p & v90d698;
assign v93f70d = BtoS_ACK6_p & v93e89f | !BtoS_ACK6_p & v930037;
assign v905d66 = jx0_p & v9081b9 | !jx0_p & !v93f888;
assign v90a6ac = jx2_p & v90a3da | !jx2_p & v93fa1e;
assign v93fa3d = StoB_REQ8_p & v87c525 | !StoB_REQ8_p & v903c81;
assign v9091c7 = StoB_REQ1_p & v905660 | !StoB_REQ1_p & v93fb00;
assign v93f73c = ENQ_p & v911a33 | !ENQ_p & v9105f4;
assign v9045e6 = jx1_p & v844f91 | !jx1_p & v93fcf1;
assign v93f71d = StoB_REQ7_p & v905ba8 | !StoB_REQ7_p & v910f4e;
assign v93f918 = EMPTY_p & v93fd19 | !EMPTY_p & v903bf8;
assign v90a8ac = jx2_p & v90e38d | !jx2_p & v907383;
assign v90a8c3 = StoB_REQ1_p & v90611f | !StoB_REQ1_p & v844f91;
assign v909366 = jx1_p & v93f1b4 | !jx1_p & v87f17d;
assign v89e108 = jx2_p & v904bd4 | !jx2_p & v86f5de;
assign v9052de = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9b;
assign v903bf8 = DEQ_p & v905ba4 | !DEQ_p & v9042d2;
assign v93f050 = BtoS_ACK8_p & v93fb66 | !BtoS_ACK8_p & v90824e;
assign v93e8d3 = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v905978;
assign v911a92 = EMPTY_p & v9097bf | !EMPTY_p & v93fa06;
assign v90ef1b = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v9052de;
assign v9104d5 = jx1_p & v91ae94 | !jx1_p & v9078b3;
assign v8b9ec2 = RtoB_ACK1_p & v93f65b | !RtoB_ACK1_p & v908ef9;
assign v903fe9 = BtoS_ACK6_p & v9096ae | !BtoS_ACK6_p & v889a9e;
assign v92fff5 = BtoS_ACK9_p & v93e168 | !BtoS_ACK9_p & v93e0fb;
assign v93f7d5 = RtoB_ACK0_p & v9049ac | !RtoB_ACK0_p & v93f75f;
assign v93fbcd = jx3_p & v93fd59 | !jx3_p & !v93fb2a;
assign v90575f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90d0b6;
assign v93facb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fc64;
assign v90a07e = jx2_p & v90a314 | !jx2_p & v87f17d;
assign v911312 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fe4c;
assign v907069 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b49ad;
assign v908000 = jx0_p & v909e2c | !jx0_p & v85f258;
assign v908d10 = jx1_p & v844f91 | !jx1_p & v88932d;
assign v93fda0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v91a771;
assign v93fb29 = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v9054c6;
assign v87283f = StoB_REQ6_p & v90f9be | !StoB_REQ6_p & v90ad77;
assign v91023b = jx0_p & v906d08 | !jx0_p & v9056ad;
assign v93f8b9 = BtoS_ACK1_p & v90da97 | !BtoS_ACK1_p & v93fcd5;
assign v93f751 = stateG12_p & v93f753 | !stateG12_p & v93fc24;
assign v90a175 = jx1_p & v844f91 | !jx1_p & v91a9b9;
assign v93fa7e = jx1_p & v93f1b4 | !jx1_p & !v93fd12;
assign v905b5d = StoB_REQ2_p & v93fdf7 | !StoB_REQ2_p & v90ad48;
assign v908d2a = jx0_p & v904f5c | !jx0_p & v844f91;
assign v905e43 = jx2_p & v906d4c | !jx2_p & !v844f91;
assign v90ef07 = EMPTY_p & v906eb2 | !EMPTY_p & v93fe15;
assign v93ebbb = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v90667f;
assign v90add9 = BtoS_ACK9_p & v8b9bd8 | !BtoS_ACK9_p & v905a88;
assign v93faf7 = jx1_p & v93fe14 | !jx1_p & v93f7fb;
assign v90aa64 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v908d1f;
assign v93fb1b = EMPTY_p & v904b8c | !EMPTY_p & v93f9ef;
assign v93fd13 = DEQ_p & v905b92 | !DEQ_p & v907685;
assign v904f76 = RtoB_ACK1_p & v90f2f8 | !RtoB_ACK1_p & v907ccf;
assign v8a8f6f = jx1_p & v9093ec | !jx1_p & v87f17d;
assign v913a39 = BtoS_ACK6_p & v93f910 | !BtoS_ACK6_p & v906c94;
assign v93f8e4 = StoB_REQ6_p & v93e7c2 | !StoB_REQ6_p & v90a1f7;
assign v90d42a = BtoS_ACK8_p & v90fe87 | !BtoS_ACK8_p & v90e62f;
assign v93ef76 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v904115;
assign v86345d = BtoS_ACK7_p & v93fc04 | !BtoS_ACK7_p & v89b107;
assign v905038 = jx0_p & v863a78 | !jx0_p & v9074ce;
assign v8a8fed = jx0_p & v93f70c | !jx0_p & v844f91;
assign v93fe6e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9105ed;
assign v910d5a = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & !v93fca7;
assign v93e819 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90515d;
assign v93f734 = BtoS_ACK8_p & v8b5f61 | !BtoS_ACK8_p & !v8bbc51;
assign v93f8a9 = jx3_p & v907c01 | !jx3_p & !v844f91;
assign v93fe5d = FULL_p & v910525 | !FULL_p & v90e361;
assign v93f6da = stateG12_p & v908325 | !stateG12_p & v93eaa6;
assign v9077f7 = ENQ_p & v910242 | !ENQ_p & v911498;
assign v93f2d9 = StoB_REQ7_p & v912fed | !StoB_REQ7_p & v913435;
assign v904d75 = jx0_p & v90f5b6 | !jx0_p & !v930109;
assign v93e948 = BtoS_ACK7_p & v93e47b | !BtoS_ACK7_p & v93e90d;
assign v93f698 = StoB_REQ9_p & v93fb5d | !StoB_REQ9_p & v91086f;
assign v93fd3a = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v863a37;
assign v904dfc = RtoB_ACK0_p & v93f9cb | !RtoB_ACK0_p & v93f6ff;
assign v859635 = jx0_p & v908e01 | !jx0_p & !v93e933;
assign v90998d = BtoS_ACK6_p & v871df8 | !BtoS_ACK6_p & v907d8b;
assign v88932d = jx0_p & v844f91 | !jx0_p & !v844f95;
assign v9097da = jx1_p & v844f91 | !jx1_p & v93f91d;
assign v8b98f1 = jx3_p & v90950c | !jx3_p & v9099a1;
assign v90e79a = jx2_p & v93fdbd | !jx2_p & v90932c;
assign v905de8 = StoB_REQ7_p & v90f0a8 | !StoB_REQ7_p & v93f779;
assign v93e549 = BtoS_ACK0_p & v90855a | !BtoS_ACK0_p & !v90df22;
assign v93f8bf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fdd4;
assign v93faef = BtoS_ACK8_p & v93fdd9 | !BtoS_ACK8_p & !v90a4bd;
assign v907a2f = BtoS_ACK7_p & v905ff9 | !BtoS_ACK7_p & v8b9c31;
assign v90f7a9 = RtoB_ACK0_p & v910525 | !RtoB_ACK0_p & v93fe5d;
assign v93e439 = BtoS_ACK6_p & v863a78 | !BtoS_ACK6_p & v93f881;
assign v8f22d0 = jx0_p & v90aeb7 | !jx0_p & !v909180;
assign v93f98c = BtoS_ACK7_p & v93e024 | !BtoS_ACK7_p & v903b9c;
assign v905ac3 = stateG7_1_p & v93faac | !stateG7_1_p & v90a5c0;
assign v905f25 = jx1_p & v8f3826 | !jx1_p & v93f12b;
assign v904603 = DEQ_p & v90acfe | !DEQ_p & v93f6fa;
assign v8ee172 = jx2_p & v93dee0 | !jx2_p & !v910403;
assign v93fc76 = RtoB_ACK0_p & v8b9b56 | !RtoB_ACK0_p & v90e958;
assign v905186 = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & v9088a3;
assign v9091b2 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fe41;
assign v93ec26 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fa81;
assign v905660 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v93fdf7;
assign v93f470 = StoB_REQ6_p & v90aeb7 | !StoB_REQ6_p & v90508f;
assign v904296 = BtoS_ACK0_p & v90deff | !BtoS_ACK0_p & v910d10;
assign v9130c9 = jx1_p & v9050a5 | !jx1_p & v844f91;
assign v93fb03 = jx0_p & v909df9 | !jx0_p & v90d6ca;
assign v9056ac = jx3_p & v844f91 | !jx3_p & v90866d;
assign v93f821 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v9120f4;
assign v90ec05 = jx1_p & v93f1cf | !jx1_p & v93e89f;
assign v93fb9a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9068c8;
assign v90ee83 = BtoS_ACK6_p & v909f04 | !BtoS_ACK6_p & v9058f3;
assign v904afe = BtoS_ACK7_p & v907fc6 | !BtoS_ACK7_p & !v86dc4b;
assign v910bb8 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v93ef1d;
assign v905460 = BtoS_ACK9_p & v93dbe9 | !BtoS_ACK9_p & v85acd3;
assign v87bae8 = jx0_p & v844f91 | !jx0_p & v90eef9;
assign v90603e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v93e602;
assign v904677 = jx3_p & v93f937 | !jx3_p & v93efb8;
assign v90a20d = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v93fcf0;
assign v93fd63 = BtoS_ACK7_p & v863b25 | !BtoS_ACK7_p & v93f085;
assign v90fc5f = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v910642;
assign v90711a = StoB_REQ9_p & v903c0d | !StoB_REQ9_p & v910289;
assign v9092a8 = EMPTY_p & v8b49bf | !EMPTY_p & v93e72a;
assign v93f695 = stateG7_1_p & v88b26d | !stateG7_1_p & v905486;
assign v93fae4 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v91086d;
assign v93f16d = jx1_p & v910e82 | !jx1_p & !v911008;
assign v93fc04 = jx2_p & v844f91 | !jx2_p & v911c6f;
assign v93f56e = ENQ_p & v90a774 | !ENQ_p & !v844f91;
assign v87c534 = StoB_REQ9_p & v90468d | !StoB_REQ9_p & v907c71;
assign v9101d0 = jx3_p & v8a921d | !jx3_p & v90adc4;
assign v93f986 = jx1_p & v93fc94 | !jx1_p & !v844f91;
assign v91325d = StoB_REQ2_p & v93fd09 | !StoB_REQ2_p & v93e188;
assign v93f760 = jx2_p & v93fbeb | !jx2_p & v93fb73;
assign v9057cb = BtoS_ACK6_p & v93e8f6 | !BtoS_ACK6_p & v844fa1;
assign v911ebf = BtoS_ACK8_p & v906046 | !BtoS_ACK8_p & v87a1d0;
assign v90653d = jx2_p & v912378 | !jx2_p & v93eaf0;
assign v93e519 = BtoS_ACK9_p & v8b5f61 | !BtoS_ACK9_p & v93fa15;
assign v913a64 = BtoS_ACK8_p & v909a21 | !BtoS_ACK8_p & v903c1f;
assign v905329 = jx1_p & v910c37 | !jx1_p & !v93ef13;
assign v90e19c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90657d;
assign v85f243 = jx1_p & v9086b7 | !jx1_p & v9099e8;
assign v93f8c1 = jx2_p & v93f2a8 | !jx2_p & !v90a149;
assign v9076a7 = BtoS_ACK6_p & v93f9af | !BtoS_ACK6_p & v9045f4;
assign v90e373 = BtoS_ACK8_p & v93ec47 | !BtoS_ACK8_p & v93fc67;
assign v93eaf0 = jx1_p & v9050a5 | !jx1_p & v907069;
assign v90a33b = BtoS_ACK6_p & v91132f | !BtoS_ACK6_p & v93fe52;
assign v872746 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v907048;
assign v90a1fd = BtoS_ACK6_p & v863a78 | !BtoS_ACK6_p & v844f91;
assign v903fee = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & v90611f;
assign v90e1dd = jx0_p & v90d6e8 | !jx0_p & !v93f685;
assign v913662 = BtoS_ACK6_p & v910230 | !BtoS_ACK6_p & v844f91;
assign v876439 = StoB_REQ1_p & v93f85e | !StoB_REQ1_p & v90da97;
assign v93e682 = jx3_p & v93fbcc | !jx3_p & v911826;
assign v93f037 = StoB_REQ7_p & v87f17d | !StoB_REQ7_p & v844f91;
assign v93f59b = jx3_p & v93fad4 | !jx3_p & v90fbad;
assign v90a2b8 = BtoS_ACK6_p & v905537 | !BtoS_ACK6_p & v8b9d49;
assign v93f7fd = jx1_p & v9082ba | !jx1_p & v9114c0;
assign v93f5b9 = BtoS_ACK7_p & v907fc6 | !BtoS_ACK7_p & !v93fa84;
assign v90fb00 = DEQ_p & v906d83 | !DEQ_p & v93ea7f;
assign v9104aa = jx1_p & v911edb | !jx1_p & v90d87f;
assign v867045 = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & v908867;
assign v904a70 = jx3_p & v93f110 | !jx3_p & v9059b8;
assign v93fc6f = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v90add6;
assign v93fb2e = BtoS_ACK1_p & v906255 | !BtoS_ACK1_p & !v9120f4;
assign v906461 = BtoS_ACK6_p & v93f1cf | !BtoS_ACK6_p & v905d73;
assign v911937 = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & !v90f9b6;
assign v93fa91 = jx1_p & v93f0a9 | !jx1_p & v844f91;
assign v911f1f = BtoS_ACK6_p & v93fc0a | !BtoS_ACK6_p & v906623;
assign v93fe1e = BtoS_ACK0_p & v9046a6 | !BtoS_ACK0_p & v90a451;
assign v871df8 = jx0_p & v844f9f | !jx0_p & v844f91;
assign v93fd1a = StoB_REQ7_p & v910f4e | !StoB_REQ7_p & v844f91;
assign v904a80 = jx2_p & v9057c9 | !jx2_p & v908d10;
assign v89e06e = BtoS_ACK9_p & v90ea51 | !BtoS_ACK9_p & v904013;
assign v910e44 = ENQ_p & v90adc4 | !ENQ_p & v90ff7e;
assign v8b7122 = EMPTY_p & v906d92 | !EMPTY_p & v909eb5;
assign v90fa18 = jx1_p & v93f085 | !jx1_p & v909c45;
assign v904632 = RtoB_ACK0_p & v904d81 | !RtoB_ACK0_p & v9051ba;
assign v90e95b = jx0_p & v9057fa | !jx0_p & !v844f91;
assign v93e3a1 = StoB_REQ8_p & v93fc04 | !StoB_REQ8_p & v93fe3f;
assign v91150c = jx0_p & v93fb6c | !jx0_p & !v904736;
assign v906fec = jx0_p & v93f793 | !jx0_p & !v93f6f0;
assign v93f9a4 = BtoS_ACK6_p & v9058f3 | !BtoS_ACK6_p & v93f681;
assign v93e853 = ENQ_p & v911a33 | !ENQ_p & v9049b2;
assign v904ef2 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v93e369;
assign v93fad7 = jx0_p & v90d4ff | !jx0_p & !v93fc06;
assign v907abc = stateG12_p & v911a33 | !stateG12_p & v93fa29;
assign v90ede1 = jx0_p & v844f97 | !jx0_p & v844f91;
assign v87a20d = BtoS_ACK6_p & v90479e | !BtoS_ACK6_p & v9300da;
assign v9099e1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fce5;
assign v90db6b = jx1_p & v8a8b0a | !jx1_p & v912679;
assign v93fa27 = BtoS_ACK9_p & v90aa42 | !BtoS_ACK9_p & v906ac6;
assign v93fbd8 = jx1_p & v913332 | !jx1_p & v909080;
assign v8b4a3a = BtoR_REQ1_p & v93fe72 | !BtoR_REQ1_p & v8660c5;
assign v90a4da = jx2_p & v88dbe7 | !jx2_p & v908d10;
assign v90d880 = jx0_p & v8b49ad | !jx0_p & v90515d;
assign v9115ae = ENQ_p & v904f0d | !ENQ_p & v906c0f;
assign v90620e = BtoS_ACK8_p & v908237 | !BtoS_ACK8_p & !v93f06e;
assign v904e2f = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v903d0c;
assign v90d651 = RtoB_ACK0_p & v909bff | !RtoB_ACK0_p & v93fbdc;
assign v93fded = BtoS_ACK8_p & v93fc5d | !BtoS_ACK8_p & v930106;
assign v93fac5 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v867045;
assign v93faec = jx0_p & v93fc65 | !jx0_p & v90815c;
assign v9049bf = jx1_p & v93f085 | !jx1_p & v844f91;
assign v90657d = BtoS_ACK1_p & v93e356 | !BtoS_ACK1_p & v85ea9a;
assign v93fddc = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v9041e4;
assign v9068ce = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v89f90b;
assign v8b9ee2 = jx2_p & v93e54b | !jx2_p & !v904755;
assign v93f098 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v90f5bd;
assign v93fce3 = StoB_REQ7_p & v908e8e | !StoB_REQ7_p & v844f91;
assign v90eaab = jx0_p & v90d6e8 | !jx0_p & v93f6fc;
assign v8d373a = jx3_p & v93fa7d | !jx3_p & !v89f830;
assign v93df06 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v93f824;
assign v905405 = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v8850b3;
assign v93fa4b = jx0_p & v90d364 | !jx0_p & v844f91;
assign v90a6f4 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8bb868;
assign v906fc1 = BtoS_ACK6_p & v8a9289 | !BtoS_ACK6_p & v90d054;
assign v91063d = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a8fda;
assign v9088ff = jx0_p & v90cc30 | !jx0_p & !v90eef9;
assign v93f41e = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v93ec83;
assign v93fc0a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v90855a;
assign v93dee2 = BtoS_ACK0_p & v9051c9 | !BtoS_ACK0_p & !v93f6c3;
assign v90fbad = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v905847;
assign v93fada = StoB_REQ7_p & v93f9c6 | !StoB_REQ7_p & v9090dd;
assign v90dcf0 = jx2_p & v910260 | !jx2_p & v844f91;
assign v90ee63 = StoB_REQ2_p & v93f6de | !StoB_REQ2_p & v87c4d9;
assign v908436 = BtoS_ACK8_p & v844fa3 | !BtoS_ACK8_p & !v907e73;
assign v904258 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910f1b;
assign v904614 = DEQ_p & v93f7ae | !DEQ_p & v906fcc;
assign v89f803 = StoB_REQ6_p & v9070e3 | !StoB_REQ6_p & v93dee2;
assign v90ad0b = BtoS_ACK9_p & v93f7d7 | !BtoS_ACK9_p & v93fb69;
assign v90fb89 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v9050d2;
assign v9115b6 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93f462;
assign v910c4e = BtoS_ACK7_p & v93fb38 | !BtoS_ACK7_p & v910dda;
assign v87a203 = FULL_p & v844f91 | !FULL_p & v93f91c;
assign v90f52f = StoB_REQ6_p & v90a0e8 | !StoB_REQ6_p & v9111cf;
assign v91071b = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93fccc;
assign v93e0c5 = StoB_REQ6_p & v912383 | !StoB_REQ6_p & v8b9e3d;
assign v93fb91 = BtoS_ACK9_p & v93e048 | !BtoS_ACK9_p & v908edf;
assign v90419d = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v90a0d7;
assign v9058e9 = StoB_REQ2_p & v93fd09 | !StoB_REQ2_p & v904d08;
assign v90d5bd = BtoS_ACK6_p & v8b9d27 | !BtoS_ACK6_p & v87f17d;
assign v90809b = jx2_p & v9049fd | !jx2_p & v906dd6;
assign v93fb83 = StoB_REQ0_p & v93f7f5 | !StoB_REQ0_p & v93f155;
assign v906534 = jx1_p & v93fdf0 | !jx1_p & v9043f4;
assign v93fe27 = BtoS_ACK6_p & v863a78 | !BtoS_ACK6_p & v904775;
assign v904221 = jx1_p & v85eacb | !jx1_p & v93f811;
assign v907e91 = jx2_p & v93f9f4 | !jx2_p & v90d22a;
assign v904b63 = StoB_REQ1_p & v90534f | !StoB_REQ1_p & v844f91;
assign v9044b1 = jx0_p & v9054b5 | !jx0_p & !v93f6fc;
assign v908e8b = BtoS_ACK8_p & v93fb78 | !BtoS_ACK8_p & v93fc7b;
assign v908e75 = BtoS_ACK7_p & v9114c9 | !BtoS_ACK7_p & !v90edca;
assign v9051ea = StoB_REQ7_p & v8b714e | !StoB_REQ7_p & v90894d;
assign v90df22 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b9c3f;
assign v90d877 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v908df7;
assign v93f0a7 = ENQ_p & v90adc4 | !ENQ_p & v93e440;
assign v87a2ae = BtoR_REQ1_p & v8f383a | !BtoR_REQ1_p & v910704;
assign v90cc57 = jx2_p & v8a8f6f | !jx2_p & v87f17d;
assign v91359a = ENQ_p & v8f2274 | !ENQ_p & v93fc97;
assign v93fd73 = jx3_p & v93fa7d | !jx3_p & !v93f82d;
assign v93f88d = StoB_REQ8_p & v907469 | !StoB_REQ8_p & v8b9884;
assign v904fd6 = DEQ_p & v913399 | !DEQ_p & v904fee;
assign v90cfda = jx1_p & v93f727 | !jx1_p & v906c66;
assign v90acfe = RtoB_ACK0_p & v93f7d6 | !RtoB_ACK0_p & v93f6fa;
assign v89f930 = jx0_p & v93ebd1 | !jx0_p & v907a13;
assign v90d00f = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v93fe04;
assign v90817e = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & v909ecc;
assign v90e341 = StoB_REQ7_p & v90998d | !StoB_REQ7_p & v90a33b;
assign v911498 = jx3_p & v844f91 | !jx3_p & v93e8cc;
assign v910d81 = jx2_p & v887bb8 | !jx2_p & v90932c;
assign v9049b2 = jx3_p & v93e137 | !jx3_p & !v908ae5;
assign v93f824 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v93fe36;
assign v93e9de = StoB_REQ7_p & v9102f4 | !StoB_REQ7_p & v93fc8d;
assign v87c9bf = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v90811c;
assign v93ee87 = jx0_p & v90d879 | !jx0_p & v844f91;
assign v90e028 = jx2_p & v93fda5 | !jx2_p & !v93fdc8;
assign v93fc84 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v908068;
assign v905a88 = StoB_REQ9_p & v90e159 | !StoB_REQ9_p & v93f9a7;
assign v912378 = jx1_p & v87c54e | !jx1_p & v906dea;
assign v93fd2e = BtoS_ACK9_p & v904c52 | !BtoS_ACK9_p & v9063b2;
assign v9040fb = jx2_p & v904c99 | !jx2_p & v844f91;
assign v907fc6 = jx2_p & v912f4e | !jx2_p & v910243;
assign v90ee4b = BtoS_ACK8_p & v93fbe4 | !BtoS_ACK8_p & v93ec28;
assign v90a2c8 = StoB_REQ1_p & v908df7 | !StoB_REQ1_p & v844f91;
assign v93e385 = jx1_p & v9090d1 | !jx1_p & v93f82e;
assign v906034 = DEQ_p & v913399 | !DEQ_p & v90f0c5;
assign v93f76b = StoB_REQ7_p & v90ec5d | !StoB_REQ7_p & v8d1873;
assign v912687 = StoB_REQ7_p & v904e70 | !StoB_REQ7_p & v910243;
assign v93e751 = EMPTY_p & v93e262 | !EMPTY_p & v90e9a1;
assign v9097c3 = jx1_p & v9093ec | !jx1_p & v9122e7;
assign v92ffd3 = jx3_p & v904590 | !jx3_p & !v87f17d;
assign v93f6c3 = StoB_REQ0_p & v906642 | !StoB_REQ0_p & v9083d3;
assign v9111a4 = StoB_REQ8_p & v907469 | !StoB_REQ8_p & v93f972;
assign v9082e4 = BtoS_ACK0_p & v86c2d0 | !BtoS_ACK0_p & v93fe20;
assign v904025 = jx3_p & v93f927 | !jx3_p & !v9097db;
assign v93f345 = BtoS_ACK6_p & v904aae | !BtoS_ACK6_p & v8a927b;
assign v93f30c = jx1_p & v93f7b0 | !jx1_p & !v89f916;
assign v8a1fe3 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v9093a9;
assign v912cf4 = jx2_p & v93fa16 | !jx2_p & !v93f860;
assign v907bfd = StoB_REQ8_p & v93e27a | !StoB_REQ8_p & v904bc1;
assign v93f6bf = jx1_p & v90f07f | !jx1_p & !v844f91;
assign v905d92 = ENQ_p & v93fa2b | !ENQ_p & v93e70e;
assign v913225 = EMPTY_p & v93f695 | !EMPTY_p & v91335a;
assign v93f856 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v93fa54;
assign v8b9bd9 = jx1_p & v8b9dff | !jx1_p & v93fdf8;
assign v907f0e = jx1_p & v90a002 | !jx1_p & !v93fb1d;
assign v905199 = jx2_p & v93f39f | !jx2_p & v90606c;
assign v8b9e12 = BtoS_ACK0_p & v9047b7 | !BtoS_ACK0_p & v90603e;
assign v909fb2 = jx2_p & v905d36 | !jx2_p & !v90ec84;
assign v903bb1 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v908346;
assign v905b62 = BtoS_ACK7_p & v911f15 | !BtoS_ACK7_p & v93f6c9;
assign v93e69c = DEQ_p & v909d90 | !DEQ_p & v906fcc;
assign v91086f = BtoS_ACK8_p & v93fde5 | !BtoS_ACK8_p & v912190;
assign v8d3791 = StoB_REQ8_p & v87a1d0 | !StoB_REQ8_p & v91229f;
assign v93ea28 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v90f36b;
assign v90749b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93e773;
assign v908106 = BtoS_ACK8_p & v93f66b | !BtoS_ACK8_p & !v904fd2;
assign v91026f = BtoS_ACK6_p & v93e89f | !BtoS_ACK6_p & v87f17d;
assign v93f91c = ENQ_p & v844f91 | !ENQ_p & v910e55;
assign v9052f0 = BtoS_ACK7_p & v93fdd2 | !BtoS_ACK7_p & v908e92;
assign v9054a8 = jx3_p & v8b9e71 | !jx3_p & v90eea6;
assign v907ccf = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8ee1a9;
assign v8a9231 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90521f;
assign v91a771 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v904b04 = jx2_p & v93f533 | !jx2_p & v90966d;
assign v8b9e6e = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v863aa0;
assign v906f1e = jx1_p & v93f8d0 | !jx1_p & v844f91;
assign v9091fe = StoB_REQ7_p & v90d22b | !StoB_REQ7_p & v905194;
assign v903e2f = ENQ_p & v93fda6 | !ENQ_p & v905da0;
assign v90faf6 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v903fc8;
assign v93fcdb = BtoS_ACK6_p & v93fcbe | !BtoS_ACK6_p & v90f2ff;
assign v93f766 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a6d8;
assign v910bd7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v906642;
assign v93fb53 = jx1_p & v90a620 | !jx1_p & !v903e94;
assign v93ee3b = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v844f91;
assign v905d36 = jx1_p & v9047cd | !jx1_p & v93f826;
assign v905972 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844fb5;
assign v89b0e5 = jx3_p & v913433 | !jx3_p & v907d8a;
assign v93fa04 = jx0_p & v844f91 | !jx0_p & v93fa6d;
assign v91038c = jx1_p & v93e819 | !jx1_p & v906dea;
assign v93f840 = StoB_REQ2_p & v93fcf0 | !StoB_REQ2_p & v93f27f;
assign v906d38 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90fcbf;
assign v90ed41 = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v93ea50;
assign v93f111 = jx0_p & v93fc0a | !jx0_p & v904725;
assign v90df4b = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v904432;
assign v8b49f1 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v909082;
assign v863a7b = ENQ_p & v93f89f | !ENQ_p & v90ec4b;
assign v905434 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v93f6ce;
assign v93faf9 = jx2_p & v904008 | !jx2_p & v863afc;
assign v93fe56 = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v8857fd;
assign v93fd85 = ENQ_p & v9083cf | !ENQ_p & v93fe38;
assign v90dc09 = StoB_REQ9_p & v93fd96 | !StoB_REQ9_p & v93fced;
assign v93f9af = jx0_p & v93fc0a | !jx0_p & v93f119;
assign v906c3f = StoB_REQ8_p & v90ddf9 | !StoB_REQ8_p & v904afe;
assign v910ffd = RtoB_ACK0_p & v93df9f | !RtoB_ACK0_p & v905d92;
assign v86344b = jx0_p & v844f9b | !jx0_p & !v844f99;
assign v906c91 = BtoS_ACK7_p & v906b57 | !BtoS_ACK7_p & v90ecba;
assign v93db10 = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v908a98;
assign v93fbee = jx3_p & v844f91 | !jx3_p & v910416;
assign v91216e = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v90636e;
assign v93e5f1 = jx3_p & v91aa04 | !jx3_p & !v93fe54;
assign v93f7b4 = BtoS_ACK7_p & v93f7f8 | !BtoS_ACK7_p & v93fa82;
assign v93f6fa = ENQ_p & v844f91 | !ENQ_p & v93fad5;
assign v90d6ca = StoB_REQ6_p & v88b9b7 | !StoB_REQ6_p & v844f91;
assign v90999b = StoB_REQ6_p & v90569e | !StoB_REQ6_p & v844f91;
assign v93db3f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v909078;
assign v904141 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v87ca8a;
assign v93e126 = jx0_p & v90ef1b | !jx0_p & v844f99;
assign v93e731 = RtoB_ACK0_p & v90809e | !RtoB_ACK0_p & v90aaa8;
assign v90a799 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v910f78;
assign v906c20 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8ee1bc;
assign v93f28b = BtoS_ACK6_p & v90a216 | !BtoS_ACK6_p & v910cda;
assign v93e68f = jx1_p & v906461 | !jx1_p & v904f32;
assign v93ea7f = RtoB_ACK0_p & v93f19b | !RtoB_ACK0_p & v9082be;
assign v87c517 = DEQ_p & v8b9d0e | !DEQ_p & v90dcca;
assign v87c525 = BtoS_ACK7_p & v93fc04 | !BtoS_ACK7_p & v905810;
assign v90612e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844fbd;
assign v9100bd = jx2_p & v93fd6d | !jx2_p & v90cb3d;
assign v9042ba = jx1_p & v89e11b | !jx1_p & v90a4f9;
assign v907bd4 = ENQ_p & v908325 | !ENQ_p & v9135f1;
assign v93fb7b = jx1_p & v844f91 | !jx1_p & v90a786;
assign v908f85 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v903d0b;
assign v8b9c4f = ENQ_p & v93f893 | !ENQ_p & v90444f;
assign v905841 = BtoS_ACK6_p & v9088ff | !BtoS_ACK6_p & !v93dac8;
assign v93f7a2 = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v91325d;
assign v904f1b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93ec0d;
assign v910260 = jx1_p & v844f91 | !jx1_p & !v906320;
assign v9067d4 = StoB_REQ9_p & v87f17f | !StoB_REQ9_p & !v90ad0a;
assign v93f87a = jx1_p & v911edb | !jx1_p & v90f3e4;
assign v93e296 = BtoS_ACK7_p & v93fc04 | !BtoS_ACK7_p & v91a992;
assign v908e92 = jx2_p & v87c51f | !jx2_p & !v863b2f;
assign BtoR_REQ1_n = !v8a9267;
assign v89f852 = jx0_p & v844f91 | !jx0_p & !v93ef46;
assign v90f0aa = StoB_REQ8_p & v90dab9 | !StoB_REQ8_p & v911167;
assign v904a61 = BtoS_ACK6_p & v91aa51 | !BtoS_ACK6_p & v844f91;
assign v91218a = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v90d7e7;
assign v93f1c8 = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & !v904f52;
assign v89f988 = StoB_REQ8_p & v9110ab | !StoB_REQ8_p & v9059d6;
assign v903db4 = StoB_REQ9_p & v93f801 | !StoB_REQ9_p & v85ef3a;
assign v907679 = jx2_p & v93f39f | !jx2_p & v93faa8;
assign v93fd84 = jx1_p & v90459f | !jx1_p & !v844f91;
assign v903fc8 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v90ea47;
assign v93fa44 = jx1_p & v90e6f1 | !jx1_p & v91879a;
assign v8b9f3e = BtoS_ACK1_p & v93dffe | !BtoS_ACK1_p & v909c0e;
assign v91a9b4 = BtoS_ACK0_p & v93e391 | !BtoS_ACK0_p & v9134fe;
assign v93f334 = BtoS_ACK9_p & v9050cc | !BtoS_ACK9_p & v93ebbb;
assign BtoS_ACK2_n = !v91aa7d;
assign v90759b = StoB_REQ1_p & v90e945 | !StoB_REQ1_p & v90d1ca;
assign v93f88a = StoB_REQ7_p & v90d22b | !StoB_REQ7_p & v90805e;
assign v907494 = RtoB_ACK0_p & v90dd67 | !RtoB_ACK0_p & v89e0d5;
assign v9134df = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93e2de;
assign v87e087 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93f69c;
assign v93fd4c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b9c3e;
assign v90aa76 = jx0_p & v93fa3c | !jx0_p & !v844f91;
assign v93dfe2 = StoB_REQ6_p & v93f32a | !StoB_REQ6_p & v85ea7f;
assign v93e335 = jx1_p & v903fef | !jx1_p & v844f91;
assign v863aa0 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v90ad69;
assign v93f058 = BtoS_ACK6_p & v863a78 | !BtoS_ACK6_p & v912405;
assign v904cc8 = stateG7_1_p & v844f91 | !stateG7_1_p & v908e7f;
assign v93f2fd = ENQ_p & v93f89f | !ENQ_p & v904bda;
assign v90ea74 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v93db4a;
assign v907e6b = jx0_p & v93fc65 | !jx0_p & v93f8d1;
assign v90cf52 = jx2_p & v90927b | !jx2_p & v93faf8;
assign v93fce6 = StoB_REQ9_p & v93f3b9 | !StoB_REQ9_p & v93fbfa;
assign v91003a = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & !v90d1ca;
assign v910f4d = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93e156;
assign v93ed29 = BtoS_ACK7_p & v910e66 | !BtoS_ACK7_p & v90f7d1;
assign v93eec4 = StoB_REQ2_p & v93ed70 | !StoB_REQ2_p & v90eef5;
assign v91090e = EMPTY_p & v93f6f9 | !EMPTY_p & !v8b9cc5;
assign v93ee22 = BtoS_ACK6_p & v90db9f | !BtoS_ACK6_p & v93fbe6;
assign v9126bb = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90748b;
assign v86335a = BtoS_ACK1_p & v93fccb | !BtoS_ACK1_p & v9104e0;
assign v91006b = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v907206;
assign v90f629 = ENQ_p & v90adc4 | !ENQ_p & v8b9972;
assign v909001 = DEQ_p & v9041a7 | !DEQ_p & v92ffd3;
assign v93efbb = jx0_p & v90ed41 | !jx0_p & v93fa90;
assign v93fb45 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v908f29;
assign v93fe57 = StoB_REQ8_p & v93ea16 | !StoB_REQ8_p & v8f223b;
assign v908fb8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93e371;
assign v90e2d7 = BtoS_ACK7_p & v90d3ff | !BtoS_ACK7_p & v90dcb3;
assign v91a796 = stateG12_p & v93f15e | !stateG12_p & v90faf6;
assign v93fa85 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v904d1a;
assign v91a9cd = StoB_REQ1_p & v90fc92 | !StoB_REQ1_p & v844f91;
assign v9049ac = ENQ_p & v90adc4 | !ENQ_p & v9135e7;
assign v93e86c = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v89f7e7;
assign v91268a = jx0_p & v93f8ca | !jx0_p & v93f8ab;
assign v909a08 = BtoR_REQ0_p & v904b1b | !BtoR_REQ0_p & v903cd1;
assign v85cca5 = StoB_REQ9_p & v86d7d1 | !StoB_REQ9_p & v93ece6;
assign v90aa8a = jx0_p & v8a927b | !jx0_p & v90515d;
assign v90aa3c = BtoS_ACK8_p & v9132eb | !BtoS_ACK8_p & !v89fd94;
assign v93fa7d = BtoS_ACK9_p & v93fd95 | !BtoS_ACK9_p & v906df1;
assign v90dedf = stateG7_1_p & v90f0bd | !stateG7_1_p & v904dc1;
assign v85eb14 = EMPTY_p & v844fcd | !EMPTY_p & !v844fcf;
assign v906b5f = jx2_p & v905618 | !jx2_p & !v91a76f;
assign v93e72a = DEQ_p & v93df9f | !DEQ_p & v93dfb4;
assign v908fba = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v90e611;
assign v93fe48 = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & !v904ba7;
assign v8f60f9 = jx1_p & v93f90a | !jx1_p & v912679;
assign v910937 = StoB_REQ9_p & v90e9f7 | !StoB_REQ9_p & v93fa93;
assign v93f7d9 = jx2_p & v904234 | !jx2_p & v844f91;
assign v905824 = BtoS_ACK0_p & v93e2de | !BtoS_ACK0_p & v93facb;
assign v87f17d = jx0_p & v844f91 | !jx0_p & !v844f91;
assign v905170 = EMPTY_p & v9061b3 | !EMPTY_p & v904603;
assign v844fa5 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v844f91;
assign v93ed70 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v90f547;
assign v90a23c = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v912fc9;
assign v93f31f = StoB_REQ7_p & v904e70 | !StoB_REQ7_p & v844f91;
assign v911318 = jx0_p & v93fdb6 | !jx0_p & v911312;
assign v90e5b9 = DEQ_p & v93fa36 | !DEQ_p & v90dc2c;
assign v93fa52 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v93e800;
assign v91364c = BtoS_ACK8_p & v93ed2a | !BtoS_ACK8_p & v93f8fa;
assign v905f24 = BtoS_ACK9_p & v90736f | !BtoS_ACK9_p & v90e988;
assign v9072b7 = stateG12_p & v93eed6 | !stateG12_p & v90f391;
assign v93f892 = jx3_p & v93fa7d | !jx3_p & !v90cbea;
assign v93faf2 = jx2_p & v93fda8 | !jx2_p & v907e86;
assign v91a757 = jx1_p & v93fd77 | !jx1_p & v9043f4;
assign v85eb28 = jx3_p & v844f91 | !jx3_p & v91066d;
assign v90985e = StoB_REQ7_p & v93fe33 | !StoB_REQ7_p & v9047f0;
assign v9051bb = StoB_REQ7_p & v9093ec | !StoB_REQ7_p & !v93f111;
assign v90470d = StoB_REQ9_p & v93f827 | !StoB_REQ9_p & v93fad2;
assign v844fb9 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f91;
assign v8b9960 = RtoB_ACK0_p & v86e277 | !RtoB_ACK0_p & v909878;
assign v903c2a = BtoS_ACK7_p & v93ed2a | !BtoS_ACK7_p & v904d89;
assign v93fc24 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v93f827;
assign v90a5a4 = DEQ_p & v93f7d6 | !DEQ_p & v863a97;
assign v863a3f = ENQ_p & v93eda4 | !ENQ_p & v907417;
assign v909e7f = StoB_REQ1_p & v906642 | !StoB_REQ1_p & v93f6a7;
assign v93f6e9 = jx2_p & v908cf4 | !jx2_p & v880314;
assign v904e47 = jx0_p & v908a2f | !jx0_p & !v93f8e4;
assign v907b84 = jx3_p & v93e105 | !jx3_p & !v93fe73;
assign v93fd93 = BtoS_ACK7_p & v93f6bd | !BtoS_ACK7_p & v93f68f;
assign v9111cf = BtoS_ACK0_p & v90534f | !BtoS_ACK0_p & v93fac2;
assign v904f5e = StoB_REQ8_p & v85ea93 | !StoB_REQ8_p & v844f91;
assign v905764 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844fa1;
assign v8a8f89 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93fe48;
assign v863b34 = StoB_REQ8_p & v91042d | !StoB_REQ8_p & v90683e;
assign v907c76 = BtoS_ACK8_p & v93f73d | !BtoS_ACK8_p & v913428;
assign v93fb1d = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & v913a60;
assign v90ba31 = BtoS_ACK9_p & v93fa54 | !BtoS_ACK9_p & !v90ef1a;
assign v911008 = StoB_REQ7_p & v866af4 | !StoB_REQ7_p & v93fabb;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v93f518 = jx1_p & v8b9eca | !jx1_p & !v907e7a;
assign v93fc68 = jx0_p & v844f91 | !jx0_p & v844fa1;
assign v93fb48 = StoB_REQ1_p & v93fc8e | !StoB_REQ1_p & !v90a233;
assign v89f97f = jx2_p & v93fa25 | !jx2_p & v90f1ab;
assign v908e52 = jx0_p & v93e589 | !jx0_p & v93e9d1;
assign v90a18c = EMPTY_p & v910c0f | !EMPTY_p & v904cc8;
assign v93fe04 = jx0_p & v907d33 | !jx0_p & v93fa40;
assign v91a76f = jx1_p & v93f31f | !jx1_p & v93fa4c;
assign v93f682 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v9054b5;
assign v87f17f = jx1_p & v844f91 | !jx1_p & !v844f91;
assign v93fca2 = BtoS_ACK6_p & v91aa51 | !BtoS_ACK6_p & v880d7e;
assign v910d62 = EMPTY_p & v93eb1d | !EMPTY_p & v91db5b;
assign v8633df = DEQ_p & v91a6e9 | !DEQ_p & v90ea21;
assign v90d543 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v903ec3;
assign v903c40 = StoB_REQ9_p & v90e9f7 | !StoB_REQ9_p & v90419d;
assign v90f1cb = BtoS_ACK6_p & v93fcc9 | !BtoS_ACK6_p & v87f17d;
assign v90d629 = jx3_p & v844f91 | !jx3_p & v903bfc;
assign v93f727 = StoB_REQ7_p & v9093ec | !StoB_REQ7_p & !v93f119;
assign v87ca3a = BtoR_REQ0_p & v91214b | !BtoR_REQ0_p & v93f9d7;
assign v93e77c = jx1_p & v93f8d0 | !jx1_p & v9046de;
assign v90a1db = jx2_p & v93f535 | !jx2_p & v9097c6;
assign v90cc4a = BtoS_ACK9_p & v93fc04 | !BtoS_ACK9_p & v90dd77;
assign v871033 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910825;
assign v911c50 = StoB_REQ1_p & v90e251 | !StoB_REQ1_p & v90ea8a;
assign v907c01 = BtoS_ACK9_p & v8b497a | !BtoS_ACK9_p & v9067d4;
assign v8b9884 = BtoS_ACK7_p & v8b9ee2 | !BtoS_ACK7_p & v93fd8c;
assign v93fd2f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9046d6;
assign v9124c5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9096fd;
assign v904b91 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v90d789;
assign v911452 = StoB_REQ9_p & v903c0d | !StoB_REQ9_p & v9063d8;
assign v913342 = BtoS_ACK7_p & v93f8c1 | !BtoS_ACK7_p & !v911815;
assign v8c8823 = BtoR_REQ1_p & v93fe1a | !BtoR_REQ1_p & !v909546;
assign v904b8c = ENQ_p & v93f15e | !ENQ_p & v910237;
assign v90e94e = jx1_p & v869aeb | !jx1_p & !v871df8;
assign v910fd8 = StoB_REQ7_p & v90998d | !StoB_REQ7_p & v90648f;
assign v93fb08 = jx0_p & v90f2ff | !jx0_p & v93fcbe;
assign v93f813 = BtoS_ACK7_p & v906c2f | !BtoS_ACK7_p & v909b10;
assign v93fdd5 = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & !v910383;
assign v9081aa = BtoS_ACK9_p & v93e048 | !BtoS_ACK9_p & v9119f8;
assign v8ee1c7 = jx0_p & v90aeb7 | !jx0_p & v90690e;
assign v906c67 = jx1_p & v844f91 | !jx1_p & !v871df8;
assign v904df8 = StoB_REQ1_p & v904ae0 | !StoB_REQ1_p & v90479a;
assign v93f6ae = RtoB_ACK0_p & v90ad6f | !RtoB_ACK0_p & v90e437;
assign v873a26 = EMPTY_p & v93fdbe | !EMPTY_p & v93f9ff;
assign v909365 = StoB_REQ9_p & v8d37d4 | !StoB_REQ9_p & v93e6c2;
assign v870d72 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v907c59;
assign v93ea3e = jx1_p & v90f5ff | !jx1_p & v90515a;
assign v87c4e7 = jx2_p & v90d634 | !jx2_p & v905dc1;
assign v90eab9 = StoB_REQ9_p & v91109f | !StoB_REQ9_p & v918724;
assign v93fd06 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v89f881;
assign v904da6 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v909367;
assign v86313d = jx0_p & v90ed41 | !jx0_p & v90a9e4;
assign v869aeb = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v87f17d;
assign v910db7 = StoB_REQ8_p & v93f444 | !StoB_REQ8_p & v90d704;
assign v906037 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v93fdd7;
assign v93fcbc = jx2_p & v904a0b | !jx2_p & v93e919;
assign v87a1d0 = BtoS_ACK7_p & v906046 | !BtoS_ACK7_p & v90da41;
assign v93f74a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v909691;
assign v8f3825 = StoB_REQ8_p & v93fdd9 | !StoB_REQ8_p & v9132eb;
assign v89f8bc = jx1_p & v844f91 | !jx1_p & !v90d7a0;
assign v9064e9 = stateG12_p & v844f91 | !stateG12_p & v93f0a6;
assign v913428 = BtoS_ACK7_p & v910fda | !BtoS_ACK7_p & v90808b;
assign v904fbb = StoB_REQ9_p & v87f17f | !StoB_REQ9_p & v8b70a3;
assign v910d6d = StoB_REQ7_p & v908e8e | !StoB_REQ7_p & v870489;
assign v93fd8f = BtoS_ACK6_p & v90df7f | !BtoS_ACK6_p & v908e52;
assign v93fa2b = jx3_p & v90aeb8 | !jx3_p & v90fbad;
assign v9045f4 = jx0_p & v906623 | !jx0_p & v93f119;
assign v90dd77 = BtoS_ACK8_p & v93fc04 | !BtoS_ACK8_p & v93e296;
assign v93fbfa = BtoS_ACK8_p & v9095b9 | !BtoS_ACK8_p & v911b47;
assign v90ff7e = jx3_p & v93e7af | !jx3_p & v90851b;
assign v904ed4 = StoB_REQ6_p & v930028 | !StoB_REQ6_p & v93fac3;
assign v93f6ec = BtoS_ACK2_p & v906cc8 | !BtoS_ACK2_p & v9058e9;
assign v908ed6 = jx1_p & v844f91 | !jx1_p & !v90ede1;
assign v93fbf8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93ef30;
assign v905d9c = jx1_p & v903cf9 | !jx1_p & v844f91;
assign v90a774 = jx3_p & v93f7a1 | !jx3_p & v844fc3;
assign v909746 = StoB_REQ8_p & v904ab4 | !StoB_REQ8_p & v93fd52;
assign v9043c7 = jx2_p & v93ec4d | !jx2_p & v91a757;
assign v9077b1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ebd28;
assign v8f37f1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90557c;
assign v93fe0e = jx0_p & v93fa4f | !jx0_p & !v844f91;
assign v93faca = BtoS_ACK9_p & v8b5f61 | !BtoS_ACK9_p & v91053d;
assign v904c38 = StoB_REQ0_p & v85eabe | !StoB_REQ0_p & v844f91;
assign v91230c = jx2_p & v93e1c0 | !jx2_p & v90cb3d;
assign v85ea5f = BtoS_ACK1_p & v9046a6 | !BtoS_ACK1_p & !v90e945;
assign v93fda5 = jx1_p & v844f91 | !jx1_p & v90a4c6;
assign v8b9dcb = BtoS_ACK7_p & v910fda | !BtoS_ACK7_p & v905168;
assign v908322 = jx1_p & v87a21e | !jx1_p & v93fd2c;
assign v90eea7 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v905ed9;
assign v90ad3d = ENQ_p & v863add | !ENQ_p & !v93f8a9;
assign v8b4a08 = BtoS_ACK6_p & v904e70 | !BtoS_ACK6_p & v93fc40;
assign v93e097 = StoB_REQ8_p & v9134bc | !StoB_REQ8_p & v93e596;
assign v8b9e97 = FULL_p & v909dec | !FULL_p & v90dcca;
assign v907b60 = ENQ_p & v93fdf6 | !ENQ_p & v93facc;
assign v89b100 = BtoS_ACK6_p & v93fcc9 | !BtoS_ACK6_p & v903e62;
assign v910cda = jx0_p & v87a979 | !jx0_p & v90cbf7;
assign v9085f5 = DEQ_p & v88bb45 | !DEQ_p & v907301;
assign v89f8b8 = StoB_REQ8_p & v93e9d8 | !StoB_REQ8_p & v844f91;
assign v908553 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v912ec8;
assign v93fbcc = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v9050ba;
assign v93f9c5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b9f3e;
assign v93f91d = jx0_p & v93fa95 | !jx0_p & v906d53;
assign v905246 = BtoS_ACK9_p & v8633ec | !BtoS_ACK9_p & v903cef;
assign v90adc4 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v93f87b;
assign v910e72 = jx0_p & v86ccf1 | !jx0_p & v903df5;
assign v903b83 = BtoS_ACK9_p & v9073c5 | !BtoS_ACK9_p & v90f7e4;
assign v93e6c2 = BtoS_ACK8_p & v905e43 | !BtoS_ACK8_p & !v93fae2;
assign v8b9d5d = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v91150c;
assign v93f94a = jx0_p & v90ea74 | !jx0_p & !v90f52f;
assign v9051d8 = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v93f8bf;
assign v912672 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v87c533;
assign v863444 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v9300af;
assign v87c51e = RtoB_ACK0_p & v905697 | !RtoB_ACK0_p & v8b9cc5;
assign v93f75c = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v9059a0;
assign v910642 = StoB_REQ3_p & v93fd8e | !StoB_REQ3_p & v90f547;
assign v93f801 = BtoS_ACK8_p & v93f73d | !BtoS_ACK8_p & v93fe4b;
assign v906201 = BtoS_ACK6_p & v910f82 | !BtoS_ACK6_p & v90ad47;
assign v93f784 = jx3_p & v93f1ad | !jx3_p & !v90490e;
assign v911d61 = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & v93e14a;
assign v90738b = EMPTY_p & v905292 | !EMPTY_p & v910fcd;
assign v93f919 = RtoB_ACK0_p & v89e0d5 | !RtoB_ACK0_p & v9133ec;
assign v90ace9 = ENQ_p & v93f89f | !ENQ_p & v87c4ee;
assign v8b4a10 = StoB_REQ9_p & v90e8f5 | !StoB_REQ9_p & v93ecf7;
assign v909f4b = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & v930037;
assign v8633ec = StoB_REQ8_p & v93e115 | !StoB_REQ8_p & v844f91;
assign v90a4f9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9096f3;
assign v87cb9e = BtoS_ACK0_p & v911102 | !BtoS_ACK0_p & v93fb37;
assign v93ec07 = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v90f864;
assign v904ecc = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v93fc27;
assign v93fc18 = StoB_REQ8_p & v90e2d7 | !StoB_REQ8_p & v905b62;
assign v93fc02 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93dffe;
assign v93f782 = jx0_p & v93f854 | !jx0_p & v90f88a;
assign v906fba = StoB_REQ9_p & v907c76 | !StoB_REQ9_p & v93f822;
assign v903fef = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93e6af;
assign v93ef57 = jx0_p & v93f70b | !jx0_p & v93fd94;
assign v93fb33 = BtoS_ACK8_p & v9132dc | !BtoS_ACK8_p & !v906c3f;
assign v8b9cc5 = ENQ_p & v8b98f1 | !ENQ_p & v93fc93;
assign v93fdd9 = jx2_p & v9057c1 | !jx2_p & v90ded0;
assign v88a51e = ENQ_p & v93fa2b | !ENQ_p & v844f91;
assign v93fd16 = jx0_p & v9133f0 | !jx0_p & v93e0c5;
assign v912172 = DEQ_p & v8b9d0e | !DEQ_p & v93f70f;
assign v90d4ff = StoB_REQ6_p & v93f8a0 | !StoB_REQ6_p & v87cb9e;
assign v910b33 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93f79a;
assign v90f07f = BtoS_ACK6_p & v93f1cf | !BtoS_ACK6_p & v90d217;
assign v911fe3 = jx1_p & v8f22ad | !jx1_p & !v908af7;
assign v93e886 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v93eb43;
assign v93faed = BtoS_ACK8_p & v93f768 | !BtoS_ACK8_p & v907799;
assign v8b9e1d = ENQ_p & v912477 | !ENQ_p & v8b495a;
assign v903b9c = jx1_p & v93e819 | !jx1_p & v870d72;
assign v907a32 = ENQ_p & v844f91 | !ENQ_p & v86ce19;
assign v90966d = jx1_p & v911724 | !jx1_p & v9043f4;
assign v907d70 = StoB_REQ7_p & v93fdea | !StoB_REQ7_p & v93fb07;
assign v8b9dbd = BtoS_ACK6_p & v910243 | !BtoS_ACK6_p & v9083d0;
assign v93e8cc = BtoS_ACK9_p & v906046 | !BtoS_ACK9_p & v911ebf;
assign v909bd3 = jx3_p & v93f749 | !jx3_p & !v93da97;
assign v883cbe = BtoS_ACK8_p & v90722c | !BtoS_ACK8_p & !v93f9bc;
assign v9093f3 = BtoS_ACK8_p & v9095b9 | !BtoS_ACK8_p & v909746;
assign v93f69a = BtoS_ACK9_p & v905d97 | !BtoS_ACK9_p & v90664c;
assign v93fd14 = jx0_p & v85eaa5 | !jx0_p & v903e8d;
assign v93f204 = ENQ_p & v93fdf6 | !ENQ_p & v8b495a;
assign v9064b4 = StoB_REQ7_p & v9043f4 | !StoB_REQ7_p & v903d01;
assign v91aa76 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85eaed;
assign v93f80a = jx3_p & v908ad9 | !jx3_p & v93fb91;
assign v911b74 = jx3_p & v93fd59 | !jx3_p & !v93e519;
assign v907897 = BtoS_ACK6_p & v905038 | !BtoS_ACK6_p & v909415;
assign v905d97 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93f6a0;
assign v93fbf3 = jx1_p & v93f6fe | !jx1_p & v9045bb;
assign v90d4c9 = StoB_REQ9_p & v911cba | !StoB_REQ9_p & v89f7e3;
assign v93fd64 = StoB_REQ9_p & v90dd77 | !StoB_REQ9_p & v9132f8;
assign v906338 = StoB_REQ8_p & v90e261 | !StoB_REQ8_p & v844f91;
assign v909ba1 = StoB_REQ7_p & v9093ec | !StoB_REQ7_p & !v844fa1;
assign v93fe36 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9d;
assign v93f838 = jx1_p & v9093ec | !jx1_p & v911509;
assign v90f1b8 = BtoS_ACK6_p & v93f9c6 | !BtoS_ACK6_p & v90e76a;
assign v8a924b = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & v93fafd;
assign v90de0e = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & !v907200;
assign v90d7d2 = EMPTY_p & v909197 | !EMPTY_p & v9085f5;
assign v90926e = RtoB_ACK0_p & v9042d2 | !RtoB_ACK0_p & v908df3;
assign v93fb5f = StoB_REQ7_p & v90479e | !StoB_REQ7_p & v93f1cf;
assign v90f7ce = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9133b0;
assign v93ef01 = BtoS_ACK6_p & v93f1cf | !BtoS_ACK6_p & v87f17d;
assign v93ea4f = jx1_p & v90d879 | !jx1_p & v844f91;
assign v93db12 = StoB_REQ8_p & v93fbe4 | !StoB_REQ8_p & v909a21;
assign v93fa6d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v90dca4;
assign v93f6e2 = jx2_p & v93f64f | !jx2_p & v87c503;
assign v91315c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8d371f;
assign v903fb0 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8f3869;
assign v93fdfb = StoB_REQ0_p & v844f97 | !StoB_REQ0_p & v844f91;
assign v93daf2 = BtoS_ACK9_p & v903b7c | !BtoS_ACK9_p & v93f2a2;
assign v907751 = jx1_p & v844f91 | !jx1_p & !v866af4;
assign v912291 = jx1_p & v9121b6 | !jx1_p & v90dcfd;
assign v93e800 = StoB_REQ8_p & v90897e | !StoB_REQ8_p & !v844f91;
assign v90a2aa = jx2_p & v90d7ce | !jx2_p & v8b9dff;
assign v93fb66 = jx1_p & v93e819 | !jx1_p & v844f91;
assign v90ed2f = BtoS_ACK1_p & v93deab | !BtoS_ACK1_p & v93fadc;
assign v8a8faa = DEQ_p & v844fa9 | !DEQ_p & !v844f91;
assign v9099e8 = StoB_REQ7_p & v906256 | !StoB_REQ7_p & v908e73;
assign v90ed6e = StoB_REQ8_p & v9071ed | !StoB_REQ8_p & v90a96f;
assign v85eacf = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93fc78;
assign v9070cb = jx1_p & v91ae94 | !jx1_p & !v912d04;
assign v9132d6 = BtoS_ACK6_p & v90630d | !BtoS_ACK6_p & v93000b;
assign v904132 = BtoS_ACK7_p & v909bbd | !BtoS_ACK7_p & !v906e04;
assign v9051da = StoB_REQ9_p & v93fd76 | !StoB_REQ9_p & v8b9c52;
assign v908a4f = StoB_REQ8_p & v908138 | !StoB_REQ8_p & v90fd1c;
assign v910d56 = jx2_p & v90cfda | !jx2_p & v8a8fdd;
assign v910416 = BtoS_ACK9_p & v90f2f4 | !BtoS_ACK9_p & v93fbc7;
assign v93e05f = StoB_REQ8_p & v93f73d | !StoB_REQ8_p & v89e122;
assign v85eb2b = BtoR_REQ1_p & v93f0bf | !BtoR_REQ1_p & v91336b;
assign v90479e = jx0_p & v844f9b | !jx0_p & !v905366;
assign v90534f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v87a979 = StoB_REQ6_p & v904765 | !StoB_REQ6_p & v93f6b8;
assign v93db1d = jx2_p & v93f30c | !jx2_p & v93f768;
assign v90cfd5 = EMPTY_p & v9081c2 | !EMPTY_p & !v86e7cf;
assign v909705 = BtoS_ACK6_p & v9058f3 | !BtoS_ACK6_p & v9044b8;
assign v9133ea = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v90919c;
assign v9094ed = StoB_REQ1_p & v90a97c | !StoB_REQ1_p & v910380;
assign v905511 = BtoS_ACK9_p & v93fd7a | !BtoS_ACK9_p & v91a9b7;
assign v93f04f = jx2_p & v9118a3 | !jx2_p & !v90cbec;
assign v9062b5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v904e16;
assign v91aa2a = RtoB_ACK0_p & v908ed2 | !RtoB_ACK0_p & v93e193;
assign v904dc1 = ENQ_p & v93f15e | !ENQ_p & v910915;
assign v889d4b = RtoB_ACK0_p & v93f959 | !RtoB_ACK0_p & v90738c;
assign v86e433 = StoB_REQ1_p & v913619 | !StoB_REQ1_p & v90fc92;
assign v863a47 = jx1_p & v913332 | !jx1_p & v93fcc9;
assign v93fbc1 = RtoB_ACK0_p & v93f899 | !RtoB_ACK0_p & v90e437;
assign v93eb1d = stateG7_1_p & v93f7d5 | !stateG7_1_p & v90ea98;
assign v90827d = StoB_REQ2_p & v8b98bd | !StoB_REQ2_p & !v93f928;
assign v90968f = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v93f825;
assign v8f3853 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v910bd7;
assign v906d2a = jx1_p & v9074ce | !jx1_p & v844f91;
assign v93fa99 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v89f82d;
assign v93e7d4 = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & !v93fc63;
assign v87a253 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v903b7d;
assign v90ee6d = StoB_REQ6_p & v8b98be | !StoB_REQ6_p & v93fc7d;
assign v9084ae = jx2_p & v909b54 | !jx2_p & v844f91;
assign v93f7f0 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v93f7b8;
assign v908d14 = jx1_p & v93e288 | !jx1_p & v93f71d;
assign v85ea4f = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v93fd4c;
assign v90474e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90f810;
assign v903b56 = ENQ_p & v91a6d3 | !ENQ_p & !v93f917;
assign v87c21e = jx1_p & v93f1b4 | !jx1_p & v908f27;
assign v93f324 = StoB_REQ7_p & v93e655 | !StoB_REQ7_p & v9102cc;
assign v909383 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v90fe49;
assign v8857fd = StoB_REQ0_p & v93f7f5 | !StoB_REQ0_p & v90e7d7;
assign v905dcf = jx1_p & v904fe6 | !jx1_p & !v86fe09;
assign v85acd3 = BtoS_ACK8_p & v93dbe9 | !BtoS_ACK8_p & v9043c2;
assign v90a241 = FULL_p & v907bd1 | !FULL_p & v91a9a2;
assign v911951 = stateG7_1_p & v844f91 | !stateG7_1_p & v909722;
assign v9102aa = jx2_p & v904bd4 | !jx2_p & v844f91;
assign v9103b5 = BtoS_ACK0_p & v93fdfe | !BtoS_ACK0_p & v8a9209;
assign v93fcc2 = jx2_p & v91143f | !jx2_p & v9119f9;
assign v93e193 = ENQ_p & v8f2274 | !ENQ_p & v844f91;
assign v93e7d1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90eef9;
assign v90d0fd = BtoS_ACK6_p & v9056bd | !BtoS_ACK6_p & v910469;
assign v93fd2c = BtoS_ACK6_p & v90630d | !BtoS_ACK6_p & !v903c43;
assign v908a2c = BtoS_ACK7_p & v90d879 | !BtoS_ACK7_p & v910e32;
assign v93e03a = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v844f91;
assign v911cba = BtoS_ACK8_p & v93e27a | !BtoS_ACK8_p & v904ab4;
assign v904ae4 = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v93f7ff;
assign v93e1c0 = jx1_p & v911edb | !jx1_p & v909b74;
assign v93e45c = BtoS_ACK6_p & v909f04 | !BtoS_ACK6_p & v903d4f;
assign v93f93c = jx1_p & v93e0b5 | !jx1_p & v844f91;
assign v907b54 = ENQ_p & v93f89f | !ENQ_p & v906c0f;
assign v93f5c0 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v9074a6;
assign v9099e3 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v907168;
assign v8a928a = BtoR_REQ1_p & v91229e | !BtoR_REQ1_p & v911328;
assign v90d8f3 = StoB_REQ9_p & v93e701 | !StoB_REQ9_p & v903c0d;
assign v93e48f = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v87b4fc;
assign v8639e7 = BtoS_ACK6_p & v9050a5 | !BtoS_ACK6_p & v93fa28;
assign v9106a7 = StoB_REQ7_p & v93fe2e | !StoB_REQ7_p & v9074ce;
assign v8b9dff = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90d879;
assign v8ee1f5 = StoB_REQ0_p & v93f7f5 | !StoB_REQ0_p & v903fee;
assign v90a314 = jx1_p & v93de80 | !jx1_p & v87f17d;
assign v93fb14 = jx0_p & v93fa4f | !jx0_p & v90690e;
assign v9109ee = StoB_REQ2_p & v907168 | !StoB_REQ2_p & v93f8f8;
assign v904303 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v909492;
assign v93fa16 = jx1_p & v9093ec | !jx1_p & !v90df7f;
assign v93eb43 = jx2_p & v93dee0 | !jx2_p & !v93fbf3;
assign v90eed7 = BtoS_ACK7_p & v87f17d | !BtoS_ACK7_p & v912481;
assign v90fbc8 = BtoS_ACK9_p & v907da6 | !BtoS_ACK9_p & v93f896;
assign v90f2f6 = BtoS_ACK9_p & v910c51 | !BtoS_ACK9_p & v93fa51;
assign v906c2f = jx2_p & v907995 | !jx2_p & v9113fb;
assign v90e6f5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v910ff7;
assign v88e55e = jx2_p & v93fac8 | !jx2_p & v90cb3d;
assign v90fa41 = StoB_REQ3_p & v904182 | !StoB_REQ3_p & v9300af;
assign v93f28c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fc46;
assign v93ebab = BtoS_ACK9_p & v9134cc | !BtoS_ACK9_p & v908fd6;
assign v9107aa = jx2_p & v93f4cd | !jx2_p & !v90ded0;
assign v90fc5e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85ea99;
assign v93e6e0 = jx0_p & v93f962 | !jx0_p & v844f91;
assign v9135db = jx1_p & v93defa | !jx1_p & v8b5f4d;
assign v93f7f6 = jx1_p & v844f91 | !jx1_p & v9096f3;
assign v93fc75 = BtoS_ACK6_p & v907ce3 | !BtoS_ACK6_p & v93f8bb;
assign v93f664 = jx0_p & v93f723 | !jx0_p & v844f91;
assign v86345c = StoB_REQ2_p & v908127 | !StoB_REQ2_p & v8b98fe;
assign v93efa3 = jx1_p & v90d81c | !jx1_p & v844f91;
assign v90ff07 = BtoS_ACK9_p & v8f3825 | !BtoS_ACK9_p & v93fd1c;
assign v909e90 = BtoS_ACK8_p & v90d3ff | !BtoS_ACK8_p & v90e2d7;
assign v93fac8 = jx1_p & v911edb | !jx1_p & v93f7e5;
assign v909a7b = StoB_REQ8_p & v93fbe4 | !StoB_REQ8_p & v93faab;
assign v906570 = EMPTY_p & v8bbc54 | !EMPTY_p & v9130c5;
assign v905486 = RtoB_ACK0_p & v93f98d | !RtoB_ACK0_p & v93f9cb;
assign v91082c = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v93f7bb;
assign v9056ad = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v906642;
assign v909312 = BtoS_ACK9_p & v8b9e96 | !BtoS_ACK9_p & v908aae;
assign v906c8b = jx1_p & v93fc94 | !jx1_p & v90d22b;
assign v93faf8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90962d;
assign v90f3f8 = BtoS_ACK8_p & v93f279 | !BtoS_ACK8_p & v90da35;
assign v90423b = jx1_p & v869aeb | !jx1_p & !v90efea;
assign v909546 = RtoB_ACK1_p & v85eb14 | !RtoB_ACK1_p & !v93fd98;
assign v89e119 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v904af3;
assign v906a5c = jx1_p & v869aeb | !jx1_p & !v93f76b;
assign v906b3d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v906d41;
assign v910490 = BtoS_ACK8_p & v87f17f | !BtoS_ACK8_p & v93fd95;
assign v8b9e96 = StoB_REQ8_p & v904b00 | !StoB_REQ8_p & v90a733;
assign v9098a3 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v93ec67;
assign v93f68c = StoB_REQ1_p & v92ffda | !StoB_REQ1_p & v93ef2e;
assign v93fc1f = BtoS_ACK8_p & v9132eb | !BtoS_ACK8_p & !v91097b;
assign v90a4e6 = StoB_REQ6_p & v90a8e9 | !StoB_REQ6_p & v8b99bb;
assign v904e48 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9062f7;
assign v8a8b0a = jx0_p & v93f738 | !jx0_p & !v904adb;
assign v93fcbf = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93f29a;
assign v907102 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v903fee;
assign v909f7e = StoB_REQ1_p & v90a20d | !StoB_REQ1_p & v912f42;
assign v904f52 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v908a34;
assign v8f22d1 = StoB_REQ7_p & v910710 | !StoB_REQ7_p & !v844f91;
assign v93fe73 = BtoS_ACK9_p & v93e85e | !BtoS_ACK9_p & v9042a0;
assign v93f155 = BtoS_ACK1_p & v93fce7 | !BtoS_ACK1_p & !v90759b;
assign v90da92 = BtoS_ACK6_p & v90a786 | !BtoS_ACK6_p & v93f90e;
assign v93e90d = jx2_p & v908a03 | !jx2_p & v93e13e;
assign v93f7e3 = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v908000;
assign v90f1b9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v912ef3;
assign v863a97 = RtoB_ACK0_p & v93f680 | !RtoB_ACK0_p & v87a203;
assign v93f731 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fb2e;
assign v85ea72 = RtoB_ACK0_p & v90e361 | !RtoB_ACK0_p & v910525;
assign v90515a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9070d5;
assign v9073c5 = StoB_REQ8_p & v93f73d | !StoB_REQ8_p & v90451f;
assign v93fae3 = jx1_p & v89e11b | !jx1_p & v844f91;
assign v90466e = StoB_REQ2_p & v93fdf7 | !StoB_REQ2_p & v9098f2;
assign v90a733 = jx2_p & v8b9bd9 | !jx2_p & v8b9dff;
assign v93e1ed = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93e439;
assign v89e08c = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v872442;
assign v93fc7d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f7ad;
assign v93f735 = jx2_p & v844f91 | !jx2_p & v93f855;
assign v907e36 = BtoS_ACK7_p & v907815 | !BtoS_ACK7_p & v8b9c55;
assign v90e978 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f9d;
assign v90e172 = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v8a9205;
assign v9054bc = StoB_REQ0_p & v910bd7 | !StoB_REQ0_p & !v91141d;
assign v910840 = BtoS_ACK9_p & v9114a0 | !BtoS_ACK9_p & v93f90d;
assign v844fa1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f91;
assign v93fa05 = BtoS_ACK8_p & v905e43 | !BtoS_ACK8_p & !v9110a7;
assign v911724 = BtoS_ACK6_p & v93f90a | !BtoS_ACK6_p & v85ea76;
assign v91093d = ENQ_p & v9093d9 | !ENQ_p & v844f91;
assign v93e281 = EMPTY_p & v904b99 | !EMPTY_p & v9114cf;
assign v93fa4c = StoB_REQ7_p & v93f9c6 | !StoB_REQ7_p & v844f91;
assign v908107 = BtoS_ACK6_p & v9047e4 | !BtoS_ACK6_p & !v90fb2b;
assign v93f7a1 = stateG12_p & v844fc3 | !stateG12_p & !v905291;
assign v906255 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v90e978;
assign v93f314 = StoB_REQ9_p & v93f8f4 | !StoB_REQ9_p & v91a73f;
assign v9091a2 = BtoR_REQ0_p & v93e037 | !BtoR_REQ0_p & v906275;
assign v93fa90 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v90a6f4;
assign v906dd6 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93ef4c;
assign v903d21 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v906024;
assign v912f42 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v93f7ce;
assign v93f6c9 = jx2_p & v904bd4 | !jx2_p & v90824f;
assign v9068b7 = jx0_p & v844f91 | !jx0_p & v863a78;
assign v90f66c = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v90ed41;
assign v910f3a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v905d28;
assign v911853 = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v93fbcf;
assign v9083cf = jx3_p & v9084d0 | !jx3_p & !v90e772;
assign v93e6fe = BtoS_ACK9_p & v93e228 | !BtoS_ACK9_p & !v93fcf9;
assign v93ebd1 = BtoS_ACK0_p & v93fccb | !BtoS_ACK0_p & v8b99b9;
assign v93e76f = jx1_p & v90980d | !jx1_p & v90db9f;
assign v93fcf3 = jx0_p & v863b25 | !jx0_p & v844f91;
assign v904fb4 = BtoS_ACK9_p & v93fcbf | !BtoS_ACK9_p & v93fb7a;
assign v8b9ecf = ENQ_p & v90adc4 | !ENQ_p & v93fafc;
assign v90f0bd = ENQ_p & v93f15e | !ENQ_p & v9104f8;
assign v8b9bd8 = StoB_REQ8_p & v93fc04 | !StoB_REQ8_p & v89e07c;
assign v930114 = BtoR_REQ1_p & v93fbec | !BtoR_REQ1_p & v93e9dd;
assign v90930e = BtoS_ACK9_p & v906338 | !BtoS_ACK9_p & v93fa69;
assign v911b4e = StoB_REQ8_p & v93fd8d | !StoB_REQ8_p & v906c91;
assign v90edd1 = EMPTY_p & v9076cf | !EMPTY_p & v93fe21;
assign v90d662 = BtoS_ACK7_p & v9133ba | !BtoS_ACK7_p & !v906cc5;
assign v93f8d1 = BtoS_ACK0_p & v90a5ef | !BtoS_ACK0_p & v93f75c;
assign v9082be = ENQ_p & v93f753 | !ENQ_p & v844f91;
assign v904f64 = jx0_p & v90549c | !jx0_p & v93fa9c;
assign v88403f = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v93fa22;
assign v904568 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ee1a3;
assign v93f28a = jx0_p & v85eaab | !jx0_p & v844f91;
assign v90d5d1 = DEQ_p & v93fb11 | !DEQ_p & v9075e7;
assign v910e82 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93eb13;
assign v93fa7c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93e391;
assign v913399 = RtoB_ACK0_p & v9096ca | !RtoB_ACK0_p & v93f56e;
assign v93fb7a = StoB_REQ9_p & v909c39 | !StoB_REQ9_p & v91a6f0;
assign v93fd9a = jx0_p & v90762a | !jx0_p & v905ffe;
assign v903f97 = jx1_p & v93fcfc | !jx1_p & !v93fb3e;
assign v9110a7 = StoB_REQ8_p & v9071ed | !StoB_REQ8_p & v93e886;
assign v93fa76 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8714f5;
assign v907995 = jx1_p & v90d880 | !jx1_p & v91a9b9;
assign v93f6fd = BtoS_ACK2_p & v906cc8 | !BtoS_ACK2_p & v93eec4;
assign v8f22ea = StoB_REQ0_p & v93db4a | !StoB_REQ0_p & v90aa64;
assign v93e9b9 = StoB_REQ8_p & v90f83a | !StoB_REQ8_p & v905461;
assign v89c580 = BtoS_ACK7_p & v90dec8 | !BtoS_ACK7_p & !v93eba3;
assign v93e4b9 = BtoS_ACK7_p & v93f8c5 | !BtoS_ACK7_p & v8b9d35;
assign v93ef13 = StoB_REQ7_p & v907da3 | !StoB_REQ7_p & v90a430;
assign v89f927 = stateG7_1_p & v880d77 | !stateG7_1_p & v907b01;
assign v93f6b6 = RtoB_ACK1_p & v909efe | !RtoB_ACK1_p & v93fb80;
assign v93fd5f = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v93f74a;
assign v905d7e = StoB_REQ7_p & v903fb2 | !StoB_REQ7_p & v93fa8f;
assign v9083c5 = BtoS_ACK8_p & v93faab | !BtoS_ACK8_p & v93fdf3;
assign v908410 = jx1_p & v8b9dff | !jx1_p & v910bf9;
assign v87b42f = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v90e76a;
assign v9045bb = StoB_REQ7_p & v905ba8 | !StoB_REQ7_p & v844f91;
assign v93f634 = jx3_p & v93fdda | !jx3_p & v906b4a;
assign v910b91 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v906492;
assign v90765f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9062b3;
assign v905775 = jx2_p & v8a8f5e | !jx2_p & v844f91;
assign v8b49bf = ENQ_p & v90fbad | !ENQ_p & v90e315;
assign v910495 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v9123a2;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v91071e = BtoS_ACK0_p & v913619 | !BtoS_ACK0_p & v88c832;
assign v90e339 = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v90d84e;
assign v9101b8 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v93e652;
assign v8b9ce2 = BtoS_ACK8_p & v909a21 | !BtoS_ACK8_p & v904eea;
assign v93f148 = jx1_p & v844f91 | !jx1_p & !v91879a;
assign v93e14f = jx0_p & v93f7b7 | !jx0_p & !v93fd94;
assign v90d46a = StoB_REQ7_p & v906320 | !StoB_REQ7_p & v903c1c;
assign v93ed1c = StoB_REQ9_p & v910490 | !StoB_REQ9_p & v90d370;
assign v93ec81 = BtoS_ACK2_p & v90854b | !BtoS_ACK2_p & v86345c;
assign v93f064 = StoB_REQ0_p & v87052e | !StoB_REQ0_p & v93eb41;
assign v90667d = BtoS_ACK6_p & v90ede1 | !BtoS_ACK6_p & v93fa4b;
assign v93fc9b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93e77b;
assign v90e612 = BtoS_ACK7_p & v93fb38 | !BtoS_ACK7_p & v90a3f5;
assign v909d9c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fa9d;
assign v93fb88 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v86337d;
assign v90a604 = BtoS_ACK7_p & v90f8d6 | !BtoS_ACK7_p & v93fcc1;
assign v908346 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v93fd9b;
assign v93f871 = jx0_p & v844f91 | !jx0_p & v93fce5;
assign v90f391 = BtoS_ACK9_p & v90dec9 | !BtoS_ACK9_p & v909c3b;
assign v908edf = StoB_REQ9_p & v909e90 | !StoB_REQ9_p & v907299;
assign v9041e6 = BtoS_ACK6_p & v9058f3 | !BtoS_ACK6_p & v93fdce;
assign v905adf = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v904182;
assign v93f9b4 = BtoS_ACK0_p & v9052de | !BtoS_ACK0_p & v90ae53;
assign v90dcca = ENQ_p & v93f89f | !ENQ_p & v906fd0;
assign v93fb93 = jx2_p & v909cea | !jx2_p & v90da8b;
assign v911c0f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b49f1;
assign v906b22 = StoB_REQ9_p & v907c76 | !StoB_REQ9_p & v913068;
assign v904fc8 = StoB_REQ1_p & v90e611 | !StoB_REQ1_p & v93ec07;
assign v93fd1b = ENQ_p & v90fe92 | !ENQ_p & v85f28b;
assign v92ffc9 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v8b9eb0;
assign v93f589 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v89f9da;
assign v909f00 = BtoS_ACK8_p & v93fe3f | !BtoS_ACK8_p & v9100b7;
assign v93fd3b = DEQ_p & v90752d | !DEQ_p & v93fb21;
assign v9080a8 = StoB_REQ3_p & v9048d7 | !StoB_REQ3_p & !v844f9f;
assign v910704 = RtoB_ACK1_p & v90561f | !RtoB_ACK1_p & v93f767;
assign v9081ef = BtoS_ACK9_p & v9044c3 | !BtoS_ACK9_p & v93e5d4;
assign v93fd43 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f812;
assign v908805 = BtoS_ACK0_p & v93fdfe | !BtoS_ACK0_p & v93f7fa;
assign v93f7fc = StoB_REQ9_p & v90620e | !StoB_REQ9_p & v844f91;
assign v906d58 = jx0_p & v90ef1b | !jx0_p & v93f6d5;
assign v93fb73 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90a1fd;
assign v90d443 = stateG7_1_p & v863359 | !stateG7_1_p & v90cf68;
assign v93f279 = jx2_p & v913592 | !jx2_p & !v904755;
assign v8b9ba5 = StoB_REQ8_p & v90ddf9 | !StoB_REQ8_p & v93f78a;
assign v90a61d = jx3_p & v90a1c6 | !jx3_p & v8a1fe3;
assign v90f2f9 = jx2_p & v8b49dc | !jx2_p & v90986f;
assign v9046a7 = StoB_REQ9_p & v903c0d | !StoB_REQ9_p & !v844f91;
assign v89f7dd = StoB_REQ8_p & v93f7f8 | !StoB_REQ8_p & v93e007;
assign v9110ab = jx1_p & v9062f7 | !jx1_p & v90468e;
assign v93fe21 = DEQ_p & v93e2a0 | !DEQ_p & v85f2b0;
assign v93e31b = BtoS_ACK9_p & v93db12 | !BtoS_ACK9_p & v9104bd;
assign v91306c = RtoB_ACK0_p & v907b54 | !RtoB_ACK0_p & v8b9e97;
assign v9087b1 = BtoS_ACK6_p & v910230 | !BtoS_ACK6_p & v93faa1;
assign v93f765 = StoB_REQ3_p & v89f840 | !StoB_REQ3_p & v844f91;
assign v93de99 = jx2_p & v93eda5 | !jx2_p & v844f91;
assign v9098ab = BtoS_ACK6_p & v8b9d27 | !BtoS_ACK6_p & v93f5e9;
assign v910221 = EMPTY_p & v9077f6 | !EMPTY_p & v8633df;
assign v90dcfd = StoB_REQ7_p & v908e8e | !StoB_REQ7_p & v9121b6;
assign v906d53 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v844f91;
assign v89f7e3 = BtoS_ACK8_p & v904bc1 | !BtoS_ACK8_p & v93ec8c;
assign v91053d = BtoS_ACK8_p & v8b5f61 | !BtoS_ACK8_p & !v91ddca;
assign v913079 = RtoB_ACK1_p & v9070f7 | !RtoB_ACK1_p & v873a26;
assign v89e07c = jx2_p & v93f389 | !jx2_p & v911c6f;
assign v93fd35 = jx1_p & v90f5ff | !jx1_p & v844f91;
assign v9067d3 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v910f5a;
assign v93eabc = BtoS_ACK7_p & v93f7f8 | !BtoS_ACK7_p & v907f0b;
assign v91267b = BtoS_ACK8_p & v90451f | !BtoS_ACK8_p & v90d6ef;
assign v93fd98 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v90cfd5;
assign v93f6c4 = EMPTY_p & v8a9250 | !EMPTY_p & v93f729;
assign v903b7b = StoB_REQ7_p & v8b4a08 | !StoB_REQ7_p & v844f91;
assign v904e00 = StoB_REQ9_p & v90a784 | !StoB_REQ9_p & v905a21;
assign v863b1a = jx1_p & v869aeb | !jx1_p & !v90ebde;
assign v9062f7 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v913435;
assign v903e94 = jx0_p & v844f9f | !jx0_p & !v844f91;
assign v90f36b = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v90deaa;
assign v93e9c7 = BtoS_ACK0_p & v9046a6 | !BtoS_ACK0_p & v90f38b;
assign v90901d = BtoS_ACK6_p & v93f63b | !BtoS_ACK6_p & v905636;
assign v93fcd0 = jx1_p & v844fa1 | !jx1_p & !v844f91;
assign v9068c8 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v8f37f1;
assign v93fa58 = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v93fb5d;
assign v93f945 = StoB_REQ0_p & v909058 | !StoB_REQ0_p & v9115b6;
assign v90e140 = EMPTY_p & v90775f | !EMPTY_p & v90575e;
assign v90a97c = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v90ba2c;
assign v911909 = StoB_REQ8_p & v93e27a | !StoB_REQ8_p & v91a799;
assign v93f6ad = StoB_REQ9_p & v909e8a | !StoB_REQ9_p & v89e086;
assign v908e7e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b8638;
assign v93fbe4 = jx2_p & v9097da | !jx2_p & v8f60f9;
assign v9086f1 = DEQ_p & v910ffd | !DEQ_p & v93fb72;
assign v93f6a2 = StoB_REQ7_p & v910243 | !StoB_REQ7_p & v844f91;
assign v908f48 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93fd32;
assign v90f16d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90d877;
assign v908209 = jx1_p & v91ae94 | !jx1_p & v90e339;
assign v93f3db = jx0_p & v904ed4 | !jx0_p & !v85f258;
assign v9132ed = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90798e;
assign v90fc6d = StoB_REQ7_p & v93f796 | !StoB_REQ7_p & v91aa06;
assign v9044c9 = jx2_p & v930083 | !jx2_p & v93fd89;
assign v90f9b6 = StoB_REQ0_p & v910bd7 | !StoB_REQ0_p & !v90aa64;
assign v903c1f = StoB_REQ8_p & v93ec28 | !StoB_REQ8_p & !v93dc87;
assign v93f8a3 = DEQ_p & v904b94 | !DEQ_p & v904c4f;
assign v91a6e9 = ENQ_p & v93e704 | !ENQ_p & v93fd73;
assign v906a84 = jx3_p & v844f91 | !jx3_p & v87c4c4;
assign v93fbaf = stateG12_p & v93f15e | !stateG12_p & v904ebe;
assign v90dcb3 = jx2_p & v90d93b | !jx2_p & v91aa3f;
assign v908aae = StoB_REQ9_p & v93f7ab | !StoB_REQ9_p & v90ccbd;
assign v93f764 = BtoS_ACK8_p & v90529c | !BtoS_ACK8_p & v93fd8a;
assign v90a0e8 = BtoS_ACK0_p & v90534f | !BtoS_ACK0_p & v909666;
assign v90f4f7 = RtoB_ACK1_p & v9100a9 | !RtoB_ACK1_p & v93fc5a;
assign v86dd54 = BtoS_ACK7_p & v9084ae | !BtoS_ACK7_p & v93fdbf;
assign v93e37e = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v90e526;
assign v8b9c31 = jx2_p & v904988 | !jx2_p & v93fcba;
assign v90561f = BtoR_REQ0_p & v93f10b | !BtoR_REQ0_p & v93dffa;
assign v909b01 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v90dc0a;
assign v904c75 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v9077a9;
assign v93fb34 = RtoB_ACK0_p & v907bd1 | !RtoB_ACK0_p & v90a241;
assign v906df1 = StoB_REQ9_p & v93f088 | !StoB_REQ9_p & v904ba4;
assign v93fc7b = BtoS_ACK7_p & v93fb78 | !BtoS_ACK7_p & v90a75f;
assign v93fd9f = jx1_p & v930047 | !jx1_p & !v844f91;
assign v90980d = jx0_p & v93fcbe | !jx0_p & v93fce5;
assign v9100a9 = BtoR_REQ0_p & v905dc0 | !BtoR_REQ0_p & v93fc42;
assign v93f6e1 = StoB_REQ6_p & v906ae9 | !StoB_REQ6_p & v93f2a0;
assign v9084ef = jx0_p & v90664a | !jx0_p & v93f6fc;
assign v9075db = StoB_REQ2_p & v87b4fc | !StoB_REQ2_p & v844f91;
assign v93f7b8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85eabe;
assign v906ce5 = EMPTY_p & v904bc0 | !EMPTY_p & v9089ef;
assign v93e8f6 = jx0_p & v844fa1 | !jx0_p & !v844f91;
assign v87ba4e = ENQ_p & v911b74 | !ENQ_p & v844f91;
assign v910b4b = BtoS_ACK7_p & v8807b1 | !BtoS_ACK7_p & !v844fa3;
assign v93fdaa = BtoS_ACK8_p & v90512d | !BtoS_ACK8_p & v90a4bf;
assign v93fb07 = BtoS_ACK6_p & v93fcfc | !BtoS_ACK6_p & v8ebce4;
assign v93f8f4 = BtoS_ACK8_p & v9134bc | !BtoS_ACK8_p & v90e2d7;
assign v9057f8 = StoB_REQ8_p & v93f769 | !StoB_REQ8_p & v904345;
assign v90536f = BtoS_ACK9_p & v844f91 | !BtoS_ACK9_p & v93f7fc;
assign v93e33e = StoB_REQ0_p & v910bd7 | !StoB_REQ0_p & !v844f91;
assign v93fe35 = jx3_p & v844f91 | !jx3_p & v904b00;
assign v907815 = jx2_p & v905408 | !jx2_p & v93fa1e;
assign v91231a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9056f9;
assign v9107e7 = BtoS_ACK8_p & v93fbe4 | !BtoS_ACK8_p & v93f960;
assign v93eadd = stateG7_1_p & v93f9e0 | !stateG7_1_p & v93f999;
assign BtoS_ACK3_n = !v91a7a5;
assign v910d28 = BtoS_ACK7_p & v93f9e3 | !BtoS_ACK7_p & v90fa18;
assign v90710d = EMPTY_p & v93fb21 | !EMPTY_p & v93eec9;
assign v90cf0e = BtoS_ACK9_p & v93e097 | !BtoS_ACK9_p & v93f314;
assign v90995e = BtoS_ACK1_p & v93fccb | !BtoS_ACK1_p & v91006b;
assign v909e99 = StoB_REQ8_p & v91a6ea | !StoB_REQ8_p & v93fb19;
assign v90861d = BtoS_ACK6_p & v91132f | !BtoS_ACK6_p & v93e6e0;
assign v906e3b = BtoS_ACK8_p & v90e893 | !BtoS_ACK8_p & v93f6b2;
assign BtoS_ACK6_n = !v8a928a;
assign v93ebb5 = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & !v93fc8e;
assign v93fbec = RtoB_ACK1_p & v90e906 | !RtoB_ACK1_p & v9113ea;
assign v909b74 = StoB_REQ7_p & v903f58 | !StoB_REQ7_p & v93f33e;
assign v9056d9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v903cf9;
assign v90edb8 = BtoS_ACK6_p & v90a786 | !BtoS_ACK6_p & v90917f;
assign v90a786 = jx0_p & v93ed91 | !jx0_p & v906ae9;
assign v9059a0 = BtoS_ACK1_p & v913348 | !BtoS_ACK1_p & v906195;
assign v910cee = StoB_REQ7_p & v9082ba | !StoB_REQ7_p & v90d5bd;
assign v91093c = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v90d71a;
assign v93fdd4 = BtoS_ACK1_p & v9052de | !BtoS_ACK1_p & v90a233;
assign v93f9f0 = jx2_p & v93f970 | !jx2_p & v93f1aa;
assign v905d68 = BtoS_ACK8_p & v93fb92 | !BtoS_ACK8_p & v9057f8;
assign v910380 = BtoS_ACK2_p & v90854b | !BtoS_ACK2_p & v93f840;
assign v909cea = jx1_p & v9099e1 | !jx1_p & v93fcd4;
assign v905292 = ENQ_p & v93eda4 | !ENQ_p & v90e3bf;
assign v93e048 = StoB_REQ8_p & v90d3ff | !StoB_REQ8_p & v93fdae;
assign v93f94b = EMPTY_p & v93fb21 | !EMPTY_p & v93fd13;
assign v90f7d6 = StoB_REQ6_p & v9081b9 | !StoB_REQ6_p & v93fb82;
assign v93faa1 = jx0_p & v93fc65 | !jx0_p & v8b4976;
assign v9117b1 = jx2_p & v90caf3 | !jx2_p & !v905718;
assign v8d371f = BtoS_ACK6_p & v93efbb | !BtoS_ACK6_p & v844f91;
assign v90583b = EMPTY_p & v91209b | !EMPTY_p & v93f8a3;
assign v93fcc8 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v93f8d3;
assign v9103bc = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8893bb;
assign v93f745 = StoB_REQ9_p & v905487 | !StoB_REQ9_p & v93fe0d;
assign v93f7c7 = jx0_p & v844f91 | !jx0_p & v90d59a;
assign v8b9f34 = BtoR_REQ0_p & v905170 | !BtoR_REQ0_p & v93f73a;
assign v93fbf9 = jx0_p & v93f9b4 | !jx0_p & v93fc0e;
assign v93f7af = BtoS_ACK0_p & v93e391 | !BtoS_ACK0_p & v906ff5;
assign v903f5a = BtoS_ACK8_p & v907eaa | !BtoS_ACK8_p & v908b06;
assign v90888d = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v93fb03;
assign v8f22bd = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v90decb;
assign v907d8a = BtoS_ACK9_p & v8b9e96 | !BtoS_ACK9_p & v911365;
assign v87c9b3 = EMPTY_p & v863a3f | !EMPTY_p & v910fcd;
assign v93fb74 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v90d59e;
assign v93f7ad = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v906255;
assign v909878 = ENQ_p & v8b98f1 | !ENQ_p & v905da0;
assign v90e433 = BtoS_ACK6_p & v90ad75 | !BtoS_ACK6_p & v93f91a;
assign v88c832 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90fe5c;
assign v911102 = StoB_REQ1_p & v9046a6 | !StoB_REQ1_p & v93fce7;
assign v85de34 = BtoS_ACK6_p & v910e72 | !BtoS_ACK6_p & v844f91;
assign v93f702 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v913619;
assign v8b6009 = BtoR_REQ0_p & v90edd1 | !BtoR_REQ0_p & v93e852;
assign v93f678 = jx1_p & v869aeb | !jx1_p & !v910fd8;
assign v93fce0 = StoB_REQ2_p & v90d9fd | !StoB_REQ2_p & v91082c;
assign v903b7d = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v93fb3a;
assign v93f1a6 = jx3_p & v93e7af | !jx3_p & v909fd6;
assign v88b9b7 = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v903c5b;
assign v905194 = jx0_p & v93f29e | !jx0_p & v87283f;
assign v93e5fc = StoB_REQ1_p & v908df7 | !StoB_REQ1_p & !v93f6a7;
assign v93f5d9 = BtoS_ACK9_p & v90f2f4 | !BtoS_ACK9_p & v87a242;
assign v93f912 = BtoS_ACK9_p & v909a7b | !BtoS_ACK9_p & v93f5db;
assign v907b21 = StoB_REQ1_p & v93fc28 | !StoB_REQ1_p & v9106af;
assign v93f860 = jx1_p & v9099ee | !jx1_p & v90ad75;
assign v93fd3d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93e2de;
assign v93f7f5 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v90fe49;
assign v89f8e5 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v89c59e;
assign v93fa2a = BtoS_ACK8_p & v90a229 | !BtoS_ACK8_p & v905653;
assign v89f840 = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v844fbb;
assign v87c533 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v90f547;
assign v93fa3c = StoB_REQ6_p & v9067d3 | !StoB_REQ6_p & v8ebcf9;
assign v93ed6a = jx1_p & v87f17d | !jx1_p & v93f6cc;
assign v90569e = BtoS_ACK0_p & v910f6e | !BtoS_ACK0_p & v906414;
assign v90fcbf = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & v9063e0;
assign v93f916 = ENQ_p & v8a1fe3 | !ENQ_p & v93fc32;
assign v9093ec = jx0_p & v844f91 | !jx0_p & !v844fa1;
assign v89f93b = BtoS_ACK0_p & v93f7ad | !BtoS_ACK0_p & v93f821;
assign v9103e5 = ENQ_p & v93f753 | !ENQ_p & !v93f784;
assign v9060c1 = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v8ee1c7;
assign v908d05 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v93e896;
assign v904f23 = RtoB_ACK0_p & v93fc6a | !RtoB_ACK0_p & v93f783;
assign v93f7fa = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f853;
assign v90e2e7 = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & v905838;
assign v8b98be = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90deff;
assign v93effa = BtoS_ACK7_p & v90eef9 | !BtoS_ACK7_p & v8b9eca;
assign v88b606 = StoB_REQ7_p & v907da3 | !StoB_REQ7_p & v844f91;
assign v85ea7f = BtoS_ACK0_p & v93f5d1 | !BtoS_ACK0_p & v90acc4;
assign v8821a1 = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v93fb14;
assign BtoS_ACK5_n = !v930114;
assign v904dd8 = StoB_REQ6_p & v93db03 | !StoB_REQ6_p & v90569e;
assign v93e80c = RtoB_ACK0_p & v93fc48 | !RtoB_ACK0_p & v905292;
assign v93df31 = jx3_p & v87ec92 | !jx3_p & v93f89f;
assign v910403 = jx1_p & v93fd1a | !jx1_p & v911880;
assign v90decb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93e95e;
assign v93f893 = jx3_p & v9072b7 | !jx3_p & v93eed6;
assign v93fa35 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v93fb9c;
assign v93fe54 = BtoS_ACK9_p & v93f9bb | !BtoS_ACK9_p & v9067ab;
assign v93f729 = DEQ_p & v912d1a | !DEQ_p & v90542e;
assign v86f729 = StoB_REQ0_p & v9071c7 | !StoB_REQ0_p & v844f91;
assign v90cbf3 = jx3_p & v908429 | !jx3_p & v93f07c;
assign v863b37 = jx1_p & v930032 | !jx1_p & v909f04;
assign v93f389 = jx1_p & v93fd9e | !jx1_p & v844f91;
assign v909eb5 = stateG7_1_p & v909722 | !stateG7_1_p & v844f91;
assign v93f9ff = DEQ_p & v87e0d8 | !DEQ_p & v93f29c;
assign v93fe07 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v93fb31 = BtoS_ACK1_p & v86c2d0 | !BtoS_ACK1_p & v93f908;
assign v90a620 = jx0_p & v844f91 | !jx0_p & v9074ce;
assign v90a4c6 = BtoS_ACK6_p & v90a786 | !BtoS_ACK6_p & v844f91;
assign v93005b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v93f70c;
assign v93f787 = jx2_p & v908209 | !jx2_p & v909661;
assign v9117db = StoB_REQ7_p & v93fc2b | !StoB_REQ7_p & v907bca;
assign v90638b = BtoS_ACK7_p & v904b00 | !BtoS_ACK7_p & v9095ec;
assign v90ae9a = jx1_p & v9051bb | !jx1_p & v906c66;
assign v87a25e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85ea4f;
assign v91035c = BtoS_ACK8_p & v9062f7 | !BtoS_ACK8_p & v93fd06;
assign v93f7ea = jx0_p & v93db03 | !jx0_p & v90a7b2;
assign v911383 = BtoS_ACK6_p & v909187 | !BtoS_ACK6_p & !v908e7c;
assign v90ad69 = jx2_p & v93f87a | !jx2_p & v908322;
assign v93ca43 = jx2_p & v93e335 | !jx2_p & v93fe75;
assign v863477 = jx0_p & v8b9c5f | !jx0_p & v906df6;
assign v93fac2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8b9e6c;
assign v93fc19 = BtoS_ACK6_p & v8ee17f | !BtoS_ACK6_p & v93fb0f;
assign v93fe45 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v85f278;
assign v93fc78 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v91305b;
assign v93fa5e = DEQ_p & v9077f7 | !DEQ_p & v9047b1;
assign v93fc26 = DEQ_p & v90744a | !DEQ_p & v93f29c;
assign v9054b6 = ENQ_p & v93df31 | !ENQ_p & v90d86f;
assign v90d6e8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v93f70c;
assign v93fb3a = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v930097;
assign v8b9e9f = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v90eab9;
assign v90a47f = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v906b66;
assign v91355f = StoB_REQ8_p & v93f769 | !StoB_REQ8_p & v910d99;
assign v908f4b = BtoS_ACK8_p & v8b9dff | !BtoS_ACK8_p & v93fc31;
assign v93f32a = BtoS_ACK0_p & v93f5d1 | !BtoS_ACK0_p & v90f16d;
assign v906b64 = BtoS_ACK8_p & v93fc15 | !BtoS_ACK8_p & !v93fdbc;
assign v909805 = jx1_p & v93f7bf | !jx1_p & v9058f3;
assign v93fa40 = StoB_REQ6_p & v93fb13 | !StoB_REQ6_p & v844f91;
assign v93fb2a = BtoS_ACK9_p & v8b5f61 | !BtoS_ACK9_p & v93f734;
assign v93f875 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v906642;
assign v89b116 = jx3_p & v9109e6 | !jx3_p & !v93fbaa;
assign v93f8b2 = BtoR_REQ0_p & v912fb2 | !BtoR_REQ0_p & v903b4e;
assign v909fd6 = BtoS_ACK9_p & v9043fc | !BtoS_ACK9_p & v93fe69;
assign v908ad9 = BtoS_ACK9_p & v93fd76 | !BtoS_ACK9_p & v908fb4;
assign v909bff = ENQ_p & v844f91 | !ENQ_p & v93fbcd;
assign v93fb1c = RtoB_ACK1_p & v93e751 | !RtoB_ACK1_p & v90e140;
assign v89f8ef = BtoS_ACK8_p & v93f768 | !BtoS_ACK8_p & v93dc29;
assign v8bbc51 = BtoS_ACK7_p & v9104ad | !BtoS_ACK7_p & !v90cf49;
assign v93e97c = BtoS_ACK0_p & v90f624 | !BtoS_ACK0_p & v93f805;
assign v93f812 = BtoS_ACK6_p & v9068b7 | !BtoS_ACK6_p & v85ea51;
assign v9132dc = jx2_p & v90caf3 | !jx2_p & !v903d5e;
assign v90949f = BtoS_ACK1_p & v93e356 | !BtoS_ACK1_p & v909f36;
assign v9112d5 = jx0_p & v844f9f | !jx0_p & !v9074ce;
assign v8baf9a = jx3_p & v93f78c | !jx3_p & !v90819e;
assign v910f4e = BtoS_ACK6_p & v910243 | !BtoS_ACK6_p & v844f91;
assign v9132b0 = StoB_REQ6_p & v863a78 | !StoB_REQ6_p & v844f91;
assign v93fe3d = BtoS_ACK6_p & v8b9b94 | !BtoS_ACK6_p & v93fb36;
assign v93f8b4 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & !v908106;
assign v93fcf2 = jx1_p & v910cee | !jx1_p & v9118f0;
assign v8f3868 = jx2_p & v9135db | !jx2_p & !v93fa80;
assign v93fdeb = StoB_REQ8_p & v93fa7e | !StoB_REQ8_p & v9049d0;
assign v93fa0d = StoB_REQ8_p & v9050e7 | !StoB_REQ8_p & v90e44c;
assign v93e829 = jx1_p & v911edb | !jx1_p & v930016;
assign v93fb5c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v906acc;
assign v9107ca = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v90d27b;
assign v90712d = BtoS_ACK8_p & v93e115 | !BtoS_ACK8_p & v93e9d8;
assign v93fcf9 = StoB_REQ9_p & v903c0d | !StoB_REQ9_p & v909c72;
assign v90d87f = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v905d66;
assign v93fc5a = BtoR_REQ0_p & v9111d3 | !BtoR_REQ0_p & v91007d;
assign v90fae7 = jx1_p & v93fc68 | !jx1_p & !v844f91;
assign v91229e = RtoB_ACK1_p & v90469d | !RtoB_ACK1_p & v90e774;
assign v90f0a1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90749b;
assign v906fbf = jx0_p & v93fb3e | !jx0_p & v913435;
assign v91334f = BtoS_ACK8_p & v93fb19 | !BtoS_ACK8_p & v93fa74;
assign v93db7f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93fd0d;
assign v87c4d9 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & !v844f91;
assign v93e162 = StoB_REQ8_p & v93ed2a | !StoB_REQ8_p & v90512d;
assign v93fd38 = StoB_REQ8_p & v93fc7b | !StoB_REQ8_p & v91143a;
assign v907299 = BtoS_ACK8_p & v93fdae | !BtoS_ACK8_p & v910101;
assign v8b9d84 = RtoB_ACK0_p & v90f304 | !RtoB_ACK0_p & v907a1b;
assign v904fcd = BtoS_ACK0_p & v9134df | !BtoS_ACK0_p & v93f69e;
assign v93f74f = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v904df8;
assign v909415 = jx0_p & v904f5c | !jx0_p & v9074ce;
assign v907110 = jx2_p & v9135db | !jx2_p & !v90cecd;
assign v9051ae = stateG7_1_p & v93e80c | !stateG7_1_p & v93fc2d;
assign v904357 = ENQ_p & v912477 | !ENQ_p & v91e95f;
assign v90e8f5 = BtoS_ACK8_p & v93fc04 | !BtoS_ACK8_p & v86345d;
assign v93f82b = BtoS_ACK1_p & v913348 | !BtoS_ACK1_p & v90a525;
assign v93f9b0 = jx0_p & v8f37ef | !jx0_p & v93f6f5;
assign v907200 = StoB_REQ9_p & v87f17f | !StoB_REQ9_p & !v844f91;
assign v90f304 = jx3_p & v93fa72 | !jx3_p & !v93f699;
assign v93fda6 = jx3_p & v90950c | !jx3_p & v903b83;
assign v93e926 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v93ed70;
assign v911946 = BtoS_ACK7_p & v844fa1 | !BtoS_ACK7_p & !v911fc7;
assign v907685 = RtoB_ACK0_p & v907bd4 | !RtoB_ACK0_p & v93fb21;
assign v93e369 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9d;
assign v90a348 = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & !v93fe46;
assign v910242 = jx3_p & v93f6db | !jx3_p & v8a1fe3;
assign v90df02 = StoB_REQ8_p & v87a1d0 | !StoB_REQ8_p & v93e948;
assign v93fdf1 = BtoS_ACK9_p & v912fad | !BtoS_ACK9_p & v910fe2;
assign v85eaa2 = stateG7_1_p & v8b9d84 | !stateG7_1_p & v906038;
assign v9135e7 = jx3_p & v93e7af | !jx3_p & v90523b;
assign v93fbd0 = jx1_p & v844f91 | !jx1_p & v909705;
assign v93f088 = BtoS_ACK8_p & v89e10d | !BtoS_ACK8_p & v93fd95;
assign v872e32 = BtoS_ACK2_p & v863a37 | !BtoS_ACK2_p & v93db3f;
assign v93f8d4 = EMPTY_p & v93f736 | !EMPTY_p & v93f9b8;
assign v90ebcd = StoB_REQ1_p & v93e926 | !StoB_REQ1_p & v93f6fd;
assign v863a2d = StoB_REQ8_p & v906915 | !StoB_REQ8_p & v93f795;
assign v907383 = jx1_p & v93ef01 | !jx1_p & v91026f;
assign v93e404 = StoB_REQ0_p & v93f7f5 | !StoB_REQ0_p & v85ea5f;
assign v93e288 = StoB_REQ7_p & v904ff8 | !StoB_REQ7_p & v910f4e;
assign v909b10 = jx2_p & v9042ba | !jx2_p & v909f68;
assign v9104ca = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91043e;
assign v93fbb9 = StoB_REQ1_p & v93def0 | !StoB_REQ1_p & v844f91;
assign v903d0b = BtoS_ACK7_p & v93f119 | !BtoS_ACK7_p & !v85eac9;
assign v91a6d5 = jx0_p & v90856f | !jx0_p & v9056ad;
assign v906209 = BtoS_ACK9_p & v8d195d | !BtoS_ACK9_p & v9117de;
assign v90ad9a = jx1_p & v8b9dff | !jx1_p & v90765f;
assign v93fcfc = jx0_p & v844f9b | !jx0_p & !v93fb3e;
assign v863afc = jx1_p & v904b4f | !jx1_p & !v90667d;
assign v90664c = StoB_REQ9_p & v9117e5 | !StoB_REQ9_p & v90dc0d;
assign v904f32 = BtoS_ACK6_p & v93e89f | !BtoS_ACK6_p & !v93f754;
assign v904a3b = DEQ_p & v8b9960 | !DEQ_p & v903e2f;
assign v93e470 = StoB_REQ7_p & v90441d | !StoB_REQ7_p & v90cbcc;
assign v90460e = jx0_p & v93ed91 | !jx0_p & v93f6e1;
assign v93f81e = jx1_p & v906461 | !jx1_p & !v844f91;
assign v93fd22 = StoB_REQ7_p & v909705 | !StoB_REQ7_p & v8f382e;
assign v906d83 = RtoB_ACK0_p & v903b56 | !RtoB_ACK0_p & v93f830;
assign v863add = jx3_p & v93fb57 | !jx3_p & v844f91;
assign v93fab8 = RtoB_ACK1_p & v93fdee | !RtoB_ACK1_p & v85eadc;
assign v90917f = jx0_p & v909157 | !jx0_p & v90932e;
assign v93fc10 = jx2_p & v903d90 | !jx2_p & !v93fa5b;
assign v90513b = DEQ_p & v9115ae | !DEQ_p & v91306c;
assign v93e148 = BtoS_ACK1_p & v90a59e | !BtoS_ACK1_p & v909c08;
assign v93fe0d = BtoS_ACK8_p & v90653d | !BtoS_ACK8_p & v93f627;
assign v93f9bc = BtoS_ACK7_p & v93f7d9 | !BtoS_ACK7_p & !v93fdb2;
assign v93eaa8 = BtoS_ACK1_p & v8bb868 | !BtoS_ACK1_p & v908c12;
assign v863abb = jx1_p & v93fc94 | !jx1_p & v844f91;
assign v9119f9 = jx1_p & v8b9ebe | !jx1_p & v8f22ce;
assign v93e23c = jx1_p & v93f768 | !jx1_p & v93fc5f;
assign v907965 = jx2_p & v90fc87 | !jx2_p & !v90a2df;
assign v93f074 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93ec47;
assign v90927a = BtoS_ACK8_p & v9074fa | !BtoS_ACK8_p & v90db9e;
assign v93f558 = jx1_p & v844f91 | !jx1_p & v9058f3;
assign v89fd8d = jx3_p & v93fdf1 | !jx3_p & !v905f24;
assign v90f9be = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v913561;
assign v87052e = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v93f9e8;
assign v91a6ea = jx2_p & v863abb | !jx2_p & !v844f91;
assign v8b9ce5 = BtoS_ACK8_p & v90451f | !BtoS_ACK8_p & !v90723b;
assign v9046a6 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v906acc = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v87c9bf;
assign v909043 = jx0_p & v93e648 | !jx0_p & v844f91;
assign v8b714e = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v93f83a;
assign v9101cc = jx1_p & v91ae94 | !jx1_p & v9060c1;
assign v93f8ab = StoB_REQ6_p & v909e9d | !StoB_REQ6_p & v93fe41;
assign v905d73 = jx0_p & v90ea74 | !jx0_p & !v90a0e8;
assign v93ec47 = jx1_p & v93ecc4 | !jx1_p & v844f91;
assign v93f8d3 = jx1_p & v844f91 | !jx1_p & v8b49f1;
assign v93fd3c = jx0_p & v90762a | !jx0_p & v90d879;
assign v905dc0 = EMPTY_p & v93f77b | !EMPTY_p & v93fa5d;
assign v93f8fa = BtoS_ACK7_p & v93ed2a | !BtoS_ACK7_p & v906541;
assign v93e896 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v911311;
assign v912d04 = BtoS_ACK6_p & v91aa51 | !BtoS_ACK6_p & v90a9c5;
assign v89fd94 = StoB_REQ8_p & v86fef2 | !StoB_REQ8_p & v89c580;
assign v911a72 = jx2_p & v909805 | !jx2_p & v844f91;
assign v908515 = BtoS_ACK8_p & v8b5f61 | !BtoS_ACK8_p & !v93f58c;
assign v85f2b0 = RtoB_ACK0_p & v93e301 | !RtoB_ACK0_p & v90539a;
assign v8f22a5 = StoB_REQ0_p & v9071c7 | !StoB_REQ0_p & v93f74f;
assign v904ba7 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v89f90b;
assign v9300af = StoB_REQ4_p & v844fbb | !StoB_REQ4_p & v904182;
assign v9134e2 = BtoS_ACK7_p & v907f25 | !BtoS_ACK7_p & v93e41f;
assign v93f714 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v93f70c;
assign v90decc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90e7d7;
assign v86c2d0 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v844f91;
assign v93e10c = jx2_p & v93f4cd | !jx2_p & !v93f75b;
assign v90526b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v93fbb9;
assign v906d77 = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & v93ebf5;
assign v91336b = RtoB_ACK1_p & v8f383c | !RtoB_ACK1_p & v908545;
assign v93fc09 = jx2_p & v93fe2d | !jx2_p & v910243;
assign v904a8a = BtoS_ACK9_p & v909e99 | !BtoS_ACK9_p & v8b9c3a;
assign v8a8f5e = jx1_p & v844f91 | !jx1_p & v93f9a4;
assign v844fa9 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v93fc98 = StoB_REQ8_p & v9071ed | !StoB_REQ8_p & v907633;
assign v93f2a4 = jx1_p & v93f63b | !jx1_p & v90ad75;
assign v93fb4a = BtoS_ACK9_p & v93e162 | !BtoS_ACK9_p & v93fd97;
assign v9097b1 = StoB_REQ0_p & v93f70c | !StoB_REQ0_p & v904e16;
assign v9124ae = jx2_p & v90e36f | !jx2_p & v93fa91;
assign v90df44 = jx2_p & v87c51f | !jx2_p & !v911090;
assign v863a00 = ENQ_p & v93f753 | !ENQ_p & v93f634;
assign v93f9dd = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v90decc;
assign v93f7bc = BtoS_ACK7_p & v907f25 | !BtoS_ACK7_p & v90921e;
assign v90a59b = BtoS_ACK8_p & v93f279 | !BtoS_ACK8_p & v93f88d;
assign v904074 = BtoS_ACK1_p & v906627 | !BtoS_ACK1_p & v907468;
assign v910710 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9093ec;
assign v93fa03 = BtoS_ACK9_p & v85ea96 | !BtoS_ACK9_p & v907ef2;
assign v93e655 = BtoS_ACK6_p & v90d22b | !BtoS_ACK6_p & v90ae6a;
assign v93eceb = BtoS_ACK0_p & v913348 | !BtoS_ACK0_p & v90a5b8;
assign v93f7ff = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fdb7;
assign v8b9f23 = jx2_p & v863a03 | !jx2_p & v93e919;
assign v90a5c0 = RtoB_ACK0_p & v907a4d | !RtoB_ACK0_p & v91a6e9;
assign v93fbfc = BtoS_ACK9_p & v91164f | !BtoS_ACK9_p & v904fbb;
assign v9089e7 = jx1_p & v90accf | !jx1_p & v93e51c;
assign v86fef2 = BtoS_ACK7_p & v9107aa | !BtoS_ACK7_p & !v904d39;
assign v904b09 = DEQ_p & v91aa2a | !DEQ_p & v90e333;
assign v87b2ea = BtoS_ACK6_p & v90ede1 | !BtoS_ACK6_p & v93f664;
assign v93fc4f = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & !v9119fd;
assign v904d40 = RtoB_ACK0_p & v93f746 | !RtoB_ACK0_p & v91a733;
assign v93f83c = jx3_p & v9073b6 | !jx3_p & v91155d;
assign jx2_n = !v8ebd2a;
assign v93fc97 = jx3_p & v844f91 | !jx3_p & !v89f894;
assign v907559 = BtoS_ACK9_p & v90a2bd | !BtoS_ACK9_p & v93fccd;
assign v904432 = jx0_p & v909e2c | !jx0_p & v93f0b0;
assign v9054a2 = jx1_p & v9105ed | !jx1_p & v909f04;
assign v93f5f6 = jx0_p & v844f91 | !jx0_p & v904de5;
assign v93f6f8 = BtoS_ACK8_p & v93f279 | !BtoS_ACK8_p & v910ebb;
assign v93fdb2 = jx2_p & v93f1c4 | !jx2_p & !v844f91;
assign v89f9da = StoB_REQ1_p & v903bb1 | !StoB_REQ1_p & v9103bc;
assign v9124bc = BtoS_ACK6_p & v93fb3e | !BtoS_ACK6_p & v9091b2;
assign v90a419 = DEQ_p & v93f8de | !DEQ_p & v90d9b7;
assign v93f9ad = StoB_REQ7_p & v910710 | !StoB_REQ7_p & v90496b;
assign v93fb2f = BtoS_ACK7_p & v93f869 | !BtoS_ACK7_p & !v89f97f;
assign v908636 = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v93ee1b;
assign v8810ad = StoB_REQ8_p & v8ee1a7 | !StoB_REQ8_p & v913342;
assign v93e773 = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v913a6f;
assign v90ed3d = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v90fe49;
assign v93faa4 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v903c65;
assign v90ad0a = BtoS_ACK8_p & v93f85d | !BtoS_ACK8_p & !v93fe49;
assign v93fc9f = jx1_p & v844f91 | !jx1_p & v90edb8;
assign v9131cb = BtoR_REQ0_p & v90d7d2 | !BtoR_REQ0_p & v908cff;
assign v910f6e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v9052de;
assign v9042fa = BtoS_ACK7_p & v910ee7 | !BtoS_ACK7_p & v910d81;
assign v93fb51 = jx3_p & v93f6da | !jx3_p & v908325;
assign v906c71 = BtoS_ACK2_p & v9076a8 | !BtoS_ACK2_p & v910b33;
assign v90a485 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v87052e;
assign v930016 = StoB_REQ7_p & v90d87f | !StoB_REQ7_p & v90d6fa;
assign v93e915 = BtoS_ACK8_p & v9095b9 | !BtoS_ACK8_p & v8cec7e;
assign v93f790 = BtoS_ACK9_p & v90a6ac | !BtoS_ACK9_p & v903c40;
assign v8f3826 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f8b1;
assign v93dab8 = jx2_p & v9135b9 | !jx2_p & v87f17d;
assign v91109f = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v907e36;
assign v87c566 = ENQ_p & v911a33 | !ENQ_p & v911a89;
assign v85e94c = jx2_p & v904fbf | !jx2_p & v93fe75;
assign v9040cd = StoB_REQ7_p & v90ebde | !StoB_REQ7_p & v90861d;
assign v9050e0 = jx0_p & v844f91 | !jx0_p & !v90eef9;
assign v911023 = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & v9068ce;
assign v908816 = StoB_REQ6_p & v908f32 | !StoB_REQ6_p & v912124;
assign v911760 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8b98bd;
assign v93fb27 = BtoS_ACK1_p & v906255 | !BtoS_ACK1_p & !v8a8f89;
assign v885188 = StoB_REQ9_p & v93fdc9 | !StoB_REQ9_p & v93fb33;
assign v844fcd = ENQ_p & v844f91 | !ENQ_p & !v844f91;
assign v9054b5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v93f70c;
assign v90456e = jx1_p & v8f22d1 | !jx1_p & !v93fe1f;
assign v90d2b7 = jx0_p & v905c01 | !jx0_p & !v93f6fc;
assign v93f6b2 = BtoS_ACK7_p & v90e893 | !BtoS_ACK7_p & v906131;
assign v90f5fc = StoB_REQ7_p & v910919 | !StoB_REQ7_p & v90d0fd;
assign v93e024 = jx1_p & v93e819 | !jx1_p & v93f739;
assign v9056f9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v90f309;
assign v93dac8 = jx0_p & v93f895 | !jx0_p & v90eef9;
assign v93ebf5 = BtoS_ACK7_p & v93f588 | !BtoS_ACK7_p & !v93fa08;
assign v8b989a = BtoS_ACK8_p & v9043e5 | !BtoS_ACK8_p & v89fe24;
assign v904b58 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v905396;
assign v908b06 = StoB_REQ8_p & v89e10d | !StoB_REQ8_p & v93f6ed;
assign v90813f = jx1_p & v9080a7 | !jx1_p & !v907b86;
assign v90d0b8 = StoB_REQ0_p & v909525 | !StoB_REQ0_p & v93fac0;
assign v85ea42 = StoB_REQ7_p & v93f7e8 | !StoB_REQ7_p & v93fbac;
assign v93fdea = BtoS_ACK6_p & v93f910 | !BtoS_ACK6_p & v8ebce4;
assign v910915 = jx3_p & v844f91 | !jx3_p & v907559;
assign v844fab = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844f91;
assign v90491c = StoB_REQ6_p & v90932e | !StoB_REQ6_p & v93f81c;
assign v910e6e = BtoS_ACK0_p & v93fb3b | !BtoS_ACK0_p & v91dd4f;
assign v912383 = BtoS_ACK0_p & v913561 | !BtoS_ACK0_p & v93ec6f;
assign v93fa17 = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v86c2d0;
assign v89f90b = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v909cb1;
assign v86d767 = jx2_p & v93f743 | !jx2_p & v90991f;
assign v91ddca = BtoS_ACK7_p & v9104ad | !BtoS_ACK7_p & !v93e8ab;
assign v91a9b9 = jx0_p & v8c737b | !jx0_p & v90414b;
assign v93fd59 = BtoS_ACK9_p & v907e3f | !BtoS_ACK9_p & v90d8f3;
assign v93f8a2 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v903e08;
assign v87a1f9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v909174;
assign v93f1cf = jx0_p & v844f9b | !jx0_p & !v905136;
assign v905d04 = BtoS_ACK6_p & v93fb08 | !BtoS_ACK6_p & v90f2ff;
assign v93e47b = jx2_p & v93f838 | !jx2_p & v90962d;
assign v905ffe = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fc22;
assign v889a9e = jx0_p & v9082e4 | !jx0_p & !v93fce2;
assign v90ea98 = RtoB_ACK0_p & v9049ac | !RtoB_ACK0_p & v90f629;
assign v93ec6f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90548c;
assign v93fcc9 = jx0_p & v8b9e82 | !jx0_p & !v906ae9;
assign v87c55f = StoB_REQ6_p & v9089bf | !StoB_REQ6_p & v9097b1;
assign v904878 = StoB_REQ8_p & v93fd86 | !StoB_REQ8_p & v90ae1b;
assign v93f6ce = StoB_REQ3_p & v904182 | !StoB_REQ3_p & !v844f91;
assign v90f38b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v91305d;
assign v90860a = jx0_p & v844f9f | !jx0_p & !v863a78;
assign v93f97f = jx0_p & v9115e3 | !jx0_p & v93e138;
assign v93dc87 = BtoS_ACK7_p & v9114c9 | !BtoS_ACK7_p & !v93edbf;
assign v911c01 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v93f865;
assign v844fb1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v93fd1c = StoB_REQ9_p & v9078a1 | !StoB_REQ9_p & v90aa3c;
assign v89c5bd = BtoS_ACK6_p & v93f63b | !BtoS_ACK6_p & v844f91;
assign v93fcb1 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93faed;
assign v906327 = StoB_REQ9_p & v91109f | !StoB_REQ9_p & v904901;
assign v903b7c = StoB_REQ8_p & v90722c | !StoB_REQ8_p & v910b7a;
assign v9077f6 = stateG7_1_p & v907292 | !stateG7_1_p & v9060e9;
assign v912178 = StoB_REQ8_p & v904ab4 | !StoB_REQ8_p & v93f7bc;
assign v93f70f = RtoB_ACK0_p & v90dcca | !RtoB_ACK0_p & v909dec;
assign v93f6df = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90eda0;
assign v86f4a3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v9095bf;
assign v9096f7 = BtoS_ACK0_p & v93f85e | !BtoS_ACK0_p & v89fdce;
assign v904779 = jx1_p & v93fd9e | !jx1_p & v93fcd4;
assign v8a8fac = StoB_REQ2_p & v905702 | !StoB_REQ2_p & !v844f91;
assign v911bb8 = StoB_REQ9_p & v90e159 | !StoB_REQ9_p & v904da8;
assign v93fe68 = StoB_REQ7_p & v9130af | !StoB_REQ7_p & v863477;
assign v90f478 = BtoS_ACK9_p & v93f074 | !BtoS_ACK9_p & v884fc2;
assign v9091b4 = jx1_p & v88d7c9 | !jx1_p & v91315c;
assign v9057c9 = jx1_p & v9056d9 | !jx1_p & v844f91;
assign v90edb9 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v91262e;
assign v8b9c3e = BtoS_ACK2_p & v87a21f | !BtoS_ACK2_p & v93ea28;
assign v9084f4 = jx1_p & v93e065 | !jx1_p & v909c15;
assign v93e9c8 = RtoB_ACK1_p & v87c9b3 | !RtoB_ACK1_p & v90738b;
assign v873bc3 = StoB_REQ9_p & v93fc35 | !StoB_REQ9_p & v93f9fa;
assign v905487 = BtoS_ACK8_p & v93ed2a | !BtoS_ACK8_p & v93f4e9;
assign v93006d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v906042;
assign v913a54 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90aa64;
assign v907bb9 = ENQ_p & v844fc3 | !ENQ_p & !v90ed80;
assign v93f68b = jx0_p & v844f91 | !jx0_p & v904f5c;
assign v90dff3 = jx3_p & v844f91 | !jx3_p & v93ed58;
assign v93f869 = jx2_p & v93ed6a | !jx2_p & !v90cbec;
assign v907e33 = ENQ_p & v911b74 | !ENQ_p & v93fbcd;
assign v912d1a = ENQ_p & v90a774 | !ENQ_p & !v93fd4a;
assign v90762a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93f7af;
assign v9084d0 = BtoS_ACK9_p & v93f979 | !BtoS_ACK9_p & v93ed1c;
assign v93e3dd = DEQ_p & v8b9960 | !DEQ_p & v8b9cc5;
assign v93fd96 = BtoS_ACK8_p & v90529c | !BtoS_ACK8_p & v93f444;
assign v93fcd6 = StoB_REQ8_p & v907adb | !StoB_REQ8_p & v909fb2;
assign v910c5b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9085ac;
assign v884481 = jx0_p & v844f9b | !jx0_p & v844f99;
assign v93eef4 = stateG7_1_p & v844f91 | !stateG7_1_p & v90d651;
assign v93f7fb = BtoS_ACK6_p & v9047e4 | !BtoS_ACK6_p & v93f722;
assign v9082a5 = BtoS_ACK7_p & v905ff9 | !BtoS_ACK7_p & v90dd28;
assign v93fe5c = jx0_p & v90f5b6 | !jx0_p & v844f91;
assign v90a20a = StoB_REQ0_p & v90a902 | !StoB_REQ0_p & v93f02c;
assign v90acaa = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90eed2;
assign v90dd1f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v9075db;
assign v903d5e = jx1_p & v910243 | !jx1_p & v93f7f1;
assign v93f689 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v9071c7;
assign v908fd6 = StoB_REQ9_p & v9103e4 | !StoB_REQ9_p & v879731;
assign v93eda5 = jx1_p & v87bae8 | !jx1_p & !v844f91;
assign v908a35 = BtoS_ACK7_p & v8b9ee2 | !BtoS_ACK7_p & v8f3868;
assign v8b9ec9 = BtoS_ACK6_p & v93fb3e | !BtoS_ACK6_p & v93f8ab;
assign v93fae2 = StoB_REQ8_p & v9071ed | !StoB_REQ8_p & v90980a;
assign v93f83f = StoB_REQ6_p & v909107 | !StoB_REQ6_p & v93fac9;
assign v93f7ae = ENQ_p & v93e704 | !ENQ_p & v90a602;
assign v89f916 = StoB_REQ7_p & v903e94 | !StoB_REQ7_p & v93fe31;
assign v90a074 = DEQ_p & v91aa2a | !DEQ_p & v93fd44;
assign v8b9d37 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8ebd0e;
assign v93f7de = StoB_REQ7_p & v903e94 | !StoB_REQ7_p & v9112d5;
assign v90f9ed = BtoS_ACK9_p & v93e136 | !BtoS_ACK9_p & v90aca4;
assign v93f2dc = jx0_p & v910fd2 | !jx0_p & !v93fd21;
assign v93fdcc = BtoS_ACK9_p & v844fa5 | !BtoS_ACK9_p & !v911452;
assign v85e7ba = jx0_p & v93fa3b | !jx0_p & !v930109;
assign v8b9ee1 = jx1_p & v844f91 | !jx1_p & !v93f6cc;
assign v909a21 = jx2_p & v90f9fc | !jx2_p & v8f60f9;
assign v9108ff = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9077b1;
assign v93fc3e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v90606d;
assign v9073b6 = BtoS_ACK9_p & v904e48 | !BtoS_ACK9_p & v9049e4;
assign v93fdde = StoB_REQ0_p & v844f97 | !StoB_REQ0_p & v90810f;
assign v90e856 = BtoS_ACK6_p & v90cc30 | !BtoS_ACK6_p & !v93f895;
assign v93f955 = jx2_p & v9080c5 | !jx2_p & !v844f91;
assign v93fbea = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v93f050;
assign v90dcf6 = BtoS_ACK7_p & v906ec1 | !BtoS_ACK7_p & v909c74;
assign v90add3 = jx0_p & v90f2de | !jx0_p & v9102bf;
assign v908c12 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v9300c0;
assign v93f8d2 = StoB_REQ6_p & v9081b9 | !StoB_REQ6_p & v911b83;
assign v904200 = BtoS_ACK6_p & v910243 | !BtoS_ACK6_p & v93f7ea;
assign v93fe6a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87a2ad;
assign v918724 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v93fdb8;
assign v90fa80 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v90968f;
assign v93ec50 = jx0_p & v93e402 | !jx0_p & !v90ee6d;
assign v93fc4c = BtoS_ACK6_p & v9100ff | !BtoS_ACK6_p & v93f895;
assign v8880f2 = StoB_REQ9_p & v86d7d1 | !StoB_REQ9_p & v8b989a;
assign v90d5b3 = EMPTY_p & v909dec | !EMPTY_p & v87c517;
assign v93f6bc = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v9052de;
assign v909e9d = BtoS_ACK0_p & v93f5d1 | !BtoS_ACK0_p & v904d38;
assign v905322 = BtoR_REQ0_p & v90f33b | !BtoR_REQ0_p & !v906570;
assign v8f22ca = RtoB_ACK0_p & v90d057 | !RtoB_ACK0_p & v93fb11;
assign v906c66 = StoB_REQ7_p & v9058f3 | !StoB_REQ7_p & v9085fc;
assign v9106af = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v93fa49;
assign v93f7c8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v87179f;
assign v93f78f = StoB_REQ8_p & v8ee1bc | !StoB_REQ8_p & v905a9e;
assign v93f8e2 = jx1_p & v89f98c | !jx1_p & !v903e94;
assign v910fcd = ENQ_p & v93eda4 | !ENQ_p & v93fa96;
assign v93fbdc = ENQ_p & v90fe92 | !ENQ_p & v93fbcd;
assign v913592 = jx1_p & v90468e | !jx1_p & v844f91;
assign v8b9c50 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v93f7f7;
assign v90e546 = stateG12_p & v93fa72 | !stateG12_p & v93e6fe;
assign v9120f4 = StoB_REQ1_p & v906642 | !StoB_REQ1_p & v93f1c8;
assign v90859f = RtoB_ACK1_p & v93e281 | !RtoB_ACK1_p & v910c29;
assign v9087d1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9087b1;
assign v8b496d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v93f2da;
assign v93ec28 = BtoS_ACK7_p & v93fbe4 | !BtoS_ACK7_p & v93df10;
assign v93fa75 = RtoB_ACK0_p & v907a32 | !RtoB_ACK0_p & v93f91c;
assign v906491 = BtoS_ACK6_p & v90df7f | !BtoS_ACK6_p & v844f91;
assign v93fa84 = jx2_p & v858fc9 | !jx2_p & !v93f9f3;
assign v903b91 = StoB_REQ9_p & v90f9f3 | !StoB_REQ9_p & v90a59b;
assign v93e356 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v91305b;
assign BtoS_ACK9_n = v89b1a4;
assign v93f29e = StoB_REQ6_p & v93e77a | !StoB_REQ6_p & v86ccf1;
assign v9056bd = jx0_p & v90eef9 | !jx0_p & !v90cc30;
assign v91305b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v93fd2b;
assign v90d5c7 = BtoS_ACK7_p & v9187aa | !BtoS_ACK7_p & v93e23c;
assign v904c99 = jx1_p & v844f91 | !jx1_p & v9041e6;
assign v907b58 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v93f7bb;
assign v9052ce = BtoS_ACK6_p & v90630d | !BtoS_ACK6_p & v93dfc7;
assign v9058c2 = StoB_REQ9_p & v93f8b5 | !StoB_REQ9_p & v89f8a9;
assign v909a7c = BtoS_ACK8_p & v911b48 | !BtoS_ACK8_p & !v93efae;
assign v8a8fb1 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v90f624;
assign v904ede = jx2_p & v93fe66 | !jx2_p & v844f91;
assign v9132f8 = BtoS_ACK8_p & v93fe3f | !BtoS_ACK8_p & v903b0f;
assign v90e251 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v91162e;
assign v9117e5 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93fcc8;
assign v93db04 = RtoB_ACK1_p & v8b9f34 | !RtoB_ACK1_p & v93fa47;
assign v93f8c3 = BtoS_ACK1_p & v8bb868 | !BtoS_ACK1_p & v91100a;
assign v93fbff = BtoS_ACK1_p & v913619 | !BtoS_ACK1_p & v90f8e7;
assign v93fe61 = EMPTY_p & v87c566 | !EMPTY_p & v90d5c3;
assign v93e037 = EMPTY_p & v90567d | !EMPTY_p & v9056e2;
assign v9046d6 = BtoS_ACK6_p & v8a9222 | !BtoS_ACK6_p & v93fce1;
assign v9130c5 = stateG7_1_p & v93f82a | !stateG7_1_p & v8b99a1;
assign v93fcf1 = BtoS_ACK6_p & v93f91d | !BtoS_ACK6_p & v844f91;
assign v912f3d = RtoB_ACK0_p & v93f6fa | !RtoB_ACK0_p & v9112d1;
assign v93fb19 = jx2_p & v93f694 | !jx2_p & !v844f91;
assign v9122e7 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v911509;
assign v93fa66 = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & !v90e1dd;
assign v90fca6 = jx1_p & v869aeb | !jx1_p & !v90ec5d;
assign v93fcba = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93faf1;
assign v884dd3 = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & v90a08d;
assign v93f68a = jx1_p & v93f0a3 | !jx1_p & v906256;
assign v93f462 = StoB_REQ1_p & v93e9cc | !StoB_REQ1_p & v90caeb;
assign v9099f2 = RtoB_ACK0_p & v886fce | !RtoB_ACK0_p & v93f6fa;
assign v908429 = BtoS_ACK9_p & v90dd2f | !BtoS_ACK9_p & v903d1e;
assign v911435 = EMPTY_p & v9082e6 | !EMPTY_p & v908ffc;
assign v9124b8 = BtoS_ACK6_p & v90df7f | !BtoS_ACK6_p & v904f64;
assign v910237 = jx3_p & v905511 | !jx3_p & v93f912;
assign v93e51c = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v93f901;
assign v844f9d = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v844f91;
assign v9057c1 = jx1_p & v93fc94 | !jx1_p & !v91aa51;
assign v9043fc = StoB_REQ8_p & v93fc04 | !StoB_REQ8_p & v93fb93;
assign v9103e4 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v910c5b;
assign v8ebd28 = StoB_REQ1_p & v872e32 | !StoB_REQ1_p & v906037;
assign v907c69 = jx3_p & v93f751 | !jx3_p & v93f753;
assign v93fb64 = BtoS_ACK0_p & v90873f | !BtoS_ACK0_p & v90acaa;
assign v910081 = StoB_REQ6_p & v93f888 | !StoB_REQ6_p & v93fbd7;
assign v93f9e8 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v9099e3;
assign v905077 = jx3_p & v91aa04 | !jx3_p & !v90a097;
assign v907684 = jx1_p & v90eef9 | !jx1_p & v90f5fc;
assign v904f0d = jx3_p & v93fcfe | !jx3_p & v93f89f;
assign v90946a = jx0_p & v90f5b6 | !jx0_p & !v90a485;
assign v8f382c = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v93fe2b;
assign v90871b = ENQ_p & v904f0d | !ENQ_p & v844f91;
assign v93f7ac = StoB_REQ7_p & v912fed | !StoB_REQ7_p & v9053de;
assign v906ff5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v92ffb9;
assign v93f75e = DEQ_p & v93f959 | !DEQ_p & v909dec;
assign v93facc = jx3_p & v93f78c | !jx3_p & !v9101c0;
assign v93fdb0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93f69e;
assign v93fa5d = DEQ_p & v90df61 | !DEQ_p & v93f899;
assign v90dcfa = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v90d42a;
assign v88de63 = StoB_REQ6_p & v909107 | !StoB_REQ6_p & v9100f8;
assign v911edb = StoB_REQ7_p & v93ef5c | !StoB_REQ7_p & !v905a80;
assign v93faeb = BtoS_ACK0_p & v90f624 | !BtoS_ACK0_p & v93e9ce;
assign v9080b4 = BtoS_ACK8_p & v8b9dff | !BtoS_ACK8_p & v93f7a8;
assign v904e13 = StoB_REQ9_p & v90e9f7 | !StoB_REQ9_p & v906b07;
assign v9091e3 = BtoS_ACK6_p & v9050a5 | !BtoS_ACK6_p & v90a3f6;
assign v90dd2f = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93f8f0;
assign v93fbe1 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v93db7f;
assign v906642 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f99;
assign v911b43 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v89f840;
assign v93e0fb = StoB_REQ9_p & v90fbfe | !StoB_REQ9_p & v93fb6e;
assign v907a13 = BtoS_ACK0_p & v90fc92 | !BtoS_ACK0_p & v93daaf;
assign v93fc8e = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v90611f;
assign v910c50 = StoB_REQ7_p & v93fc2b | !StoB_REQ7_p & v93f3a8;
assign v93fba0 = EMPTY_p & v93f736 | !EMPTY_p & v90e027;
assign v90f88e = BtoS_ACK0_p & v93f6bc | !BtoS_ACK0_p & v906a51;
assign v910e66 = jx2_p & v910e84 | !jx2_p & v93fe75;
assign v909bdf = ENQ_p & v91a6d3 | !ENQ_p & !v93ed15;
assign v93f7d3 = StoB_REQ9_p & v9110a9 | !StoB_REQ9_p & v93f7dd;
assign v93f6cb = jx2_p & v90a214 | !jx2_p & v911c82;
assign v93f917 = jx3_p & v90ba31 | !jx3_p & !v844f91;
assign v90575e = DEQ_p & v93e3f1 | !DEQ_p & v90926e;
assign v90980a = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8ee172;
assign v93ecc4 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v863b25;
assign v91a71d = DEQ_p & v8b9c4f | !DEQ_p & v90ad6f;
assign v9049d0 = BtoS_ACK7_p & v89f983 | !BtoS_ACK7_p & v87c21e;
assign v93f913 = BtoS_ACK7_p & v907965 | !BtoS_ACK7_p & v8b9e4f;
assign v9054c9 = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & !v904757;
assign v908f32 = BtoS_ACK0_p & v86e433 | !BtoS_ACK0_p & v904654;
assign v89f80d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f692;
assign v9045fa = BtoS_ACK6_p & v90ede1 | !BtoS_ACK6_p & !v90752a;
assign v9062d9 = StoB_REQ1_p & v913348 | !StoB_REQ1_p & v8bb868;
assign v93fac1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9104ca;
assign v905168 = jx2_p & v863a03 | !jx2_p & v90eaad;
assign v908073 = jx2_p & v93fa16 | !jx2_p & !v93f2a4;
assign v908df3 = FULL_p & v9082be | !FULL_p & v93f19b;
assign v90a6d8 = BtoS_ACK6_p & v90a926 | !BtoS_ACK6_p & v93f69b;
assign v9050ba = StoB_REQ9_p & v89e10d | !StoB_REQ9_p & v844f91;
assign v905397 = ENQ_p & v844f91 | !ENQ_p & v90d629;
assign v90d250 = StoB_REQ9_p & v908fe9 | !StoB_REQ9_p & v93fc4f;
assign v90451f = jx2_p & v90423b | !jx2_p & v90cbec;
assign v93fa7b = BtoS_ACK7_p & v90408b | !BtoS_ACK7_p & v85ead8;
assign v91214b = EMPTY_p & v9076cf | !EMPTY_p & v93e4b4;
assign v904988 = jx1_p & v87a20b | !jx1_p & v93f84d;
assign v909b02 = BtoS_ACK7_p & v906c2f | !BtoS_ACK7_p & v93f6cb;
assign v90ed7e = ENQ_p & v844fc3 | !ENQ_p & !v93ef38;
assign v93fb8d = jx1_p & v90fb54 | !jx1_p & !v844f91;
assign v93fd51 = BtoS_ACK6_p & v910f82 | !BtoS_ACK6_p & v9070e2;
assign v93dc15 = jx1_p & v93f0a9 | !jx1_p & v90a876;
assign v90ed80 = jx3_p & v93f937 | !jx3_p & v90536f;
assign v9062ae = StoB_REQ8_p & v93fe4b | !StoB_REQ8_p & v93fd04;
assign v903d0c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90893a;
assign v93fb8a = EMPTY_p & v911b68 | !EMPTY_p & v904614;
assign v93f77a = BtoS_ACK8_p & v89f988 | !BtoS_ACK8_p & v90f7ce;
assign v90611f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v90fe49;
assign v906623 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v909637;
assign v905d0a = BtoS_ACK9_p & v90dec9 | !BtoS_ACK9_p & v93fbea;
assign v9055bd = BtoS_ACK6_p & v884481 | !BtoS_ACK6_p & v91023b;
assign v93fd18 = BtoS_ACK8_p & v90a4da | !BtoS_ACK8_p & v904878;
assign v87179f = BtoS_ACK6_p & v905971 | !BtoS_ACK6_p & v93fd9a;
assign v93debb = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v90432c;
assign v906d92 = stateG7_1_p & v90d651 | !stateG7_1_p & v844f91;
assign v90aaca = BtoS_ACK0_p & v910825 | !BtoS_ACK0_p & v9073c3;
assign v911b68 = ENQ_p & v93e704 | !ENQ_p & v90f819;
assign v93f6ac = StoB_REQ7_p & v87a20d | !StoB_REQ7_p & v89f938;
assign v93fdd7 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93f765;
assign v93fb5d = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v93fbb6;
assign v91247f = jx2_p & v904b51 | !jx2_p & v93faa7;
assign v9300da = jx0_p & v90ea74 | !jx0_p & !v904521;
assign v90e333 = ENQ_p & v911a33 | !ENQ_p & v904ba3;
assign v90e4ec = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v908df7;
assign v905da3 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93e48f;
assign v909c15 = StoB_REQ7_p & v93f9a4 | !StoB_REQ7_p & v93e45c;
assign v90931a = StoB_REQ8_p & v93e296 | !StoB_REQ8_p & v910c4e;
assign v93f492 = jx3_p & v910840 | !jx3_p & v909312;
assign v911c73 = jx0_p & v90515d | !jx0_p & v844f91;
assign v904b45 = jx1_p & v90515d | !jx1_p & v904809;
assign v93ef46 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v90729a;
assign v90a5c1 = jx1_p & v906fbf | !jx1_p & v90460e;
assign v93f82a = DEQ_p & v93fd1b | !DEQ_p & !v904f93;
assign v86345f = jx3_p & v93f110 | !jx3_p & v90a4b7;
assign v93fe34 = BtoS_ACK0_p & v90a5ef | !BtoS_ACK0_p & v872746;
assign v9083f0 = StoB_REQ8_p & v90722c | !StoB_REQ8_p & v9132dc;
assign v911b50 = jx0_p & v844f91 | !jx0_p & v93f8bb;
assign v93ec0d = BtoS_ACK1_p & v90a59e | !BtoS_ACK1_p & v93fbf8;
assign v9124a6 = StoB_REQ0_p & v93fc1a | !StoB_REQ0_p & v93fc38;
assign v90cbf6 = jx0_p & v93fc0a | !jx0_p & v8d37c1;
assign v93fa9d = BtoS_ACK6_p & v93f91d | !BtoS_ACK6_p & v93fbb3;
assign v8f383a = RtoB_ACK1_p & v9092a8 | !RtoB_ACK1_p & v93fcb2;
assign v90dc9c = jx1_p & v844f91 | !jx1_p & !v93fcc9;
assign v93fd1d = StoB_REQ7_p & v910710 | !StoB_REQ7_p & !v93fbe5;
assign v90f0c5 = RtoB_ACK0_p & v904fee | !RtoB_ACK0_p & v904c4f;
assign v9098e3 = BtoS_ACK7_p & v93e47b | !BtoS_ACK7_p & v910644;
assign v903df5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9062d9;
assign v93f6f5 = StoB_REQ6_p & v93f7c4 | !StoB_REQ6_p & v9133d2;
assign v93f9cb = ENQ_p & v908325 | !ENQ_p & v90f2da;
assign v91a6dc = EMPTY_p & v910525 | !EMPTY_p & v9102bb;
assign v90d9b7 = RtoB_ACK0_p & v908751 | !RtoB_ACK0_p & v93dfb4;
assign v904da8 = BtoS_ACK8_p & v93fe3f | !BtoS_ACK8_p & v93f6a6;
assign v93f87c = BtoS_ACK9_p & v93e3a1 | !BtoS_ACK9_p & v911bb8;
assign v93fc1a = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v93fc28;
assign v906b07 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & v913265;
assign v9065d3 = jx2_p & v911fe3 | !jx2_p & v905329;
assign v85f268 = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v88036c;
assign v93faf0 = BtoS_ACK9_p & v9056a4 | !BtoS_ACK9_p & v903b91;
assign v904b9e = BtoS_ACK9_p & v90f947 | !BtoS_ACK9_p & v8d37d4;
assign v93e681 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93fc02;
assign v904bcb = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v90d972;
assign v90508f = BtoS_ACK0_p & v93fb3b | !BtoS_ACK0_p & v91a6f7;
assign v93fc4e = StoB_REQ0_p & v907c8c | !StoB_REQ0_p & v844f91;
assign v904b51 = jx1_p & v93f7c8 | !jx1_p & v90fc6d;
assign v8ee1d1 = jx1_p & v844f91 | !jx1_p & v908546;
assign v87c4fa = BtoS_ACK6_p & v844f95 | !BtoS_ACK6_p & !v904de5;
assign v8a9205 = jx0_p & v90cfa8 | !jx0_p & !v905619;
assign v904d56 = FULL_p & v904c4f | !FULL_p & v904fee;
assign v93fdc0 = stateG12_p & v844fc3 | !stateG12_p & !v90f4dd;
assign v907d8b = jx0_p & v9081b9 | !jx0_p & v844f91;
assign v90ded0 = jx1_p & v8b9b9f | !jx1_p & !v844f91;
assign v87c54e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90d880;
assign v93e4c1 = StoB_REQ7_p & v93e655 | !StoB_REQ7_p & v844f91;
assign v9087d2 = jx1_p & v9091e3 | !jx1_p & v844f91;
assign v87c503 = jx1_p & v906495 | !jx1_p & v9064b4;
assign v910243 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910f6e;
assign v93f797 = StoB_REQ1_p & v905660 | !StoB_REQ1_p & v93fb5a;
assign v93fce8 = BtoS_ACK6_p & v90a6d6 | !BtoS_ACK6_p & v93fdc4;
assign v888002 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v903d21;
assign v90e4f2 = BtoS_ACK7_p & v9104ad | !BtoS_ACK7_p & !v93f787;
assign v905ed9 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v93faa4;
assign v90fe92 = jx3_p & v87f17f | !jx3_p & !v844f91;
assign v8c7343 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v93e356;
assign v89b1a0 = jx1_p & v93f293 | !jx1_p & v93f6c6;
assign v8f3874 = BtoS_ACK7_p & v8633c3 | !BtoS_ACK7_p & !v93f80d;
assign v87c4d2 = BtoS_ACK7_p & v90541b | !BtoS_ACK7_p & !v93f9bb;
assign v9085b3 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v93fde4;
assign v909d71 = jx2_p & v9101cc | !jx2_p & v89b1a0;
assign v93f899 = ENQ_p & v93eed6 | !ENQ_p & v93fcbd;
assign v93f19b = ENQ_p & v93f753 | !ENQ_p & v93e189;
assign v91262e = BtoS_ACK7_p & v93ea4f | !BtoS_ACK7_p & v93f02f;
assign v8b9c00 = stateG12_p & v90a9cc | !stateG12_p & v93e4f9;
assign v91042d = jx1_p & v8b9dff | !jx1_p & v93f7bf;
assign v907ef2 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v8b9d25;
assign v905b81 = ENQ_p & v93f89f | !ENQ_p & v93fe44;
assign v882135 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90e304;
assign v93e903 = BtoS_ACK6_p & v90860a | !BtoS_ACK6_p & v90e95b;
assign v9102f4 = BtoS_ACK6_p & v8a9289 | !BtoS_ACK6_p & v90e32f;
assign v9109dc = jx2_p & v93fc9f | !jx2_p & !v93fa70;
assign v93f535 = jx1_p & v913332 | !jx1_p & v89b100;
assign v90a1c0 = BtoR_REQ0_p & v9094f2 | !BtoR_REQ0_p & v910b22;
assign v904f14 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v89f79e;
assign v93fe06 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v9109ee;
assign v93fa1b = jx0_p & v90515d | !jx0_p & v8a927b;
assign v907c85 = BtoS_ACK7_p & v93dbf1 | !BtoS_ACK7_p & v93fae3;
assign v903eef = BtoS_ACK8_p & v93f73d | !BtoS_ACK8_p & v90dab9;
assign jx3_n = !v9384b0;
assign v93eaca = jx1_p & v93e7d1 | !jx1_p & v93fa86;
assign v90927b = jx1_p & v844f91 | !jx1_p & v9122e7;
assign v87ca35 = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v89e10d;
assign v904ee9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f91d;
assign v93e86e = jx0_p & v90d4cc | !jx0_p & v89f9bc;
assign v93fbfe = jx2_p & v93fe55 | !jx2_p & v90f1ab;
assign v909be8 = BtoS_ACK9_p & v9083f0 | !BtoS_ACK9_p & v885188;
assign v903f58 = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v90468f;
assign v90798e = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & !v9126bb;
assign v87a28e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93fcf1;
assign v93e9d1 = BtoS_ACK0_p & v93e2de | !BtoS_ACK0_p & v8b9e17;
assign v908fe9 = BtoS_ACK8_p & v90a6ac | !BtoS_ACK8_p & !v90d866;
assign v85eaed = StoB_REQ2_p & v93fdf7 | !StoB_REQ2_p & v90fc5f;
assign v93fc34 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v90712c;
assign v9043ec = BtoS_ACK6_p & v910f82 | !BtoS_ACK6_p & v909043;
assign v8b9c1e = StoB_REQ7_p & v93f910 | !StoB_REQ7_p & v93fcfc;
assign v93fd4e = jx0_p & v93005b | !jx0_p & v844f91;
assign v93fbe5 = BtoS_ACK6_p & v87f17d | !BtoS_ACK6_p & v93fc68;
assign v903d12 = stateG7_1_p & v906226 | !stateG7_1_p & v93fe47;
assign v90e906 = EMPTY_p & v90ace9 | !EMPTY_p & v93f75e;
assign v905dd8 = BtoS_ACK6_p & v93f910 | !BtoS_ACK6_p & v87f17d;
assign v90d4cc = BtoS_ACK0_p & v86c2d0 | !BtoS_ACK0_p & v907840;
assign v8ee17f = jx0_p & v906623 | !jx0_p & v8d37c1;
assign v906d4c = jx1_p & v90879a | !jx1_p & !v844f91;
assign v93def0 = BtoS_ACK2_p & v9123a2 | !BtoS_ACK2_p & v870fb9;
assign v90a7ea = StoB_REQ7_p & v903f58 | !StoB_REQ7_p & v8b9d5d;
assign v90df61 = RtoB_ACK0_p & v8b9c4f | !RtoB_ACK0_p & v90567c;
assign v8f2274 = jx3_p & v93fde9 | !jx3_p & v911a33;
assign v93edc8 = BtoS_ACK0_p & v90deff | !BtoS_ACK0_p & v906717;
assign v911c82 = jx1_p & v93f92c | !jx1_p & v908fb8;
assign v87a20b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93eb70;
assign v8a8fa0 = jx0_p & v93f83f | !jx0_p & !v904736;
assign v9119f8 = StoB_REQ9_p & v909e90 | !StoB_REQ9_p & v93fc0b;
assign v904b77 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v90fb89;
assign v93fa36 = RtoB_ACK0_p & v89f966 | !RtoB_ACK0_p & v91093d;
assign v93f743 = jx1_p & v93f28c | !jx1_p & v9109e5;
assign v906c0f = jx3_p & v844f91 | !jx3_p & v93f708;
assign v90fb5d = jx0_p & v844f9f | !jx0_p & !v844f9d;
assign v9110fe = jx3_p & v844f91 | !jx3_p & v903db7;
assign v905467 = BtoS_ACK7_p & v907684 | !BtoS_ACK7_p & v8b9eca;
assign v904f88 = StoB_REQ7_p & v93f8a6 | !StoB_REQ7_p & v93f307;
assign v93f3a8 = BtoS_ACK6_p & v910243 | !BtoS_ACK6_p & v904dd8;
assign v93f7b9 = ENQ_p & v93f15e | !ENQ_p & v9054a8;
assign v93fe55 = jx1_p & v869aeb | !jx1_p & !v90441d;
assign v90a4bf = StoB_REQ8_p & v93f8fa | !StoB_REQ8_p & v909b02;
assign v90e770 = EMPTY_p & v904357 | !EMPTY_p & !v93fc45;
assign v93e137 = BtoS_ACK9_p & v912fad | !BtoS_ACK9_p & v93f8b4;
assign v93fdb7 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v91aa52;
assign v904115 = StoB_REQ8_p & v911a00 | !StoB_REQ8_p & v8b9e60;
assign v90824f = jx1_p & v90e25e | !jx1_p & !v905de8;
assign v909637 = BtoS_ACK0_p & v90855a | !BtoS_ACK0_p & !v9062b5;
assign v90d0f9 = BtoS_ACK6_p & v93fcfc | !BtoS_ACK6_p & v91a9e1;
assign v9132d2 = jx0_p & v844f91 | !jx0_p & v93f6fc;
assign v90dd67 = ENQ_p & v93f15e | !ENQ_p & v93fc53;
assign v907f0b = jx2_p & v90cbfc | !jx2_p & !v93f6bf;
assign v93f8b1 = BtoS_ACK6_p & v89f84e | !BtoS_ACK6_p & v93f51c;
assign v910644 = jx2_p & v87a1f0 | !jx2_p & v93e13e;
assign v91066d = BtoS_ACK9_p & v9044c3 | !BtoS_ACK9_p & v93fce6;
assign v93f811 = StoB_REQ7_p & v9043f4 | !StoB_REQ7_p & v93f28b;
assign v93fb26 = BtoS_ACK9_p & v93e85e | !BtoS_ACK9_p & v93f6ad;
assign v90d634 = jx1_p & v93f766 | !jx1_p & v90f1b9;
assign v93e5d4 = StoB_REQ9_p & v911cba | !StoB_REQ9_p & v85eb17;
assign v90a07b = ENQ_p & v93fb51 | !ENQ_p & v90f2da;
assign v904f5c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v904fcd;
assign v909357 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v908574;
assign v8839a7 = BtoS_ACK6_p & v909f4c | !BtoS_ACK6_p & !v93f941;
assign v907122 = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & v93f5c0;
assign v90a334 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93f345;
assign v90f500 = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v93f81b;
assign v906b57 = jx1_p & v93ecc4 | !jx1_p & v9124cb;
assign v908083 = jx0_p & v9082e4 | !jx0_p & !v93fa56;
assign v93fc27 = StoB_REQ0_p & v906642 | !StoB_REQ0_p & !v844f91;
assign v90cc7a = BtoS_ACK6_p & v93f90a | !BtoS_ACK6_p & v93f782;
assign v91091b = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v93effa;
assign v8b9dfa = BtoS_ACK3_p & v91058e | !BtoS_ACK3_p & v911b78;
assign v9134c0 = StoB_REQ1_p & v904e53 | !StoB_REQ1_p & v906bf5;
assign v93f687 = jx1_p & v910710 | !jx1_p & v905252;
assign v90df7f = jx0_p & v93ed00 | !jx0_p & v93fd3d;
assign v910543 = jx3_p & v904b7f | !jx3_p & v93fb4a;
assign v90fe7e = jx3_p & v8b9c00 | !jx3_p & v844f91;
assign v909666 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v908096;
assign v91aa06 = BtoS_ACK6_p & v9058f3 | !BtoS_ACK6_p & v93f3db;
assign v90e36f = jx1_p & v844f91 | !jx1_p & v906042;
assign v8b9de1 = StoB_REQ0_p & v93fd87 | !StoB_REQ0_p & v90ed2f;
assign v93f7dc = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v88946f;
assign v93fc81 = BtoS_ACK8_p & v90776b | !BtoS_ACK8_p & v90adef;
assign v90e6b0 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85eacf;
assign v9080f5 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v905adf;
assign v903d90 = jx1_p & v8b4990 | !jx1_p & v93e898;
assign v907f74 = RtoB_ACK0_p & v93fb21 | !RtoB_ACK0_p & v93f6ff;
assign v93f67b = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v93fe01;
assign v909174 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v93fc8e;
assign v90529c = jx2_p & v844f91 | !jx2_p & v93fe75;
assign v844fcf = DEQ_p & v844f91 | !DEQ_p & !v844f91;
assign v93fb3b = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v93deab;
assign v905425 = jx0_p & v93f665 | !jx0_p & !v89e0b4;
assign v912384 = BtoS_ACK6_p & v9099fa | !BtoS_ACK6_p & v91a75e;
assign v910f62 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v906642;
assign v910515 = jx2_p & v9104d5 | !jx2_p & v930005;
assign v905285 = BtoS_ACK2_p & v9123a2 | !BtoS_ACK2_p & v911ec2;
assign v93f965 = StoB_REQ0_p & v93db4a | !StoB_REQ0_p & v844f91;
assign v93f6fb = jx2_p & v913169 | !jx2_p & v844f91;
assign v844fa3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844f91;
assign v93f6c6 = BtoS_ACK6_p & v9047e4 | !BtoS_ACK6_p & !v90eaab;
assign v930047 = BtoS_ACK6_p & v93f1cf | !BtoS_ACK6_p & v906c94;
assign v93e156 = StoB_REQ0_p & v93fc1a | !StoB_REQ0_p & v844f91;
assign v9040a9 = StoB_REQ7_p & v906fc1 | !StoB_REQ7_p & v93fdb4;
assign v90d52b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v911f1f;
assign v93f994 = jx0_p & v910e17 | !jx0_p & v90d21a;
assign v908f73 = StoB_REQ8_p & v90e2d7 | !StoB_REQ8_p & v93fdd1;
assign v90824e = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v907c85;
assign v907e73 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v9112e1;
assign v8b9b71 = jx1_p & v93f136 | !jx1_p & v904ee9;
assign v9101be = jx2_p & v90a53b | !jx2_p & !v8b4a12;
assign v85eaa5 = StoB_REQ6_p & v911005 | !StoB_REQ6_p & v93f9b4;
assign v9187aa = jx1_p & v93f768 | !jx1_p & v9106a7;
assign v93fc77 = jx1_p & v9056b0 | !jx1_p & v844f91;
assign v90f2f4 = StoB_REQ8_p & v904b00 | !StoB_REQ8_p & v911a72;
assign v90839e = EMPTY_p & v93eadd | !EMPTY_p & v90da38;
assign v91209b = ENQ_p & v844fc3 | !ENQ_p & !v93f3f2;
assign v8b9972 = jx3_p & v844f91 | !jx3_p & v90de74;
assign v93fd54 = StoB_REQ8_p & v93fc85 | !StoB_REQ8_p & v93fda2;
assign v930083 = jx1_p & v93fd1d | !jx1_p & v8b714e;
assign v93f2bd = BtoS_ACK9_p & v93f73d | !BtoS_ACK9_p & v93f801;
assign v90630d = jx0_p & v844f97 | !jx0_p & !v844f95;
assign v90d8d5 = RtoB_ACK0_p & v844fcd | !RtoB_ACK0_p & v844f91;
assign v93f7ab = BtoS_ACK8_p & v904b00 | !BtoS_ACK8_p & v903c4d;
assign v909367 = jx1_p & v844fa3 | !jx1_p & !v844f91;
assign v905eaa = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93ef1d;
assign v844fb7 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v87c558 = BtoS_ACK8_p & v905461 | !BtoS_ACK8_p & !v93f282;
assign v93fe3f = jx2_p & v93fc77 | !jx2_p & v911c6f;
assign v90598f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f61e;
assign v904eba = BtoS_ACK6_p & v93fb3e | !BtoS_ACK6_p & v93fe41;
assign v904de5 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93f6fc;
assign v93f89e = BtoS_ACK6_p & v93e126 | !BtoS_ACK6_p & v844f91;
assign v906915 = BtoS_ACK7_p & v93e27a | !BtoS_ACK7_p & v93e672;
assign v90f947 = jx2_p & v93fb3f | !jx2_p & !v844f91;
assign v904e70 = jx0_p & v910243 | !jx0_p & v93fc9b;
assign v8b98b7 = BtoS_ACK8_p & v9117b1 | !BtoS_ACK8_p & !v8b9bb4;
assign v906e3d = BtoS_ACK6_p & v90ede1 | !BtoS_ACK6_p & v90e76a;
assign v93fdc9 = BtoS_ACK8_p & v90722c | !BtoS_ACK8_p & !v90ddf9;
assign v93f76d = jx1_p & v8b9eca | !jx1_p & !v93f324;
assign v9082fc = jx0_p & v93ee82 | !jx0_p & v90a30e;
assign v90ea47 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v904abe;
assign v86f60a = BtoS_ACK7_p & v904b00 | !BtoS_ACK7_p & v9040fb;
assign v89f948 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v904ae4;
assign v8ee1bc = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v90628f;
assign v910c37 = StoB_REQ7_p & v93f977 | !StoB_REQ7_p & v90e1d0;
assign v90fa03 = StoB_REQ9_p & v90748c | !StoB_REQ9_p & v844f91;
assign v907e8f = jx3_p & v908ad9 | !jx3_p & v9081aa;
assign v93fb61 = jx0_p & v9082e4 | !jx0_p & !v90f7d3;
assign v93f61e = BtoS_ACK1_p & v90534f | !BtoS_ACK1_p & !v90e4ec;
assign v93fb71 = BtoS_ACK7_p & v93e27a | !BtoS_ACK7_p & v90dcf0;
assign v90501e = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v93fc8e;
assign v93fdf7 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v93fd8e;
assign v93fb92 = jx2_p & v85cd12 | !jx2_p & !v844f91;
assign v93fdfe = StoB_REQ1_p & v906627 | !StoB_REQ1_p & v844f91;
assign v90834a = jx3_p & v93fdc0 | !jx3_p & v844fc3;
assign v905252 = BtoS_ACK6_p & v9096ae | !BtoS_ACK6_p & v908083;
assign v910e2d = jx1_p & v90a334 | !jx1_p & v93006d;
assign v90cc30 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f6bc;
assign v9041e4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90a233;
assign v904809 = StoB_REQ7_p & v911c73 | !StoB_REQ7_p & v90fc7f;
assign v90a149 = jx1_p & v93ec50 | !jx1_p & v859635;
assign v9104e0 = BtoS_ACK2_p & v93f9a9 | !BtoS_ACK2_p & v91063d;
assign v93f7f1 = StoB_REQ7_p & v93f9c6 | !StoB_REQ7_p & v910243;
assign v904bc0 = stateG7_1_p & v93f5d7 | !stateG7_1_p & v904852;
assign v903c0d = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v907e3f;
assign v903cda = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8f22e3;
assign SLC0_n = !v863478;
assign v91071c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8f22a2;
assign v90faaf = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93e2c2;
assign v906e08 = jx1_p & v906d3f | !jx1_p & !v904f85;
assign v93fbb8 = BtoS_ACK6_p & v93f90a | !BtoS_ACK6_p & v93f990;
assign v911833 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v90e8fa;
assign v9056a0 = StoB_REQ8_p & v93f769 | !StoB_REQ8_p & v93fd42;
assign v910d70 = BtoS_ACK6_p & v9096ae | !BtoS_ACK6_p & v93fb61;
assign v93fd40 = BtoS_ACK0_p & v93dfc0 | !BtoS_ACK0_p & v93db10;
assign v908a98 = BtoS_ACK1_p & v93dfc0 | !BtoS_ACK1_p & v93fdba;
assign v909197 = stateG7_1_p & v90f8ce | !stateG7_1_p & v904632;
assign v91162e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v93fd5c;
assign v93ece6 = BtoS_ACK8_p & v9043e5 | !BtoS_ACK8_p & v93f86a;
assign v93fb6e = BtoS_ACK8_p & v910d56 | !BtoS_ACK8_p & !v8810ad;
assign v91a6f0 = BtoS_ACK8_p & v93f29a | !BtoS_ACK8_p & v93fe57;
assign v93f541 = jx2_p & v93fd23 | !jx2_p & v93f68a;
assign v9098f2 = BtoS_ACK3_p & v93fd2b | !BtoS_ACK3_p & v93df39;
assign v90ef0d = RtoB_ACK1_p & v90a1c0 | !RtoB_ACK1_p & v93e0e6;
assign v906b71 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v93f6f3;
assign v8a927b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v90d21a;
assign v93f75b = jx1_p & v93e126 | !jx1_p & !v844f91;
assign v909dd5 = EMPTY_p & v93dfb4 | !EMPTY_p & v90a419;
assign v872187 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v93f945;
assign v88c2af = RtoB_ACK0_p & v904c4f | !RtoB_ACK0_p & v904d56;
assign v906131 = jx2_p & v87f17f | !jx2_p & v93f852;
assign v90f0a2 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v905791;
assign v8ee173 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86335a;
assign v93fd67 = ENQ_p & v93eed6 | !ENQ_p & v911013;
assign v93f696 = jx1_p & v844f91 | !jx1_p & !v904f32;
assign v87bf0e = StoB_REQ6_p & v91a6e7 | !StoB_REQ6_p & v909637;
assign v93fb86 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9046de;
assign v8f3849 = StoB_REQ7_p & v93f989 | !StoB_REQ7_p & v93fcda;
assign v904852 = RtoB_ACK0_p & v90494f | !RtoB_ACK0_p & v93fc6c;
assign v910226 = BtoS_ACK8_p & v93e819 | !BtoS_ACK8_p & v90567a;
assign v93ed96 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f906;
assign v93e85e = StoB_REQ8_p & v93f955 | !StoB_REQ8_p & v93fb92;
assign v9061b3 = stateG7_1_p & v93df15 | !stateG7_1_p & v9099f2;
assign v93fd7a = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v93ecc4;
assign v91016c = BtoS_ACK0_p & v90855a | !BtoS_ACK0_p & !v8b9c2c;
assign v90f8ce = RtoB_ACK0_p & v904d81 | !RtoB_ACK0_p & v90cf68;
assign v93ee84 = StoB_REQ0_p & v908fba | !StoB_REQ0_p & v89f844;
assign v911b9a = StoB_REQ8_p & v907e36 | !StoB_REQ8_p & v93f5ae;
assign v90f8d6 = jx1_p & v90eef9 | !jx1_p & v844f91;
assign jx0_n = !v85eb2b;
assign v93f627 = StoB_REQ8_p & v93f4e9 | !StoB_REQ8_p & v907e88;
assign v90df59 = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v844f91;
assign v90dc2c = RtoB_ACK0_p & v90a2f1 | !RtoB_ACK0_p & v90ad6f;
assign v93ed09 = RtoB_ACK0_p & v90444d | !RtoB_ACK0_p & v90ad03;
assign v93f85e = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v93f9a9;
assign v910fd2 = StoB_REQ6_p & v93fbd4 | !StoB_REQ6_p & v906d63;
assign v90a2b9 = jx1_p & v9051bb | !jx1_p & v87f17d;
assign v90a181 = StoB_REQ7_p & v93f796 | !StoB_REQ7_p & v90ad02;
assign v9086d9 = jx1_p & v8f22d1 | !jx1_p & !v93e4c1;
assign v90815c = StoB_REQ6_p & v93fe34 | !StoB_REQ6_p & v90a29a;
assign v93e41f = jx2_p & v904f4d | !jx2_p & v93fb73;
assign v8ebd2a = BtoR_REQ1_p & v93e9c8 | !BtoR_REQ1_p & v93fbce;
assign v8d1873 = BtoS_ACK6_p & v9099fa | !BtoS_ACK6_p & v88e6c4;
assign SLC2_n = !v87cb21;
assign v907adb = jx2_p & v93fb7b | !jx2_p & !v904755;
assign v93fcdc = StoB_REQ8_p & v913428 | !StoB_REQ8_p & v9115a9;
assign v85ea79 = BtoS_ACK1_p & v8bb868 | !BtoS_ACK1_p & v9133ea;
assign v911c6f = jx1_p & v844f91 | !jx1_p & !v93e89f;
assign v93fd4f = StoB_REQ9_p & v909995 | !StoB_REQ9_p & v8b9ce2;
assign v93e77a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v876439;
assign v909f68 = jx1_p & v9091e3 | !jx1_p & v908fb8;
assign v93f91a = jx0_p & v93f682 | !jx0_p & !v93f6fc;
assign v90d64c = ENQ_p & v93eed6 | !ENQ_p & v904bdb;
assign v910820 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v9082d3;
assign v90f5f8 = BtoS_ACK9_p & v93e162 | !BtoS_ACK9_p & v9091dd;
assign v93e2fa = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v90936b;
assign v93f652 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v90decf;
assign v87a242 = StoB_REQ9_p & v904b00 | !StoB_REQ9_p & v90f161;
assign v93e610 = jx1_p & v93fd1d | !jx1_p & v9051ea;
assign v90a6d6 = jx0_p & v93f119 | !jx0_p & v93fc0a;
assign v909e8a = BtoS_ACK8_p & v93f955 | !BtoS_ACK8_p & v93f769;
assign v93e259 = jx2_p & v90a62c | !jx2_p & v911c6f;
assign v905aa1 = EMPTY_p & v93e853 | !EMPTY_p & v93f8b8;
assign v90671f = jx0_p & v904de5 | !jx0_p & !v844f95;
assign v90894d = BtoS_ACK6_p & v90fb5d | !BtoS_ACK6_p & v8f22d0;
assign v912334 = jx3_p & v93f78c | !jx3_p & !v93f2bd;
assign v91aa7d = BtoR_REQ1_p & v93fab8 | !BtoR_REQ1_p & v90f4f7;
assign v911f15 = jx2_p & v93eda5 | !jx2_p & v908ed6;
assign v93fbb7 = BtoS_ACK6_p & v93f91d | !BtoS_ACK6_p & v93fe64;
assign v93e596 = jx2_p & v90ef16 | !jx2_p & v908ed6;
assign v9058f1 = BtoS_ACK0_p & v913561 | !BtoS_ACK0_p & v93fab0;
assign v904b7f = BtoS_ACK9_p & v93f8e0 | !BtoS_ACK9_p & v87a98d;
assign v90805e = jx0_p & v93f29e | !jx0_p & v93ec44;
assign v907d33 = StoB_REQ6_p & v90ff24 | !StoB_REQ6_p & v844f91;
assign v9062b3 = BtoS_ACK6_p & v930032 | !BtoS_ACK6_p & v93fd3c;
assign v906717 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v907add;
assign v9071f8 = BtoS_ACK6_p & v863a78 | !BtoS_ACK6_p & v904f5c;
assign v90a229 = jx2_p & v863476 | !jx2_p & !v90fc9a;
assign v93fb43 = jx2_p & v9057c1 | !jx2_p & v93f75b;
assign v913619 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9d;
assign v9053de = BtoS_ACK6_p & v93f8cf | !BtoS_ACK6_p & v904ae8;
assign v90479c = jx0_p & v906f44 | !jx0_p & v89f803;
assign v87575e = StoB_REQ9_p & v844f91 | !StoB_REQ9_p & v90f787;
assign v93f533 = jx1_p & v844f91 | !jx1_p & v863363;
assign v9074fa = jx2_p & v87c51f | !jx2_p & !v907e86;
assign v8b9b9f = jx0_p & v90ef1b | !jx0_p & v903c46;
assign v91086d = StoB_REQ1_p & v93e926 | !StoB_REQ1_p & v904808;
assign v909016 = StoB_REQ2_p & v93fdf7 | !StoB_REQ2_p & v904c75;
assign v907c59 = BtoS_ACK6_p & v90d880 | !BtoS_ACK6_p & v90aa8a;
assign v93e648 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v93fd5f;
assign v93dbf1 = jx1_p & v90515d | !jx1_p & v844f91;
assign v90500e = DEQ_p & v909878 | !DEQ_p & v87c51e;
assign v91267e = BtoS_ACK4_p & v844f9f | !BtoS_ACK4_p & v844f9d;
assign v90a75f = jx2_p & v90d93b | !jx2_p & v844f91;
assign v93f7e9 = jx1_p & v93f1cf | !jx1_p & !v910bea;
assign v93fbe6 = jx0_p & v93fbd6 | !jx0_p & v93fb64;
assign v90fa8a = StoB_REQ7_p & v903e94 | !StoB_REQ7_p & v93e903;
assign v91335a = DEQ_p & v9043bd | !DEQ_p & v93f9cb;
assign v9044c6 = jx0_p & v909e2c | !jx0_p & !v844f91;
assign v93fb09 = jx1_p & v86f4a3 | !jx1_p & v911451;
assign v93fe01 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v90631b;
assign v905539 = BtoS_ACK9_p & v87f17f | !BtoS_ACK9_p & v908fb4;
assign v93e3a5 = DEQ_p & v90567c | !DEQ_p & v93fbc1;
assign v9095ec = jx2_p & v93fbd0 | !jx2_p & v844f91;
assign v90a451 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85ea5f;
assign v93f7b3 = BtoS_ACK7_p & v93fd84 | !BtoS_ACK7_p & v93fb8d;
assign v910473 = StoB_REQ6_p & v93f682 | !StoB_REQ6_p & v90f88e;
assign v904bbf = BtoS_ACK8_p & v93ec47 | !BtoS_ACK8_p & v903cda;
assign v93f0bf = RtoB_ACK1_p & v93fb8a | !RtoB_ACK1_p & v910221;
assign v85cd12 = jx1_p & v909dde | !jx1_p & v844f91;
assign v90fa0b = jx1_p & v9047cd | !jx1_p & v844f91;
assign v910be8 = BtoS_ACK1_p & v93dffe | !BtoS_ACK1_p & v90efe2;
assign v904f2e = BtoS_ACK1_p & v93e2de | !BtoS_ACK1_p & v90631b;
assign v907633 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v903c6e;
assign v93fe1f = StoB_REQ7_p & v8821a1 | !StoB_REQ7_p & v844f91;
assign v9133d9 = BtoS_ACK1_p & v93f85e | !BtoS_ACK1_p & v90914c;
assign v904eea = StoB_REQ8_p & v90944f | !StoB_REQ8_p & !v90477e;
assign v93e996 = StoB_REQ9_p & v93f2c6 | !StoB_REQ9_p & v93f584;
assign v8850b3 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v9095d0;
assign v90950c = stateG12_p & v908ad9 | !stateG12_p & !v93dfc2;
assign v9045df = jx2_p & v93fda7 | !jx2_p & v93e68f;
assign v93eb41 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v90dc28;
assign v90add6 = StoB_REQ9_p & v91a7a3 | !StoB_REQ9_p & v93ef76;
assign v90a44f = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v93f7bb;
assign v93fe69 = StoB_REQ9_p & v90dd77 | !StoB_REQ9_p & v8f381e;
assign v8b8638 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v93f702;
assign v91007f = RtoB_ACK0_p & v904b94 | !RtoB_ACK0_p & v912d1a;
assign v93f9c7 = jx1_p & v913a39 | !jx1_p & !v844f91;
assign v906eb2 = stateG7_1_p & v93ecad | !stateG7_1_p & v93e2b8;
assign v90490e = BtoS_ACK9_p & v93fcc4 | !BtoS_ACK9_p & v90fa80;
assign v90fd1c = BtoS_ACK7_p & v911f15 | !BtoS_ACK7_p & v93faff;
assign v910ebb = StoB_REQ8_p & v904838 | !StoB_REQ8_p & v93e810;
assign v93fd3e = FULL_p & v87e0d8 | !FULL_p & v92ffd3;
assign v908a03 = jx1_p & v90804e | !jx1_p & v909222;
assign v93f444 = BtoS_ACK7_p & v90529c | !BtoS_ACK7_p & v90ebe8;
assign v93fce5 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v93fcbe;
assign v93e3f1 = ENQ_p & v907c69 | !ENQ_p & v90e5b4;
assign v9113ea = EMPTY_p & v905355 | !EMPTY_p & v90513b;
assign v93e60f = StoB_REQ7_p & v93ee3b | !StoB_REQ7_p & v844f91;
assign v90edca = jx2_p & v870dd6 | !jx2_p & v880314;
assign v86dde6 = BtoS_ACK8_p & v93f7f8 | !BtoS_ACK8_p & v93f7b4;
assign v93fe75 = jx1_p & v90787b | !jx1_p & v844f91;
assign v90656f = BtoS_ACK9_p & v90d78b | !BtoS_ACK9_p & !v9051da;
assign v90738d = jx2_p & v93f678 | !jx2_p & v863afc;
assign v905461 = jx2_p & v90ae9a | !jx2_p & v8a8fdd;
assign v910c51 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v93e7d1;
assign v870fb9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v908d05;
assign v90505e = RtoB_ACK0_p & v907bb9 | !RtoB_ACK0_p & v93f6d0;
assign v91a73f = BtoS_ACK8_p & v93e596 | !BtoS_ACK8_p & v908f73;
assign v904b99 = jx3_p & v93fa3a | !jx3_p & !v93daf2;
assign v93fbd2 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v908eea;
assign v89f938 = BtoS_ACK6_p & v93f1cf | !BtoS_ACK6_p & v93f94a;
assign v93f9d7 = EMPTY_p & v93e301 | !EMPTY_p & v904b09;
assign v8a8fda = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v906c10;
assign v86e831 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v888002;
assign v93f0a9 = BtoS_ACK6_p & v9050a5 | !BtoS_ACK6_p & v93fca3;
assign v93eece = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v9047b7;
assign v90a20e = BtoS_ACK1_p & v90da97 | !BtoS_ACK1_p & v9094ed;
assign v93f738 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v9046a6;
assign v93ec83 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v90f500;
assign v9083d3 = StoB_REQ1_p & v906642 | !StoB_REQ1_p & !v90a233;
assign v90d364 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v91a771;
assign v9059b7 = jx0_p & v9054b5 | !jx0_p & !v90664a;
assign v90e027 = DEQ_p & v8f22ca | !DEQ_p & v904dc1;
assign v93ec9d = BtoS_ACK6_p & v86344b | !BtoS_ACK6_p & v90fa5e;
assign v90fa88 = ENQ_p & v9101d0 | !ENQ_p & v8b9972;
assign v93f822 = BtoS_ACK8_p & v90451f | !BtoS_ACK8_p & v904610;
assign v90ba2c = StoB_REQ2_p & v93fcf0 | !StoB_REQ2_p & v8a8fda;
assign v87261e = RtoB_ACK0_p & v907bb9 | !RtoB_ACK0_p & v904e3a;
assign v90d698 = BtoS_ACK2_p & v90854b | !BtoS_ACK2_p & v905d37;
assign v93faab = jx2_p & v8b9b71 | !jx2_p & v8f60f9;
assign v908574 = StoB_REQ1_p & v90636e | !StoB_REQ1_p & v91093c;
assign v93fae1 = BtoS_ACK9_p & v9114a0 | !BtoS_ACK9_p & v93f5cb;
assign v90e6f8 = BtoS_ACK7_p & v90f575 | !BtoS_ACK7_p & v93f91f;
assign v93e065 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v93ebe6;
assign v93f5d7 = RtoB_ACK0_p & v90494f | !RtoB_ACK0_p & v93fd85;
assign v93ef2e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v93fce0;
assign v93f02f = jx1_p & v906dd6 | !jx1_p & v844f91;
assign v93fe5b = BtoS_ACK2_p & v90e978 | !BtoS_ACK2_p & v93ef30;
assign ENQ_n = (BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((RtoB_ACK0_n) | (!RtoB_ACK0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!DEQ_n & ((RtoB_ACK0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((BtoR_REQ0_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))) | (!DEQ_n & ((BtoR_REQ0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_1_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!stateG7_1_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n) | (!RtoB_ACK0_n & ((stateG7_0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!stateG7_0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((BtoR_REQ0_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))) | (!DEQ_n & ((BtoR_REQ0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))))) | (!jx3_n & ((jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((StoB_REQ9_n))) | (!BtoS_ACK9_n & ((jx0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))) | (!StoB_REQ6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))))))))))))))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!SLC0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))))))) | (!SLC1_n & ((SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!SLC2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n)))))))))))))))))))))))))))))))))))))))))))))));
assign SLC3_n = (BtoR_REQ1_n & ((EMPTY_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!DEQ_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((BtoR_REQ0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!BtoR_REQ0_n & ((stateG7_0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG7_0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((BtoR_REQ0_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!stateG7_1_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!DEQ_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((BtoR_REQ0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!BtoR_REQ0_n & ((stateG7_0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG7_0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((BtoR_REQ0_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!stateG7_1_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!DEQ_n & ((BtoR_REQ0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!RtoB_ACK0_n & ((stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))) | (!stateG12_n & ((jx3_n & ((jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx1_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((jx0_n & ((StoB_REQ9_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!StoB_REQ9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))) | (!jx0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))))))))))) | (!jx3_n & ((BtoS_ACK9_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK9_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC1_n) | (!SLC1_n & ((SLC2_n)))))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  StoB_REQ4_p = 0;
  StoB_REQ5_p = 0;
  StoB_REQ6_p = 0;
  StoB_REQ7_p = 0;
  StoB_REQ8_p = 0;
  StoB_REQ9_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoS_ACK4_p = 0;
  BtoS_ACK5_p = 0;
  BtoS_ACK6_p = 0;
  BtoS_ACK7_p = 0;
  BtoS_ACK8_p = 0;
  BtoS_ACK9_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  SLC2_p = 0;
  SLC3_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
  jx3_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  StoB_REQ4_p = StoB_REQ4_n;
  StoB_REQ5_p = StoB_REQ5_n;
  StoB_REQ6_p = StoB_REQ6_n;
  StoB_REQ7_p = StoB_REQ7_n;
  StoB_REQ8_p = StoB_REQ8_n;
  StoB_REQ9_p = StoB_REQ9_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoS_ACK4_p = BtoS_ACK4_n;
  BtoS_ACK5_p = BtoS_ACK5_n;
  BtoS_ACK6_p = BtoS_ACK6_n;
  BtoS_ACK7_p = BtoS_ACK7_n;
  BtoS_ACK8_p = BtoS_ACK8_n;
  BtoS_ACK9_p = BtoS_ACK9_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  SLC2_p = SLC2_n;
  SLC3_p = SLC3_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
  jx3_p = jx3_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
