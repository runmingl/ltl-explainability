module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, StoB_REQ4_n, StoB_REQ5_n, StoB_REQ6_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoS_ACK4_n, BtoS_ACK5_n, BtoS_ACK6_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, SLC2_n, jx0_n, jx1_n, jx2_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844fb7;
  wire v8fd879;
  wire v844fa1;
  wire v882006;
  wire v8944a2;
  wire v892417;
  wire v8fd1ea;
  wire v8b6040;
  wire v882c70;
  wire v884a9c;
  wire v88483c;
  wire v8fd5cd;
  wire v887b60;
  wire v8fd398;
  wire v887f6f;
  wire v8fd755;
  wire v887a78;
  wire v8fd7e9;
  wire v86ed7e;
  wire v883d82;
  wire v844f9f;
  wire v88576e;
  wire v8fd646;
  wire v8fd932;
  wire v885dfd;
  wire v8fd6d6;
  wire v8fd2a7;
  wire v8841f8;
  wire v8ad074;
  wire v88fa1c;
  wire v887d49;
  wire v8c4cf8;
  wire v8fd8a4;
  wire v88234e;
  wire v8879eb;
  wire v8802a9;
  wire v8fc7c3;
  wire v8fd443;
  wire v8811aa;
  wire v844f9d;
  wire v8fd5ad;
  wire v88219e;
  wire v884ac0;
  wire v8c2e72;
  wire v88eb82;
  wire v887f3a;
  wire v8fd6b3;
  wire v88786f;
  wire v891077;
  wire v88618b;
  wire v8fd8a5;
  wire v89fadb;
  wire v884dd2;
  wire v844f9b;
  wire v882bdd;
  wire v8fd764;
  wire v880fd1;
  wire v8fd5dc;
  wire v881f1a;
  wire v8fd775;
  wire v8dacbf;
  wire v8850d3;
  wire v880b56;
  wire v882473;
  wire v844f99;
  wire v88eb87;
  wire v8836c4;
  wire v8ad0e2;
  wire v882fc1;
  wire v88f1b0;
  wire v8fcc5a;
  wire v8b6053;
  wire v887dc2;
  wire v8972fa;
  wire v887d9a;
  wire v844f97;
  wire v8fd5c9;
  wire v853f24;
  wire v880717;
  wire v880616;
  wire v88945f;
  wire v8fd84e;
  wire v8fd1ac;
  wire v8c2ecf;
  wire v88401d;
  wire v8830a5;
  wire v88386a;
  wire v8fd62e;
  wire v8c2df5;
  wire v8fd197;
  wire v885c13;
  wire v8fd327;
  wire v8836b1;
  wire v887924;
  wire v884b2b;
  wire v8830ac;
  wire v887f47;
  wire v88a2df;
  wire v8a88c6;
  wire v883706;
  wire v880c71;
  wire v8fd88a;
  wire v8f2abd;
  wire v8879f2;
  wire v8fc19e;
  wire v8fc986;
  wire v880383;
  wire v8fd86a;
  wire v8fcd32;
  wire v884531;
  wire v8819d6;
  wire v8822d4;
  wire v883c14;
  wire v884171;
  wire v887b14;
  wire v88289d;
  wire v8fd819;
  wire v8fd5ab;
  wire v8fd83e;
  wire v895b93;
  wire v8fd2ab;
  wire v881e67;
  wire v8fd588;
  wire v892c48;
  wire v8fd4c4;
  wire v883879;
  wire v8fd63c;
  wire v880f9a;
  wire v8b60ca;
  wire v8fd810;
  wire v85582e;
  wire v8b89cf;
  wire v8fc46b;
  wire v88576c;
  wire v885fe4;
  wire v8dabe8;
  wire v854be6;
  wire v88429a;
  wire v8fd1f1;
  wire v883f90;
  wire v8fc651;
  wire v887f13;
  wire v8fd1cd;
  wire v885867;
  wire v8c48b6;
  wire v88802b;
  wire v887f97;
  wire v8fc688;
  wire v8ce150;
  wire v882d19;
  wire v8dac3a;
  wire v8828b1;
  wire v8fd6f9;
  wire v8fd71e;
  wire v87fee2;
  wire v882f43;
  wire v8fd78b;
  wire v8fd7cc;
  wire v883ea8;
  wire v885660;
  wire v883cf0;
  wire v8fd8f3;
  wire v890d96;
  wire v8c2eb4;
  wire v8842ac;
  wire v885c06;
  wire v881f61;
  wire v8825e6;
  wire v8fc810;
  wire v88225a;
  wire v883817;
  wire v884497;
  wire v897c49;
  wire v8f2aa9;
  wire v8846bf;
  wire v85839b;
  wire v880933;
  wire v887734;
  wire v8daca2;
  wire v8876bb;
  wire v8fd704;
  wire v891da3;
  wire v8876d0;
  wire v8a88d6;
  wire v844faf;
  wire v8fd866;
  wire v8fd6ec;
  wire v8fcdd0;
  wire v884e81;
  wire v8fd7c7;
  wire v87fee8;
  wire v8fd6d3;
  wire v883ee4;
  wire v887adb;
  wire v883bb8;
  wire v8f2a3f;
  wire v88271c;
  wire v8947da;
  wire v88404f;
  wire v8fd6cd;
  wire v882d86;
  wire v880d9c;
  wire v8fd54e;
  wire v882c77;
  wire v8fd5b7;
  wire v8fd79c;
  wire v885d96;
  wire v891109;
  wire v885be7;
  wire v8fd7cb;
  wire v8fd8cf;
  wire v8811a0;
  wire v885f78;
  wire v897405;
  wire v884a91;
  wire v88193e;
  wire v8fd8c7;
  wire v8fd70d;
  wire v8fd587;
  wire v8fd163;
  wire v8c2e4a;
  wire v887e01;
  wire v8fd85f;
  wire v885077;
  wire v8c2ea3;
  wire v882d6b;
  wire v8fd315;
  wire v8fd7b7;
  wire v88c127;
  wire v887d74;
  wire v8588b1;
  wire v891114;
  wire v885694;
  wire v895d61;
  wire v8fc312;
  wire v8fd5ed;
  wire v875145;
  wire v8dabff;
  wire v882505;
  wire v8841eb;
  wire v8fd7e8;
  wire v8fd782;
  wire v882d8f;
  wire v8825e5;
  wire v8842b7;
  wire v8fd3b5;
  wire v8fd8ff;
  wire v884216;
  wire v8fd202;
  wire v8fc77f;
  wire v8fd8e2;
  wire v8fd5a6;
  wire v881686;
  wire v895b31;
  wire v897cf5;
  wire v8808eb;
  wire v8811e6;
  wire v895d68;
  wire v8fd172;
  wire v8831c8;
  wire v8fd8cd;
  wire v885ffa;
  wire v8fd1a8;
  wire v8fd8b9;
  wire v8fd797;
  wire v8dacfc;
  wire v885c4b;
  wire v8fd6e3;
  wire v8a87f2;
  wire v8823d8;
  wire v8fd94e;
  wire v87a65f;
  wire v8fd33e;
  wire v8fd881;
  wire v866b82;
  wire v86ecdb;
  wire v8fd66c;
  wire v8fd90f;
  wire v8fc1f9;
  wire v88052d;
  wire v8f2a19;
  wire v8fd4f5;
  wire v895abb;
  wire v895b24;
  wire v8dac30;
  wire v88a63c;
  wire v897358;
  wire v8fd895;
  wire v884d49;
  wire v8ac1f3;
  wire v8c2e6c;
  wire v8fd739;
  wire v8859ec;
  wire v8ac9bd;
  wire v8fcfe7;
  wire v8fd75d;
  wire v882a93;
  wire v8847be;
  wire v8fd8b4;
  wire v880e79;
  wire v8fd8dd;
  wire v8fc2b2;
  wire v8fc182;
  wire v8fc691;
  wire v8ad047;
  wire v8fd5f2;
  wire v883d9e;
  wire v884335;
  wire v887d86;
  wire v882c31;
  wire v8fd873;
  wire v8fd22d;
  wire v88e2d2;
  wire v883fee;
  wire v8fd58e;
  wire v8ac9e4;
  wire v8a87de;
  wire v8849ea;
  wire v896e20;
  wire v8fd596;
  wire v858501;
  wire v879b9f;
  wire v883cf7;
  wire v890b45;
  wire v885ec1;
  wire v8fd260;
  wire v89735b;
  wire v884d94;
  wire v881fe6;
  wire v88372b;
  wire v884adf;
  wire v86ed40;
  wire v8824dc;
  wire v8817c2;
  wire v8a7071;
  wire v8fd607;
  wire v8fd86e;
  wire v88044e;
  wire v8fd185;
  wire v880dba;
  wire v8845c3;
  wire v8879aa;
  wire v882e00;
  wire v887b5e;
  wire v88565e;
  wire v8861a4;
  wire v8830bd;
  wire v880403;
  wire v8ed1a5;
  wire v8fc1f8;
  wire v8876cd;
  wire v8fd5e5;
  wire v8fd8ac;
  wire v88582f;
  wire v89facc;
  wire v8fd698;
  wire v8fd6e7;
  wire v8816be;
  wire v88621e;
  wire v88616c;
  wire v880fe9;
  wire v8fd727;
  wire v876115;
  wire v89fac8;
  wire v87943e;
  wire v8fd7d3;
  wire v8fd636;
  wire v8816e8;
  wire v881923;
  wire v8fd5e8;
  wire v88772e;
  wire v895d4e;
  wire v8fd710;
  wire v8fd7bf;
  wire v883c3b;
  wire v8fd71c;
  wire v8f2abf;
  wire v844fa3;
  wire v8676b7;
  wire v8fd5df;
  wire v8fd967;
  wire v8fd088;
  wire v88e5f0;
  wire v8fd8af;
  wire v87d10c;
  wire v8fd6f3;
  wire v8851dd;
  wire v8fd6fc;
  wire v88093b;
  wire v883ddb;
  wire v8fd8d8;
  wire v8563aa;
  wire v8846ff;
  wire v887f44;
  wire v8fd6a6;
  wire v887fa9;
  wire v883f65;
  wire v844f95;
  wire v8ce165;
  wire v8fd77b;
  wire v8fd356;
  wire v8fd916;
  wire v8fc7f4;
  wire v854113;
  wire v880a21;
  wire v885cf3;
  wire v8fd690;
  wire v8f29f1;
  wire v8fd28e;
  wire v8fd8d1;
  wire v8fd014;
  wire v8fd658;
  wire v882a63;
  wire v89484f;
  wire v87bb99;
  wire v8972d8;
  wire v884b56;
  wire v885da7;
  wire v844fb1;
  wire v882b6f;
  wire v887bf3;
  wire v88800a;
  wire v886176;
  wire v8fd76a;
  wire v88fa9e;
  wire v887d85;
  wire v88565d;
  wire v88ebbe;
  wire v887913;
  wire v89110a;
  wire v8fd7fb;
  wire v86ed36;
  wire v8fd947;
  wire v878328;
  wire v880760;
  wire v8fd667;
  wire v8fd576;
  wire v8fd8cc;
  wire v8840b0;
  wire v8821b5;
  wire v887a24;
  wire v8c48b3;
  wire v8fd5eb;
  wire v8fd5da;
  wire v85cf4b;
  wire v883852;
  wire v8562b0;
  wire v8fc3e8;
  wire v8b6088;
  wire v8fd204;
  wire v8fc7cc;
  wire v8540de;
  wire v884b89;
  wire v8fd1ce;
  wire v8fd830;
  wire v8fd760;
  wire v8818a8;
  wire v8809c4;
  wire v885863;
  wire v8fd084;
  wire v8f2a03;
  wire v8824d4;
  wire v8fd921;
  wire v8fd585;
  wire v8fd94b;
  wire v880982;
  wire v8973aa;
  wire v885bcf;
  wire v880fa6;
  wire v891ac4;
  wire v8cd9c1;
  wire v8fcd47;
  wire v884203;
  wire v887abb;
  wire v885733;
  wire v8fd832;
  wire v88fcc6;
  wire v885c0e;
  wire v88784a;
  wire v885f76;
  wire v8fd952;
  wire v8fd908;
  wire v8b5fbd;
  wire v887904;
  wire v8fcb34;
  wire v8fd672;
  wire v885723;
  wire v88fa48;
  wire v8ce184;
  wire v8fd745;
  wire v8fd74b;
  wire v88086e;
  wire v8fd7cf;
  wire v88497c;
  wire v882136;
  wire v8795bb;
  wire v883e9b;
  wire v881fdb;
  wire v8fc8ad;
  wire v895b52;
  wire v85872e;
  wire v8dabf0;
  wire v8fcae9;
  wire v88810b;
  wire v853f4e;
  wire v8fd5a5;
  wire v8876ed;
  wire v8fd5a1;
  wire v887f70;
  wire v8fd595;
  wire v8ed1f7;
  wire v844fa5;
  wire v8ac9d6;
  wire v8fd94f;
  wire v8fce18;
  wire v887906;
  wire v8fc862;
  wire v883824;
  wire v8fd8fe;
  wire v8bb760;
  wire v8817bd;
  wire v8fd6d7;
  wire v882276;
  wire v8b6045;
  wire v8fd848;
  wire v88058c;
  wire v880cff;
  wire v880f9f;
  wire v8fd18d;
  wire v8fd58c;
  wire v8fc1c0;
  wire v8591df;
  wire v8fd4e5;
  wire v884f1f;
  wire v8d6a33;
  wire v88096f;
  wire v884049;
  wire v88033b;
  wire v884fdd;
  wire v8859f7;
  wire v88164d;
  wire v8fd179;
  wire v8830a3;
  wire v8fd777;
  wire v88190c;
  wire v885bba;
  wire v8dac46;
  wire v881113;
  wire v8c2eb8;
  wire v8fd899;
  wire v8fd8bc;
  wire v8fd65a;
  wire v879486;
  wire v8fd0e6;
  wire v8fcc2e;
  wire v884256;
  wire v8fd221;
  wire v883762;
  wire v8824a9;
  wire v881fa4;
  wire v8820f2;
  wire v8fd285;
  wire v8fd95a;
  wire v887680;
  wire v884b78;
  wire v8c4d26;
  wire v8fccf0;
  wire v8fca9c;
  wire v8878a5;
  wire v8dac78;
  wire v88507a;
  wire v8fd664;
  wire v892b90;
  wire v8fd6ea;
  wire v8840c7;
  wire v8fd57d;
  wire v88402c;
  wire v8fc1cf;
  wire v8fd8df;
  wire v87653c;
  wire v8c2e5d;
  wire v8fd1e1;
  wire v8588ba;
  wire v8fca9d;
  wire v884dec;
  wire v885e24;
  wire v8fd72e;
  wire v884fc8;
  wire v881630;
  wire v884767;
  wire v884476;
  wire v8fd8c0;
  wire v8843d1;
  wire v8fd24f;
  wire v8fd856;
  wire v884b6c;
  wire v88496e;
  wire v894620;
  wire v898f1a;
  wire v882431;
  wire v8fd6f2;
  wire v884d67;
  wire v883ad4;
  wire v88fdf5;
  wire v87b523;
  wire v88264d;
  wire v8fd1e2;
  wire v88785e;
  wire v8fd7c8;
  wire v88807f;
  wire v8fd1da;
  wire v895c65;
  wire v883752;
  wire v8fd243;
  wire v8fd922;
  wire v8fd809;
  wire v868d2b;
  wire v89488f;
  wire v8cd9b9;
  wire v88837d;
  wire v8c2eaf;
  wire v8fd818;
  wire v885fda;
  wire v8881bb;
  wire v8fd812;
  wire v8fd841;
  wire v8fd7af;
  wire v8837c5;
  wire v8816f3;
  wire v8fd379;
  wire v885fe3;
  wire v8fd6d8;
  wire v8fc21f;
  wire v8fc237;
  wire v883a94;
  wire v8838dc;
  wire v8fd7e6;
  wire v8dac8a;
  wire v897374;
  wire v887fd5;
  wire v854c1c;
  wire v8831e6;
  wire v854d5c;
  wire v8880b3;
  wire v88397d;
  wire v88315a;
  wire v882066;
  wire v8fd592;
  wire v8fd849;
  wire v8fd254;
  wire v8a8734;
  wire v88265b;
  wire v8809b9;
  wire v8822bf;
  wire v8878b5;
  wire v8fc762;
  wire v8fd6b6;
  wire v8fd90c;
  wire v888057;
  wire v8fd5ff;
  wire v887c3e;
  wire v8fcefb;
  wire v887ad8;
  wire v887d78;
  wire v885185;
  wire v8fd3ee;
  wire v885fe8;
  wire v8818ad;
  wire v8856f5;
  wire v884c7a;
  wire v8fd0b7;
  wire v8fd353;
  wire v884882;
  wire v8810dc;
  wire v88107d;
  wire v8fd58b;
  wire v892c64;
  wire v86a020;
  wire v8dac82;
  wire v8948c3;
  wire v88029d;
  wire v887bbb;
  wire v883710;
  wire v883700;
  wire v8fd00a;
  wire v892c36;
  wire v8ad0d9;
  wire v887c2f;
  wire v89fb49;
  wire v880665;
  wire v8fd8f8;
  wire v88040b;
  wire v8fd7e3;
  wire v882b15;
  wire v8878da;
  wire v89fb74;
  wire v8fc19f;
  wire v8817cc;
  wire v8810a6;
  wire v8fd67c;
  wire v8fd746;
  wire v87af07;
  wire v881840;
  wire v8fc78f;
  wire v885695;
  wire v8d4bf0;
  wire v8fd6a5;
  wire v8fd917;
  wire v88084d;
  wire v8fc982;
  wire v8fd700;
  wire v89471b;
  wire v88f618;
  wire v883a7f;
  wire v8fc68e;
  wire v894636;
  wire v880931;
  wire v881e80;
  wire v883c48;
  wire v88186b;
  wire v885d25;
  wire v885b17;
  wire v883759;
  wire v8fd78e;
  wire v884796;
  wire v895c47;
  wire v88369c;
  wire v8876c3;
  wire v8947e0;
  wire v8fd1bc;
  wire v8fd906;
  wire v884834;
  wire v88f9d2;
  wire v880e82;
  wire v883ed8;
  wire v8fc2b8;
  wire v884206;
  wire v8fd6b2;
  wire v880ed2;
  wire v880ccb;
  wire v8fca41;
  wire v8fd953;
  wire v8fd74e;
  wire v882baa;
  wire v884919;
  wire v8fc6a5;
  wire v8fcbc7;
  wire v8857e5;
  wire v8839d5;
  wire v8fd75c;
  wire v880ac1;
  wire v895b2a;
  wire v88578e;
  wire v887d16;
  wire v8fc1a7;
  wire v8821ba;
  wire v8f11a7;
  wire v8fd817;
  wire v880ab4;
  wire v882d4e;
  wire v8811ca;
  wire v881172;
  wire v8fc732;
  wire v8806c7;
  wire v883f1b;
  wire v8fd20e;
  wire v8fc61e;
  wire v8fd738;
  wire v8cecad;
  wire v8fd1d7;
  wire v884ba1;
  wire v8877e9;
  wire v882a0a;
  wire v886048;
  wire v858985;
  wire v8793ad;
  wire v8876f2;
  wire v8fd1a1;
  wire v8fcc77;
  wire v876549;
  wire v8fd8ab;
  wire v8819b3;
  wire v87afd1;
  wire v884421;
  wire v8831ee;
  wire v8fd7ff;
  wire v8881fb;
  wire v8fd23e;
  wire v8fd3cb;
  wire v895b92;
  wire v8fd70f;
  wire v8826bd;
  wire v89fb10;
  wire v88e7c3;
  wire v8fd17b;
  wire v8fd5b3;
  wire v8fc1d2;
  wire v8fd600;
  wire v884031;
  wire v8fd7ba;
  wire v86ed35;
  wire v8fd75f;
  wire v8819ce;
  wire v880934;
  wire v8846a5;
  wire v8fd8b1;
  wire v8fd0a4;
  wire v88299b;
  wire v8b605d;
  wire v882a61;
  wire v89fb1e;
  wire v88808a;
  wire v858320;
  wire v880abb;
  wire v8fd678;
  wire v8fd7a0;
  wire v8fd734;
  wire v8fd1d8;
  wire v8fd864;
  wire v887ab9;
  wire v8fd813;
  wire v882f82;
  wire v895aff;
  wire v885f26;
  wire v8fd652;
  wire v884f8c;
  wire v8684ff;
  wire v88808c;
  wire v88a5d1;
  wire v88963d;
  wire v8fd230;
  wire v88fc61;
  wire v88089e;
  wire v8877c1;
  wire v858678;
  wire v890ce8;
  wire v885b96;
  wire v884cd5;
  wire v8fd741;
  wire v8ad078;
  wire v885836;
  wire v895b02;
  wire v882459;
  wire v8b607f;
  wire v8fc73e;
  wire v895ccc;
  wire v88254c;
  wire v8ad0bf;
  wire v8fc35c;
  wire v8846d2;
  wire v880f76;
  wire v882b85;
  wire v8fd95f;
  wire v886092;
  wire v8fd1af;
  wire v8fd7b3;
  wire v8840af;
  wire v8ac9d2;
  wire v8fc99d;
  wire v8fceeb;
  wire v8fccca;
  wire v8972a7;
  wire v8fd581;
  wire v879e64;
  wire v8808f4;
  wire v895d6d;
  wire v8837af;
  wire v8f2a07;
  wire v8fd95c;
  wire v8880e0;
  wire v884197;
  wire v88112b;
  wire v8fd231;
  wire v885713;
  wire v8fd6cc;
  wire v8fd5b1;
  wire v8a705e;
  wire v8fd4a9;
  wire v88172f;
  wire v8fd5b6;
  wire v87fed4;
  wire v887b15;
  wire v8fd568;
  wire v894b33;
  wire v8fd882;
  wire v86f4d0;
  wire v882563;
  wire v8ad115;
  wire v884976;
  wire v883a4d;
  wire v895ceb;
  wire v8766ed;
  wire v898f2f;
  wire v882417;
  wire v854d12;
  wire v88097a;
  wire v883776;
  wire v880dc0;
  wire v880952;
  wire v8fd1de;
  wire v892416;
  wire v8fd1c9;
  wire v8fd724;
  wire v8c2ee6;
  wire v88464a;
  wire v891ab3;
  wire v8fd6ff;
  wire v8ceca9;
  wire v8fd19b;
  wire v8fd8e5;
  wire v8847f1;
  wire v8fd8c5;
  wire v8fc729;
  wire v8dab8a;
  wire v8fd490;
  wire v879570;
  wire v8c2de4;
  wire v884f4a;
  wire v8dacf2;
  wire v8fd24d;
  wire v8fd1b8;
  wire v88201b;
  wire v884de8;
  wire v885e9b;
  wire v8fd24e;
  wire v895bb9;
  wire v88363c;
  wire v88251e;
  wire v882d4a;
  wire v8f2a5f;
  wire v88489f;
  wire v8794e0;
  wire v8fd0b4;
  wire v883791;
  wire v8fd1f3;
  wire v889dee;
  wire v884a33;
  wire v8fd796;
  wire v880cf5;
  wire v882fda;
  wire v885e59;
  wire v8fd93c;
  wire v880a73;
  wire v8fd620;
  wire v8539e7;
  wire v8fd5d1;
  wire v8fd3c6;
  wire v8b605e;
  wire v8857fb;
  wire v86ec4a;
  wire v8fcba5;
  wire v8fce0d;
  wire v8ac9ad;
  wire v880b2d;
  wire v8fd893;
  wire v8fd786;
  wire v854bb9;
  wire v8fd6c5;
  wire v8fd589;
  wire v8fd67e;
  wire v883105;
  wire v8fca4a;
  wire v887b09;
  wire v8fd2b1;
  wire v8c4d01;
  wire v8837ba;
  wire v8fc2e4;
  wire v8fc295;
  wire v88579b;
  wire v8fd87f;
  wire v89386c;
  wire v8fd1f9;
  wire v8fd655;
  wire v88bc53;
  wire v8fd610;
  wire v88ea5a;
  wire v8fcbb4;
  wire v8dab62;
  wire v85e9fa;
  wire v87954a;
  wire v882a5a;
  wire v880c8a;
  wire v8ac1f8;
  wire v8a87b1;
  wire v882ae8;
  wire v8819fb;
  wire v8fd5d3;
  wire v8805be;
  wire v880c81;
  wire v8fd91b;
  wire v8856d5;
  wire v8fce44;
  wire v8fce83;
  wire v8fd6c6;
  wire v8849d3;
  wire v8fd6f1;
  wire v887fec;
  wire v8fcb1c;
  wire v887c6e;
  wire v8fd570;
  wire v8fd244;
  wire v887dff;
  wire v884df7;
  wire v880750;
  wire v8fd82b;
  wire v8fd281;
  wire v88ea40;
  wire v8fd1a3;
  wire v8fd92f;
  wire v884f00;
  wire v89fb02;
  wire v8fc2d4;
  wire v8861c8;
  wire v8fd649;
  wire v88fb91;
  wire v8fd7a1;
  wire v8fd572;
  wire v8850dd;
  wire v8fd633;
  wire v8fd2d5;
  wire v887d67;
  wire v880bb6;
  wire v88318b;
  wire v885d0d;
  wire v8fd7f0;
  wire v8fd08a;
  wire v88280d;
  wire v8fd383;
  wire v885d0a;
  wire v884cea;
  wire v8818e1;
  wire v885eba;
  wire v8fc495;
  wire v885a16;
  wire v88fa9a;
  wire v8fd5d5;
  wire v86edd5;
  wire v8fd8d0;
  wire v8fd8e0;
  wire v887bbe;
  wire v88096b;
  wire v88101f;
  wire v8825fc;
  wire v8878bd;
  wire v8b5fc7;
  wire v8fd236;
  wire v8fd930;
  wire v8dac5d;
  wire v8fd255;
  wire v8fd6a7;
  wire v884c5a;
  wire v8daba0;
  wire v8fd1fe;
  wire v884da1;
  wire v884464;
  wire v890ce6;
  wire v8844ce;
  wire v8829eb;
  wire v883046;
  wire v88774e;
  wire v8fd209;
  wire v8fd6a1;
  wire v88795b;
  wire v8878c8;
  wire v88068f;
  wire v859713;
  wire v8fce7b;
  wire v8fd965;
  wire v8838c5;
  wire v882788;
  wire v8ed953;
  wire v884136;
  wire v8fd36d;
  wire v866229;
  wire v88294d;
  wire v8c2eb0;
  wire v8840e1;
  wire v8b5fca;
  wire v88580d;
  wire v8fd665;
  wire v884329;
  wire v858564;
  wire v858acb;
  wire v8fd7a7;
  wire v885947;
  wire v8fd95d;
  wire v8fc1fa;
  wire v8583a8;
  wire v882de0;
  wire v880626;
  wire v854c61;
  wire v8809df;
  wire v8fc644;
  wire v894671;
  wire v8877fe;
  wire v8fd7ca;
  wire v8fd7be;
  wire v8dad1a;
  wire v8fd6d4;
  wire v8fd5c7;
  wire v887c1e;
  wire v844fa0;
  wire v8fd17e;
  wire v8fd816;
  wire v8861f9;
  wire v885fb3;
  wire v8816ff;
  wire v8fcd29;
  wire v844f9e;
  wire v881099;
  wire v8c48b7;
  wire v8fd790;
  wire v8fd484;
  wire v881649;
  wire v8fd5d7;
  wire v8fd68b;
  wire v87bbad;
  wire v88496c;
  wire v887d06;
  wire v88254d;
  wire v887a7c;
  wire v844fbb;
  wire v895d16;
  wire v8c48b2;
  wire v844fbf;
  wire v8fd886;
  wire v8fd869;
  wire v884842;
  wire v858a41;
  wire v889757;
  wire v884735;
  wire v8fd877;
  wire v8a8729;
  wire v887cd8;
  wire v8fd72c;
  wire v887c95;
  wire v8fd467;
  wire v8587ba;
  wire v8ac1fa;
  wire v844fab;
  wire v8fd72b;
  wire v882c16;
  wire v88394f;
  wire v8880da;
  wire v8fd918;
  wire v882db5;
  wire v8810f4;
  wire v887ad9;
  wire v8fd7c2;
  wire v884a73;
  wire v8fd4f0;
  wire v87734f;
  wire v880f23;
  wire v882c83;
  wire v8dacfe;
  wire v887abd;
  wire v87949d;
  wire v8fd736;
  wire v880c4c;
  wire v8fd907;
  wire v8fd768;
  wire v882c78;
  wire v882186;
  wire v8827e5;
  wire v8fd85c;
  wire v881982;
  wire v88567a;
  wire v8fcbe3;
  wire v868a24;
  wire v8fd79f;
  wire v891b69;
  wire v883f96;
  wire v8fd242;
  wire v85f322;
  wire v892c49;
  wire v8ed1d1;
  wire v8fd51b;
  wire v8fd661;
  wire v8fd770;
  wire v880a3a;
  wire v8f29ed;
  wire v885215;
  wire v85397b;
  wire v8fd6c2;
  wire v884d11;
  wire v8fd296;
  wire v8fd957;
  wire v890cdc;
  wire v881ee1;
  wire v885d67;
  wire v87adc8;
  wire v884262;
  wire v88407b;
  wire v8fcf21;
  wire v854139;
  wire v880752;
  wire v8fd5b2;
  wire v88a4a0;
  wire v887b46;
  wire v8fd696;
  wire v88e5f1;
  wire v884577;
  wire v887b68;
  wire v884448;
  wire v8824d8;
  wire v885cc5;
  wire v894e08;
  wire v881ef6;
  wire v8880d8;
  wire v88313d;
  wire v882ea3;
  wire v8fce5e;
  wire v88083d;
  wire v881944;
  wire v8fd63e;
  wire v8a7085;
  wire v8ed1d8;
  wire v8881bd;
  wire v8ce0f4;
  wire v8fd7e4;
  wire v879433;
  wire v858ace;
  wire v8fd65f;
  wire v88454a;
  wire v8809eb;
  wire v88506d;
  wire v887ca3;
  wire v8fd714;
  wire v8fd752;
  wire v8587ee;
  wire v883928;
  wire v8fd7b5;
  wire v8fd64a;
  wire v8fd8ed;
  wire v881faf;
  wire v882f72;
  wire v88275b;
  wire v8fd958;
  wire v8fc296;
  wire v8fcc49;
  wire v8fce9e;
  wire v883c09;
  wire v895abe;
  wire v882d68;
  wire v8fd79b;
  wire v882402;
  wire v8a8783;
  wire v8fd857;
  wire v8fd7a5;
  wire v8fd8c9;
  wire v8fd1f8;
  wire v884292;
  wire v887fc7;
  wire v88fc7a;
  wire v8fd799;
  wire v8d4782;
  wire v8fd7b1;
  wire v8878e0;
  wire v880769;
  wire v8fd651;
  wire v8cd9ef;
  wire v880660;
  wire v8fd7f7;
  wire v8fd15f;
  wire v883b45;
  wire v8877a0;
  wire v8843d0;
  wire v882214;
  wire v8fd002;
  wire v885ab0;
  wire v882e12;
  wire v8fd1a0;
  wire v8fd64c;
  wire v8fd80f;
  wire v8fd1b9;
  wire v89475e;
  wire v882093;
  wire v8827ac;
  wire v880240;
  wire v88100b;
  wire v8fd182;
  wire v887f32;
  wire v895d18;
  wire v89243a;
  wire v88499a;
  wire v8fd29a;
  wire v87feab;
  wire v8844a9;
  wire v8fd71b;
  wire v8821d3;
  wire v89476c;
  wire v8879ab;
  wire v8fd1bd;
  wire v887ac6;
  wire v8f2a2c;
  wire v8fc970;
  wire v88783d;
  wire v85b247;
  wire v88186f;
  wire v887657;
  wire v858a9b;
  wire v8ed18b;
  wire v884cc3;
  wire v8ad08b;
  wire v8fd77a;
  wire v8594cb;
  wire v883c24;
  wire v8821e0;
  wire v880ac4;
  wire v88d4df;
  wire v895afe;
  wire v882b4a;
  wire v884718;
  wire v881022;
  wire v883050;
  wire v8fd8f6;
  wire v883158;
  wire v8810ca;
  wire v8fd6b5;
  wire v8fd1d0;
  wire v882302;
  wire v884953;
  wire v8858bb;
  wire v8880e4;
  wire v844fb3;
  wire v859c5b;
  wire v858acd;
  wire v8b5ff4;
  wire v8f2a80;
  wire v881018;
  wire v87dfe7;
  wire v8fcf97;
  wire v8743a1;
  wire v8fcb01;
  wire v8fd6f7;
  wire v8842de;
  wire v880263;
  wire v8fd23a;
  wire v86e414;
  wire v8fd65b;
  wire v884a25;
  wire v8fcd77;
  wire v885f1e;
  wire v8fc844;
  wire v882f33;
  wire v885b21;
  wire v882699;
  wire v883b18;
  wire v8807a6;
  wire v8fc18e;
  wire v885b36;
  wire v884d47;
  wire v879581;
  wire v885d66;
  wire v8fccac;
  wire v882b84;
  wire v880e0b;
  wire v887de8;
  wire v8810bc;
  wire v8fca7a;
  wire v885692;
  wire v8fd608;
  wire v8fcd8f;
  wire v882b41;
  wire v87bba1;
  wire v8fce87;
  wire v8fd740;
  wire v8fc484;
  wire v8fd63d;
  wire v8fd6db;
  wire v88e43b;
  wire v88235e;
  wire v8fd5f5;
  wire v882719;
  wire v8947e2;
  wire v887b69;
  wire v88770c;
  wire v8fc85b;
  wire v89fb26;
  wire v8806f0;
  wire v885d03;
  wire v887827;
  wire v8fce6a;
  wire v89faf7;
  wire v883e92;
  wire v8fd7d5;
  wire v8ad009;
  wire v8fd90b;
  wire v8946de;
  wire v8fd5c8;
  wire v8fd859;
  wire v8fd631;
  wire v8830bf;
  wire v880f35;
  wire v885beb;
  wire v887f67;
  wire v8ed93d;
  wire v8fd669;
  wire v8859f1;
  wire v882048;
  wire v8fd1dd;
  wire v8fd80d;
  wire v882569;
  wire v880bc8;
  wire v881f4a;
  wire v8f2a14;
  wire v8fd77e;
  wire v8fd1e9;
  wire v884d53;
  wire v884143;
  wire v8fd428;
  wire v880cd6;
  wire v882fd7;
  wire v88785b;
  wire v8fd1ba;
  wire v88234f;
  wire v8857e9;
  wire v8fd7c9;
  wire v89737b;
  wire v8f2a0b;
  wire v885119;
  wire v8fd5f6;
  wire v8fd349;
  wire v880638;
  wire v887627;
  wire v8860d7;
  wire v85b93e;
  wire v8dac53;
  wire v8fd5ae;
  wire v8fd358;
  wire v87bb5f;
  wire v8fd176;
  wire v887d22;
  wire v8847d3;
  wire v8fcfa9;
  wire v8586ec;
  wire v8fd641;
  wire v8fd75b;
  wire v882fd1;
  wire v8896fc;
  wire v8a707e;
  wire v884dca;
  wire v879434;
  wire v89830f;
  wire v888015;
  wire v8fce12;
  wire v8fd1bb;
  wire v8c2de8;
  wire v8821dc;
  wire v8fd683;
  wire v8818fb;
  wire v8881d6;
  wire v895a9c;
  wire v8fd232;
  wire v8dac0f;
  wire v8770c9;
  wire v8fd808;
  wire v884147;
  wire v892c5b;
  wire v880834;
  wire v882908;
  wire v8fd1e0;
  wire v8fd5e0;
  wire v8fc6b2;
  wire v8ce0f7;
  wire v885f7b;
  wire v8c008e;
  wire v8fd90d;
  wire v8fd852;
  wire v8fd035;
  wire v8587eb;
  wire v882ac1;
  wire v876f96;
  wire v883c1a;
  wire v8fc193;
  wire v8896a5;
  wire v8fd84a;
  wire v8fd823;
  wire v88595e;
  wire v8946bb;
  wire v8fce77;
  wire v8fd22e;
  wire v8fcfe8;
  wire v8947b9;
  wire v880648;
  wire v8806a9;
  wire v8fd87b;
  wire v8fd7de;
  wire v880bb1;
  wire v880643;
  wire v8fd7ee;
  wire v88258c;
  wire v8802a4;
  wire v882841;
  wire v8948bb;
  wire v895cb4;
  wire v8c2e6b;
  wire v895cb0;
  wire v8fcabb;
  wire v887656;
  wire v8846bb;
  wire v8c2ef2;
  wire v844fad;
  wire v8fd20b;
  wire v8846ba;
  wire v8fc5ad;
  wire v8861ed;
  wire v886129;
  wire v8817a3;
  wire v880341;
  wire v8f2aa3;
  wire v8fd5c4;
  wire v882490;
  wire v88380c;
  wire v887cf6;
  wire v8f29e2;
  wire v8ed983;
  wire v8fcd00;
  wire v884b64;
  wire v8861df;
  wire v880a2a;
  wire v885963;
  wire v887d93;
  wire v8fd24b;
  wire v8fd629;
  wire v8fd23f;
  wire v8fc934;
  wire v8fd744;
  wire v8847a4;
  wire v8fd729;
  wire v884d32;
  wire v87bb4b;
  wire v8fd853;
  wire v883fd7;
  wire v868e18;
  wire v897377;
  wire v8fca05;
  wire v888205;
  wire v8860a7;
  wire v8ce142;
  wire v8a8786;
  wire v8fcaa8;
  wire v885063;
  wire v888056;
  wire v881fdc;
  wire v8825d5;
  wire v8fd795;
  wire v892156;
  wire v8824ae;
  wire v8fd7b6;
  wire v8fc8a5;
  wire v88055d;
  wire v883f8f;
  wire v8fd871;
  wire v8fcbd7;
  wire v8fd717;
  wire v8fd926;
  wire v887adf;
  wire v8a0a29;
  wire v880294;
  wire v883890;
  wire v8fc2dd;
  wire v8fd969;
  wire v885c76;
  wire v8fd1c5;
  wire v8861c0;
  wire v8fc48c;
  wire v8fd68d;
  wire v8879a7;
  wire v883719;
  wire v8fcff6;
  wire v8811ad;
  wire v8fc802;
  wire v885f5a;
  wire v8fd659;
  wire v88295b;
  wire v8848b0;
  wire v8fd7d4;
  wire v888046;
  wire v87d828;
  wire v8fd599;
  wire v8fd8d6;
  wire v880b75;
  wire v883cd2;
  wire v882300;
  wire v887a17;
  wire v887fc2;
  wire v8dace1;
  wire v885ee9;
  wire v8808da;
  wire v883c0c;
  wire v8829ee;
  wire v88fdb7;
  wire v85879a;
  wire v8fd478;
  wire v8fd88e;
  wire v8fd180;
  wire v885b81;
  wire v8fd8b8;
  wire v881048;
  wire v8fd6c1;
  wire v8fd868;
  wire v8fd6b4;
  wire v884ada;
  wire v897386;
  wire v8fc246;
  wire v88b623;
  wire v887cde;
  wire v883d79;
  wire v887f3f;
  wire v8fd5fa;
  wire v88ed82;
  wire v88486a;
  wire v885931;
  wire v8fd70b;
  wire v8fc68f;
  wire v888a80;
  wire v88436d;
  wire v8831a1;
  wire v8818d7;
  wire v86ef5c;
  wire v880f84;
  wire v8820a0;
  wire v89dbce;
  wire v882ea6;
  wire v882bf5;
  wire v891e93;
  wire v8fce85;
  wire v8cd9e5;
  wire v881e54;
  wire v8a0b36;
  wire v883a3f;
  wire v8fc67a;
  wire v881f75;
  wire v8fd829;
  wire v887a90;
  wire v887c60;
  wire v883aae;
  wire v8fd7ed;
  wire v883c46;
  wire v8fd936;
  wire v8dabdf;
  wire v8fd955;
  wire v89463b;
  wire v8ad131;
  wire v884258;
  wire v8ce14d;
  wire v887f2c;
  wire v8fd81c;
  wire v8fd19d;
  wire v8588b8;
  wire v895cec;
  wire v8fd571;
  wire v88366d;
  wire v8ed1e2;
  wire v885ee1;
  wire v8859bf;
  wire v8fd847;
  wire v8fd234;
  wire v88f395;
  wire v8773cf;
  wire v8ed1ce;
  wire v88e3ec;
  wire v8819df;
  wire v880af8;
  wire v886012;
  wire v8fd747;
  wire v8fd218;
  wire v887baf;
  wire v8fd55c;
  wire v8fcc72;
  wire v8948c2;
  wire v887b03;
  wire v8fc1fe;
  wire v8851ef;
  wire v8fc1dc;
  wire v8fd78d;
  wire v8fc5e1;
  wire v88383e;
  wire v8fc938;
  wire v87948e;
  wire v884b4e;
  wire v8859af;
  wire v8fd611;
  wire v88588a;
  wire v8795c1;
  wire v884904;
  wire v8ac9cb;
  wire v8fd865;
  wire v888096;
  wire v8fc6fe;
  wire v884565;
  wire v8818e8;
  wire v8fc692;
  wire v8fd66a;
  wire v880816;
  wire v8f1f45;
  wire v884034;
  wire v8fcedb;
  wire v887c98;
  wire v8fd54b;
  wire v8fc8ca;
  wire v883677;
  wire v8fcd0e;
  wire v889be1;
  wire v881e44;
  wire v895ce3;
  wire v887a69;
  wire v8ed1c6;
  wire v8fd284;
  wire v887bef;
  wire v8fd6aa;
  wire v885144;
  wire v8fd538;
  wire v8fd5ea;
  wire v8827ef;
  wire v8c2de5;
  wire v8fc7b1;
  wire v881a1a;
  wire v87dfc7;
  wire v8fd1d6;
  wire v8fd4e0;
  wire v894924;
  wire v884d85;
  wire v8858e2;
  wire v887629;
  wire v8fd1db;
  wire v88108f;
  wire v8843b6;
  wire v883f84;
  wire v8fcba4;
  wire v89fb46;
  wire v8fc9d9;
  wire v8fd6a0;
  wire v8802a2;
  wire v8fcd75;
  wire v890fe3;
  wire v8fd88d;
  wire v8940fc;
  wire v887aee;
  wire v8818f6;
  wire v880d6b;
  wire v883968;
  wire v8846fc;
  wire v895a39;
  wire v8803e6;
  wire v8569e0;
  wire v887c9a;
  wire v8fd1ca;
  wire v880821;
  wire v883de0;
  wire v8859d2;
  wire v882024;
  wire v8972bc;
  wire v8fd5fc;
  wire v884941;
  wire v8828f5;
  wire v895d4b;
  wire v8972ae;
  wire v8fd18f;
  wire v881985;
  wire v8fd65e;
  wire v8dacc2;
  wire v883bef;
  wire v8fd903;
  wire v854830;
  wire v882673;
  wire v895a71;
  wire v88d29b;
  wire v880507;
  wire v884bdc;
  wire v885a06;
  wire v88e73e;
  wire v882bb8;
  wire v8fc5a3;
  wire v8fd011;
  wire v8861bc;
  wire v88417e;
  wire v8fd2f7;
  wire v885102;
  wire v885b44;
  wire v883837;
  wire v881e33;
  wire v8fd637;
  wire v8ad079;
  wire v890631;
  wire v8dad14;
  wire v882910;
  wire v8810d4;
  wire v880a70;
  wire v8fc679;
  wire v884ccb;
  wire v891594;
  wire v897303;
  wire v881720;
  wire v88391f;
  wire v884afb;
  wire v885d0f;
  wire v884f6d;
  wire v883b53;
  wire v8584ff;
  wire v898e5c;
  wire v887f4e;
  wire v887a7a;
  wire v86b3d4;
  wire v8fd96b;
  wire v8ad12a;
  wire v8fd56f;
  wire v8845a2;
  wire v8fd60b;
  wire v880d42;
  wire v8816ab;
  wire v887c6c;
  wire v8fd794;
  wire v8849ca;
  wire v8fd150;
  wire v887a7f;
  wire v8839ba;
  wire v860216;
  wire v882cf9;
  wire v88f397;
  wire v881117;
  wire v8fd6de;
  wire v8827e6;
  wire v8fc6ea;
  wire v885b62;
  wire v874ed6;
  wire v883eb1;
  wire v858422;
  wire v8fd579;
  wire v8fd68f;
  wire v8fd5cc;
  wire v880d40;
  wire v8fd5d4;
  wire v88315b;
  wire v88e6e1;
  wire v86ef60;
  wire v8806a6;
  wire v883d20;
  wire v8c98e7;
  wire v8fc4c0;
  wire v8fcc62;
  wire v8fd6bf;
  wire v887d9c;
  wire v8fd83c;
  wire v87bb76;
  wire v8fd966;
  wire v8fd5e2;
  wire v8fd96a;
  wire v88442a;
  wire v8b606c;
  wire v8946a5;
  wire v888162;
  wire v887a00;
  wire v8845a8;
  wire v883833;
  wire v88fbd1;
  wire v880b8e;
  wire v887868;
  wire v8a704c;
  wire v885a43;
  wire v88769d;
  wire v883781;
  wire v880804;
  wire v882e16;
  wire v88426c;
  wire v8fc606;
  wire v8fd623;
  wire v885c69;
  wire v88579e;
  wire v8fd7a8;
  wire v895c60;
  wire v8827b2;
  wire v887b5a;
  wire v8805c4;
  wire v887f56;
  wire v87eaaf;
  wire v8881d4;
  wire v8ad053;
  wire v8fd7aa;
  wire v8fd851;
  wire v883035;
  wire v884867;
  wire v883d66;
  wire v8fd950;
  wire v8fd25a;
  wire v8844d6;
  wire v8fd556;
  wire v8830a2;
  wire v8fd1d9;
  wire v8fd57a;
  wire v8fce04;
  wire v8fd8db;
  wire v8fd2cf;
  wire v8ad133;
  wire v887768;
  wire v8fd8f4;
  wire v885d08;
  wire v889498;
  wire v8b5feb;
  wire v880614;
  wire v8fd196;
  wire v8f2a5a;
  wire v885f69;
  wire v8fd8a2;
  wire v88174e;
  wire v8fd17d;
  wire v8fd1c7;
  wire v88478b;
  wire v884cad;
  wire v884a6e;
  wire v8fd5a2;
  wire v8fd657;
  wire v8fd788;
  wire v8fd5a8;
  wire v8587bf;
  wire v880e00;
  wire v885a6c;
  wire v844fb5;
  wire v888182;
  wire v885b89;
  wire v8fd186;
  wire v884170;
  wire v8fd951;
  wire v8ce111;
  wire v8878ac;
  wire v858796;
  wire v880323;
  wire v8fcf25;
  wire v8860bd;
  wire v88310a;
  wire v8829b5;
  wire v88118b;
  wire v8fd341;
  wire v8836e8;
  wire v88fdb8;
  wire v8fd6ae;
  wire v8896ed;
  wire v880c0e;
  wire v8897a6;
  wire v887644;
  wire v8e1d28;
  wire v8fd455;
  wire v884482;
  wire v883d05;
  wire v882a64;
  wire v894850;
  wire v880565;
  wire v8fd7a4;
  wire v883f7a;
  wire v8974c9;
  wire v8ce1ae;
  wire v8dab99;
  wire v88f0b3;
  wire v8fd686;
  wire v88232b;
  wire v8fd82a;
  wire v87ff04;
  wire v895a65;
  wire v8b78a2;
  wire v884359;
  wire v8fd6c3;
  wire v88793c;
  wire v875cbc;
  wire v882905;
  wire v885909;
  wire v8820ed;
  wire v890fd8;
  wire v88319e;
  wire v8fd174;
  wire v8dac2c;
  wire v8fd8e4;
  wire v88079c;
  wire v8fd64d;
  wire v888bbe;
  wire v888a7f;
  wire v8c2ed0;
  wire v8fd90e;
  wire v887f88;
  wire v8820d8;
  wire v89fb1c;
  wire v895bb6;
  wire v88369f;
  wire v8fc719;
  wire v8822fe;
  wire v885dc6;
  wire v8b5ff5;
  wire v89736f;
  wire v8fd872;
  wire v881975;
  wire v8809d1;
  wire v882772;
  wire v884cde;
  wire v8fd6e6;
  wire v8fcf73;
  wire v8ce1b0;
  wire v8fd91d;
  wire v87001c;
  wire v8841cd;
  wire v8fd896;
  wire v8fc9c2;
  wire v8947ee;
  wire v8fd7f2;
  wire v883a54;
  wire v8fd6d9;
  wire v880d9a;
  wire v88251a;
  wire v8856e4;
  wire v885d31;
  wire v8fd5b0;
  wire v887881;
  wire v894722;
  wire v8fce28;
  wire v8fd69d;
  wire v884d3b;
  wire v884585;
  wire v882d42;
  wire v8fc9fd;
  wire v884984;
  wire v8fd6e0;
  wire v8802ff;
  wire v8fd6d1;
  wire v88786b;
  wire v895c31;
  wire v8fd913;
  wire v880620;
  wire v8ed1d3;
  wire v880236;
  wire v884626;
  wire v8a87bc;
  wire v8fd8eb;
  wire v890cff;
  wire v8fd923;
  wire v88ec29;
  wire v8fd627;
  wire v8fd843;
  wire v882a37;
  wire v88bb79;
  wire v8fd92a;
  wire v87feba;
  wire v8894e3;
  wire v8fd7b2;
  wire v887d8f;
  wire v8fcd6f;
  wire v8762d1;
  wire v88376e;
  wire v8823c2;
  wire v8830c5;
  wire v88ea59;
  wire v8fd914;
  wire v883e2e;
  wire v8fc5c1;
  wire v8fd876;
  wire v854a91;
  wire v882e65;
  wire v8fd51f;
  wire v88bb4f;
  wire v895b58;
  wire v882764;
  wire v883c06;
  wire v88e1fb;
  wire v883071;
  wire v882bb2;
  wire v8837fe;
  wire v887c92;
  wire v85bfad;
  wire v8fd24a;
  wire v8fd25d;
  wire v8fd594;
  wire v8fd215;
  wire v886188;
  wire v888143;
  wire v8fd705;
  wire v8fc42f;
  wire v8879a4;
  wire v8810de;
  wire v87bacb;
  wire v882bee;
  wire v8fd3c8;
  wire v887ce9;
  wire v882b96;
  wire v881e4b;
  wire v8fd18b;
  wire v880d0c;
  wire v8f2abb;
  wire v884036;
  wire v88602f;
  wire v8fd1d2;
  wire v8642ea;
  wire v8fd83b;
  wire v8848a0;
  wire v8ed1b3;
  wire v8896c7;
  wire v8fcb09;
  wire v887d31;
  wire v8dac95;
  wire v8fd850;
  wire v8fc1cd;
  wire v8fd726;
  wire v86bd4d;
  wire v881edd;
  wire v8fd183;
  wire v8fd8fa;
  wire v8fcfaa;
  wire v8fd2a3;
  wire v8fc8f1;
  wire v8fd5ac;
  wire v885149;
  wire v8fd842;
  wire v883f9f;
  wire v88514d;
  wire v8f2a50;
  wire v887cca;
  wire v8fd20a;
  wire v88777d;
  wire v887846;
  wire v8fd5f9;
  wire v882e37;
  wire v8fc98c;
  wire v8fd693;
  wire v8fd662;
  wire v8fc708;
  wire v881963;
  wire v884539;
  wire v8fd6a9;
  wire v890fdd;
  wire v8fd7f4;
  wire v88e2ce;
  wire v86deca;
  wire v8fd7fd;
  wire v8fca66;
  wire v8fd597;
  wire v8fd8d5;
  wire v8881e7;
  wire v8910ad;
  wire v883012;
  wire v882217;
  wire v8fc1bf;
  wire v8881f0;
  wire v8fd773;
  wire v8fc61c;
  wire v87945a;
  wire v88306a;
  wire v88390f;
  wire v882603;
  wire v88212e;
  wire v8fd793;
  wire v8843ba;
  wire v884013;
  wire v885026;
  wire v883e11;
  wire v885fb8;
  wire v89726c;
  wire v8808cf;
  wire v884a26;
  wire v8fd20f;
  wire v8fd689;
  wire v8fd612;
  wire v88589c;
  wire v885d73;
  wire v8856c1;
  wire v884d5a;
  wire v8fd5dd;
  wire v8c4d03;
  wire v8881be;
  wire v8847e5;
  wire v8fd805;
  wire v8fd5a4;
  wire v880b07;
  wire v8fd713;
  wire v8c0098;
  wire v887aed;
  wire v8fcdd5;
  wire v883089;
  wire v87b4e7;
  wire v8a87b9;
  wire v884fa4;
  wire v8587e6;
  wire v885ddd;
  wire v895b0b;
  wire v884920;
  wire v882484;
  wire v883e1c;
  wire v8826ea;
  wire v8fd836;
  wire v8fd5d2;
  wire v8fd59f;
  wire v8fc942;
  wire v854d37;
  wire v8989c5;
  wire v896f10;
  wire v8818b7;
  wire v88a2de;
  wire v884d5e;
  wire v8fd60e;
  wire v88259e;
  wire v8fd82e;
  wire v88ec23;
  wire v8808c9;
  wire v8fd860;
  wire v8f2a18;
  wire v8837de;
  wire v8fd113;
  wire v887ccd;
  wire v8805b9;
  wire v8886e1;
  wire v8b5fc6;
  wire v8838cd;
  wire v8fd80a;
  wire v8c2ebb;
  wire v8805d7;
  wire v8fd928;
  wire v8fd761;
  wire v8b60d1;
  wire v8816cc;
  wire v88023c;
  wire v890d28;
  wire v8fc2e5;
  wire v8fd688;
  wire v8847e2;
  wire v8fccad;
  wire v8ad0c2;
  wire v88112f;
  wire v88fd1c;
  wire v8cd9cd;
  wire v8fd1a4;
  wire v8fd039;
  wire v88085d;
  wire v8805dc;
  wire v880db3;
  wire v89488c;
  wire v887a4a;
  wire v883cd1;
  wire v8fd8b2;
  wire v88791d;
  wire v8fc57a;
  wire v8fd8a0;
  wire v8cadd9;
  wire v88ec21;
  wire v8fd77d;
  wire v8fd7c3;
  wire v8b5ffa;
  wire v8fd1e7;
  wire v8822cf;
  wire v898e61;
  wire v8fd1a6;
  wire v881ec5;
  wire v8816aa;
  wire v87102d;
  wire v881657;
  wire v8811b3;
  wire v880e69;
  wire v884e03;
  wire v885e81;
  wire v882852;
  wire v882c30;
  wire v8b6054;
  wire v8fd58f;
  wire v88397a;
  wire v8fd256;
  wire v8fc945;
  wire v880e10;
  wire v885f4a;
  wire v887887;
  wire v8fd920;
  wire v8fd59c;
  wire v8fc9ca;
  wire v8fd7ac;
  wire v8fd7fc;
  wire v8fd5db;
  wire v8fd880;
  wire v8fc5f2;
  wire v87fe68;
  wire v8fce5c;
  wire v8fd251;
  wire v88064f;
  wire v895d15;
  wire v882b76;
  wire v884035;
  wire v8fd6be;
  wire v89241d;
  wire v8fd22a;
  wire v8fd84d;
  wire v8856f6;
  wire v880eda;
  wire v8fd12b;
  wire v882d74;
  wire v887f83;
  wire v897323;
  wire v8c4d0d;
  wire v887efe;
  wire v88599b;
  wire v884bdd;
  wire v885fbe;
  wire v8fd452;
  wire v8fccd5;
  wire v85841e;
  wire v882e64;
  wire v887d0a;
  wire v8fd8d7;
  wire v8fd222;
  wire v883e34;
  wire v8fcb76;
  wire v8fcac6;
  wire v883c78;
  wire v8fd5f7;
  wire v885b3a;
  wire v8f2a7d;
  wire v894703;
  wire v886197;
  wire v8fd8fb;
  wire v8fd7e7;
  wire v8fc76f;
  wire v895ce5;
  wire v8ed1ca;
  wire v884782;
  wire v884875;
  wire v8fc67f;
  wire v8fd8c4;
  wire v8fd18e;
  wire v8843ae;
  wire v8fcf10;
  wire v8fd598;
  wire v892325;
  wire v8fd6bd;
  wire v8fd19f;
  wire v8fd863;
  wire v88604b;
  wire v8fd929;
  wire v887fe2;
  wire v89fb88;
  wire v8fd833;
  wire v8fd3fc;
  wire v8fd7f3;
  wire v883b2a;
  wire v8fd751;
  wire v8a7063;
  wire v8fd89a;
  wire v88574b;
  wire v8fd6e1;
  wire v8fd6e2;
  wire v8846f7;
  wire v8fc325;
  wire v8878c5;
  wire v887bfb;
  wire v888662;
  wire v8fced0;
  wire v8859e8;
  wire v8fd648;
  wire v8fd457;
  wire v8fd8d4;
  wire v8877c5;
  wire v8fd837;
  wire v88305d;
  wire v887cfa;
  wire v883cfc;
  wire v8fca32;
  wire v880741;
  wire v8fd614;
  wire v8947ed;
  wire v8fd62f;
  wire v88367e;
  wire v8fc6aa;
  wire v895b2f;
  wire v8fd2b7;
  wire v882034;
  wire v8825da;
  wire v881141;
  wire v885684;
  wire v8fcecd;
  wire v8fd733;
  wire v8f2a57;
  wire v8fd91a;
  wire v8fcfce;
  wire v894637;
  wire v887ade;
  wire v8fc801;
  wire v8ac9b2;
  wire v88bc54;
  wire v8fc64f;
  wire v8fd846;
  wire v88498b;
  wire v885ea9;
  wire v8c2e51;
  wire v885ab1;
  wire v8fd6d0;
  wire v88c103;
  wire v8f29e5;
  wire v887ac3;
  wire v8fd654;
  wire v8fd701;
  wire v8ad05f;
  wire v85fc7a;
  wire v8850e9;
  wire v8fd609;
  wire v8fd685;
  wire v8a88d5;
  wire v8fce1f;
  wire v882507;
  wire v8a70a6;
  wire v885e84;
  wire v88241f;
  wire v870c76;
  wire v8807d3;
  wire v87bb66;
  wire v8fd73a;
  wire v8fd8ba;
  wire v88493b;
  wire v89726a;
  wire v8ad097;
  wire v894dfc;
  wire v8fd73b;
  wire v8fd4e2;
  wire v884bc5;
  wire v882bc8;
  wire v8fd6ab;
  wire v8fd5e3;
  wire v8896fd;
  wire v884a6d;
  wire v8fd666;
  wire v887966;
  wire v854ae6;
  wire v8823f5;
  wire v8fd1fd;
  wire v884747;
  wire v8fd63f;
  wire v8fd5b4;
  wire v8fd7dc;
  wire v8fce55;
  wire v8fd939;
  wire v885b87;
  wire v8f2aa5;
  wire v8841bc;
  wire v885df9;
  wire v8fcd1f;
  wire v890676;
  wire v8939a7;
  wire v880544;
  wire v8fd238;
  wire v887879;
  wire v8fc9d3;
  wire v88fbfc;
  wire v8fd85b;
  wire v864119;
  wire v8fc5a6;
  wire v887c44;
  wire v885de9;
  wire v88fb6f;
  wire v880487;
  wire v8857aa;
  wire v8850ab;
  wire v8805ad;
  wire v885fce;
  wire v880231;
  wire v8fd6bc;
  wire v88fcc8;
  wire v882d0f;
  wire v8fd742;
  wire v885d65;
  wire v897301;
  wire v87debc;
  wire v8fd5fd;
  wire v8915ef;
  wire v8fd5d6;
  wire v87ff08;
  wire v8fcfc3;
  wire v882170;
  wire v8b60af;
  wire v8b603b;
  wire v8fd574;
  wire v8fd8aa;
  wire v884316;
  wire v8ce18c;
  wire v8fd6a8;
  wire v8fd239;
  wire v894721;
  wire v885ea3;
  wire v8fd195;
  wire v8fd8ea;
  wire v8fd716;
  wire v880674;
  wire v882a2c;
  wire v885748;
  wire v885bee;
  wire v869327;
  wire v8fd214;
  wire v854bab;
  wire v8fd584;
  wire v88284b;
  wire v8fc8d5;
  wire v88ed0c;
  wire v8823a0;
  wire v884bcc;
  wire v8fd84f;
  wire v8fd6c9;
  wire v8fd577;
  wire v8840d5;
  wire v8fd8c1;
  wire v8fd64f;
  wire v895a56;
  wire v880763;
  wire v884f81;
  wire v882bbf;
  wire v88170c;
  wire v884870;
  wire v882f45;
  wire v8fd536;
  wire v8fd1aa;
  wire v880eac;
  wire v880d66;
  wire v8d4e0d;
  wire v8fd87d;
  wire v885bf2;
  wire v884b83;
  wire v8fc9f1;
  wire v88237c;
  wire v884f8e;
  wire v8fc28a;
  wire v869e2c;
  wire v894828;
  wire v885e9f;
  wire v8fd5ee;
  wire v8fcd30;
  wire v887897;
  wire v882d73;
  wire v883a2e;
  wire v882859;
  wire v8fd7c6;
  wire v8838a3;
  wire v880f66;
  wire v8fd642;
  wire v882ae0;
  wire v8fc3cf;
  wire v8fd8c3;
  wire v880bf2;
  wire v88770f;
  wire v8850da;
  wire v880c3a;
  wire v883685;
  wire v887dae;
  wire v884907;
  wire v887d5b;
  wire v8fd5bf;
  wire v8fc7b7;
  wire v885b2d;
  wire v86ecd4;
  wire v884058;
  wire v883b0e;
  wire v87fb41;
  wire v88055f;
  wire v8840c5;
  wire v880599;
  wire v887def;
  wire v88257d;
  wire v887765;
  wire v8fd940;
  wire v8841f9;
  wire v8fc290;
  wire v88046c;
  wire v888062;
  wire v8878bb;
  wire v880b5b;
  wire v8972d7;
  wire v8d477f;
  wire v8fd602;
  wire v88810f;
  wire v8fd8b7;
  wire v880b78;
  wire v85397c;
  wire v8fd715;
  wire v8c993e;
  wire v8fd71a;
  wire v884a71;
  wire v892ca3;
  wire v882002;
  wire v89fb95;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg StoB_REQ4_p;
  input StoB_REQ4_n;
  reg StoB_REQ5_p;
  input StoB_REQ5_n;
  reg StoB_REQ6_p;
  input StoB_REQ6_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoS_ACK4_p;
  output BtoS_ACK4_n;
  reg BtoS_ACK5_p;
  output BtoS_ACK5_n;
  reg BtoS_ACK6_p;
  output BtoS_ACK6_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg SLC2_p;
  output SLC2_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  wire SLC0_n;
  wire ENQ_n;
  wire SLC2_n;

assign v8fcfce = RtoB_ACK1_p & v8f2a57 | !RtoB_ACK1_p & v8fce5c;
assign v883fd7 = StoB_REQ1_p & v88eb82 | !StoB_REQ1_p & v844f91;
assign v8fd84a = BtoR_REQ1_p & v8896a5 | !BtoR_REQ1_p & v844f91;
assign v8fcf25 = StoB_REQ2_p & v8fd951 | !StoB_REQ2_p & v880323;
assign v8857e5 = StoB_REQ6_p & v8fcbc7 | !StoB_REQ6_p & v8878da;
assign v8fd689 = jx0_p & v88390f | !jx0_p & !v882e37;
assign v8849ca = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd794;
assign v8fd923 = StoB_REQ2_p & v8fd196 | !StoB_REQ2_p & v890cff;
assign v8fd5f5 = StoB_REQ1_p & v8fd15f | !StoB_REQ1_p & v88235e;
assign v8859d2 = stateG7_1_p & v883de0 | !stateG7_1_p & v8fc6fe;
assign v88234f = jx1_p & v880cd6 | !jx1_p & v8fd1ba;
assign v8837fe = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v882bb2;
assign v8fd296 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd1b8;
assign v8766ed = RtoB_ACK1_p & v87fed4 | !RtoB_ACK1_p & v895ceb;
assign v880d42 = BtoS_ACK1_p & v88219e | !BtoS_ACK1_p & v8fd60b;
assign v885ab0 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd002;
assign v8fcecd = RtoB_ACK0_p & v8fce5c | !RtoB_ACK0_p & v885684;
assign v88e6e1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v88315b;
assign v8fce83 = jx0_p & v8810a6 | !jx0_p & v8fce44;
assign v8fd6a6 = jx0_p & v844f9b | !jx0_p & v895d61;
assign v8fd683 = BtoS_ACK0_p & v8a707e | !BtoS_ACK0_p & v8821dc;
assign v844fad = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v885f5a = jx1_p & v8811ad | !jx1_p & !v8fc802;
assign v8fd58e = jx1_p & v8dabff | !jx1_p & v883fee;
assign v8fd917 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd6a5;
assign v884767 = BtoS_ACK0_p & v88402c | !BtoS_ACK0_p & v881630;
assign v884049 = EMPTY_p & v8b6045 | !EMPTY_p & !v8fd848;
assign v8fd895 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & !v8822d4;
assign v8ac9bd = BtoS_ACK0_p & v8fd70d | !BtoS_ACK0_p & v8859ec;
assign v895b93 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd83e;
assign v884d49 = StoB_REQ2_p & v8fd895 | !StoB_REQ2_p & v844f91;
assign v885d25 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v88367e = BtoR_REQ1_p & v8816aa | !BtoR_REQ1_p & v8fd62f;
assign v8fd65b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86e414;
assign v8fd87f = StoB_REQ6_p & v8fc2e4 | !StoB_REQ6_p & v88579b;
assign v884d94 = jx0_p & v885ec1 | !jx0_p & !v89735b;
assign v882d8f = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v844f91;
assign v8fd1de = EMPTY_p & v8fd231 | !EMPTY_p & v880952;
assign v887b5e = jx2_p & v882e00 | !jx2_p & v8fd596;
assign v8841f9 = jx1_p & v8fd940 | !jx1_p & !v844f91;
assign v8fd5a5 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v853f4e;
assign v887f4e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v898e5c;
assign v8830bf = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8fd1b9;
assign v8946de = RtoB_ACK0_p & v880e0b | !RtoB_ACK0_p & v8fd90b;
assign v8806a9 = RtoB_ACK1_p & v8947b9 | !RtoB_ACK1_p & v844f91;
assign v8fd63d = RtoB_ACK0_p & v880e0b | !RtoB_ACK0_p & v8fc484;
assign v87948e = RtoB_ACK0_p & v887baf | !RtoB_ACK0_p & v8fc938;
assign v882f33 = StoB_REQ1_p & v8fd15f | !StoB_REQ1_p & v8fc844;
assign v8fd163 = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v8fd587;
assign v8fc8a5 = jx1_p & v8fd795 | !jx1_p & !v8fd7b6;
assign v844fb3 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f91;
assign v8818e8 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd6b3;
assign v8fd833 = BtoS_ACK0_p & v8fd1a3 | !BtoS_ACK0_p & v89fb88;
assign v8fd966 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87bb76;
assign v8fd1d7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cecad;
assign v8dabdf = BtoS_ACK6_p & v885d25 | !BtoS_ACK6_p & !v8fd78e;
assign v8fd8df = StoB_REQ3_p & v8fc1cf | !StoB_REQ3_p & v844f9d;
assign v8fd597 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fca66;
assign v8fd7fb = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v89110a;
assign v8fd5ac = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fc8f1;
assign v88083d = stateG7_1_p & v8fce5e | !stateG7_1_p & v85f322;
assign v883bb8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v887adb;
assign v883105 = BtoS_ACK6_p & v884476 | !BtoS_ACK6_p & v8fd67e;
assign v8c993e = RtoB_ACK0_p & v88046c | !RtoB_ACK0_p & v8fd715;
assign v884d32 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd729;
assign v885fe4 = BtoS_ACK0_p & v8836c4 | !BtoS_ACK0_p & v88576c;
assign v8fd24a = StoB_REQ3_p & v88e1fb | !StoB_REQ3_p & v882673;
assign v880b56 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8850d3;
assign v8fd6b6 = RtoB_ACK1_p & v8fd812 | !RtoB_ACK1_p & v8878b5;
assign v894721 = RtoB_ACK0_p & v87bb66 | !RtoB_ACK0_p & v8fd239;
assign v8fd6fc = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8851dd;
assign v89dbce = jx0_p & v8fd926 | !jx0_p & v8820a0;
assign v8fd85c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8827e5;
assign v881ec5 = jx1_p & v844f91 | !jx1_p & !v8fd1a6;
assign v886048 = RtoB_ACK0_p & v880ed2 | !RtoB_ACK0_p & v882a0a;
assign v8fce77 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8946bb;
assign v8587ee = RtoB_ACK1_p & v88506d | !RtoB_ACK1_p & v8fd752;
assign v88784a = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v885c0e;
assign v883833 = jx2_p & v8fd6bf | !jx2_p & v8845a8;
assign v8fd704 = FULL_p & v8f2aa9 | !FULL_p & v8876bb;
assign v8fd84f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd73a;
assign v8ad12a = jx0_p & v844f9f | !jx0_p & !v8fd96b;
assign v86ed7e = BtoS_ACK0_p & v844fa1 | !BtoS_ACK0_p & !v882006;
assign v8fd8a2 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v885f69;
assign v880e79 = jx0_p & v8588b1 | !jx0_p & !v8fd8b4;
assign v887d22 = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v8fd176;
assign v8fd733 = jx1_p & v8676b7 | !jx1_p & v8fd614;
assign v8cadd9 = StoB_REQ2_p & v885909 | !StoB_REQ2_p & v8fd8a0;
assign v8ce142 = jx1_p & v880341 | !jx1_p & v8860a7;
assign v884f00 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8fd92f;
assign v8fca32 = stateG7_1_p & v883cfc | !stateG7_1_p & v8fc945;
assign v8fd6a1 = BtoR_REQ1_p & v8fd8e0 | !BtoR_REQ1_p & v8fd209;
assign v883d66 = RtoB_ACK1_p & v8fc7b1 | !RtoB_ACK1_p & v87eaaf;
assign v8a707e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd764;
assign v8859f1 = jx1_p & v887f67 | !jx1_p & v8fd669;
assign v884316 = jx2_p & v8fd8aa | !jx2_p & v87bb66;
assign v8fd847 = jx1_p & v883f8f | !jx1_p & v8859bf;
assign v8fd17e = StoB_REQ4_n & v844f91 | !StoB_REQ4_n & v844fa0;
assign v88ea5a = BtoS_ACK6_p & v885b17 | !BtoS_ACK6_p & v8fd610;
assign v8fd94b = RtoB_ACK1_p & v8f2a03 | !RtoB_ACK1_p & v8fd585;
assign v882302 = stateG7_1_p & v8fd1d0 | !stateG7_1_p & v8810ca;
assign v888bbe = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v8fd64d;
assign v8b605e = BtoS_ACK0_p & v8fd3c6 | !BtoS_ACK0_p & !v8fc2b8;
assign v883ee4 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8fd6d3;
assign v88777d = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd20a;
assign v8586ec = jx0_p & v8fd358 | !jx0_p & v8fcfa9;
assign v8743a1 = StoB_REQ0_p & v8877a0 | !StoB_REQ0_p & v8fcf97;
assign v881113 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8dac46;
assign v887f70 = EMPTY_p & v885723 | !EMPTY_p & v8fd5a1;
assign v880c8a = stateG7_1_p & v882a5a | !stateG7_1_p & v882a0a;
assign v882d42 = jx2_p & v884585 | !jx2_p & !v88793c;
assign v887c44 = StoB_REQ6_p & v892c36 | !StoB_REQ6_p & v8fd939;
assign v887f2c = jx2_p & v8ce142 | !jx2_p & v8ce14d;
assign v88810f = stateG7_1_p & v8fd602 | !stateG7_1_p & v8fc290;
assign v8fc5a6 = jx0_p & v844f91 | !jx0_p & v882bc8;
assign v887a69 = stateG12_p & v8fc6fe | !stateG12_p & v895ce3;
assign v8fc68f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8fd70b;
assign v8fd823 = BtoR_REQ0_p & v8896fc | !BtoR_REQ0_p & v8fd84a;
assign v8fc1a7 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v887d16;
assign v894b33 = stateG7_1_p & v8fd568 | !stateG7_1_p & v87fed4;
assign v864119 = jx2_p & v8fc9d3 | !jx2_p & !v8fd85b;
assign v880d9a = BtoR_REQ1_p & v8fd896 | !BtoR_REQ1_p & v8fd6d9;
assign v8842b7 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8825e5;
assign v882d74 = BtoR_REQ0_p & v8856f6 | !BtoR_REQ0_p & v8fd12b;
assign v86ed35 = jx1_p & v8fd922 | !jx1_p & !v8fd7ba;
assign v8fd744 = StoB_REQ1_p & v8fc934 | !StoB_REQ1_p & v844f91;
assign v8fcc5a = StoB_REQ6_p & v88f1b0 | !StoB_REQ6_p & v844f91;
assign v8fd1e7 = BtoS_ACK6_p & v882baa | !BtoS_ACK6_p & v8b5ffa;
assign v882093 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v89475e;
assign v8fd7a4 = StoB_REQ0_p & v8e1d28 | !StoB_REQ0_p & v880565;
assign v8fd7f4 = jx1_p & v884539 | !jx1_p & v890fdd;
assign v88772e = BtoR_REQ1_p & v8fd5e8 | !BtoR_REQ1_p & v8fd727;
assign v882569 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd80d;
assign v883781 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88769d;
assign v885b81 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd180;
assign v880e82 = StoB_REQ6_p & v853f24 | !StoB_REQ6_p & v887ad8;
assign v88602f = StoB_REQ0_p & v887ce9 | !StoB_REQ0_p & v884036;
assign v892c5b = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v884147;
assign v8a8783 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v882402;
assign v8ad0e2 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f99;
assign v858564 = RtoB_ACK1_p & v866229 | !RtoB_ACK1_p & v884329;
assign v88a2de = RtoB_ACK1_p & v894722 | !RtoB_ACK1_p & v882d42;
assign v8896a5 = stateG7_1_p & v8fc193 | !stateG7_1_p & v8fd75b;
assign v8fd150 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v887f3a;
assign v8d477f = BtoR_REQ0_p & v88055f | !BtoR_REQ0_p & v8972d7;
assign v8fd19f = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v882217;
assign v884ada = BtoS_ACK0_p & v8fd853 | !BtoS_ACK0_p & v8fd6b4;
assign v88265b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a8734;
assign v87bb4b = BtoS_ACK0_p & v8fd629 | !BtoS_ACK0_p & v884d32;
assign v880c81 = StoB_REQ6_p & v8fc78f | !StoB_REQ6_p & v8805be;
assign v887887 = jx1_p & v8676b7 | !jx1_p & v887a4a;
assign v8808c9 = RtoB_ACK0_p & v88ec23 | !RtoB_ACK0_p & v882d42;
assign v889be1 = stateG7_1_p & v8fcd0e | !stateG7_1_p & v8fc8ca;
assign v882bbf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v884f81;
assign v8fd7c6 = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v8fd92f;
assign v884782 = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v8ed1ca;
assign v8fd2d5 = StoB_REQ6_p & v88fb91 | !StoB_REQ6_p & v8fd633;
assign v885fce = BtoS_ACK6_p & v885df9 | !BtoS_ACK6_p & v8805ad;
assign v8fd1aa = stateG7_1_p & v8fd536 | !stateG7_1_p & v8fd5fd;
assign v8fc67a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v887fa9;
assign v887d85 = jx1_p & v8fd76a | !jx1_p & v88fa9e;
assign v884058 = BtoR_REQ0_p & v880eac | !BtoR_REQ0_p & v86ecd4;
assign v8fd490 = StoB_REQ6_p & v8fc729 | !StoB_REQ6_p & v8dab8a;
assign v883a54 = jx1_p & v885a6c | !jx1_p & v8fd7f2;
assign BtoS_ACK0_n = v8cd9ef;
assign v8840c5 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8850ab;
assign v887d93 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9f;
assign v895abe = jx2_p & v8fcc49 | !jx2_p & v883c09;
assign v8fd1b8 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8fd895;
assign v898f2f = stateG7_1_p & v8766ed | !stateG7_1_p & v895ceb;
assign v885fda = jx0_p & v88837d | !jx0_p & !v8fd818;
assign v8808eb = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v897cf5;
assign v8840af = StoB_REQ6_p & v8fc21f | !StoB_REQ6_p & v885b96;
assign v8861a4 = stateG7_1_p & v88565e | !stateG7_1_p & v887b5e;
assign v85f322 = jx2_p & v8fd242 | !jx2_p & v8fd79f;
assign v869327 = jx0_p & v885bee | !jx0_p & v8fd238;
assign v8fd5b4 = stateG12_p & v87bb66 | !stateG12_p & v8fd63f;
assign v88514d = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v883f9f;
assign v8fd78b = BtoS_ACK0_p & v880fd1 | !BtoS_ACK0_p & v882f43;
assign v88791d = jx1_p & v8fc1c0 | !jx1_p & !v8fd8b2;
assign v885d0f = jx0_p & v884afb | !jx0_p & v880816;
assign v8fd51b = stateG7_1_p & v8ed1d1 | !stateG7_1_p & v85f322;
assign v88299b = StoB_REQ6_p & v8fd7af | !StoB_REQ6_p & v8fd0a4;
assign v8843b6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v88108f;
assign v8fd231 = BtoR_REQ0_p & v88fc61 | !BtoR_REQ0_p & v88112b;
assign v885b17 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v882bdd;
assign v8fd1cd = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v887f13;
assign v8fd751 = RtoB_ACK1_p & v8fd6bd | !RtoB_ACK1_p & v883b2a;
assign v8fd5da = BtoS_ACK0_p & v86ed36 | !BtoS_ACK0_p & v8fd5eb;
assign v883c24 = jx2_p & v8594cb | !jx2_p & v8827ac;
assign v8fc938 = BtoR_REQ1_p & v88383e | !BtoR_REQ1_p & v8fcc72;
assign v8fd8fa = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fd183;
assign v88257d = jx0_p & v8c2eb0 | !jx0_p & v887def;
assign v8fd1f9 = StoB_REQ0_p & v8fc295 | !StoB_REQ0_p & v89386c;
assign v8fd760 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8fd830;
assign v890d28 = jx0_p & v8809c4 | !jx0_p & !v844f91;
assign v8fd6f1 = StoB_REQ6_p & v8849d3 | !StoB_REQ6_p & v882bdd;
assign v8fd928 = EMPTY_p & v884920 | !EMPTY_p & !v8805d7;
assign v880f84 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86ef5c;
assign v884b6c = StoB_REQ3_p & v8822d4 | !StoB_REQ3_p & !v844f91;
assign v8fd204 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8b6088;
assign v8ac1fa = DEQ_p & v887a7c | !DEQ_p & v8587ba;
assign v884170 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8fd186;
assign v8c2de5 = jx1_p & v885144 | !jx1_p & v8827ef;
assign v8fd7af = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd841;
assign v880f35 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8830bf;
assign v87fed4 = jx2_p & v8fd5b6 | !jx2_p & !v844f91;
assign v88417e = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v8861bc;
assign v87734f = stateG12_p & v844fab | !stateG12_p & !v8fd4f0;
assign v8fd842 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v885149;
assign v882b41 = jx1_p & v8843d0 | !jx1_p & v8fcd8f;
assign v8fcba5 = jx1_p & v8fd5d1 | !jx1_p & v86ec4a;
assign v8fd871 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8847a4;
assign v8fd8d4 = jx1_p & v8676b7 | !jx1_p & v8fd457;
assign v885c76 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fc68e;
assign v87adc8 = jx1_p & v8dacfe | !jx1_p & v885d67;
assign v891109 = stateG12_p & v8fcdd0 | !stateG12_p & v885d96;
assign v8d4bf0 = StoB_REQ6_p & v8fc78f | !StoB_REQ6_p & v885695;
assign v8fd1a6 = jx0_p & v898e61 | !jx0_p & v844f91;
assign v8fce44 = BtoS_ACK0_p & v882ae8 | !BtoS_ACK0_p & v8856d5;
assign v880f76 = BtoS_ACK0_p & v8fd7c8 | !BtoS_ACK0_p & v8846d2;
assign v858796 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8878ac;
assign v88366d = BtoS_ACK6_p & v8fd629 | !BtoS_ACK6_p & v8fd571;
assign v88429a = jx1_p & v8dabe8 | !jx1_p & !v854be6;
assign v8fd7e8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8841eb;
assign v8fd91a = BtoR_REQ1_p & v8fc9ca | !BtoR_REQ1_p & v8f2a57;
assign v8fd66a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc692;
assign v8fd7f7 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v880660;
assign v8b60ca = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v880f9a;
assign v8fd6bc = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v880231;
assign v8fd7a5 = BtoR_REQ0_p & v882f72 | !BtoR_REQ0_p & v8fd857;
assign v8fd62f = jx2_p & v8947ed | !jx2_p & v88791d;
assign v883158 = jx1_p & v883050 | !jx1_p & v8fd8f6;
assign v86bd4d = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8fd726;
assign v8fd2b1 = jx0_p & v880ac1 | !jx0_p & v887b09;
assign v8856c1 = StoB_REQ3_p & v8fd726 | !StoB_REQ3_p & v89736f;
assign v887ac6 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8fca41;
assign v884497 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v88225a;
assign v8fd727 = stateG7_1_p & v880fe9 | !stateG7_1_p & v844f91;
assign v884f6d = jx1_p & v881720 | !jx1_p & v885d0f;
assign v884f8c = jx0_p & v887ab9 | !jx0_p & v8fd652;
assign v8fd611 = EMPTY_p & v88e3ec | !EMPTY_p & v8859af;
assign v8fd852 = jx2_p & v8770c9 | !jx2_p & v8fd90d;
assign v8591df = jx1_p & v8fc1c0 | !jx1_p & v844f91;
assign v85397b = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v885215;
assign v8fc9fd = BtoR_REQ1_p & v884d3b | !BtoR_REQ1_p & v882d42;
assign v882772 = StoB_REQ1_p & v8ce111 | !StoB_REQ1_p & v8809d1;
assign v8830ac = BtoR_REQ1_p & v8fd879 | !BtoR_REQ1_p & v884b2b;
assign v88e7c3 = jx1_p & v88265b | !jx1_p & v8809b9;
assign v8540de = jx1_p & v85cf4b | !jx1_p & v8fc7cc;
assign v8fc78f = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v881840;
assign v8876cd = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8fc1f8;
assign v885d96 = BtoR_REQ0_p & v8fd54e | !BtoR_REQ0_p & v8fd79c;
assign v8fc810 = RtoB_ACK1_p & v88386a | !RtoB_ACK1_p & v844f91;
assign v8f29f1 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd690;
assign v8dac2c = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd174;
assign v8fd813 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v881f1a;
assign v858acb = stateG7_1_p & v858564 | !stateG7_1_p & v884329;
assign v8860bd = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fcf25;
assign v8972d7 = RtoB_ACK0_p & v88046c | !RtoB_ACK0_p & v880b5b;
assign v8fd60b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8845a2;
assign v88f0b3 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v8dab99;
assign v8a704c = BtoS_ACK1_p & v8fd5d4 | !BtoS_ACK1_p & v887868;
assign v890fdd = jx0_p & v8fd6a9 | !jx0_p & !v884359;
assign v884c5a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd6a7;
assign v8fd82b = jx0_p & v8fc2b8 | !jx0_p & !v8857fb;
assign v8fd698 = jx1_p & v844f91 | !jx1_p & v89facc;
assign v883b18 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v882699;
assign v8794e0 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v88489f;
assign v8fd90f = EMPTY_p & v8fcdd0 | !EMPTY_p & v8fd66c;
assign v8896fd = jx2_p & v8fd5e3 | !jx2_p & v87bb66;
assign v8fc2e5 = jx1_p & v8817bd | !jx1_p & v890d28;
assign v8878e0 = FULL_p & v8fd7a5 | !FULL_p & v8fd7b1;
assign v88068f = RtoB_ACK1_p & v882a0a | !RtoB_ACK1_p & v8878c8;
assign v8fcf73 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fd6e6;
assign v883d20 = BtoS_ACK6_p & v88315b | !BtoS_ACK6_p & v8806a6;
assign v88786b = StoB_REQ3_p & v8fd6d1 | !StoB_REQ3_p & !v844f91;
assign v8fc708 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8fd662;
assign v885102 = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v8fd2f7;
assign v885ea9 = RtoB_ACK1_p & v8fc945 | !RtoB_ACK1_p & v8fd62f;
assign v882136 = jx0_p & v88497c | !jx0_p & !v844f91;
assign v8795c1 = DEQ_p & v8fd599 | !DEQ_p & v88588a;
assign v88306a = StoB_REQ0_p & v8881e7 | !StoB_REQ0_p & v87945a;
assign v8879eb = BtoS_ACK1_p & v8fd932 | !BtoS_ACK1_p & v88234e;
assign v8807d3 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v870c76;
assign v8fd183 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v881edd;
assign v88201b = StoB_REQ1_p & v8fd24d | !StoB_REQ1_p & v8fd1b8;
assign v88369c = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & !v895c47;
assign v892c36 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd00a;
assign v8fd947 = BtoS_ACK3_p & v88576e | !BtoS_ACK3_p & v844f91;
assign v8fc651 = BtoS_ACK3_p & v88576e | !BtoS_ACK3_p & v8841f8;
assign v8fd83b = jx1_p & v8856e4 | !jx1_p & !v8642ea;
assign v887bef = jx2_p & v8fd284 | !jx2_p & v880816;
assign v884292 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8fd1f8;
assign v8850da = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88770f;
assign v8fd8c7 = BtoS_ACK0_p & v885be7 | !BtoS_ACK0_p & v88193e;
assign v89386c = BtoS_ACK6_p & v882bdd | !BtoS_ACK6_p & v8fd87f;
assign v8fccd5 = stateG12_p & v8fd452 | !stateG12_p & !v882d74;
assign v887a7f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd150;
assign v8fd6c2 = StoB_REQ0_p & v85397b | !StoB_REQ0_p & v844f91;
assign v8fd587 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8fd70d;
assign v8fc19e = BtoS_ACK2_p & v8fd646 | !BtoS_ACK2_p & v8879f2;
assign v88258c = stateG7_1_p & v8fd7ee | !stateG7_1_p & v8947b9;
assign v8cd9c1 = jx2_p & v891ac4 | !jx2_p & !v8fd084;
assign v8fd4f0 = BtoR_REQ0_p & v8810f4 | !BtoR_REQ0_p & v884a73;
assign v880931 = StoB_REQ6_p & v8fc68e | !StoB_REQ6_p & v894636;
assign v895a71 = StoB_REQ3_p & v881985 | !StoB_REQ3_p & !v882673;
assign v8fd17d = jx0_p & v880614 | !jx0_p & !v88174e;
assign v8fd7cf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88086e;
assign v883ddb = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v88093b;
assign v8fd8f8 = StoB_REQ2_p & v887c2f | !StoB_REQ2_p & v88576e;
assign v884b89 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v882b6f;
assign v880dc0 = BtoR_REQ0_p & v8fd882 | !BtoR_REQ0_p & v883776;
assign v8840c7 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v844f91;
assign v8fc1c0 = jx0_p & v8fd58c | !jx0_p & v844f91;
assign v8fd906 = BtoS_ACK0_p & v883759 | !BtoS_ACK0_p & v8fd1bc;
assign v8fd536 = jx2_p & v882d0f | !jx2_p & !v882f45;
assign v882bee = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v87bacb;
assign v887aed = jx2_p & v8c0098 | !jx2_p & !v8fd7f4;
assign v880d40 = jx0_p & v880816 | !jx0_p & v8fd5cc;
assign v880752 = jx0_p & v88407b | !jx0_p & v854139;
assign v883f1b = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8806c7;
assign v8fd94e = jx2_p & v8823d8 | !jx2_p & v8fcdd0;
assign v89fb46 = StoB_REQ0_p & v888096 | !StoB_REQ0_p & v8fcba4;
assign v881720 = jx0_p & v8810d4 | !jx0_p & v897303;
assign v8a87b9 = jx1_p & v8856e4 | !jx1_p & !v87b4e7;
assign v8fd256 = jx1_p & v844f91 | !jx1_p & !v88397a;
assign v8818a8 = jx0_p & v8fd760 | !jx0_p & v8fd8b4;
assign v885d31 = jx1_p & v8856e4 | !jx1_p & !v8974c9;
assign v88808a = jx0_p & v89fb1e | !jx0_p & v8fd7e6;
assign v8fd33e = stateG7_1_p & v87a65f | !stateG7_1_p & v8fd94e;
assign v8fd77d = StoB_REQ1_p & v8820ed | !StoB_REQ1_p & v88ec21;
assign v8fd36d = jx1_p & v8fd6a6 | !jx1_p & !v844f91;
assign v888182 = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & v844fb5;
assign v8fd623 = RtoB_ACK1_p & v883833 | !RtoB_ACK1_p & v8fc606;
assign v8861bc = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd819;
assign v880cff = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v88058c;
assign v884464 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v884da1;
assign v8fcae9 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8fd967;
assign v8b605d = BtoS_ACK6_p & v88402c | !BtoS_ACK6_p & v88299b;
assign v89110a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v887913;
assign v8fc9c2 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v858796;
assign v884ac0 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v88219e;
assign v8fd5fc = RtoB_ACK0_p & v8972bc | !RtoB_ACK0_p & v8fc6fe;
assign v895d18 = jx1_p & v887f32 | !jx1_p & v8843d0;
assign v8fd82e = jx2_p & v88259e | !jx2_p & !v88793c;
assign v8811ad = jx0_p & v8fc48c | !jx0_p & v8fcff6;
assign v8820a0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v880f84;
assign v895ceb = jx2_p & v883a4d | !jx2_p & !v844f91;
assign v8fca9d = StoB_REQ2_p & v8fd8df | !StoB_REQ2_p & v8588ba;
assign v895d6d = BtoR_REQ1_p & v88808c | !BtoR_REQ1_p & v8808f4;
assign v8fd793 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v88212e;
assign v8843d0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8877a0;
assign v887924 = RtoB_ACK1_p & v8fd879 | !RtoB_ACK1_p & v8fd5cd;
assign v884d11 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd6c2;
assign v8fd93c = StoB_REQ6_p & v884796 | !StoB_REQ6_p & v885e59;
assign v8fd5df = jx1_p & v8676b7 | !jx1_p & !v844f91;
assign v8827ef = jx0_p & v885144 | !jx0_p & v844f91;
assign v8fd696 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v887b46;
assign v8896fc = RtoB_ACK0_p & v8857e9 | !RtoB_ACK0_p & v882fd1;
assign v88394f = jx2_p & v882c16 | !jx2_p & !v844fab;
assign v8fd3ee = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v885185;
assign v884143 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v884d53;
assign v8fd6e3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd866;
assign v887b46 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8fd5f2;
assign v8fd6b3 = BtoS_ACK1_p & v88219e | !BtoS_ACK1_p & v887f3a;
assign v8fd1e2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88264d;
assign v880383 = BtoS_ACK1_p & v8fd932 | !BtoS_ACK1_p & v8fc986;
assign v8fce04 = FULL_p & v884867 | !FULL_p & v8fd57a;
assign v8819fb = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v884476;
assign v890ce8 = StoB_REQ1_p & v8843d1 | !StoB_REQ1_p & v858678;
assign v8fd58f = stateG7_1_p & v8b6054 | !stateG7_1_p & v8816aa;
assign v8b6045 = jx2_p & v8fd5df | !jx2_p & v8fd6d7;
assign v8cd9ef = DEQ_p & v880a3a | !DEQ_p & v8fd651;
assign v880bb6 = StoB_REQ0_p & v8fc2d4 | !StoB_REQ0_p & v887d67;
assign v87d828 = BtoR_REQ0_p & v88295b | !BtoR_REQ0_p & v888046;
assign v895ce5 = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v8fc76f;
assign v887c6c = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v8816ab;
assign v887de8 = StoB_REQ3_p & v8fd7f7 | !StoB_REQ3_p & !v880660;
assign v887906 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v8fce18;
assign v8fd28e = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8f29f1;
assign v883837 = jx1_p & v8fd18f | !jx1_p & !v885b44;
assign v8fcf97 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v87dfe7;
assign v8fd23e = StoB_REQ6_p & v8831ee | !StoB_REQ6_p & v8881fb;
assign v8fd6e0 = stateG12_p & v88251a | !stateG12_p & !v884984;
assign v882859 = jx2_p & v869e2c | !jx2_p & !v883a2e;
assign v8fd5a2 = jx2_p & v8fd1c7 | !jx2_p & v884a6e;
assign v8861c0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd1c5;
assign v8fd7b3 = jx2_p & v882459 | !jx2_p & !v8fd1af;
assign v883b2a = jx2_p & v8fd7f3 | !jx2_p & !v8f2a7d;
assign v895a56 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ad097;
assign v8fd936 = BtoS_ACK0_p & v89471b | !BtoS_ACK0_p & v883c46;
assign v8818b7 = BtoR_REQ0_p & v8826ea | !BtoR_REQ0_p & v896f10;
assign v880a3a = ENQ_p & v87734f | !ENQ_p & !v8fd770;
assign v885fb3 = BtoS_ACK1_p & v8fd17e | !BtoS_ACK1_p & v8861f9;
assign v88305d = BtoR_REQ1_p & v8fd648 | !BtoR_REQ1_p & v8fd837;
assign v8fd64c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd1a0;
assign v888057 = BtoR_REQ0_p & v8fc762 | !BtoR_REQ0_p & v8fd90c;
assign v881686 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd7b7;
assign v8859f7 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v884fdd;
assign v8fd209 = stateG7_1_p & v883046 | !stateG7_1_p & v88774e;
assign v88ed82 = jx0_p & v8809c4 | !jx0_p & v8fd5fa;
assign v8847a4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd744;
assign v87954a = jx1_p & v85e9fa | !jx1_p & !v884ba1;
assign v884919 = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v882baa;
assign v8fd7aa = stateG7_1_p & v8ad053 | !stateG7_1_p & v844f91;
assign v887a24 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8821b5;
assign v8fd251 = BtoR_REQ1_p & v8fc5f2 | !BtoR_REQ1_p & v8fce5c;
assign v885fe8 = BtoS_ACK0_p & v887c3e | !BtoS_ACK0_p & !v8fd3ee;
assign v8ed1d1 = RtoB_ACK1_p & v891b69 | !RtoB_ACK1_p & v85f322;
assign v8fc1f9 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & v88576e;
assign v882b6f = StoB_REQ3_p & v844fb1 | !StoB_REQ3_p & v844f91;
assign v8840b0 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd8cc;
assign v8fd5d6 = RtoB_ACK1_p & v864119 | !RtoB_ACK1_p & v8fd5fd;
assign v885b36 = jx0_p & v8fc18e | !jx0_p & v8fcb01;
assign v8ce0f7 = BtoS_ACK0_p & v882e12 | !BtoS_ACK0_p & v8fc6b2;
assign v883de0 = RtoB_ACK1_p & v880821 | !RtoB_ACK1_p & v8fc6fe;
assign v8fcd30 = BtoS_ACK0_p & v88493b | !BtoS_ACK0_p & v8fd5ee;
assign v87d10c = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd8cf;
assign v880d6b = StoB_REQ1_p & v8ac9cb | !StoB_REQ1_p & v8818f6;
assign v884953 = BtoR_REQ1_p & v882302 | !BtoR_REQ1_p & v844f91;
assign v8fce7b = RtoB_ACK0_p & v8878c8 | !RtoB_ACK0_p & v859713;
assign v8fcf10 = jx1_p & v8676b7 | !jx1_p & v8843ae;
assign v8820d8 = StoB_REQ6_p & v8fd8e4 | !StoB_REQ6_p & v887f88;
assign v858a41 = stateG12_p & v884842 | !stateG12_p & v8c48b2;
assign v879486 = RtoB_ACK0_p & v8fd777 | !RtoB_ACK0_p & v8fd65a;
assign v884bdc = StoB_REQ1_p & v883bef | !StoB_REQ1_p & v880507;
assign v887f47 = RtoB_ACK0_p & v8fd879 | !RtoB_ACK0_p & v8830ac;
assign v883968 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v880d6b;
assign v884256 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8fcc2e;
assign v88b623 = BtoS_ACK6_p & v89471b | !BtoS_ACK6_p & v8fd1f3;
assign v8a88d5 = FULL_p & v88bc54 | !FULL_p & v8fd685;
assign v8fceeb = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fc99d;
assign v8880b3 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v88807f;
assign v882fd7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd002;
assign v8a87de = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8ac9e4;
assign v8809eb = jx1_p & v88454a | !jx1_p & v868a24;
assign v8ed18b = BtoS_ACK6_p & v8fd1bd | !BtoS_ACK6_p & v858a9b;
assign v8fd8b1 = StoB_REQ1_p & v87653c | !StoB_REQ1_p & v8846a5;
assign v880ac1 = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v8fd75c;
assign v88397d = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8880b3;
assign v8c2e51 = stateG7_1_p & v885ea9 | !stateG7_1_p & v8fd62f;
assign v894703 = jx2_p & v8fd5f7 | !jx2_p & !v8f2a7d;
assign v8880e0 = RtoB_ACK1_p & v8fd95c | !RtoB_ACK1_p & v8fd581;
assign v8fd94f = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v8ac9d6;
assign v8a7085 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fd63e;
assign v8fd568 = RtoB_ACK1_p & v887b15 | !RtoB_ACK1_p & v87fed4;
assign v8fd379 = StoB_REQ0_p & v8fd1e1 | !StoB_REQ0_p & v8816f3;
assign v883752 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v895c65;
assign v885d73 = RtoB_ACK1_p & v8fd20f | !RtoB_ACK1_p & v88589c;
assign v8fd1f8 = stateG7_1_p & v8fd8c9 | !stateG7_1_p & v895abe;
assign v8fd882 = RtoB_ACK0_p & v87fed4 | !RtoB_ACK0_p & v894b33;
assign v8588ba = StoB_REQ3_p & v8fc1cf | !StoB_REQ3_p & v844f91;
assign v8fcd47 = stateG7_1_p & v8cd9c1 | !stateG7_1_p & v844f91;
assign v8563aa = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd8d8;
assign v870c76 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v88241f;
assign v88e3ec = BtoR_REQ0_p & v883aae | !BtoR_REQ0_p & v8ed1ce;
assign v887ad9 = RtoB_ACK1_p & v88394f | !RtoB_ACK1_p & v882db5;
assign v8fd8b7 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v88810f;
assign v880665 = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v89fb49;
assign v887d16 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88578e;
assign v8817c2 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8824dc;
assign v891ac4 = jx1_p & v88401d | !jx1_p & !v8fc7cc;
assign v882bb2 = StoB_REQ3_p & v88e1fb | !StoB_REQ3_p & v883071;
assign v8fd08a = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v8fd7f0;
assign v882563 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8fca9c;
assign v8fd7a1 = StoB_REQ3_p & v86ed40 | !StoB_REQ3_p & v8824dc;
assign v88f9d2 = StoB_REQ6_p & v844f97 | !StoB_REQ6_p & v8fd5ff;
assign v895c31 = StoB_REQ2_p & v8fd8f4 | !StoB_REQ2_p & v88786b;
assign v883c09 = jx1_p & v844f91 | !jx1_p & v8fce9e;
assign v885fb8 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v883e11;
assign v8fd738 = BtoS_ACK6_p & v8fd5ff | !BtoS_ACK6_p & v8fc61e;
assign v8fd736 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v844f91;
assign v880674 = BtoS_ACK1_p & v8fd7dc | !BtoS_ACK1_p & v8fd716;
assign v880c0e = StoB_REQ3_p & v8fd6ae | !StoB_REQ3_p & v8896ed;
assign v8fd741 = BtoS_ACK6_p & v88089e | !BtoS_ACK6_p & v884cd5;
assign v8fd6d3 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v87fee8;
assign v8cecad = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd738;
assign v883050 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v882093;
assign v8fd809 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v882bdd;
assign v883890 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v880294;
assign v885b87 = BtoS_ACK6_p & v8fd7dc | !BtoS_ACK6_p & v8fd939;
assign v8fd455 = StoB_REQ2_p & v880c0e | !StoB_REQ2_p & v8fd6ae;
assign v8dac53 = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v85b93e;
assign v8fd816 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8fd17e;
assign v88576c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc46b;
assign v88052d = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8fc1f9;
assign v885b3a = jx0_p & v8fd6a9 | !jx0_p & v844f91;
assign v8846fc = StoB_REQ6_p & v8fd865 | !StoB_REQ6_p & v883968;
assign v88096b = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v887bbe;
assign v8fd1bd = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8879ab;
assign v8fd1fe = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8daba0;
assign v895b31 = BtoS_ACK6_p & v882d6b | !BtoS_ACK6_p & v881686;
assign v8802a2 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd6a0;
assign v885ddd = jx2_p & v8a87b9 | !jx2_p & !v8587e6;
assign v8848b0 = RtoB_ACK1_p & v88055d | !RtoB_ACK1_p & v8fd659;
assign v8c2eaf = StoB_REQ6_p & v844f97 | !StoB_REQ6_p & v8fd764;
assign v880ed2 = jx2_p & v8fd700 | !jx2_p & v8fd6b2;
assign v881141 = RtoB_ACK1_p & v8fc9ca | !RtoB_ACK1_p & v8fce5c;
assign v8fd612 = jx1_p & v8856e4 | !jx1_p & !v8fd689;
assign v8c2de8 = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v8fd1bb;
assign v8fd8d8 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v883ddb;
assign v88186f = BtoS_ACK2_p & v89476c | !BtoS_ACK2_p & v85b247;
assign v8fc67f = BtoS_ACK6_p & v88402c | !BtoS_ACK6_p & v884875;
assign v885d08 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd8f4;
assign v8569e0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8803e6;
assign v8fc495 = jx2_p & v885eba | !jx2_p & v87954a;
assign v8fd24e = StoB_REQ6_p & v884de8 | !StoB_REQ6_p & v885e9b;
assign v8fd7f0 = StoB_REQ1_p & v8fd6c5 | !StoB_REQ1_p & v885d0d;
assign v8fd2a7 = StoB_REQ5_n & v844f9f | !StoB_REQ5_n & !v844f91;
assign v8841cd = jx1_p & v885a6c | !jx1_p & v87001c;
assign v8f2a2c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v887ac6;
assign v8881d4 = BtoR_REQ1_p & v8fc7b1 | !BtoR_REQ1_p & v87eaaf;
assign v88372b = jx1_p & v884d94 | !jx1_p & v881fe6;
assign v881649 = BtoS_ACK0_p & v844f9e | !BtoS_ACK0_p & v8fd484;
assign v8fd218 = jx2_p & v844f91 | !jx2_p & v8fd747;
assign v880fa6 = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v885bcf;
assign v8fd68f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd579;
assign v8fd1b9 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd80f;
assign v8fd6bf = jx1_p & v880d40 | !jx1_p & !v8fcc62;
assign v8c4d26 = DEQ_p & v88096f | !DEQ_p & !v884b78;
assign v8fc98c = jx0_p & v8fd5ac | !jx0_p & !v882e37;
assign v8fd284 = jx1_p & v880816 | !jx1_p & !v8ed1c6;
assign v884a71 = FULL_p & v8d477f | !FULL_p & v8fd71a;
assign v8fcb34 = stateG7_1_p & v887904 | !stateG7_1_p & v844f91;
assign v895c60 = RtoB_ACK1_p & v8fc7b1 | !RtoB_ACK1_p & v844f91;
assign v8fd95f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cd9b9;
assign v88058c = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844fb1;
assign v895c65 = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & !v8fd1da;
assign v885de9 = BtoS_ACK6_p & v8fd7dc | !BtoS_ACK6_p & v887c44;
assign v8fce28 = RtoB_ACK0_p & v8fd5b0 | !RtoB_ACK0_p & v894722;
assign v89fb02 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v884f00;
assign v8878bb = stateG7_1_p & v888062 | !stateG7_1_p & v844f91;
assign v8fcaa8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a8786;
assign v8fd60e = RtoB_ACK0_p & v882d42 | !RtoB_ACK0_p & v884d5e;
assign v8fd478 = StoB_REQ1_p & v85879a | !StoB_REQ1_p & v844f91;
assign v8fd796 = BtoS_ACK6_p & v882bdd | !BtoS_ACK6_p & v884a33;
assign v885eba = jx1_p & v880ccb | !jx1_p & !v8818e1;
assign v8fd701 = RtoB_ACK1_p & v8fce5c | !RtoB_ACK1_p & v8f2a57;
assign v8860d7 = BtoS_ACK1_p & v8fd002 | !BtoS_ACK1_p & v887627;
assign v884476 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v882d8f;
assign v8fd585 = jx2_p & v8fd921 | !jx2_p & v8fd084;
assign v854a91 = RtoB_ACK0_p & v8fd5a2 | !RtoB_ACK0_p & v8fd876;
assign v887879 = jx0_p & v8841bc | !jx0_p & v8fd238;
assign v88599b = RtoB_ACK0_p & v8fd688 | !RtoB_ACK0_p & v887efe;
assign v8fd8f4 = StoB_REQ3_p & v887768 | !StoB_REQ3_p & !v844f91;
assign v8fd627 = StoB_REQ1_p & v8f2a5a | !StoB_REQ1_p & v88ec29;
assign v88383e = stateG7_1_p & v8fc5e1 | !stateG7_1_p & v8fd218;
assign v8fc46b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v8b89cf;
assign v883e92 = jx2_p & v89faf7 | !jx2_p & v8843d0;
assign v8fd484 = BtoS_ACK6_p & v844f9e | !BtoS_ACK6_p & v8fd790;
assign v896f10 = RtoB_ACK0_p & v8989c5 | !RtoB_ACK0_p & v8fd6d9;
assign v8947ee = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8e1d28;
assign v874ed6 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v885b62;
assign v895aff = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v882f82;
assign v8562b0 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v883852;
assign v885a16 = RtoB_ACK1_p & v88ea40 | !RtoB_ACK1_p & v8fc495;
assign v8fd764 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v882bdd;
assign v8fcd1f = BtoS_ACK2_p & v882d8f | !BtoS_ACK2_p & v885df9;
assign v8fd7cb = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v88576e;
assign v885c69 = stateG7_1_p & v8fd623 | !stateG7_1_p & v8fd6de;
assign v880403 = BtoR_REQ0_p & v883cf7 | !BtoR_REQ0_p & v8830bd;
assign v8ad053 = RtoB_ACK1_p & v87eaaf | !RtoB_ACK1_p & v844f91;
assign v87943e = BtoR_REQ0_p & v8876cd | !BtoR_REQ0_p & v89fac8;
assign v8fd1ca = jx1_p & v8fd88d | !jx1_p & v887c9a;
assign v8ce165 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v894828 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8ad097;
assign v88498b = RtoB_ACK0_p & v8fc945 | !RtoB_ACK0_p & v8fd846;
assign v885185 = BtoS_ACK6_p & v8fd5ff | !BtoS_ACK6_p & !v887d78;
assign v885be7 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v844f91;
assign v8fd57a = BtoR_REQ0_p & v8fd25a | !BtoR_REQ0_p & v8fd1d9;
assign v868a24 = jx0_p & v8fcbe3 | !jx0_p & v8ce165;
assign v88380c = jx0_p & v844f91 | !jx0_p & v8846ba;
assign v85bfad = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v887c92;
assign v8fd82a = jx0_p & v8fd58c | !jx0_p & !v88232b;
assign v86f4d0 = BtoR_REQ1_p & v887b15 | !BtoR_REQ1_p & v87fed4;
assign v8fcbb4 = StoB_REQ0_p & v8a87de | !StoB_REQ0_p & v88ea5a;
assign v8ac9b2 = BtoR_REQ0_p & v8fcecd | !BtoR_REQ0_p & v8fc801;
assign v885c13 = BtoR_REQ1_p & v8fd197 | !BtoR_REQ1_p & !v844f91;
assign v884a6d = jx0_p & v844f91 | !jx0_p & v87bb66;
assign v892156 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v887fa9;
assign v8fd8ed = RtoB_ACK1_p & v85f322 | !RtoB_ACK1_p & v844f91;
assign v8fd1ba = jx0_p & v88785b | !jx0_p & v8827ac;
assign v8896ed = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v8fd6ae;
assign v88e73e = StoB_REQ6_p & v8fd903 | !StoB_REQ6_p & v885a06;
assign v884b78 = ENQ_p & v884049 | !ENQ_p & v887680;
assign v8fd745 = BtoS_ACK1_p & v8fd932 | !BtoS_ACK1_p & v8ce184;
assign v882a64 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v883d05;
assign v8851ef = RtoB_ACK1_p & v8fd659 | !RtoB_ACK1_p & v8fd218;
assign v8fd356 = jx1_p & v8fd6a6 | !jx1_p & v8fd77b;
assign v8805dc = BtoS_ACK6_p & v882baa | !BtoS_ACK6_p & v88085d;
assign v8fd6d7 = jx1_p & v8817bd | !jx1_p & v844f91;
assign v887656 = EMPTY_p & v8fd823 | !EMPTY_p & v8fcabb;
assign v885b21 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v882f33;
assign v8821ba = jx0_p & v880ac1 | !jx0_p & v8fc1a7;
assign v88ebbe = stateG7_1_p & v88565d | !stateG7_1_p & v844f91;
assign v854bb9 = StoB_REQ2_p & v8fd5f2 | !StoB_REQ2_p & v882d8f;
assign v8fd8cc = BtoS_ACK2_p & v8fd646 | !BtoS_ACK2_p & v8fd576;
assign v8594cb = jx1_p & v8827ac | !jx1_p & v8fd77a;
assign v885b44 = jx0_p & v8fd011 | !jx0_p & !v885102;
assign v883c46 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd7ed;
assign v887b5a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8827b2;
assign v8fd70d = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v844f91;
assign v8fd24d = BtoS_ACK2_p & v882d8f | !BtoS_ACK2_p & v8dacf2;
assign v8c2e6c = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v8ac1f3;
assign v881f1a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd5dc;
assign v8fd940 = jx0_p & v844f9b | !jx0_p & !v844f91;
assign v8fd6de = jx2_p & v8fd56f | !jx2_p & v881117;
assign v8948c3 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v88576e;
assign v8ad047 = jx2_p & v8fd75d | !jx2_p & v8fc691;
assign v8fd896 = jx2_p & v8841cd | !jx2_p & v88793c;
assign v8fd899 = jx1_p & v8c2eb8 | !jx1_p & v844f91;
assign v8fd5b0 = jx2_p & v885d31 | !jx2_p & !v88793c;
assign v8fd775 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v881f1a;
assign v8fd80d = BtoS_ACK1_p & v8fd002 | !BtoS_ACK1_p & v8fd1dd;
assign v8fd913 = BtoS_ACK2_p & v8fd953 | !BtoS_ACK2_p & v895c31;
assign v8dabf0 = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v85872e;
assign v8fd59c = jx1_p & v8676b7 | !jx1_p & v8fd1a6;
assign v8fd95a = BtoR_REQ0_p & v879486 | !BtoR_REQ0_p & v8fd285;
assign v8fd1dd = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v882048;
assign v8fc844 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v885f1e;
assign v885f76 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88784a;
assign v880f66 = StoB_REQ6_p & v89fb02 | !StoB_REQ6_p & v8838a3;
assign v885909 = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v882905;
assign v876549 = StoB_REQ6_p & v892c36 | !StoB_REQ6_p & v8fcc77;
assign v8fd63c = StoB_REQ6_p & v883879 | !StoB_REQ6_p & v844f91;
assign v8dac8a = jx0_p & v885fe3 | !jx0_p & v8fd7e6;
assign v8fd3b5 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8842b7;
assign v8fd74b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd745;
assign v880ccb = jx0_p & v88507a | !jx0_p & v86a020;
assign v8fd866 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844faf;
assign v886012 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v880af8;
assign v858985 = RtoB_ACK1_p & v880ed2 | !RtoB_ACK1_p & v882a0a;
assign v880804 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v883781;
assign v8fd96b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86b3d4;
assign v88264d = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v883879;
assign v8830a5 = jx1_p & v88401d | !jx1_p & v844f91;
assign v8829b5 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v88310a;
assign v884d3b = jx2_p & v8fd69d | !jx2_p & !v88793c;
assign v86ecdb = BtoR_REQ0_p & v8fcdd0 | !BtoR_REQ0_p & v866b82;
assign v87dfc7 = RtoB_ACK1_p & v887bef | !RtoB_ACK1_p & v8fc7b1;
assign v8fd72e = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v885e24;
assign v8846bf = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v88386a;
assign v885063 = BtoS_ACK0_p & v89471b | !BtoS_ACK0_p & v8fcaa8;
assign v88391f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v88219e;
assign v8fd315 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v882d6b;
assign v880d66 = StoB_REQ1_p & v885df9 | !StoB_REQ1_p & v844f91;
assign v8946a5 = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v8b606c;
assign v8fc182 = jx0_p & v8fc2b2 | !jx0_p & v8f2a3f;
assign v88567a = StoB_REQ0_p & v887fa9 | !StoB_REQ0_p & v844f91;
assign v8881bb = jx1_p & v8fd922 | !jx1_p & !v885fda;
assign v880620 = StoB_REQ1_p & v885d08 | !StoB_REQ1_p & v8fd913;
assign v882a93 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ad0e2;
assign v8810f4 = RtoB_ACK0_p & v88394f | !RtoB_ACK0_p & v882db5;
assign v8819df = RtoB_ACK1_p & v8fd659 | !RtoB_ACK1_p & v844f91;
assign v8587ba = ENQ_p & v889757 | !ENQ_p & v8fd467;
assign v8773cf = stateG7_1_p & v88f395 | !stateG7_1_p & v8fd234;
assign v8fc5f2 = stateG7_1_p & v8fd880 | !stateG7_1_p & v8fc9ca;
assign v88079c = StoB_REQ4_p & v888182 | !StoB_REQ4_p & v844f91;
assign v885da7 = jx1_p & v88401d | !jx1_p & !v884b56;
assign v882908 = BtoS_ACK0_p & v882e12 | !BtoS_ACK0_p & v880834;
assign v87bbad = jx2_p & v8fd68b | !jx2_p & !v8fd356;
assign v882db5 = jx2_p & v8fd918 | !jx2_p & !v844fab;
assign v88fa48 = BtoS_ACK2_p & v8fd646 | !BtoS_ACK2_p & v8fd932;
assign v895b24 = BtoS_ACK1_p & v885be7 | !BtoS_ACK1_p & v895abb;
assign v85872e = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v895b52;
assign v88289d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v887b14;
assign v885ab1 = BtoR_REQ1_p & v8c2e51 | !BtoR_REQ1_p & v895b2f;
assign v8947da = jx1_p & v88271c | !jx1_p & v8fcdd0;
assign v887c92 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8837fe;
assign v885f69 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8f2a5a;
assign v8fd4f5 = StoB_REQ2_p & v8f2a19 | !StoB_REQ2_p & v844f91;
assign v86ecd4 = BtoR_REQ1_p & v885b2d | !BtoR_REQ1_p & v844f91;
assign v8fd25d = StoB_REQ2_p & v882bb2 | !StoB_REQ2_p & v8fd24a;
assign v887cfa = BtoR_REQ0_p & v8fd8fb | !BtoR_REQ0_p & v88305d;
assign v8587e6 = jx1_p & v884fa4 | !jx1_p & v8808cf;
assign v8826ea = RtoB_ACK0_p & v8fd6d9 | !RtoB_ACK0_p & v883e1c;
assign v8fca4a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883105;
assign v8fd67e = StoB_REQ6_p & v8fd786 | !StoB_REQ6_p & v8fd589;
assign v88fa9a = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v880bb6;
assign BtoS_ACK4_n = !v8c2ef2;
assign v88783d = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fc970;
assign v883c06 = StoB_REQ4_p & v888182 | !StoB_REQ4_p & !v844f91;
assign v8823c2 = BtoR_REQ1_p & v887d8f | !BtoR_REQ1_p & v8fd788;
assign v8838c5 = StoB_REQ0_p & v8fd8d8 | !StoB_REQ0_p & v844f9d;
assign v8fd5bf = jx1_p & v8fc5a6 | !jx1_p & v887d5b;
assign v8fd8e4 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8dac2c;
assign v884904 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844fb3;
assign BtoR_REQ1_n = !v8ac1fa;
assign v88774e = jx2_p & v89fb10 | !jx2_p & !v8829eb;
assign v8fd7b7 = BtoS_ACK1_p & v882d6b | !BtoS_ACK1_p & v8fd315;
assign v8fd7b2 = jx1_p & v8824d4 | !jx1_p & !v8894e3;
assign v879581 = jx2_p & v884d47 | !jx2_p & v8fcb01;
assign v8fd819 = BtoS_ACK1_p & v88219e | !BtoS_ACK1_p & v88289d;
assign v885a06 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v884bdc;
assign BtoS_ACK2_n = !v8f2abf;
assign v8684ff = jx1_p & v884f8c | !jx1_p & v8809b9;
assign v86deca = stateG7_1_p & v88e2ce | !stateG7_1_p & v894722;
assign v891594 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v884ccb;
assign v8c2eb0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ad0d9;
assign v881e44 = BtoR_REQ1_p & v889be1 | !BtoR_REQ1_p & v8fc8ca;
assign v885b89 = StoB_REQ4_p & v888182 | !StoB_REQ4_p & v844f9f;
assign v8972ae = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v895d4b;
assign v8821dc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c2de8;
assign v8817bd = jx0_p & v8fd760 | !jx0_p & v844f91;
assign v881923 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v88621e;
assign v882e65 = BtoR_REQ1_p & v883e2e | !BtoR_REQ1_p & v8fd5a2;
assign v8ed1b3 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & !v8848a0;
assign v887baf = BtoR_REQ1_p & v8fd659 | !BtoR_REQ1_p & v8fd218;
assign v895cb0 = BtoR_REQ0_p & v8802a4 | !BtoR_REQ0_p & v8c2e6b;
assign v85b247 = StoB_REQ2_p & v887ac6 | !StoB_REQ2_p & v8fca41;
assign v8c48b6 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v885867;
assign v8861ed = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v853f24;
assign v888056 = BtoS_ACK6_p & v885d25 | !BtoS_ACK6_p & v884796;
assign v8fd3c6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v882bdd;
assign v8a8786 = BtoS_ACK6_p & v89471b | !BtoS_ACK6_p & v8fc68e;
assign v8fd690 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & !v844f91;
assign v8fd75c = StoB_REQ0_p & v8ad0d9 | !StoB_REQ0_p & v8839d5;
assign v882de0 = RtoB_ACK0_p & v884329 | !RtoB_ACK0_p & v8583a8;
assign v88bb4f = BtoR_REQ0_p & v854a91 | !BtoR_REQ0_p & v8fd51f;
assign v884842 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v8fd869;
assign v8fd58b = stateG12_p & v888057 | !stateG12_p & v88107d;
assign v887fe2 = BtoS_ACK6_p & v88402c | !BtoS_ACK6_p & v8fd929;
assign v885df9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v882d8f;
assign v8fd244 = BtoS_ACK6_p & v885b17 | !BtoS_ACK6_p & !v8fd570;
assign v884013 = jx0_p & v88390f | !jx0_p & !v8843ba;
assign v8fcd8f = jx0_p & v8fd608 | !jx0_p & v8843d0;
assign v8fd195 = stateG12_p & v885ea3 | !stateG12_p & v87bb66;
assign v8947e2 = StoB_REQ6_p & v883b45 | !StoB_REQ6_p & v882719;
assign v8972bc = BtoR_REQ1_p & v880821 | !BtoR_REQ1_p & v8fc6fe;
assign v89726a = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v8fd73a;
assign v885119 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8f2a0b;
assign v8ed1d8 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8a7085;
assign v8fd932 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8fd646;
assign v8c4d01 = jx1_p & v880ccb | !jx1_p & !v8fd2b1;
assign v8fc5ad = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f97;
assign v8fd805 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8847e5;
assign v883a7f = StoB_REQ1_p & v8fd5dc | !StoB_REQ1_p & v844f91;
assign v8fd1ea = jx0_p & v892417 | !jx0_p & !v8fd879;
assign v8fd25a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8fd950;
assign v8c2ebb = stateG12_p & v8805b9 | !stateG12_p & !v8fd80a;
assign v8fd734 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd7a0;
assign v882d73 = jx0_p & v884bc5 | !jx0_p & v882bc8;
assign v895bb6 = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v89fb1c;
assign v880a2a = BtoR_REQ0_p & v8ed983 | !BtoR_REQ0_p & v8861df;
assign v8878bd = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v8825fc;
assign v8816e8 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8fd636;
assign v859c5b = StoB_REQ3_p & v8fd7f7 | !StoB_REQ3_p & !v844fb3;
assign v882b76 = ENQ_p & v8ad0c2 | !ENQ_p & v895d15;
assign v88295b = RtoB_ACK0_p & v88055d | !RtoB_ACK0_p & v8fd659;
assign v8fd950 = stateG7_1_p & v883d66 | !stateG7_1_p & v87eaaf;
assign v8a705e = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fc21f;
assign v8fd7ff = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v87af07;
assign v8fd846 = stateG7_1_p & v8fc64f | !stateG7_1_p & v8fd62f;
assign v8fd63e = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8817c2;
assign v8fc2b2 = BtoS_ACK0_p & v8fd8dd | !BtoS_ACK0_p & v883bb8;
assign v8fd6a0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8843b6;
assign v8818fb = jx0_p & v8827ac | !jx0_p & v8fd683;
assign v895b92 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v8fd3cb;
assign v887fec = BtoS_ACK6_p & v882bdd | !BtoS_ACK6_p & v8fd6f1;
assign v8c4d03 = StoB_REQ1_p & v8fd597 | !StoB_REQ1_p & v8fd5dd;
assign v8ac9e4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8ad0e2;
assign v887a7a = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v887f4e;
assign v8a87b1 = StoB_REQ1_p & v884476 | !StoB_REQ1_p & v8fd70d;
assign v854139 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fcf21;
assign v88100b = jx1_p & v880240 | !jx1_p & v8843d0;
assign v844fa5 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844f91;
assign v884dec = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v8fca9d;
assign v887abb = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v884203;
assign v8f2a14 = BtoS_ACK0_p & v882e12 | !BtoS_ACK0_p & v881f4a;
assign v88eb82 = BtoS_ACK2_p & v8fd5ad | !BtoS_ACK2_p & v88219e;
assign v8f29e2 = jx2_p & v887cf6 | !jx2_p & v8846ba;
assign v88837d = BtoS_ACK0_p & v8fd809 | !BtoS_ACK0_p & !v8cd9b9;
assign v8fd5a6 = jx1_p & v8dabff | !jx1_p & v8fd8e2;
assign v8fd715 = BtoR_REQ1_p & v85397c | !BtoR_REQ1_p & v8878bb;
assign v880717 = StoB_REQ6_p & v853f24 | !StoB_REQ6_p & !v844f91;
assign v8fd5ea = jx1_p & v8fd6aa | !jx1_p & !v8fd538;
assign v885694 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v891114;
assign v8fd576 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8fd667;
assign v878328 = StoB_REQ4_p & v844f9f | !StoB_REQ4_p & !v844f91;
assign v882006 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844fa1;
assign v8fd646 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v88576e;
assign v88fdf5 = jx0_p & v884767 | !jx0_p & v883ad4;
assign v8dacfe = jx0_p & v8ce165 | !jx0_p & v882c83;
assign v890fd8 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8820ed;
assign v88588a = ENQ_p & v8829ee | !ENQ_p & v8fd611;
assign v88604b = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v8fd863;
assign v8ac9ad = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v8fd5f2;
assign v888205 = BtoS_ACK0_p & v8fd853 | !BtoS_ACK0_p & v8fca05;
assign v8ce0f4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8881bd;
assign v887768 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v844f91;
assign v881f75 = jx0_p & v8fc67a | !jx0_p & !v844f91;
assign v8fd66c = stateG12_p & v86ecdb | !stateG12_p & v8fcdd0;
assign v8fd5b3 = BtoR_REQ1_p & v8793ad | !BtoR_REQ1_p & v8fd17b;
assign v882459 = jx1_p & v8fd6ea | !jx1_p & v895b02;
assign v884da1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd1fe;
assign v886129 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & !v8861ed;
assign v8b607f = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8fd7a0;
assign v884577 = StoB_REQ0_p & v88e5f1 | !StoB_REQ0_p & v844f91;
assign v895afe = StoB_REQ0_p & v88783d | !StoB_REQ0_p & v88d4df;
assign v89471b = StoB_REQ1_p & v882bdd | !StoB_REQ1_p & v844f91;
assign v8fd868 = BtoS_ACK6_p & v8fd853 | !BtoS_ACK6_p & v8fd6c1;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v885f7b = jx0_p & v882908 | !jx0_p & v8ce0f7;
assign v8fc2dd = jx0_p & v8fd926 | !jx0_p & v883890;
assign v887b69 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8947e2;
assign v8fd810 = BtoS_ACK0_p & v880fd1 | !BtoS_ACK0_p & v8b60ca;
assign v88044e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd86e;
assign v882ae8 = StoB_REQ6_p & v8fd67c | !StoB_REQ6_p & v8a87b1;
assign v882a37 = StoB_REQ6_p & v885f69 | !StoB_REQ6_p & v8fd843;
assign v884735 = jx0_p & v844f9b | !jx0_p & v89735b;
assign v8818ad = jx0_p & v885fe8 | !jx0_p & v892b90;
assign v882c70 = jx2_p & v8b6040 | !jx2_p & !v8fd879;
assign v8fd596 = jx1_p & v896e20 | !jx1_p & v8fd172;
assign v884fa4 = jx0_p & v884256 | !jx0_p & !v885fb8;
assign v8fc18e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8807a6;
assign v8fd5d3 = StoB_REQ1_p & v87af07 | !StoB_REQ1_p & v8819fb;
assign v884870 = jx0_p & v8fd64f | !jx0_p & !v88170c;
assign v8fd88e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd478;
assign v8fc6fe = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v888096;
assign v894722 = jx2_p & v887881 | !jx2_p & !v88793c;
assign v882490 = jx2_p & v8fd5c4 | !jx2_p & v8846ba;
assign v8fd6d6 = StoB_REQ6_p & v885dfd | !StoB_REQ6_p & v844f91;
assign v8816f3 = BtoS_ACK6_p & v88402c | !BtoS_ACK6_p & v8837c5;
assign v8fd851 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fd7aa;
assign v88bb79 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v882a37;
assign v87653c = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd8df;
assign v8ad097 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v89726a;
assign v8845c3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v880dba;
assign v8831c8 = jx1_p & v8811e6 | !jx1_p & v8fd172;
assign v881fdb = RtoB_ACK1_p & v883e9b | !RtoB_ACK1_p & v844f91;
assign v8fd654 = RtoB_ACK0_p & v8fce5c | !RtoB_ACK0_p & v887ac3;
assign v888046 = BtoR_REQ1_p & v8fd7d4 | !BtoR_REQ1_p & v844f91;
assign v887fa9 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & !v853f24;
assign v8fd768 = jx1_p & v8dacfe | !jx1_p & v8fd907;
assign v8fc73e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b607f;
assign v8fc85b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88770c;
assign v8859ec = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd739;
assign v8fd398 = RtoB_ACK1_p & v882c70 | !RtoB_ACK1_p & !v8fd5cd;
assign v88770f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v880bf2;
assign v8ac9cb = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v884904;
assign v8a8734 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd254;
assign v880763 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v895a56;
assign v885a6c = jx0_p & v844f91 | !jx0_p & !v880e00;
assign v895b0b = BtoR_REQ1_p & v8fcdd5 | !BtoR_REQ1_p & v885ddd;
assign v884147 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd808;
assign v88d4df = BtoS_ACK6_p & v8fd1bd | !BtoS_ACK6_p & v880ac4;
assign v8fd893 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v880b2d;
assign v8fd8c9 = RtoB_ACK1_p & v85f322 | !RtoB_ACK1_p & v895abe;
assign v88580d = jx0_p & v8c2eb0 | !jx0_p & v8b5fca;
assign v884adf = jx2_p & v8c2ea3 | !jx2_p & v88372b;
assign v880fd1 = StoB_REQ6_p & v8fd764 | !StoB_REQ6_p & v844f91;
assign v884a73 = BtoR_REQ1_p & v8fd7c2 | !BtoR_REQ1_p & v882db5;
assign v8fc644 = RtoB_ACK0_p & v88294d | !RtoB_ACK0_p & v8809df;
assign v886197 = stateG7_1_p & v894703 | !stateG7_1_p & v8fc9ca;
assign v85cf4b = jx0_p & v8fd5da | !jx0_p & v86ed7e;
assign v8857e9 = jx2_p & v8859f1 | !jx2_p & v88234f;
assign v866b82 = RtoB_ACK0_p & v8fcdd0 | !RtoB_ACK0_p & v8fd881;
assign v8fd1e1 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8c2e5d;
assign v8850e9 = RtoB_ACK0_p & v8fd91a | !RtoB_ACK0_p & v85fc7a;
assign v8fd56f = jx1_p & v8fd6aa | !jx1_p & !v8ad12a;
assign v8cd9e5 = BtoS_ACK6_p & v89471b | !BtoS_ACK6_p & v8fce85;
assign v892ca3 = EMPTY_p & v884058 | !EMPTY_p & v884a71;
assign v8c4cf8 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v887d49;
assign v8fd8c0 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v884476;
assign v88363c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v895bb9;
assign v887a00 = jx0_p & v8fd66a | !jx0_p & v880816;
assign v8fd79f = jx1_p & v881982 | !jx1_p & v868a24;
assign v883c14 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v8822d4;
assign v882b15 = BtoS_ACK1_p & v88029d | !BtoS_ACK1_p & v8fd7e3;
assign v8939a7 = BtoS_ACK6_p & v885df9 | !BtoS_ACK6_p & v890676;
assign v8a87bc = StoB_REQ0_p & v8b5feb | !StoB_REQ0_p & v884626;
assign v8fc2e4 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8837ba;
assign v8808cf = jx0_p & v895a65 | !jx0_p & !v884359;
assign v895d16 = RtoB_ACK0_p & v844fbb | !RtoB_ACK0_p & !v8fd5c7;
assign v8879ab = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v89476c;
assign v885e24 = StoB_REQ1_p & v87653c | !StoB_REQ1_p & v884dec;
assign v8fd865 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ac9cb;
assign v88234e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd8a4;
assign v8fd18d = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v880f9f;
assign v87fb41 = stateG7_1_p & v883b0e | !stateG7_1_p & v844f91;
assign v8877c5 = jx1_p & v8fd221 | !jx1_p & !v8fd598;
assign v882f72 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v881faf;
assign v8fd907 = jx0_p & v87949d | !jx0_p & v880c4c;
assign v88496c = stateG7_1_p & v844f91 | !stateG7_1_p & v87bbad;
assign v887627 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v880638;
assign v8fd83e = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd5ab;
assign v8fcfa9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8847d3;
assign v8828f5 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8818e8;
assign v8fc290 = jx2_p & v887765 | !jx2_p & !v8841f9;
assign v8fd90e = StoB_REQ1_p & v8820ed | !StoB_REQ1_p & v8c2ed0;
assign v8811e6 = jx0_p & v8808eb | !jx0_p & !v895d61;
assign v8fd5e3 = jx1_p & v8fd6ab | !jx1_p & v87bb66;
assign v882e16 = jx0_p & v844f9f | !jx0_p & !v880804;
assign v8762d1 = stateG7_1_p & v8fcd6f | !stateG7_1_p & v8fd788;
assign v8fd886 = BtoR_REQ1_p & v8ac9d6 | !BtoR_REQ1_p & v844fbf;
assign v8fd8a5 = BtoS_ACK0_p & v8c2e72 | !BtoS_ACK0_p & v88618b;
assign v882c83 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v880f23;
assign v883a2e = jx1_p & v887897 | !jx1_p & !v882d73;
assign v8fd6c9 = BtoS_ACK0_p & v8fd84f | !BtoS_ACK0_p & v884bc5;
assign v885a43 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8a704c;
assign v887aee = StoB_REQ2_p & v884904 | !StoB_REQ2_p & v8940fc;
assign v8fd664 = StoB_REQ0_p & v882006 | !StoB_REQ0_p & v8878a5;
assign v88096f = ENQ_p & v8fd848 | !ENQ_p & v8d6a33;
assign v8811ca = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v882d4e;
assign v8f2abb = StoB_REQ6_p & v8fd3c8 | !StoB_REQ6_p & v880d0c;
assign v8fd71c = ENQ_p & v8fd90f | !ENQ_p & v883c3b;
assign v8bb760 = DEQ_p & v844f91 | !DEQ_p & v8fd8fe;
assign v8fd89a = StoB_REQ2_p & v8fca66 | !StoB_REQ2_p & v8a7063;
assign v8fd214 = jx1_p & v882bc8 | !jx1_p & v869327;
assign v8972d8 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v87bb99;
assign v8fd795 = jx0_p & v885063 | !jx0_p & v8825d5;
assign v880834 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v892c5b;
assign v882d6b = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v844faf = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v8fd6cd = jx0_p & v844f91 | !jx0_p & v8fcdd0;
assign v885c0e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8ad0e2;
assign v882852 = jx1_p & v844f91 | !jx1_p & !v885e81;
assign v8fd7bf = FULL_p & v87943e | !FULL_p & v8fd710;
assign v8ce184 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v88fa48;
assign v88376e = RtoB_ACK0_p & v8fd788 | !RtoB_ACK0_p & v8762d1;
assign v882a5a = jx2_p & v8c4d01 | !jx2_p & v87954a;
assign v897386 = jx0_p & v8fd8b8 | !jx0_p & v884ada;
assign v8fc325 = BtoS_ACK6_p & v882baa | !BtoS_ACK6_p & v8846f7;
assign v895d61 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v885694;
assign v8fd5db = jx2_p & v8fd7fc | !jx2_p & !v88791d;
assign v8fce5c = jx2_p & v87fe68 | !jx2_p & !v88791d;
assign v8850ab = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8857aa;
assign v88254d = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v887d06;
assign v8fd6a9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v895a65;
assign v8fd8bc = jx2_p & v8fd5df | !jx2_p & v8fd899;
assign v881099 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9e;
assign v894637 = stateG7_1_p & v8fcfce | !stateG7_1_p & v8fce5c;
assign v8fcc2e = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8fd0e6;
assign v8ac9d2 = BtoS_ACK6_p & v88089e | !BtoS_ACK6_p & v8840af;
assign v883824 = EMPTY_p & v844f91 | !EMPTY_p & v8fc862;
assign v8fd80a = BtoR_REQ0_p & v8838cd | !BtoR_REQ0_p & v8808c9;
assign v86b3d4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v887a7a;
assign v883c48 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v881e80;
assign v880741 = RtoB_ACK0_p & v8fc945 | !RtoB_ACK0_p & v8fca32;
assign v880323 = StoB_REQ3_p & v8fd186 | !StoB_REQ3_p & v882673;
assign v892c64 = StoB_REQ0_p & v882006 | !StoB_REQ0_p & v885185;
assign v889dee = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & !v892c48;
assign v8fd85b = jx1_p & v88fbfc | !jx1_p & !v882bc8;
assign v8816aa = jx2_p & v881ec5 | !jx2_p & v88791d;
assign v87af07 = BtoS_ACK2_p & v882d8f | !BtoS_ACK2_p & v884476;
assign v892416 = StoB_REQ3_p & v8fc1f9 | !StoB_REQ3_p & v844f91;
assign v887d67 = BtoS_ACK6_p & v8fd57d | !BtoS_ACK6_p & v8fd2d5;
assign v8fd5e5 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd3b5;
assign v88033b = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v88058c;
assign BtoR_REQ0_n = !v8ed1f7;
assign v884036 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8f2abb;
assign v885bcf = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8973aa;
assign v8fd84d = stateG7_1_p & v8fd22a | !stateG7_1_p & v8fccad;
assign v8fc982 = jx0_p & v8810a6 | !jx0_p & v88084d;
assign v88193e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v884a91;
assign v880b78 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8fc290;
assign v8a0b36 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v881e54;
assign v8ac9d6 = stateG7_1_p & v844fa5 | !stateG7_1_p & !v844f91;
assign v884df7 = BtoS_ACK0_p & v883759 | !BtoS_ACK0_p & v887dff;
assign v8fd2b7 = BtoR_REQ1_p & v8fc945 | !BtoR_REQ1_p & v895b2f;
assign v882276 = jx2_p & v844f91 | !jx2_p & !v8fd6d7;
assign v88eb87 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v844f99;
assign v883700 = StoB_REQ3_p & v88576e | !StoB_REQ3_p & v844f91;
assign v8f29ed = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8f2a19;
assign v888a80 = BtoS_ACK2_p & v8fd5ad | !BtoS_ACK2_p & v8fc68f;
assign v881117 = jx1_p & v88f397 | !jx1_p & v8827ef;
assign v887f97 = StoB_REQ6_p & v88802b | !StoB_REQ6_p & v844f91;
assign v8fd91b = BtoS_ACK6_p & v8a87b1 | !BtoS_ACK6_p & v880c81;
assign v8fd92a = StoB_REQ0_p & v8fd8a2 | !StoB_REQ0_p & v88bb79;
assign v8807a6 = StoB_REQ0_p & v8877a0 | !StoB_REQ0_p & v883b18;
assign v844f9f = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & !v844f91;
assign v876115 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fd727;
assign v8fd1a4 = StoB_REQ1_p & v8820ed | !StoB_REQ1_p & v8cd9cd;
assign v883cf0 = BtoS_ACK0_p & v8836c4 | !BtoS_ACK0_p & v885660;
assign v8fd7dc = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8840c7;
assign v8fce0d = jx2_p & v8f2a5f | !jx2_p & v8fcba5;
assign v8fd035 = jx0_p & v844f91 | !jx0_p & v8fd683;
assign v882bdd = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9b;
assign v8fc2d4 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v89fb02;
assign v87b4e7 = jx0_p & v883089 | !jx0_p & !v8843ba;
assign v8827e5 = StoB_REQ0_p & v885694 | !StoB_REQ0_p & v844f91;
assign v887913 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v88ebbe;
assign v885e9b = BtoS_ACK1_p & v884476 | !BtoS_ACK1_p & v8fd24d;
assign v8830a2 = BtoR_REQ1_p & v8fd556 | !BtoR_REQ1_p & v8fd7aa;
assign v8fd182 = jx2_p & v88100b | !jx2_p & v8843d0;
assign v89476c = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8fca41;
assign v8fd7e7 = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v887ac6;
assign v880952 = stateG12_p & v88097a | !stateG12_p & v880dc0;
assign v8fc606 = jx2_p & v88426c | !jx2_p & v881117;
assign v882214 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f9d;
assign v8820f2 = stateG7_1_p & v881fa4 | !stateG7_1_p & v8fd8bc;
assign v882505 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v897405;
assign v882d0f = jx1_p & v8fc5a6 | !jx1_p & v88fcc8;
assign v8b5fca = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8840e1;
assign v880240 = jx0_p & v8827ac | !jx0_p & v8843d0;
assign v88507a = BtoS_ACK0_p & v8fccf0 | !BtoS_ACK0_p & !v8dac78;
assign v885748 = StoB_REQ0_p & v8c2ee6 | !StoB_REQ0_p & v882a2c;
assign v88618b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v891077;
assign v88fcc8 = jx0_p & v880487 | !jx0_p & v8fd6bc;
assign v884d53 = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v8fd1e9;
assign v8fd95d = BtoR_REQ0_p & v8fce7b | !BtoR_REQ0_p & v885947;
assign v8810d4 = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v882910;
assign v8843ae = jx0_p & v8fd18e | !jx0_p & v844f91;
assign v8fd755 = BtoR_REQ1_p & v887f6f | !BtoR_REQ1_p & !v8fd5cd;
assign v887765 = jx1_p & v844f91 | !jx1_p & v88257d;
assign v895b2a = StoB_REQ6_p & v844f9d | !StoB_REQ6_p & v885695;
assign v8879a7 = BtoS_ACK6_p & v885d25 | !BtoS_ACK6_p & v8fd68d;
assign v854113 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fc7f4;
assign v887b09 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fca4a;
assign v8fd726 = BtoS_ACK4_p & v88079c | !BtoS_ACK4_p & v888182;
assign v887ca3 = jx0_p & v8ce0f4 | !jx0_p & v887b68;
assign v8825fc = BtoS_ACK6_p & v88089e | !BtoS_ACK6_p & v88101f;
assign v8fce87 = RtoB_ACK1_p & v87bba1 | !RtoB_ACK1_p & v8843d0;
assign v887ad8 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & !v8fcefb;
assign v8877a0 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v883b45;
assign v8fd6a5 = BtoS_ACK6_p & v884476 | !BtoS_ACK6_p & v8d4bf0;
assign v8fd739 = BtoS_ACK6_p & v8fd70d | !BtoS_ACK6_p & v8c2e6c;
assign v884bdd = BtoR_REQ1_p & v897323 | !BtoR_REQ1_p & v8fd688;
assign v8fd594 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd25d;
assign v8ed1e2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88366d;
assign v8948c2 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fcc72;
assign v8fd73a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v8fd7fc = jx1_p & v8676b7 | !jx1_p & v885e81;
assign v8583a8 = stateG7_1_p & v8fc1fa | !stateG7_1_p & v866229;
assign v88186b = BtoS_ACK0_p & v88f618 | !BtoS_ACK0_p & v883c48;
assign v8fd659 = jx2_p & v8fd969 | !jx2_p & v885f5a;
assign v8fd234 = jx2_p & v8fd847 | !jx2_p & v8fd829;
assign v8b606c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88442a;
assign v8ce14d = jx1_p & v8ad131 | !jx1_p & !v884258;
assign v8846ff = jx0_p & v8fd6fc | !jx0_p & v8563aa;
assign v881edd = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v86bd4d;
assign v8fd174 = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v884170;
assign v884136 = jx1_p & v885713 | !jx1_p & !v8ed953;
assign v882baa = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v8fd74e;
assign v8fd642 = BtoS_ACK6_p & v8fd7dc | !BtoS_ACK6_p & v880f66;
assign v8dac30 = BtoS_ACK6_p & v885be7 | !BtoS_ACK6_p & v895b24;
assign v888143 = StoB_REQ6_p & v887c92 | !StoB_REQ6_p & v886188;
assign v8dab99 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f99;
assign v884bc5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd4e2;
assign v895c47 = StoB_REQ1_p & v8ad0e2 | !StoB_REQ1_p & !v8fd5dc;
assign v8fd8fb = RtoB_ACK0_p & v8fd8d7 | !RtoB_ACK0_p & v886197;
assign v8947ed = jx1_p & v844f91 | !jx1_p & !v8fd614;
assign v8ad115 = BtoS_ACK0_p & v8fccf0 | !BtoS_ACK0_p & !v882563;
assign v884875 = StoB_REQ6_p & v890fd8 | !StoB_REQ6_p & v884782;
assign v8817a3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v886129;
assign v8dac5d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd6f9;
assign v887d9a = jx0_p & v882473 | !jx0_p & v8972fa;
assign v887a4a = jx0_p & v89488c | !jx0_p & v844f91;
assign v882f43 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87fee2;
assign v885660 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883ea8;
assign v8b89cf = StoB_REQ6_p & v85582e | !StoB_REQ6_p & !v844f91;
assign v854d12 = RtoB_ACK0_p & v86f4d0 | !RtoB_ACK0_p & v882417;
assign v885bba = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v88190c;
assign v8811b3 = BtoS_ACK6_p & v882baa | !BtoS_ACK6_p & v881657;
assign v88f618 = StoB_REQ6_p & v89471b | !StoB_REQ6_p & v882bdd;
assign v8fd8d7 = jx2_p & v887887 | !jx2_p & !v887d0a;
assign v884206 = BtoS_ACK0_p & v88f9d2 | !BtoS_ACK0_p & v8fc2b8;
assign v8fd176 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v87bb5f;
assign v8b5ff5 = RtoB_ACK0_p & v875cbc | !RtoB_ACK0_p & v885dc6;
assign v8fd65f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v858ace;
assign v8851dd = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fd6f3;
assign v885dfd = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd932;
assign v882417 = BtoR_REQ1_p & v87fed4 | !BtoR_REQ1_p & v898f2f;
assign v8fd817 = StoB_REQ6_p & v844f9b | !StoB_REQ6_p & v894636;
assign v887d5b = jx0_p & v8fc3cf | !jx0_p & v8fd6bc;
assign v8f2a5f = jx1_p & v8dac82 | !jx1_p & !v882d4a;
assign v8fd64f = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8fc295;
assign v8fd770 = BtoR_REQ0_p & v892c49 | !BtoR_REQ0_p & v8fd661;
assign v89facc = jx0_p & v844f91 | !jx0_p & v88582f;
assign v8fc688 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v887f97;
assign v882e00 = jx1_p & v8dabff | !jx1_p & v8879aa;
assign v882a2c = BtoS_ACK6_p & v8fd7dc | !BtoS_ACK6_p & v880674;
assign v88f395 = RtoB_ACK1_p & v887f2c | !RtoB_ACK1_p & v8fd234;
assign v8fd1ac = jx1_p & v887d9a | !jx1_p & v8fd84e;
assign v881fa4 = RtoB_ACK1_p & v8824a9 | !RtoB_ACK1_p & v8fd8bc;
assign v89fadb = jx0_p & v8811aa | !jx0_p & v8fd8a5;
assign v8fd916 = jx2_p & v887f44 | !jx2_p & !v8fd356;
assign v884747 = BtoR_REQ1_p & v8fd1fd | !BtoR_REQ1_p & v887966;
assign v8fd6b2 = jx1_p & v884834 | !jx1_p & !v884206;
assign v8fcac6 = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v8fcb76;
assign v8822bf = jx1_p & v8fd592 | !jx1_p & v8809b9;
assign v8fd5ff = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v882bdd;
assign v8fc61e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v887ad8;
assign v87eaaf = jx2_p & v887f56 | !jx2_p & v844f91;
assign v880d0c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd18b;
assign v8fd7ee = RtoB_ACK1_p & v8810ca | !RtoB_ACK1_p & v8947b9;
assign v8fce6a = jx0_p & v887827 | !jx0_p & v8843d0;
assign v8fd5c4 = jx1_p & v8f2aa3 | !jx1_p & v8846ba;
assign v8fd7d5 = RtoB_ACK1_p & v885d03 | !RtoB_ACK1_p & v883e92;
assign v88506d = jx2_p & v879433 | !jx2_p & v8809eb;
assign v8819ce = StoB_REQ3_p & v8fd5f2 | !StoB_REQ3_p & v844f91;
assign v8fd85f = BtoS_ACK0_p & v8fd70d | !BtoS_ACK0_p & v887e01;
assign v88319e = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v890fd8;
assign v880616 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v880717;
assign v858320 = jx1_p & v8fd6ea | !jx1_p & v88808a;
assign jx1_n = v8a70a6;
assign v8fd7b6 = jx0_p & v883f65 | !jx0_p & v8824ae;
assign v8843d1 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8822d4;
assign v8fd631 = EMPTY_p & v8fd6db | !EMPTY_p & v8fd859;
assign v8825d5 = BtoS_ACK0_p & v885d25 | !BtoS_ACK0_p & v881fdc;
assign v885ec1 = BtoS_ACK0_p & v882d6b | !BtoS_ACK0_p & v890b45;
assign v8fd538 = jx0_p & v844f9f | !jx0_p & !v885144;
assign v887c2f = StoB_REQ3_p & v88576e | !StoB_REQ3_p & v8fd7cb;
assign v8fd86a = StoB_REQ6_p & v880383 | !StoB_REQ6_p & v844f91;
assign v8fd5ee = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v885e9f;
assign v882673 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8fca41;
assign v8fd700 = jx1_p & v8dac82 | !jx1_p & !v8fc982;
assign v8b78a2 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v895a65;
assign v8880e4 = ENQ_p & v8821d3 | !ENQ_p & v8858bb;
assign v88464a = StoB_REQ3_p & v8fc1f9 | !StoB_REQ3_p & v88052d;
assign v8fc934 = BtoS_ACK2_p & v887d93 | !BtoS_ACK2_p & v8fd23f;
assign v884335 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v883d9e;
assign v88315b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd5d4;
assign v890631 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8ad079;
assign v8876ed = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v8fd5a5;
assign v8fc1fe = BtoR_REQ0_p & v886012 | !BtoR_REQ0_p & v887b03;
assign v87fee8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8ad0e2;
assign v88232b = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8fd686;
assign v88275b = StoB_REQ0_p & v8840e1 | !StoB_REQ0_p & v844f91;
assign v8830c5 = RtoB_ACK0_p & v8823c2 | !RtoB_ACK0_p & v8fd788;
assign v8ac1f8 = RtoB_ACK0_p & v8fce0d | !RtoB_ACK0_p & v880c8a;
assign v8fd6d9 = jx2_p & v883a54 | !jx2_p & v88793c;
assign v8fd1e0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd64c;
assign v884c7a = jx2_p & v8856f5 | !jx2_p & !v8881bb;
assign v887a90 = jx2_p & v882ea6 | !jx2_p & v8fd829;
assign v8fd19d = BtoS_ACK2_p & v887d93 | !BtoS_ACK2_p & v8fd81c;
assign v885836 = BtoS_ACK0_p & v8877c1 | !BtoS_ACK0_p & v8ad078;
assign v8f2aa3 = jx0_p & v880341 | !jx0_p & v8846ba;
assign v8847f1 = BtoS_ACK2_p & v8948c3 | !BtoS_ACK2_p & v8fd8e5;
assign v887c1e = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8fd5c7;
assign v8fd782 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd7e8;
assign v883e34 = BtoS_ACK6_p & v882baa | !BtoS_ACK6_p & v8fd222;
assign v887d31 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v895a65;
assign v8fd830 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8fd1ce;
assign v882e37 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd5f9;
assign v8fd8db = EMPTY_p & v8fd7a8 | !EMPTY_p & v8fce04;
assign v8818f6 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v887aee;
assign v885e84 = StoB_REQ3_p & v844fb1 | !StoB_REQ3_p & !v844f91;
assign v8fd260 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & !v8ad0e2;
assign v882905 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v888182;
assign v868d2b = StoB_REQ6_p & v853f24 | !StoB_REQ6_p & !v8fd775;
assign v884421 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v882d8f;
assign v8fd6b5 = RtoB_ACK0_p & v883c24 | !RtoB_ACK0_p & v8810ca;
assign v8fd7c9 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8ac9ad;
assign v8f2abf = DEQ_p & v885c4b | !DEQ_p & v8fd71c;
assign v8fd6ff = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v891ab3;
assign v8fccac = stateG7_1_p & v885d66 | !stateG7_1_p & v8843d0;
assign v8fd90b = BtoR_REQ1_p & v8843d0 | !BtoR_REQ1_p & v8ad009;
assign v88565e = RtoB_ACK1_p & v884adf | !RtoB_ACK1_p & v887b5e;
assign v8fd7a8 = BtoR_REQ0_p & v8fc6ea | !BtoR_REQ0_p & v88579e;
assign v895d68 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v883bb8;
assign v887fd5 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v883879;
assign v884fc8 = BtoS_ACK6_p & v88402c | !BtoS_ACK6_p & v8fd72e;
assign v88172f = jx0_p & v8fd5b1 | !jx0_p & v8fd4a9;
assign v8847e5 = StoB_REQ6_p & v8fd8d5 | !StoB_REQ6_p & v8881be;
assign v8fc7f4 = stateG7_1_p & v8fd916 | !stateG7_1_p & v844f91;
assign v885692 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fca7a;
assign v890b45 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v882d6b;
assign v8878da = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v880665;
assign v8fd8e0 = stateG7_1_p & v885a16 | !stateG7_1_p & v8fd8d0;
assign v8fd5cd = jx2_p & v88483c | !jx2_p & v8fd879;
assign v8808f4 = stateG7_1_p & v879e64 | !stateG7_1_p & v88a5d1;
assign v8fd6e2 = BtoS_ACK1_p & v8fd74e | !BtoS_ACK1_p & v8fd6e1;
assign v88bc53 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v895c47;
assign v884f4a = BtoS_ACK0_p & v883710 | !BtoS_ACK0_p & v8c2de4;
assign v8816be = jx1_p & v8fd6e7 | !jx1_p & v844f91;
assign v8fc42f = StoB_REQ0_p & v85bfad | !StoB_REQ0_p & v8fd705;
assign v897303 = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v891594;
assign v8fd75f = jx2_p & v87b523 | !jx2_p & !v86ed35;
assign v887abd = StoB_REQ0_p & v8851dd | !StoB_REQ0_p & v844f91;
assign v8fd71b = BtoR_REQ0_p & v88499a | !BtoR_REQ0_p & v8844a9;
assign v8878c8 = jx2_p & v89fb10 | !jx2_p & !v844f91;
assign v8828b1 = jx1_p & v883d82 | !jx1_p & !v8dac3a;
assign v8fd5f9 = StoB_REQ0_p & v88514d | !StoB_REQ0_p & v887846;
assign v8f2a18 = stateG12_p & v8818b7 | !stateG12_p & !v8fd860;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v88770c = StoB_REQ0_p & v8877a0 | !StoB_REQ0_p & v887b69;
assign v8839d5 = BtoS_ACK6_p & v8fd57d | !BtoS_ACK6_p & v8857e5;
assign v85879a = BtoS_ACK2_p & v887d93 | !BtoS_ACK2_p & v88fdb7;
assign v844fa1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f91;
assign v8588b1 = BtoS_ACK0_p & v882d6b | !BtoS_ACK0_p & v887d74;
assign v897405 = BtoS_ACK1_p & v885be7 | !BtoS_ACK1_p & v885f78;
assign v887cca = StoB_REQ2_p & v885149 | !StoB_REQ2_p & v8f2a50;
assign v8f2a07 = jx1_p & v8fd6ea | !jx1_p & v8837af;
assign v8fd6c5 = BtoS_ACK2_p & v882d8f | !BtoS_ACK2_p & v854bb9;
assign v880982 = stateG7_1_p & v8fd94b | !stateG7_1_p & !v844f91;
assign v883d9e = StoB_REQ2_p & v8fd5f2 | !StoB_REQ2_p & v844f91;
assign v86a020 = BtoS_ACK0_p & v887c3e | !BtoS_ACK0_p & !v892c64;
assign v885b62 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8fc68f;
assign v8fd1a3 = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v88402c;
assign v8822cf = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v8fd1e7;
assign v8859e8 = jx2_p & v8fced0 | !jx2_p & !v8f2a7d;
assign v898e5c = BtoS_ACK1_p & v88219e | !BtoS_ACK1_p & v8584ff;
assign v8fd74e = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8fd953;
assign v8fd685 = stateG12_p & v88c103 | !stateG12_p & !v8fd609;
assign v85582e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v882fc1;
assign v8876c3 = StoB_REQ6_p & v884796 | !StoB_REQ6_p & v88369c;
assign v8810dc = BtoR_REQ1_p & v884882 | !BtoR_REQ1_p & v8fd90c;
assign v8fcabb = FULL_p & v880643 | !FULL_p & v895cb0;
assign v8fcd6f = RtoB_ACK1_p & v887d8f | !RtoB_ACK1_p & v8fd788;
assign v8fcfe7 = jx0_p & v897358 | !jx0_p & v8ac9bd;
assign v8fd957 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8fd296;
assign v885144 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd66a;
assign v88386a = jx2_p & v8830a5 | !jx2_p & v844f91;
assign v8fcd0e = RtoB_ACK1_p & v8fcedb | !RtoB_ACK1_p & v8fc8ca;
assign v8fd68b = jx1_p & v88401d | !jx1_p & !v8fd5d7;
assign v88040b = BtoS_ACK2_p & v8948c3 | !BtoS_ACK2_p & v8fd8f8;
assign v897358 = BtoS_ACK0_p & v885be7 | !BtoS_ACK0_p & v88a63c;
assign v8fd5ad = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9d;
assign v8fd8c4 = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v8fc67f;
assign v883b0e = RtoB_ACK1_p & v8fd5fd | !RtoB_ACK1_p & v844f91;
assign v868e18 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v883fd7;
assign v8ad05f = stateG7_1_p & v8fd701 | !stateG7_1_p & v8f2a57;
assign v883852 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8fd658;
assign v8c2de4 = StoB_REQ0_p & v8c2ee6 | !StoB_REQ0_p & v879570;
assign v884d67 = StoB_REQ0_p & v8fd856 | !StoB_REQ0_p & v8fd6f2;
assign v885963 = stateG12_p & v8846ba | !stateG12_p & v880a2a;
assign v8fd8b9 = stateG7_1_p & v8fd1a8 | !stateG7_1_p & v8fd8cd;
assign v8a88c6 = stateG12_p & v88a2df | !stateG12_p & v8fd879;
assign v887ac3 = stateG7_1_p & v8f29e5 | !stateG7_1_p & v8f2a57;
assign v8972a7 = jx1_p & v8fd6ea | !jx1_p & v8fccca;
assign v8fd939 = BtoS_ACK1_p & v8fd7dc | !BtoS_ACK1_p & v8fce55;
assign v881a1a = RtoB_ACK0_p & v887bef | !RtoB_ACK0_p & v8fc7b1;
assign v8fd818 = BtoS_ACK0_p & v8c2eaf | !BtoS_ACK0_p & v8cd9b9;
assign v8fd869 = RtoB_ACK0_p & v844fbb | !RtoB_ACK0_p & !v8fd886;
assign v882603 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8fd6ae;
assign SLC1_n = v8dad1a;
assign v8850dd = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v8fd572;
assign v887868 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v880b8e;
assign v8fd6ab = jx0_p & v882bc8 | !jx0_p & v87bb66;
assign v8fd1c7 = jx1_p & v88401d | !jx1_p & v8fd17d;
assign v880507 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v88d29b;
assign v895b58 = stateG12_p & v88bb4f | !stateG12_p & !v88ea59;
assign v88d29b = StoB_REQ2_p & v8dacc2 | !StoB_REQ2_p & v895a71;
assign v89737b = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd7c9;
assign v8fd8c3 = StoB_REQ6_p & v8850ab | !StoB_REQ6_p & v885bf2;
assign v8fc9d3 = jx1_p & v882bc8 | !jx1_p & v887879;
assign v8ed983 = RtoB_ACK0_p & v882490 | !RtoB_ACK0_p & v8f29e2;
assign v8825e5 = StoB_REQ2_p & v882d8f | !StoB_REQ2_p & v844f91;
assign v880bc8 = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v882569;
assign v88089e = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8fd70d;
assign v88785e = BtoS_ACK0_p & v8fd764 | !BtoS_ACK0_p & v8fd1e2;
assign v8817cc = StoB_REQ0_p & v8ad0d9 | !StoB_REQ0_p & v8fc19f;
assign v890676 = BtoS_ACK1_p & v885df9 | !BtoS_ACK1_p & v8fcd1f;
assign v89faf7 = jx1_p & v8fce6a | !jx1_p & v8843d0;
assign v8846bb = ENQ_p & v8fd631 | !ENQ_p & v887656;
assign v88478b = jx0_p & v8fd760 | !jx0_p & !v8fd8b4;
assign v8fc48c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8861c0;
assign v85fc7a = BtoR_REQ1_p & v8ad05f | !BtoR_REQ1_p & v894637;
assign v8fd428 = BtoS_ACK0_p & v882e12 | !BtoS_ACK0_p & v884143;
assign v88f1b0 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v882fc1;
assign v88fdb7 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8f2a19;
assign v88271c = jx0_p & v8f2a3f | !jx0_p & v8fcdd0;
assign v883071 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v88e1fb;
assign v882a0a = jx2_p & v8f11a7 | !jx2_p & v8877e9;
assign v8fd7f2 = jx0_p & v8fc9c2 | !jx0_p & !v8947ee;
assign v8845a8 = jx1_p & v888162 | !jx1_p & v887a00;
assign v8fd5e0 = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v8fd1e0;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v8878ac = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8ce111;
assign v8dac46 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v885bba;
assign v8fd221 = jx0_p & v884256 | !jx0_p & v844f91;
assign v887def = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v880599;
assign v8fd584 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8ad097;
assign v892c48 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v882bdd;
assign v886092 = jx0_p & v8fd95f | !jx0_p & !v884031;
assign v8fd18b = StoB_REQ1_p & v882bee | !StoB_REQ1_p & v881e4b;
assign v8fd921 = jx1_p & v8824d4 | !jx1_p & v8fc7cc;
assign v8ac1f3 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v884d49;
assign v89fb88 = StoB_REQ0_p & v8881e7 | !StoB_REQ0_p & v887fe2;
assign v8880d8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v881ef6;
assign v8fd8a0 = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v88079c;
assign v8fd6f2 = BtoS_ACK6_p & v8fd8c0 | !BtoS_ACK6_p & v882431;
assign v885d67 = jx0_p & v884d11 | !jx0_p & v881ee1;
assign v8fce18 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8ac9d6;
assign v8fd799 = BtoR_REQ1_p & v88fc7a | !BtoR_REQ1_p & v882402;
assign v8a88d6 = DEQ_p & v8836b1 | !DEQ_p & v8876d0;
assign v882066 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88315a;
assign v8fc1cf = BtoS_ACK3_p & v88576e | !BtoS_ACK3_p & v844f9d;
assign v875145 = jx2_p & v8c2ea3 | !jx2_p & v8fd5ed;
assign v888015 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v89830f;
assign v885e9f = BtoS_ACK6_p & v8fd8ba | !BtoS_ACK6_p & v894828;
assign v844fb5 = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & !v844f91;
assign v8fd238 = BtoS_ACK0_p & v885df9 | !BtoS_ACK0_p & v880544;
assign v8fd8cd = jx2_p & v8fd5a6 | !jx2_p & v8831c8;
assign v8fc8ca = jx2_p & v8fd54b | !jx2_p & v8fc6fe;
assign v885d0a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd383;
assign v8fcd29 = BtoS_ACK0_p & v8fd17e | !BtoS_ACK0_p & v8816ff;
assign v8a7071 = StoB_REQ2_p & v8817c2 | !StoB_REQ2_p & v844f91;
assign v880236 = StoB_REQ6_p & v889498 | !StoB_REQ6_p & v8ed1d3;
assign v8fd7cc = StoB_REQ6_p & v882fc1 | !StoB_REQ6_p & v844f91;
assign v87bb76 = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v8fd83c;
assign v8fd742 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v884bc5;
assign v884cde = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v882772;
assign v883f65 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v887fa9;
assign v87fe68 = jx1_p & v8676b7 | !jx1_p & v88397a;
assign v8fd7e4 = jx0_p & v8ce0f4 | !jx0_p & v880c4c;
assign v883c0c = stateG12_p & v8808da | !stateG12_p & v8846ba;
assign v883776 = RtoB_ACK0_p & v86f4d0 | !RtoB_ACK0_p & v87fed4;
assign v88ec21 = BtoS_ACK2_p & v8fd953 | !BtoS_ACK2_p & v8cadd9;
assign v8fc942 = jx1_p & v885a6c | !jx1_p & v8fd59f;
assign v8fd649 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8861c8;
assign v8fd7ed = BtoS_ACK6_p & v89471b | !BtoS_ACK6_p & v8849d3;
assign v8fcb01 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8743a1;
assign v897c49 = RtoB_ACK0_p & v88386a | !RtoB_ACK0_p & v884497;
assign v882217 = StoB_REQ2_p & v8fca66 | !StoB_REQ2_p & v883012;
assign v8fd955 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dabdf;
assign v884882 = stateG7_1_p & v8fd353 | !stateG7_1_p & v8878b5;
assign v8587eb = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88783d;
assign v885026 = jx1_p & v8856e4 | !jx1_p & !v884013;
assign v880294 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a0a29;
assign v880dba = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd185;
assign v8842de = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd6f7;
assign v8fd76a = jx0_p & v886176 | !jx0_p & v89735b;
assign v8fd752 = jx2_p & v8fd714 | !jx2_p & v882ea3;
assign v884a33 = StoB_REQ6_p & v8fd1f3 | !StoB_REQ6_p & v889dee;
assign v8819d6 = BtoS_ACK0_p & v8fd6d6 | !BtoS_ACK0_p & v884531;
assign v8fd6cc = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd7af;
assign v8fd2f7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88417e;
assign v8fd92f = StoB_REQ3_p & v86ed40 | !StoB_REQ3_p & v844f91;
assign v8fc8f1 = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v8fd2a3;
assign v880565 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v894850;
assign v887b14 = BtoS_ACK2_p & v8fd5ad | !BtoS_ACK2_p & v884171;
assign v8fc1bf = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v882217;
assign v892c49 = RtoB_ACK0_p & v891b69 | !RtoB_ACK0_p & v85f322;
assign v883706 = EMPTY_p & v8fd879 | !EMPTY_p & v8a88c6;
assign v8fd8f6 = jx0_p & v883050 | !jx0_p & v844f91;
assign v8fd78d = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8fc1dc;
assign v8fd773 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8881f0;
assign v8fd6f3 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v87d10c;
assign v88404f = jx2_p & v8947da | !jx2_p & v8fcdd0;
assign v88436d = StoB_REQ1_p & v888a80 | !StoB_REQ1_p & v844f91;
assign v87bb66 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8807d3;
assign v891114 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v8ad0e2;
assign v8fd202 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v884216;
assign v890fe3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fcd75;
assign v8ceca9 = BtoS_ACK3_p & v88576e | !BtoS_ACK3_p & v8fc1f9;
assign v897374 = jx1_p & v8fd6ea | !jx1_p & v8dac8a;
assign v883f90 = RtoB_ACK0_p & v8fd1f1 | !RtoB_ACK0_p & !v88386a;
assign v8830bd = BtoR_REQ1_p & v8861a4 | !BtoR_REQ1_p & v844f91;
assign v8fd113 = stateG7_1_p & v8837de | !stateG7_1_p & v854d37;
assign v8847d3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v887d22;
assign v8fd7ba = jx0_p & v88837d | !jx0_p & v884031;
assign v87bacb = StoB_REQ3_p & v8fd6ae | !StoB_REQ3_p & !v8810de;
assign v858501 = jx2_p & v8fd58e | !jx2_p & v8fd596;
assign v8811aa = BtoS_ACK0_p & v8fd6d6 | !BtoS_ACK0_p & v8fd443;
assign v884262 = StoB_REQ0_p & v8fd0b4 | !StoB_REQ0_p & v844f91;
assign v854d37 = jx2_p & v8fc942 | !jx2_p & v88793c;
assign v8fd2a3 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fcfaa;
assign v8fd20f = jx2_p & v885026 | !jx2_p & !v884a26;
assign v88795b = BtoR_REQ0_p & v8ac1f8 | !BtoR_REQ0_p & v8fd6a1;
assign v8881bd = StoB_REQ0_p & v8ed1d8 | !StoB_REQ0_p & v844f91;
assign v8fd5dc = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v882bdd;
assign v883c3b = EMPTY_p & v880403 | !EMPTY_p & v8fd7bf;
assign v8fc6b2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd5e0;
assign v8fd7d3 = RtoB_ACK1_p & v8fd8cd | !RtoB_ACK1_p & v88621e;
assign v885723 = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v8fd672;
assign v8fd349 = jx1_p & v8821e0 | !jx1_p & v8fd5f6;
assign v889757 = EMPTY_p & v8c48b2 | !EMPTY_p & v858a41;
assign v8fd51f = RtoB_ACK0_p & v882e65 | !RtoB_ACK0_p & v8fd5a2;
assign v8fd864 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd1d8;
assign v8fc729 = BtoS_ACK1_p & v88029d | !BtoS_ACK1_p & v8fd8c5;
assign v88164d = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8859f7;
assign v882c78 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v844f91;
assign v880643 = BtoR_REQ0_p & v8fce77 | !BtoR_REQ0_p & v880bb1;
assign v8fd88d = jx0_p & v8fc9d9 | !jx0_p & v890fe3;
assign v88055d = jx2_p & v8ce142 | !jx2_p & v8fc8a5;
assign v8b60d1 = DEQ_p & v8802ff | !DEQ_p & !v8fd761;
assign v885149 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8fd6ae;
assign v883677 = RtoB_ACK0_p & v8fcedb | !RtoB_ACK0_p & v8fc8ca;
assign v844f91 = 1;
assign v8fd5b6 = jx1_p & v885713 | !jx1_p & v88172f;
assign v844fbb = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v844f91;
assign v8fc1fa = RtoB_ACK1_p & v882a0a | !RtoB_ACK1_p & v866229;
assign v8fd7e6 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8838dc;
assign v880487 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88fb6f;
assign v8823a0 = BtoS_ACK0_p & v88493b | !BtoS_ACK0_p & v88ed0c;
assign v8fd667 = StoB_REQ3_p & v8fd947 | !StoB_REQ3_p & v880760;
assign v88107d = BtoR_REQ0_p & v8fd0b7 | !BtoR_REQ0_p & v8810dc;
assign v8d4e0d = StoB_REQ6_p & v885df9 | !StoB_REQ6_p & v880d66;
assign v8fd8ac = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd5e5;
assign v882ea3 = jx1_p & v88313d | !jx1_p & v868a24;
assign v883f84 = StoB_REQ6_p & v8fd865 | !StoB_REQ6_p & v8843b6;
assign v88407b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v884262;
assign v887fc2 = stateG7_1_p & v887a17 | !stateG7_1_p & v882300;
assign v8fd880 = RtoB_ACK1_p & v8fd920 | !RtoB_ACK1_p & v8fd5db;
assign v8fd5e2 = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v8fd966;
assign v8827e6 = stateG7_1_p & v8fd6de | !stateG7_1_p & v8fc7b1;
assign v883759 = StoB_REQ6_p & v885d25 | !StoB_REQ6_p & v885b17;
assign v887f32 = jx0_p & v844f91 | !jx0_p & v8843d0;
assign v884203 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fcd47;
assign v880760 = BtoS_ACK4_p & v878328 | !BtoS_ACK4_p & v844f9d;
assign v8fd8fe = ENQ_p & v8fc862 | !ENQ_p & v883824;
assign v883035 = RtoB_ACK0_p & v8881d4 | !RtoB_ACK0_p & v8fd851;
assign v8fd452 = BtoR_REQ0_p & v88599b | !BtoR_REQ0_p & v885fbe;
assign v884976 = jx0_p & v8ad115 | !jx0_p & v844f91;
assign v885733 = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v887abb;
assign v884a25 = jx0_p & v8fcb01 | !jx0_p & v8fd65b;
assign BtoS_ACK3_n = !v89fb95;
assign v881fdc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v888056;
assign v8810a6 = BtoS_ACK0_p & v883710 | !BtoS_ACK0_p & v8817cc;
assign v8805ad = StoB_REQ6_p & v8850ab | !StoB_REQ6_p & v890676;
assign v884ccb = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v8fc679;
assign BtoS_ACK6_n = !v8a88d6;
assign v853f24 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v884b64 = stateG7_1_p & v8fcd00 | !stateG7_1_p & v8f29e2;
assign v8fd215 = StoB_REQ1_p & v8837fe | !StoB_REQ1_p & v8fd594;
assign v8fd70b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8fd5f2;
assign v8fd5c7 = BtoR_REQ1_p & v8ac9d6 | !BtoR_REQ1_p & v8fd6d4;
assign v8809d1 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v881975;
assign v882170 = BtoR_REQ0_p & v8915ef | !BtoR_REQ0_p & v8fcfc3;
assign v885713 = jx0_p & v88507a | !jx0_p & v844f91;
assign v8dac95 = jx0_p & v887d31 | !jx0_p & v884359;
assign v8c2ed0 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v888a7f;
assign v8fd75b = jx2_p & v8fd349 | !jx2_p & v8fd641;
assign v8f2a5a = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8fd196;
assign v8fc7c3 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8802a9;
assign v844f9e = StoB_REQ4_n & v844f91 | !StoB_REQ4_n & !v844f91;
assign v882d86 = jx1_p & v8fd6cd | !jx1_p & v8fcdd0;
assign v883cd2 = jx1_p & v880b75 | !jx1_p & v8846ba;
assign v8836e8 = StoB_REQ0_p & v858796 | !StoB_REQ0_p & v8fd341;
assign v89fb1e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v882a61;
assign v880c4c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd736;
assign v8fd908 = jx0_p & v844f9b | !jx0_p & v8fd952;
assign v8fd8c1 = jx2_p & v8fd214 | !jx2_p & !v8840d5;
assign v8dacf2 = StoB_REQ2_p & v8fd895 | !StoB_REQ2_p & v882d8f;
assign v8fc312 = jx0_p & v8588b1 | !jx0_p & !v895d61;
assign v88ea59 = BtoR_REQ0_p & v88376e | !BtoR_REQ0_p & v8830c5;
assign v8830a3 = jx1_p & v8fd179 | !jx1_p & v844f91;
assign v8fd7c3 = BtoS_ACK1_p & v8fd74e | !BtoS_ACK1_p & v8fd77d;
assign v882764 = EMPTY_p & v88ea59 | !EMPTY_p & !v895b58;
assign v880c71 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & v8841f8;
assign v885dc6 = jx2_p & v8822fe | !jx2_p & v88793c;
assign v887c6e = BtoS_ACK0_p & v88f618 | !BtoS_ACK0_p & v8fcb1c;
assign v8fd577 = jx0_p & v8fd6c9 | !jx0_p & v882bc8;
assign v8fcbc7 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fc6a5;
assign v885f1e = StoB_REQ2_p & v8fd7f7 | !StoB_REQ2_p & v8fcd77;
assign v8ad133 = DEQ_p & v884d85 | !DEQ_p & v8fd2cf;
assign v8fd8b4 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8847be;
assign v8fd4c4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v892c48;
assign v8fd608 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v885692;
assign v88807f = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v881f1a;
assign v8fd850 = jx1_p & v8fcb09 | !jx1_p & !v8dac95;
assign v8fcfaa = StoB_REQ6_p & v8fd8fa | !StoB_REQ6_p & v887f88;
assign v8f1f45 = jx0_p & v880816 | !jx0_p & v8fc6fe;
assign v881985 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9f;
assign v882910 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dad14;
assign v89488f = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & !v868d2b;
assign v887bbb = StoB_REQ1_p & v8fd57d | !StoB_REQ1_p & v88029d;
assign v8f2aa9 = BtoR_REQ0_p & v883817 | !BtoR_REQ0_p & v897c49;
assign v88280d = StoB_REQ6_p & v8fd786 | !StoB_REQ6_p & v8fd08a;
assign v89fb95 = DEQ_p & v8b60af | !DEQ_p & v882002;
assign v88486a = jx1_p & v887f3f | !jx1_p & v88ed82;
assign v8fce85 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v891e93;
assign v8879aa = jx0_p & v8845c3 | !jx0_p & v88e2d2;
assign v885beb = BtoS_ACK0_p & v882e12 | !BtoS_ACK0_p & v880f35;
assign v887b60 = RtoB_ACK0_p & v882c70 | !RtoB_ACK0_p & !v8fd5cd;
assign v8fc7b7 = jx2_p & v8fd5bf | !jx2_p & !v882f45;
assign v882c30 = jx2_p & v882852 | !jx2_p & v88791d;
assign v883d82 = jx0_p & v892417 | !jx0_p & v86ed7e;
assign v8876bb = BtoR_REQ0_p & v8846bf | !BtoR_REQ0_p & v8daca2;
assign v884de8 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v88201b;
assign v88310a = StoB_REQ1_p & v8ce111 | !StoB_REQ1_p & v8860bd;
assign v8839ba = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v887a7f;
assign v884a6e = jx1_p & v88478b | !jx1_p & !v884cad;
assign v87102d = RtoB_ACK0_p & v8fc57a | !RtoB_ACK0_p & v8816aa;
assign v8816ff = BtoS_ACK6_p & v8fd17e | !BtoS_ACK6_p & v885fb3;
assign v885f4a = BtoR_REQ0_p & v87102d | !BtoR_REQ0_p & v880e10;
assign v8fd786 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd893;
assign v880626 = RtoB_ACK1_p & v884329 | !RtoB_ACK1_p & v866229;
assign v882e64 = jx0_p & v887d31 | !jx0_p & !v844f91;
assign v895a9c = StoB_REQ0_p & v88783d | !StoB_REQ0_p & v8881d6;
assign v8fd794 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v887c6c;
assign v883046 = jx2_p & v8fd930 | !jx2_p & !v8829eb;
assign v8ad0c2 = stateG12_p & v8fd688 | !stateG12_p & !v8fccad;
assign v884035 = jx0_p & v8fd8eb | !jx0_p & v844f91;
assign v880f23 = StoB_REQ0_p & v882006 | !StoB_REQ0_p & !v844f91;
assign v883cfc = RtoB_ACK1_p & v8816aa | !RtoB_ACK1_p & v8fc945;
assign v8fd77b = jx0_p & v883f65 | !jx0_p & !v8ce165;
assign v8fd63f = BtoR_REQ0_p & v854ae6 | !BtoR_REQ0_p & v884747;
assign v860216 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8839ba;
assign v8fd5eb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c48b3;
assign v88785b = BtoS_ACK0_p & v882fd7 | !BtoS_ACK0_p & v882093;
assign v8fd657 = jx1_p & v8824d4 | !jx1_p & !v8fd17d;
assign BtoS_ACK5_n = !v8ad133;
assign v8fd6a8 = stateG7_1_p & v8ce18c | !stateG7_1_p & v884316;
assign v894924 = BtoR_REQ0_p & v881a1a | !BtoR_REQ0_p & v8fd4e0;
assign v8846ba = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd20b;
assign v8824dc = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v86ed40;
assign v884448 = jx0_p & v87949d | !jx0_p & v887b68;
assign v88ed0c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc8d5;
assign v8fd6aa = jx0_p & v844f91 | !jx0_p & v880816;
assign v8802a4 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v88258c;
assign v8fced0 = jx1_p & v8676b7 | !jx1_p & v888662;
assign v885d03 = jx2_p & v8806f0 | !jx2_p & v8843d0;
assign v887e01 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c2e4a;
assign v8821e0 = jx0_p & v844f91 | !jx0_p & v8827ac;
assign v884585 = jx1_p & v8856e4 | !jx1_p & !v8fd7f2;
assign v882d4a = jx0_p & v884f4a | !jx0_p & v88251e;
assign v8816ab = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v880d42;
assign v894671 = BtoR_REQ0_p & v882de0 | !BtoR_REQ0_p & v8fc644;
assign v883fee = jx0_p & v8fd782 | !jx0_p & v88e2d2;
assign v8fd7c8 = StoB_REQ6_p & v88eb87 | !StoB_REQ6_p & v8fd764;
assign v8fd20a = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v887cca;
assign v8ce1ae = jx1_p & v885a6c | !jx1_p & v8974c9;
assign v8fd556 = stateG7_1_p & v8844d6 | !stateG7_1_p & v87eaaf;
assign v885e59 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v895c47;
assign v8584ff = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v888a80;
assign v88574b = BtoS_ACK2_p & v8fd953 | !BtoS_ACK2_p & v8fd89a;
assign v8fd467 = EMPTY_p & v887c95 | !EMPTY_p & v858a41;
assign v8805d7 = FULL_p & v8f2a18 | !FULL_p & v8c2ebb;
assign v8803e6 = StoB_REQ0_p & v888096 | !StoB_REQ0_p & v895a39;
assign v8840e1 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8831ee;
assign v8c2eb8 = jx0_p & v881113 | !jx0_p & v844f91;
assign v883b45 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd15f;
assign v8fd574 = jx0_p & v8b603b | !jx0_p & v87bb66;
assign v8fd6e7 = jx0_p & v844f91 | !jx0_p & !v895d61;
assign v8910ad = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v88079c;
assign v8fc5e1 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8fd218;
assign v8fd1e9 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd77e;
assign v8d6a33 = stateG12_p & v8fd4e5 | !stateG12_p & !v884f1f;
assign v8fd84e = BtoS_ACK0_p & v8fd5c9 | !BtoS_ACK0_p & v88945f;
assign v87feab = stateG7_1_p & v8fd29a | !stateG7_1_p & v89243a;
assign v8fce12 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v888015;
assign v886176 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v88800a;
assign v88f397 = jx0_p & v8849ca | !jx0_p & v882cf9;
assign v890cdc = StoB_REQ0_p & v8fd957 | !StoB_REQ0_p & v844f91;
assign v887d8f = jx2_p & v8fd7b2 | !jx2_p & !v884a6e;
assign v887b68 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v884577;
assign v8fd002 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v882214;
assign v8fd633 = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v8850dd;
assign v8fd69d = jx1_p & v8856e4 | !jx1_p & !v87001c;
assign v8fd8dd = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f99;
assign v85397c = stateG7_1_p & v880b78 | !stateG7_1_p & v8fc290;
assign v8b6088 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8fc3e8;
assign v8fd6b4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd868;
assign v882a61 = StoB_REQ0_p & v8fd1e1 | !StoB_REQ0_p & v8b605d;
assign v880750 = jx0_p & v887c6e | !jx0_p & v884df7;
assign v8fd7b1 = BtoR_REQ0_p & v884292 | !BtoR_REQ0_p & v8d4782;
assign v8876f2 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fcbc7;
assign v8fd15f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8fd7f7;
assign v8fd22e = jx0_p & v8587eb | !jx0_p & !v844f9d;
assign v8819b3 = StoB_REQ0_p & v8876f2 | !StoB_REQ0_p & v8fd8ab;
assign v880eac = RtoB_ACK0_p & v8fd8c1 | !RtoB_ACK0_p & v8fd1aa;
assign v853f4e = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v88810b;
assign v8fd6ea = jx0_p & v88507a | !jx0_p & v892b90;
assign v883ea8 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd7cc;
assign v895d4e = RtoB_ACK0_p & v88616c | !RtoB_ACK0_p & v88772e;
assign v8897a6 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v880c0e;
assign v86ed40 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v88576e;
assign v8fd655 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8fd1f9;
assign v8ad0d9 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v892c36;
assign v87bb99 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v89484f;
assign v8823f5 = RtoB_ACK1_p & v8896fd | !RtoB_ACK1_p & v887966;
assign v8fca41 = StoB_REQ4_p & v844f9f | !StoB_REQ4_p & v844f91;
assign v8848a0 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8dab99;
assign v884941 = BtoR_REQ0_p & v882024 | !BtoR_REQ0_p & v8fd5fc;
assign v8879a4 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fc42f;
assign v8fc19f = BtoS_ACK6_p & v8fd57d | !BtoS_ACK6_p & v89fb74;
assign v895bb9 = BtoS_ACK6_p & v884476 | !BtoS_ACK6_p & v8fd24e;
assign v887f3f = jx0_p & v883d79 | !jx0_p & v8825d5;
assign v8fcbd7 = BtoS_ACK6_p & v8fd629 | !BtoS_ACK6_p & v8fd871;
assign v88fc61 = RtoB_ACK0_p & v8fd75f | !RtoB_ACK0_p & v8fd230;
assign v8fd6be = jx1_p & v8676b7 | !jx1_p & v884035;
assign v8fd8e5 = StoB_REQ2_p & v88464a | !StoB_REQ2_p & v8fd19b;
assign v8fd6c1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v881048;
assign v8dab8a = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v8fd6ff;
assign v8fd930 = jx1_p & v8fd6ea | !jx1_p & v8fd236;
assign v8fd873 = BtoS_ACK6_p & v8fd70d | !BtoS_ACK6_p & v882c31;
assign v8fd967 = jx2_p & v8fd5df | !jx2_p & !v844f91;
assign v884f1f = jx2_p & v8fd5df | !jx2_p & v8591df;
assign v895b52 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8fc8ad;
assign v890cff = StoB_REQ3_p & v883852 | !StoB_REQ3_p & v844fb3;
assign v8fcfc3 = BtoR_REQ1_p & v87ff08 | !BtoR_REQ1_p & v844f91;
assign v883e11 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8dab99;
assign v8fd951 = StoB_REQ3_p & v8fd186 | !StoB_REQ3_p & v884170;
assign v880e10 = BtoR_REQ1_p & v8fd58f | !BtoR_REQ1_p & v8fc945;
assign v8fd665 = jx1_p & v885713 | !jx1_p & v88580d;
assign v854c61 = stateG7_1_p & v880626 | !stateG7_1_p & v866229;
assign v89475e = BtoS_ACK6_p & v885ab0 | !BtoS_ACK6_p & v8fd1b9;
assign v8fd849 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd775;
assign v8838dc = StoB_REQ0_p & v8fd856 | !StoB_REQ0_p & v883a94;
assign v882cf9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v860216;
assign v8fd5d1 = jx0_p & v882fda | !jx0_p & v8539e7;
assign v880cd6 = jx0_p & v8f2a14 | !jx0_p & v8fd428;
assign v882b4a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v895afe;
assign v8fcdd0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd6ec;
assign v8858e2 = StoB_REQ3_p & v884904 | !StoB_REQ3_p & v844fb3;
assign v8fd29a = RtoB_ACK1_p & v8fd182 | !RtoB_ACK1_p & v89243a;
assign v88190c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v88058c;
assign v884197 = stateG7_1_p & v8880e0 | !stateG7_1_p & v88a5d1;
assign v8fd777 = jx2_p & v8fd5df | !jx2_p & v8830a3;
assign v8fd1bb = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fce12;
assign v8fd71e = StoB_REQ6_p & v8fd6f9 | !StoB_REQ6_p & v844f91;
assign v87afd1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8819b3;
assign v8c48b7 = BtoS_ACK2_p & v844f9e | !BtoS_ACK2_p & v881099;
assign v8fd8a4 = BtoS_ACK2_p & v8fd646 | !BtoS_ACK2_p & v8c4cf8;
assign v8770c9 = jx1_p & v8818fb | !jx1_p & v8dac0f;
assign v8fd746 = StoB_REQ6_p & v8fd67c | !StoB_REQ6_p & v884476;
assign v887f6f = stateG7_1_p & v8fd398 | !stateG7_1_p & !v8fd5cd;
assign v8fd54e = RtoB_ACK0_p & v88404f | !RtoB_ACK0_p & v880d9c;
assign v8f2a03 = jx2_p & v8540de | !jx2_p & v8fd084;
assign v8f29e5 = RtoB_ACK1_p & v8fc9ca | !RtoB_ACK1_p & v8f2a57;
assign v882b84 = RtoB_ACK0_p & v8843d0 | !RtoB_ACK0_p & v8fccac;
assign v8fd714 = jx1_p & v883f96 | !jx1_p & v887ca3;
assign v8844a9 = BtoR_REQ1_p & v87feab | !BtoR_REQ1_p & v89243a;
assign v88ea40 = jx2_p & v8fd6c6 | !jx2_p & v8fd281;
assign v887cf6 = jx1_p & v88380c | !jx1_p & v8846ba;
assign v883685 = jx1_p & v8fc5a6 | !jx1_p & v880c3a;
assign v8844ce = jx0_p & v8a8734 | !jx0_p & v844f91;
assign v8821b5 = BtoS_ACK1_p & v8fd932 | !BtoS_ACK1_p & v8840b0;
assign v8809df = BtoR_REQ1_p & v854c61 | !BtoR_REQ1_p & v858acb;
assign v887bbe = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8819fb;
assign v885d66 = RtoB_ACK1_p & v879581 | !RtoB_ACK1_p & v8843d0;
assign v8fd23f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8fd8cf;
assign v887846 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v88777d;
assign v88fdb8 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8836e8;
assign v880263 = StoB_REQ6_p & v8842de | !StoB_REQ6_p & v881018;
assign v8b5fbd = jx1_p & v8fd908 | !jx1_p & v88fa9e;
assign v88fbfc = jx0_p & v844f9b | !jx0_p & !v882bc8;
assign v88489f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f9b;
assign v884718 = jx0_p & v882b4a | !jx0_p & !v844f9d;
assign v8c008e = jx0_p & v882093 | !jx0_p & v8827ac;
assign v8816cc = jx0_p & v880614 | !jx0_p & v844f91;
assign v8fd5e8 = stateG7_1_p & v881923 | !stateG7_1_p & v88621e;
assign DEQ_n = !v8bb760;
assign v8b5ffa = StoB_REQ6_p & v8fd8e4 | !StoB_REQ6_p & v8fd7c3;
assign v854d5c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8831e6;
assign v882699 = StoB_REQ6_p & v883b45 | !StoB_REQ6_p & v885b21;
assign v86ef5c = BtoS_ACK6_p & v8fd853 | !BtoS_ACK6_p & v8818d7;
assign v88237c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc9f1;
assign v881f61 = BtoR_REQ1_p & v885c06 | !BtoR_REQ1_p & !v844f91;
assign v8fc295 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8fc2e4;
assign v881ef6 = StoB_REQ0_p & v8a87de | !StoB_REQ0_p & v844f91;
assign v8fd620 = StoB_REQ0_p & v8847be | !StoB_REQ0_p & v880a73;
assign v87b523 = jx1_p & v8fd6ea | !jx1_p & v88fdf5;
assign v8b5fc7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8878bd;
assign v8fd788 = jx2_p & v8fd657 | !jx2_p & !v884a6e;
assign v8973aa = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v880982;
assign v8802a9 = StoB_REQ6_p & v8879eb | !StoB_REQ6_p & v844f91;
assign v8fc1d2 = BtoR_REQ0_p & v886048 | !BtoR_REQ0_p & v8fd5b3;
assign v8842ac = RtoB_ACK1_p & v8c2eb4 | !RtoB_ACK1_p & !v88386a;
assign v8ed1ca = StoB_REQ1_p & v8820ed | !StoB_REQ1_p & v895ce5;
assign v8fd62e = RtoB_ACK0_p & v8c2ecf | !RtoB_ACK0_p & !v88386a;
assign v892417 = BtoS_ACK0_p & v844fa1 | !BtoS_ACK0_p & !v8944a2;
assign v8fd443 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc7c3;
assign v8fd7e3 = StoB_REQ1_p & v880665 | !StoB_REQ1_p & v88040b;
assign v8fd678 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v880abb;
assign v880a70 = BtoS_ACK1_p & v8fd5ad | !BtoS_ACK1_p & v887f3a;
assign v880a73 = BtoS_ACK6_p & v885b17 | !BtoS_ACK6_p & v8fd93c;
assign v88241f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v885e84;
assign v88093b = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8fd5ad;
assign v8fcc77 = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v8fd1a1;
assign v8fd86e = BtoS_ACK1_p & v885be7 | !BtoS_ACK1_p & v8fd607;
assign v8fd629 = StoB_REQ1_p & v8fd24b | !StoB_REQ1_p & v844f91;
assign v8fd91d = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8ce1b0;
assign v8fc5c1 = RtoB_ACK1_p & v883e2e | !RtoB_ACK1_p & v8fd5a2;
assign v87001c = jx0_p & v8fd91d | !jx0_p & !v883f7a;
assign v88499a = RtoB_ACK0_p & v8fd182 | !RtoB_ACK0_p & v89243a;
assign v881657 = StoB_REQ6_p & v8fd8e4 | !StoB_REQ6_p & v8fd039;
assign v8fd7c7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v884e81;
assign v8fd83c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v887d9c;
assign v882f82 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd813;
assign v887c95 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8fd72c;
assign v880af8 = stateG7_1_p & v8819df | !stateG7_1_p & v844f91;
assign v8dac78 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8878a5;
assign v8fd589 = BtoS_ACK1_p & v884476 | !BtoS_ACK1_p & v8fd6c5;
assign v8fc1f8 = stateG7_1_p & v8ed1a5 | !stateG7_1_p & v844f91;
assign v881e4b = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v882b96;
assign v8fd7a7 = BtoR_REQ1_p & v8878c8 | !BtoR_REQ1_p & v858acb;
assign v8fd5b7 = stateG7_1_p & v882c77 | !stateG7_1_p & v880d9c;
assign v882300 = jx2_p & v883cd2 | !jx2_p & v8846ba;
assign v8fd6d1 = BtoS_ACK3_p & v8fca41 | !BtoS_ACK3_p & !v844f91;
assign v866229 = jx2_p & v884136 | !jx2_p & v8fd36d;
assign v8fd602 = RtoB_ACK1_p & v8fd5fd | !RtoB_ACK1_p & v8fc290;
assign v883719 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8879a7;
assign v8fc484 = BtoR_REQ1_p & v8843d0 | !BtoR_REQ1_p & v8fd740;
assign v8fd6d8 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v884b6c;
assign v88ec29 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8fd923;
assign v8847e2 = jx1_p & v8676b7 | !jx1_p & v8816cc;
assign v8fcefb = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8fd5dc;
assign v8fd00a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v883700;
assign v8fd71a = BtoR_REQ0_p & v8fd8b7 | !BtoR_REQ0_p & v8c993e;
assign v8fd609 = BtoR_REQ0_p & v8fd654 | !BtoR_REQ0_p & v8850e9;
assign v8947b9 = jx2_p & v8fcfe8 | !jx2_p & v844f91;
assign v89241d = jx2_p & v8fd6be | !jx2_p & !v8fc2e5;
assign v88294d = BtoR_REQ1_p & v882a0a | !BtoR_REQ1_p & v866229;
assign v881e67 = jx0_p & v8819d6 | !jx0_p & v8fd2ab;
assign v885cf3 = ENQ_p & v8fd8af | !ENQ_p & v880a21;
assign v88108f = StoB_REQ1_p & v8ac9cb | !StoB_REQ1_p & v8fd1db;
assign v89830f = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v879434;
assign v8837de = RtoB_ACK1_p & v885dc6 | !RtoB_ACK1_p & v854d37;
assign v8b6040 = jx1_p & v8fd1ea | !jx1_p & !v8fd879;
assign v895a39 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8846fc;
assign v88800a = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v887bf3;
assign v8dace1 = BtoR_REQ1_p & v8846ba | !BtoR_REQ1_p & v887fc2;
assign v880d9c = jx2_p & v882d86 | !jx2_p & v8fcdd0;
assign v8827ac = BtoS_ACK0_p & v882e12 | !BtoS_ACK0_p & v882093;
assign v8fd1f3 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v883791;
assign v8fc801 = RtoB_ACK0_p & v8fd91a | !RtoB_ACK0_p & v887ade;
assign v8f2a50 = StoB_REQ3_p & v8fd6ae | !StoB_REQ3_p & v885149;
assign v8fd358 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd5ae;
assign v887f56 = jx1_p & v844f91 | !jx1_p & !v8805c4;
assign v8fd011 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fc5a3;
assign v8b5ff4 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v858acd;
assign v889498 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v885d08;
assign jx2_n = v8c4d26;
assign v887adb = BtoS_ACK6_p & v884e81 | !BtoS_ACK6_p & v883ee4;
assign v884796 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8fd78e;
assign v88793c = jx1_p & v8fd82a | !jx1_p & v8fd6c3;
assign v8f2aa5 = StoB_REQ0_p & v8ad0d9 | !StoB_REQ0_p & v885b87;
assign v8f2a57 = jx2_p & v8fd733 | !jx2_p & !v88791d;
assign v885ea3 = BtoR_REQ0_p & v87bb66 | !BtoR_REQ0_p & v894721;
assign v8fd836 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fd8e4;
assign v8fd18e = BtoS_ACK0_p & v8fd1a3 | !BtoS_ACK0_p & v8fd8c4;
assign v8fd5ae = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dac53;
assign v8676b7 = jx0_p & v844f91 | !jx0_p & !v844f91;
assign v887a17 = RtoB_ACK1_p & v8846ba | !RtoB_ACK1_p & v882300;
assign v87dfe7 = StoB_REQ6_p & v883b45 | !StoB_REQ6_p & v881018;
assign v8fd72c = BtoR_REQ1_p & v8ac9d6 | !BtoR_REQ1_p & v887cd8;
assign v8fc9f1 = BtoS_ACK6_p & v880d66 | !BtoS_ACK6_p & v884b83;
assign v879433 = jx1_p & v8dacfe | !jx1_p & v8fd7e4;
assign v8fd8b8 = BtoS_ACK0_p & v8fd629 | !BtoS_ACK0_p & v885b81;
assign v885931 = jx2_p & v8fc246 | !jx2_p & v88486a;
assign v885f78 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8811a0;
assign v883e1c = stateG7_1_p & v882484 | !stateG7_1_p & v8fd6d9;
assign v8e1d28 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v887644;
assign v8fc6aa = RtoB_ACK1_p & v8fd62f | !RtoB_ACK1_p & v8fc945;
assign v88101f = StoB_REQ6_p & v8831ee | !StoB_REQ6_p & v88096b;
assign v883c78 = jx0_p & v8fcac6 | !jx0_p & v844f91;
assign v885fe3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd379;
assign v8fd185 = BtoS_ACK6_p & v885be7 | !BtoS_ACK6_p & v88044e;
assign v885ee1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ed1e2;
assign v8fd5d4 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9d;
assign v883791 = StoB_REQ1_p & v892c48 | !StoB_REQ1_p & !v844f91;
assign v880b5b = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8878bb;
assign v8fd17b = jx2_p & v89fb10 | !jx2_p & !v88e7c3;
assign v8fd55c = RtoB_ACK1_p & v8fd218 | !RtoB_ACK1_p & v844f91;
assign v880e00 = BtoS_ACK0_p & v844fa1 | !BtoS_ACK0_p & v8587bf;
assign v8ce111 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8fd951;
assign v8fd95c = jx2_p & v8f2a07 | !jx2_p & !v8fd1af;
assign v8fd8c5 = StoB_REQ1_p & v8fd6ff | !StoB_REQ1_p & v8847f1;
assign v844fa0 = StoB_REQ5_n & v844f91 | !StoB_REQ5_n & !v844f91;
assign v8c2eb4 = jx2_p & v8828b1 | !jx2_p & !v890d96;
assign v885947 = RtoB_ACK0_p & v88294d | !RtoB_ACK0_p & v8fd7a7;
assign v8825e6 = BtoR_REQ0_p & v883f90 | !BtoR_REQ0_p & v881f61;
assign v88212e = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v882603;
assign v883817 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v88225a;
assign v882048 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8fd002;
assign v885d0d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v854bb9;
assign v8fd70f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v895b92;
assign v883762 = jx1_p & v8fd221 | !jx1_p & v844f91;
assign v8fd7be = ENQ_p & v8fd1de | !ENQ_p & v8fd7ca;
assign v88284b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8fd584;
assign v8fd0b4 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8794e0;
assign v8fd5a4 = StoB_REQ0_p & v8881e7 | !StoB_REQ0_p & v8fd805;
assign v8fd651 = ENQ_p & v844fab | !ENQ_p & !v880769;
assign v8fd285 = BtoR_REQ1_p & v8820f2 | !BtoR_REQ1_p & v8824a9;
assign v8fcfe8 = jx1_p & v844f91 | !jx1_p & v8fd22e;
assign v8c2e4a = BtoS_ACK6_p & v8fd70d | !BtoS_ACK6_p & v8fd163;
assign v8fd5b2 = jx1_p & v880752 | !jx1_p & v868a24;
assign v8daca2 = RtoB_ACK0_p & v88386a | !RtoB_ACK0_p & v887734;
assign v8fcc62 = jx0_p & v844f9f | !jx0_p & !v8fc4c0;
assign v887d06 = BtoR_REQ1_p & v8ac9d6 | !BtoR_REQ1_p & v88496c;
assign v8857aa = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v885df9;
assign v88254c = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v882fc1;
assign v8a87f2 = jx0_p & v8fd6e3 | !jx0_p & v8fcdd0;
assign v887fc7 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v895abe;
assign v8a70a6 = DEQ_p & v882b76 | !DEQ_p & !v882507;
assign v884031 = BtoS_ACK0_p & v8fccf0 | !BtoS_ACK0_p & !v8cd9b9;
assign v883f8f = jx0_p & v844f91 | !jx0_p & v880341;
assign v88174e = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd8a2;
assign v858422 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v883eb1;
assign v883e2e = jx2_p & v8fd914 | !jx2_p & v884a6e;
assign v882507 = ENQ_p & v85841e | !ENQ_p & v8fce1f;
assign v844fab = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v8894e3 = jx0_p & v8fd8eb | !jx0_p & !v87feba;
assign v85b93e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8860d7;
assign v8fcbe3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88567a;
assign v884bcc = jx0_p & v854bab | !jx0_p & !v8823a0;
assign v8fd1db = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v887629;
assign v884e03 = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v880e69;
assign v8fd79b = RtoB_ACK1_p & v895abe | !RtoB_ACK1_p & v844f91;
assign v8ad074 = BtoS_ACK4_p & v88576e | !BtoS_ACK4_p & v8841f8;
assign v8fd922 = jx0_p & v88785e | !jx0_p & v8fd243;
assign v887a78 = BtoR_REQ0_p & v887b60 | !BtoR_REQ0_p & v8fd755;
assign v8837c5 = StoB_REQ6_p & v8fd7af | !StoB_REQ6_p & v8fd72e;
assign v8fc237 = StoB_REQ6_p & v8fc21f | !StoB_REQ6_p & v882431;
assign v887ccd = RtoB_ACK0_p & v8fd6d9 | !RtoB_ACK0_p & v8fd113;
assign v8820ed = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v885909;
assign v86e414 = StoB_REQ0_p & v8877a0 | !StoB_REQ0_p & v8fd23a;
assign v884d47 = jx1_p & v884a25 | !jx1_p & v885b36;
assign v8fd599 = ENQ_p & v885963 | !ENQ_p & v87d828;
assign v8fd570 = StoB_REQ6_p & v8fd78e | !StoB_REQ6_p & v895c47;
assign v88fb6f = StoB_REQ0_p & v8ad0d9 | !StoB_REQ0_p & v885de9;
assign v888162 = jx0_p & v8fd5e2 | !jx0_p & v8946a5;
assign v8fd7fd = RtoB_ACK0_p & v8fc1cd | !RtoB_ACK0_p & v86deca;
assign v8c2e5d = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v87653c;
assign v882fda = BtoS_ACK0_p & v88f618 | !BtoS_ACK0_p & v880cf5;
assign v85e9fa = jx0_p & v8fd655 | !jx0_p & v8dab62;
assign v887cde = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88b623;
assign v884f81 = BtoS_ACK6_p & v8fd8ba | !BtoS_ACK6_p & v880763;
assign v885ffa = RtoB_ACK0_p & v875145 | !RtoB_ACK0_p & v8fd8cd;
assign v883f96 = jx0_p & v844f91 | !jx0_p & v882c83;
assign v8fd0b7 = RtoB_ACK0_p & v884c7a | !RtoB_ACK0_p & v8878b5;
assign v8818d7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8831a1;
assign v88e2d2 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd22d;
assign v8fd7b5 = BtoR_REQ1_p & v883928 | !BtoR_REQ1_p & v844f91;
assign v8fd637 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v881e33;
assign v844fb1 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v887d49 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v88fa1c;
assign v8fd1c5 = BtoS_ACK6_p & v89471b | !BtoS_ACK6_p & v885c76;
assign v8806f0 = jx1_p & v89fb26 | !jx1_p & v8fcd8f;
assign v8fd222 = StoB_REQ6_p & v8fd8fa | !StoB_REQ6_p & v8fd7c3;
assign v8fd1af = jx1_p & v882b85 | !jx1_p & v886092;
assign v884cea = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v885d0a;
assign v88e1fb = BtoS_ACK4_p & v883c06 | !BtoS_ACK4_p & v888182;
assign v88ec23 = BtoR_REQ1_p & v894722 | !BtoR_REQ1_p & v8fd82e;
assign v8fd243 = BtoS_ACK0_p & v8fd7c8 | !BtoS_ACK0_p & v883752;
assign v880933 = stateG7_1_p & v85839b | !stateG7_1_p & v88386a;
assign v885695 = BtoS_ACK1_p & v884476 | !BtoS_ACK1_p & v87af07;
assign v8861c8 = StoB_REQ3_p & v86ed40 | !StoB_REQ3_p & v8fd7cb;
assign v88483c = jx1_p & v884a9c | !jx1_p & v8fd879;
assign v880599 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8840c5;
assign v858678 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v88496e;
assign v880e69 = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v8811b3;
assign v885e81 = jx0_p & v884e03 | !jx0_p & v844f91;
assign v8fd196 = StoB_REQ3_p & v883852 | !StoB_REQ3_p & v8fd658;
assign v887a7c = ENQ_p & v887c1e | !ENQ_p & v88254d;
assign v8809b9 = jx0_p & v88265b | !jx0_p & v844f91;
assign v8fd859 = stateG12_p & v8fd5c8 | !stateG12_p & v8fd6db;
assign v88369f = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v895bb6;
assign v8fd87d = StoB_REQ1_p & v8fcd1f | !StoB_REQ1_p & v8857aa;
assign v880f9f = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v880cff;
assign v8fd64a = BtoR_REQ0_p & v881944 | !BtoR_REQ0_p & v8fd7b5;
assign v89fb10 = jx1_p & v8fd6ea | !jx1_p & v8826bd;
assign v885684 = stateG7_1_p & v881141 | !stateG7_1_p & v8fce5c;
assign v880cf5 = StoB_REQ0_p & v8fd0b4 | !StoB_REQ0_p & v8fd796;
assign v8831a1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v88436d;
assign v887f88 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fd90e;
assign v8fd58c = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8fd18d;
assign v8dac0f = jx0_p & v8fd232 | !jx0_p & !v885119;
assign v8fd4e5 = jx2_p & v844f91 | !jx2_p & !v8591df;
assign v8fccf0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8fd764;
assign v869e2c = jx1_p & v882bc8 | !jx1_p & v8fc28a;
assign v8fc986 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fc19e;
assign v882fc1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8ad0e2;
assign v882719 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd5f5;
assign v88493b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8fd8ba;
assign v88576e = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v844f9f;
assign v882d4e = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v880ab4;
assign v8fd7d4 = stateG7_1_p & v8848b0 | !stateG7_1_p & v8fd659;
assign v884b56 = jx0_p & v8fd014 | !jx0_p & v8972d8;
assign v895b02 = jx0_p & v885fe3 | !jx0_p & v885836;
assign v88315a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88397d;
assign v8fd8ea = EMPTY_p & v87bb66 | !EMPTY_p & v8fd195;
assign v8fccad = jx2_p & v8847e2 | !jx2_p & !v8fc2e5;
assign v88085d = StoB_REQ6_p & v890fd8 | !StoB_REQ6_p & v8fd039;
assign v8fd5dd = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v884d5a;
assign v8fcd32 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd86a;
assign v8915ef = RtoB_ACK0_p & v864119 | !RtoB_ACK0_p & v8fd5fd;
assign v8fd90d = jx1_p & v885f7b | !jx1_p & v8c008e;
assign v884dca = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v8fd5f2;
assign v8880da = jx0_p & v844f91 | !jx0_p & !v844fab;
assign v8c48b2 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v895d16;
assign v884cad = jx0_p & v8809c4 | !jx0_p & !v8ce165;
assign v885f26 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v895aff;
assign v884cd5 = StoB_REQ6_p & v882431 | !StoB_REQ6_p & v885b96;
assign v8fd571 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v895cec;
assign v8fd860 = BtoR_REQ0_p & v8fd60e | !BtoR_REQ0_p & v8808c9;
assign v8818e1 = jx0_p & v88318b | !jx0_p & v884cea;
assign v854830 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fd903;
assign v88bc54 = stateG12_p & v8825da | !stateG12_p & !v8ac9b2;
assign v888a7f = StoB_REQ2_p & v885909 | !StoB_REQ2_p & v888bbe;
assign v8f2abd = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8fd88a;
assign v885fbe = RtoB_ACK0_p & v884bdd | !RtoB_ACK0_p & v8fd688;
assign v8ce18c = RtoB_ACK1_p & v87bb66 | !RtoB_ACK1_p & v884316;
assign v883f9f = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd842;
assign v8fd20e = jx0_p & v8811ca | !jx0_p & v883f1b;
assign v88565d = jx2_p & v885da7 | !jx2_p & !v887d85;
assign v8fd8d6 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fad;
assign v88235e = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v88e43b;
assign v8fd5d7 = jx0_p & v8fcd29 | !jx0_p & v881649;
assign v8881d6 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v858a9b;
assign v89fac8 = RtoB_ACK0_p & v88616c | !RtoB_ACK0_p & v876115;
assign v8fd039 = BtoS_ACK1_p & v8fd74e | !BtoS_ACK1_p & v8fd1a4;
assign v8fd8ab = BtoS_ACK6_p & v88402c | !BtoS_ACK6_p & v876549;
assign v895d4b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8828f5;
assign v85841e = EMPTY_p & v882d74 | !EMPTY_p & !v8fccd5;
assign v8fc9d9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v89fb46;
assign v8a8729 = jx2_p & v8fd68b | !jx2_p & !v8fd877;
assign v8fd22d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd873;
assign v887adf = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v868e18;
assign v8fd710 = BtoR_REQ0_p & v8816e8 | !BtoR_REQ0_p & v895d4e;
assign v8fd958 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88275b;
assign v8fd7ac = RtoB_ACK0_p & v8fd920 | !RtoB_ACK0_p & v8fc9ca;
assign v88029d = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8948c3;
assign v8fd73b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v894dfc;
assign v8fca66 = StoB_REQ3_p & v8fd726 | !StoB_REQ3_p & v86bd4d;
assign v8fd1a8 = RtoB_ACK1_p & v875145 | !RtoB_ACK1_p & v8fd8cd;
assign v884258 = jx0_p & v887fa9 | !jx0_p & !v8fd5fa;
assign v887c60 = stateG7_1_p & v887a90 | !stateG7_1_p & v8fd659;
assign v881982 = jx0_p & v882186 | !jx0_p & v8fd85c;
assign v8fd717 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fcbd7;
assign v884531 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fcd32;
assign v8fd641 = jx1_p & v8586ec | !jx1_p & v8fd8f6;
assign v88802b = BtoS_ACK1_p & v8fd932 | !BtoS_ACK1_p & v8c48b6;
assign v8fd1d8 = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8fd734;
assign v8fc9ca = jx2_p & v8fd59c | !jx2_p & !v88791d;
assign v8fd857 = RtoB_ACK0_p & v882d68 | !RtoB_ACK0_p & v8a8783;
assign v8a7063 = StoB_REQ3_p & v8fd726 | !StoB_REQ3_p & v88079c;
assign v887904 = jx2_p & v887f44 | !jx2_p & !v8b5fbd;
assign v892b90 = BtoS_ACK0_p & v8fccf0 | !BtoS_ACK0_p & !v8fd664;
assign v884907 = RtoB_ACK1_p & v882859 | !RtoB_ACK1_p & v887dae;
assign v8fd1da = StoB_REQ6_p & v85582e | !StoB_REQ6_p & !v88807f;
assign v8fd4e0 = BtoR_REQ1_p & v8fd1d6 | !BtoR_REQ1_p & v844f91;
assign v8831ee = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v884421;
assign v895a65 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & v87ff04;
assign v880c3a = jx0_p & v8fc3cf | !jx0_p & v8850da;
assign v8fd903 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v883bef;
assign v88589c = jx2_p & v8fd612 | !jx2_p & !v8fd7f4;
assign v8539e7 = BtoS_ACK0_p & v883759 | !BtoS_ACK0_p & v8fd620;
assign v880769 = EMPTY_p & v8fd64a | !EMPTY_p & v8878e0;
assign v881963 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8fc708;
assign v8dac3a = jx0_p & v882d19 | !jx0_p & v8fd8a5;
assign v8fd829 = jx1_p & v883a3f | !jx1_p & !v881f75;
assign v8836c4 = StoB_REQ6_p & v88eb87 | !StoB_REQ6_p & v844f91;
assign v858ace = StoB_REQ0_p & v8fd260 | !StoB_REQ0_p & v844f91;
assign v88fc7a = stateG7_1_p & v887fc7 | !stateG7_1_p & v895abe;
assign v8806a6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v86ef60;
assign v8fd929 = StoB_REQ6_p & v8fd8d5 | !StoB_REQ6_p & v88604b;
assign v880648 = BtoR_REQ1_p & v8810ca | !BtoR_REQ1_p & v8947b9;
assign v887ce9 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8fd3c8;
assign v8fd661 = BtoR_REQ1_p & v8fd51b | !BtoR_REQ1_p & v844f91;
assign v881018 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8f2a80;
assign v8b5feb = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v889498;
assign v8fc6ea = RtoB_ACK0_p & v883b53 | !RtoB_ACK0_p & v8827e6;
assign v887dc2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b6053;
assign v8fd6ae = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9d;
assign v88e2ce = jx2_p & v8fd693 | !jx2_p & !v8fd7f4;
assign v88578e = BtoS_ACK6_p & v884476 | !BtoS_ACK6_p & v895b2a;
assign v8fd877 = jx1_p & v884735 | !jx1_p & v88fa9e;
assign v8810ca = jx2_p & v881022 | !jx2_p & v883158;
assign v8fc719 = jx0_p & v88369f | !jx0_p & !v883f7a;
assign v880abb = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v882bdd;
assign v8fcb09 = jx0_p & v88164d | !jx0_p & !v8896c7;
assign v8fc970 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8f2a2c;
assign v887827 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v883b45;
assign v8fd68d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v884796;
assign v887bfb = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v8878c5;
assign v8fd729 = BtoS_ACK6_p & v8fd629 | !BtoS_ACK6_p & v8847a4;
assign v89488c = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v880db3;
assign v8810de = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8fd6ae;
assign v885863 = jx0_p & v8809c4 | !jx0_p & v8ce165;
assign v88fa9e = jx0_p & v887fa9 | !jx0_p & !v8ce165;
assign v881e54 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cd9e5;
assign v887d0a = jx1_p & v8fd179 | !jx1_p & v882e64;
assign v883ad4 = BtoS_ACK0_p & v8fd8c0 | !BtoS_ACK0_p & v884d67;
assign v887dff = StoB_REQ0_p & v8fd260 | !StoB_REQ0_p & v8fd244;
assign v885b96 = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v890ce8;
assign v86ed36 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v885dfd;
assign v8fd180 = BtoS_ACK6_p & v8fd629 | !BtoS_ACK6_p & v8fd88e;
assign v883ed8 = BtoS_ACK6_p & v8fd5ff | !BtoS_ACK6_p & !v880e82;
assign v884d5a = StoB_REQ2_p & v8fca66 | !StoB_REQ2_p & v8856c1;
assign v87bb5f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd64c;
assign v883710 = StoB_REQ6_p & v887bbb | !StoB_REQ6_p & v8fd57d;
assign v879434 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v884dca;
assign v885c06 = stateG7_1_p & v8842ac | !stateG7_1_p & !v88386a;
assign v844f9d = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v844f91;
assign v8fd5c8 = BtoR_REQ0_p & v882b84 | !BtoR_REQ0_p & v8946de;
assign v887dae = jx2_p & v883685 | !jx2_p & !v882f45;
assign v880231 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v885fce;
assign v8ad078 = StoB_REQ0_p & v8fd856 | !StoB_REQ0_p & v8fd741;
assign v8fd636 = stateG7_1_p & v8fd7d3 | !stateG7_1_p & v88621e;
assign v88769d = BtoS_ACK6_p & v88315b | !BtoS_ACK6_p & v885a43;
assign v8fd6ec = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd866;
assign v887f44 = jx1_p & v88401d | !jx1_p & !v8846ff;
assign v8829eb = jx1_p & v890ce6 | !jx1_p & v8844ce;
assign v8daba0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v881f1a;
assign v8fd666 = jx1_p & v884a6d | !jx1_p & v87bb66;
assign v8fd843 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8fd627;
assign v88fd1c = StoB_REQ2_p & v885909 | !StoB_REQ2_p & v88112f;
assign v887ade = BtoR_REQ1_p & v8fce5c | !BtoR_REQ1_p & v894637;
assign v8fcba4 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v883f84;
assign v8877fe = FULL_p & v8fd95d | !FULL_p & v894671;
assign v8fd12b = RtoB_ACK0_p & v880eda | !RtoB_ACK0_p & v8fccad;
assign v880638 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8fd002;
assign v8f2a19 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v88052d;
assign v891ab3 = StoB_REQ2_p & v88464a | !StoB_REQ2_p & v892416;
assign v882c16 = jx1_p & v8fd72b | !jx1_p & !v844fab;
assign v8fd0e6 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v88058c;
assign v8fd5c9 = StoB_REQ6_p & v844f97 | !StoB_REQ6_p & v844f91;
assign v8fc246 = jx1_p & v880341 | !jx1_p & v897386;
assign v887c98 = jx0_p & v844f91 | !jx0_p & v8fc6fe;
assign v8fcb76 = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v883e34;
assign v887efe = stateG7_1_p & v8c4d0d | !stateG7_1_p & v8fd688;
assign v882788 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8838c5;
assign v8fc8d5 = BtoS_ACK6_p & v8fd8ba | !BtoS_ACK6_p & v88284b;
assign v8ce150 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc688;
assign v8fd0a4 = BtoS_ACK1_p & v8fd57d | !BtoS_ACK1_p & v8fd8b1;
assign v88496e = StoB_REQ2_p & v8822d4 | !StoB_REQ2_p & v884b6c;
assign v8ed1ce = BtoR_REQ1_p & v8773cf | !BtoR_REQ1_p & v844f91;
assign v8fcc72 = stateG7_1_p & v8fd55c | !stateG7_1_p & v844f91;
assign v8944a2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v882006;
assign v8989c5 = BtoR_REQ1_p & v885dc6 | !BtoR_REQ1_p & v854d37;
assign v88390f = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v88306a;
assign v883d79 = BtoS_ACK0_p & v89471b | !BtoS_ACK0_p & v887cde;
assign v88084d = BtoS_ACK0_p & v8fd746 | !BtoS_ACK0_p & v8fd917;
assign v854c1c = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v887fd5;
assign v8841bc = BtoS_ACK0_p & v8fd7dc | !BtoS_ACK0_p & v8f2aa5;
assign v8fd1c9 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v892416;
assign v887734 = BtoR_REQ1_p & v880933 | !BtoR_REQ1_p & v88225a;
assign v884329 = jx2_p & v8fd665 | !jx2_p & !v844f91;
assign v8850d3 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8dacbf;
assign v8fd77e = BtoS_ACK1_p & v882214 | !BtoS_ACK1_p & v8fd64c;
assign v887d86 = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v884335;
assign v894dfc = BtoS_ACK1_p & v8fd73a | !BtoS_ACK1_p & v8ad097;
assign v8fc732 = BtoS_ACK6_p & v885b17 | !BtoS_ACK6_p & v881172;
assign v8fd2ab = BtoS_ACK0_p & v8c2e72 | !BtoS_ACK0_p & v895b93;
assign v883bef = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v8dacc2;
assign v854bab = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8fd0b4;
assign v88fb91 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fd649;
assign v885bf2 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd87d;
assign v8fd255 = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8dac5d;
assign v8fce1f = EMPTY_p & v887cfa | !EMPTY_p & !v8a88d5;
assign v8fd327 = BtoR_REQ0_p & v8fd62e | !BtoR_REQ0_p & v885c13;
assign v887881 = jx1_p & v8856e4 | !jx1_p & !v8fc719;
assign v8fd179 = jx0_p & v88164d | !jx0_p & v844f91;
assign v858a9b = BtoS_ACK1_p & v8879ab | !BtoS_ACK1_p & v887657;
assign v88219e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8fd5ad;
assign v8fd7f3 = jx1_p & v8676b7 | !jx1_p & v8fd3fc;
assign v8fd341 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v88118b;
assign v8fd088 = stateG7_1_p & v8fd967 | !stateG7_1_p & v844f91;
assign v8fd600 = ENQ_p & v8fd58b | !ENQ_p & v8fc1d2;
assign v8fd353 = RtoB_ACK1_p & v884c7a | !RtoB_ACK1_p & v8878b5;
assign v8824d8 = jx1_p & v883f96 | !jx1_p & v884448;
assign v884867 = BtoR_REQ0_p & v887b5a | !BtoR_REQ0_p & v883035;
assign v8811a0 = StoB_REQ2_p & v8fd8cf | !StoB_REQ2_p & v844f91;
assign v8c2ee6 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd724;
assign v8972fa = BtoS_ACK0_p & v8836c4 | !BtoS_ACK0_p & v887dc2;
assign v882186 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v882c78;
assign v882c77 = RtoB_ACK1_p & v88404f | !RtoB_ACK1_p & v880d9c;
assign v897323 = jx2_p & v887f83 | !jx2_p & v8fc2e5;
assign v8881be = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8c4d03;
assign v8f2a80 = StoB_REQ1_p & v8fd15f | !StoB_REQ1_p & v8b5ff4;
assign v8946bb = stateG7_1_p & v88595e | !stateG7_1_p & v844f91;
assign v89463b = BtoS_ACK0_p & v885d25 | !BtoS_ACK0_p & v8fd955;
assign v887bf3 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v882b6f;
assign v884cc3 = StoB_REQ0_p & v88783d | !StoB_REQ0_p & v8ed18b;
assign v880544 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8939a7;
assign v881ee1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v890cdc;
assign v887b15 = jx2_p & v858320 | !jx2_p & !v8822bf;
assign v8fd5f6 = jx0_p & v882b4a | !jx0_p & !v885119;
assign v88579b = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v880abb;
assign v8fd7e9 = stateG12_p & v8fd879 | !stateG12_p & !v887a78;
assign v887629 = StoB_REQ2_p & v884904 | !StoB_REQ2_p & v8858e2;
assign v8fd6c3 = jx0_p & v8b78a2 | !jx0_p & !v884359;
assign v8fce5e = jx2_p & v8824d8 | !jx2_p & v882ea3;
assign v8fc77f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd202;
assign v881048 = StoB_REQ1_p & v887b14 | !StoB_REQ1_p & v844f91;
assign v879b9f = stateG7_1_p & v858501 | !stateG7_1_p & v8fd8cd;
assign v8845a2 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v88219e;
assign v8fd80f = BtoS_ACK1_p & v8fd002 | !BtoS_ACK1_p & v8fd64c;
assign v8fd232 = BtoS_ACK0_p & v8fd1bd | !BtoS_ACK0_p & v895a9c;
assign v8fd90c = stateG7_1_p & v8fd6b6 | !stateG7_1_p & v8878b5;
assign v8fd8ff = StoB_REQ6_p & v8fd3b5 | !StoB_REQ6_p & v8fd163;
assign v88c127 = BtoS_ACK6_p & v882d6b | !BtoS_ACK6_p & v8fd7b7;
assign v8cd9b9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v89488f;
assign v8fc862 = BtoR_REQ0_p & v8fd94f | !BtoR_REQ0_p & !v887906;
assign v886188 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fd215;
assign v8c2e6b = RtoB_ACK0_p & v880648 | !RtoB_ACK0_p & v895cb4;
assign v8859bf = jx0_p & v885ee1 | !jx0_p & v8820a0;
assign v8846f7 = StoB_REQ6_p & v8fd8d5 | !StoB_REQ6_p & v8fd6e2;
assign v8fc5a3 = StoB_REQ0_p & v854830 | !StoB_REQ0_p & v882bb8;
assign v88046c = BtoR_REQ1_p & v8fd5fd | !BtoR_REQ1_p & v8fc290;
assign v8fc1cd = jx2_p & v8fd83b | !jx2_p & !v8fd850;
assign v8821d3 = stateG12_p & v8843d0 | !stateG12_p & v8fd71b;
assign v8fc1dc = stateG7_1_p & v8851ef | !stateG7_1_p & v8fd218;
assign v8fce55 = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v883700;
assign v8858bb = BtoR_REQ0_p & v8fd6b5 | !BtoR_REQ0_p & v884953;
assign v89fb26 = jx0_p & v8fc85b | !jx0_p & v8843d0;
assign v88426c = jx1_p & v88fbd1 | !jx1_p & !v882e16;
assign v854be6 = BtoS_ACK0_p & v844fa1 | !BtoS_ACK0_p & !v88945f;
assign v86ef60 = BtoS_ACK1_p & v8fd5d4 | !BtoS_ACK1_p & v8fd637;
assign v8fd812 = jx2_p & v87b523 | !jx2_p & !v8881bb;
assign v8fcb1c = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v887fec;
assign v884a26 = jx1_p & v89726c | !jx1_p & v8808cf;
assign v8806c7 = StoB_REQ0_p & v885694 | !StoB_REQ0_p & v8fc732;
assign v8fd761 = ENQ_p & v882764 | !ENQ_p & v8fd928;
assign v8fd1d6 = stateG7_1_p & v87dfc7 | !stateG7_1_p & v8fc7b1;
assign v883b53 = jx2_p & v883837 | !jx2_p & v884f6d;
assign v8fd239 = BtoR_REQ1_p & v87bb66 | !BtoR_REQ1_p & v8fd6a8;
assign v880816 = BtoS_ACK0_p & v884565 | !BtoS_ACK0_p & v8fd66a;
assign v8c2ea3 = jx1_p & v8f2a3f | !jx1_p & v885077;
assign v8881e7 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fd8d5;
assign v88e5f0 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fd088;
assign v8fd3fc = jx0_p & v8fd833 | !jx0_p & v844f91;
assign v8fcc49 = jx1_p & v844f91 | !jx1_p & v8fc296;
assign v8fd24b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v887d93;
assign v8877e9 = jx1_p & v8fd20e | !jx1_p & !v884ba1;
assign v8b6054 = RtoB_ACK1_p & v8fc57a | !RtoB_ACK1_p & v882c30;
assign v895ce3 = BtoR_REQ0_p & v883677 | !BtoR_REQ0_p & v881e44;
assign v88318b = BtoS_ACK0_p & v8fd1a3 | !BtoS_ACK0_p & v880bb6;
assign v88595e = RtoB_ACK1_p & v8810ca | !RtoB_ACK1_p & v844f91;
assign v8fd713 = jx0_p & v880b07 | !jx0_p & !v882e37;
assign v8fd6bd = jx2_p & v8fcf10 | !jx2_p & !v892325;
assign v88112f = StoB_REQ3_p & v888182 | !StoB_REQ3_p & v8fca41;
assign v880b07 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fd5a4;
assign v8fd705 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v888143;
assign v8859af = FULL_p & v8fc1fe | !FULL_p & v884b4e;
assign v8dab62 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8fcbb4;
assign v859713 = stateG7_1_p & v88068f | !stateG7_1_p & v8878c8;
assign v8fd607 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a7071;
assign v880b2d = StoB_REQ2_p & v8fd5f2 | !StoB_REQ2_p & v8ac9ad;
assign v882ac1 = jx0_p & v8587eb | !jx0_p & !v885119;
assign v8fc68e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v883a7f;
assign v8fc21f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd6d8;
assign v882473 = BtoS_ACK0_p & v880fd1 | !BtoS_ACK0_p & v880b56;
assign v8c2e72 = StoB_REQ6_p & v884ac0 | !StoB_REQ6_p & v844f91;
assign v8fd57d = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8840c7;
assign v8fd952 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v885f76;
assign v8fd648 = stateG7_1_p & v8fd751 | !stateG7_1_p & v8859e8;
assign v8fc76f = StoB_REQ2_p & v885909 | !StoB_REQ2_p & v8fd7e7;
assign v8826bd = jx0_p & v87afd1 | !jx0_p & v8fd70f;
assign v8fd953 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v8fca41;
assign v88fa1c = BtoS_ACK3_p & v88576e | !BtoS_ACK3_p & v8ad074;
assign v8fd965 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8876f2;
assign v880ab4 = BtoS_ACK6_p & v882bdd | !BtoS_ACK6_p & v8fd817;
assign v8861f9 = BtoS_ACK2_p & v8fd17e | !BtoS_ACK2_p & v8fd816;
assign v8d4782 = RtoB_ACK0_p & v882d68 | !RtoB_ACK0_p & v8fd799;
assign v883aae = RtoB_ACK0_p & v885931 | !RtoB_ACK0_p & v887c60;
assign v88251a = BtoR_REQ0_p & v8b5ff5 | !BtoR_REQ0_p & v880d9a;
assign v882484 = RtoB_ACK1_p & v885dc6 | !RtoB_ACK1_p & v8fd6d9;
assign v887cd8 = stateG7_1_p & v844f91 | !stateG7_1_p & v8a8729;
assign v8fd5d2 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fd836;
assign v883eb1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v874ed6;
assign v887897 = jx0_p & v8fd64f | !jx0_p & !v8fcd30;
assign v8fd8af = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v88e5f0;
assign v8fd808 = BtoS_ACK1_p & v8fd002 | !BtoS_ACK1_p & v885ab0;
assign v8f2a7d = jx1_p & v8c2eb8 | !jx1_p & !v885b3a;
assign v8856d5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd91b;
assign v882d19 = BtoS_ACK0_p & v8fd6d6 | !BtoS_ACK0_p & v8ce150;
assign v888062 = RtoB_ACK1_p & v8fc290 | !RtoB_ACK1_p & v844f91;
assign v898e61 = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v8822cf;
assign v8fd1a1 = StoB_REQ1_p & v8fc6a5 | !StoB_REQ1_p & v880665;
assign v887c3e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8fd5ff;
assign v8827b2 = stateG7_1_p & v895c60 | !stateG7_1_p & v844f91;
assign v895abb = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8fd4f5;
assign v8836b1 = ENQ_p & v8fd7e9 | !ENQ_p & !v8fd327;
assign v8fd588 = jx1_p & v883d82 | !jx1_p & !v881e67;
assign v882f45 = jx1_p & v884870 | !jx1_p & !v897301;
assign v880614 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8b5feb;
assign v8fd848 = stateG12_p & v882276 | !stateG12_p & !v8b6045;
assign v882c31 = StoB_REQ6_p & v8fd3b5 | !StoB_REQ6_p & v887d86;
assign v8fd879 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fb7;
assign v883d05 = StoB_REQ1_p & v8897a6 | !StoB_REQ1_p & v884482;
assign v8fd686 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v88f0b3;
assign v8fd6e6 = StoB_REQ6_p & v8878ac | !StoB_REQ6_p & v884cde;
assign v89726c = jx0_p & v881113 | !jx0_p & !v885fb8;
assign v8f2a0b = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v89737b;
assign v8ce1b0 = StoB_REQ0_p & v858796 | !StoB_REQ0_p & v8fcf73;
assign v87fee2 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd71e;
assign v8fd6d4 = stateG7_1_p & v844f91 | !stateG7_1_p & v8fd967;
assign v881172 = StoB_REQ6_p & v891114 | !StoB_REQ6_p & v88369c;
assign v86ec4a = jx0_p & v8b605e | !jx0_p & v8857fb;
assign v8fc691 = jx1_p & v880e79 | !jx1_p & v8fc182;
assign v8856f6 = RtoB_ACK0_p & v8fccad | !RtoB_ACK0_p & v8fd84d;
assign v8fd5cc = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd68f;
assign v8fd197 = stateG7_1_p & v8c2df5 | !stateG7_1_p & !v88386a;
assign v8fd4a9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a705e;
assign v8840d5 = jx1_p & v884bcc | !jx1_p & !v8fd577;
assign v890ce6 = jx0_p & v884c5a | !jx0_p & v884464;
assign v8856e4 = jx0_p & v844f91 | !jx0_p & v880e00;
assign v890d96 = jx1_p & v8fd8f3 | !jx1_p & !v854be6;
assign v8fd242 = jx1_p & v883f96 | !jx1_p & v8fd907;
assign v882b85 = jx0_p & v895ccc | !jx0_p & v880f76;
assign v8fd87b = stateG7_1_p & v8806a9 | !stateG7_1_p & v844f91;
assign v8fd918 = jx1_p & v8880da | !jx1_p & !v844fab;
assign v8fd7a0 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v8fd678;
assign v8fd1ce = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v884b89;
assign v8fd5fa = BtoS_ACK0_p & v8fc5ad | !BtoS_ACK0_p & v892156;
assign v8841f8 = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v8fd2a7;
assign v8856f5 = jx1_p & v8818ad | !jx1_p & v88fdf5;
assign v883cf7 = RtoB_ACK0_p & v8ad047 | !RtoB_ACK0_p & v879b9f;
assign v8fd658 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9d;
assign v8843ba = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd793;
assign v8878c5 = StoB_REQ0_p & v8881e7 | !StoB_REQ0_p & v8fc325;
assign v8881fb = BtoS_ACK1_p & v884476 | !BtoS_ACK1_p & v8fd7ff;
assign v8825da = BtoR_REQ0_p & v880741 | !BtoR_REQ0_p & v882034;
assign v8fd3cb = BtoS_ACK6_p & v8fd8c0 | !BtoS_ACK6_p & v8fd23e;
assign v8fd6f7 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844fb1;
assign v88963d = RtoB_ACK1_p & v88808c | !RtoB_ACK1_p & v88a5d1;
assign v887b03 = RtoB_ACK0_p & v887baf | !RtoB_ACK0_p & v8948c2;
assign v891b69 = jx2_p & v8fd768 | !jx2_p & v8fd79f;
assign v887f83 = jx1_p & v844f91 | !jx1_p & !v884035;
assign v8fd747 = jx1_p & v844f91 | !jx1_p & !v8fc802;
assign v880bf2 = BtoS_ACK6_p & v880d66 | !BtoS_ACK6_p & v8fd8c3;
assign v8642ea = jx0_p & v8879a4 | !jx0_p & !v8fd1d2;
assign v8fd595 = ENQ_p & v88fcc6 | !ENQ_p & v887f70;
assign v8ed1a5 = RtoB_ACK1_p & v8fd8cd | !RtoB_ACK1_p & v844f91;
assign v892325 = jx1_p & v8c2eb8 | !jx1_p & !v8fd598;
assign v885215 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8f29ed;
assign v8fd5fd = jx2_p & v882d0f | !jx2_p & !v87debc;
assign v881f4a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v880bc8;
assign v8fd22a = RtoB_ACK1_p & v89241d | !RtoB_ACK1_p & v8fccad;
assign v8fd5a8 = stateG12_p & v8fd5a2 | !stateG12_p & !v8fd788;
assign v8fd6e1 = StoB_REQ1_p & v8fd597 | !StoB_REQ1_p & v88574b;
assign v89243a = jx2_p & v895d18 | !jx2_p & v8843d0;
assign v8ed1f7 = DEQ_p & v885cf3 | !DEQ_p & v8fd595;
assign v8c98e7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883d20;
assign v8fd1f1 = jx2_p & v8fd588 | !jx2_p & !v88429a;
assign v8896c7 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8ed1b3;
assign v88497c = BtoS_ACK0_p & v86ed36 | !BtoS_ACK0_p & v8fd7cf;
assign v8824a9 = jx2_p & v8fd5df | !jx2_p & v883762;
assign v8857fb = BtoS_ACK0_p & v887c3e | !BtoS_ACK0_p & !v8fc2b8;
assign v89735b = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8fd260;
assign v88582f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd8ac;
assign v887f13 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8fc651;
assign v8fca7a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8810bc;
assign v8fd853 = StoB_REQ1_p & v88219e | !StoB_REQ1_p & v844f91;
assign v883089 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v88319e;
assign v8fd610 = StoB_REQ6_p & v8ac9e4 | !StoB_REQ6_p & v88bc53;
assign v8fd8d1 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fd28e;
assign v8fcff6 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v883719;
assign v8824ae = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v892156;
assign v880bb1 = RtoB_ACK0_p & v880648 | !RtoB_ACK0_p & v8fd7de;
assign v8fd920 = jx2_p & v887887 | !jx2_p & !v88791d;
assign v880f9a = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd63c;
assign v880341 = BtoS_ACK0_p & v8fc5ad | !BtoS_ACK0_p & v8817a3;
assign v8fd872 = StoB_REQ3_p & v8fd186 | !StoB_REQ3_p & v89736f;
assign v8849ea = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8a87de;
assign v8fcedb = jx2_p & v884034 | !jx2_p & v8fc6fe;
assign v8fd926 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd717;
assign v8fd6f9 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v8fd764;
assign v895cec = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8588b8;
assign v8808da = BtoR_REQ0_p & v8846ba | !BtoR_REQ0_p & v885ee9;
assign v8fd65e = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v881985;
assign v8841eb = BtoS_ACK6_p & v885be7 | !BtoS_ACK6_p & v882505;
assign v8dad1a = DEQ_p & v8fd600 | !DEQ_p & v8fd7be;
assign v8dacc2 = StoB_REQ3_p & v881985 | !StoB_REQ3_p & !v8fd65e;
assign v8f2a3f = BtoS_ACK0_p & v8fd7c7 | !BtoS_ACK0_p & v883bb8;
assign v887f67 = jx0_p & v8827ac | !jx0_p & v885beb;
assign v882402 = stateG7_1_p & v8fd79b | !stateG7_1_p & v844f91;
assign v882bf5 = StoB_REQ1_p & v880abb | !StoB_REQ1_p & v844f91;
assign v884ba1 = jx0_p & v8fd1d7 | !jx0_p & v844f91;
assign v880db3 = StoB_REQ0_p & v88319e | !StoB_REQ0_p & v8805dc;
assign v882024 = RtoB_ACK0_p & v8fc6fe | !RtoB_ACK0_p & v8859d2;
assign v854ae6 = RtoB_ACK0_p & v8896fd | !RtoB_ACK0_p & v887966;
assign v8fd881 = BtoR_REQ1_p & v8fcdd0 | !BtoR_REQ1_p & v8fd33e;
assign v884920 = BtoR_REQ0_p & v8fd7fd | !BtoR_REQ0_p & v895b0b;
assign v887d74 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88c127;
assign v891da3 = EMPTY_p & v8825e6 | !EMPTY_p & !v8fd704;
assign v894636 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v8fd5dc;
assign v8fd77a = jx0_p & v8ad08b | !jx0_p & !v844f9d;
assign v8948bb = stateG7_1_p & v882841 | !stateG7_1_p & v8947b9;
assign v8823d8 = jx1_p & v8a87f2 | !jx1_p & v8fcdd0;
assign v8587bf = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v844fa1;
assign v881944 = RtoB_ACK0_p & v88a4a0 | !RtoB_ACK0_p & v88083d;
assign v880fe9 = RtoB_ACK1_p & v88621e | !RtoB_ACK1_p & v844f91;
assign v883e9b = jx2_p & v8795bb | !jx2_p & !v844f91;
assign v88064f = BtoR_REQ0_p & v8fd7ac | !BtoR_REQ0_p & v8fd251;
assign v89484f = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v882a63;
assign v8fc692 = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v8818e8;
assign v8fd014 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fd8d1;
assign v8fd81c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8817c2;
assign v8cd9cd = BtoS_ACK2_p & v8fd953 | !BtoS_ACK2_p & v88fd1c;
assign v87feba = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd92a;
assign v883a94 = BtoS_ACK6_p & v8fd8c0 | !BtoS_ACK6_p & v8fc237;
assign v8c4d0d = RtoB_ACK1_p & v897323 | !RtoB_ACK1_p & v8fd688;
assign v88808c = jx2_p & v858320 | !jx2_p & !v8684ff;
assign v8dacfc = BtoR_REQ0_p & v885ffa | !BtoR_REQ0_p & v8fd797;
assign v882d68 = BtoR_REQ1_p & v85f322 | !BtoR_REQ1_p & v895abe;
assign v8c2ef2 = DEQ_p & v8880e4 | !DEQ_p & v8846bb;
assign v8fd4e2 = BtoS_ACK6_p & v8fd8ba | !BtoS_ACK6_p & v8fd73b;
assign v88225a = stateG7_1_p & v8fc810 | !stateG7_1_p & v844f91;
assign v88454a = jx0_p & v882186 | !jx0_p & v8fd65f;
assign v844fa3 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v8974c9 = jx0_p & v88fdb8 | !jx0_p & !v883f7a;
assign v880e0b = BtoR_REQ1_p & v879581 | !BtoR_REQ1_p & v8843d0;
assign v885ee9 = RtoB_ACK0_p & v8846ba | !RtoB_ACK0_p & v8dace1;
assign v895ccc = BtoS_ACK0_p & v8fd764 | !BtoS_ACK0_p & v8fc73e;
assign v8fc193 = RtoB_ACK1_p & v8fd852 | !RtoB_ACK1_p & v883c1a;
assign v88401d = jx0_p & v844f91 | !jx0_p & !v86ed7e;
assign v881e80 = BtoS_ACK6_p & v882bdd | !BtoS_ACK6_p & v880931;
assign v884216 = BtoS_ACK6_p & v8fd70d | !BtoS_ACK6_p & v8fd8ff;
assign v895d15 = stateG12_p & v885f4a | !stateG12_p & !v88064f;
assign v8838cd = RtoB_ACK0_p & v882d42 | !RtoB_ACK0_p & v8b5fc6;
assign v87bba1 = jx2_p & v882b41 | !jx2_p & v8843d0;
assign v882bc8 = BtoS_ACK0_p & v88493b | !BtoS_ACK0_p & v884bc5;
assign v8fd5b1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd6cc;
assign v8fc57a = jx2_p & v883cd1 | !jx2_p & v88791d;
assign v8fd20b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844fad;
assign v88086e = BtoS_ACK6_p & v885dfd | !BtoS_ACK6_p & v8fd74b;
assign v883f7a = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd7a4;
assign v888662 = jx0_p & v887bfb | !jx0_p & v844f91;
assign v882b96 = StoB_REQ2_p & v87bacb | !StoB_REQ2_p & v8fd6ae;
assign v885d65 = jx0_p & v844f9b | !jx0_p & !v8fd742;
assign v8fd2cf = ENQ_p & v884941 | !ENQ_p & v8fd8db;
assign v8fd672 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fcb34;
assign v8fd6db = BtoR_REQ0_p & v882b84 | !BtoR_REQ0_p & v8fd63d;
assign v8829ee = EMPTY_p & v8846ba | !EMPTY_p & v883c0c;
assign v8940fc = StoB_REQ3_p & v884904 | !StoB_REQ3_p & !v844f91;
assign v8fd96a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v887f3a;
assign v88402c = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v8fd57d;
assign v881faf = stateG7_1_p & v8fd8ed | !stateG7_1_p & v844f91;
assign v891e93 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v882bf5;
assign v884034 = jx1_p & v8f1f45 | !jx1_p & v8fc6fe;
assign v88945f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v880616;
assign v8fd1d0 = RtoB_ACK1_p & v883c24 | !RtoB_ACK1_p & v8810ca;
assign v884171 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v883c14;
assign v8fd837 = jx2_p & v8fd8d4 | !jx2_p & !v8877c5;
assign v8fc7cc = jx0_p & v8fd014 | !jx0_p & v8fd204;
assign v8fd5a1 = stateG12_p & v8dabf0 | !stateG12_p & v8876ed;
assign v884539 = jx0_p & v881113 | !jx0_p & !v881963;
assign v8947e0 = BtoS_ACK6_p & v885b17 | !BtoS_ACK6_p & v8876c3;
assign v884b83 = StoB_REQ6_p & v890676 | !StoB_REQ6_p & v885bf2;
assign v8fd662 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8dab99;
assign v88a5d1 = jx2_p & v897374 | !jx2_p & !v8684ff;
assign v8fc2b8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883ed8;
assign v8fd084 = jx1_p & v8818a8 | !jx1_p & !v885863;
assign v8fd7de = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v8fd87b;
assign v844fb7 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844f91;
assign v8fd863 = StoB_REQ1_p & v8fd597 | !StoB_REQ1_p & v8fd19f;
assign v8849d3 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v89471b;
assign v8fd79c = BtoR_REQ1_p & v8fd5b7 | !BtoR_REQ1_p & v880d9c;
assign v884d5e = stateG7_1_p & v88a2de | !stateG7_1_p & v882d42;
assign v8877c1 = StoB_REQ6_p & v8fd8c0 | !StoB_REQ6_p & v88089e;
assign BtoS_ACK1_n = !v8795c1;
assign v887644 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8897a6;
assign v8fc28a = jx0_p & v8841bc | !jx0_p & v884f8e;
assign v8fd457 = jx0_p & v883089 | !jx0_p & v844f91;
assign v8fd8cf = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8fd7cb;
assign v8860a7 = jx0_p & v87bb4b | !jx0_p & v888205;
assign v8b603b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v870c76;
assign v8fc945 = jx2_p & v8fd256 | !jx2_p & v88791d;
assign v883c1a = jx2_p & v876f96 | !jx2_p & v8fd641;
assign v8fcd77 = StoB_REQ3_p & v8fd7f7 | !StoB_REQ3_p & v844f91;
assign v897377 = BtoS_ACK6_p & v8fd853 | !BtoS_ACK6_p & v868e18;
assign v88579e = BtoR_REQ1_p & v885c69 | !BtoR_REQ1_p & v844f91;
assign v8c2ecf = jx2_p & v884dd2 | !jx2_p & !v8fd1ac;
assign v8fd5f2 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9d;
assign v8c0098 = jx1_p & v8856e4 | !jx1_p & !v8fd713;
assign v884afb = BtoS_ACK0_p & v88391f | !BtoS_ACK0_p & v8fd66a;
assign v898f1a = StoB_REQ1_p & v8843d1 | !StoB_REQ1_p & v894620;
assign v8dabff = jx0_p & v844f91 | !jx0_p & v8f2a3f;
assign v880eda = BtoR_REQ1_p & v89241d | !BtoR_REQ1_p & v8fccad;
assign v8fc99d = StoB_REQ0_p & v8fd856 | !StoB_REQ0_p & v8ac9d2;
assign v8fca05 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v897377;
assign v87a65f = RtoB_ACK1_p & v8fcdd0 | !RtoB_ACK1_p & v8fd94e;
assign v8fd8f3 = jx0_p & v8fd78b | !jx0_p & v883cf0;
assign v885c4b = ENQ_p & v891109 | !ENQ_p & v8dacfc;
assign v8a0a29 = BtoS_ACK6_p & v8fd853 | !BtoS_ACK6_p & v887adf;
assign v8fc35c = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8ad0bf;
assign v8dacbf = StoB_REQ6_p & v8fd775 | !StoB_REQ6_p & v844f91;
assign v8b6053 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fcc5a;
assign v884e81 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v8846a5 = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v880934;
assign v881fe6 = jx0_p & v883bb8 | !jx0_p & v8f2a3f;
assign v88810b = stateG7_1_p & v8fcae9 | !stateG7_1_p & v844f91;
assign v88097a = BtoR_REQ0_p & v8fd882 | !BtoR_REQ0_p & v854d12;
assign v8588b8 = StoB_REQ1_p & v8fd19d | !StoB_REQ1_p & v844f91;
assign v8ed1c6 = jx0_p & v844f9f | !jx0_p & !v880816;
assign v8fd740 = stateG7_1_p & v8fce87 | !stateG7_1_p & v8843d0;
assign v880934 = StoB_REQ2_p & v8fd8df | !StoB_REQ2_p & v8819ce;
assign v8805b9 = BtoR_REQ0_p & v887ccd | !BtoR_REQ0_p & v896f10;
assign v88259e = jx1_p & v8856e4 | !jx1_p & !v8fd59f;
assign v88a63c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dac30;
assign v88c103 = BtoR_REQ0_p & v88498b | !BtoR_REQ0_p & v8fd6d0;
assign v883cd1 = jx1_p & v844f91 | !jx1_p & !v887a4a;
assign v8795bb = jx1_p & v882136 | !jx1_p & !v844f91;
assign v8fc762 = RtoB_ACK0_p & v8fd812 | !RtoB_ACK0_p & v8878b5;
assign v882034 = RtoB_ACK0_p & v88367e | !RtoB_ACK0_p & v8fd2b7;
assign v85839b = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v88386a;
assign v8fd7ca = EMPTY_p & v88795b | !EMPTY_p & v8877fe;
assign v885867 = BtoS_ACK2_p & v8fd646 | !BtoS_ACK2_p & v8fd1cd;
assign v888096 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8fd865;
assign v8fd1bc = StoB_REQ0_p & v885694 | !StoB_REQ0_p & v8947e0;
assign v884fdd = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v88033b;
assign v887657 = StoB_REQ1_p & v8f2a2c | !StoB_REQ1_p & v88186f;
assign v894620 = BtoS_ACK2_p & v882d8f | !BtoS_ACK2_p & !v88496e;
assign v884d85 = ENQ_p & v887a69 | !ENQ_p & v894924;
assign v8fc3cf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v882ae0;
assign v88616c = BtoR_REQ1_p & v8fd8cd | !BtoR_REQ1_p & v88621e;
assign v881630 = StoB_REQ0_p & v8fd1e1 | !StoB_REQ0_p & v884fc8;
assign v882841 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8947b9;
assign v8b5fc6 = stateG7_1_p & v8886e1 | !stateG7_1_p & v8fd82e;
assign v883012 = StoB_REQ3_p & v8fd726 | !StoB_REQ3_p & v8910ad;
assign v882a63 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8fd658;
assign v8fd614 = jx0_p & v8fd5d2 | !jx0_p & v844f91;
assign v8ad009 = stateG7_1_p & v8fd7d5 | !stateG7_1_p & v883e92;
assign v8fd18f = jx0_p & v880816 | !jx0_p & v8972ae;
assign v87ff08 = stateG7_1_p & v8fd5d6 | !stateG7_1_p & v8fd5fd;
assign v88a4a0 = jx2_p & v87adc8 | !jx2_p & v8fd5b2;
assign v880a21 = BtoR_REQ0_p & v844fa3 | !BtoR_REQ0_p & v854113;
assign v880b8e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8fc68f;
assign v8822fe = jx1_p & v885a6c | !jx1_p & v8fc719;
assign v8fd581 = jx2_p & v8972a7 | !jx2_p & !v8684ff;
assign v8fd7c2 = stateG7_1_p & v887ad9 | !stateG7_1_p & v882db5;
assign v8fd969 = jx1_p & v883f8f | !jx1_p & v8fc2dd;
assign v89fb74 = StoB_REQ6_p & v882b15 | !StoB_REQ6_p & v8878da;
assign v8fd383 = BtoS_ACK6_p & v8a87b1 | !BtoS_ACK6_p & v88280d;
assign v88786f = StoB_REQ6_p & v8fd6b3 | !StoB_REQ6_p & v844f91;
assign v8fc679 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v880a70;
assign v8b60af = ENQ_p & v8fd5b4 | !ENQ_p & v882170;
assign v8f11a7 = jx1_p & v880ccb | !jx1_p & !v8821ba;
assign v8fd5ed = jx1_p & v8fc312 | !jx1_p & v8f2a3f;
assign v8fd236 = jx0_p & v87afd1 | !jx0_p & v8b5fc7;
assign jx0_n = v8b60d1;
assign v897cf5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v895b31;
assign v879570 = BtoS_ACK6_p & v8fd57d | !BtoS_ACK6_p & v8fd490;
assign v8881f0 = StoB_REQ1_p & v8fd597 | !StoB_REQ1_p & v8fc1bf;
assign v8fd8d5 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8fd597;
assign v880ac4 = StoB_REQ6_p & v8fc970 | !StoB_REQ6_p & v858a9b;
assign v8824d4 = jx0_p & v844f91 | !jx0_p & v86ed7e;
assign v881e33 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v88219e;
assign v88a2df = BtoR_REQ0_p & v8fd879 | !BtoR_REQ0_p & v887f47;
assign v895b2f = stateG7_1_p & v8fc6aa | !stateG7_1_p & v8fc945;
assign v8ad08b = BtoS_ACK0_p & v8fd1bd | !BtoS_ACK0_p & v884cc3;
assign v8fc802 = jx0_p & v883f65 | !jx0_p & !v844f91;
assign v887f3a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v88eb82;
assign v8fcd00 = RtoB_ACK1_p & v882490 | !RtoB_ACK1_p & v8f29e2;
assign v884834 = jx0_p & v88186b | !jx0_p & v8fd906;
assign v8fd8b2 = jx0_p & v8b78a2 | !jx0_p & v844f91;
assign v88fcc6 = EMPTY_p & v8fd7fb | !EMPTY_p & v8fd832;
assign v8fd716 = BtoS_ACK2_p & v8840c7 | !BtoS_ACK2_p & v892416;
assign v87debc = jx1_p & v885d65 | !jx1_p & !v897301;
assign v875cbc = jx2_p & v8ce1ae | !jx2_p & v88793c;
assign v8fd186 = BtoS_ACK4_p & v885b89 | !BtoS_ACK4_p & v888182;
assign v8dabe8 = jx0_p & v8fd810 | !jx0_p & v885fe4;
assign v8fd75d = jx1_p & v8f2a3f | !jx1_p & v8fcfe7;
assign v8fd72b = jx0_p & v8ce165 | !jx0_p & !v844fab;
assign v8886e1 = RtoB_ACK1_p & v894722 | !RtoB_ACK1_p & v8fd82e;
assign v884626 = BtoS_ACK6_p & v882baa | !BtoS_ACK6_p & v880236;
assign v8fd6c6 = jx1_p & v8dac82 | !jx1_p & !v8fce83;
assign v8fd8aa = jx1_p & v8fd574 | !jx1_p & v87bb66;
assign v894850 = StoB_REQ6_p & v887644 | !StoB_REQ6_p & v882a64;
assign v884984 = BtoR_REQ0_p & v8fce28 | !BtoR_REQ0_p & v8fc9fd;
assign v8fc4c0 = BtoS_ACK0_p & v88e6e1 | !BtoS_ACK0_p & v8c98e7;
assign v8ad131 = jx0_p & v8fd936 | !jx0_p & v89463b;
assign v8fd790 = BtoS_ACK1_p & v844f9e | !BtoS_ACK1_p & v8c48b7;
assign v884a91 = BtoS_ACK6_p & v885be7 | !BtoS_ACK6_p & v897405;
assign v8fd1d9 = RtoB_ACK0_p & v8881d4 | !RtoB_ACK0_p & v8830a2;
assign v88112b = RtoB_ACK0_p & v895d6d | !RtoB_ACK0_p & v884197;
assign v8fd8d0 = jx2_p & v86edd5 | !jx2_p & v87954a;
assign v8fce9e = jx0_p & v844f91 | !jx0_p & v8ce165;
assign v88397a = jx0_p & v8fc9c2 | !jx0_p & v844f91;
assign v8847be = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & !v882a93;
assign v8fd24f = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8843d1;
assign v87949d = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v887abd;
assign v885b2d = stateG7_1_p & v884907 | !stateG7_1_p & v8fc7b7;
assign v8fc8ad = stateG7_1_p & v881fdb | !stateG7_1_p & !v844f91;
assign v858acd = StoB_REQ2_p & v8fd7f7 | !StoB_REQ2_p & v859c5b;
assign v8fc6a5 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v887c2f;
assign v8878a5 = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & !v8fca9c;
assign v89fb1c = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8820d8;
assign v8844d6 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v87eaaf;
assign v880b75 = jx0_p & v8fd8d6 | !jx0_p & v8846ba;
assign v8837af = jx0_p & v884767 | !jx0_p & v885836;
assign v884a9c = jx0_p & v844f91 | !jx0_p & v8fd879;
assign v8fd6a7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fd255;
assign v881022 = jx1_p & v8821e0 | !jx1_p & v884718;
assign v8878b5 = jx2_p & v897374 | !jx2_p & !v8822bf;
assign v8fd54b = jx1_p & v887c98 | !jx1_p & v8fc6fe;
assign v8fd172 = jx0_p & v895d68 | !jx0_p & v844f91;
assign v8ed953 = jx0_p & v8fd965 | !jx0_p & v882788;
assign v88055f = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v87fb41;
assign v8fd1fd = stateG7_1_p & v8823f5 | !stateG7_1_p & v887966;
assign v8879f2 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8f2abd;
assign v88170c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v882bbf;
assign v89fb49 = StoB_REQ2_p & v887c2f | !StoB_REQ2_p & v883700;
assign v8fc3e8 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8562b0;
assign v8fc296 = jx0_p & v844f91 | !jx0_p & v8fd958;
assign v8fd1d2 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v88602f;
assign v86edd5 = jx1_p & v880ccb | !jx1_p & !v8fd5d5;
assign v8fd19b = StoB_REQ3_p & v8fc1f9 | !StoB_REQ3_p & v8ceca9;
assign v8fd914 = jx1_p & v88401d | !jx1_p & v8894e3;
assign v8fd67c = StoB_REQ1_p & v884476 | !StoB_REQ1_p & v844f9d;
assign v8fd3c8 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v882bee;
assign v8fd876 = stateG7_1_p & v8fc5c1 | !stateG7_1_p & v8fd5a2;
assign v896e20 = jx0_p & v8808eb | !jx0_p & !v8849ea;
assign v88621e = jx2_p & v8fd698 | !jx2_p & v8816be;
assign v8809c4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v887fa9;
assign v8fc64f = RtoB_ACK1_p & v8816aa | !RtoB_ACK1_p & v8fd62f;
assign v88313d = jx0_p & v894e08 | !jx0_p & v8880d8;
assign v8838a3 = BtoS_ACK1_p & v8fd7dc | !BtoS_ACK1_p & v8fd7c6;
assign v882431 = BtoS_ACK1_p & v884476 | !BtoS_ACK1_p & v898f1a;
assign v880821 = jx2_p & v8fd1ca | !jx2_p & v8fc9d9;
assign v881975 = StoB_REQ2_p & v8fd951 | !StoB_REQ2_p & v8fd872;
assign v882ea6 = jx1_p & v883f8f | !jx1_p & v89dbce;
assign v8802ff = ENQ_p & v8fd5a8 | !ENQ_p & v8fd6e0;
assign v884dd2 = jx1_p & v883d82 | !jx1_p & !v89fadb;
assign v88e5f1 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8fd696;
assign v887d9c = BtoS_ACK1_p & v88219e | !BtoS_ACK1_p & v884ac0;
assign v8822d4 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9d;
assign v882e12 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v885ab0;
assign v88442a = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v8fd96a;
assign v8876d0 = ENQ_p & v883706 | !ENQ_p & !v891da3;
assign v8fd693 = jx1_p & v8856e4 | !jx1_p & !v8fc98c;
assign v894e08 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v885cc5;
assign v883a4d = jx1_p & v884976 | !jx1_p & v88172f;
assign v879e64 = RtoB_ACK1_p & v8fd7b3 | !RtoB_ACK1_p & v8fd581;
assign v895cb4 = BtoR_REQ1_p & v8948bb | !BtoR_REQ1_p & v8fd87b;
assign v884b4e = BtoR_REQ0_p & v8fd78d | !BtoR_REQ0_p & v87948e;
assign v8fd5f7 = jx1_p & v8676b7 | !jx1_p & v883c78;
assign v884359 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v844f95;
assign v8c2df5 = RtoB_ACK1_p & v8c2ecf | !RtoB_ACK1_p & !v88386a;
assign v8fd598 = jx0_p & v895a65 | !jx0_p & v844f91;
assign v8ed1d3 = BtoS_ACK1_p & v8fd74e | !BtoS_ACK1_p & v880620;
assign v881840 = StoB_REQ1_p & v87af07 | !StoB_REQ1_p & v844f9d;
assign v882bb8 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v88e73e;
assign v883879 = BtoS_ACK1_p & v882bdd | !BtoS_ACK1_p & v8fd4c4;
assign v8831e6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v854c1c;
assign v8fd841 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8588ba;
assign v887d78 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v887ad8;
assign v8fca9c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8fd775;
assign v8fd88a = BtoS_ACK3_p & v88576e | !BtoS_ACK3_p & v880c71;
assign v883928 = stateG7_1_p & v8587ee | !stateG7_1_p & v8fd752;
assign v885bee = BtoS_ACK0_p & v8fd7dc | !BtoS_ACK0_p & v885748;
assign v8fd281 = jx1_p & v880750 | !jx1_p & !v8fd82b;
assign v8fc7b1 = jx2_p & v8fd5ea | !jx2_p & v8c2de5;
assign v8fd8ba = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8fd73a;
assign v8fcd75 = StoB_REQ0_p & v888096 | !StoB_REQ0_p & v8802a2;
assign v887c9a = jx0_p & v8569e0 | !jx0_p & v8fc9d9;
assign v8fd579 = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v858422;
assign v884565 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v884ac0;
assign v8fd797 = BtoR_REQ1_p & v8fd8b9 | !BtoR_REQ1_p & v844f91;
assign v8dac82 = jx0_p & v885fe8 | !jx0_p & v86a020;
assign v882fd1 = stateG7_1_p & v8fd75b | !stateG7_1_p & v8810ca;
assign v8fd688 = jx2_p & v88023c | !jx2_p & v8fc2e5;
assign v887680 = EMPTY_p & v8fd95a | !EMPTY_p & !v8d6a33;
assign v8fccca = jx0_p & v885fe3 | !jx0_p & v8fceeb;
assign v8fd254 = BtoS_ACK6_p & v8fd764 | !BtoS_ACK6_p & v8fd849;
assign v8fd5ab = StoB_REQ6_p & v8fd819 | !StoB_REQ6_p & v844f91;
assign v8fd64d = BtoS_ACK3_p & v8fca41 | !BtoS_ACK3_p & v88079c;
assign v8805c4 = jx0_p & v844f9f | !jx0_p & !v844f91;
assign v8fd65a = stateG7_1_p & v8fd8bc | !stateG7_1_p & v884f1f;
assign v8ad079 = BtoS_ACK1_p & v88219e | !BtoS_ACK1_p & v8fd637;
assign v884f8e = BtoS_ACK0_p & v8d4e0d | !BtoS_ACK0_p & v88237c;
assign v8fd230 = stateG7_1_p & v88963d | !stateG7_1_p & v8878b5;
assign v8fd652 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v885f26;
assign v8fd78e = StoB_REQ1_p & v8ad0e2 | !StoB_REQ1_p & !v844f91;
assign v844fbf = stateG7_1_p & v844f91 | !stateG7_1_p & !v844f91;
assign v8793ad = stateG7_1_p & v858985 | !stateG7_1_p & v882a0a;
assign v8fd856 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8fd24f;
assign v8fd6d0 = RtoB_ACK0_p & v88367e | !RtoB_ACK0_p & v885ab1;
assign v88118b = StoB_REQ6_p & v8878ac | !StoB_REQ6_p & v8829b5;
assign v887ab9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fd864;
assign v8837ba = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f9b;
assign v88251e = BtoS_ACK0_p & v8fd746 | !BtoS_ACK0_p & v88363c;
assign v885cc5 = StoB_REQ0_p & v8fc295 | !StoB_REQ0_p & v844f91;
assign v885077 = jx0_p & v8fd8c7 | !jx0_p & v8fd85f;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v8fd1a0 = BtoS_ACK2_p & v882214 | !BtoS_ACK2_p & v8fd002;
assign v8861df = BtoR_REQ1_p & v884b64 | !BtoR_REQ1_p & v8f29e2;
assign v8fd23a = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v880263;
assign v88fbd1 = jx0_p & v844f91 | !jx0_p & v8fd5cc;
assign v8fc61c = StoB_REQ6_p & v8fd8d5 | !StoB_REQ6_p & v8fd773;
assign v884482 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8fd455;
assign v8810bc = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v887de8;
assign v8dad14 = BtoS_ACK6_p & v884ac0 | !BtoS_ACK6_p & v890631;
assign v8fd59f = jx0_p & v8fd5d2 | !jx0_p & !v8947ee;
assign v8fd8eb = BtoS_ACK0_p & v884919 | !BtoS_ACK0_p & v8a87bc;
assign v88023c = jx1_p & v844f91 | !jx1_p & !v8816cc;
assign v8fd5d5 = jx0_p & v88fa9a | !jx0_p & v887b09;
assign v88e43b = StoB_REQ2_p & v8fd7f7 | !StoB_REQ2_p & v887de8;
assign v876f96 = jx1_p & v8fd035 | !jx1_p & v882ac1;
assign v89736f = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v88079c;
assign v8fd8e2 = jx0_p & v8fd782 | !jx0_p & v8fc77f;
assign v8805be = BtoS_ACK1_p & v8fd70d | !BtoS_ACK1_p & v8fd5d3;
assign v8846d2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fc35c;
assign v8c48b3 = BtoS_ACK6_p & v885dfd | !BtoS_ACK6_p & v887a24;
assign v87ff04 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v8fcdd5 = stateG7_1_p & v885d73 | !stateG7_1_p & v887aed;
assign v882002 = ENQ_p & v8fd8ea | !ENQ_p & v892ca3;
assign v882ae0 = StoB_REQ0_p & v8fc2d4 | !StoB_REQ0_p & v8fd642;
assign v880660 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & !v844f91;
assign v87945a = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8fc61c;
assign v891077 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v88786f;
assign v884b2b = stateG7_1_p & v887924 | !stateG7_1_p & v8fd5cd;
assign v897301 = jx0_p & v8fd742 | !jx0_p & v844f91;
assign v887966 = jx2_p & v8fd666 | !jx2_p & v87bb66;
assign v8ad0bf = StoB_REQ6_p & v88254c | !StoB_REQ6_p & v8fd813;
assign v8fcf21 = StoB_REQ0_p & v8847be | !StoB_REQ0_p & v844f91;
assign v8fd724 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8fd1c9;
assign v8fd572 = StoB_REQ2_p & v8fd7a1 | !StoB_REQ2_p & v8fd92f;
assign v883a3f = jx0_p & v8a0b36 | !jx0_p & v8fcff6;
assign v8ed93d = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8fd856;
assign v8fd669 = jx0_p & v8ad08b | !jx0_p & !v8ed93d;
assign v8fd592 = jx0_p & v854d5c | !jx0_p & v882066;
assign v8fd832 = stateG12_p & v880fa6 | !stateG12_p & v885733;
assign SLC0_n = (DEQ_n & ((FULL_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!FULL_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))))) | (!DEQ_n & ((EMPTY_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!BtoR_REQ1_n & ((!BtoS_ACK0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC1_n))) | (!jx2_n & ((jx1_n & ((SLC1_n))) | (!jx1_n & ((!jx0_n & ((SLC1_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC1_n))) | (!jx2_n & ((jx1_n & ((SLC1_n))) | (!jx1_n & ((!jx0_n & ((SLC1_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC1_n))) | (!jx2_n & ((jx1_n & ((SLC1_n))) | (!jx1_n & ((!jx0_n & ((SLC1_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC1_n))) | (!jx2_n & ((jx1_n & ((SLC1_n))) | (!jx1_n & ((!jx0_n & ((SLC1_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((!BtoS_ACK0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!RtoB_ACK1_n & ((!BtoS_ACK0_n & ((!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC1_n))) | (!jx2_n & ((jx1_n & ((SLC1_n))) | (!jx1_n & ((!jx0_n & ((SLC1_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((stateG12_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n))) | (!jx0_n & ((!StoB_REQ6_n & ((SLC1_n))))))) | (!jx1_n & ((!StoB_REQ6_n & ((SLC1_n))))))) | (!jx2_n & ((!StoB_REQ6_n & ((SLC1_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n))) | (!jx0_n & ((!StoB_REQ6_n & ((SLC1_n))))))) | (!jx1_n & ((!StoB_REQ6_n & ((SLC1_n))))))) | (!jx2_n & ((!StoB_REQ6_n & ((SLC1_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!stateG12_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((!StoB_REQ6_n & ((SLC1_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n))))) | (!StoB_REQ2_n & ((SLC1_n))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n & ((SLC1_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n)))))))))))))))))))))))))))))))))))))));
assign ENQ_n = (DEQ_n & ((stateG12_n & ((BtoR_REQ0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((!jx0_n & ((StoB_REQ6_n))))) | (!jx1_n & ((StoB_REQ6_n))))) | (!jx2_n & ((StoB_REQ6_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n) | (!stateG7_1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))) | (!SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n) | (!RtoB_ACK1_n & ((jx2_n) | (!jx2_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))) | (!SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))))))))))))) | (!EMPTY_n & ((!FULL_n & ((stateG12_n & ((BtoR_REQ0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((!jx0_n & ((StoB_REQ6_n))))) | (!jx1_n & ((StoB_REQ6_n))))) | (!jx2_n & ((StoB_REQ6_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((!jx0_n & ((StoB_REQ6_n))))) | (!jx1_n & ((StoB_REQ6_n))))) | (!jx2_n & ((StoB_REQ6_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))))))))))))))) | (!stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((SLC2_n & ((!SLC1_n))) | (!SLC2_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC2_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((SLC2_n)))))))))))))))))))))));
assign SLC2_n = (DEQ_n & ((FULL_n & ((stateG12_n & ((BtoR_REQ0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC0_n))) | (!jx0_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx1_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx2_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC0_n))) | (!jx0_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx1_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx2_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!stateG12_n & ((SLC0_n))))) | (!FULL_n & ((stateG12_n & ((BtoR_REQ0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC0_n))) | (!jx0_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx1_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx2_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!stateG12_n & ((SLC0_n))))))) | (!DEQ_n & ((EMPTY_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((!BtoS_ACK0_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))) | (!jx0_n & ((StoB_REQ6_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((!BtoS_ACK0_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))) | (!jx0_n & ((StoB_REQ6_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC0_n))) | (!jx2_n & ((jx1_n & ((SLC0_n))) | (!jx1_n & ((!jx0_n & ((SLC0_n))))))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC0_n))) | (!jx2_n & ((jx1_n & ((SLC0_n))) | (!jx1_n & ((!jx0_n & ((SLC0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC0_n))) | (!jx2_n & ((jx1_n & ((SLC0_n))) | (!jx1_n & ((!jx0_n & ((SLC0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC0_n))) | (!jx2_n & ((jx1_n & ((SLC0_n))) | (!jx1_n & ((!jx0_n & ((SLC0_n))))))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!RtoB_ACK1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((!BtoS_ACK0_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))) | (!jx0_n & ((StoB_REQ6_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))))) | (!RtoB_ACK1_n & ((!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n) | (!jx2_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))) | (!jx0_n & ((StoB_REQ6_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx2_n & ((SLC0_n))) | (!jx2_n & ((jx1_n & ((SLC0_n))) | (!jx1_n & ((!jx0_n & ((SLC0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((SLC0_n))) | (!FULL_n & ((stateG12_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC0_n))) | (!jx0_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx1_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx2_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC0_n))) | (!jx0_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx1_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!jx2_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!stateG12_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!jx2_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC0_n))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((SLC0_n))))) | (!BtoS_ACK6_n & ((jx2_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx0_n & ((StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC0_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n)))))))))))))))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  StoB_REQ4_p = 0;
  StoB_REQ5_p = 0;
  StoB_REQ6_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoS_ACK4_p = 0;
  BtoS_ACK5_p = 0;
  BtoS_ACK6_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  SLC2_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  StoB_REQ4_p = StoB_REQ4_n;
  StoB_REQ5_p = StoB_REQ5_n;
  StoB_REQ6_p = StoB_REQ6_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoS_ACK4_p = BtoS_ACK4_n;
  BtoS_ACK5_p = BtoS_ACK5_n;
  BtoS_ACK6_p = BtoS_ACK6_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  SLC2_p = SLC2_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
