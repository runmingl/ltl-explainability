module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hbusreq2, hlock2, hbusreq3, hlock3, hbusreq4, hlock4, hburst0, hburst1, hmaster0, hmaster1, hmaster2, hmastlock, start, decide, locked, hgrant0, hgrant1, hgrant2, hgrant3, hgrant4, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, stateG10_2, stateG10_3, stateG10_4, jx0, jx1, jx2);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v845542;
  wire v845578;
  wire v84555e;
  wire v889629;
  wire c3d667;
  wire c3d668;
  wire c3d669;
  wire c3d66a;
  wire c3d66b;
  wire c3d66c;
  wire v84557a;
  wire c3d66d;
  wire c3d66e;
  wire c3d66f;
  wire c3d670;
  wire c3d671;
  wire c3d672;
  wire c3d673;
  wire c3d674;
  wire c3d675;
  wire c3d676;
  wire c3d677;
  wire c3d678;
  wire c3d679;
  wire c3d67a;
  wire c3d67b;
  wire c3d67c;
  wire c3d67d;
  wire c3d67e;
  wire c3d67f;
  wire c3d680;
  wire c3d681;
  wire c3d682;
  wire c3d683;
  wire c3d684;
  wire c3d685;
  wire c3d686;
  wire c3d687;
  wire c3d688;
  wire c3d689;
  wire c3d68a;
  wire c3d68b;
  wire c3d68c;
  wire c3d68d;
  wire c3d68e;
  wire c3d68f;
  wire c3d690;
  wire c3d691;
  wire c3d692;
  wire c3d693;
  wire c3d694;
  wire c3d695;
  wire c3d696;
  wire c3d697;
  wire c3d698;
  wire c3d699;
  wire c3d69a;
  wire c3d69b;
  wire c3d69c;
  wire c3d69d;
  wire c3d69e;
  wire c3d69f;
  wire c3d6a0;
  wire c3d6a1;
  wire c3d6a2;
  wire c3d6a3;
  wire c3d6a4;
  wire c3d6a5;
  wire c3d6a6;
  wire c3d6a7;
  wire c3d6a8;
  wire c3d6a9;
  wire c3d6aa;
  wire c3d6ab;
  wire c3d6ac;
  wire c3d6ad;
  wire c3d6ae;
  wire c3d6af;
  wire c3d6b0;
  wire c3d6b1;
  wire c3d6b2;
  wire c3d6b3;
  wire c3d6b4;
  wire c3d6b5;
  wire c3d6b6;
  wire c3d6b7;
  wire c3d6b8;
  wire c3d6b9;
  wire c3d6ba;
  wire c3d6bb;
  wire c3d6bc;
  wire c3d6bd;
  wire c3d6be;
  wire c3d6bf;
  wire c3d6c0;
  wire c3d6c1;
  wire c3d6c2;
  wire c3d6c3;
  wire c3d6c4;
  wire c3d6c5;
  wire c3d6c6;
  wire c3d6c7;
  wire c3d6c8;
  wire c3d6c9;
  wire c3d6ca;
  wire c3d6cb;
  wire c3d6cc;
  wire c3d6cd;
  wire c3d6ce;
  wire c3d6cf;
  wire c3d6d0;
  wire c3d6d1;
  wire c3d6d2;
  wire c3d6d3;
  wire c3d6d4;
  wire c3d6d5;
  wire c3d6d6;
  wire c3d6d7;
  wire c3d6d8;
  wire c3d6d9;
  wire c3d6da;
  wire c3d6db;
  wire c3d6dc;
  wire c3d6dd;
  wire c3d6de;
  wire c3d6df;
  wire c3d6e0;
  wire c3d6e1;
  wire c3d6e2;
  wire c3d6e3;
  wire c3d6e4;
  wire c3d6e5;
  wire c3d6e6;
  wire c3d6e7;
  wire c3d6e8;
  wire c3d6e9;
  wire c3d6ea;
  wire c3d6eb;
  wire c3d6ec;
  wire c3d6ed;
  wire c3d6ee;
  wire c3d6ef;
  wire c3d6f0;
  wire c3d6f1;
  wire c3d6f2;
  wire c3d6f3;
  wire c3d6f4;
  wire c3d6f5;
  wire c3d6f6;
  wire c3d6f7;
  wire c3d6f8;
  wire c3d6f9;
  wire c3d6fa;
  wire c3d6fb;
  wire c3d6fc;
  wire c3d6fd;
  wire c3d6fe;
  wire c3d6ff;
  wire c3d700;
  wire c3d701;
  wire c3d702;
  wire c3d703;
  wire c3d704;
  wire c3d705;
  wire c3d706;
  wire c3d707;
  wire c3d708;
  wire c3d709;
  wire c3d70a;
  wire c3d70b;
  wire c3d70c;
  wire c3d70d;
  wire c3d70e;
  wire c3d70f;
  wire c3d710;
  wire c3d711;
  wire c3d712;
  wire c3d713;
  wire c3d714;
  wire c3d715;
  wire c3d716;
  wire c3d717;
  wire c3d718;
  wire c3d719;
  wire c3d71a;
  wire c3d71b;
  wire c3d71c;
  wire c3d71d;
  wire c3d71e;
  wire c3d71f;
  wire c3d720;
  wire c3d721;
  wire c3d722;
  wire c3d723;
  wire c3d724;
  wire c3d725;
  wire c3d726;
  wire c3d727;
  wire c3d728;
  wire c3d729;
  wire c3d72a;
  wire c3d72b;
  wire c3d72c;
  wire c3d72d;
  wire c3d72e;
  wire c3d72f;
  wire c3d730;
  wire c3d731;
  wire c3d732;
  wire c3d733;
  wire c3d734;
  wire c3d735;
  wire c3d736;
  wire c3d737;
  wire c3d738;
  wire c3d739;
  wire c3d73a;
  wire c3d73b;
  wire c3d73c;
  wire c3d73d;
  wire c3d73e;
  wire c3d73f;
  wire c3d740;
  wire c3d741;
  wire c3d742;
  wire c3d743;
  wire c3d744;
  wire c3d745;
  wire c3d746;
  wire c3d747;
  wire c3d748;
  wire c3d749;
  wire c3d74a;
  wire c3d74b;
  wire c3d74c;
  wire c3d74d;
  wire c3d74e;
  wire c3d74f;
  wire c3d750;
  wire c3d751;
  wire c3d752;
  wire c3d753;
  wire c3d754;
  wire c3d755;
  wire c3d756;
  wire c3d757;
  wire c3d758;
  wire c3d759;
  wire c3d75a;
  wire c3d75b;
  wire c3d75c;
  wire c3d75d;
  wire c3d75e;
  wire c3d75f;
  wire c3d760;
  wire c3d761;
  wire c3d762;
  wire c3d763;
  wire v84554c;
  wire ad13df;
  wire ad13e0;
  wire ad13e1;
  wire ad13e2;
  wire ad13e3;
  wire ad13e4;
  wire ad13e5;
  wire v845550;
  wire v845572;
  wire ba05cd;
  wire ba05ce;
  wire ba05cf;
  wire ba05d0;
  wire v845558;
  wire v9041a4;
  wire v898970;
  wire v85746e;
  wire aa425c;
  wire aa425d;
  wire v845564;
  wire v8587b7;
  wire v86cea1;
  wire v857463;
  wire aa425e;
  wire aa425f;
  wire aa4260;
  wire v845580;
  wire bbbcd6;
  wire bb9c5a;
  wire bbbcd8;
  wire v8ccb66;
  wire v8ccb67;
  wire v8ccb68;
  wire v8ccb69;
  wire v8ccb6a;
  wire v8ccb6b;
  wire v8ccb6d;
  wire v8ccb6e;
  wire v8ccb72;
  wire v8ccb74;
  wire v8d29f8;
  wire v8d29f9;
  wire v8d29fa;
  wire v8ccb75;
  wire v8ccb76;
  wire v8ccb78;
  wire v8ccb79;
  wire v8ccb7b;
  wire v8ccb7e;
  wire v8ccb80;
  wire v8ccb81;
  wire v8ccb82;
  wire v8ccb83;
  wire v8ccb84;
  wire v8ccb87;
  wire v8ccb88;
  wire v8ccb89;
  wire v8ccb8c;
  wire v8ccb8d;
  wire v8ccb8f;
  wire v8ccbd6;
  wire v8ccbd7;
  wire v8d2b2b;
  wire v8ccbd8;
  wire v8ccbd9;
  wire v8ccbda;
  wire v8ccbdb;
  wire v8ccbdc;
  wire v8ccbdd;
  wire v8ccbde;
  wire v8ccbe1;
  wire v8ccbe2;
  wire v8ccbe3;
  wire v8ccbe5;
  wire v8ccbe6;
  wire v8ccbe7;
  wire v8ccbe8;
  wire v8ccbeb;
  wire v8ccbec;
  wire v8ccbee;
  wire v8ccbf0;
  wire v8ccbf2;
  wire v8ccbf3;
  wire v8ccbf4;
  wire v8ccbf6;
  wire v8ccbf7;
  wire v8ccbf8;
  wire v8ccbf9;
  wire v8ccbfa;
  wire v8ccbfb;
  wire v8cc434;
  wire v8cc435;
  wire v8cc436;
  wire v8cc437;
  wire v8cc438;
  wire v8cc439;
  wire v8cc43a;
  wire v8cc43b;
  wire v8cc43d;
  wire v8cc43f;
  wire v8cc455;
  wire v8cc470;
  wire v8cc472;
  wire v8d2b2e;
  wire v8cc473;
  wire v8cc474;
  wire v8cc475;
  wire v8cc476;
  wire v8cc479;
  wire v8cc47a;
  wire v8cc47b;
  wire v8cc47c;
  wire v8cc47d;
  wire v8cc47f;
  wire v8cc481;
  wire v8cc482;
  wire v8cc483;
  wire v8cc484;
  wire v8cc487;
  wire v8cc488;
  wire v8cc489;
  wire v8cc48a;
  wire v8cc48c;
  wire v8cc48d;
  wire v8cc48e;
  wire v8cc48f;
  wire v8cc491;
  wire v8cc492;
  wire v8cc493;
  wire v8cc494;
  wire v8cc496;
  wire v8cc497;
  wire v8cc498;
  wire v8cc499;
  wire v8cc49a;
  wire v8cc49c;
  wire v8cc49d;
  wire v8cc49e;
  wire v8cc49f;
  wire v8cc4a0;
  wire v8cc4a1;
  wire v8cc4a2;
  wire v8cc4a3;
  wire v8cc4a4;
  wire v8cc4a5;
  wire v8cc4a6;
  wire v8cc4a7;
  wire v8cc4a8;
  wire v8cc4a9;
  wire v8cc4aa;
  wire v8cc4ab;
  wire v8cc4ac;
  wire v8cc4ad;
  wire v8cc4ae;
  wire v8cc4af;
  wire v8cc4b0;
  wire v8cc4b1;
  wire v8cc4b2;
  wire v8cc4b3;
  wire v8cc4b4;
  wire v8cc4b6;
  wire v8cc4b8;
  wire v8cc4b9;
  wire v8cc4ba;
  wire v8cc4bb;
  wire v8cc4da;
  wire v8cc4db;
  wire v8cc4dc;
  wire v8cc4dd;
  wire v8cc4df;
  wire v8cc4e0;
  wire v8d29fb;
  wire v8cc4ed;
  wire v8cc4ee;
  wire v8cc4f0;
  wire v8cc4f1;
  wire v8cc4f2;
  wire v8cc4f3;
  wire v8cc4f4;
  wire v8cc4f6;
  wire v8cc4f7;
  wire v8cc4f9;
  wire v8cc4fa;
  wire v8cc4fc;
  wire v8cc4fd;
  wire v8cc4fe;
  wire v8cc500;
  wire v8cc501;
  wire v8cc502;
  wire v8cc503;
  wire v8cc504;
  wire v8cc506;
  wire v8cc507;
  wire v8cc508;
  wire v8cc509;
  wire v8cc50a;
  wire v8cc50c;
  wire v8cc50d;
  wire v8cc50e;
  wire v8cc50f;
  wire v8cc58f;
  wire v8cc590;
  wire v8cc592;
  wire v8cc593;
  wire v8cc595;
  wire v8cc598;
  wire v8cc599;
  wire v8cc59b;
  wire v8cc59c;
  wire v8cc59e;
  wire v8cc59f;
  wire v8cc5a0;
  wire v8cc5a4;
  wire v8cc5a5;
  wire v8cc5a6;
  wire v8cc5a7;
  wire v8cc5a8;
  wire v8cc5a9;
  wire v8cc5aa;
  wire v8cc5ab;
  wire v8cc5ac;
  wire v8cc5b0;
  wire v8cc5b1;
  wire v8cc5b2;
  wire v8cc5b3;
  wire v8cc5b4;
  wire v8cc5b5;
  wire v8cc5b9;
  wire v8cc5ba;
  wire v8cc5bb;
  wire v8cc5bd;
  wire v8cc5be;
  wire v8cc5bf;
  wire v8cc5c0;
  wire v8cc5c1;
  wire v8cc5c2;
  wire v8cc5c4;
  wire v8cc5c5;
  wire v8cc5c6;
  wire v8cc5c7;
  wire v8cc5c8;
  wire v8cc5c9;
  wire v8cc5f8;
  wire v8cc5f9;
  wire v8cc5fb;
  wire v8cc5fd;
  wire v8cc5fe;
  wire v8cc5ff;
  wire v8cc600;
  wire v8cc601;
  wire v8cc602;
  wire v8cc603;
  wire v8cc604;
  wire v8cc619;
  wire v8cc61a;
  wire v8cc61c;
  wire v8cc61e;
  wire v8cc620;
  wire v8cc621;
  wire v8cc623;
  wire v8cc624;
  wire v8cc625;
  wire v8cc626;
  wire v8cc627;
  wire v8cc628;
  wire v8cc629;
  wire v8cc62b;
  wire v8cc62c;
  wire v8cc62d;
  wire v8cc62e;
  wire v8cc62f;
  wire v8cc630;
  wire v8cc633;
  wire v8cc634;
  wire v8cc6b3;
  wire v8cc6b4;
  wire v8cc6b5;
  wire v8cc6b6;
  wire v8cc6b7;
  wire v8cc6b8;
  wire v8cc757;
  wire v8cc758;
  wire v8cc759;
  wire v8cc75b;
  wire v8cc75c;
  wire v8cc75e;
  wire v8cc75f;
  wire v8cc760;
  wire v8cc761;
  wire v8cc762;
  wire v8cc763;
  wire v8cc765;
  wire v8cc766;
  wire v8cc768;
  wire v8cc769;
  wire v8cc76b;
  wire v8cc76c;
  wire v8cc76e;
  wire v8cc781;
  wire v8cc782;
  wire v8cc783;
  wire v8cc784;
  wire v8cc785;
  wire v8cc786;
  wire v8cc787;
  wire v8cc788;
  wire v8cc789;
  wire v8cc78a;
  wire v8cc78b;
  wire v8cc78d;
  wire v8cc78e;
  wire v8cc78f;
  wire v8cc790;
  wire v8cc791;
  wire v8cc792;
  wire v8cc793;
  wire v8cc796;
  wire v8cc797;
  wire v8cc798;
  wire v8cc799;
  wire v8cc79a;
  wire v8cc79b;
  wire v8cc79c;
  wire v8cc79d;
  wire v8cc79e;
  wire v8cc79f;
  wire v8cc7a0;
  wire v8cc7a1;
  wire v8cc7a2;
  wire v8cc7a5;
  wire v8cc7a6;
  wire v8cc7a7;
  wire v8cc7a8;
  wire v8cc7aa;
  wire v8cc7ab;
  wire v8cc7ad;
  wire v8cc7b0;
  wire v8cc7b1;
  wire v8cc7b2;
  wire v8cc7b4;
  wire v8cc7b5;
  wire v8cc7b6;
  wire v8cc7b8;
  wire v8cc7b9;
  wire v8cc7ba;
  wire v8cc7bb;
  wire v8cc7bc;
  wire v8cc7bd;
  wire v8cc7bf;
  wire v8cc7c0;
  wire v8cc7c1;
  wire v8cc7c2;
  wire v8cc7c3;
  wire v8cc7c4;
  wire v8cc7c5;
  wire v8cc7c8;
  wire v8cc7c9;
  wire v8cc7ca;
  wire v8cc7cb;
  wire v8cc7cc;
  wire v8cc7cd;
  wire v8cc7ce;
  wire v8cc7cf;
  wire v8cc7d0;
  wire v8cc7d2;
  wire v8cc7d3;
  wire v8cc7d5;
  wire v8cc7d7;
  wire v8cc7d8;
  wire v8cc7d9;
  wire v8cc7da;
  wire v8cc7db;
  wire v8cc7dc;
  wire v8cc7dd;
  wire v8cc7de;
  wire v8cc7df;
  wire v8cc7e1;
  wire v8cc7e2;
  wire v8cc7e3;
  wire v8cc7e4;
  wire v8cc7e5;
  wire v8cc7e6;
  wire v8cc7e7;
  wire v8cc7e8;
  wire v8cc7e9;
  wire v8cc7ea;
  wire v8cc7eb;
  wire v8cc7ee;
  wire v8cc7ef;
  wire v8cc7f0;
  wire v8cc7f1;
  wire v8cc7f4;
  wire v8cc7f7;
  wire v8cc7f8;
  wire v8cc7f9;
  wire v8cc7fa;
  wire v8cc7fc;
  wire v8cc7fd;
  wire v8cc7fe;
  wire v8cc7ff;
  wire v8cc800;
  wire v8cc801;
  wire v8cc802;
  wire v8cc803;
  wire v8cc805;
  wire v8cc806;
  wire v8cc807;
  wire v8cc808;
  wire v8cc809;
  wire v8cc80a;
  wire v8cc80b;
  wire v8cc80c;
  wire v8cc80d;
  wire v8cc80f;
  wire v8cc810;
  wire v8cc812;
  wire v8cc813;
  wire v8cc815;
  wire v8cc816;
  wire v8cc818;
  wire v8cc819;
  wire v8cc81a;
  wire v8cc81c;
  wire v8cc81d;
  wire v8cc81e;
  wire v8cc81f;
  wire v8cc820;
  wire v8cc821;
  wire v8cc822;
  wire v8cc825;
  wire v8cc826;
  wire v8cc827;
  wire v8cc829;
  wire v8cc82a;
  wire v8cc82c;
  wire v8cc82e;
  wire v8cc031;
  wire v8cc034;
  wire v8cc035;
  wire v8cc036;
  wire v8cc038;
  wire v8cc0c2;
  wire v8cc0c3;
  wire v8cc0c4;
  wire v8cc0c5;
  wire v8cc0c9;
  wire v8cc0ca;
  wire v8cc0ce;
  wire v8cc0cf;
  wire v8cc0d0;
  wire v8cc0d1;
  wire v8cc0d2;
  wire v8cc0d3;
  wire v8cc0d4;
  wire v8cc0d5;
  wire v8cc0d6;
  wire v8cc0d7;
  wire v8cc0d8;
  wire v8cc0d9;
  wire v8cc0da;
  wire v8cc0db;
  wire v8cc0dc;
  wire v8cc0dd;
  wire v8cc0de;
  wire v8cc0df;
  wire v8cc0e0;
  wire v8cc0e1;
  wire v8cc0e2;
  wire v8cc0e4;
  wire v8cc0e6;
  wire v8cc0e7;
  wire v8cc0e8;
  wire v8cc0e9;
  wire v8cc0eb;
  wire v8cc0ec;
  wire v8cc0ee;
  wire v8cc0f0;
  wire v8cc0f1;
  wire v8cc0f2;
  wire v8cc0f4;
  wire v8cc0f5;
  wire v8cc11e;
  wire v8cc11f;
  wire v8cc120;
  wire v8cc121;
  wire v8cc122;
  wire v8cc125;
  wire v8cc126;
  wire v8cc127;
  wire v8cc128;
  wire v8cc129;
  wire v8cc12a;
  wire v8cc12b;
  wire v8cc12d;
  wire v8cc12f;
  wire v8cc130;
  wire v8cc132;
  wire v8cc167;
  wire v8cc169;
  wire v8cc16a;
  wire v8cc16c;
  wire v8cc16f;
  wire v8cc170;
  wire v845560;
  wire d6ebc9;
  wire v845570;
  wire d6ebca;
  wire d6ebcb;
  wire d6ebcc;
  wire v845568;
  wire bb9bdc;
  wire bb9bdd;
  wire c5c88b;
  wire c5c88c;
  wire c5c88d;
  wire c5c88e;
  wire c5c88f;
  wire c5c890;
  wire c5c891;
  wire c5c892;
  wire c5c893;
  wire c5c894;
  wire c5c895;
  wire c5c896;
  wire c5c897;
  wire c5c898;
  wire c5c899;
  wire c5c89a;
  wire c5c89b;
  wire c5c89c;
  wire c5c89d;
  wire c5c89e;
  wire c5c89f;
  wire c5c8a0;
  wire c5c8a1;
  wire c5c8a2;
  wire c5c8a3;
  wire c5c8a4;
  wire c5c8a5;
  wire c5c8a6;
  wire c5c8a7;
  wire c5c8a8;
  wire c5c8e0;
  wire c5c8e1;
  wire c5c8e2;
  wire c5c8e3;
  wire c5c8e4;
  wire c5c8e5;
  wire c5c8e6;
  wire c5c8e7;
  wire c5c8e8;
  wire c5c8e9;
  wire c5c8ea;
  wire c5c8eb;
  wire c5c8ec;
  wire c5c8ed;
  wire c5c8ee;
  wire c5c8ef;
  wire c5c8f0;
  wire c5c8f1;
  wire c5c8f2;
  wire c5c8f3;
  wire c5c8f4;
  wire c5c8f5;
  wire c5c8f6;
  wire c5c8f7;
  wire c5c8f8;
  wire c5c8f9;
  wire c5c8fa;
  wire c5c8fb;
  wire c5c8fc;
  wire c5c8fd;
  wire c5c8fe;
  wire c5c8ff;
  wire c5c900;
  wire c5c901;
  wire c5c902;
  wire c5c903;
  wire c5c904;
  wire c5c905;
  wire c5c92c;
  wire c5c92d;
  wire c5c92e;
  wire c5c92f;
  wire c5c930;
  wire c5c931;
  wire c5c932;
  wire c5c933;
  wire c5c934;
  wire c5c935;
  wire c5c936;
  wire c5c937;
  wire c5c938;
  wire c5c939;
  wire c5c93a;
  wire c5c93b;
  wire c5c93c;
  wire c5c93d;
  wire c5c93e;
  wire c5c93f;
  wire c5c940;
  wire c5c951;
  wire c5c952;
  wire c5c953;
  wire c5c966;
  wire c5c967;
  wire c5c968;
  wire c5c969;
  wire c5c96a;
  wire c5c96b;
  wire c5c96c;
  wire c5c96d;
  wire c5c96e;
  wire c5c96f;
  wire c5c970;
  wire c5c971;
  wire c5c972;
  wire c5c973;
  wire c5c974;
  wire c5c975;
  wire c5c976;
  wire c5c977;
  wire c5c978;
  wire c5c979;
  wire c5c97a;
  wire c5c97b;
  wire c5c97c;
  wire c5c999;
  wire c5c99a;
  wire c5c99b;
  wire c5c99c;
  wire c5c99d;
  wire c5c99e;
  wire c5c99f;
  wire c5c9a0;
  wire c5c9a8;
  wire c5c9a9;
  wire c5c9aa;
  wire c5c9ab;
  wire c5c9ac;
  wire c5c9ad;
  wire c5c9ae;
  wire c5c9af;
  wire c5c9b0;
  wire c5c9b1;
  wire c5c9b2;
  wire c5c9b3;
  wire c5c9b4;
  wire c5c9b5;
  wire c5c9b6;
  wire c5c3b5;
  wire c5c3b6;
  wire c5c3b7;
  wire c5c3be;
  wire c5c3bf;
  wire c5bed6;
  wire v857b36;
  wire c74a04;
  wire v8f2540;
  wire adea85;
  wire adea86;
  wire adea87;
  wire adea88;
  wire adea89;
  wire adea8a;
  wire adea8b;
  wire adea8c;
  wire adea8d;
  wire adea8f;
  wire adea90;
  wire v84556c;
  wire adea92;
  wire adea93;
  wire adea94;
  wire adea95;
  wire adea96;
  wire adea97;
  wire adea98;
  wire adea99;
  wire adea9a;
  wire adea9b;
  wire adea9c;
  wire adea9d;
  wire adea9e;
  wire adea9f;
  wire adeaa0;
  wire adeaa1;
  wire adeaa2;
  wire v845576;
  wire adeaa4;
  wire adeaa5;
  wire adeaa6;
  wire adeaa7;
  wire adeaa8;
  wire adeaab;
  wire adeaac;
  wire adeaad;
  wire v845566;
  wire adeaae;
  wire adeaaf;
  wire adeab0;
  wire adeab1;
  wire adeab2;
  wire adeab3;
  wire adeab4;
  wire adeab5;
  wire adeab6;
  wire adeab7;
  wire adeab8;
  wire adeab9;
  wire adec89;
  wire adec8a;
  wire bbbcd9;
  wire adec8b;
  wire adec8c;
  wire adec8d;
  wire adec8e;
  wire adec8f;
  wire adec90;
  wire adec91;
  wire adec92;
  wire adec93;
  wire adec94;
  wire adec95;
  wire adec96;
  wire adec97;
  wire adec98;
  wire adec99;
  wire adec9a;
  wire adec9b;
  wire adec9c;
  wire adec9d;
  wire adec9e;
  wire adec9f;
  wire adeca0;
  wire adeca1;
  wire adeca2;
  wire ade4a6;
  wire ade4a7;
  wire ade4a8;
  wire ade4a9;
  wire ade4aa;
  wire ade4ab;
  wire ade4ac;
  wire ade4ad;
  wire ade4ae;
  wire ade4af;
  wire ade4b0;
  wire ade4b1;
  wire ade4b2;
  wire ade4b3;
  wire ade4b4;
  wire ade4b5;
  wire ade4b6;
  wire ade4b7;
  wire ade4b8;
  wire ade4b9;
  wire v8f96d9;
  wire ade4ba;
  wire ade4bb;
  wire ade4bc;
  wire ade4bd;
  wire ade4be;
  wire ade4bf;
  wire ade4c0;
  wire ade4c1;
  wire ade4c2;
  wire ade4c3;
  wire ade4c4;
  wire ade4c5;
  wire ade4c6;
  wire ade4c7;
  wire ade4c8;
  wire c74620;
  wire c74621;
  wire ade4c9;
  wire ade4ca;
  wire ade4cb;
  wire ade4cc;
  wire ade4cd;
  wire ade4ce;
  wire ade4cf;
  wire ade4d0;
  wire ade4d1;
  wire ade4d2;
  wire ade4d3;
  wire ade4d4;
  wire ade4d5;
  wire ade4d6;
  wire ade4d7;
  wire ade4d8;
  wire ade4d9;
  wire ade4da;
  wire ade4db;
  wire ade4dc;
  wire ade4dd;
  wire ade4de;
  wire ade4df;
  wire ade4e0;
  wire ade4e1;
  wire ade4e2;
  wire ade4e3;
  wire ade4e4;
  wire ade4e5;
  wire ade4e6;
  wire ade4e7;
  wire ade4e8;
  wire ade4e9;
  wire ade4ea;
  wire ade4eb;
  wire ade4ec;
  wire ade4ed;
  wire ade4ee;
  wire ade4ef;
  wire ade4f0;
  wire ade4f1;
  wire ade4f2;
  wire ade4f3;
  wire ade540;
  wire ade541;
  wire ade542;
  wire ade543;
  wire ade544;
  wire ade545;
  wire ade546;
  wire ade547;
  wire ade548;
  wire ade549;
  wire ade54a;
  wire ade54b;
  wire ade54c;
  wire ade54d;
  wire ade54e;
  wire ade54f;
  wire ade550;
  wire ade551;
  wire ade552;
  wire ade553;
  wire ade554;
  wire ade555;
  wire ade556;
  wire ade557;
  wire ade558;
  wire ade559;
  wire ade55b;
  wire ade55c;
  wire ade55d;
  wire ade55e;
  wire ade55f;
  wire ade560;
  wire ade561;
  wire ade562;
  wire ade563;
  wire ade564;
  wire ade565;
  wire ade566;
  wire ade567;
  wire ade568;
  wire ade569;
  wire ade56a;
  wire ade56b;
  wire ade56c;
  wire ade56d;
  wire ade56e;
  wire ade56f;
  wire ade570;
  wire ade571;
  wire ade572;
  wire ade573;
  wire ade574;
  wire ade575;
  wire ade576;
  wire ade578;
  wire ade579;
  wire ade57a;
  wire ade57b;
  wire ade57c;
  wire ade57d;
  wire ade57e;
  wire ade57f;
  wire ade580;
  wire ade581;
  wire ade582;
  wire ade583;
  wire ade584;
  wire ade585;
  wire ade586;
  wire ade587;
  wire ade588;
  wire ade589;
  wire ade58a;
  wire ade58b;
  wire ade58c;
  wire ade58d;
  wire ade58e;
  wire ade58f;
  wire ade590;
  wire ade591;
  wire ade592;
  wire ade593;
  wire ade594;
  wire ade595;
  wire ade596;
  wire ade597;
  wire ade598;
  wire ade599;
  wire ade59a;
  wire ade59b;
  wire ade59c;
  wire ade59d;
  wire ade59e;
  wire ade59f;
  wire ade5a0;
  wire ade5a1;
  wire ade5a2;
  wire ade5a3;
  wire ade5a4;
  wire ade5a5;
  wire ade5a6;
  wire ade5a7;
  wire ade5a8;
  wire ade5a9;
  wire ade5aa;
  wire ade5ab;
  wire ade5ac;
  wire ade5ad;
  wire ade5ae;
  wire ade5af;
  wire ade5b0;
  wire ade5b1;
  wire ade5b2;
  wire ade5b3;
  wire ade5b4;
  wire ade5b5;
  wire ade5b6;
  wire ade5b7;
  wire ade5b8;
  wire ade5b9;
  wire ade5ba;
  wire ade5bb;
  wire ade5bc;
  wire ade5bd;
  wire ade5be;
  wire ade5bf;
  wire ade5c0;
  wire ade5c1;
  wire ade5c2;
  wire ade5c3;
  wire ade5c4;
  wire ade5c5;
  wire ade5c6;
  wire ade5c7;
  wire ade5c8;
  wire ade5c9;
  wire ade5ca;
  wire ade5cb;
  wire ade5cc;
  wire ade5cd;
  wire ade5ce;
  wire ade5cf;
  wire ade5d0;
  wire ade5d1;
  wire ade5d2;
  wire ade5d3;
  wire ade5d4;
  wire ade5d5;
  wire ade5d6;
  wire ade5d7;
  wire ade5d8;
  wire ade5d9;
  wire ade5da;
  wire ade5db;
  wire ade5dc;
  wire ade5dd;
  wire ade5de;
  wire ade5df;
  wire ade615;
  wire ade616;
  wire ade617;
  wire ade618;
  wire ade619;
  wire ade61a;
  wire ade61b;
  wire ade61c;
  wire ade61d;
  wire ade61e;
  wire ade61f;
  wire ade620;
  wire ade621;
  wire ade622;
  wire ade623;
  wire ade624;
  wire ade625;
  wire ade626;
  wire ade627;
  wire ade628;
  wire ade629;
  wire ade63c;
  wire ade63d;
  wire ade63e;
  wire ade64d;
  wire ade64e;
  wire ade64f;
  wire ade650;
  wire ade651;
  wire ade652;
  wire ade653;
  wire ade654;
  wire ade655;
  wire ade656;
  wire ade657;
  wire ade658;
  wire ade659;
  wire ade65a;
  wire ade65b;
  wire ade65c;
  wire ade65d;
  wire ade65e;
  wire ade65f;
  wire ade660;
  wire ade661;
  wire ade662;
  wire ade665;
  wire ade666;
  wire ade667;
  wire c749e5;
  wire c74b29;
  wire v9c81a4;
  wire v9f21c4;
  wire v9f21c5;
  wire v9ea3e1;
  wire v9ea3e2;
  wire v9ea3e3;
  wire v845582;
  wire c6d405;
  wire c6d406;
  wire c6d407;
  wire b06719;
  wire v9f20a1;
  wire v9ea3e4;
  wire v9ea3e5;
  wire v9ea3e6;
  wire v9ea3e7;
  wire v9ea3e8;
  wire v9ea3e9;
  wire v9ea3ea;
  wire v9ea3eb;
  wire v9ea3ec;
  wire v9ea3ed;
  wire v9ea3ee;
  wire v9ea3ef;
  wire v9ea3f0;
  wire v9ea3f1;
  wire v9ea3f2;
  wire v9ea3f3;
  wire v9ea3f4;
  wire v9ea3f5;
  wire v9ea3f6;
  wire v9ea3f7;
  wire v9ea3f8;
  wire v9ea3f9;
  wire v9ea3fa;
  wire v9ea3fb;
  wire v9ea3fc;
  wire v9ea3fd;
  wire v9ea3fe;
  wire v9ea3ff;
  wire v9ea400;
  wire v9ea401;
  wire v9ea402;
  wire v9ea403;
  wire v9ea404;
  wire v9ea405;
  wire v9ea406;
  wire v9ea407;
  wire v9ea408;
  wire v9ea409;
  wire v9ea40a;
  wire v9ea40b;
  wire v9ea40c;
  wire v9ea40d;
  wire v9f21c6;
  wire v9ea40e;
  wire v9ea40f;
  wire v9ea410;
  wire v84557e;
  wire v9ea411;
  wire v9ea412;
  wire v9ea413;
  wire v9ea414;
  wire v9ea415;
  wire v9ea416;
  wire v9ea417;
  wire v9ea418;
  wire v9ea419;
  wire v9ea41a;
  wire v9ea41b;
  wire v9ea41c;
  wire v9ea41d;
  wire v9ea41e;
  wire v9ea41f;
  wire v9ea420;
  wire v9ea421;
  wire v9ea422;
  wire v9ea423;
  wire v9ea424;
  wire v9ea425;
  wire v9ea426;
  wire v9ea427;
  wire v9ea428;
  wire v9ea429;
  wire v9ea42a;
  wire v9ea42b;
  wire v9ea42d;
  wire v9ea42e;
  wire v9ea42f;
  wire v9ea430;
  wire v9ea431;
  wire v9ea432;
  wire v9ea433;
  wire v9ea434;
  wire v9ea435;
  wire v9ea436;
  wire v9ea437;
  wire v9ea438;
  wire v9ea439;
  wire v9ea43a;
  wire v9ea43b;
  wire v9ea43c;
  wire v9ea43d;
  wire v9ea43e;
  wire v9ea43f;
  wire v9ea440;
  wire v9ea441;
  wire v9ea442;
  wire v9ea443;
  wire v9ea444;
  wire v9ea445;
  wire v9ea446;
  wire v9ea447;
  wire v9ea448;
  wire v9ea449;
  wire v9ea44a;
  wire v9ea44b;
  wire v9ea44c;
  wire v9ea44d;
  wire v9ea44e;
  wire v9ea44f;
  wire v9ea450;
  wire v9ea451;
  wire v9ea452;
  wire v9ea453;
  wire v9ea454;
  wire v9ea455;
  wire v9ea456;
  wire v9ea457;
  wire v9ea458;
  wire v9ea459;
  wire v9ea45a;
  wire v9ea45b;
  wire v9ea45c;
  wire v9ea45d;
  wire v9ea45e;
  wire v9ea45f;
  wire v9ea460;
  wire v9ea461;
  wire v9ea462;
  wire v9ea463;
  wire v9ea464;
  wire v9ea465;
  wire v9ea466;
  wire v9ea467;
  wire v9ea46a;
  wire v9ea46b;
  wire v9ea46c;
  wire v9ea46d;
  wire v9ea46e;
  wire v9ea46f;
  wire v9ea470;
  wire v9ea471;
  wire v9ea472;
  wire v9ea473;
  wire v9ea474;
  wire v9ea475;
  wire v9ea476;
  wire v9ea477;
  wire v9ea478;
  wire v9ea479;
  wire v9ea47a;
  wire v9ea47b;
  wire v9ea47c;
  wire v9ea47d;
  wire v9ea47e;
  wire v9ea47f;
  wire v9ea480;
  wire v9ea481;
  wire v9ea482;
  wire v9ea483;
  wire v9ea484;
  wire v9ea485;
  wire v9ea486;
  wire v9ea487;
  wire v9ea488;
  wire v9ea489;
  wire v9ea48a;
  wire v9ea48b;
  wire v9ea48c;
  wire v9ea48d;
  wire v9ea48e;
  wire v9ea48f;
  wire v9ea490;
  wire v9ea491;
  wire v9ea492;
  wire v9ea493;
  wire v9ea494;
  wire v9ea495;
  wire v9ea496;
  wire v9ea497;
  wire v9ea498;
  wire v9ea499;
  wire v9ea49a;
  wire v9ea49b;
  wire v9ea49c;
  wire v9ea49d;
  wire v9ea49e;
  wire v9ea49f;
  wire v9ea4a0;
  wire v9ea4a1;
  wire v9ea4a2;
  wire v9ea4a3;
  wire v9ea4a4;
  wire v9ea4a5;
  wire v9ea4a6;
  wire v9ea4a7;
  wire v9ea4a8;
  wire v9ea4a9;
  wire v9ea4aa;
  wire v9ea4ab;
  wire v9ea4ac;
  wire v9ea4ad;
  wire v9ea4ae;
  wire v9ea4af;
  wire v9ea4b0;
  wire v9ea4b1;
  wire v9ea4b2;
  wire v9ea4b3;
  wire v9ea4b4;
  wire v9ea4b5;
  wire v9ea4b6;
  wire v9ea4b7;
  wire v9ea4b8;
  wire v9ea4b9;
  wire v9ea4ba;
  wire v9ea4bb;
  wire v9ea4bc;
  wire v9ea4bd;
  wire v9ea4be;
  wire v9ea4bf;
  wire v9ea4c0;
  wire v9ea4c1;
  wire v9ea4c2;
  wire v9ea4c3;
  wire v9ea4c4;
  wire v9ea4c5;
  wire v9ea4c6;
  wire v9ea4c7;
  wire v9ea4c8;
  wire v9ea4c9;
  wire v9ea4ca;
  wire v9ea4cb;
  wire v9ea4cc;
  wire v9ea4cd;
  wire v9ea4ce;
  wire v9ea4cf;
  wire v9ea4d0;
  wire v9ea4d1;
  wire v9ea4d2;
  wire v9ea4d3;
  wire v9ea4d4;
  wire v9ea4d5;
  wire v9ea4d6;
  wire v9ea4d7;
  wire v9ea4d8;
  wire v9ea4d9;
  wire v9ea4da;
  wire v9ea4db;
  wire v9ea4dc;
  wire v9ea4dd;
  wire v9ea4de;
  wire v9ea4df;
  wire v9ea4e0;
  wire v9ea4e1;
  wire v9ea4e2;
  wire v9ea4e3;
  wire v9ea4e4;
  wire v9ea4e5;
  wire v9ea4e6;
  wire v9ea566;
  wire v9ea567;
  wire v9ea568;
  wire v9ea569;
  wire v9ea56a;
  wire v9ea56b;
  wire v9ea56c;
  wire v9ea56d;
  wire v9ea56e;
  wire v9ea56f;
  wire v9ea570;
  wire v9ea571;
  wire v9ea572;
  wire v9ea573;
  wire v9ea574;
  wire v9ea575;
  wire v9ea576;
  wire v9ea577;
  wire v9ea578;
  wire v9ea579;
  wire v9ea57a;
  wire v9ea57b;
  wire v9ea57c;
  wire v9ea57d;
  wire v9ea57e;
  wire v9ea57f;
  wire v9ea580;
  wire v9ea581;
  wire v9ea582;
  wire v9ea583;
  wire v9ea584;
  wire v9ea585;
  wire v9ea586;
  wire v9ea587;
  wire v9ea588;
  wire v9ea589;
  wire v9ea58a;
  wire v9ea58b;
  wire v9ea58c;
  wire v9ea58d;
  wire v9ea58e;
  wire v9ea58f;
  wire v9ea590;
  wire v9ea591;
  wire v9ea592;
  wire v9ea593;
  wire v9ea594;
  wire v9ea595;
  wire v9ea596;
  wire v9ea597;
  wire v9ea598;
  wire v9ea599;
  wire v9ea59a;
  wire v9ea59b;
  wire v9ea59c;
  wire v9ea59d;
  wire v9ea59e;
  wire v9ea59f;
  wire v9ea5a0;
  wire v9ea5a1;
  wire v9ea5a2;
  wire v9ea5a3;
  wire v9ea5a4;
  wire v9ea5a5;
  wire v9ea5a6;
  wire v9ea5a7;
  wire v9ea5a8;
  wire v9ea5a9;
  wire v9ea5aa;
  wire v9ea5ab;
  wire v9ea5ac;
  wire v9ea5ad;
  wire v9ea5ae;
  wire v9ea5af;
  wire v9ea5b0;
  wire v9ea5b1;
  wire v9ea5b2;
  wire v9ea5b3;
  wire v9ea5b4;
  wire v9ea5b5;
  wire v9ea5b6;
  wire v9ea5b7;
  wire v9ea5b8;
  wire v9ea5b9;
  wire v9ea5ba;
  wire v9ea5bb;
  wire v9ea5bc;
  wire v9ea5bd;
  wire v9ea5be;
  wire v9ea5ca;
  wire v9ea5cb;
  wire v9ea5cc;
  wire v9ea5cd;
  wire v9ea5ce;
  wire v9ea5cf;
  wire v9ea5d0;
  wire v9ea5d1;
  wire v9ea5d2;
  wire v9ea5d3;
  wire v9ea5d4;
  wire v9ea5d5;
  wire v9ea5d6;
  wire v9ea5d7;
  wire v9ea5d8;
  wire v9ea5d9;
  wire v9ea5da;
  wire v9ea5db;
  wire v9ea5dc;
  wire v9ea5dd;
  wire v9ea5de;
  wire v9ea5df;
  wire v9ea5e0;
  wire v9ea5e1;
  wire v9ea5e2;
  wire v9ea5e3;
  wire v9ea5e4;
  wire v9ea5e5;
  wire v9ea5e6;
  wire v9ea5e7;
  wire v9ea5e8;
  wire v9ea5e9;
  wire v9ea5ea;
  wire v9ea5eb;
  wire v9ea5f3;
  wire v9ea5f4;
  wire v9ea5f5;
  wire v9ea5f6;
  wire v9ea5f7;
  wire v9ea5f8;
  wire v9ea5f9;
  wire v9ea5fa;
  wire v9ea602;
  wire v9ea603;
  wire v9ea604;
  wire v9ea605;
  wire v9ea606;
  wire v9ea607;
  wire v9ea608;
  wire v9ea609;
  wire v9ea60a;
  wire v9ea60b;
  wire v9ea60c;
  wire v9ea60d;
  wire v9ea60e;
  wire v9ea60f;
  wire v9ea610;
  wire v9ea611;
  wire v9ea612;
  wire v9ea613;
  wire v9ea614;
  wire v9ea615;
  wire v9ea616;
  wire v9ea617;
  wire v9ea618;
  wire v9ea619;
  wire v9ea61a;
  wire v9ea61b;
  wire v9ea61c;
  wire v9ea61d;
  wire v9ea61e;
  wire v9ea61f;
  wire v9ea620;
  wire v9ea621;
  wire v9ea622;
  wire v9ea623;
  wire v9ea624;
  wire v9ea625;
  wire v9ea626;
  wire v9ea627;
  wire v9ea628;
  wire v9e9e67;
  wire v9e9e68;
  wire v9e9e69;
  wire v9e9e6a;
  wire v9e9e6b;
  wire v9e9e6c;
  wire v9e9e6d;
  wire v9e9e6e;
  wire v9e9e6f;
  wire v9e9e70;
  wire v9e9e71;
  wire v9e9e72;
  wire v9e9e73;
  wire v9e9e74;
  wire v9e9e75;
  wire v9e9e76;
  wire v9e9e77;
  wire v9e9e78;
  wire v9e9e79;
  wire v9e9e7a;
  wire v9e9e7b;
  wire v9e9e7c;
  wire v9e9e7d;
  wire v9e9e7e;
  wire v9e9e9a;
  wire v9e9e9b;
  wire v9e9e9c;
  wire v9e9e9d;
  wire v9e9e9e;
  wire v9e9e9f;
  wire v9e9ea0;
  wire v9e9ea1;
  wire v9e9ea2;
  wire v9e9ea3;
  wire v9e9ea4;
  wire v9e9ea5;
  wire v9e9ea6;
  wire v9e9ea7;
  wire v9e9ea8;
  wire v9e9ea9;
  wire v9e9eaa;
  wire v9e9eab;
  wire v9e9eac;
  wire v9e9ead;
  wire v9e9eae;
  wire v9e9eaf;
  wire v9e9eb0;
  wire v9e9eb1;
  wire v9e9eb2;
  wire v9e9eb3;
  wire v9e9eb4;
  wire v9e9eb5;
  wire v9e9eb6;
  wire v9e9eb7;
  wire v9e9eb8;
  wire v9e9eb9;
  wire v9e9eba;
  wire v9e9ebb;
  wire v9e9ebc;
  wire v9e9ebd;
  wire v9e9ebe;
  wire v9e9ebf;
  wire v9e9ec0;
  wire v9e9ec1;
  wire v9e9ec2;
  wire v9e9ec3;
  wire v9e9ec4;
  wire v9e9ec5;
  wire v9e9ec6;
  wire v9e9ec7;
  wire v9e9ec8;
  wire v9e9ec9;
  wire v9e9eca;
  wire v9e9ecb;
  wire v9e9ecc;
  wire v9e9ecd;
  wire v9e9ece;
  wire v9e9ecf;
  wire v9e9ed0;
  wire v9e9ed1;
  wire v9e9ed2;
  wire v9e9ed3;
  wire v9e9ed4;
  wire v9e9ed5;
  wire v9e9ed6;
  wire v9e9ed7;
  wire v9e9ed8;
  wire v9e9ed9;
  wire v9e9eda;
  wire v9e9edb;
  wire v9e9edc;
  wire v9e9edd;
  wire v9e9ede;
  wire v9e9edf;
  wire v9e9ee0;
  wire v9e9ee1;
  wire v9e9ee2;
  wire v9e9ee3;
  wire v9e9ee4;
  wire v9e9ee5;
  wire v9e9ee6;
  wire v9e9ee7;
  wire v9e9ee8;
  wire v9e9ee9;
  wire v9e9eea;
  wire v9e9eeb;
  wire v9e9eec;
  wire v9e9eed;
  wire v9e9eee;
  wire v9e9eef;
  wire v9e9ef0;
  wire v9e9ef1;
  wire v9e9ef2;
  wire v9e9ef3;
  wire v9e9ef4;
  wire v9e9ef5;
  wire v9e9ef6;
  wire v9e9ef7;
  wire v9e9f49;
  wire v9e9f4a;
  wire v9e9f4c;
  wire v9e9f4d;
  wire v9e9f4e;
  wire v9e9f4f;
  wire v9e9f50;
  wire v9e9f51;
  wire v9e9f52;
  wire v9e9f53;
  wire v9e9f54;
  wire v9e9f55;
  wire v9e9f56;
  wire v9e9f57;
  wire v9e9f58;
  wire v9e9f59;
  wire v9e9f5a;
  wire v9e9f5b;
  wire v9e9f5c;
  wire v9e9f5d;
  wire v9e9f5e;
  wire v9e9f5f;
  wire v9e9f60;
  wire v9e9f61;
  wire v9e9f62;
  wire v9e9f63;
  wire v9e9f64;
  wire v9e9f65;
  wire v9e9f66;
  wire v9e9f67;
  wire v9e9f68;
  wire v9e9f69;
  wire v9e9f6a;
  wire v9e9f6b;
  wire v9e9f6c;
  wire v9e9f6d;
  wire v9e9f6e;
  wire v9e9f6f;
  wire v9e9f70;
  wire v9e9f71;
  wire v9e9f72;
  wire v9e9f73;
  wire v9e9f74;
  wire v9e9f75;
  wire v9e9f76;
  wire v9e9f77;
  wire v9e9f78;
  wire v9e9f79;
  wire v9e9f7a;
  wire v9e9f7b;
  wire v9e9f7c;
  wire v9e9f7d;
  wire v9e9f7e;
  wire v9e9f7f;
  wire v9e9f80;
  wire v9e9f81;
  wire v9e9f82;
  wire v9e9f83;
  wire v9e9f84;
  wire v9e9f85;
  wire v9e9f86;
  wire v9e9f87;
  wire v9e9f88;
  wire v9e9f89;
  wire v9e9f8a;
  wire v9e9f8b;
  wire v9e9f8c;
  wire v9e9f8d;
  wire v9e9f8e;
  wire v9e9f8f;
  wire v9e9f90;
  wire v9e9f91;
  wire v9e9f92;
  wire v9e9f93;
  wire v9e9f94;
  wire v9e9f95;
  wire v9e9f96;
  wire v9e9f97;
  wire v9e9f98;
  wire v9e9f99;
  wire v9e9f9a;
  wire v9e9f9b;
  wire v9e9f9c;
  wire v9e9f9d;
  wire v9e9f9e;
  wire v9e9f9f;
  wire v9e9fa0;
  wire v9e9fa1;
  wire v9e9fa2;
  wire v9e9fa3;
  wire v9e9fa4;
  wire v9e9fa5;
  wire v9e9fa6;
  wire v9e9fa7;
  wire v9e9fa8;
  wire v9e9fa9;
  wire v9e9faa;
  wire v9e9fab;
  wire v9e9fac;
  wire v9e9fad;
  wire v9e9fae;
  wire v9e9faf;
  wire v9e9fb0;
  wire v9e9fb1;
  wire v9e9fb2;
  wire v9e9fb3;
  wire v9e9fb4;
  wire v9e9fb5;
  wire v9e9fb6;
  wire v9e9fb7;
  wire v9e9fb8;
  wire v9e9fb9;
  wire v9e9fba;
  wire v9e9fbb;
  wire v9e9fbc;
  wire v9e9fbd;
  wire v9e9fbe;
  wire v9e9fbf;
  wire v9e9fc0;
  wire v9e9fc1;
  wire v9e9fc2;
  wire v9e9fc3;
  wire v9e9fc4;
  wire v9e9fc5;
  wire v9e9fc6;
  wire v9e9fc7;
  wire v9e9fc8;
  wire v9e9fc9;
  wire v9e9fca;
  wire v9e9fcb;
  wire v9e9fcc;
  wire v9e9fcd;
  wire v9e9fce;
  wire v9e9fcf;
  wire v9e9fd0;
  wire v9e9fd1;
  wire v9e9fd2;
  wire v9e9fd3;
  wire v9e9fd4;
  wire v9e9fd5;
  wire v9e9fd6;
  wire v9e9fd7;
  wire v9e9fd8;
  wire v9e9fd9;
  wire v9e9fda;
  wire v9e9fdb;
  wire v9e9fdc;
  wire v9e9fdd;
  wire v9e9fde;
  wire v9e9fdf;
  wire v9e9fe0;
  wire v9e9fe1;
  wire v9e9fe2;
  wire v9e9fe3;
  wire v9e9fe4;
  wire v9e9fe5;
  wire v9e9fe6;
  wire v9e9fe7;
  wire v9e9fe8;
  wire v9e9fe9;
  wire v8da59e;
  wire v84556e;
  wire v8da59f;
  wire v8da5a0;
  wire v8da5a1;
  wire v8da5a4;
  wire v8da5a6;
  wire v8da603;
  wire v8da604;
  wire dc4f61;
  wire dc4f62;
  wire dc4f63;
  wire dc4f64;
  wire dc4f66;
  wire dc4f67;
  wire dc4f68;
  wire dc4f69;
  wire dc4f6a;
  wire dc4f6b;
  wire dc4f6c;
  wire dc4f6d;
  wire dc4f6e;
  wire dc4f6f;
  wire dc4f70;
  wire dc4f71;
  wire dc4f72;
  wire dc4f73;
  wire dc4f74;
  wire dc4f75;
  wire dc4f76;
  wire dc4f77;
  wire dc4f78;
  wire bbb7c6;
  wire bbb7c7;
  wire dc4f79;
  wire dc4f7a;
  wire dc4f7b;
  wire dc4f7c;
  wire dc4f7d;
  wire dc4f7e;
  wire dc4f7f;
  wire dc4f80;
  wire dc4f81;
  wire dc4f82;
  wire dc4f83;
  wire dc4f84;
  wire dc4f85;
  wire dc4f86;
  wire dc4f87;
  wire dc4f88;
  wire dc4f89;
  wire dc4f8a;
  wire dc4f8b;
  wire dc4f8c;
  wire dc4f8d;
  wire dc4f8e;
  wire dc4f8f;
  wire dc4f90;
  wire dc4f91;
  wire dc4f92;
  wire dc4f93;
  wire dc4f94;
  wire dc4f96;
  wire dc4f97;
  wire dc4f98;
  wire dc4f9a;
  wire dc4f9b;
  wire dc4f9c;
  wire dc4f9d;
  wire dc4f9e;
  wire dc4f9f;
  wire dc4fa0;
  wire dc4fa1;
  wire dc4fa2;
  wire dc4fa3;
  wire dc4fa4;
  wire dc4fa5;
  wire dc4fa6;
  wire dc4fa7;
  wire dc4fa8;
  wire dc4fa9;
  wire dc4faa;
  wire dc4fab;
  wire dc4fac;
  wire dc4fad;
  wire dc4fae;
  wire dc4faf;
  wire dc4fb0;
  wire dc4fb1;
  wire dc4fb2;
  wire dc4fb3;
  wire dc4fb4;
  wire dc4fb5;
  wire dc4fb6;
  wire dc4fb7;
  wire dc4fb8;
  wire dc4fb9;
  wire dc4fba;
  wire dc4fbb;
  wire dc4fbc;
  wire dc4fbd;
  wire dc4fbe;
  wire dc4fbf;
  wire dc4fc0;
  wire dc4fc1;
  wire dc4fc3;
  wire dc4fc4;
  wire dc4fc5;
  wire dc4fc6;
  wire dc4fc7;
  wire dc4fc8;
  wire dc4fc9;
  wire dc4fca;
  wire dc4fcb;
  wire dc4fcc;
  wire dc4fcd;
  wire dc4fce;
  wire dc4fcf;
  wire dc4fd0;
  wire dc4fd1;
  wire dc4fd2;
  wire dc4fd3;
  wire dc4fd4;
  wire dc4fd5;
  wire dc4fd6;
  wire dc4fd7;
  wire dc4fd8;
  wire dc4fd9;
  wire dc4fda;
  wire dc4fdb;
  wire dc4fdc;
  wire dc4fdd;
  wire dc4fdf;
  wire dc4fe0;
  wire dc4fe1;
  wire dc4fe2;
  wire dc4fe3;
  wire dc4fe4;
  wire dc4fe5;
  wire dc4fe6;
  wire dc4fe7;
  wire dc4fe8;
  wire dc4fe9;
  wire dc4fea;
  wire dc4feb;
  wire dc4fec;
  wire dc4fed;
  wire dc4fee;
  wire dc4fef;
  wire dc4ff0;
  wire dc4ff1;
  wire dc4ff2;
  wire dc4ff3;
  wire dc4ff4;
  wire dc4ff5;
  wire dc4ff6;
  wire dc4ff7;
  wire dc4ff8;
  wire dc4ff9;
  wire dc4ffa;
  wire dc4ffb;
  wire dc4ffc;
  wire dc4ffd;
  wire dc4ffe;
  wire dc4fff;
  wire dc5000;
  wire dc5001;
  wire dc5002;
  wire dc5003;
  wire dc5004;
  wire dc5005;
  wire dc5006;
  wire dc5007;
  wire dc5008;
  wire dc5009;
  wire dc500a;
  wire dc500b;
  wire dc500c;
  wire dc500d;
  wire dc500e;
  wire dc500f;
  wire dc5010;
  wire dc5011;
  wire dc5012;
  wire dc5013;
  wire dc5014;
  wire dc5015;
  wire dc5016;
  wire dc5017;
  wire dc5018;
  wire dc5019;
  wire dc501a;
  wire dc501b;
  wire dc501c;
  wire dc501d;
  wire dc501e;
  wire dc501f;
  wire dc5020;
  wire dc5021;
  wire dc5022;
  wire dc5023;
  wire dc5024;
  wire dc5025;
  wire dc5026;
  wire dc5027;
  wire dc5028;
  wire dc5029;
  wire dc502a;
  wire dc502b;
  wire dc502c;
  wire dc502d;
  wire dc502e;
  wire dc502f;
  wire dc5030;
  wire dc5031;
  wire dc5032;
  wire dc5033;
  wire dc5034;
  wire dc5035;
  wire dc5036;
  wire dc5037;
  wire dc5038;
  wire dc503a;
  wire dc503b;
  wire dc503c;
  wire dc503d;
  wire dc503e;
  wire dc503f;
  wire dc5040;
  wire dc5041;
  wire dc5042;
  wire dc5043;
  wire dc5044;
  wire dc5045;
  wire dc5046;
  wire dc5047;
  wire dc5048;
  wire dc5049;
  wire dc504a;
  wire dc504b;
  wire bbbe35;
  wire bbbe36;
  wire dc504c;
  wire dc504d;
  wire dc504e;
  wire dc504f;
  wire dc5050;
  wire dc5051;
  wire dc5052;
  wire dc5053;
  wire dc5054;
  wire dc5055;
  wire dc5056;
  wire dc5057;
  wire dc5058;
  wire dc5059;
  wire dc505a;
  wire dc505b;
  wire dc505c;
  wire dc505d;
  wire dc505e;
  wire dc505f;
  wire dc5060;
  wire dc5061;
  wire dc5062;
  wire dc5063;
  wire dc5064;
  wire dc5065;
  wire dc5066;
  wire dc5067;
  wire dc5068;
  wire dc5069;
  wire dc506a;
  wire dc506b;
  wire dc506c;
  wire dc506d;
  wire dc506e;
  wire dc506f;
  wire dc5070;
  wire dc5071;
  wire dc5072;
  wire dc5073;
  wire dc5074;
  wire dc5075;
  wire dc5076;
  wire dc5077;
  wire dc5079;
  wire dc507a;
  wire dc507b;
  wire dc507c;
  wire dc507d;
  wire dc507e;
  wire dc507f;
  wire dc5080;
  wire dc5081;
  wire dc5082;
  wire dc5085;
  wire dc5086;
  wire dc5087;
  wire v84556a;
  wire dc5088;
  wire dc5089;
  wire dc52f8;
  wire dc52f9;
  wire dc52fa;
  wire dc52fb;
  wire dc52fc;
  wire dc52fd;
  wire dc52fe;
  wire dc52ff;
  wire dc5300;
  wire dc5301;
  wire dc5302;
  wire dc5303;
  wire dc5307;
  wire dc5311;
  wire dc5314;
  wire dc5315;
  wire dc5316;
  wire dc5317;
  wire dc5318;
  wire dc5319;
  wire dc531a;
  wire dc531b;
  wire dc531c;
  wire dc531d;
  wire dc531e;
  wire dc531f;
  wire dc5320;
  wire dc5385;
  wire dc5386;
  wire dc5387;
  wire dc5388;
  wire dc5389;
  wire dc538a;
  wire dc538b;
  wire dc538c;
  wire dc538d;
  wire dc538e;
  wire dc538f;
  wire dc5390;
  wire dc5391;
  wire dc5392;
  wire dc5393;
  wire dc5394;
  wire dc539c;
  wire dc539d;
  wire dc539e;
  wire dc539f;
  wire dc53a0;
  wire dc53a1;
  wire dc53a2;
  wire dc53a3;
  wire dc53a4;
  wire dc53a5;
  wire dc53a6;
  wire dc53a7;
  wire dc53a8;
  wire dc53a9;
  wire dc53aa;
  wire dc53b2;
  wire dc53b3;
  wire dc53b4;
  wire dc53b5;
  wire dc53b6;
  wire dc53b7;
  wire dc53b8;
  wire dc53b9;
  wire dc53ba;
  wire dc53bb;
  wire dc53bc;
  wire dc53bd;
  wire dc53be;
  wire dc53bf;
  wire dc53c0;
  wire dc53c1;
  wire dc53c2;
  wire dc53c3;
  wire dc53c4;
  wire dc53c5;
  wire dc53c6;
  wire dc53c7;
  wire dc53c8;
  wire dc53c9;
  wire dc53ca;
  wire dc53cb;
  wire dc53cc;
  wire dc53cd;
  wire dc53ce;
  wire dc53cf;
  wire dc53d0;
  wire dc53d1;
  wire dc53d2;
  wire dc53d5;
  wire dc53d6;
  wire dc53d7;
  wire dc53d8;
  wire dc53d9;
  wire dc53da;
  wire dc53db;
  wire dc53dc;
  wire dc53dd;
  wire dc53de;
  wire dc53df;
  wire dc53e0;
  wire df54d6;
  wire df54d7;
  wire df54d8;
  wire df54d9;
  wire df54da;
  wire df54db;
  wire df54dc;
  wire df54dd;
  wire e0edf9;
  wire df54de;
  wire df54df;
  wire df54e0;
  wire df54e1;
  wire df54e2;
  wire df54e3;
  wire df54e4;
  wire df54e5;
  wire df54e6;
  wire df54e7;
  wire df54e8;
  wire df54e9;
  wire df54ea;
  wire df54eb;
  wire df54ed;
  wire df54ee;
  wire df54ef;
  wire df54f0;
  wire df54f2;
  wire df54f3;
  wire df54f4;
  wire df54f5;
  wire df54f6;
  wire df54f7;
  wire df54f8;
  wire df54f9;
  wire df54fa;
  wire df54fb;
  wire df54fc;
  wire df54fd;
  wire df54ff;
  wire df552b;
  wire df552c;
  wire df552d;
  wire df552e;
  wire df552f;
  wire df5530;
  wire df5531;
  wire df5532;
  wire df5533;
  wire df5534;
  wire df5535;
  wire df5536;
  wire df5537;
  wire df5538;
  wire df5539;
  wire df553a;
  wire df553b;
  wire df553c;
  wire df553d;
  wire df553e;
  wire df553f;
  wire df5540;
  wire df5541;
  wire df5542;
  wire df5543;
  wire df5544;
  wire df5078;
  wire df5079;
  wire df507a;
  wire df507b;
  wire df507c;
  wire df507d;
  wire df507e;
  wire df50cb;
  wire df50cc;
  wire df50cd;
  wire df50ce;
  wire df50cf;
  wire df50d0;
  wire df50d1;
  wire df50d2;
  wire df50d3;
  wire df50d4;
  wire df50d5;
  wire df50d6;
  wire df50d7;
  wire df50d8;
  wire df50d9;
  wire df50da;
  wire df50db;
  wire df50dc;
  wire df50dd;
  wire df50de;
  wire df5114;
  wire df5115;
  wire df5116;
  wire df5117;
  wire df5118;
  wire df5119;
  wire df511a;
  wire df511b;
  wire df511c;
  wire df511d;
  wire df5124;
  wire df5125;
  wire df5126;
  wire df5127;
  wire df5128;
  wire df5129;
  wire df512a;
  wire df512b;
  wire df512c;
  wire df512d;
  wire df512e;
  wire df512f;
  wire df5130;
  wire df5131;
  wire df5132;
  wire df5133;
  wire df5134;
  wire df5135;
  wire df5136;
  wire df5137;
  wire df5138;
  wire df5139;
  wire df513a;
  wire df513b;
  wire df513c;
  wire df513d;
  wire df513e;
  wire df513f;
  wire df5140;
  wire df5141;
  wire df5142;
  wire df5143;
  wire df5144;
  wire df5145;
  wire df5146;
  wire df5147;
  wire df5148;
  wire df5149;
  wire df514a;
  wire df514b;
  wire df514c;
  wire df514d;
  wire df514e;
  wire df514f;
  wire df5150;
  wire df5151;
  wire df5152;
  wire df5153;
  wire df5154;
  wire df5155;
  wire df5156;
  wire df5157;
  wire df5158;
  wire df5159;
  wire df515a;
  wire df515b;
  wire df515c;
  wire df515d;
  wire df515e;
  wire df515f;
  wire df5160;
  wire df5161;
  wire df5162;
  wire df5163;
  wire df5164;
  wire df5165;
  wire df5166;
  wire df5167;
  wire df5168;
  wire df5169;
  wire df516a;
  wire df516b;
  wire df516c;
  wire df516d;
  wire df516e;
  wire df516f;
  wire df5170;
  wire df5171;
  wire df5172;
  wire df5173;
  wire df5174;
  wire df5175;
  wire df5176;
  wire df5177;
  wire df5178;
  wire df5179;
  wire df517a;
  wire df517b;
  wire df517c;
  wire df517d;
  wire df517e;
  wire df517f;
  wire df5182;
  wire df5183;
  wire df5184;
  wire df5185;
  wire df5186;
  wire df5187;
  wire df5188;
  wire df5189;
  wire df518a;
  wire df518b;
  wire df518c;
  wire df518d;
  wire df518e;
  wire df518f;
  wire df5190;
  wire df5191;
  wire df5192;
  wire df5193;
  wire df5194;
  wire df5195;
  wire df5196;
  wire df5197;
  wire df5198;
  wire df5199;
  wire df519a;
  wire df519b;
  wire df519c;
  wire df519d;
  wire df519e;
  wire df519f;
  wire df51a0;
  wire df51a1;
  wire df51a2;
  wire df51a3;
  wire df51a4;
  wire df51a5;
  wire df51a6;
  wire df51a7;
  wire df51a8;
  wire df51a9;
  wire df51aa;
  wire df51ab;
  wire df51ac;
  wire df51ad;
  wire df51ae;
  wire df51af;
  wire df51b0;
  wire df51b1;
  wire df51b2;
  wire df51b3;
  wire df51b4;
  wire df51b5;
  wire df51b6;
  wire df51b7;
  wire df51b8;
  wire df51b9;
  wire df51ba;
  wire df51bb;
  wire df51bc;
  wire df51bd;
  wire df51be;
  wire df51bf;
  wire df51c0;
  wire df51c1;
  wire df51c2;
  wire df51c3;
  wire df51c4;
  wire df51c5;
  wire df51c6;
  wire df51c7;
  wire df51c8;
  wire df51c9;
  wire df51ca;
  wire df51cb;
  wire df51cc;
  wire df51cd;
  wire df51ce;
  wire df51cf;
  wire df51d0;
  wire df51d1;
  wire df51d2;
  wire df51d3;
  wire df51d4;
  wire df51d5;
  wire df51da;
  wire df51db;
  wire df51dc;
  wire df51dd;
  wire df51de;
  wire df51df;
  wire df51e0;
  wire v845556;
  wire d358e8;
  wire d358ea;
  wire d358eb;
  wire d358ec;
  wire d358ed;
  wire d358ee;
  wire d358ef;
  wire d358f0;
  wire d358f1;
  wire d358f2;
  wire d358f3;
  wire d358f4;
  wire d358f5;
  wire d358f6;
  wire d358f8;
  wire d358f9;
  wire d358fa;
  wire d358fb;
  wire d358fc;
  wire d358fd;
  wire d358fe;
  wire d358ff;
  wire d35900;
  wire d35902;
  wire d35903;
  wire d35905;
  wire d35906;
  wire d35907;
  wire d35908;
  wire d35909;
  wire d3590a;
  wire d3590b;
  wire d3590c;
  wire d3590d;
  wire d3590e;
  wire d3590f;
  wire d35910;
  wire d35911;
  wire d35912;
  wire d35913;
  wire d35914;
  wire d35915;
  wire d35916;
  wire d35917;
  wire d35918;
  wire d35919;
  wire d3591a;
  wire d3591b;
  wire d3591c;
  wire d3591d;
  wire d3591e;
  wire d35920;
  wire d35921;
  wire d35949;
  wire d3594a;
  wire d3594b;
  wire d3594c;
  wire d3594d;
  wire d3594e;
  wire d3594f;
  wire d35950;
  wire d35951;
  wire d35952;
  wire d35953;
  wire d35954;
  wire d35955;
  wire d35956;
  wire d35957;
  wire d35958;
  wire d35959;
  wire d3595a;
  wire d3595b;
  wire d3597a;
  wire d3597b;
  wire d3597c;
  wire d3597d;
  wire d3597e;
  wire d3597f;
  wire d35980;
  wire d35981;
  wire d35982;
  wire d35983;
  wire d35984;
  wire d35985;
  wire d35986;
  wire d35987;
  wire d35988;
  wire d35989;
  wire d3598a;
  wire d3598b;
  wire d3598c;
  wire d3598d;
  wire d3598e;
  wire d3598f;
  wire d35991;
  wire d35992;
  wire d35993;
  wire d35994;
  wire d35995;
  wire d35996;
  wire d35997;
  wire d35998;
  wire d35999;
  wire d3599a;
  wire d3599b;
  wire d3599c;
  wire d3599d;
  wire d3599e;
  wire d3599f;
  wire d359a0;
  wire d359a1;
  wire d359a2;
  wire d359a3;
  wire d359a4;
  wire d359a5;
  wire d359a6;
  wire d359a7;
  wire d359a8;
  wire d359a9;
  wire d359aa;
  wire d359ab;
  wire d359ac;
  wire d359ad;
  wire d359ae;
  wire d359af;
  wire d359b0;
  wire d359b1;
  wire d359b2;
  wire d359b3;
  wire bbb31e;
  wire d359b4;
  wire d359b5;
  wire d359b6;
  wire d359b7;
  wire d359b8;
  wire d359b9;
  wire d359ba;
  wire d359bb;
  wire d359bc;
  wire d359bd;
  wire d359be;
  wire d359bf;
  wire d359c0;
  wire d359c1;
  wire d359c2;
  wire d359c3;
  wire d359c4;
  wire d359c5;
  wire d359c6;
  wire d359c7;
  wire d359c8;
  wire d359c9;
  wire d359ca;
  wire d359cb;
  wire d359cc;
  wire d359cd;
  wire d359ce;
  wire d359cf;
  wire d359d0;
  wire d359d1;
  wire d359d2;
  wire d359d3;
  wire d359d4;
  wire d359d5;
  wire d359d6;
  wire d359d7;
  wire d359d8;
  wire d359d9;
  wire d359da;
  wire d359db;
  wire d359dc;
  wire d359dd;
  wire d359de;
  wire d359df;
  wire d359e0;
  wire d359e1;
  wire d359e2;
  wire d359e3;
  wire d359e4;
  wire d359e5;
  wire d359e6;
  wire d359e7;
  wire d359e8;
  wire d359e9;
  wire d359ea;
  wire d359eb;
  wire d359ec;
  wire d359ed;
  wire d359ee;
  wire d359ef;
  wire d359f0;
  wire d359f1;
  wire d359f2;
  wire d359f3;
  wire d359f4;
  wire d359f5;
  wire d359f6;
  wire d359f7;
  wire d359f8;
  wire d359f9;
  wire d359fa;
  wire d359fb;
  wire d359fc;
  wire d359fd;
  wire d359fe;
  wire d359ff;
  wire d35a00;
  wire d35a01;
  wire d35a02;
  wire d35a03;
  wire d35a04;
  wire d35a05;
  wire d35a06;
  wire d35a07;
  wire d35a08;
  wire d35a09;
  wire d35a0a;
  wire d35a0b;
  wire d35a0c;
  wire d35a0d;
  wire d35a0e;
  wire d35a0f;
  wire d35a10;
  wire d35a11;
  wire d35a12;
  wire d35a13;
  wire d35a14;
  wire d35a15;
  wire d35a16;
  wire d35a17;
  wire d35a18;
  wire d35a19;
  wire d35a1a;
  wire d35a1b;
  wire d35a1c;
  wire d35a1d;
  wire d35a1e;
  wire d35a1f;
  wire d35a20;
  wire d35a21;
  wire d35a22;
  wire d35a23;
  wire d35a24;
  wire d35a25;
  wire d35a26;
  wire d35a27;
  wire d35a28;
  wire d35a29;
  wire d35a2a;
  wire d35a2b;
  wire d35a2d;
  wire d35a2e;
  wire d35a2f;
  wire d35a30;
  wire d35a31;
  wire d35a32;
  wire d35a33;
  wire d35a34;
  wire d35a35;
  wire d35a36;
  wire d35a37;
  wire d35a38;
  wire d35a39;
  wire d35a3a;
  wire d35a3b;
  wire d35a3c;
  wire d35a3d;
  wire d35a3e;
  wire d35a3f;
  wire d35a40;
  wire d35a41;
  wire d35a42;
  wire d35a43;
  wire d35a44;
  wire d35a45;
  wire d35a46;
  wire d35a47;
  wire d35a48;
  wire d35a49;
  wire d35a4a;
  wire d35a4b;
  wire d35a4c;
  wire d35a4d;
  wire d35a4e;
  wire d35a4f;
  wire d35a50;
  wire d35a51;
  wire d35a52;
  wire d35a53;
  wire d35a54;
  wire d35a55;
  wire d35a56;
  wire d35a57;
  wire d35a58;
  wire d35a59;
  wire d35a5a;
  wire d35a5b;
  wire d35a5c;
  wire d35a5d;
  wire d35a5e;
  wire d35a5f;
  wire d35a60;
  wire d35a61;
  wire d35a62;
  wire d35a63;
  wire d35a64;
  wire d35a65;
  wire d35a66;
  wire d35a67;
  wire d35a68;
  wire d35a69;
  wire d35a6a;
  wire d35a6b;
  wire d35a6c;
  wire d35a6d;
  wire d35a6e;
  wire d35a6f;
  wire d35a70;
  wire d35a71;
  wire d35a72;
  wire d35a73;
  wire d35a74;
  wire d35a75;
  wire d35a76;
  wire d35a77;
  wire d35a78;
  wire d35a79;
  wire d35a7a;
  wire d35a7b;
  wire d35a92;
  wire d35a93;
  wire d35a94;
  wire v84555a;
  wire d35a95;
  wire d35a96;
  wire d35a97;
  wire v845548;
  wire d35a98;
  wire d35a99;
  wire d35a9a;
  wire d35a9b;
  wire v84554a;
  wire d35a9c;
  wire d35a9d;
  wire d35a9e;
  wire d35a9f;
  wire d35aa0;
  wire d35aa1;
  wire d35aa2;
  wire d35aa3;
  wire v84554e;
  wire d35aa4;
  wire d35aa5;
  wire d35aa6;
  wire d35aa7;
  wire d35aa8;
  wire d35aa9;
  wire d35aaa;
  wire d35aab;
  wire d35aac;
  wire d35aad;
  wire d35aae;
  wire d35aaf;
  wire d35ab0;
  wire d35ab1;
  wire d35ab2;
  wire d35ab3;
  wire d35ab4;
  wire d35ab5;
  wire d35ab6;
  wire d35ab7;
  wire d35ab8;
  wire d35ab9;
  wire d35aba;
  wire d35abb;
  wire d35abc;
  wire d35abd;
  wire d35be2;
  wire d35be3;
  wire d35be4;
  wire d35be5;
  wire d35be6;
  wire d35be7;
  wire d35be8;
  wire d35be9;
  wire d35bea;
  wire d35beb;
  wire d35bec;
  wire d35bed;
  wire d35bee;
  wire d35bef;
  wire d35bf0;
  wire d35bf1;
  wire d35bf2;
  wire d35bf3;
  wire d35bf4;
  wire d35bf5;
  wire d35bf6;
  wire d35bf7;
  wire d35bf8;
  wire d35bf9;
  wire d35bfa;
  wire d35bfb;
  wire d35bfc;
  wire d35bfd;
  wire d35bfe;
  wire d35bff;
  wire d35c00;
  wire d35c01;
  wire d35c02;
  wire d35c03;
  wire d35c04;
  wire d35c05;
  wire d35c06;
  wire d35c07;
  wire d35c08;
  wire d35c09;
  wire d35c0a;
  wire d35c0b;
  wire d3540f;
  wire d35410;
  wire d35411;
  wire d35412;
  wire d35413;
  wire d35414;
  wire d35415;
  wire d35416;
  wire d35417;
  wire d35418;
  wire d35419;
  wire d3541a;
  wire d3541b;
  wire d3541c;
  wire d3541e;
  wire d3541f;
  wire d35420;
  wire d35421;
  wire d35422;
  wire d35423;
  wire d35424;
  wire d35425;
  wire d35426;
  wire d35427;
  wire d35428;
  wire d35429;
  wire d3542a;
  wire d3542b;
  wire d3542c;
  wire d3542d;
  wire d3542e;
  wire d3542f;
  wire d35430;
  wire d35431;
  wire d35432;
  wire d35433;
  wire d35434;
  wire d35435;
  wire d35436;
  wire d35437;
  wire d35438;
  wire d35439;
  wire d3543a;
  wire d3543b;
  wire d3543c;
  wire d3543d;
  wire d3543e;
  wire d3543f;
  wire d35440;
  wire d35441;
  wire d35442;
  wire d35443;
  wire d35444;
  wire d35445;
  wire d35492;
  wire d35493;
  wire d35494;
  wire d35495;
  wire d35496;
  wire d35497;
  wire d35498;
  wire d35499;
  wire d3549a;
  wire d3549b;
  wire d3549c;
  wire d3549d;
  wire d3549e;
  wire d3549f;
  wire d354a0;
  wire d354a1;
  wire d354a2;
  wire d354a3;
  wire d354a4;
  wire d354a5;
  wire d354a6;
  wire d354a7;
  wire d354a8;
  wire d354a9;
  wire d354aa;
  wire d354ab;
  wire d354ac;
  wire d354ad;
  wire d354ae;
  wire d354af;
  wire d354b0;
  wire d354b1;
  wire d354b2;
  wire d354b3;
  wire d354b4;
  wire d354b5;
  wire d354b6;
  wire d354b7;
  wire d354b8;
  wire d354b9;
  wire d354ba;
  wire d354bb;
  wire d354bc;
  wire d354bd;
  wire d354be;
  wire d354bf;
  wire d354c0;
  wire d354c1;
  wire d354c2;
  wire d354c3;
  wire d354c4;
  wire d354c5;
  wire d354c6;
  wire d354c7;
  wire d354c8;
  wire d354c9;
  wire d354ca;
  wire d354cb;
  wire d354cc;
  wire d354cd;
  wire d354ce;
  wire d354cf;
  wire d354d0;
  wire d354d1;
  wire d354d2;
  wire d354d3;
  wire d354d4;
  wire d354d5;
  wire d354d6;
  wire d354d7;
  wire d354d8;
  wire d354d9;
  wire d354da;
  wire d354db;
  wire d354dc;
  wire d354dd;
  wire d354de;
  wire d354df;
  wire d354e0;
  wire d354e1;
  wire d354e2;
  wire d354e3;
  wire d354e4;
  wire d354e5;
  wire d354e6;
  wire d354e7;
  wire d354e8;
  wire d354e9;
  wire d354ea;
  wire d354eb;
  wire d354ec;
  wire d354ed;
  wire d354ee;
  wire d354ef;
  wire d354f0;
  wire d354f1;
  wire d354f2;
  wire d354f3;
  wire d354f4;
  wire d354f5;
  wire d354f6;
  wire d354f7;
  wire d354f8;
  wire d354f9;
  wire d354fa;
  wire d354fb;
  wire d354fc;
  wire d354fd;
  wire d354fe;
  wire d354ff;
  wire d35500;
  wire d35501;
  wire d35502;
  wire d35503;
  wire d35504;
  wire d35505;
  wire d35506;
  wire d35507;
  wire d35508;
  wire d35509;
  wire d3550a;
  wire d3550b;
  wire d3550c;
  wire d3550d;
  wire d3550e;
  wire d3550f;
  wire d35510;
  wire d35511;
  wire d35512;
  wire d35513;
  wire d35514;
  wire d35515;
  wire d35516;
  wire d35517;
  wire d35518;
  wire d35519;
  wire d3551a;
  wire d3551b;
  wire d3551c;
  wire d3551d;
  wire d3551e;
  wire d3551f;
  wire d35520;
  wire d35521;
  wire d35522;
  wire d35523;
  wire d35524;
  wire d35525;
  wire d35526;
  wire d35527;
  wire d35528;
  wire d35529;
  wire d3552a;
  wire d3552b;
  wire d3552c;
  wire d3552d;
  wire d3552e;
  wire d3552f;
  wire d35565;
  wire d35566;
  wire d35567;
  wire d35568;
  wire d35569;
  wire d3556a;
  wire d3556b;
  wire d3556c;
  wire d3556d;
  wire d3556e;
  wire d3556f;
  wire d35570;
  wire d35571;
  wire d35572;
  wire d35573;
  wire d35574;
  wire d35575;
  wire d35576;
  wire d35577;
  wire d35578;
  wire d35579;
  wire d3557a;
  wire d3557b;
  wire d3557c;
  wire d3557d;
  wire d3557e;
  wire d3557f;
  wire d35580;
  wire d35581;
  wire d35582;
  wire d35583;
  wire d35584;
  wire d35585;
  wire d35586;
  wire d35587;
  wire d35588;
  wire d35589;
  wire d3558a;
  wire d3558b;
  wire d3558c;
  wire d3558d;
  wire d3558e;
  wire d3558f;
  wire d35590;
  wire d35591;
  wire d35592;
  wire d35593;
  wire d35594;
  wire d35595;
  wire d35596;
  wire d35597;
  wire d35598;
  wire d35599;
  wire d3559a;
  wire d3559b;
  wire d3559c;
  wire d3559d;
  wire d3559e;
  wire d3559f;
  wire d355a0;
  wire d355a1;
  wire d355a2;
  wire d355a3;
  wire d355a4;
  wire d355a5;
  wire d355a6;
  wire d355a7;
  wire d355a8;
  wire d355a9;
  wire d355aa;
  wire d355ab;
  wire d355ac;
  wire d355ad;
  wire d355ae;
  wire v845552;
  wire d355af;
  wire d355b0;
  wire d3560e;
  wire d35616;
  wire d35617;
  wire d35618;
  wire d35619;
  wire d3561a;
  wire d3561b;
  wire d3561c;
  wire d3561d;
  wire d3561e;
  wire d3561f;
  wire d35620;
  wire d35621;
  wire d35622;
  wire d35623;
  wire d35624;
  wire d35625;
  wire d35626;
  wire d35627;
  wire d35628;
  wire d35629;
  wire d3562a;
  wire d3562b;
  wire d3562c;
  wire d3562d;
  wire d3562e;
  wire d3562f;
  wire d35630;
  wire d35631;
  wire d35632;
  wire d35633;
  wire d3563b;
  wire d3563c;
  wire d3563d;
  wire d3563e;
  wire d3563f;
  wire d35640;
  wire d35641;
  wire d35642;
  wire d35643;
  wire d35644;
  wire d35645;
  wire d35646;
  wire d35647;
  wire d35648;
  wire d35649;
  wire d3564a;
  wire d3564b;
  wire d3564c;
  wire d3564d;
  wire d3564e;
  wire d3564f;
  wire d35650;
  wire d35651;
  wire d35652;
  wire d35653;
  wire d35654;
  wire d35655;
  wire d35656;
  wire d35657;
  wire d35658;
  wire d35659;
  wire d3565a;
  wire d3565b;
  wire d3565c;
  wire d3565d;
  wire d3565e;
  wire d35687;
  wire d35688;
  wire d35689;
  wire d3568a;
  wire d3568b;
  wire d3568c;
  wire d3568d;
  wire d3568e;
  wire d3568f;
  wire d35690;
  wire d35691;
  wire d35692;
  wire d35693;
  wire d35694;
  wire d35695;
  wire d35696;
  wire d35697;
  wire d35698;
  wire d35699;
  wire d3569a;
  wire d3569b;
  wire d3569c;
  wire d3569d;
  wire d3569e;
  wire d3569f;
  wire d356a0;
  wire d356a1;
  wire d356a2;
  wire d356a3;
  wire d356a4;
  wire d356a5;
  wire d356a6;
  wire d356a7;
  wire d356a8;
  wire d356a9;
  wire d356aa;
  wire d356ab;
  wire d356ac;
  wire d356ad;
  wire d356ae;
  wire d356af;
  wire d356b0;
  wire d356b1;
  wire d356b2;
  wire d356b3;
  wire d356b4;
  wire d356b5;
  wire d356b6;
  wire d356b7;
  wire d356b8;
  wire d356b9;
  wire d356ba;
  wire d356bb;
  wire d356bc;
  wire d356bd;
  wire d356be;
  wire d356bf;
  wire d356c0;
  wire d356c1;
  wire d356c2;
  wire d356c3;
  wire d356c4;
  wire d356c5;
  wire d356c6;
  wire d356c7;
  wire d356c8;
  wire d356c9;
  wire d356ca;
  wire d356cb;
  wire d356cc;
  wire d356cd;
  wire d356ce;
  wire d356cf;
  wire d356d0;
  wire d356d1;
  wire d356d2;
  wire d356d3;
  wire d356d4;
  wire d356d5;
  wire d356d6;
  wire d356d7;
  wire d356d8;
  wire d356d9;
  wire d356da;
  wire d356db;
  wire d356dc;
  wire d356dd;
  wire d356de;
  wire d356df;
  wire d356e0;
  wire d356e1;
  wire d356e2;
  wire d356e3;
  wire d356e4;
  wire d356e5;
  wire d356e6;
  wire d356e7;
  wire d356e8;
  wire d356e9;
  wire d356ea;
  wire d356eb;
  wire d356ec;
  wire d356ed;
  wire d356ee;
  wire d356ef;
  wire d356f0;
  wire d356f1;
  wire d356f2;
  wire d356f3;
  wire d356f4;
  wire d356f5;
  wire d356f6;
  wire d356f7;
  wire d356f8;
  wire d356f9;
  wire d356fa;
  wire d356fb;
  wire d356fc;
  wire d356fd;
  wire d356fe;
  wire d356ff;
  wire d35700;
  wire d35701;
  wire d35702;
  wire d35703;
  wire d35704;
  wire d35705;
  wire d35706;
  wire d35707;
  wire d35708;
  wire d35709;
  wire d3570a;
  wire d3570b;
  wire d3570c;
  wire d3570d;
  wire d3570e;
  wire d3570f;
  wire d35710;
  wire d35711;
  wire d35712;
  wire d35713;
  wire d35714;
  wire d35715;
  wire d35716;
  wire d35717;
  wire d35718;
  wire d35719;
  wire d3571a;
  wire d3571b;
  wire d3571c;
  wire d3571d;
  wire d3571e;
  wire d3571f;
  wire d35720;
  wire d35721;
  wire d35722;
  wire d35723;
  wire d35724;
  wire d35725;
  wire d35726;
  wire d35727;
  wire d35728;
  wire d35729;
  wire d3572a;
  wire d3572b;
  wire d3572c;
  wire d3572d;
  wire d3572e;
  wire d3572f;
  wire d35730;
  wire d35731;
  wire d35732;
  wire d35733;
  wire d35734;
  wire d35735;
  wire d35736;
  wire d35737;
  wire d35738;
  wire d35739;
  wire d3573a;
  wire d3573b;
  wire d3573c;
  wire d3573d;
  wire d3573e;
  wire d3573f;
  wire d35740;
  wire d35741;
  wire d35742;
  wire d35743;
  wire d35744;
  wire d35745;
  wire d35746;
  wire d35747;
  wire d35748;
  wire d35749;
  wire d3574a;
  wire d3574b;
  wire d3574c;
  wire d3574d;
  wire d3574e;
  wire d3574f;
  wire d35750;
  wire d35751;
  wire d35752;
  wire d35753;
  wire d35754;
  wire d35755;
  wire d35756;
  wire d35757;
  wire d35758;
  wire d35759;
  wire d3575a;
  wire d3575b;
  wire d3575c;
  wire d3575d;
  wire d3575e;
  wire d3575f;
  wire d35760;
  wire d35761;
  wire d35762;
  wire d35763;
  wire d35764;
  wire d35765;
  wire d35766;
  wire d35767;
  wire d35768;
  wire d35769;
  wire d3576a;
  wire d3576b;
  wire d3576e;
  wire d3576f;
  wire d35770;
  wire d35771;
  wire d35774;
  wire d35775;
  wire d35776;
  wire d35777;
  wire d35778;
  wire d35779;
  wire d3577a;
  wire d3577b;
  wire d3577c;
  wire d3577d;
  wire d3577e;
  wire d3577f;
  wire d3578a;
  wire d3578b;
  wire d3578c;
  wire d3578d;
  wire d3578e;
  wire d3578f;
  wire d35790;
  wire d35791;
  wire d35792;
  wire d35793;
  wire d35794;
  wire d35795;
  wire d35796;
  wire d35797;
  wire d35798;
  wire d35799;
  wire d3579a;
  wire d3579b;
  wire d3579c;
  wire d3579d;
  wire d3579e;
  wire d3579f;
  wire d357a0;
  wire d357a1;
  wire d357a2;
  wire d357a3;
  wire d357a4;
  wire d357a5;
  wire d357a6;
  wire d357a7;
  wire d357a8;
  wire d357a9;
  wire d357aa;
  wire d357ab;
  wire d357ac;
  wire d357ad;
  wire d357ae;
  wire d357af;
  wire d357b0;
  wire d357b1;
  wire d357b2;
  wire d357b3;
  wire d357b6;
  wire d357b7;
  wire d357b8;
  wire d357b9;
  wire d357ba;
  wire d357bb;
  wire d357bc;
  wire d357bd;
  wire d357be;
  wire d357bf;
  wire d357c0;
  wire d357c1;
  wire d357c2;
  wire d357c3;
  wire d357c4;
  wire d357c5;
  wire d357c6;
  wire d357c8;
  wire d357c9;
  wire d357ca;
  wire d357cb;
  wire d357cc;
  wire d357cd;
  wire d357ce;
  wire d357cf;
  wire d357d0;
  wire d357d1;
  wire d357d3;
  wire d357d4;
  wire d357d5;
  wire d357d6;
  wire d357d7;
  wire d357da;
  wire d357db;
  wire d357dc;
  wire d357dd;
  wire d357de;
  wire d357df;
  wire d357e0;
  wire d357e1;
  wire d357e2;
  wire d357e3;
  wire d357e4;
  wire d357e7;
  wire d357e8;
  wire d357e9;
  wire d357ea;
  wire d357eb;
  wire d357ec;
  wire d357ed;
  wire d357ee;
  wire d357ef;
  wire d357f0;
  wire d357f1;
  wire d357f2;
  wire d357f3;
  wire d357f4;
  wire d357f5;
  wire d357f6;
  wire d357f7;
  wire d357f8;
  wire d357f9;
  wire d357fa;
  wire d357fb;
  wire d357fc;
  wire d357fd;
  wire d357fe;
  wire d357ff;
  wire d35800;
  wire d35801;
  wire d35802;
  wire d35803;
  wire d35804;
  wire d35805;
  wire d35806;
  wire d35807;
  wire d35808;
  wire d35809;
  wire d3580a;
  wire d3580b;
  wire d3580c;
  wire d3500f;
  wire d35010;
  wire d35011;
  wire d35012;
  wire d35013;
  wire d35014;
  wire d35015;
  wire d35016;
  wire d35017;
  wire d35018;
  wire d35019;
  wire d3501a;
  wire d3501b;
  wire d3501c;
  wire d3501d;
  wire d3501e;
  wire d3501f;
  wire d35020;
  wire d35021;
  wire d35022;
  wire d35023;
  wire d35024;
  wire d35025;
  wire d35026;
  wire d35027;
  wire d35028;
  wire cc36b8;
  wire cc36b9;
  wire cc36ba;
  wire cc36bb;
  wire cc36bc;
  wire cc36bd;
  wire cc36be;
  wire cc36bf;
  wire cc36c0;
  wire cc36c1;
  wire cc36c2;
  wire cc36c3;
  wire cc36c4;
  wire cc36c5;
  wire cc36c6;
  wire cc36c7;
  wire cc36c8;
  wire cc36c9;
  wire cc36ca;
  wire cc36cb;
  wire cc36cc;
  wire cc36cd;
  wire cc36ce;
  wire cc36cf;
  wire cc36d0;
  wire cc36d1;
  wire cc36d2;
  wire cc36d3;
  wire cc36d4;
  wire cc36d5;
  wire cc36d6;
  wire cc36d7;
  wire cc36d8;
  wire cc36d9;
  wire cc36da;
  wire cc36db;
  wire cc36dc;
  wire cc36dd;
  wire cc36de;
  wire cc36df;
  wire cc36e0;
  wire cc36e1;
  wire cc36e2;
  wire cc36e3;
  wire cc36e4;
  wire cc36e5;
  wire cc36e6;
  wire cc36e7;
  wire cc36e8;
  wire cc36e9;
  wire cc36ea;
  wire cc36eb;
  wire cc36ec;
  wire cc36ed;
  wire cc36ee;
  wire cc36ef;
  wire cc36f0;
  wire cc36f1;
  wire cc36f2;
  wire cc36f3;
  wire cc36f4;
  wire cc36f5;
  wire cc36f6;
  wire cc36f7;
  wire cc36f8;
  wire cc36f9;
  wire cc36fa;
  wire cc36fb;
  wire cc36fc;
  wire cc36fd;
  wire cc36fe;
  wire cc36ff;
  wire cc3700;
  wire cc3701;
  wire cc3702;
  wire cc3703;
  wire cc3704;
  wire cc3705;
  wire cc3706;
  wire cc3707;
  wire cc3708;
  wire cc3709;
  wire cc370a;
  wire cc370b;
  wire v845555;
  wire v84557c;
  wire c3d2ad;
  wire c3d2ae;
  wire c3d2af;
  wire c3d2b0;
  wire c3d2b1;
  wire c3d2b2;
  wire c3d2b3;
  wire c3d2b4;
  wire c3d2b5;
  wire c3d2b6;
  wire c3d2b7;
  wire c3d2b8;
  wire c3d2b9;
  wire c3d2ba;
  wire v84554d;
  wire c3d2bb;
  wire c3d2bc;
  wire c3d2bd;
  wire c3d2be;
  wire c3d2bf;
  wire c3d2c0;
  wire c3d2c4;
  wire c3d2c5;
  wire c3d2c6;
  wire c3d2c7;
  wire c3d2c8;
  wire c3d2c9;
  wire c3d2ca;
  wire c3d2cb;
  wire c3d2cc;
  wire c3d2cd;
  wire c3d2ce;
  wire c3d2cf;
  wire c3d2d0;
  wire c3d2d1;
  wire c3d2d2;
  wire c3d2d5;
  wire c3d2d6;
  wire c3d2d7;
  wire c3d2d8;
  wire c3d2d9;
  wire c3d2da;
  wire c3d2db;
  wire c3d2dc;
  wire c3d2dd;
  wire c3d2de;
  wire c3d2df;
  wire c3d2e0;
  wire c3d2e1;
  wire c3d2e2;
  wire c3d2e3;
  wire v845551;
  wire c3d2e5;
  wire c3d2e6;
  wire c3d2e7;
  wire c3d2e8;
  wire c3d2e9;
  wire c3d2ea;
  wire c3d2eb;
  wire c3d2ec;
  wire c3d2ed;
  wire c3d2ee;
  wire c3d2ef;
  wire c3d2f0;
  wire c3d2f1;
  wire c3d2f2;
  wire c3d2f3;
  wire c3d2f4;
  wire c3d2f5;
  wire c3d2f6;
  wire c3d2f7;
  wire c3d2f8;
  wire c3d2f9;
  wire c3d2fa;
  wire c3d2fb;
  wire c3d2fc;
  wire c3d2fd;
  wire c3d2fe;
  wire c3d2ff;
  wire c3d300;
  wire c3d301;
  wire c3d302;
  wire c3d303;
  wire c3d304;
  wire c3d305;
  wire c3d306;
  wire c3d307;
  wire c3d308;
  wire c3d309;
  wire c3d30a;
  wire c3d30b;
  wire c3d30c;
  wire c3d30d;
  wire c3d30e;
  wire c3d30f;
  wire c3d310;
  wire c3d311;
  wire c3d312;
  wire c3d313;
  wire c3d314;
  wire c3d315;
  wire c3d316;
  wire c3d317;
  wire c3d318;
  wire c3d319;
  wire c3d31a;
  wire c3d31b;
  wire c3d31c;
  wire c3d31d;
  wire c3d31e;
  wire c3d31f;
  wire c3d320;
  wire c3d321;
  wire c3d322;
  wire c3d323;
  wire c3d324;
  wire c3d325;
  wire c3d326;
  wire c3d327;
  wire c3d328;
  wire c3d329;
  wire c3d32a;
  wire c3d32b;
  wire c3d32c;
  wire c3d32d;
  wire c3d32e;
  wire c3d32f;
  wire c3d330;
  wire c3d331;
  wire c3d332;
  wire c3d333;
  wire c3d336;
  wire c3d337;
  wire c3d338;
  wire c3d339;
  wire c3d33a;
  wire c3d33b;
  wire c3d33c;
  wire c3d33d;
  wire c3d33e;
  wire c3d33f;
  wire c3d340;
  wire c3d341;
  wire c3d342;
  wire c3d343;
  wire c3d344;
  wire c3d345;
  wire c3d346;
  wire c3d347;
  wire c3d348;
  wire c3d349;
  wire c3d34a;
  wire c3d34b;
  wire c3d34c;
  wire c3d34d;
  wire c3d34e;
  wire c3d34f;
  wire c3d350;
  wire c3d351;
  wire c3d352;
  wire c3d353;
  wire c3d354;
  wire c3d355;
  wire c3d356;
  wire c3d357;
  wire c3d359;
  wire c3d35b;
  wire c3d35c;
  wire c3d35d;
  wire c3d35e;
  wire c3d35f;
  wire c3d360;
  wire c3d361;
  wire c3d362;
  wire c3d364;
  wire c3d368;
  wire c3d369;
  wire c3d36a;
  wire c3d36b;
  wire c3d36c;
  wire c3d36e;
  wire c3d36f;
  wire c3d370;
  wire c3d371;
  wire c3d372;
  wire c3d373;
  wire c3d374;
  wire c3d375;
  wire c3d376;
  wire c3d377;
  wire c3d378;
  wire c3d379;
  wire c3d37a;
  wire c3d37b;
  wire c3d37c;
  wire c3d37d;
  wire c3d37e;
  wire c3d37f;
  wire c3d380;
  wire c3d381;
  wire c3d382;
  wire c3d383;
  wire c3d385;
  wire c3d386;
  wire c3d387;
  wire c3d388;
  wire c3d389;
  wire c3d38a;
  wire c3d38b;
  wire c3d38c;
  wire c3d38d;
  wire c3d38e;
  wire c3d38f;
  wire c3d390;
  wire c3d391;
  wire c3d392;
  wire c3d393;
  wire c3d394;
  wire c3d395;
  wire c3d396;
  wire c3d397;
  wire c3d398;
  wire c3d399;
  wire c3d39a;
  wire c3d39b;
  wire c3d39c;
  wire c3d39d;
  wire c3d39e;
  wire c3d39f;
  wire c3d3a0;
  wire c3d3a1;
  wire c3d3a2;
  wire c3d3a3;
  wire c3d3a4;
  wire c3d3a5;
  wire c3d3a6;
  wire c3d3a7;
  wire c3d3a8;
  wire c3d3a9;
  wire c3d3aa;
  wire c3d3ab;
  wire c3d3ac;
  wire c3d3ad;
  wire c3d478;
  wire c3d479;
  wire c3d47a;
  wire c3d47b;
  wire c3d47c;
  wire c3d47d;
  wire c3d47e;
  wire c3d47f;
  wire c3d480;
  wire c3d481;
  wire c3d482;
  wire c3d483;
  wire c3d484;
  wire c3d4db;
  wire c3d4dc;
  wire c3d4dd;
  wire c3d4de;
  wire c3d4df;
  wire c3d4e0;
  wire c3d4e1;
  wire c3d4e2;
  wire c3d4e3;
  wire c3d4f0;
  wire c3d4f1;
  wire c3d4f2;
  wire c3d4f3;
  wire c3d4f4;
  wire c3d4f5;
  wire c3d4f6;
  wire c3d4f7;
  wire c3d4f8;
  wire c3d4f9;
  wire c3d4fa;
  wire c3d4fb;
  wire c3d4fc;
  wire c3d4fd;
  wire c3d4fe;
  wire c3d4ff;
  wire c3d500;
  wire c3d501;
  wire c3d502;
  wire c3d503;
  wire c3d504;
  wire c3d505;
  wire c3d506;
  wire c3d507;
  wire c3d508;
  wire c3d509;
  wire c3d50a;
  wire c3d50b;
  wire c3d50c;
  wire c3d50d;
  wire c3d50e;
  wire c3d50f;
  wire c3d510;
  wire c3d511;
  wire c3d512;
  wire c3d513;
  wire c3d514;
  wire c3d515;
  wire c3d516;
  wire c3d517;
  wire c3d518;
  wire c3d519;
  wire c3d51a;
  wire c3d51b;
  wire c3d51c;
  wire c3d51d;
  wire c3d51e;
  wire c3d51f;
  wire c3d520;
  wire c3d521;
  wire c3d522;
  wire c3d523;
  wire c3d524;
  wire c3d525;
  wire c3d526;
  wire c3d527;
  wire c3d528;
  wire c3d529;
  wire c3d52a;
  wire c3d52b;
  wire c3d52c;
  wire c3d52d;
  wire c3d52e;
  wire c3d52f;
  wire c3d530;
  wire c3d531;
  wire c3d532;
  wire c3d533;
  wire c3d534;
  wire c3d535;
  wire c3d578;
  wire c3d579;
  wire c3d57a;
  wire c3d57b;
  wire c3d57c;
  wire c3d57d;
  wire c3d57e;
  wire c3d57f;
  wire c3d580;
  wire c3d581;
  wire c3d582;
  wire c3d583;
  wire c3d584;
  wire c3d585;
  wire c3d586;
  wire c3d587;
  wire c3d588;
  wire c3d589;
  wire c3d58a;
  wire c3d58e;
  wire c3d58f;
  wire c3d590;
  wire c3d591;
  wire c3d592;
  wire c3d594;
  wire c3d595;
  wire c3d596;
  wire c3d597;
  wire c3d598;
  wire c3d599;
  wire c3d59a;
  wire c3d59d;
  wire c3d59e;
  wire c3d59f;
  wire c3d5a0;
  wire c3d5a1;
  wire c3d5a2;
  wire c3d5a3;
  wire c3d5a6;
  wire c3d5a7;
  wire c3d5a8;
  wire c3d5a9;
  wire c3d5aa;
  wire c3d5ab;
  wire c3d5ac;
  wire c3d5ad;
  wire c3d5ae;
  wire c3d5af;
  wire c3d5b0;
  wire c3d5b1;
  wire c3d5b2;
  wire c3d5b3;
  wire c3d5b4;
  wire c3d5b5;
  wire c3d5b6;
  wire c3d5b7;
  wire c3d5b8;
  wire c3d5b9;
  wire c3d5ba;
  wire c3d5bb;
  wire c3d5bc;
  wire c3d5bd;
  wire c3d5be;
  wire c3d5bf;
  wire c3d5c0;
  wire c3d5c1;
  wire c3d5c2;
  wire c3d5c3;
  wire c3d5c4;
  wire c3d5c5;
  wire c3d5c6;
  wire c3d5c7;
  wire c3d5c8;
  wire c3d5c9;
  wire c3d5ca;
  wire c3d5cb;
  wire c3d5cc;
  wire c3d5cd;
  wire c3d5ce;
  wire c3d5cf;
  wire c3d5d0;
  wire c3d5d1;
  wire c3d5d2;
  wire c3d5d3;
  wire c3d5d4;
  wire c3d5d5;
  wire c3d5d6;
  wire c3d5d7;
  wire c3d5d8;
  wire c3d5d9;
  wire c3d5da;
  wire c3d5db;
  wire c3d5dc;
  wire c3d5dd;
  wire c3d5de;
  wire c3d5df;
  wire c3d5e0;
  wire c3d5e1;
  wire c3d5e2;
  wire c3d5e3;
  wire c3d5e4;
  wire c3d5e5;
  wire c3d5e6;
  wire c3d5e7;
  wire c3d5e8;
  wire c3d5e9;
  wire c3d5ea;
  wire c3d5eb;
  wire c3d5ec;
  wire c3d5ed;
  wire c3d5ee;
  wire c3d5ef;
  wire c3d5f0;
  wire c3d5f1;
  wire c3d5f2;
  wire c3d5f3;
  wire c3d5f4;
  wire c3d5f5;
  wire c3cdf9;
  wire c3cdfa;
  wire c3cdfb;
  wire c3cdfc;
  wire c3cdfd;
  wire c3cdfe;
  wire c3cdff;
  wire c3ce00;
  wire c3ce01;
  wire c3ce02;
  wire c3ce03;
  wire c3ce04;
  wire c3ce05;
  wire c3ce06;
  wire c3ce07;
  wire c3ce08;
  wire c3ce09;
  wire c3ce0a;
  wire c3ce13;
  wire c3ce14;
  wire c3ce15;
  wire c3ce16;
  wire c3ce17;
  wire c3ce18;
  wire c3ce19;
  wire c3ce1a;
  wire c3ce1b;
  wire c3ce1c;
  wire c3ce1d;
  wire c3ce1e;
  wire c3ce1f;
  wire c3ce20;
  wire c3ce21;
  wire c3ce22;
  wire c3ce23;
  wire c3ce24;
  wire c3ce25;
  wire c3ce26;
  wire c3ce27;
  wire c3ce28;
  wire c3ce29;
  wire c3ce2a;
  wire c3ce2b;
  wire c3ce2c;
  wire c3ce2d;
  wire c3ce2e;
  wire c3ce2f;
  wire c3ce30;
  wire c3ce31;
  wire c3ce32;
  wire c3ce33;
  wire c3ce34;
  wire c3ce35;
  wire c3ce36;
  wire c3ce37;
  wire c3ce38;
  wire c3ce39;
  wire c3ce3a;
  wire c3ce3b;
  wire c3ce3c;
  wire c3ce3d;
  wire c3ce3e;
  wire c3ce3f;
  wire c3ce40;
  wire c3ce41;
  wire c3ce42;
  wire c3ce43;
  wire c3ce44;
  wire c3ce45;
  wire c3ce46;
  wire c3ce47;
  wire c3ce48;
  wire c3ce49;
  wire c3ce4a;
  wire c3ce4b;
  wire c3ce4c;
  wire c3ce4d;
  wire c3ce4e;
  wire c3ce4f;
  wire c3ce50;
  wire c3ce51;
  wire c3ce52;
  wire c3ce53;
  wire c3ce54;
  wire c3ce55;
  wire c3ce56;
  wire c3ce57;
  wire c3ce58;
  wire c3ce59;
  wire c3ce5a;
  wire c3ce5b;
  wire c3ce5c;
  wire c3ce5d;
  wire c3ce5e;
  wire c3ce5f;
  wire c3ce60;
  wire c3ce61;
  wire c3ce62;
  wire c3ce63;
  wire c3ce64;
  wire c3ce65;
  wire c3ce66;
  wire c3ce67;
  wire c3ce68;
  wire c3ce69;
  wire c3ce6a;
  wire c3ce6b;
  wire c3ce6c;
  wire c3ce6d;
  wire c3ce6e;
  wire c3ce6f;
  wire c3ce70;
  wire c3ce71;
  wire c3ce72;
  wire c3ce73;
  wire c3ce74;
  wire c3ce75;
  wire c3ce76;
  wire c3ce77;
  wire c3ce78;
  wire c3ce79;
  wire c3ce7a;
  wire c3ce7b;
  wire c3ce7c;
  wire c3ce7d;
  wire c3ce7e;
  wire c3ce7f;
  wire c3ce80;
  wire c3ce81;
  wire c3ce82;
  wire c3ce83;
  wire c3ce84;
  wire c3ce85;
  wire c3ce86;
  wire c3ce87;
  wire c3ce88;
  wire c3ce89;
  wire c3ce8a;
  wire c3ce8b;
  wire c3ce8c;
  wire c3ce8d;
  wire c3ce8e;
  wire c3ce8f;
  wire c3ce90;
  wire c3ce91;
  wire c3ce92;
  wire c3ce93;
  wire c3ce94;
  wire c3ce95;
  wire c3ce96;
  wire c3ce97;
  wire c3ce98;
  wire c3ce99;
  wire c3ce9a;
  wire c3ce9b;
  wire c3ce9c;
  wire c3ce9d;
  wire c3ce9e;
  wire c3ce9f;
  wire c3cea0;
  wire c3cea1;
  wire c3cea2;
  wire c3cea3;
  wire c3cea4;
  wire c3cea5;
  wire c3cea6;
  wire c3cea7;
  wire c3cea8;
  wire c3cea9;
  wire c3ceaa;
  wire c3ceab;
  wire c3ceac;
  wire c3cead;
  wire c3ceae;
  wire c3ceaf;
  wire c3ceb0;
  wire c3ceb1;
  wire c3ceb2;
  wire c3ceb3;
  wire c3ceb4;
  wire c3ceb5;
  wire c3ceb6;
  wire c3ceb7;
  wire c3ceb8;
  wire c3ceb9;
  wire c3ceba;
  wire c3cebb;
  wire c3cebc;
  wire c3cebd;
  wire c3cebe;
  wire c3cebf;
  wire c3cec0;
  wire c3cec2;
  wire c3cec3;
  wire c3cec4;
  wire c3cec5;
  wire c3cec6;
  wire c3cec7;
  wire c3cec8;
  wire c3cec9;
  wire c3ceca;
  wire c3cecb;
  wire c3cecc;
  wire c3cecd;
  wire c3cece;
  wire c3cecf;
  wire c3ced0;
  wire c3ced1;
  wire c3ced2;
  wire c3ced3;
  wire c3ced4;
  wire c3ced5;
  wire c3ced6;
  wire c3ced7;
  wire c3ced8;
  wire c3ced9;
  wire c3ceda;
  wire c3cedb;
  wire c3cedc;
  wire c3cedd;
  wire c3cede;
  wire c3cedf;
  wire c3cee0;
  wire c3cee1;
  wire c3cee2;
  wire c3cee3;
  wire c3cee4;
  wire c3cee5;
  wire c3cee6;
  wire c3cee7;
  wire c3cee8;
  wire c3cee9;
  wire c3ceea;
  wire c3ceeb;
  wire c3ceec;
  wire c3ceed;
  wire c3ceee;
  wire c3ceef;
  wire c3cef0;
  wire c3cef1;
  wire c3cef2;
  wire c3cef3;
  wire c3cef4;
  wire c3cef5;
  wire c3cef6;
  wire c3cef7;
  wire c3cef8;
  wire c3cef9;
  wire c3cefa;
  wire c3cefb;
  wire c3cefc;
  wire c3cefd;
  wire c3cefe;
  wire c3ceff;
  wire c3cf00;
  wire c3cf01;
  wire c3cf02;
  wire c3cf03;
  wire c3cf04;
  wire c3cf05;
  wire c3cf06;
  wire c3cf07;
  wire c3cf08;
  wire c3cf09;
  wire c3cf0a;
  wire c3cf0b;
  wire c3cf0c;
  wire c3cf0d;
  wire c3cf0e;
  wire c3cf0f;
  wire c3cf10;
  wire c3cf11;
  wire c3cf12;
  wire c3cf13;
  wire c3cf14;
  wire c3cf15;
  wire c3cf16;
  wire c3cf17;
  wire c3cf18;
  wire c3cf19;
  wire c3cf1a;
  wire c3cf1b;
  wire c3cf1c;
  wire c3cf1d;
  wire c3cf1e;
  wire c3cf1f;
  wire c3cf20;
  wire c3cf21;
  wire c3cf22;
  wire c3cf23;
  wire c3cf24;
  wire c3cf25;
  wire c3cf26;
  wire c3cf27;
  wire c3cf28;
  wire c3cf29;
  wire c3cf2a;
  wire c3cf2b;
  wire c3cf2c;
  wire c3cf2d;
  wire c3cf2e;
  wire c3cf2f;
  wire c3cf30;
  wire c3cf31;
  wire c3cf32;
  wire c3cf33;
  wire c3cf34;
  wire bd5b69;
  wire bd5b6a;
  wire bd5b6b;
  wire bd5b6c;
  wire bd5b6d;
  wire bd5b6e;
  wire bd5b6f;
  wire bd5b70;
  wire bd5b71;
  wire bd5b72;
  wire bd5b73;
  wire bd5b74;
  wire bd5b75;
  wire bd5b77;
  wire bd5b78;
  wire bd5b79;
  wire bd5b7a;
  wire bd5b7b;
  wire bd5b7c;
  wire bd5b7d;
  wire bd5b7e;
  wire bd5b7f;
  wire bd5b80;
  wire bd5b81;
  wire bd5b82;
  wire bd5b83;
  wire bd5b84;
  wire bd5b85;
  wire bd5b86;
  wire bd5b87;
  wire bd5b88;
  wire bd5b89;
  wire bd5b8a;
  wire bd5b8b;
  wire bd5b8c;
  wire bd5b8d;
  wire bd5b8e;
  wire bd5b8f;
  wire bd5b90;
  wire bd5b91;
  wire bd5b92;
  wire bd5b93;
  wire bd5b94;
  wire bd5b95;
  wire bd5b96;
  wire bd5b97;
  wire bd5b98;
  wire bd5b99;
  wire bd5b9a;
  wire bd5b9b;
  wire bd5b9c;
  wire bd5b9d;
  wire bd5b9f;
  wire bd5ba0;
  wire bd5ba1;
  wire bd5ba2;
  wire bd5ba3;
  wire bd5ba4;
  wire bd5ba5;
  wire bd5ba6;
  wire bd5ba7;
  wire bd5ba8;
  wire bd5ba9;
  wire bd5baa;
  wire bd5bab;
  wire bd5bac;
  wire bd5bad;
  wire bd5bae;
  wire bd5baf;
  wire bd5bb0;
  wire bd5bb1;
  wire bd5bb2;
  wire bd5bb3;
  wire bd5e1b;
  wire bd5e1c;
  wire bd5e1d;
  wire bd5e1e;
  wire bd5e1f;
  wire bd5e20;
  wire bd5e21;
  wire bd5e22;
  wire bd5e25;
  wire bd5e26;
  wire bd5e29;
  wire bd5e99;
  wire bd5e9a;
  wire bd5e9b;
  wire bd5e9c;
  wire bd5e9d;
  wire bd5e9e;
  wire bd5e9f;
  wire bd5ea0;
  wire bd5ea1;
  wire bd5ea2;
  wire bd5ea3;
  wire bd5ea4;
  wire bd5ea5;
  wire bd5ea6;
  wire bd5ea7;
  wire bd5ea8;
  wire bd5ea9;
  wire bd56cb;
  wire bd56cc;
  wire bd56cd;
  wire bd56ce;
  wire bd56cf;
  wire bd56d0;
  wire bd56d1;
  wire bd56d2;
  wire bd56d3;
  wire bd56d4;
  wire bd56d5;
  wire bd56d6;
  wire bd56d7;
  wire bd56d8;
  wire bd56d9;
  wire bd56da;
  wire bd56db;
  wire bd56dc;
  wire bd56dd;
  wire bd56de;
  wire bd56df;
  wire bd56e0;
  wire bd5728;
  wire bd572c;
  wire bd572e;
  wire bd572f;
  wire bd5733;
  wire bd5735;
  wire bd5736;
  wire bd5737;
  wire bd5738;
  wire bd5739;
  wire bd573d;
  wire bd573f;
  wire bd5740;
  wire bd5744;
  wire bd5746;
  wire bd5747;
  wire bd5748;
  wire bd5749;
  wire bd574a;
  wire bd574b;
  wire bd574c;
  wire bd574d;
  wire bd574e;
  wire bd574f;
  wire bd5750;
  wire bd5752;
  wire bd5754;
  wire bd5755;
  wire bd5756;
  wire bd5757;
  wire bd5758;
  wire bd5759;
  wire bd575a;
  wire bd575b;
  wire bd575c;
  wire bd575d;
  wire bd575e;
  wire bd575f;
  wire bd5760;
  wire bd5761;
  wire bd5762;
  wire bd5765;
  wire bd5766;
  wire bd5767;
  wire bd5768;
  wire bd5769;
  wire bd576a;
  wire bd576b;
  wire bd576c;
  wire bd576d;
  wire bd576e;
  wire bd5771;
  wire bd5772;
  wire bd5773;
  wire bd5774;
  wire bd5775;
  wire bd5776;
  wire bd5777;
  wire bd5778;
  wire bd5779;
  wire bd577a;
  wire bd577b;
  wire bd577e;
  wire bd577f;
  wire bd5780;
  wire bd5781;
  wire bd5782;
  wire bd5783;
  wire bd5784;
  wire bd5785;
  wire bd5786;
  wire bd5787;
  wire bd5788;
  wire bd5789;
  wire bd578a;
  wire bd578b;
  wire bd578c;
  wire bd578d;
  wire bd578e;
  wire bd578f;
  wire bd5790;
  wire bd5791;
  wire bd5792;
  wire bd5793;
  wire bd5794;
  wire bd5795;
  wire bd5796;
  wire bd5797;
  wire bd5798;
  wire bd5799;
  wire bd579a;
  wire bd579b;
  wire bd579c;
  wire bd579d;
  wire bd579e;
  wire bd579f;
  wire bd57a0;
  wire bd57a1;
  wire bd57a2;
  wire bd57ae;
  wire bd57af;
  wire bd57b0;
  wire bd57b1;
  wire bd57b2;
  wire bd57ba;
  wire bd57bb;
  wire bd57bc;
  wire bd57bd;
  wire bd57be;
  wire bd57bf;
  wire bd57c0;
  wire bd57c1;
  wire bd57c2;
  wire bd57c3;
  wire bd57c4;
  wire bd57c5;
  wire bd57c7;
  wire bd57c8;
  wire bd57c9;
  wire bd57ca;
  wire bd57cb;
  wire bd57cc;
  wire bd57cd;
  wire bd57ce;
  wire bd57cf;
  wire bd57d0;
  wire bd57d1;
  wire bd57d2;
  wire bd57de;
  wire bd57df;
  wire bd57e0;
  wire bd57e1;
  wire bd57e2;
  wire bd57e3;
  wire bd57e4;
  wire bd57e5;
  wire bd57e6;
  wire bd57e7;
  wire bd57e8;
  wire bd57e9;
  wire bd57ea;
  wire bd57eb;
  wire bd57ec;
  wire bd57ed;
  wire bd57ee;
  wire bd57ef;
  wire bd57f0;
  wire bd57f1;
  wire bd57f2;
  wire bd57f3;
  wire bd57f4;
  wire bd57f5;
  wire bd57f6;
  wire bd57f7;
  wire bd57f8;
  wire bd57f9;
  wire bd57fa;
  wire bd57fb;
  wire bd57fc;
  wire bd57fd;
  wire bd57fe;
  wire bd57ff;
  wire bd5800;
  wire bd5801;
  wire bd5802;
  wire bd5803;
  wire bd5804;
  wire bd5805;
  wire bd5806;
  wire bd5807;
  wire bd5808;
  wire bd5809;
  wire bd580a;
  wire bd580b;
  wire bd580c;
  wire bd580d;
  wire bd580e;
  wire bd580f;
  wire bd5810;
  wire bd5811;
  wire bd5812;
  wire bd5813;
  wire bd5814;
  wire bd5815;
  wire bd5816;
  wire bd5817;
  wire bd5818;
  wire bd5819;
  wire bd581a;
  wire bd581b;
  wire bd581c;
  wire bd581d;
  wire bd581e;
  wire bd581f;
  wire bd5820;
  wire bd5821;
  wire bd5822;
  wire bd5823;
  wire bd5824;
  wire bd5825;
  wire bd5826;
  wire bd5827;
  wire bd5828;
  wire bd5829;
  wire bd582a;
  wire bd582b;
  wire bd582c;
  wire bd582d;
  wire bd582e;
  wire bd582f;
  wire bd5830;
  wire bd5831;
  wire bd5832;
  wire bd5833;
  wire bd5834;
  wire bd5835;
  wire bd5836;
  wire bd5837;
  wire bd5838;
  wire bd5839;
  wire bd583a;
  wire bd583b;
  wire bd583c;
  wire bd583d;
  wire bd583e;
  wire bd583f;
  wire bd5840;
  wire bd5841;
  wire bd5842;
  wire bd5843;
  wire bd5844;
  wire bd5845;
  wire bd5846;
  wire bd5847;
  wire bd5848;
  wire bd5849;
  wire bd584a;
  wire bd584b;
  wire bd584c;
  wire bd584d;
  wire bd584e;
  wire bd584f;
  wire bd5850;
  wire bd5851;
  wire bd5852;
  wire bd5853;
  wire bd5854;
  wire bd5855;
  wire bd5856;
  wire bd5857;
  wire bd5858;
  wire bd5859;
  wire bd585a;
  wire bd585b;
  wire bd585c;
  wire bd585d;
  wire bd585e;
  wire bd585f;
  wire bd5860;
  wire bd5861;
  wire bd5862;
  wire bd5863;
  wire bd5864;
  wire bd5865;
  wire bd5866;
  wire bd5867;
  wire bd5868;
  wire bd5869;
  wire bd586a;
  wire bd586b;
  wire bd586c;
  wire bd586d;
  wire bd586e;
  wire bd586f;
  wire bd5870;
  wire bd5871;
  wire bd5872;
  wire bd5873;
  wire bd5874;
  wire bd5875;
  wire bd5876;
  wire bd5877;
  wire bd5878;
  wire bd5879;
  wire bd587a;
  wire bd587b;
  wire bd587c;
  wire bd587d;
  wire bd587e;
  wire bd587f;
  wire bd5880;
  wire bd5881;
  wire bd5882;
  wire bd5883;
  wire bd5884;
  wire bd5885;
  wire bd5886;
  wire bd5887;
  wire bd5888;
  wire bd5889;
  wire bd588a;
  wire bd588b;
  wire bd588c;
  wire bd588d;
  wire bd588e;
  wire bd588f;
  wire bd5890;
  wire bd5891;
  wire bd5892;
  wire bd5893;
  wire bd5894;
  wire bd5895;
  wire bd5896;
  wire bd5897;
  wire bd5898;
  wire bd5899;
  wire bd589a;
  wire bd589b;
  wire bd589c;
  wire bd589d;
  wire bd589e;
  wire bd589f;
  wire bd58a0;
  wire bd58a1;
  wire bd58a2;
  wire bd58a3;
  wire bd58a4;
  wire bd58a5;
  wire bd58a6;
  wire bd58a7;
  wire bd58a8;
  wire bd58a9;
  wire bd58aa;
  wire bd58ab;
  wire bd58ac;
  wire bd58ad;
  wire bd58ae;
  wire bd58af;
  wire bd58b0;
  wire bd58b1;
  wire bd58b2;
  wire bd58b3;
  wire bd58b4;
  wire bd58b5;
  wire bd58b6;
  wire bd58b7;
  wire bd58b8;
  wire bd58b9;
  wire bd58ba;
  wire bd58bb;
  wire bd58bc;
  wire bd58bd;
  wire bd58be;
  wire bd58bf;
  wire bd58c0;
  wire bd58c1;
  wire bd58c2;
  wire bd58c3;
  wire bd58c4;
  wire bd58c5;
  wire bd58c6;
  wire bd58c7;
  wire bd58c8;
  wire bd58c9;
  wire bd58ca;
  wire bd58cb;
  wire bd58cc;
  wire bd58cd;
  wire bd58ce;
  wire bd58cf;
  wire bd58d0;
  wire bd58d1;
  wire bd58d2;
  wire bd58d3;
  wire bd58d4;
  wire bd58d5;
  wire bd58d6;
  wire bd58d7;
  wire bd58d8;
  wire bd58d9;
  wire bd58da;
  wire bd58db;
  wire bd58e4;
  wire bd58e5;
  wire bd58e6;
  wire bd58e7;
  wire bd58e8;
  wire bd58e9;
  wire bd58ea;
  wire bd58eb;
  wire bd58ec;
  wire bd58ed;
  wire bd58ee;
  wire bd58ef;
  wire bd58f0;
  wire bd58f1;
  wire bd58f2;
  wire bd58f3;
  wire bd58f4;
  wire bd58f5;
  wire bd58f6;
  wire bd58f7;
  wire bd58f8;
  wire bd58f9;
  wire bd58fa;
  wire bd58fb;
  wire bd58fc;
  wire bd58fd;
  wire bd58fe;
  wire bd58ff;
  wire bd5900;
  wire bd5901;
  wire bd5902;
  wire bd5903;
  wire bd5904;
  wire bd5905;
  wire bd5906;
  wire bd5907;
  wire bd5908;
  wire bd5909;
  wire bd590a;
  wire bd590b;
  wire bd590c;
  wire bd590d;
  wire bd590e;
  wire bd590f;
  wire bd5910;
  wire bd5911;
  wire bd5912;
  wire bd5913;
  wire bd5914;
  wire bd5915;
  wire bd5916;
  wire bd5917;
  wire bd5918;
  wire bd5919;
  wire bd591a;
  wire bd591b;
  wire bd591c;
  wire bd591d;
  wire bd591e;
  wire bd591f;
  wire bd5920;
  wire bd5921;
  wire bd5922;
  wire bd5923;
  wire bd5924;
  wire bd5925;
  wire bd5926;
  wire bd5927;
  wire bd5928;
  wire bd5929;
  wire bd592a;
  wire bd592b;
  wire bd592c;
  wire bd592d;
  wire bd592e;
  wire bd592f;
  wire bd5930;
  wire bd5931;
  wire bd5932;
  wire bd5933;
  wire bd5934;
  wire bd5935;
  wire bd5936;
  wire bd5937;
  wire bd5938;
  wire bd5939;
  wire bd593a;
  wire bd593b;
  wire bd593c;
  wire bd593d;
  wire bd593e;
  wire bd593f;
  wire bd5940;
  wire bd5941;
  wire bd5942;
  wire v845574;
  wire bcd5a7;
  wire v845562;
  wire b8f6e0;
  wire b8f6e1;
  wire b8f6e2;
  wire b8f6e3;
  wire b8f6e4;
  wire b8f6e5;
  wire b8f6e6;
  wire b8f6e7;
  wire b8f743;
  wire b8f744;
  wire b8f745;
  wire b8f746;
  wire b8f747;
  wire b8f748;
  wire b8f749;
  wire b8f74a;
  wire b8f74b;
  wire b8f74c;
  wire b8f74d;
  wire b8ef50;
  wire b8ef51;
  wire b8ef52;
  wire b8ef53;
  wire ba7c64;
  wire ba7c65;
  wire ba7c66;
  wire ba7c67;
  wire ba7c68;
  wire ba7c69;
  wire ba7c6a;
  wire ba7c6b;
  wire ba7c6c;
  wire ba7c6d;
  wire ba7c6e;
  wire ba7c6f;
  wire ba7c70;
  wire ba7c71;
  wire ba7c72;
  wire ba7c73;
  wire ba7c74;
  wire ba7c75;
  wire ba7c76;
  wire ba7c77;
  wire ba7c78;
  wire ba7c79;
  wire ba7c7a;
  wire ba7c7b;
  wire ba7c7c;
  wire ba7c7d;
  wire ba7c7e;
  wire ba7c7f;
  wire ba7c80;
  wire ba7c81;
  wire c74198;
  wire c74202;
  wire b0ed8b;
  wire b5b407;
  wire b5b408;
  wire b578f1;
  wire b578f2;
  wire b578f3;
  wire b578f4;
  wire b578f5;
  wire v8b08c1;
  wire b578f6;
  wire b578f7;
  wire b578f8;
  wire b578f9;
  wire b578fa;
  wire b578fb;
  wire b578fc;
  wire b578fd;
  wire b578fe;
  wire b578ff;
  wire b57900;
  wire b57901;
  wire b57902;
  wire b57903;
  wire b57904;
  wire b57905;
  wire b57906;
  wire b57907;
  wire b57908;
  wire b57909;
  wire b5790a;
  wire b5793f;
  wire b57940;
  wire b57941;
  wire b57942;
  wire b57943;
  wire b57944;
  wire b57945;
  wire b57946;
  wire b57947;
  wire b57948;
  wire b5b409;
  wire b57949;
  wire b5794a;
  wire b5794b;
  wire b5794c;
  wire b5794d;
  wire b5794e;
  wire b5794f;
  wire b57950;
  wire b57951;
  wire b57952;
  wire b57953;
  wire b57954;
  wire b57955;
  wire b57956;
  wire b57957;
  wire b57958;
  wire b57959;
  wire b5795a;
  wire b5795b;
  wire b57982;
  wire b57983;
  wire b57984;
  wire b57985;
  wire b57986;
  wire b57987;
  wire b57988;
  wire b57989;
  wire b5798a;
  wire b5798b;
  wire b5799c;
  wire b579af;
  wire b579b0;
  wire b579b1;
  wire b579b2;
  wire b579b3;
  wire b579b4;
  wire b579b5;
  wire b579b6;
  wire b579b7;
  wire b579b8;
  wire b579b9;
  wire b579ba;
  wire b579bb;
  wire b579bc;
  wire b579bd;
  wire b579be;
  wire b579bf;
  wire b579c0;
  wire b579c1;
  wire b579c2;
  wire b579c3;
  wire b579c4;
  wire b579c5;
  wire b579c6;
  wire b579c7;
  wire b579c8;
  wire b579c9;
  wire b579ca;
  wire b579cb;
  wire b579cc;
  wire b579cd;
  wire b579ce;
  wire b579cf;
  wire b579d0;
  wire b579d1;
  wire b579d2;
  wire b579d3;
  wire b579d4;
  wire b579d5;
  wire b579d6;
  wire b579d7;
  wire b579d8;
  wire b579d9;
  wire b579da;
  wire b579db;
  wire b579dc;
  wire b579dd;
  wire b579de;
  wire b579df;
  wire b579e0;
  wire b579e1;
  wire b579e2;
  wire b579e3;
  wire b579e4;
  wire b579e5;
  wire b579e6;
  wire b579e7;
  wire b579e8;
  wire b579e9;
  wire b579ea;
  wire b579eb;
  wire b579ec;
  wire b579ed;
  wire b579ee;
  wire b579ef;
  wire b579f0;
  wire b579f1;
  wire b57a0d;
  wire b57a0e;
  wire b57a0f;
  wire b57a10;
  wire b57a11;
  wire b57a12;
  wire b57a1a;
  wire b57a1b;
  wire b57a1c;
  wire b57a1d;
  wire b57a1e;
  wire b57a1f;
  wire b57a20;
  wire b57a21;
  wire b57a22;
  wire b57a23;
  wire b5b40a;
  wire b5b4ef;
  wire b57a25;
  wire b57a26;
  wire b57a27;
  wire b57a28;
  wire b57a29;
  wire b57a2a;
  wire b57a2b;
  wire b57a2c;
  wire b57a2d;
  wire b57a2e;
  wire b57a2f;
  wire b57a30;
  wire b57a31;
  wire b57a32;
  wire b57a33;
  wire b57a34;
  wire b57a35;
  wire b57a66;
  wire b57a67;
  wire b57a68;
  wire b57a69;
  wire b57a6a;
  wire b57a6b;
  wire b57a6c;
  wire b57a6d;
  wire b57a6e;
  wire b57a6f;
  wire b57a70;
  wire b57a71;
  wire b57a72;
  wire b57a73;
  wire b57a74;
  wire b57a75;
  wire b57a76;
  wire b57a77;
  wire b57a78;
  wire b57a79;
  wire b57a7a;
  wire b57a7b;
  wire b57a7c;
  wire b57a7d;
  wire b57a7e;
  wire b57a7f;
  wire b57a80;
  wire b57a81;
  wire b57a82;
  wire b57a83;
  wire b57a84;
  wire b57a85;
  wire b57a86;
  wire b57a87;
  wire b57a88;
  wire b57a89;
  wire b57a8a;
  wire b57a8b;
  wire b57a8c;
  wire b57a8d;
  wire b57a8e;
  wire b57a8f;
  wire b57ab2;
  wire b57ab3;
  wire b57ab4;
  wire b57ab5;
  wire b57ab6;
  wire b57ab7;
  wire b57ab8;
  wire b57ab9;
  wire b57aba;
  wire b57abb;
  wire b57abc;
  wire b57abd;
  wire b57abe;
  wire b57abf;
  wire b57ac0;
  wire b57ac1;
  wire b57ac2;
  wire b57ac3;
  wire b57ac4;
  wire b57ac5;
  wire b57ac6;
  wire b57ac7;
  wire b57ac8;
  wire b57ac9;
  wire b57aca;
  wire b57acb;
  wire b57acc;
  wire b57acd;
  wire b57ace;
  wire b57acf;
  wire b57ad0;
  wire b57ad1;
  wire b57ad2;
  wire b57ad3;
  wire b57adf;
  wire b57ae0;
  wire b57ae1;
  wire b57ae2;
  wire b57ae3;
  wire b57ae4;
  wire b57ae5;
  wire b57ae6;
  wire b57ae7;
  wire b57ae8;
  wire b57ae9;
  wire b57aea;
  wire b57aeb;
  wire b57aec;
  wire b57aed;
  wire b57aee;
  wire b57af0;
  wire b57af1;
  wire b57af2;
  wire b57af3;
  wire b57af4;
  wire b57af5;
  wire b57af6;
  wire b57af7;
  wire b57b57;
  wire b57b58;
  wire b57b59;
  wire b57b5a;
  wire b57b5b;
  wire b57b5c;
  wire b573d7;
  wire b573d8;
  wire b573d9;
  wire b573da;
  wire b573db;
  wire b573dc;
  wire b573dd;
  wire b573de;
  wire b573df;
  wire b573e0;
  wire b573e1;
  wire b573e2;
  wire b573e3;
  wire b573e4;
  wire b573e5;
  wire b573e6;
  wire b573e7;
  wire b573e8;
  wire b573f6;
  wire b573f7;
  wire b573f8;
  wire b573f9;
  wire b573fa;
  wire b573fb;
  wire b573fc;
  wire b573fd;
  wire b573fe;
  wire b573ff;
  wire b57400;
  wire b57401;
  wire b57402;
  wire b57403;
  wire b57404;
  wire b57405;
  wire b57406;
  wire b57407;
  wire b57408;
  wire b57409;
  wire b5740a;
  wire b5740b;
  wire b5740c;
  wire b5740d;
  wire b5740e;
  wire b5740f;
  wire b57410;
  wire b57411;
  wire b57412;
  wire b57413;
  wire b57414;
  wire b57415;
  wire b57416;
  wire b57417;
  wire b57418;
  wire b57419;
  wire b5741a;
  wire b5741b;
  wire b5741c;
  wire b5741d;
  wire b5741e;
  wire b5741f;
  wire b57420;
  wire b57421;
  wire b57422;
  wire b57423;
  wire b57424;
  wire b57425;
  wire b57426;
  wire b57427;
  wire b57428;
  wire b57429;
  wire b5742a;
  wire b5742b;
  wire b5742c;
  wire b5742d;
  wire b5742e;
  wire b5742f;
  wire b57430;
  wire b57431;
  wire b57432;
  wire b57433;
  wire b57434;
  wire b57435;
  wire b57436;
  wire b57437;
  wire b57438;
  wire b57439;
  wire b5743a;
  wire b5743b;
  wire b5743c;
  wire b5743d;
  wire b5743e;
  wire b5743f;
  wire b57440;
  wire b57441;
  wire b57442;
  wire b57443;
  wire b57444;
  wire b57445;
  wire b57446;
  wire b57447;
  wire b57448;
  wire b57449;
  wire b5744a;
  wire b5744b;
  wire b5744c;
  wire b5744d;
  wire b5744e;
  wire b5744f;
  wire b57450;
  wire b574b1;
  wire b574b2;
  wire b574b3;
  wire b574b4;
  wire b574b5;
  wire b574b6;
  wire b574b7;
  wire b574b8;
  wire b574b9;
  wire b574ba;
  wire b574bb;
  wire b574bc;
  wire b574bd;
  wire b574be;
  wire b574bf;
  wire b574c0;
  wire b574c1;
  wire b574c2;
  wire b574c3;
  wire b574c4;
  wire b574c5;
  wire b574c6;
  wire b574c7;
  wire b574c8;
  wire b574c9;
  wire b574ca;
  wire b574cb;
  wire b574cc;
  wire b574cd;
  wire b574ce;
  wire b574cf;
  wire b574d0;
  wire b574d1;
  wire b574d2;
  wire b574d3;
  wire b574d4;
  wire b574d5;
  wire b574d6;
  wire b574d7;
  wire b574d8;
  wire b574f9;
  wire b574fa;
  wire b574fb;
  wire b574fc;
  wire b574fd;
  wire b574fe;
  wire b574ff;
  wire b57500;
  wire b57501;
  wire b57502;
  wire b57503;
  wire b57504;
  wire b57506;
  wire b57507;
  wire b57508;
  wire b57509;
  wire b57532;
  wire b57533;
  wire b57534;
  wire b57535;
  wire b57536;
  wire b57537;
  wire b57538;
  wire v8a9702;
  wire v92e9d9;
  wire v85746a;
  wire v91784a;
  wire v882b8e;
  wire v857467;
  wire v9f7c93;
  wire v9f7c94;
  wire v9f7c95;
  wire v9f7c96;
  wire v9f7c97;
  wire v9f7c98;
  wire v9f7c99;
  wire v9f7c9a;
  wire v9f7c9b;
  wire v9f7c9c;
  wire v93a916;
  wire v857440;
  wire c6d44d;
  wire v9f7c9d;
  wire v9f7c9e;
  wire v9f7c9f;
  wire v9f7ca0;
  wire v9f7ca1;
  wire v9f7ca2;
  wire v9f7ca3;
  wire v9f7ca4;
  wire v9f7ca5;
  wire v9f7ca6;
  wire v9f7ca7;
  wire v9f7ca8;
  wire v9f7ca9;
  wire v9f7caa;
  wire v9f7cab;
  wire v9f7cac;
  wire v9f7cad;
  wire v9f7cae;
  wire v9f7caf;
  wire v9f7cb0;
  wire v9f7cb1;
  wire v9f7cb2;
  wire v9f7cb3;
  wire v9f7cb4;
  wire v9f7cb5;
  wire v9f7cb6;
  wire v9f7cb7;
  wire v9f7cb8;
  wire v9f7cb9;
  wire v9f7cba;
  wire v9f7cbb;
  wire v9f7cbc;
  wire v9f7cbd;
  wire v9f7cbe;
  wire v9f7cbf;
  wire v9f7cc0;
  wire v9f7cc1;
  wire v9f7cc2;
  wire v9f7cc3;
  wire v9f7cc4;
  wire v9f7cc5;
  wire v9f7cc6;
  wire v9f7cc7;
  wire v9f7cc8;
  wire v9f7cc9;
  wire v9f7cca;
  wire v9f7ccb;
  wire v9f7ccc;
  wire v9f7ccd;
  wire v9f7cce;
  wire v9f7ccf;
  wire v9f7cd0;
  wire v9f7cd1;
  wire v9f7cd2;
  wire v9f7cd3;
  wire v9f7cd4;
  wire v9f7cd5;
  wire v9f7cd6;
  wire v9f7cd7;
  wire v9f7cd8;
  wire v9f7cd9;
  wire v9f7cda;
  wire v9f7cdb;
  wire v9f7cdc;
  wire v9f7cdd;
  wire v9f7cde;
  wire v9f7cdf;
  wire v9f7ce0;
  wire v9f7ce1;
  wire v9f7ce2;
  wire v9f7ce3;
  wire v9f7ce4;
  wire v9f7ce5;
  wire v9f7ce6;
  wire v9f7ce7;
  wire v9f7ce8;
  wire v9f7ce9;
  wire v9f7cea;
  wire v9f7ceb;
  wire v9f7cec;
  wire v9f7ced;
  wire v9f7cee;
  wire v9f7cef;
  wire v9f7cf0;
  wire v9f7cf1;
  wire v9fa31b;
  wire v9f7cf2;
  wire v9f7cf3;
  wire v9f7cf4;
  wire v9f7cf5;
  wire v9f7cf6;
  wire v9f7cf7;
  wire v9f7cf8;
  wire v9f7cf9;
  wire v9f7cfa;
  wire v9f7cfb;
  wire v9f7cfc;
  wire v9f7cfd;
  wire v9f7cfe;
  wire v9f7cff;
  wire v9f7d00;
  wire v9f7d01;
  wire v9f7d02;
  wire v9f7d03;
  wire v9f7d04;
  wire v9f7d05;
  wire v9f7d06;
  wire v9f7d07;
  wire v9f7d08;
  wire v9f7d09;
  wire v9f7d0a;
  wire v9f7d0b;
  wire v9f7d0c;
  wire v9f7d0d;
  wire v9f7d0e;
  wire v9f7d0f;
  wire v9f7d10;
  wire v9f7d11;
  wire v9f7d12;
  wire v9f7d13;
  wire v9f7d14;
  wire v9f7d15;
  wire v9f7d16;
  wire v9f7d17;
  wire v9f7d18;
  wire v9f7d19;
  wire v9f7d1a;
  wire v9f7d1b;
  wire v9f7d1c;
  wire v9f7d1d;
  wire v9f7d1e;
  wire v9f7d1f;
  wire v9f7d20;
  wire v9f7d21;
  wire v9f7d22;
  wire v9f7d23;
  wire v9f7d24;
  wire v9f7d25;
  wire v9f7d26;
  wire v9f7d27;
  wire v9f7d28;
  wire v9f7d29;
  wire v9f7d2a;
  wire v9f7d2b;
  wire v9f7d2c;
  wire v9f7d2d;
  wire v9f7d2e;
  wire v9f7d2f;
  wire v9f7d30;
  wire v9f7d31;
  wire v9f7d32;
  wire v9f7d33;
  wire v9f7d34;
  wire v9f7d35;
  wire v9f7d36;
  wire v9f7d37;
  wire v9f7d38;
  wire v9f7d39;
  wire b06735;
  wire v9f7d3a;
  wire v9f7d3b;
  wire v9f7d3c;
  wire v9f7d3d;
  wire v9f7d3e;
  wire v9f7d3f;
  wire v9f7d40;
  wire v9f7d41;
  wire v9f7d42;
  wire v9f7d43;
  wire v9f7d44;
  wire v9f7d45;
  wire v9f7d46;
  wire v9f7d47;
  wire v9f7d48;
  wire v9f7d49;
  wire v9f7d4a;
  wire v9f7d4b;
  wire v9f7d4c;
  wire v9f7d4d;
  wire v9f7d4e;
  wire v9f7d4f;
  wire v9f7d50;
  wire v9f7d51;
  wire v9f7d52;
  wire v9f7d53;
  wire v9f7d54;
  wire v9f7d55;
  wire v9f7d56;
  wire v9f7d57;
  wire v9f7d58;
  wire v9f7d59;
  wire v9f7d5a;
  wire v9f7d5b;
  wire v9f7d5c;
  wire v9f7d5d;
  wire v9f7d5e;
  wire v9f7d5f;
  wire v9f7d60;
  wire v9f7d61;
  wire v9f7d62;
  wire v9f7d63;
  wire v9f7d64;
  wire v9f7d65;
  wire v9f7d66;
  wire v9f7d67;
  wire v9f7d68;
  wire v9f7d69;
  wire v9f7d6a;
  wire v9f7d6b;
  wire v9f7d6c;
  wire v9f7d6d;
  wire v9f7d6e;
  wire v9f7d6f;
  wire v9f7d70;
  wire v9f7d71;
  wire v9f7d72;
  wire v9f7d73;
  wire v9f7d74;
  wire v9f7d75;
  wire v9f7d76;
  wire v9f7d77;
  wire v9f7d78;
  wire v9f7d79;
  wire v9f7d7a;
  wire v9f7d7b;
  wire v9f7d7c;
  wire v9f7d7d;
  wire v9f7d7e;
  wire v9f7d7f;
  wire v9f7d80;
  wire v9f7d81;
  wire v9f7d82;
  wire v9f7d83;
  wire v9f7d84;
  wire v9f7d85;
  wire v9f7d86;
  wire v9f7d87;
  wire v9f7d88;
  wire v9f7d89;
  wire v9f7d8a;
  wire v9f7d8b;
  wire v9f7d8c;
  wire v9f7d8d;
  wire v9f7d8e;
  wire v9f7d8f;
  wire v9f7d90;
  wire v9f7d91;
  wire v9f7d92;
  wire v9f7d93;
  wire v9f7d94;
  wire v9f7d95;
  wire v9f7d96;
  wire v9f7d97;
  wire v9f7d98;
  wire v9f7d99;
  wire v9f7d9a;
  wire v9f7d9b;
  wire v9f7d9c;
  wire v9f7d9d;
  wire v9f7d9e;
  wire v9f7d9f;
  wire v9f7da0;
  wire v9f7da1;
  wire v9f7da2;
  wire v9f7da3;
  wire v9f7da4;
  wire v9f7da5;
  wire v9f7da6;
  wire v9f7da7;
  wire v9f7da8;
  wire v9f7da9;
  wire v9f7daa;
  wire v9f7dab;
  wire v9f7dac;
  wire v9f7dad;
  wire v9f7dae;
  wire v9f7daf;
  wire v9f7db0;
  wire v9f7db1;
  wire v9f7db2;
  wire v9f7db3;
  wire v9f7db4;
  wire v9f7db5;
  wire v9f7db6;
  wire v9f7db7;
  wire v9f7db8;
  wire v9f7db9;
  wire v9f7dba;
  wire v9f7dbb;
  wire v9f7dbc;
  wire v9f7dbd;
  wire v9f7dbe;
  wire v9f7dbf;
  wire v9f7dc0;
  wire v9f7dc1;
  wire v9f7dc2;
  wire v9f7dc3;
  wire v9f7dc4;
  wire v9f7dc5;
  wire v9f7dc6;
  wire v9f7dc7;
  wire v9f7dc8;
  wire v9f7dc9;
  wire v9f7dca;
  wire v9f7dcb;
  wire v9f7dcc;
  wire v9f7dcd;
  wire v9f7dce;
  wire v9f7dcf;
  wire v9f7dd0;
  wire v9f7dd1;
  wire v9f7dd2;
  wire v9f7dd3;
  wire v9f7dd4;
  wire v9f7dd5;
  wire v9f7dd6;
  wire v9f7dd7;
  wire v9f7dd8;
  wire v9f7dd9;
  wire v9f7dda;
  wire v9f7ddb;
  wire v9f7ddc;
  wire v9f7ddd;
  wire v9f7dde;
  wire v9f7ddf;
  wire v9f7de0;
  wire v9f7de1;
  wire v9f7de2;
  wire v9f7de3;
  wire v9f7de4;
  wire v9f7de5;
  wire v9f7de6;
  wire v9f7de7;
  wire v9f7de8;
  wire v9f7de9;
  wire v9f7dea;
  wire v9f7deb;
  wire v9f7dec;
  wire v9f7ded;
  wire v9f7dee;
  wire v9f7def;
  wire v9f7df0;
  wire v9f7df1;
  wire v9f7df2;
  wire v9f7df3;
  wire v9f7df4;
  wire v9f7df5;
  wire v9f7df6;
  wire v9f7df7;
  wire v9f7df8;
  wire v9f7df9;
  wire v9f7dfa;
  wire v9f7dfb;
  wire v9f7dfc;
  wire v9f7dfd;
  wire v9f7dfe;
  wire v9f7dff;
  wire v9f7e00;
  wire v9f7e01;
  wire v9f7e02;
  wire v9f7e03;
  wire v9f7e04;
  wire v9f7e05;
  wire v9f7e06;
  wire v9f7e07;
  wire v9f7e08;
  wire v9f7e09;
  wire v9f7e0a;
  wire v9f7e0b;
  wire v9f7e0c;
  wire v9f7e0d;
  wire v9f7e0e;
  wire v9f7e0f;
  wire v9f7e10;
  wire v9f7e11;
  wire v9f7e12;
  wire v9f7e13;
  wire v9f7e14;
  wire v9f7e15;
  wire v9f7e16;
  wire v9f7e17;
  wire v9f7e18;
  wire v9f7e19;
  wire v9f7e1a;
  wire v9f7e1b;
  wire v9f7e1c;
  wire v9f7e1d;
  wire v9f7e1e;
  wire v9f7e1f;
  wire v9f7e20;
  wire v9f7e21;
  wire v9f7e22;
  wire v9f7e23;
  wire v9f7e24;
  wire v9f7e25;
  wire v9f7e26;
  wire v9f7e27;
  wire v9f7e28;
  wire v9f7e29;
  wire v9f7e2a;
  wire v9f7e2b;
  wire v9f7e2c;
  wire v9f7e2d;
  wire v9f7e2e;
  wire v9f7e2f;
  wire v9f7e30;
  wire v9f7e31;
  wire v9f7e32;
  wire v9f7e33;
  wire v9f7e34;
  wire v9f7e35;
  wire v9f7e36;
  wire v9f7e37;
  wire v9f7e38;
  wire v9f7e39;
  wire v9f7e3a;
  wire v9f7e3b;
  wire v9f7e3c;
  wire v9f7e3d;
  wire v9f7e3e;
  wire v9f7e3f;
  wire v9f7e40;
  wire v9f7e41;
  wire v9f7e42;
  wire v9f7645;
  wire v9f7646;
  wire v9f7647;
  wire v9f7648;
  wire v9f7649;
  wire v9f764a;
  wire v9f764b;
  wire v9f764c;
  wire v9f764d;
  wire v9f764e;
  wire v9f764f;
  wire v9f7650;
  wire v9f7651;
  wire v9f7652;
  wire v9f7653;
  wire v9f7654;
  wire v9f7655;
  wire v9f7656;
  wire v9f7657;
  wire v9f7658;
  wire v9f7659;
  wire v9f765a;
  wire v9f765b;
  wire v9f765c;
  wire v9f765d;
  wire v9f765e;
  wire v9f765f;
  wire v9f7660;
  wire v9f7661;
  wire v9f7662;
  wire v9f7663;
  wire v9f7664;
  wire v9f7665;
  wire v9f7666;
  wire v9f7667;
  wire v9f7668;
  wire v9f7669;
  wire v9f766a;
  wire v9f766b;
  wire v9f766c;
  wire v9f766d;
  wire v9f766e;
  wire v9f766f;
  wire v9f7670;
  wire v9f7671;
  wire v9f7672;
  wire v9f7673;
  wire v9f7674;
  wire v9f7675;
  wire v9f7676;
  wire v9f7677;
  wire v9f7678;
  wire v9f7679;
  wire v9f767a;
  wire v9f767b;
  wire v9f767c;
  wire v9f767d;
  wire v9f767e;
  wire v9f767f;
  wire v9f7680;
  wire v9f7681;
  wire v9f7682;
  wire v9f7683;
  wire v9f7684;
  wire v9f7685;
  wire v9f7686;
  wire v9f7687;
  wire v9f7688;
  wire v9f7689;
  wire v9f768a;
  wire v9f768b;
  wire v9f768c;
  wire v9f768d;
  wire v9f768e;
  wire v9f768f;
  wire v9f7690;
  wire v9f7691;
  wire v9f7692;
  wire v9f7693;
  wire v9f7694;
  wire v9f7695;
  wire v9f7696;
  wire v9f7697;
  wire v9f7698;
  wire v9f7699;
  wire v9f769a;
  wire v9f769b;
  wire v9f769c;
  wire v9f769d;
  wire v9f769e;
  wire v9f769f;
  wire v9f76a0;
  wire v9f76a1;
  wire v9f76a2;
  wire v9f76a3;
  wire v9f76a4;
  wire v9f76a5;
  wire v9f76a6;
  wire v9f76a7;
  wire v9f76a8;
  wire v9f76a9;
  wire v9f76aa;
  wire v9f76ab;
  wire v9f76ac;
  wire v9f76ad;
  wire v9f76ae;
  wire v9f76af;
  wire v9f76b0;
  wire v9f76b1;
  wire v9f76b2;
  wire v9f76b3;
  wire v9f76b4;
  wire v9f76b5;
  wire v9f76b6;
  wire v9f76b7;
  wire v9f76b8;
  wire v9f76b9;
  wire v9f76ba;
  wire v9f76bb;
  wire v9f76bc;
  wire v9f76bd;
  wire v9f76be;
  wire v9f76bf;
  wire v9f76c0;
  wire v9f76c1;
  wire v9f76c2;
  wire v9f76c3;
  wire v9f76c4;
  wire v9f76c5;
  wire v9f76c6;
  wire v9f76c7;
  wire v9f76c8;
  wire v9f76c9;
  wire v9f76ca;
  wire v9f76cb;
  wire v9f76cc;
  wire v9f76cd;
  wire v9f76ce;
  wire v9f76cf;
  wire v9f76d0;
  wire v9f76d1;
  wire v9f76d2;
  wire v9f76d3;
  wire v9f76d4;
  wire v9f76d5;
  wire v9f76d6;
  wire v9f76d7;
  wire v9f76d8;
  wire v9f76d9;
  wire v9f76da;
  wire v9f76db;
  wire v9f76dc;
  wire v9f76dd;
  wire v9f76de;
  wire v9f76df;
  wire v9f76e0;
  wire v9f76e1;
  wire v9f76e2;
  wire v9f76e3;
  wire v9f76e4;
  wire v9f76e5;
  wire v9f76e6;
  wire v9f76e7;
  wire v9f76e8;
  wire v9f76e9;
  wire v9f76ea;
  wire v9f76eb;
  wire v9f76ec;
  wire v9f76ed;
  wire v9f76ee;
  wire v9f76ef;
  wire v9f76f0;
  wire v9f76f1;
  wire v9f76f2;
  wire v9f76f3;
  wire v9f76f4;
  wire v9f76f5;
  wire v9f76f6;
  wire v9f76f7;
  wire v9f76f8;
  wire v9f76f9;
  wire v9f76fa;
  wire v9f76fb;
  wire v9f76fc;
  wire v9f76fd;
  wire v9f76fe;
  wire v9f76ff;
  wire v9f7700;
  wire v9f7701;
  wire v9f7702;
  wire v9f7703;
  wire v9f7704;
  wire v9f7705;
  wire v9f7706;
  wire v9f7707;
  wire v9f7708;
  wire v9f7709;
  wire v9f770a;
  wire v9f770b;
  wire v9f770c;
  wire v9f770d;
  wire v9f770e;
  wire v9f770f;
  wire v9f7710;
  wire v9f7711;
  wire v9f7712;
  wire v9f7713;
  wire v9f7714;
  wire v9f7715;
  wire v9f7716;
  wire v9f7717;
  wire v9f7718;
  wire v9f7719;
  wire v9f771a;
  wire v9f771b;
  wire v9f771c;
  wire v9f771d;
  wire v9f771e;
  wire v9f771f;
  wire v9f7720;
  wire v9f7721;
  wire v9f7722;
  wire v9f7723;
  wire v9f7724;
  wire v9f7725;
  wire v9f7726;
  wire v9f7727;
  wire v9f7728;
  wire v9f772a;
  wire v9f772b;
  wire v9f772c;
  wire v9f772d;
  wire v9f772e;
  wire v9f772f;
  wire v9f7730;
  wire v9f7731;
  wire v9f7732;
  wire v9f7733;
  wire v9f7734;
  wire v9f7735;
  wire v9f7736;
  wire v9f7737;
  wire v9f7738;
  wire v9f7739;
  wire v9f773a;
  wire v9f773b;
  wire v9f773c;
  wire v9f773d;
  wire v9f773e;
  wire v9f773f;
  wire v9f7740;
  wire v9f7741;
  wire v9f7742;
  wire v9f7743;
  wire v9f7744;
  wire v9f7745;
  wire v9f7746;
  wire v9f7747;
  wire v9f7748;
  wire v9f7749;
  wire v9f774a;
  wire v9f774b;
  wire v9f774c;
  wire v9f774d;
  wire v9f774e;
  wire v9f774f;
  wire v9f7750;
  wire v9f7751;
  wire v9f7752;
  wire v9f7753;
  wire v9f7754;
  wire v9f7755;
  wire v9f7756;
  wire v9f7757;
  wire v9f7758;
  wire v9f7759;
  wire v9f775a;
  wire v9f775b;
  wire v9f775c;
  wire v9f775d;
  wire v9f775e;
  wire v9f775f;
  wire v9f7760;
  wire v9f7761;
  wire v9f7762;
  wire v9f7763;
  wire v9f7764;
  wire v9f7765;
  wire v9f7766;
  wire v9f7767;
  wire v9f7768;
  wire v9f7769;
  wire v9f776a;
  wire v9f776b;
  wire v9f776c;
  wire v9f776d;
  wire v9f776e;
  wire v9f776f;
  wire v9f7770;
  wire v9f7771;
  wire v9f7772;
  wire v9f7773;
  wire v9f7774;
  wire v9f7775;
  wire v9f7776;
  wire v9f7777;
  wire v9f7778;
  wire v9f7779;
  wire v9f777a;
  wire v9f777b;
  wire v9f777c;
  wire v9f777d;
  wire v9f777e;
  wire v9f777f;
  wire v9f7780;
  wire v9f7781;
  wire v9f7782;
  wire v9f7783;
  wire v9f7784;
  wire v9f7785;
  wire v9f7786;
  wire v9f7787;
  wire v9f7788;
  wire v9f7789;
  wire v9f778a;
  wire v9f778b;
  wire v9f778c;
  wire v9f778d;
  wire v9f778e;
  wire v9f778f;
  wire v9f7790;
  wire v9f7791;
  wire v9f7792;
  wire v9f7793;
  wire v9f7794;
  wire v9f7795;
  wire v9f7796;
  wire v9f7797;
  wire v9f7798;
  wire v9f7799;
  wire v9f779a;
  wire v9f779b;
  wire v9f779c;
  wire v9f779d;
  wire v9f779e;
  wire v9f779f;
  wire v9f77a0;
  wire v9f77a1;
  wire v9f77a2;
  wire v9f77a3;
  wire v9f77a4;
  wire v9f77a5;
  wire v9f77a6;
  wire v9f77a7;
  wire v9f77a8;
  wire v9f77a9;
  wire v9f77aa;
  wire v9f77ab;
  wire v9f77ac;
  wire v9f77ad;
  wire v9f77ae;
  wire v9f77af;
  wire v9f77b0;
  wire v9f77b1;
  wire v9f77b2;
  wire v9f77b3;
  wire v9f77b4;
  wire v9f77b5;
  wire v9f77b6;
  wire v9f77b7;
  wire v9f77b8;
  wire v9f77b9;
  wire v9f77ba;
  wire v9f77bb;
  wire v9f77bc;
  wire v9f77bd;
  wire v9f77be;
  wire v9f77bf;
  wire v9f77c0;
  wire v9f77c1;
  wire v9f77c2;
  wire v9f77c3;
  wire v9f77c4;
  wire v9f77c5;
  wire v9f77c6;
  wire v9f77c7;
  wire v9f77c8;
  wire v9f77c9;
  wire v9f77ca;
  wire v9f77cb;
  wire v9f77cc;
  wire v9f77cd;
  wire v9f77ce;
  wire v9f77cf;
  wire v9f77d0;
  wire v9f77d1;
  wire v9f77d2;
  wire v9f77d3;
  wire v9f77d4;
  wire v9f77d5;
  wire v9f77d6;
  wire v9f77d7;
  wire v9f77d8;
  wire v9f77d9;
  wire v9f77da;
  wire v9f77db;
  wire v9f77dc;
  wire v9f77dd;
  wire v9f77de;
  wire v9f77df;
  wire v9f77e0;
  wire v9f77e1;
  wire v9f77e2;
  wire v9f77e3;
  wire v9f77e4;
  wire v9f77e5;
  wire v9f77e6;
  wire v9f77e7;
  wire v9f77e8;
  wire v9f77e9;
  wire v9f77ea;
  wire v9f77eb;
  wire v9f77ec;
  wire v9f77ed;
  wire v9f77ee;
  wire v9f77ef;
  wire v9f77f0;
  wire v9f77f1;
  wire v9f77f2;
  wire v9f77f3;
  wire v9f77f4;
  wire v9f77f5;
  wire v9f77f6;
  wire v9f77f7;
  wire v9f77f8;
  wire v9f77f9;
  wire v9f77fa;
  wire v9f77fb;
  wire v9f77fc;
  wire v9f77fd;
  wire v9f77fe;
  wire v9f77ff;
  wire v9f7800;
  wire v9f7801;
  wire v9f7802;
  wire v9f7803;
  wire v9f7804;
  wire v9f7805;
  wire v9f7806;
  wire v9f7807;
  wire v9f7808;
  wire v9f7809;
  wire v9f780a;
  wire v9f780b;
  wire v9f780c;
  wire v9f780d;
  wire v9f780e;
  wire v9f780f;
  wire v9f7810;
  wire v9f7811;
  wire v9f7812;
  wire v9f7813;
  wire v9f7814;
  wire v9f7815;
  wire v9f7816;
  wire v9f7817;
  wire v9f7818;
  wire v9f7819;
  wire v9f781a;
  wire v9f781b;
  wire v9f781c;
  wire v9f781d;
  wire v9f781e;
  wire v9f781f;
  wire v9f7820;
  wire v9f7821;
  wire v9f7822;
  wire v9f7823;
  wire v9f7824;
  wire v9f7825;
  wire v9f7826;
  wire v9f7827;
  wire v9f7828;
  wire v9f7829;
  wire v9f782a;
  wire v9f782b;
  wire v9f782c;
  wire v9f782d;
  wire v9f782e;
  wire v9f782f;
  wire v9f7830;
  wire v9f7831;
  wire v9f7832;
  wire v9f7833;
  wire v9f7834;
  wire v9f7835;
  wire v9f7836;
  wire v9f7837;
  wire v9f7838;
  wire v9f7839;
  wire v9f783a;
  wire v9f783b;
  wire v9f783c;
  wire v9f783d;
  wire v9f783e;
  wire v9f783f;
  wire v9f7840;
  wire v9f7841;
  wire v9f7842;
  wire v9f7843;
  wire v9f7844;
  wire v9f7845;
  wire v9f7846;
  wire v9f7847;
  wire v9f7848;
  wire v9f7849;
  wire v9f784a;
  wire v9f784b;
  wire v9f784c;
  wire v9f784d;
  wire v9f784e;
  wire v9f784f;
  wire v9f7850;
  wire v9f7851;
  wire v9f7852;
  wire v9f7853;
  wire v9f7854;
  wire v9f7855;
  wire v9f7856;
  wire v9f7857;
  wire v9f7858;
  wire v9f7859;
  wire v9f785a;
  wire v9f785b;
  wire v9f785c;
  wire v9f785d;
  wire v9f785e;
  wire v9f785f;
  wire v9f7860;
  wire v9f7861;
  wire v9f7862;
  wire v9f7863;
  wire v9f7864;
  wire v9f7865;
  wire v9f7866;
  wire v9f7867;
  wire v9f7868;
  wire v9f7869;
  wire v9f786a;
  wire v9f786b;
  wire v9f786c;
  wire v9f786d;
  wire v9f786e;
  wire v9f786f;
  wire v9f7870;
  wire v9f7871;
  wire v9f7872;
  wire v9f7873;
  wire v9f7874;
  wire v9f7875;
  wire v9f7876;
  wire v9f7877;
  wire v9f7878;
  wire v9f7879;
  wire v9f787a;
  wire v9f787b;
  wire v9f787c;
  wire v9f787d;
  wire v9f787e;
  wire v9f787f;
  wire v9f7880;
  wire v9f7881;
  wire v9f7882;
  wire v9f7883;
  wire v9f7884;
  wire v9f7885;
  wire v9f7886;
  wire v9f7887;
  wire v9f7888;
  wire v9f7889;
  wire v9f788a;
  wire v9f788b;
  wire v9f788c;
  wire v9f788d;
  wire v9f788e;
  wire v9f788f;
  wire v9f7890;
  wire v9f7891;
  wire v9f7892;
  wire v9f7893;
  wire v9f7894;
  wire v9f7895;
  wire v9f7896;
  wire v9f7897;
  wire v9f7898;
  wire v9f7899;
  wire v9f789a;
  wire v9f789b;
  wire v9f789c;
  wire v9f789d;
  wire v9f789e;
  wire v9f789f;
  wire v9f78a0;
  wire v9f78a1;
  wire v9f78a2;
  wire v9f78a3;
  wire v9f78a4;
  wire v9f78a5;
  wire v9f78a6;
  wire v9f78a7;
  wire v9f78a8;
  wire v9f78a9;
  wire v9f78aa;
  wire v9f78ab;
  wire v9f78ac;
  wire v9f78ad;
  wire v9f78ae;
  wire v9f78af;
  wire v9f78b0;
  wire v9f78b1;
  wire b1cf24;
  wire b1cf25;
  wire b1cf26;
  wire b1cf27;
  wire b1cf28;
  wire b1cf29;
  wire b1cf2a;
  wire b1cf2b;
  wire b1cf2c;
  wire b1cf2d;
  wire b1cf2e;
  wire b1cf2f;
  wire b1cf30;
  wire b1cf31;
  wire b1cf32;
  wire b1cf33;
  wire b1cf34;
  wire b1cf35;
  wire b1cf37;
  wire b1cf38;
  wire b1cf3a;
  wire b1cf3b;
  wire b1cf3c;
  wire b1cf3d;
  wire b1cf3e;
  wire b1cf3f;
  wire b1cf40;
  wire b1cf41;
  wire b1cf42;
  wire b1cf43;
  wire b1cf45;
  wire b1cf46;
  wire b1cf47;
  wire b1cf48;
  wire b1cf49;
  wire b1cfb6;
  wire b1cfb7;
  wire b1cfb8;
  wire b1cfbe;
  wire b1cfbf;
  wire b1cfc0;
  wire b1cfc1;
  wire b1cfc2;
  wire b1cfc3;
  wire b1cfc4;
  wire b1cfc5;
  wire b1cfc6;
  wire b1cfc7;
  wire b1cfc8;
  wire b1cfc9;
  wire b1cfca;
  wire b1cfcb;
  wire b1cfcc;
  wire b1cfcd;
  wire b1cfce;
  wire b1cfcf;
  wire b1cfd0;
  wire b1cfd1;
  wire b1cfd2;
  wire b1cfd3;
  wire b1cfd4;
  wire b1cfd5;
  wire b1cff4;
  wire b1cff5;
  wire b1cff6;
  wire b1cff7;
  wire b1cff8;
  wire b1cff9;
  wire b1cffa;
  wire b1cffb;
  wire b1cffc;
  wire b1cffd;
  wire b1cffe;
  wire b1cfff;
  wire b1d000;
  wire b1d001;
  wire b1d002;
  wire b1d003;
  wire b1d004;
  wire b1d005;
  wire b1d006;
  wire b1d007;
  wire b1d00d;
  wire b1d00e;
  wire b1d00f;
  wire b1d010;
  wire b1d011;
  wire b1d012;
  wire b1d013;
  wire b1d014;
  wire b1d017;
  wire b1d018;
  wire b1d019;
  wire b1d01a;
  wire b1c82c;
  wire b1c82d;
  wire b1c82e;
  wire b1c82f;
  wire b1c840;
  wire b1c841;
  wire b1c842;
  wire b1c843;
  wire b1c844;
  wire b1c845;
  wire b1c846;
  wire b1c847;
  wire b1c848;
  wire b1c849;
  wire b1c84a;
  wire b1c84b;
  wire b1c84d;
  wire b1c84e;
  wire b1c84f;
  wire b1c850;
  wire b1c851;
  wire b1c852;
  wire b1c853;
  wire b1c854;
  wire b1c855;
  wire b1c856;
  wire b1c857;
  wire b1c858;
  wire b1c859;
  wire b1c85a;
  wire b1c85b;
  wire b1c85c;
  wire b1c85d;
  wire b1c85e;
  wire b1c85f;
  wire b1c860;
  wire b1c861;
  wire b1c862;
  wire b1c863;
  wire b1c864;
  wire b1c865;
  wire b1c866;
  wire b1c867;
  wire b1c868;
  wire b1c869;
  wire b1c86a;
  wire b1c86b;
  wire b1cae9;
  wire b1caea;
  wire b1caeb;
  wire b1caec;
  wire b1caed;
  wire b1caee;
  wire b1caf4;
  wire b1caf5;
  wire b1caf6;
  wire b1caf7;
  wire b1caf8;
  wire b1caf9;
  wire b1cafd;
  wire b1cafe;
  wire b1caff;
  wire b1cb00;
  wire b1cbf0;
  wire b1cbf1;
  wire b1cbf2;
  wire b1cbf3;
  wire b1cbf4;
  wire b1cbf5;
  wire b1cbf6;
  wire b1cbf9;
  wire b1cbfa;
  wire b1cbfd;
  wire b1cbfe;
  wire b1cbff;
  wire b1cc00;
  wire b1cc01;
  wire b1cc02;
  wire b1cc03;
  wire b1cc04;
  wire b1cc05;
  wire b1c45c;
  wire b1c45d;
  wire b1c45e;
  wire b1c495;
  wire b1c496;
  wire b1c497;
  wire b1c498;
  wire b1c4a3;
  wire b1c4a4;
  wire b1c4a5;
  wire b1c4a6;
  wire b1c4a7;
  wire b1c4ae;
  wire b1c4af;
  wire b1c4c3;
  wire b1c4c4;
  wire b1c4c5;
  wire b1c4c6;
  wire b1c4c7;
  wire b1c4c8;
  wire b1c4c9;
  wire b1c4ca;
  wire b1c4cb;
  wire b1c4cc;
  wire b1c4cd;
  wire b1c4ce;
  wire b1c4cf;
  wire b1c4d0;
  wire b1c50c;
  wire b1c50d;
  wire b1c50e;
  wire b1c55d;
  wire b1c55e;
  wire b1c55f;
  wire b1c560;
  wire b1c561;
  wire b1c562;
  wire b1c563;
  wire b1c564;
  wire b1c565;
  wire b1c566;
  wire b1c567;
  wire b1c568;
  wire b1c569;
  wire b1c56a;
  wire b1c56b;
  wire b1c56c;
  wire b1c56d;
  wire b1c56e;
  wire b1c57b;
  wire b1c57c;
  wire b1c57d;
  wire b1c57e;
  wire b1c57f;
  wire b1c580;
  wire b1c581;
  wire b1c582;
  wire b1c583;
  wire b1c584;
  wire b1c585;
  wire b1c586;
  wire b1c587;
  wire b1c588;
  wire b1c589;
  wire b1c58a;
  wire b1c58b;
  wire b1c5b3;
  wire b1c5b4;
  wire b1c5b5;
  wire b1c5b6;
  wire b1c5b7;
  wire b1c5b8;
  wire b1c5b9;
  wire b1c5ba;
  wire b1c5bb;
  wire b1c5bc;
  wire b1c5bd;
  wire b1c5be;
  wire b1c5bf;
  wire b1c5d7;
  wire b1c5d8;
  wire b1c5d9;
  wire b1c5da;
  wire b1c5db;
  wire b1c5dc;
  wire b1c5dd;
  wire b1c5de;
  wire b1c5df;
  wire b1c5e0;
  wire b1c5e1;
  wire b1c5e2;
  wire b1c5e3;
  wire b1c5e4;
  wire b1c5e5;
  wire b1c5e6;
  wire b1c5e7;
  wire b1c5e8;
  wire b1c5e9;
  wire b1c5ea;
  wire b1c5eb;
  wire b1c5ec;
  wire b1c5ed;
  wire b1c5ee;
  wire b1c5ef;
  wire b1c5f0;
  wire b1c5f1;
  wire b1c5f2;
  wire b1c5f3;
  wire b1c5f4;
  wire b1c5f5;
  wire b1c5f6;
  wire b1c5f7;
  wire b1c5f8;
  wire b1c5fc;
  wire b1c5fd;
  wire b1c5fe;
  wire b1c5ff;
  wire b1c600;
  wire b1c610;
  wire b1c611;
  wire b1c612;
  wire b1c613;
  wire b1c614;
  wire b1c615;
  wire b1c616;
  wire b1c617;
  wire b1c618;
  wire b1c619;
  wire b1c61a;
  wire b1c61b;
  wire b1c61c;
  wire b1c6b7;
  wire b1c6b8;
  wire b1c6b9;
  wire b1c6ba;
  wire b1c6bb;
  wire b1c6bc;
  wire b1c6bd;
  wire b1c6be;
  wire b1c6c7;
  wire b1c6c8;
  wire b1c6c9;
  wire b1c6ca;
  wire b1c6cb;
  wire b1c6cc;
  wire b1c6cd;
  wire b1c6ce;
  wire b1c6cf;
  wire b1c6da;
  wire b1c6db;
  wire b1c6dc;
  wire b1c6de;
  wire b1c6df;
  wire b1c6e0;
  wire b1c6f8;
  wire b1c6f9;
  wire b1c6fa;
  wire b1c6fb;
  wire b1c6fc;
  wire b1c6fd;
  wire b1c6fe;
  wire b1c700;
  wire b1c701;
  wire b1c702;
  wire b1c703;
  wire b1c704;
  wire b1c705;
  wire b1c706;
  wire b1c707;
  wire b1c708;
  wire b1c709;
  wire b1c70c;
  wire b1c70d;
  wire b1c70e;
  wire b1c70f;
  wire b1c710;
  wire b1c711;
  wire b1c712;
  wire b1c713;
  wire b1c714;
  wire b1c715;
  wire b1c716;
  wire b1c717;
  wire b1c718;
  wire b1c719;
  wire b1c71a;
  wire b1c71b;
  wire b1c71c;
  wire b1c71d;
  wire b1c71e;
  wire b1c71f;
  wire b1c720;
  wire b1c721;
  wire b1c722;
  wire b1c723;
  wire b1c724;
  wire b1c725;
  wire b1c726;
  wire b1c727;
  wire b1c728;
  wire b1c729;
  wire b1c72a;
  wire b1c72b;
  wire b1c72c;
  wire b1c72d;
  wire b1c72e;
  wire b1c72f;
  wire b1c730;
  wire b1c731;
  wire b1c732;
  wire b1c733;
  wire b1c734;
  wire b1c735;
  wire b1c736;
  wire b1c737;
  wire b1c738;
  wire b1c739;
  wire b1c73a;
  wire b1c73b;
  wire b1c73c;
  wire b1c73d;
  wire b1c73e;
  wire b1c73f;
  wire b1c740;
  wire b1c741;
  wire b1c742;
  wire b1c743;
  wire b1c744;
  wire b1c745;
  wire b1c746;
  wire b1c747;
  wire b1c748;
  wire b1c749;
  wire b1c74a;
  wire b1c74b;
  wire b1c74c;
  wire b1c74d;
  wire b1c74e;
  wire b1c74f;
  wire b1c750;
  wire b1c751;
  wire b1c752;
  wire b1c753;
  wire b1c754;
  wire b1c755;
  wire b1c756;
  wire b1c757;
  wire b1c758;
  wire b1c759;
  wire b1c75a;
  wire b1c75b;
  wire b1c75c;
  wire b1c75d;
  wire b1c75e;
  wire b1c75f;
  wire b1c760;
  wire b1c761;
  wire b1c762;
  wire b1c763;
  wire b1c764;
  wire b1c765;
  wire b1c766;
  wire b1c767;
  wire b1c768;
  wire b1c769;
  wire b1c76a;
  wire b1c76b;
  wire b1c76c;
  wire b1c76d;
  wire b1c76e;
  wire b1c76f;
  wire b1c770;
  wire b1c771;
  wire b1c772;
  wire b1c773;
  wire b1c774;
  wire b1c775;
  wire b1c776;
  wire b1c777;
  wire b1c778;
  wire b1c779;
  wire b1c77a;
  wire b1c77b;
  wire b1c77c;
  wire b1c77d;
  wire b1c77e;
  wire b1c77f;
  wire b1c780;
  wire b1c781;
  wire b1c782;
  wire b1c783;
  wire b1c784;
  wire b1c785;
  wire b1c786;
  wire b1c787;
  wire b1c788;
  wire b1c789;
  wire b1c78a;
  wire b1c78b;
  wire b1c78c;
  wire b1c78d;
  wire b1c78e;
  wire b1c78f;
  wire b1c790;
  wire b1c791;
  wire b1c792;
  wire b1c793;
  wire b1c794;
  wire b1c795;
  wire b1c796;
  wire b1c797;
  wire b1c798;
  wire b1c799;
  wire b1c79a;
  wire b1c79b;
  wire b1c79c;
  wire b1c79d;
  wire b1c79e;
  wire b1c79f;
  wire b1c7a0;
  wire b1c7a1;
  wire b1c7a2;
  wire b1c7a3;
  wire b1c7a4;
  wire b1c7a5;
  wire b1c7a6;
  wire b1c7a7;
  wire b1c7a8;
  wire b1c7a9;
  wire b1c7aa;
  wire b1c7ab;
  wire b1c7ac;
  wire b1c7ad;
  wire b1c7ae;
  wire b1c7af;
  wire b1c7b0;
  wire b1c7b1;
  wire b1c7b2;
  wire b1c7b3;
  wire b1c7b4;
  wire b1c7b5;
  wire b1c7b6;
  wire b1c7b7;
  wire b1c7b8;
  wire b1c7b9;
  wire b1c7ba;
  wire b1c7bb;
  wire b1c7bc;
  wire b1c7bd;
  wire b1c7be;
  wire b1c7bf;
  wire b1c7c0;
  wire b1c7c1;
  wire b1c7c2;
  wire b1c7c3;
  wire b1c7c4;
  wire b1c7c5;
  wire b1c7c6;
  wire b1c7c7;
  wire b1c7c8;
  wire b1c7c9;
  wire b1c7ca;
  wire b1c7cb;
  wire b1c7cc;
  wire b1c7cd;
  wire b1c7ce;
  wire b1c7cf;
  wire b1c7d0;
  wire b1c7d1;
  wire b1c7d2;
  wire b1c7d3;
  wire b1c7d4;
  wire b1c7d5;
  wire b1c7d6;
  wire b1c7d7;
  wire b1c7d8;
  wire b1c7d9;
  wire b1c7da;
  wire b1c7db;
  wire b1c7dc;
  wire b1c7dd;
  wire b1c7de;
  wire b1c7df;
  wire b1c7e0;
  wire b1c7e1;
  wire b1c7e2;
  wire b1c7e3;
  wire b1c7e4;
  wire b1c7e5;
  wire b1c7e6;
  wire b1c7e7;
  wire b1c7e8;
  wire b1c7e9;
  wire b1c7ea;
  wire b1c7eb;
  wire b1c7ec;
  wire b1c7ed;
  wire b1c7ee;
  wire b1c7ef;
  wire b1c7f0;
  wire b1c7f1;
  wire b1c7f2;
  wire b1c7f3;
  wire b1c7f4;
  wire b1c7f5;
  wire b1c7f6;
  wire b1c7f7;
  wire b1c7f8;
  wire b1c7f9;
  wire b1c7fa;
  wire b1c7fc;
  wire b1c7fd;
  wire b1c7fe;
  wire b1c7ff;
  wire b1c800;
  wire b1c801;
  wire b1c802;
  wire b1c803;
  wire b1c804;
  wire b1c805;
  wire b1c806;
  wire b1c807;
  wire b1c808;
  wire b1c809;
  wire b1c80a;
  wire b1c80b;
  wire b1c80c;
  wire b1c80d;
  wire b1c80e;
  wire b1c80f;
  wire b1c81b;
  wire b1c81c;
  wire b1c81d;
  wire b1c81e;
  wire b1c81f;
  wire b1c820;
  wire b1c821;
  wire b1c822;
  wire b1c823;
  wire b1c824;
  wire b1c825;
  wire b1c826;
  wire b1c827;
  wire b1c828;
  wire b1c829;
  wire b1c02d;
  wire b1c02e;
  wire b1c02f;
  wire b1c030;
  wire b1c031;
  wire b1c032;
  wire b1c033;
  wire b1c034;
  wire b1c035;
  wire b1c036;
  wire b1c037;
  wire b1c038;
  wire b1c039;
  wire b1c03a;
  wire b1c03b;
  wire b1c03c;
  wire b1c03d;
  wire b1c03e;
  wire b1c03f;
  wire b1c040;
  wire b1c041;
  wire b1c042;
  wire b1c043;
  wire b1c044;
  wire b1c045;
  wire b1c046;
  wire b1c047;
  wire b1c048;
  wire b1c049;
  wire b1c04a;
  wire b1c04b;
  wire b1c04c;
  wire b1c04d;
  wire b1c04e;
  wire b1c04f;
  wire b1c050;
  wire b1c051;
  wire b1c052;
  wire b1c053;
  wire b1c054;
  wire b1c055;
  wire b1c056;
  wire b1c057;
  wire b1c058;
  wire b1c059;
  wire b1c05a;
  wire b1c05b;
  wire b1c05c;
  wire b1c05d;
  wire b1c05e;
  wire b1c05f;
  wire b1c060;
  wire b1c061;
  wire b1c062;
  wire b1c063;
  wire b1c064;
  wire b1c065;
  wire b1c066;
  wire b1c067;
  wire b1c068;
  wire b1c069;
  wire b1c06a;
  wire b1c06b;
  wire b1c06c;
  wire b1c06d;
  wire b1c06e;
  wire b1c06f;
  wire b1c070;
  wire b1c071;
  wire b1c072;
  wire b1c073;
  wire b1c074;
  wire b1c075;
  wire b1c076;
  wire b1c077;
  wire b1c078;
  wire b1c079;
  wire b1c07a;
  wire b1c07b;
  wire b1c07c;
  wire b1c07d;
  wire b1c07e;
  wire b1c07f;
  wire b1c080;
  wire b1c081;
  wire b1c082;
  wire b1c083;
  wire b1c084;
  wire b1c085;
  wire b1c086;
  wire b1c087;
  wire b1c088;
  wire b1c089;
  wire b1c08a;
  wire b1c08b;
  wire b1c08c;
  wire b1c08d;
  wire b1c08e;
  wire b1c08f;
  wire b1c090;
  wire b1c091;
  wire b1c092;
  wire b1c093;
  wire b1c094;
  wire b1c095;
  wire b1c096;
  wire b1c097;
  wire b1c098;
  wire b1c0a6;
  wire b1c0a7;
  wire b1c0a8;
  wire b1c0a9;
  wire b1c0aa;
  wire b1c0ab;
  wire b1c0ac;
  wire b1c0b0;
  wire b1c0b1;
  wire b1c0b2;
  wire b1c0b3;
  wire b1c0b4;
  wire b1c0b5;
  wire b0589e;
  wire b0589f;
  wire b058a0;
  wire b058a1;
  wire b058a2;
  wire b058a3;
  wire b058a4;
  wire b058a5;
  wire b058a6;
  wire b058a7;
  wire b058a8;
  wire b058a9;
  wire b058aa;
  wire b058ab;
  wire b058ac;
  wire b058ad;
  wire b058ae;
  wire b058af;
  wire b058b0;
  wire b058b1;
  wire b058b2;
  wire b058b3;
  wire b058b4;
  wire b058b5;
  wire b058b6;
  wire b058b7;
  wire b058b8;
  wire b058b9;
  wire b058ba;
  wire b058bb;
  wire b058bc;
  wire b058bd;
  wire b058be;
  wire b058c1;
  wire b058c2;
  wire b058c3;
  wire b058c4;
  wire b058c5;
  wire b058c6;
  wire b058c7;
  wire b058c8;
  wire b058c9;
  wire b058ca;
  wire b058cb;
  wire b058cc;
  wire b058cd;
  wire b058ce;
  wire b058cf;
  wire b058d0;
  wire b058d1;
  wire b058d2;
  wire b058d3;
  wire b058d4;
  wire b058d5;
  wire b058d6;
  wire b058d7;
  wire b058d8;
  wire b058d9;
  wire b058da;
  wire b058db;
  wire b058dc;
  wire b058dd;
  wire b058de;
  wire b058df;
  wire b058e0;
  wire b058e1;
  wire b058e2;
  wire b058e3;
  wire b058e4;
  wire b058e5;
  wire b058e6;
  wire b058e7;
  wire b058e8;
  wire b058e9;
  wire b058ea;
  wire b058eb;
  wire b058ec;
  wire b058ed;
  wire b058ee;
  wire b058ef;
  wire b058f0;
  wire b058f1;
  wire b058f2;
  wire b058f3;
  wire b058f5;
  wire b058f6;
  wire b058f7;
  wire b058f8;
  wire b058f9;
  wire b058fa;
  wire b058fb;
  wire b058fc;
  wire b058fd;
  wire b058fe;
  wire b058ff;
  wire b05900;
  wire b05901;
  wire b05902;
  wire b05903;
  wire b05904;
  wire b05905;
  wire b05906;
  wire b05907;
  wire b05908;
  wire b05909;
  wire b0590a;
  wire b0590b;
  wire b0590c;
  wire b0590d;
  wire b0590e;
  wire b0590f;
  wire b05910;
  wire b05911;
  wire b05912;
  wire b05913;
  wire b05914;
  wire b05915;
  wire b05916;
  wire b05917;
  wire b05918;
  wire b0591b;
  wire b0591c;
  wire b0591d;
  wire b0591e;
  wire b0591f;
  wire b05920;
  wire b05921;
  wire b05922;
  wire b05923;
  wire b05924;
  wire b05925;
  wire b05926;
  wire b05927;
  wire b05928;
  wire b05929;
  wire b0592a;
  wire b0592b;
  wire b0592c;
  wire b0592d;
  wire b0592e;
  wire b0592f;
  wire b05930;
  wire b05931;
  wire b05932;
  wire b05933;
  wire b05934;
  wire b05935;
  wire b05936;
  wire b05937;
  wire b05938;
  wire b05939;
  wire b0593a;
  wire b0593b;
  wire b0593c;
  wire b0593d;
  wire b0593e;
  wire b0593f;
  wire b05940;
  wire b05941;
  wire b05942;
  wire b05943;
  wire b05944;
  wire b05945;
  wire b05946;
  wire b05947;
  wire b05948;
  wire b05949;
  wire b0594a;
  wire b0594b;
  wire b0594c;
  wire b0594d;
  wire b0594e;
  wire b0594f;
  wire b05950;
  wire b05951;
  wire b05952;
  wire b05953;
  wire b05954;
  wire b05955;
  wire b05956;
  wire b05957;
  wire b05958;
  wire b05959;
  wire b0595a;
  wire b0595b;
  wire b0595c;
  wire b0595d;
  wire b0595e;
  wire b0595f;
  wire b05960;
  wire b05961;
  wire b05962;
  wire b05963;
  wire b05964;
  wire b05965;
  wire b05966;
  wire b05967;
  wire b05968;
  wire b05969;
  wire b0596a;
  wire b0596b;
  wire b0596c;
  wire b0596d;
  wire b0596e;
  wire b0596f;
  wire b05970;
  wire b05971;
  wire b05972;
  wire b05973;
  wire b05974;
  wire b05975;
  wire b05976;
  wire b05977;
  wire b05978;
  wire b05979;
  wire b0597a;
  wire b0597b;
  wire b0597c;
  wire b0597d;
  wire b0597e;
  wire b0597f;
  wire b05980;
  wire b05981;
  wire b05982;
  wire b05983;
  wire b05984;
  wire b05985;
  wire b05986;
  wire b05987;
  wire b05988;
  wire b05989;
  wire b0598a;
  wire b0598b;
  wire b0598c;
  wire b0598d;
  wire b0598e;
  wire b0598f;
  wire b05990;
  wire b05991;
  wire b05992;
  wire b05993;
  wire b05994;
  wire b05995;
  wire b05996;
  wire b05997;
  wire b05998;
  wire b05999;
  wire b0599a;
  wire b0599b;
  wire b0599c;
  wire b0599d;
  wire b0599e;
  wire b0599f;
  wire b059a0;
  wire b059a1;
  wire b059a2;
  wire b059a3;
  wire b059a4;
  wire b059a5;
  wire b059a6;
  wire b059a7;
  wire b059a8;
  wire b059a9;
  wire b059aa;
  wire b059ab;
  wire b059ac;
  wire b059ad;
  wire b059ae;
  wire b059af;
  wire b059b0;
  wire b059b1;
  wire b059b2;
  wire b059b3;
  wire b059b4;
  wire b059b5;
  wire b059b6;
  wire b059b7;
  wire b059b8;
  wire b059b9;
  wire b059ba;
  wire b059bb;
  wire b059bc;
  wire b059bd;
  wire b059be;
  wire b059bf;
  wire b059c0;
  wire b059c1;
  wire b059c2;
  wire b059c3;
  wire b059c4;
  wire b059c5;
  wire b059c6;
  wire b059c7;
  wire b059c8;
  wire b059c9;
  wire b059ca;
  wire b059cb;
  wire b059cc;
  wire b059cd;
  wire b059ce;
  wire b059cf;
  wire b059d0;
  wire b059d1;
  wire b059d2;
  wire b059d3;
  wire b059d4;
  wire b059d5;
  wire b059d6;
  wire b059d7;
  wire b059d8;
  wire b059d9;
  wire b059da;
  wire b059db;
  wire b059dc;
  wire b059dd;
  wire b059de;
  wire b059df;
  wire b059e0;
  wire b059e1;
  wire b059e2;
  wire b059e3;
  wire b059e4;
  wire b059e5;
  wire b059e6;
  wire b059e7;
  wire b059e8;
  wire b059e9;
  wire b059ea;
  wire b059eb;
  wire b059ec;
  wire b059ed;
  wire b059ee;
  wire b059ef;
  wire b059f0;
  wire b059f1;
  wire b059f2;
  wire b059f3;
  wire b059f4;
  wire b059f5;
  wire b059f6;
  wire b059f7;
  wire b059f8;
  wire b059f9;
  wire b059fa;
  wire b059fb;
  wire b059fc;
  wire b059fd;
  wire b059fe;
  wire b059ff;
  wire b05a00;
  wire b05a01;
  wire b05a02;
  wire b05a03;
  wire b05a04;
  wire b05a05;
  wire b05a06;
  wire b05a07;
  wire b05a08;
  wire b05a09;
  wire b05a0a;
  wire b05a0b;
  wire b05a0c;
  wire b05a0d;
  wire b05a0e;
  wire b05a0f;
  wire b05a10;
  wire b05a11;
  wire b05a12;
  wire b05a13;
  wire b05a14;
  wire b05a15;
  wire b05a16;
  wire b05a17;
  wire b05a18;
  wire b05a19;
  wire b05a1a;
  wire b05a1b;
  wire b05a1c;
  wire b05a1d;
  wire b05a1e;
  wire b05a1f;
  wire b05a20;
  wire b05a21;
  wire b05a22;
  wire b05a23;
  wire b05a24;
  wire b05a25;
  wire b05a26;
  wire b05a27;
  wire b05a28;
  wire b05a29;
  wire b05a2a;
  wire b05a2b;
  wire b05a2c;
  wire b05a2d;
  wire b05a2e;
  wire b05a2f;
  wire b05a30;
  wire b05a31;
  wire b05a32;
  wire b05a33;
  wire b05a34;
  wire b05a35;
  wire b05a36;
  wire b05a37;
  wire b05a38;
  wire b05a39;
  wire b05a3a;
  wire b05a3b;
  wire b05a3c;
  wire b05a3d;
  wire b05a3e;
  wire b05a3f;
  wire b05a40;
  wire b05a41;
  wire b05a42;
  wire b05a43;
  wire b05a44;
  wire b05a45;
  wire b05a46;
  wire b05a47;
  wire b05a48;
  wire b05a49;
  wire b05a4a;
  wire b05a4b;
  wire b05a4c;
  wire b05a4d;
  wire b05a4e;
  wire b05a4f;
  wire b05a50;
  wire b05a51;
  wire b05a52;
  wire b05a53;
  wire b05a54;
  wire b05a55;
  wire b05a56;
  wire b05a57;
  wire b05a58;
  wire b05a59;
  wire b05a5a;
  wire b05a5b;
  wire b05a5c;
  wire b05a5d;
  wire b05a5e;
  wire b05a5f;
  wire b05a60;
  wire b05a61;
  wire b05a62;
  wire b05a63;
  wire b05a64;
  wire b05a65;
  wire b05a66;
  wire b05a67;
  wire b05a68;
  wire b05a69;
  wire b05a6a;
  wire b05a6b;
  wire b05a6c;
  wire b05a6d;
  wire b05a6e;
  wire b05a6f;
  wire b05a70;
  wire b05a71;
  wire b05a72;
  wire b05a73;
  wire b05a74;
  wire b05a75;
  wire b05a76;
  wire b05a77;
  wire b05a78;
  wire b05a79;
  wire b05a7a;
  wire b05a7b;
  wire b05a7c;
  wire b05a7d;
  wire b05a7e;
  wire b05a7f;
  wire b05a80;
  wire b05a81;
  wire b05a82;
  wire b05a83;
  wire b05a84;
  wire b05a85;
  wire b05a86;
  wire b05a87;
  wire b05a88;
  wire b05a89;
  wire b05a8a;
  wire b05a8b;
  wire b05a8c;
  wire b05a8d;
  wire b05a8e;
  wire b05a8f;
  wire b05a90;
  wire b05a91;
  wire b05a92;
  wire b05a93;
  wire b05a94;
  wire b05a95;
  wire b05a96;
  wire b05a97;
  wire b05a98;
  wire b05a99;
  wire b05a9a;
  wire b05a9b;
  wire b05a9c;
  wire v867d75;
  wire b05a9d;
  wire b05a9e;
  wire ac144e;
  wire ac144f;
  wire ac1450;
  wire ac1451;
  wire ac1452;
  wire ac1453;
  wire ac1454;
  wire ac1455;
  wire ac1456;
  wire ac1458;
  wire ac1459;
  wire ac145a;
  wire ac145b;
  wire ac145c;
  wire ac145d;
  wire ac145e;
  wire ac145f;
  wire ac1460;
  wire ac1461;
  wire ac1462;
  wire ac1463;
  wire ac1464;
  wire ac1465;
  wire ac1466;
  wire ac1467;
  wire ac1468;
  wire ac1469;
  wire ac146a;
  wire ac146b;
  wire ac146c;
  wire ac146d;
  wire ac146e;
  wire ac146f;
  wire ac1470;
  wire ac1472;
  wire ac1474;
  wire ac1475;
  wire ac1476;
  wire ac1477;
  wire ac1478;
  wire ac1479;
  wire ac147a;
  wire ac147b;
  wire ac147c;
  wire ac147d;
  wire ac147e;
  wire ac1480;
  wire ac1481;
  wire ac1482;
  wire ac1483;
  wire ac1484;
  wire ac1485;
  wire ac1486;
  wire ac1487;
  wire ac1488;
  wire ac1489;
  wire ac148a;
  wire ac148b;
  wire ac148c;
  wire ac148d;
  wire ac148e;
  wire ac148f;
  wire ac1490;
  wire ac1491;
  wire ac1492;
  wire ac1493;
  wire ac1494;
  wire ac1495;
  wire ad4d8e;
  wire ad4d8f;
  wire ad4d90;
  wire ad4d91;
  wire ad4d92;
  wire ad4d93;
  wire ad4d94;
  wire ad4d96;
  wire ad4d97;
  wire ad4d98;
  wire ad4d99;
  wire ad4d9a;
  wire ad4d9b;
  wire ad4d9c;
  wire ad4d9d;
  wire ad4d9e;
  wire ad4d9f;
  wire ad4da0;
  wire ad4da1;
  wire ad4da2;
  wire ad4da3;
  wire ad4da4;
  wire ad4da8;
  wire ad4da9;
  wire ad4daa;
  wire ad4dab;
  wire ad4dac;
  wire ad4dad;
  wire ad4dae;
  wire ad4daf;
  wire ad4db0;
  wire ad4db1;
  wire ad4db2;
  wire ad4db3;
  wire ad4db4;
  wire ad4db5;
  wire ad4db6;
  wire ad4db7;
  wire ad4db8;
  wire ad4db9;
  wire ad4dba;
  wire ad4dbc;
  wire ad4dbd;
  wire ad4dbe;
  wire ad4dbf;
  wire ad4dc0;
  wire ad4dc1;
  wire ad4dc2;
  wire ad4dc3;
  wire ad4dc4;
  wire ad4dc5;
  wire ad4dc6;
  wire ad4dc7;
  wire ad4dc8;
  wire ad4dc9;
  wire ad4dca;
  wire ad4dce;
  wire ad4dcf;
  wire ad4dd0;
  wire ad4dd1;
  wire ad4dd2;
  wire ad4dd3;
  wire ad4dd4;
  wire ad4dd5;
  wire ad4dd6;
  wire ad4dd7;
  wire ad4dd9;
  wire ad4dda;
  wire ad4ddb;
  wire ad4ddd;
  wire ad4dde;
  wire ad4ddf;
  wire ad4de0;
  wire ad4de1;
  wire ad4de2;
  wire ad4de3;
  wire ad4de4;
  wire ad4de5;
  wire ad4de6;
  wire ad4de7;
  wire ad4de8;
  wire ad4de9;
  wire ad4dea;
  wire ad4deb;
  wire ad4dec;
  wire ad4ded;
  wire ad4dee;
  wire ad4def;
  wire ad4df0;
  wire ad4df1;
  wire ad4df2;
  wire ad4df3;
  wire ad4df5;
  wire ad4df6;
  wire ad4df7;
  wire ad4df8;
  wire ad4e0b;
  wire ad4e1f;
  wire ad4e20;
  wire ad4e21;
  wire v845547;
  wire ad4e22;
  wire ad4e23;
  wire ad4e24;
  wire ad4e40;
  wire ad4e41;
  wire ad4e42;
  wire ad4e43;
  wire ad4e44;
  wire af7f59;
  wire af7f5a;
  wire ad4e45;
  wire ad4e46;
  wire ad4e47;
  wire ad4e48;
  wire ad4e49;
  wire ad4e4a;
  wire ad4e4b;
  wire ad4e4c;
  wire ad4e4d;
  wire ad4e4e;
  wire ad4e4f;
  wire ad4e50;
  wire ad4e51;
  wire ad4e52;
  wire ad4e53;
  wire ad4e54;
  wire ad4e55;
  wire ad4e56;
  wire ad4e57;
  wire ad4e58;
  wire ad4e59;
  wire ad4e5a;
  wire ad4e5b;
  wire ad4e5c;
  wire ad4e5d;
  wire ad4e5e;
  wire ad4e5f;
  wire ad4e60;
  wire ad4e61;
  wire ad4e62;
  wire ad4e64;
  wire ad4e65;
  wire ad4e66;
  wire ad4e67;
  wire ad4e68;
  wire ad4e69;
  wire ad4e6a;
  wire ad4e6b;
  wire ad4e6c;
  wire ad4e6d;
  wire ad4e6e;
  wire ad4e6f;
  wire ad4e70;
  wire ad4e71;
  wire ad4e72;
  wire ad4e73;
  wire ad4e74;
  wire ad4e75;
  wire ad4e76;
  wire ad4e77;
  wire ad4e78;
  wire ad4e79;
  wire ad4e7a;
  wire ad4e7b;
  wire ad4e7c;
  wire ad4e7d;
  wire ad4e7e;
  wire ad4e7f;
  wire ad4e80;
  wire ad4e81;
  wire ad4e82;
  wire ad4e83;
  wire ad4e84;
  wire ad4e85;
  wire ad4e86;
  wire ad4e87;
  wire ad4e88;
  wire ad4e89;
  wire ad4e8a;
  wire ad4e8b;
  wire ad4e8c;
  wire ad4e8d;
  wire ad4e8e;
  wire ad4e8f;
  wire ad4e90;
  wire ad4e91;
  wire ad4e92;
  wire ad4e93;
  wire ad4e94;
  wire ad4e95;
  wire ad4e96;
  wire ad4e97;
  wire ad4e98;
  wire ad4e99;
  wire ad4e9a;
  wire ad4e9b;
  wire ad4e9c;
  wire ad4e9d;
  wire ad4e9e;
  wire ad4e9f;
  wire ad4ea0;
  wire ad4ea1;
  wire ad4ea2;
  wire ad4ea3;
  wire ad4ea4;
  wire ad4ea5;
  wire ad4ea6;
  wire ad4ea7;
  wire ad4ea8;
  wire ad4ea9;
  wire ad4eaa;
  wire ad4eab;
  wire ad4eac;
  wire ad4ead;
  wire ad4eae;
  wire ad4eaf;
  wire ad4eb0;
  wire ad4eb1;
  wire ad4eb2;
  wire ad4eb3;
  wire ad4eb4;
  wire ad4eb5;
  wire ad4eb6;
  wire ad4eb7;
  wire ad4eb8;
  wire ad4eb9;
  wire ad4eba;
  wire ad4ebb;
  wire ad4ebc;
  wire ad4ebd;
  wire ad4ebe;
  wire ad4ebf;
  wire ad4ec0;
  wire ad4ec1;
  wire ad4ec2;
  wire ad4ec3;
  wire ad4ec4;
  wire ad4ec5;
  wire ad4ec6;
  wire ad4ec7;
  wire ad4ec8;
  wire ad4ec9;
  wire ad4eca;
  wire ad4ecb;
  wire ad4ecc;
  wire ad4ecd;
  wire ad4ece;
  wire ad4ecf;
  wire ad4ed0;
  wire ad4ed1;
  wire ad4ed2;
  wire ad4ed3;
  wire ad4ed4;
  wire ad4ed5;
  wire ad4ed6;
  wire ad4ed7;
  wire ad4ed8;
  wire ad4ed9;
  wire ad4eda;
  wire ad4edb;
  wire ad4edc;
  wire ad4edd;
  wire ad4ede;
  wire ad4edf;
  wire ad4ee0;
  wire ad4ee1;
  wire ad4ee2;
  wire ad4ee3;
  wire ad4ee4;
  wire ad4ee5;
  wire ad4ee6;
  wire ad4ee7;
  wire ad4ee8;
  wire ad4ee9;
  wire ad4eea;
  wire ad4eeb;
  wire ad4eec;
  wire ad4eed;
  wire ad4eee;
  wire ad4eef;
  wire ad4ef0;
  wire ad4ef1;
  wire ad4ef2;
  wire ad4ef3;
  wire ad4ef4;
  wire ad4ef5;
  wire ad4ef6;
  wire ad4ef7;
  wire ad4ef8;
  wire ad4ef9;
  wire ad4efa;
  wire ad4efb;
  wire ad4efc;
  wire ad4efd;
  wire ad4efe;
  wire ad4eff;
  wire ad4f00;
  wire ad4f01;
  wire ad4f02;
  wire ad4f03;
  wire ad4f04;
  wire ad4f05;
  wire ad4f06;
  wire ad4f07;
  wire ad4f08;
  wire ad4f09;
  wire ad4f0a;
  wire ad4f0b;
  wire ad4f0c;
  wire ad4f0d;
  wire ad4f0e;
  wire ad4f0f;
  wire ad4f10;
  wire ad4f11;
  wire ad4f12;
  wire ad4f13;
  wire ad4f14;
  wire ad4f15;
  wire ad4f16;
  wire ad4f17;
  wire ad4f18;
  wire ad4f19;
  wire ad4f1a;
  wire ad4f1b;
  wire ad4f1c;
  wire ad4f1d;
  wire ad4f1e;
  wire ad4f1f;
  wire ad4f20;
  wire ad4f21;
  wire ad4f22;
  wire ad4f23;
  wire ad4f24;
  wire ad4f25;
  wire ad4f26;
  wire ad4f27;
  wire ad4f28;
  wire ad4f2a;
  wire ad4f2b;
  wire ad4f2c;
  wire ad4f2d;
  wire ad4f2e;
  wire ad4f2f;
  wire ad4f30;
  wire ad4f31;
  wire ad4f32;
  wire ad4f33;
  wire v8b08c2;
  wire ad4f34;
  wire ad4f35;
  wire ad4f36;
  wire ad4f37;
  wire ad4f38;
  wire ad4f39;
  wire ad4f3a;
  wire ad4f3b;
  wire ad4f3c;
  wire ad4f3d;
  wire ad4f3e;
  wire ad4f3f;
  wire ad4f40;
  wire ad4f41;
  wire ad4f42;
  wire ad4f43;
  wire ad4f44;
  wire ad4f45;
  wire ad4f46;
  wire ad4f47;
  wire ad4f48;
  wire ad4f49;
  wire ad4f4a;
  wire ad4f4b;
  wire ad4f4c;
  wire ad4f4d;
  wire ad4f4e;
  wire ad4f4f;
  wire ad4f50;
  wire ad4f52;
  wire ad4f53;
  wire ad4f54;
  wire ad4f55;
  wire ad4f56;
  wire ad4f57;
  wire ad4f58;
  wire ad4f59;
  wire ad4f5a;
  wire ad4f5b;
  wire ad4f5c;
  wire ad4f5d;
  wire ad4f5e;
  wire ad4f5f;
  wire ad4f60;
  wire ad4f61;
  wire ad4f62;
  wire ad4f63;
  wire ad4f64;
  wire ad4f65;
  wire ad4f66;
  wire ad4f67;
  wire ad4f68;
  wire ad4f69;
  wire ad4f6a;
  wire ad4f6b;
  wire ad4f6c;
  wire ad4f6d;
  wire ad4f6e;
  wire ad4f6f;
  wire ad4f70;
  wire ad4f71;
  wire ad4f72;
  wire ad4f73;
  wire ad4f74;
  wire ad4f75;
  wire ad4f76;
  wire ad4f77;
  wire ad4f78;
  wire ad4f79;
  wire ad4f7a;
  wire ad4f7b;
  wire ad4f7c;
  wire ad4f7d;
  wire ad4f7e;
  wire ad4f7f;
  wire ad4f80;
  wire ad4f81;
  wire ad4f82;
  wire ad4f83;
  wire ad4f84;
  wire ad4f85;
  wire ad4f86;
  wire ad4f87;
  wire ad4f88;
  wire ad4f89;
  wire ad4f8a;
  wire ad4f8b;
  wire ad4f8c;
  wire ad4f8d;
  wire ad4f8e;
  wire ad4f8f;
  wire ad4f90;
  wire ad4f91;
  wire ad4f92;
  wire ad4f93;
  wire ad4f94;
  wire ad4f95;
  wire ad4f96;
  wire ad4f97;
  wire ad4f98;
  wire ad4f99;
  wire ad4f9a;
  wire ad4f9b;
  wire ad4f9c;
  wire ad4f9d;
  wire ad4f9e;
  wire ad4f9f;
  wire ad4fa0;
  wire ad4fa1;
  wire ad4fa2;
  wire ad4fa4;
  wire ad4fa5;
  wire ad4fa6;
  wire ad4fa7;
  wire ad4fa8;
  wire ad4fa9;
  wire ad4faa;
  wire c76645;
  wire c73a9a;
  wire c76647;
  wire e199ba;
  wire ad4fab;
  wire ad4fac;
  wire ad4fad;
  wire ad4fae;
  wire ad4faf;
  wire ad4fb0;
  wire ad4fb1;
  wire ad4fb2;
  wire ad4fb3;
  wire ad4fb4;
  wire ad4fb5;
  wire ad4fb6;
  wire ad4fb7;
  wire ad4fb8;
  wire ad4fb9;
  wire ad4fbb;
  wire ad4fbc;
  wire ad4fbd;
  wire ad4fbe;
  wire ad4fbf;
  wire ad4fc0;
  wire ad4fc1;
  wire ad4fc2;
  wire ad4fc3;
  wire ad4fc4;
  wire ad4fc5;
  wire ad4fc6;
  wire ad4fc7;
  wire ad4fc8;
  wire ad4fc9;
  wire ad4fca;
  wire ad4fcb;
  wire ad4fcc;
  wire ad4fcd;
  wire ad4fce;
  wire ad4fcf;
  wire ad4fd0;
  wire ad4fd1;
  wire ad4fd2;
  wire ad4fd3;
  wire ad4fd4;
  wire ad4fd5;
  wire ad4fd6;
  wire ad4fd7;
  wire ad4fd8;
  wire ad4fd9;
  wire ad4fda;
  wire ad4fdb;
  wire ad4fdc;
  wire ad4fdd;
  wire ad4fde;
  wire ad4fdf;
  wire ad4fe0;
  wire ad4fe1;
  wire ad4fe2;
  wire ad4fe3;
  wire ad4fe4;
  wire ad4fe5;
  wire ad4fe6;
  wire ad4fe7;
  wire ad4fe8;
  wire ad4fe9;
  wire ad4fea;
  wire ad4feb;
  wire ad4fec;
  wire ad4fed;
  wire ad4fee;
  wire ad4fef;
  wire ad4ff0;
  wire ad4ff1;
  wire ad4ff2;
  wire ad4ff3;
  wire ad4ff5;
  wire ad4ff6;
  wire ad4ff7;
  wire ad4ff8;
  wire ad4ff9;
  wire ad4ffa;
  wire ad4ffb;
  wire ad5012;
  wire ad5013;
  wire ad5014;
  wire ad5015;
  wire ad5016;
  wire ad5017;
  wire ad5018;
  wire ad5019;
  wire ad501a;
  wire ad501b;
  wire ad501c;
  wire ad501d;
  wire ad501e;
  wire ad501f;
  wire ad5021;
  wire ad5022;
  wire ad5023;
  wire ad5024;
  wire ad5025;
  wire ad5026;
  wire ad5027;
  wire ad5028;
  wire ad5029;
  wire ad502a;
  wire ad502b;
  wire ad502c;
  wire ad502d;
  wire ad502e;
  wire ad502f;
  wire ad5030;
  wire ad5031;
  wire ad5032;
  wire ad5033;
  wire ad5034;
  wire ad5035;
  wire ad5036;
  wire ad5037;
  wire ad5038;
  wire ad5039;
  wire ad503a;
  wire ad503b;
  wire ad503c;
  wire ad503d;
  wire ad503e;
  wire ad503f;
  wire ad5040;
  wire ad5041;
  wire ad5042;
  wire ad5043;
  wire ad5044;
  wire ad5045;
  wire ad5046;
  wire ad5047;
  wire ad5048;
  wire ad5049;
  wire ad504a;
  wire ad504b;
  wire ad504c;
  wire ad504d;
  wire ad504e;
  wire ad504f;
  wire ad5050;
  wire ad5051;
  wire ad5052;
  wire ad5053;
  wire ad5054;
  wire ad5055;
  wire ad5056;
  wire ad5057;
  wire ad5058;
  wire ad5059;
  wire ad505a;
  wire ad505b;
  wire ad505d;
  wire ad505e;
  wire ad505f;
  wire ad5060;
  wire ad5061;
  wire ad5062;
  wire ad5063;
  wire ad5064;
  wire ad5065;
  wire ad5066;
  wire ad5067;
  wire ad5068;
  wire ad5069;
  wire ad506a;
  wire ad506b;
  wire ad506d;
  wire ad506e;
  wire ad506f;
  wire ad5070;
  wire ad5071;
  wire ad508d;
  wire ad508e;
  wire ad508f;
  wire ad5090;
  wire ad48c5;
  wire ad48c6;
  wire ad48c7;
  wire ad48c8;
  wire ad48c9;
  wire ad48ca;
  wire ad48cb;
  wire ad4554;
  wire ad4555;
  wire ad4556;
  wire ad4557;
  wire ad4558;
  wire ad4559;
  wire ad455a;
  wire ad455b;
  wire ad455c;
  wire ad455d;
  wire ad455e;
  wire ad455f;
  wire ad4560;
  wire ad4561;
  wire ad4562;
  wire ad4563;
  wire ad4564;
  wire ad4565;
  wire ad4566;
  wire ad4567;
  wire ad4568;
  wire ad4569;
  wire ad456a;
  wire ad456b;
  wire ad456c;
  wire ad456d;
  wire ad456e;
  wire ad456f;
  wire ad4570;
  wire ad4571;
  wire ad4572;
  wire ad4573;
  wire ad4574;
  wire ad4575;
  wire ad4576;
  wire ad4577;
  wire ad4578;
  wire ad4579;
  wire ad457a;
  wire ad457b;
  wire ad457c;
  wire ad457d;
  wire ad457e;
  wire ad457f;
  wire ad4580;
  wire ad4581;
  wire ad4582;
  wire ad4583;
  wire ad4584;
  wire ad4585;
  wire ad4586;
  wire ad4587;
  wire ad4588;
  wire ad4589;
  wire ad458a;
  wire ad458b;
  wire ad458c;
  wire ad458d;
  wire ad458e;
  wire ad458f;
  wire ad4590;
  wire ad4591;
  wire ad4592;
  wire ad4593;
  wire ad4594;
  wire ad4595;
  wire ad4596;
  wire ad4597;
  wire ad4598;
  wire ad4599;
  wire ad459a;
  wire ad459b;
  wire ad459c;
  wire ad459d;
  wire ad459e;
  wire ad459f;
  wire ad45a0;
  wire ad45a1;
  wire ad45a2;
  wire ad45a3;
  wire ad45a4;
  wire ad45a5;
  wire ad45a6;
  wire ad45a7;
  wire ad45a8;
  wire ad45a9;
  wire ad45aa;
  wire ad45ab;
  wire ad45ac;
  wire ad45ad;
  wire ad45ae;
  wire ad45af;
  wire ad45b0;
  wire ad45b1;
  wire ad45b2;
  wire ad45b3;
  wire ad45b4;
  wire ad45b5;
  wire ad45b6;
  wire ad45b7;
  wire ad45b8;
  wire ad45b9;
  wire ad45ba;
  wire ad45bb;
  wire ad45bc;
  wire ad45bd;
  wire ad45be;
  wire ad45bf;
  wire ad45c0;
  wire ad45c1;
  wire ad45c2;
  wire ad45c3;
  wire ad45c4;
  wire ad45c5;
  wire ad45c6;
  wire ad45c7;
  wire ad45c8;
  wire ad45c9;
  wire ad45ca;
  wire ad45cb;
  wire ad45cc;
  wire ad45df;
  wire ad45e0;
  wire ad45e1;
  wire ad45e2;
  wire ad45e3;
  wire ad45e4;
  wire ad45e5;
  wire ad45e6;
  wire ad45e7;
  wire ad45e8;
  wire ad45e9;
  wire ad45ea;
  wire ad45eb;
  wire ad45ec;
  wire ad45ed;
  wire ad45ee;
  wire ad45ef;
  wire ad45f0;
  wire ad45f1;
  wire ad45f2;
  wire ad45f3;
  wire ad45f4;
  wire ad45f8;
  wire ad45f9;
  wire ad45fa;
  wire ad45fb;
  wire ad45fc;
  wire ad45fd;
  wire ad45fe;
  wire ad45ff;
  wire ad4600;
  wire ad4601;
  wire ad4602;
  wire ad4603;
  wire ad4604;
  wire ad4605;
  wire ad4606;
  wire ad4607;
  wire ad4608;
  wire ad4609;
  wire ad460a;
  wire ad460b;
  wire ad460c;
  wire ad460d;
  wire ad460e;
  wire ad460f;
  wire ad4610;
  wire ad4611;
  wire ad4687;
  wire ad4688;
  wire ad4689;
  wire ad468a;
  wire ad468b;
  wire ad468c;
  wire ad468d;
  wire ad468e;
  wire ad468f;
  wire ad4690;
  wire ad4691;
  wire ad4692;
  wire ad4693;
  wire ad4694;
  wire ad4695;
  wire ad4696;
  wire ad4697;
  wire ad4698;
  wire ad4699;
  wire ad469a;
  wire ad469b;
  wire ad469c;
  wire ad469d;
  wire ad469e;
  wire ad469f;
  wire ad46a0;
  wire ad46a1;
  wire ad46a2;
  wire ad46a3;
  wire ad46a4;
  wire ad46a5;
  wire ad46a6;
  wire ad46a7;
  wire ad46a8;
  wire ad46a9;
  wire ad46aa;
  wire ad46ab;
  wire ad46ac;
  wire ad46ad;
  wire ad46ae;
  wire ad46af;
  wire ad46b0;
  wire ad46b1;
  wire ad46b2;
  wire ad46b3;
  wire ad46b4;
  wire ad46b5;
  wire ad46b6;
  wire ad46b7;
  wire ad46b8;
  wire ad46b9;
  wire ad46ba;
  wire ad46bb;
  wire ad46bc;
  wire ad46bd;
  wire ad46be;
  wire ad46bf;
  wire ad46c0;
  wire ad46c1;
  wire ad46c2;
  wire ad46c3;
  wire ad46c4;
  wire ad46c5;
  wire ad46c6;
  wire ad46c7;
  wire ad46c8;
  wire ad46c9;
  wire ad46ca;
  wire ad46cb;
  wire ad46cc;
  wire ad46cd;
  wire ad46ce;
  wire ad46cf;
  wire ad46d0;
  wire ad46d1;
  wire ad46d2;
  wire ad46d3;
  wire ad46d4;
  wire ad46d5;
  wire ad46d6;
  wire ad46d7;
  wire ad46d8;
  wire ad46d9;
  wire ad46da;
  wire ad46db;
  wire ad46dc;
  wire ad46dd;
  wire ad46de;
  wire ad46df;
  wire ad46e0;
  wire ad46e1;
  wire ad46e2;
  wire ad46e3;
  wire ad46e4;
  wire ad46e5;
  wire ad46e6;
  wire ad46e7;
  wire ad46e8;
  wire ad46e9;
  wire ad46ea;
  wire ad46eb;
  wire ad46ec;
  wire ad46ed;
  wire ad46ee;
  wire ad46ef;
  wire ad46f0;
  wire ad46f1;
  wire ad46f2;
  wire ad46f3;
  wire ad46f4;
  wire ad46f5;
  wire ad46f6;
  wire ad46f7;
  wire ad46f8;
  wire ad46f9;
  wire ad46fa;
  wire ad46fb;
  wire ad46fc;
  wire ad46fd;
  wire ad46fe;
  wire ad46ff;
  wire ad4700;
  wire ad4701;
  wire ad4702;
  wire ad4703;
  wire ad4704;
  wire ad4705;
  wire ad4706;
  wire ad4707;
  wire ad4708;
  wire ad4709;
  wire ad470a;
  wire ad470b;
  wire ad470c;
  wire ad470d;
  wire ad470e;
  wire ad470f;
  wire ad4710;
  wire ad4711;
  wire ad4712;
  wire ad4713;
  wire ad4714;
  wire ad4715;
  wire ad4716;
  wire ad4717;
  wire ad4718;
  wire ad4719;
  wire ad471a;
  wire ad471b;
  wire ad471c;
  wire ad471d;
  wire ad471e;
  wire ad471f;
  wire ad4720;
  wire ad4721;
  wire ad4722;
  wire ad4723;
  wire ad4724;
  wire ad4725;
  wire ad472c;
  wire ad472d;
  wire ad472e;
  wire ad472f;
  wire ad4730;
  wire ad4731;
  wire ad4732;
  wire ad4733;
  wire ad4734;
  wire ad4735;
  wire ad4736;
  wire ad4737;
  wire ad4738;
  wire ad4739;
  wire ad473a;
  wire ad473b;
  wire ad473c;
  wire ad473d;
  wire ad473e;
  wire ad473f;
  wire ad4740;
  wire ad4741;
  wire ad4742;
  wire ad4743;
  wire ad4744;
  wire ad4745;
  wire ad4746;
  wire ad4747;
  wire ad4748;
  wire ad4749;
  wire ad474a;
  wire ad474b;
  wire ad474c;
  wire ad474d;
  wire ad474e;
  wire ad474f;
  wire ad4750;
  wire ad4751;
  wire ad4752;
  wire ad4753;
  wire ad4754;
  wire ad4755;
  wire ad4756;
  wire ad4757;
  wire ad4758;
  wire ad4759;
  wire ad475a;
  wire ad475b;
  wire ad475c;
  wire ad475d;
  wire ad475e;
  wire ad475f;
  wire ad4760;
  wire ad4761;
  wire ad4762;
  wire ad4763;
  wire ad4764;
  wire ad4765;
  wire ad4766;
  wire ad4767;
  wire ad4768;
  wire ad4769;
  wire ad476a;
  wire ad476b;
  wire ad476c;
  wire ad476d;
  wire ad476e;
  wire ad476f;
  wire ad4770;
  wire ad4774;
  wire ad4775;
  wire ad4776;
  wire ad4777;
  wire ad4778;
  wire ad4779;
  wire ad477a;
  wire ad477b;
  wire ad477c;
  wire ad477d;
  wire ad4781;
  wire ad4782;
  wire ad4783;
  wire ad4784;
  wire ad4785;
  wire ad4786;
  wire ad4787;
  wire ad4788;
  wire ad4789;
  wire ad47e8;
  wire ad47e9;
  wire ad47ea;
  wire ad47eb;
  wire ad47ec;
  wire ad47ed;
  wire ad47ee;
  wire ad47ef;
  wire ad47f0;
  wire ad47f1;
  wire ad47f2;
  wire ad47f3;
  wire ad47f4;
  wire ad47f5;
  wire ad47f6;
  wire ad47f7;
  wire ad47f8;
  wire ad47f9;
  wire ad47fa;
  wire ad47fb;
  wire ad47fc;
  wire ad47fd;
  wire ad47fe;
  wire ad47ff;
  wire ad4800;
  wire ad4801;
  wire ad4802;
  wire ad4803;
  wire ad4804;
  wire ad4805;
  wire ad4806;
  wire ad4807;
  wire ad4808;
  wire ad4809;
  wire ad480a;
  wire ad480b;
  wire ad480c;
  wire ad480d;
  wire ad480e;
  wire ad480f;
  wire ad4810;
  wire ad4811;
  wire ad4812;
  wire ad4813;
  wire ad4814;
  wire ad4815;
  wire ad4816;
  wire ad4817;
  wire ad4818;
  wire ad4819;
  wire ad481a;
  wire ad481b;
  wire ad481c;
  wire ad481d;
  wire ad481e;
  wire ad481f;
  wire ad4820;
  wire ad4821;
  wire ad4822;
  wire ad4823;
  wire ad4824;
  wire ad4825;
  wire ad4826;
  wire ad4827;
  wire ad4828;
  wire ad4844;
  wire ad4845;
  wire ad4846;
  wire ad4847;
  wire ad4848;
  wire ad4849;
  wire ad484a;
  wire ad484b;
  wire ad484c;
  wire ad484d;
  wire ad484e;
  wire ad484f;
  wire ad4850;
  wire ad4851;
  wire ad4894;
  wire ad4895;
  wire ad4896;
  wire ad4897;
  wire ad4898;
  wire ad48a5;
  wire ad48a6;
  wire ad48b0;
  wire ad48b1;
  wire ad48b2;
  wire ad48b3;
  wire ad48b4;
  wire ad48b5;
  wire ad48b6;
  wire ad48b7;
  wire ad40ba;
  wire ad40e6;
  wire ad40e7;
  wire ad40e8;
  wire ad40e9;
  wire ad40ea;
  wire ad40eb;
  wire ad40ec;
  wire ad40ed;
  wire ad40ee;
  wire ad40ef;
  wire ad40f0;
  wire ad40f1;
  wire ad40f2;
  wire ad40f3;
  wire ad40f4;
  wire ad40f5;
  wire ad40f6;
  wire ad40f7;
  wire ad40f8;
  wire ad40fa;
  wire ad40fb;
  wire ad40fc;
  wire ad40fd;
  wire ad40fe;
  wire ad40ff;
  wire ad4100;
  wire ad4101;
  wire ad4102;
  wire ad4103;
  wire ad4104;
  wire ad4105;
  wire ad4106;
  wire ad4107;
  wire ad4108;
  wire ad4109;
  wire ad410a;
  wire ad410b;
  wire ad410c;
  wire ad410d;
  wire ad410e;
  wire ad410f;
  wire ad4110;
  wire ad4111;
  wire ad4131;
  wire ad4132;
  wire ad4133;
  wire ad4134;
  wire ad4135;
  wire ad4136;
  wire ad4137;
  wire ad4138;
  wire ad4139;
  wire ad413a;
  wire ad413b;
  wire ad413c;
  wire ad413d;
  wire ad413e;
  wire ad413f;
  wire ad4140;
  wire ad4141;
  wire ad4142;
  wire ad4143;
  wire ad4144;
  wire ad4145;
  wire ad4146;
  wire ad4147;
  wire ad4148;
  wire ad4149;
  wire ad414a;
  wire ad414b;
  wire ad414c;
  wire ad414d;
  wire ad414e;
  wire ad414f;
  wire ad4150;
  wire ad4151;
  wire ad4152;
  wire ad4153;
  wire ad4154;
  wire ad4155;
  wire ad4156;
  wire ad4157;
  wire ad4158;
  wire ad4159;
  wire ad415a;
  wire ad415b;
  wire ad415c;
  wire ad415d;
  wire ad415e;
  wire ad415f;
  wire ad4160;
  wire ad4161;
  wire ad4162;
  wire ad4163;
  wire ad4164;
  wire ad4165;
  wire ad4166;
  wire ad4167;
  wire ad4168;
  wire ad4169;
  wire ad416a;
  wire ad416b;
  wire ad416c;
  wire ad416d;
  wire ad416e;
  wire ad416f;
  wire ad419d;
  wire ad419e;
  wire ad419f;
  wire ad41a0;
  wire ad41a1;
  wire ad41a2;
  wire ad41a3;
  wire ad41a4;
  wire ad41a5;
  wire ad41a6;
  wire ad41a7;
  wire ad41a8;
  wire ad41a9;
  wire ad41ab;
  wire ad41ac;
  wire ad41ad;
  wire ad41ae;
  wire ad41af;
  wire ad41b0;
  wire ad41b1;
  wire ad41b2;
  wire ad41b3;
  wire ad41b4;
  wire ad41b5;
  wire ad41b6;
  wire ad41b7;
  wire ad41b8;
  wire ad41b9;
  wire ad4257;
  wire ad4258;
  wire ad4259;
  wire ad425a;
  wire ad425b;
  wire ad425c;
  wire ad425e;
  wire ad425f;
  wire ad4260;
  wire ad4261;
  wire ad4262;
  wire ad4263;
  wire ad4264;
  wire ad4265;
  wire ad4266;
  wire ad4267;
  wire ad4268;
  wire ad4269;
  wire ad426a;
  wire ad426b;
  wire ad426c;
  wire ad426d;
  wire ad426e;
  wire ad426f;
  wire ad4270;
  wire ad4271;
  wire ad4272;
  wire ad4273;
  wire ad4274;
  wire ad4275;
  wire ad4276;
  wire ad4277;
  wire ad4278;
  wire ad4279;
  wire ad427a;
  wire ad427b;
  wire ad427c;
  wire ad427d;
  wire ad427e;
  wire ad427f;
  wire ad4280;
  wire ad4281;
  wire ad4282;
  wire ad4283;
  wire ad4284;
  wire ad4285;
  wire ad4286;
  wire ad4287;
  wire ad4288;
  wire ad4289;
  wire ad428a;
  wire ad428b;
  wire ad428c;
  wire ad428d;
  wire ad428e;
  wire ad428f;
  wire ad4290;
  wire ad4291;
  wire ad4292;
  wire ad4293;
  wire ad4294;
  wire ad4295;
  wire ad4296;
  wire ad4297;
  wire ad4298;
  wire ad4299;
  wire ad429a;
  wire ad429b;
  wire ad429c;
  wire ad429d;
  wire ad429e;
  wire ad429f;
  wire ad42a0;
  wire ad42a1;
  wire ad42a2;
  wire ad42a3;
  wire ad42a4;
  wire ad42a5;
  wire ad42a6;
  wire ad42a7;
  wire ad42a8;
  wire ad42a9;
  wire ad42aa;
  wire ad42ab;
  wire ad42af;
  wire ad42b0;
  wire ad42b1;
  wire ad42b2;
  wire ad42b3;
  wire ad42b4;
  wire ad42b5;
  wire ad42b6;
  wire ad42b7;
  wire ad42b8;
  wire ad42b9;
  wire ad42ba;
  wire ad42bb;
  wire ad42bc;
  wire ad42bd;
  wire ad42be;
  wire ad42bf;
  wire ad42c0;
  wire ad42c1;
  wire ad42c2;
  wire ad42c3;
  wire ad42c4;
  wire ad42c5;
  wire ad42c6;
  wire ad42c7;
  wire ad42c8;
  wire ad42c9;
  wire ad42ca;
  wire ad42cb;
  wire ad42cc;
  wire ad42cd;
  wire ad42ce;
  wire ad42cf;
  wire ad42d0;
  wire ad42d1;
  wire ad42d2;
  wire ad42d3;
  wire ad42d4;
  wire ad42d5;
  wire ad42d6;
  wire ad42d7;
  wire ad42d8;
  wire ad42d9;
  wire ad42da;
  wire ad42db;
  wire ad42dc;
  wire ad42dd;
  wire ad42de;
  wire ad42df;
  wire ad42e0;
  wire ad42e1;
  wire ad42e2;
  wire ad42e3;
  wire ad42e4;
  wire ad42e5;
  wire ad42e6;
  wire ad42e7;
  wire ad42e8;
  wire ad42e9;
  wire ad42ea;
  wire ad42eb;
  wire ad42ec;
  wire ad42ed;
  wire ad42ee;
  wire ad42ef;
  wire ad42f0;
  wire ad42f1;
  wire ad42f2;
  wire ad42f3;
  wire ad42f4;
  wire ad42f5;
  wire ad42f6;
  wire ad42f7;
  wire ad42f8;
  wire ad42f9;
  wire ad42fa;
  wire ad42fb;
  wire ad42fc;
  wire ad42fd;
  wire ad42fe;
  wire ad42ff;
  wire ad4300;
  wire ad4301;
  wire ad4302;
  wire ad4303;
  wire ad4304;
  wire ad4305;
  wire ad4306;
  wire ad4307;
  wire ad4308;
  wire ad4309;
  wire ad430a;
  wire ad430b;
  wire ad430c;
  wire ad430d;
  wire ad430e;
  wire ad430f;
  wire ad4310;
  wire ad4311;
  wire ad4312;
  wire ad4313;
  wire ad4314;
  wire ad4315;
  wire ad4316;
  wire ad4317;
  wire ad4318;
  wire ad4319;
  wire ad431a;
  wire ad431b;
  wire ad431c;
  wire ad431d;
  wire ad431e;
  wire ad431f;
  wire ad4320;
  wire ad4321;
  wire ad4322;
  wire ad4323;
  wire ad4324;
  wire ad4325;
  wire ad4326;
  wire ad4327;
  wire ad4328;
  wire ad4329;
  wire ad432a;
  wire ad432b;
  wire ad432c;
  wire ad432d;
  wire ad432e;
  wire ad432f;
  wire ad4330;
  wire ad4331;
  wire ad4332;
  wire ad4333;
  wire ad4334;
  wire ad4335;
  wire ad4336;
  wire ad4337;
  wire ad4338;
  wire ad4339;
  wire ad433a;
  wire ad433b;
  wire ad433c;
  wire ad433d;
  wire ad433e;
  wire ad433f;
  wire ad4340;
  wire ad4341;
  wire ad4342;
  wire ad4343;
  wire ad4344;
  wire ad4345;
  wire ad4346;
  wire ad4347;
  wire ad4348;
  wire ad4349;
  wire ad434a;
  wire ad434b;
  wire ad434c;
  wire ad434d;
  wire ad434e;
  wire ad434f;
  wire ad4350;
  wire ad4351;
  wire ad4352;
  wire ad4353;
  wire ad4354;
  wire ad4355;
  wire ad4356;
  wire ad4357;
  wire ad4358;
  wire ad4359;
  wire ad435a;
  wire ad435b;
  wire ad435c;
  wire ad435d;
  wire ad435e;
  wire ad435f;
  wire ad4360;
  wire ad4361;
  wire ad4362;
  wire ad4363;
  wire ad4364;
  wire ad4365;
  wire ad4366;
  wire ad4367;
  wire ad4368;
  wire ad4369;
  wire ad436a;
  wire ad436b;
  wire ad436c;
  wire ad436d;
  wire ad436e;
  wire ad436f;
  wire ad4370;
  wire ad4371;
  wire ad4372;
  wire ad4373;
  wire ad4374;
  wire ad4375;
  wire ad4376;
  wire ad4377;
  wire ad4378;
  wire ad4379;
  wire ad437a;
  wire ad437b;
  wire ad437d;
  wire ad437e;
  wire ad437f;
  wire ad4380;
  wire ad4381;
  wire ad4382;
  wire ad4383;
  wire ad4384;
  wire ad4385;
  wire ad4387;
  wire ad4388;
  wire ad4389;
  wire ad438a;
  wire ad438b;
  wire ad438c;
  wire ad438d;
  wire ad438e;
  wire ad438f;
  wire ad4390;
  wire ad4391;
  wire ad4392;
  wire ad4393;
  wire ad4394;
  wire ad4395;
  wire ad4396;
  wire ad4397;
  wire ad4398;
  wire ad4399;
  wire ad439a;
  wire ad439b;
  wire ad439c;
  wire ad439d;
  wire ad439e;
  wire ad439f;
  wire ad43a0;
  wire ad43a1;
  wire ad43a2;
  wire ad43a3;
  wire ad43a4;
  wire ad43a5;
  wire ad43a6;
  wire ad43a7;
  wire ad43a8;
  wire ad43a9;
  wire ad43aa;
  wire ad43ab;
  wire ad43ac;
  wire ad43b5;
  wire ad43b6;
  wire ad43b7;
  wire ad43b8;
  wire ad43b9;
  wire ad43ba;
  wire ad43bb;
  wire ad43bc;
  wire ad43bd;
  wire ad43be;
  wire ad43bf;
  wire ad43c0;
  wire ad43c1;
  wire ad43c2;
  wire ad43c3;
  wire ad43c4;
  wire ad43c6;
  wire ad43c7;
  wire ad43c8;
  wire ad43c9;
  wire ad43ca;
  wire ad43cb;
  wire ad43cc;
  wire ad43cd;
  wire ad43cf;
  wire ad43d0;
  wire ad43d1;
  wire ad43d2;
  wire ad43d3;
  wire ad43d4;
  wire ad43d7;
  wire ad43d8;
  wire ad43d9;
  wire ad43da;
  wire ad43db;
  wire ad43dc;
  wire v845549;
  wire ad43dd;
  wire ad43de;
  wire ad43df;
  wire ad43e0;
  wire ad43ef;
  wire ad43f0;
  wire ad43f1;
  wire ad43f2;
  wire ad43f3;
  wire ad43f4;
  wire ad43f5;
  wire ad43f6;
  wire ad43f7;
  wire ad43f8;
  wire ad43f9;
  wire ad43fa;
  wire ad43fb;
  wire ad43fc;
  wire ad43fd;
  wire ad43fe;
  wire ad43ff;
  wire ad4400;
  wire ad4401;
  wire ad4402;
  wire ad4403;
  wire ad4404;
  wire ad4405;
  wire ad4406;
  wire ad4407;
  wire ad4408;
  wire ad4409;
  wire ad440a;
  wire ad440b;
  wire ad440c;
  wire ad440d;
  wire ad440e;
  wire ad440f;
  wire ad4410;
  wire ad4411;
  wire ad4412;
  wire ad4413;
  wire ad4414;
  wire ad4415;
  wire ad4416;
  wire ad4417;
  wire ad4418;
  wire ad4419;
  wire ad441a;
  wire ad441b;
  wire ad441c;
  wire ad441d;
  wire ad441e;
  wire ad441f;
  wire ad4420;
  wire ad4421;
  wire ad4422;
  wire ad4423;
  wire ad4424;
  wire ad4425;
  wire ad4426;
  wire ad4427;
  wire ad4428;
  wire ad4429;
  wire ad442a;
  wire ad442b;
  wire ad442c;
  wire ad442d;
  wire ad442e;
  wire ad442f;
  wire ad4430;
  wire ad4431;
  wire ad4432;
  wire ad4433;
  wire ad4434;
  wire ad4435;
  wire ad4436;
  wire ad4437;
  wire ad4438;
  wire ad4439;
  wire ad443a;
  wire ad443b;
  wire ad443c;
  wire ad443d;
  wire ad443e;
  wire ad443f;
  wire ad4440;
  wire ad4456;
  wire ad4457;
  wire ad4458;
  wire ad4459;
  wire ad445a;
  wire ad445b;
  wire ad445c;
  wire ad445d;
  wire ad445e;
  wire ad445f;
  wire ad4460;
  wire ad4461;
  wire ad4462;
  wire ad4463;
  wire ad4464;
  wire ad4465;
  wire ad4466;
  wire ad4467;
  wire ad4468;
  wire ad4469;
  wire ad446a;
  wire ad446b;
  wire ad446c;
  wire ad446d;
  wire ad446e;
  wire ad446f;
  wire ad4470;
  wire ad4471;
  wire ad4472;
  wire ad4473;
  wire ad4474;
  wire ad4475;
  wire ad4476;
  wire ad4477;
  wire ad4478;
  wire ad4479;
  wire ad447a;
  wire ad447b;
  wire ad4480;
  wire ad4481;
  wire ad4482;
  wire ad4483;
  wire ad4484;
  wire ad4485;
  wire ad4486;
  wire ad4487;
  wire ad4488;
  wire ad4489;
  wire ad448a;
  wire ad448b;
  wire ad448c;
  wire ad448d;
  wire ad448e;
  wire ad448f;
  wire ad4490;
  wire ad4499;
  wire ad449a;
  wire ad44a3;
  wire ad44a4;
  wire ad44a5;
  wire ad44a6;
  wire ad44a7;
  wire ad44a8;
  wire ad44b1;
  wire ad44b2;
  wire ad44b3;
  wire ad44b4;
  wire ad44b5;
  wire ad44b6;
  wire ad44b7;
  wire ad3cbb;
  wire ad3cbc;
  wire ad3cbd;
  wire ad3cbe;
  wire ad3cbf;
  wire ad3cc0;
  wire ad3cc1;
  wire ad3cc2;
  wire ad3cc3;
  wire ad3cc4;
  wire ad3cc5;
  wire ad3cc8;
  wire ad3cc9;
  wire ad3cca;
  wire ad3ccb;
  wire ad3ccc;
  wire ad3ccd;
  wire ad3cce;
  wire ad3ccf;
  wire ad3cd0;
  wire ad3cd5;
  wire ad3cd6;
  wire ad3cd7;
  wire ad3cd8;
  wire ad3cd9;
  wire ad3cda;
  wire ad3cdb;
  wire ad3cdc;
  wire ad3cdd;
  wire ad3cde;
  wire ad3cdf;
  wire ad3ce0;
  wire ad3ce1;
  wire ad3ce2;
  wire ad3ce3;
  wire ad3ce4;
  wire ad3ce5;
  wire ad3ce6;
  wire ad3ce7;
  wire ad3ce8;
  wire ad3ce9;
  wire ad3cea;
  wire ad3ceb;
  wire ad3cec;
  wire ad3ced;
  wire ad3cee;
  wire ad3cef;
  wire ad3cf0;
  wire ad3cf1;
  wire ad3cf6;
  wire ad3cf7;
  wire ad3cf8;
  wire ad3cf9;
  wire ad3cfa;
  wire ad3cfb;
  wire ad3cfc;
  wire ad3cfd;
  wire ad3cfe;
  wire ad3cff;
  wire ad3d00;
  wire ad3d01;
  wire ad3d02;
  wire ad3d03;
  wire ad3d04;
  wire ad3d05;
  wire ad3d06;
  wire ad3d07;
  wire ad3d08;
  wire ad3d09;
  wire ad3d0a;
  wire ad3d0b;
  wire ad3d0c;
  wire ad3d0d;
  wire ad3d0e;
  wire ad3d0f;
  wire ad3d10;
  wire ad3d11;
  wire ad3d12;
  wire ad3d13;
  wire ad3d14;
  wire ad3d15;
  wire ad3d16;
  wire ad3d17;
  wire ad3d18;
  wire ad3d19;
  wire ad3d1a;
  wire ad3d1b;
  wire ad3d1c;
  wire ad3d1d;
  wire ad3d1e;
  wire ad3d1f;
  wire ad3d20;
  wire ad3d21;
  wire ad3d22;
  wire ad3d23;
  wire ad3d24;
  wire ad3d25;
  wire ad3d26;
  wire ad3d27;
  wire ad3d2b;
  wire ad3d2c;
  wire ad3d2d;
  wire ad3d2e;
  wire ad3d2f;
  wire ad3d30;
  wire ad3d31;
  wire ad3d32;
  wire ad3d33;
  wire ad3d34;
  wire ad3d35;
  wire ad3d36;
  wire ad3d37;
  wire ad3d38;
  wire ad3d39;
  wire ad3d3a;
  wire ad3d3e;
  wire ad3d3f;
  wire ad3d40;
  wire ad3d41;
  wire ad3d42;
  wire ad3d43;
  wire ad3d44;
  wire ad3d45;
  wire ad3d46;
  wire ad3d47;
  wire ad3d48;
  wire ad3d49;
  wire ad3d4a;
  wire ad3d4b;
  wire ad3d4e;
  wire ad3d4f;
  wire ad3d50;
  wire ad3d51;
  wire ad3d52;
  wire ad3d53;
  wire ad3d54;
  wire ad3d55;
  wire ad3d56;
  wire ad3d57;
  wire ad3d58;
  wire ad3d59;
  wire ad3d5a;
  wire ad3d5b;
  wire ad3d5c;
  wire ad3d5d;
  wire ad3d5e;
  wire ad3d5f;
  wire ad3d60;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hbusreq2_p;
  input hbusreq2;
  reg hlock2_p;
  input hlock2;
  reg hbusreq3_p;
  input hbusreq3;
  reg hlock3_p;
  input hlock3;
  reg hbusreq4_p;
  input hbusreq4;
  reg hlock4_p;
  input hlock4;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmaster1_p;
  output hmaster1;
  reg hmaster2_p;
  output hmaster2;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg hgrant2_p;
  output hgrant2;
  reg hgrant3_p;
  output hgrant3;
  reg hgrant4_p;
  output hgrant4;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg stateG10_2_p;
  output stateG10_2;
  reg stateG10_3_p;
  output stateG10_3;
  reg stateG10_4_p;
  output stateG10_4;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;
  reg jx2_p;
  output jx2;

assign ade658 = hready_p & v845542 | !hready_p & ade657;
assign df54f8 = hlock1_p & df54f7 | !hlock1_p & !v845542;
assign ad3ce8 = hbusreq1 & ad3ce5 | !hbusreq1 & ad3ce7;
assign cc36f8 = hgrant1_p & cc36c6 | !hgrant1_p & cc36f6;
assign v9f77d0 = hgrant1_p & v9f772d | !hgrant1_p & v9f77c8;
assign b058e1 = hmaster0_p & b058cd | !hmaster0_p & b058e0;
assign b058d2 = hbusreq4_p & v9ea3e9 | !hbusreq4_p & v9f7d42;
assign ade576 = hbusreq1_p & ade56a | !hbusreq1_p & ade575;
assign bd5b92 = hburst0 & v8ccb69 | !hburst0 & bd5b91;
assign v9f7cab = hbusreq4 & v9f7ca9 | !hbusreq4 & v9f7caa;
assign bd587f = hgrant4_p & bd576b | !hgrant4_p & !adec89;
assign v9f7e03 = hmaster1_p & v9f7e02 | !hmaster1_p & v9f7d2f;
assign dc53cc = decide_p & dc53cb | !decide_p & !v845542;
assign d356c6 = hbusreq3 & d356c5 | !hbusreq3 & !v84554e;
assign v9ea43c = hmaster0_p & v9ea43a | !hmaster0_p & v9ea43b;
assign ad4e8e = hmaster2_p & ad4e8d | !hmaster2_p & v845542;
assign dc5015 = hgrant1_p & dc4ffe | !hgrant1_p & dc5014;
assign v9e9f5d = hbusreq1 & v9e9f5b | !hbusreq1 & v9e9f5c;
assign ade553 = hlock0_p & ade551 | !hlock0_p & ade552;
assign v9ea456 = hbusreq1_p & v9ea3fa | !hbusreq1_p & v9ea455;
assign b1d007 = hgrant2_p & v845542 | !hgrant2_p & b1d006;
assign c3d5b5 = hbusreq4_p & c3d5b3 | !hbusreq4_p & c3d5b4;
assign ad4439 = hmaster2_p & ad442b | !hmaster2_p & ad4438;
assign v9f7e12 = hgrant4_p & v9f7c9c | !hgrant4_p & v9f7d70;
assign ad4e5f = hbusreq3 & ad4e5e | !hbusreq3 & v845542;
assign ad4e64 = hbusreq1 & ad4e42 | !hbusreq1 & v845542;
assign ad457f = hmaster0_p & ad4578 | !hmaster0_p & ad457e;
assign v9f7db4 = hmaster2_p & v9f7d88 | !hmaster2_p & v9f7db3;
assign ade4d5 = hbusreq4_p & ade4d4 | !hbusreq4_p & !v845542;
assign df51b9 = hready_p & df51b1 | !hready_p & df51b8;
assign c74621 = hburst0_p & v845542 | !hburst0_p & c74620;
assign ad4f50 = hmaster1_p & ad4f43 | !hmaster1_p & ad4f4f;
assign ad4e66 = hbusreq1 & ad4e65 | !hbusreq1 & !v845542;
assign b1cff8 = hgrant0_p & d35a4f | !hgrant0_p & v845542;
assign bd58c2 = hmaster2_p & bd58bb | !hmaster2_p & bd58c1;
assign d359c9 = locked_p & d359c8 | !locked_p & adeca0;
assign v9f76d7 = hgrant2_p & v9f76d4 | !hgrant2_p & v9f76d6;
assign bd5791 = hmaster2_p & bd5786 | !hmaster2_p & !bd5790;
assign c3cf2c = hready_p & v845555 | !hready_p & !c3d36c;
assign aa425f = jx0_p & aa425e | !jx0_p & v845542;
assign v9f7cac = hready & v9f7cab | !hready & v9f7ca7;
assign bd5b7b = hbusreq2_p & bd5b7a | !hbusreq2_p & v845542;
assign d356a4 = locked_p & d356a3 | !locked_p & !v845542;
assign ade545 = hmaster0_p & ade543 | !hmaster0_p & ade544;
assign ade4df = hburst0 & c3d66d | !hburst0 & ade4de;
assign d3559b = hbusreq1_p & d35437 | !hbusreq1_p & d3559a;
assign b57446 = decide_p & v845542 | !decide_p & b57445;
assign v8cc0ca = hbusreq4 & v8cc0c5 | !hbusreq4 & v8cc0c9;
assign v9f76cf = hmaster1_p & v9f76ce | !hmaster1_p & v9f7d64;
assign df51af = hmaster1_p & df51ae | !hmaster1_p & df51a9;
assign b57a30 = hmaster1_p & b579b4 | !hmaster1_p & b57a2f;
assign b1c787 = hbusreq2_p & b1c784 | !hbusreq2_p & b1c786;
assign ad43c6 = hbusreq0_p & v9f21c4 | !hbusreq0_p & v845542;
assign ade65a = hgrant1_p & v845542 | !hgrant1_p & !ade659;
assign df54f3 = hbusreq1_p & df54f2 | !hbusreq1_p & !v845542;
assign c3ced2 = hgrant1_p & v84554d | !hgrant1_p & c3ced1;
assign v9f7d97 = hbusreq1 & v9f7d95 | !hbusreq1 & v9f7d96;
assign c3d3ad = hbusreq3_p & c3d387 | !hbusreq3_p & c3d3ac;
assign d35a5e = hgrant4_p & v84556c | !hgrant4_p & d35a5d;
assign d3578c = hmaster2_p & d3578a | !hmaster2_p & d3578b;
assign b1c754 = hburst0 & b1c74f | !hburst0 & b1c753;
assign b0594d = hbusreq1_p & b0594c | !hbusreq1_p & b058fd;
assign c3d684 = hmaster0_p & c3d682 | !hmaster0_p & c3d683;
assign bd586e = hgrant4_p & bd5838 | !hgrant4_p & !bd5842;
assign bd5b86 = hburst1 & adea98 | !hburst1 & bd5b85;
assign ad46cf = hbusreq4_p & ad46ce | !hbusreq4_p & v845542;
assign dc4fb6 = hbusreq1 & dc4f9e | !hbusreq1 & dc4f89;
assign v8cc62b = hlock3 & v8ccbd8 | !hlock3 & v8cc4b4;
assign b1c75a = hlock0_p & bd578b | !hlock0_p & b1c759;
assign ad440b = hbusreq0_p & ad5016 | !hbusreq0_p & v845542;
assign ad458a = hbusreq4 & ad4f1d | !hbusreq4 & !v845542;
assign v8cc0d9 = hbusreq4_p & v8cc48e | !hbusreq4_p & v8cc0d8;
assign c3d696 = hmaster2_p & c3d669 | !hmaster2_p & c3d66e;
assign ad484f = hlock1_p & ad484e | !hlock1_p & ad4da1;
assign ad45cb = hlock1_p & ad45c4 | !hlock1_p & ad45ca;
assign v9ea60a = hbusreq2 & v9ea609 | !hbusreq2 & v9ea607;
assign b059f4 = hbusreq2 & b059f2 | !hbusreq2 & b059f3;
assign v8cc7d7 = hbusreq2_p & v8cc7d5 | !hbusreq2_p & v8cc7d3;
assign ac1483 = decide_p & cc36ba | !decide_p & ac1451;
assign v9f7d5c = hmaster0_p & v9f7d5a | !hmaster0_p & v9f7d5b;
assign v9f773e = hbusreq2_p & v9f773b | !hbusreq2_p & v9f773d;
assign dc5046 = hgrant4_p & ade4aa | !hgrant4_p & ade59c;
assign bd5920 = hready_p & bd591e | !hready_p & !bd591f;
assign d35429 = hbusreq2 & d35421 | !hbusreq2 & d35428;
assign ad4141 = hmaster2_p & ad4140 | !hmaster2_p & ad4f0f;
assign c3ce54 = hbusreq1 & c3d300 | !hbusreq1 & c3d305;
assign ac1480 = decide_p & ac1472 | !decide_p & ac147e;
assign d3551b = hmaster1_p & d3550e | !hmaster1_p & d3551a;
assign ad4827 = hbusreq2_p & ad4826 | !hbusreq2_p & v845542;
assign v9ea615 = hgrant2_p & v9ea612 | !hgrant2_p & v9ea614;
assign bd5831 = hbusreq2 & bd5830 | !hbusreq2 & v845542;
assign v92e9d9 = hmaster1_p & v8a9702 | !hmaster1_p & v845542;
assign ad456a = hbusreq4 & ad4565 | !hbusreq4 & ad4569;
assign bd5756 = hbusreq0_p & adec89 | !hbusreq0_p & bd574e;
assign v9ea628 = hready_p & v9ea4a4 | !hready_p & v9ea627;
assign v9f7d92 = hbusreq0 & v9f7d7f | !hbusreq0 & v9f7d91;
assign c3ce9f = hready & c3ce9e | !hready & !v845564;
assign b1cf26 = hlock0_p & bd5b6e | !hlock0_p & v845542;
assign b1c091 = hgrant3_p & b1c04c | !hgrant3_p & b1c090;
assign v9f784f = hmaster0_p & v9f7829 | !hmaster0_p & v9f784e;
assign bd5853 = hbusreq0 & bd584d | !hbusreq0 & bd5852;
assign v9ea416 = hbusreq1_p & v9ea3e1 | !hbusreq1_p & v9ea415;
assign b0598d = hbusreq0_p & b0598c | !hbusreq0_p & b0597f;
assign b57948 = hmaster1_p & b57947 | !hmaster1_p & v845542;
assign dc52fd = hmastlock_p & v8cc7d9 | !hmastlock_p & v845542;
assign adea9e = hmaster2_p & adea9d | !hmaster2_p & adea94;
assign ade5de = decide_p & ade5dd | !decide_p & v845542;
assign b1c81d = hmaster2_p & v845542 | !hmaster2_p & !d35a9c;
assign v845552 = hlock2_p & v845542 | !hlock2_p & !v845542;
assign ad3d2f = hmaster1_p & ad3d2e | !hmaster1_p & ad4419;
assign bd590d = hlock2_p & bd590c | !hlock2_p & v845542;
assign cc36f5 = hmaster2_p & d35a49 | !hmaster2_p & cc36f4;
assign v8cc80c = hlock3 & v8ccb6b | !hlock3 & v8cc7e6;
assign dc53da = decide_p & dc53d7 | !decide_p & v845542;
assign v9f764d = hgrant1_p & v9f764b | !hgrant1_p & v9f764c;
assign c3d5de = hbusreq0 & c3d5d8 | !hbusreq0 & c3d5dd;
assign ade4e3 = hmaster2_p & adeaae | !hmaster2_p & !ade4e2;
assign v9e9e9c = hgrant4_p & v9ea3e6 | !hgrant4_p & v9e9e9b;
assign v9f7734 = hlock0_p & v845542 | !hlock0_p & v9f7733;
assign c3cf32 = jx1_p & c3cf2b | !jx1_p & c3cf31;
assign ad4db2 = hbusreq4_p & adea85 | !hbusreq4_p & v845542;
assign b1c824 = decide_p & b1c823 | !decide_p & v845542;
assign b05a6a = hlock0 & b05a69 | !hlock0 & b05a61;
assign v9f7d5e = hmaster2_p & v9f7d59 | !hmaster2_p & !v9f7d5d;
assign b05a7b = hbusreq1_p & b0595b | !hbusreq1_p & b05a69;
assign b57a6e = hbusreq1_p & b57942 | !hbusreq1_p & b57a6d;
assign v9e9fd9 = hmaster1_p & v9ea3e7 | !hmaster1_p & v9ea3f0;
assign v9e9fd2 = hgrant2_p & v9ea602 | !hgrant2_p & v9e9fd1;
assign ad45c3 = hmaster0_p & ad45c1 | !hmaster0_p & ad45c2;
assign d359d4 = hmaster2_p & d3599c | !hmaster2_p & d359d3;
assign d35a54 = hgrant1_p & d35a53 | !hgrant1_p & d35a4a;
assign stateG3_0 = !b57538;
assign c3ce00 = hmaster1_p & c3d306 | !hmaster1_p & c3cdff;
assign c5c99d = hgrant3_p & c5c8ee | !hgrant3_p & c5c99c;
assign b57acc = hmaster1_p & b57acb | !hmaster1_p & b57901;
assign v9f7d6d = hlock1_p & v9f7cbe | !hlock1_p & v9f7d0c;
assign cc36db = hgrant4_p & cc36bd | !hgrant4_p & cc36da;
assign ad442a = hgrant4_p & ad4380 | !hgrant4_p & b1cfcb;
assign dc4fa8 = hmaster2_p & dc4fa6 | !hmaster2_p & dc4fa7;
assign b059fa = hlock2 & b058a8 | !hlock2 & b059f9;
assign b1c80d = hbusreq1_p & b1c739 | !hbusreq1_p & b1c807;
assign v9f76da = hgrant2_p & v9f76d9 | !hgrant2_p & v9f76d6;
assign d35a37 = hbusreq2 & df54f5 | !hbusreq2 & df54f6;
assign df50da = hbusreq1_p & df50d9 | !hbusreq1_p & v845542;
assign d359bf = hburst1 & d359bc | !hburst1 & d359be;
assign v9ea451 = hlock4 & v9ea3fa | !hlock4 & v9ea450;
assign d359aa = hbusreq4 & d359a4 | !hbusreq4 & d359a9;
assign b1c76d = hbusreq4_p & b1c756 | !hbusreq4_p & !ade4d4;
assign b57a88 = hbusreq2 & b57a87 | !hbusreq2 & b57942;
assign d35be5 = hbusreq4_p & d35be4 | !hbusreq4_p & v845542;
assign v9ea4d8 = hbusreq4_p & v9ea4d6 | !hbusreq4_p & v9ea4d7;
assign b1c5de = decide_p & b1c5dd | !decide_p & v845542;
assign ade626 = decide_p & ade625 | !decide_p & adeaa7;
assign ade4c1 = stateA1_p & v845542 | !stateA1_p & !ade4ba;
assign ad4dc3 = stateA1_p & ad4dc2 | !stateA1_p & adea85;
assign c3d5a1 = hmaster2_p & c3d59e | !hmaster2_p & v845542;
assign d3556b = hbusreq2 & d35c08 | !hbusreq2 & !v84555a;
assign b57952 = hgrant0_p & b5b408 | !hgrant0_p & v845542;
assign c3ce13 = hbusreq3 & c3d2d6 | !hbusreq3 & c3d2d9;
assign b1c56b = hmaster1_p & b1c85a | !hmaster1_p & b1c56a;
assign v9ea4b0 = hmaster1_p & v9ea4a8 | !hmaster1_p & v9ea4af;
assign ade589 = locked_p & ade588 | !locked_p & c3d66d;
assign d35a6b = hgrant1_p & df54f3 | !hgrant1_p & d35a6a;
assign d356e7 = hmaster0_p & d356da | !hmaster0_p & d356e2;
assign v9ea4ba = hbusreq0_p & v9ea3fb | !hbusreq0_p & v9ea4b6;
assign c5c8a3 = hlock2_p & c5c8a0 | !hlock2_p & c5c8a2;
assign b1c097 = hready_p & b1c096 | !hready_p & b1c707;
assign ad4280 = hbusreq2_p & ad427b | !hbusreq2_p & ad427f;
assign c3d34d = hbusreq0 & c3d342 | !hbusreq0 & c3d34c;
assign b05a32 = hmaster0_p & b059fb | !hmaster0_p & b058c5;
assign b57425 = hbusreq1 & b57423 | !hbusreq1 & b57424;
assign ad4fb3 = hready & v84556c | !hready & dc4fcb;
assign c3d6c2 = hgrant4_p & c3d681 | !hgrant4_p & !c3d6ac;
assign stateG2 = !c5bed6;
assign v9f7811 = hmaster0_p & v9f7808 | !hmaster0_p & !v9f7810;
assign v9f765c = hmaster2_p & v9f7655 | !hmaster2_p & v9f765b;
assign c3ceb1 = hbusreq3 & c3ceae | !hbusreq3 & c3ceb0;
assign b05926 = hmaster0_p & b05921 | !hmaster0_p & b05925;
assign b57ac6 = hbusreq1_p & b578f9 | !hbusreq1_p & b57ac5;
assign b1c731 = hlock0_p & c3d669 | !hlock0_p & !v845542;
assign bd574e = locked_p & v845542 | !locked_p & !c3d674;
assign ad428d = hmaster1_p & ad428c | !hmaster1_p & ad4289;
assign v9f7853 = decide_p & v9f7784 | !decide_p & v9f7852;
assign ad4384 = hbusreq0 & ad4383 | !hbusreq0 & v845542;
assign b1d000 = hgrant4_p & v845542 | !hgrant4_p & b1cfff;
assign b57905 = hlock2_p & b57902 | !hlock2_p & b57904;
assign bd57d2 = hbusreq2 & bd57d1 | !hbusreq2 & !v845542;
assign dc538e = hbusreq3 & dc5389 | !hbusreq3 & dc538d;
assign bd5728 = hgrant3_p & bd56e0 | !hgrant3_p & !bd56cc;
assign hgrant3 = dc53e0;
assign ad4270 = hbusreq3 & ad4269 | !hbusreq3 & ad426f;
assign b1c84d = hbusreq2_p & b1c82f | !hbusreq2_p & b1c84b;
assign b1cf37 = hgrant2_p & b1cf35 | !hgrant2_p & b1cf2f;
assign c3cf05 = hmaster2_p & c3cf00 | !hmaster2_p & v845542;
assign v9ea5d1 = hlock1 & v9ea5cb | !hlock1 & v9ea5d0;
assign adec90 = locked_p & adec8f | !locked_p & c3d66d;
assign bbbcd8 = start_p & v845542 | !start_p & !bbbcd6;
assign c3d4f3 = hbusreq4 & c3d4e3 | !hbusreq4 & !c3d4f2;
assign d35bfe = hmaster1_p & d35bfd | !hmaster1_p & d35bfa;
assign dc5065 = hgrant1_p & dc5035 | !hgrant1_p & dc5064;
assign v9f774a = hlock1 & v9f7745 | !hlock1 & v9f7749;
assign b573dd = hbusreq2 & b573db | !hbusreq2 & b573dc;
assign b1caf6 = hbusreq4_p & d3591a | !hbusreq4_p & !v84554a;
assign b1c03f = hbusreq1_p & b1c766 | !hbusreq1_p & b1c03e;
assign d359c6 = hbusreq1 & d359ad | !hbusreq1 & !d359c5;
assign bd589a = hgrant2_p & bd5bab | !hgrant2_p & !bd5899;
assign v9f7690 = hmaster2_p & v9f768f | !hmaster2_p & !v9ea448;
assign v9f7ca6 = locked_p & v9f7c9d | !locked_p & v9ea3ec;
assign v9ea4b6 = locked_p & v845542 | !locked_p & v9ea4a6;
assign v8cc7c4 = hbusreq4 & v8cc7c2 | !hbusreq4 & v8cc7c3;
assign df54e5 = hbusreq1_p & df54e4 | !hbusreq1_p & v845542;
assign b1c50d = decide_p & b1c50c | !decide_p & v845542;
assign b1cfbf = hbusreq4_p & b1cfb7 | !hbusreq4_p & !b1cfbe;
assign dc4f9e = hmaster2_p & ade4bf | !hmaster2_p & dc4f9d;
assign ade588 = hburst0 & c3d66b | !hburst0 & ade587;
assign b1c4cd = hbusreq4 & b1c4c7 | !hbusreq4 & b1c4cc;
assign ad4dbc = hbusreq3 & ad4da1 | !hbusreq3 & v845542;
assign v9ea4aa = stateG10_4_p & v9ea3e9 | !stateG10_4_p & !v9ea4a6;
assign c3d5c8 = hmaster2_p & c3d5bf | !hmaster2_p & v845542;
assign c3d4f7 = hready & c3d4f3 | !hready & c3d4f6;
assign dc506d = hbusreq3 & dc501a | !hbusreq3 & !v845542;
assign d356cc = hbusreq3 & d356cb | !hbusreq3 & !v84554e;
assign df5125 = hlock1_p & df5124 | !hlock1_p & !v845542;
assign b05a27 = hmaster1_p & b05a26 | !hmaster1_p & b05a20;
assign c3ceaf = hready & d35a99 | !hready & v845564;
assign bd5883 = hbusreq4_p & bd5880 | !hbusreq4_p & bd5882;
assign d357a8 = hmaster0_p & d35791 | !hmaster0_p & d35799;
assign bd5868 = stateG10_4_p & bd5865 | !stateG10_4_p & bd5867;
assign c3d52f = hbusreq1 & c3d526 | !hbusreq1 & c3d52a;
assign ad4f15 = hbusreq3 & ad4f14 | !hbusreq3 & v845542;
assign adeaa8 = decide_p & adeaa2 | !decide_p & adeaa7;
assign ad4289 = hmaster0_p & ad4286 | !hmaster0_p & !ad4288;
assign c5c8fd = hlock0_p & c5c8fc | !hlock0_p & !v845542;
assign b8f6e7 = hgrant3_p & b8f6e0 | !hgrant3_p & b8f6e6;
assign b059f8 = hlock3 & b058a8 | !hlock3 & b059ca;
assign b1c5e3 = hgrant2_p & v845542 | !hgrant2_p & b1c5e2;
assign ad3cdf = hmaster2_p & b1c714 | !hmaster2_p & !ad3cde;
assign ad48c9 = hready_p & v845542 | !hready_p & ad48c8;
assign ad3d3f = hgrant2_p & ad446d | !hgrant2_p & ad3d3e;
assign v9e9fa9 = hgrant1_p & v9e9eed | !hgrant1_p & v9e9f7f;
assign c3d4e2 = hmaster2_p & c3d4df | !hmaster2_p & c3d4e1;
assign ad4108 = hbusreq1_p & ad4107 | !hbusreq1_p & ad40fe;
assign v8cc475 = hgrant1_p & v845542 | !hgrant1_p & v8cc474;
assign v9f787c = hmaster1_p & v9f787b | !hmaster1_p & v9f7736;
assign ad4e4d = hmaster2_p & v845542 | !hmaster2_p & ad4e4c;
assign v9f7897 = hlock2 & v9f77e2 | !hlock2 & v9f7896;
assign ad44a5 = stateG10_4_p & c3cec2 | !stateG10_4_p & !ad44a4;
assign bd592f = hlock0_p & adea9a | !hlock0_p & bd592e;
assign c3ce05 = hmaster0_p & c3ce03 | !hmaster0_p & c3ce04;
assign dc4f7a = hmastlock_p & dc4f79 | !hmastlock_p & !v845542;
assign v9ea4cc = hmaster0_p & v9ea4cb | !hmaster0_p & v9ea44a;
assign d3558b = hbusreq4_p & d354cb | !hbusreq4_p & !d35aab;
assign busreq = c3cf34;
assign bd5840 = hgrant0_p & v84556c | !hgrant0_p & bd574e;
assign c5c93a = hmaster2_p & c5c935 | !hmaster2_p & !c5c939;
assign ad448e = hbusreq0 & ad448d | !hbusreq0 & v845542;
assign cc36e7 = hmaster2_p & cc36e3 | !hmaster2_p & !cc36e6;
assign v8cc7b5 = hbusreq3 & v8cc7b2 | !hbusreq3 & v8cc7b4;
assign b0595c = hlock0 & b0595b | !hlock0 & b0595a;
assign d3550c = hbusreq4 & d3550a | !hbusreq4 & d3550b;
assign ad474c = hready & ad4748 | !hready & ad474b;
assign b1c868 = decide_p & b1c84d | !decide_p & b1d013;
assign v9f7d8d = hlock4_p & v9f7d8b | !hlock4_p & v9f7d8c;
assign b1d00f = hmaster2_p & v8da5a1 | !hmaster2_p & v8da59f;
assign d359ba = hburst0_p & v845542 | !hburst0_p & !v845568;
assign ade4e7 = hbusreq0_p & ade4e6 | !hbusreq0_p & ade4d9;
assign adeaa2 = hgrant2_p & v845542 | !hgrant2_p & adeaa1;
assign b1c032 = hbusreq4_p & ade4d4 | !hbusreq4_p & b1c031;
assign c3d675 = locked_p & v845542 | !locked_p & c3d674;
assign v9ea4c2 = decide_p & v9ea4b2 | !decide_p & v9ea4c1;
assign ad429c = decide_p & ad428f | !decide_p & ad429b;
assign b1c0aa = hgrant2_p & b1d01a | !hgrant2_p & b1c0a9;
assign b1c58a = hbusreq1_p & b1cf28 | !hbusreq1_p & b1cf32;
assign ad4ef0 = hmaster2_p & ad4eee | !hmaster2_p & ad4eef;
assign bd58f8 = hbusreq1_p & bd58f6 | !hbusreq1_p & bd58f7;
assign df51de = jx1_p & df51dd | !jx1_p & df51d2;
assign ad427f = hmaster1_p & ad427e | !hmaster1_p & ad427a;
assign bd57f7 = stateG2_p & v845542 | !stateG2_p & v889629;
assign b1c725 = hbusreq4_p & b1c71a | !hbusreq4_p & b1c720;
assign ad471d = hgrant2_p & ad46fc | !hgrant2_p & ad471c;
assign v9ea4db = hmaster0_p & v9ea4cf | !hmaster0_p & v9ea4da;
assign bd56cb = decide_p & bd5e25 | !decide_p & !v845572;
assign v9f770d = hbusreq2_p & v9f76db | !hbusreq2_p & v9f770c;
assign d357c9 = hlock4_p & d3576e | !hlock4_p & d357c8;
assign v9f7da1 = stateA1_p & v845542 | !stateA1_p & !v9f7cf2;
assign ad4f34 = hburst0_p & v84557e | !hburst0_p & v8b08c2;
assign v9f7da2 = locked_p & v9f7da1 | !locked_p & v9f7cc6;
assign b57506 = decide_p & b57a21 | !decide_p & b574fa;
assign c3d6f1 = hgrant4_p & c3d66e | !hgrant4_p & !c3d6ab;
assign ad46f5 = hbusreq1_p & ad46f3 | !hbusreq1_p & !ad46f4;
assign c3d305 = hbusreq4 & c3d303 | !hbusreq4 & !c3d304;
assign ad425b = hbusreq2_p & ad425a | !hbusreq2_p & v845542;
assign c3ce33 = jx0_p & c3d3ad | !jx0_p & c3ce32;
assign bd5765 = hmaster1_p & bd5762 | !hmaster1_p & bd5ba9;
assign v9ea59e = hlock0 & v9ea59b | !hlock0 & v9ea59d;
assign c5c8a7 = hmaster1_p & c5c898 | !hmaster1_p & c5c89f;
assign dc53a0 = hbusreq3 & dc5394 | !hbusreq3 & dc539f;
assign b1caed = hmaster2_p & v845542 | !hmaster2_p & b1caec;
assign v9f7e15 = hgrant4_p & v9f7cb4 | !hgrant4_p & v9f7d78;
assign ad3cee = hbusreq4_p & ad3cec | !hbusreq4_p & ad3ced;
assign b05a59 = stateA1_p & v845542 | !stateA1_p & !b05a58;
assign b1c081 = hbusreq0 & b1c080 | !hbusreq0 & b1c85e;
assign d35734 = hbusreq2_p & d35728 | !hbusreq2_p & d35733;
assign d357c2 = hgrant4_p & d3576e | !hgrant4_p & d357c1;
assign d35a0b = hgrant4_p & d359c4 | !hgrant4_p & !v845542;
assign ad4585 = hbusreq4 & d359ad | !hbusreq4 & !v845542;
assign v8cc5fd = hmaster0_p & v8cc5fb | !hmaster0_p & v845542;
assign cc36d6 = hbusreq2_p & cc36d5 | !hbusreq2_p & !cc36d4;
assign d3573e = hmaster0_p & d3573d | !hmaster0_p & d356f8;
assign dc4fc1 = hmaster1_p & dc4fb5 | !hmaster1_p & dc4fc0;
assign df50cb = hbusreq1 & dc52fc | !hbusreq1 & dc5302;
assign ad446e = hgrant2_p & ad446d | !hgrant2_p & ad446a;
assign bd5895 = hbusreq4 & bd587b | !hbusreq4 & bd5894;
assign ad4e7e = hgrant4_p & v845542 | !hgrant4_p & ad4e75;
assign v9f7824 = hbusreq1 & v9f7822 | !hbusreq1 & v9f7823;
assign b1c05d = hmaster0_p & b1c05b | !hmaster0_p & b1c05c;
assign v9f7dc4 = hlock2 & v9f7dc1 | !hlock2 & v9f7dc3;
assign v9ea4a5 = stateA1_p & v9ea3e5 | !stateA1_p & v9ea3e4;
assign b1c728 = hmaster2_p & b1c714 | !hmaster2_p & v845542;
assign b1c5f8 = hgrant3_p & b1c5df | !hgrant3_p & b1c5f7;
assign v9ea442 = hgrant4_p & v9ea3e6 | !hgrant4_p & v9ea441;
assign d3598b = hmaster2_p & d35988 | !hmaster2_p & d3598a;
assign v8cc805 = hlock3 & v8cc43a | !hlock3 & v8cc803;
assign v9f7d7e = hbusreq4_p & v9f7d7c | !hbusreq4_p & v9f7d7d;
assign c3ce3c = hbusreq1 & c3d2c7 | !hbusreq1 & !v845542;
assign ad4e76 = hgrant4_p & d3597f | !hgrant4_p & ad4e75;
assign d35a2e = hbusreq1 & d35a21 | !hbusreq1 & !v845542;
assign d358fb = hbusreq1 & v845542 | !hbusreq1 & d358fa;
assign v9f7cf5 = locked_p & v9f7cf4 | !locked_p & v9f7c9f;
assign ac1475 = stateG10_4_p & v845542 | !stateG10_4_p & !ac1461;
assign v9e9f4a = hmaster1_p & v9e9f49 | !hmaster1_p & v9e9ef1;
assign v9e9f7f = hbusreq1 & v9e9f7d | !hbusreq1 & v9e9f7e;
assign b579cf = hgrant0_p & b579ba | !hgrant0_p & v845542;
assign v8cc4aa = hlock1 & v8cc494 | !hlock1 & v8cc4a9;
assign ad4279 = hbusreq3 & ad4278 | !hbusreq3 & v845542;
assign bd5878 = stateG10_4_p & bd5875 | !stateG10_4_p & bd5877;
assign ad4367 = hmaster0_p & ad4362 | !hmaster0_p & ad4305;
assign ad4f7f = hbusreq4_p & ad4f7e | !hbusreq4_p & b1cfbe;
assign dc4f61 = hbusreq3 & v84556c | !hbusreq3 & v845542;
assign ad4476 = hbusreq2_p & ad446f | !hbusreq2_p & ad4475;
assign ad4f89 = hgrant4_p & v84556c | !hgrant4_p & ad4f88;
assign b1c6e0 = hready_p & b1c82d | !hready_p & b1c6df;
assign b1c7a4 = hgrant4_p & b1c714 | !hgrant4_p & !b1c797;
assign v9f7cb4 = locked_p & v9f7cb3 | !locked_p & !v9f7c9f;
assign c3d75a = hgrant2_p & c3d757 | !hgrant2_p & c3d759;
assign bd58ca = hbusreq4_p & bd58c7 | !hbusreq4_p & bd58c9;
assign bd58bc = hgrant0_p & bd575d | !hgrant0_p & v84556c;
assign ad4407 = hmaster1_p & ad4406 | !hmaster1_p & ad43fc;
assign ad4812 = hbusreq2 & ad4811 | !hbusreq2 & v845542;
assign b5742f = hbusreq3 & b57410 | !hbusreq3 & b5742e;
assign df5144 = hmaster0_p & df513f | !hmaster0_p & df5143;
assign bd57b1 = hmaster0_p & bd57a2 | !hmaster0_p & bd57b0;
assign v8cc0e9 = hmaster1_p & v8cc475 | !hmaster1_p & v8cc0e8;
assign d35a10 = hbusreq4_p & d35a0e | !hbusreq4_p & d35a0f;
assign ad4415 = hbusreq4_p & b1c70e | !hbusreq4_p & b1c714;
assign bd5939 = hgrant2_p & bd5938 | !hgrant2_p & !v845542;
assign b05a3f = hbusreq4_p & b0591c | !hbusreq4_p & b05a3e;
assign df51d4 = decide_p & df511a | !decide_p & v845542;
assign v9ea575 = hmaster2_p & v9ea570 | !hmaster2_p & v9ea574;
assign c5c88b = stateG2_p & v845542 | !stateG2_p & !bb9bdd;
assign b058b3 = hbusreq3 & b058b1 | !hbusreq3 & b058b2;
assign b05905 = hbusreq3 & b05903 | !hbusreq3 & b05904;
assign ad4458 = hbusreq4_p & ad4457 | !hbusreq4_p & v845542;
assign b05995 = hlock4 & b05992 | !hlock4 & b05994;
assign b1c845 = hmaster2_p & d35a9c | !hmaster2_p & !b1c844;
assign v9f76c5 = hbusreq4_p & v9f7d3a | !hbusreq4_p & v9f76c4;
assign d356ba = hlock1_p & d35a2d | !hlock1_p & v84556c;
assign v8cc47a = locked_p & v8cc479 | !locked_p & v845542;
assign c3d5bd = hgrant4_p & v845542 | !hgrant4_p & !c3d5b2;
assign b1d014 = decide_p & b1d00d | !decide_p & b1d013;
assign b1c57e = hbusreq4_p & d3591a | !hbusreq4_p & !v845542;
assign df5164 = hmaster1_p & df515c | !hmaster1_p & df5163;
assign c5c89e = hmaster2_p & c5c89c | !hmaster2_p & c5c89d;
assign v9ea40e = hgrant4_p & v845542 | !hgrant4_p & v9f21c6;
assign dc5085 = decide_p & dc4fc6 | !decide_p & v845542;
assign dc4fe9 = hgrant4_p & c3d66d | !hgrant4_p & ade557;
assign ad473a = hbusreq4_p & ad5032 | !hbusreq4_p & !v845542;
assign ad46a2 = hbusreq4_p & ad46a1 | !hbusreq4_p & v845542;
assign c3d71a = hready_p & c3d706 | !hready_p & !c3d719;
assign b1cfd5 = hgrant2_p & v845542 | !hgrant2_p & b1cfd4;
assign b57412 = hgrant1_p & b57411 | !hgrant1_p & b5794a;
assign v9f7e38 = hlock1 & v9f7e32 | !hlock1 & v9f7e37;
assign df5198 = hmaster1_p & df5190 | !hmaster1_p & df5197;
assign c3d5d1 = hmaster1_p & c3d5ce | !hmaster1_p & c3d5d0;
assign v9f77ab = hbusreq2 & v9f77a9 | !hbusreq2 & v9f77aa;
assign v8cc59b = hbusreq1 & v8cc599 | !hbusreq1 & v8ccbd8;
assign ad470f = hbusreq1_p & ad4705 | !hbusreq1_p & ad4702;
assign v9f7731 = hbusreq1_p & v9f772d | !hbusreq1_p & v9f7730;
assign ad43ab = hready & ad43aa | !hready & ad43a8;
assign c3cebb = hbusreq0_p & v845542 | !hbusreq0_p & v84556e;
assign adea90 = hready_p & v845542 | !hready_p & adea8f;
assign b1c74c = decide_p & b1c74b | !decide_p & v845542;
assign ad3d25 = hmaster1_p & ad3d24 | !hmaster1_p & ad43ba;
assign v9e9f52 = hbusreq4_p & v9e9f50 | !hbusreq4_p & v9e9f51;
assign ad4e5a = hbusreq4_p & v845542 | !hbusreq4_p & ad4e54;
assign ad48b2 = hbusreq3 & ad48a6 | !hbusreq3 & ad48b1;
assign v9f764c = hbusreq1_p & v9f7e1f | !hbusreq1_p & v9f7e3f;
assign dc4fd9 = hmaster2_p & dc4fd8 | !hmaster2_p & ade4aa;
assign b8ef52 = jx0_p & b8ef51 | !jx0_p & b8f745;
assign ad4f69 = hgrant4_p & v845542 | !hgrant4_p & !ad4f67;
assign v9f779c = hmaster0_p & v9f7790 | !hmaster0_p & v9f779b;
assign df512f = hgrant3_p & df511d | !hgrant3_p & df512e;
assign ad4e6b = hmastlock_p & ad4e6a | !hmastlock_p & !v845542;
assign v9ea473 = hbusreq4_p & v9ea471 | !hbusreq4_p & v9ea472;
assign c5c92c = hbusreq2_p & c5c905 | !hbusreq2_p & c5c904;
assign b05942 = hmaster2_p & b0593f | !hmaster2_p & b05941;
assign b05a4b = decide_p & b05a45 | !decide_p & !b05a4a;
assign bd57ed = hbusreq2_p & bd57ec | !hbusreq2_p & v845542;
assign v9f7e37 = hready & v9f7e36 | !hready & v9f7e32;
assign c3d6eb = hgrant4_p & c3d675 | !hgrant4_p & c3d6b7;
assign d359b7 = locked_p & d359b6 | !locked_p & v845542;
assign ad45fd = hlock2_p & ad45f9 | !hlock2_p & ad45fc;
assign ad4e86 = hbusreq4_p & ad4e85 | !hbusreq4_p & b1cfcd;
assign v8cc7cb = hlock3 & v8ccbf6 | !hlock3 & v8cc7ca;
assign ade4ad = hmaster2_p & v845542 | !hmaster2_p & adec93;
assign ad42fd = hbusreq2 & ad4281 | !hbusreq2 & !ad4282;
assign v8b08c1 = start_p & v845542 | !start_p & v84557e;
assign v8cc500 = hgrant1_p & v845542 | !hgrant1_p & v8cc4fe;
assign ad13df = hgrant1_p & v845542 | !hgrant1_p & v84554c;
assign c3ce40 = hmaster1_p & c3ce3a | !hmaster1_p & c3ce3f;
assign d359cd = hgrant0_p & adeca0 | !hgrant0_p & d35983;
assign ad4390 = hbusreq3 & ad438f | !hbusreq3 & v845542;
assign bd5919 = hmaster0_p & v84556c | !hmaster0_p & bd5918;
assign ade562 = hgrant0_p & v845542 | !hgrant0_p & !v84556c;
assign b1c584 = hmaster1_p & b1c842 | !hmaster1_p & b1c583;
assign v9f7661 = hgrant0_p & v9f7e31 | !hgrant0_p & !v9f7cc6;
assign v8cc793 = hmastlock_p & v8cc792 | !hmastlock_p & v845542;
assign d354c1 = hbusreq4_p & d354c0 | !hbusreq4_p & v845542;
assign c3cec4 = stateG10_4_p & c3cec2 | !stateG10_4_p & !c3cec3;
assign d35913 = hmaster0_p & d3590b | !hmaster0_p & d35912;
assign c3d6dc = hgrant1_p & c3d6db | !hgrant1_p & c3d6bd;
assign v9e9fb1 = hgrant2_p & v9e9fa8 | !hgrant2_p & v9e9fb0;
assign v8cc0c2 = hbusreq0_p & v8cc47a | !hbusreq0_p & v8d2b2b;
assign ad430b = hbusreq1_p & ad430a | !hbusreq1_p & v845542;
assign d35722 = hbusreq2_p & d35716 | !hbusreq2_p & !d35721;
assign b1cff7 = hmaster2_p & b1cfbf | !hmaster2_p & b1cff6;
assign v9ea5cc = hmaster2_p & v9ea570 | !hmaster2_p & v9ea587;
assign ad4360 = hmaster1_p & ad435f | !hmaster1_p & ad42f9;
assign ac148e = hmaster0_p & ac148d | !hmaster0_p & ac146b;
assign ade5a0 = hbusreq4_p & ade59f | !hbusreq4_p & !v845542;
assign b574b6 = hbusreq4 & b574b4 | !hbusreq4 & b574b5;
assign b8f747 = jx0_p & b8f6e7 | !jx0_p & b8f746;
assign v8cc434 = hbusreq2_p & v8ccbfb | !hbusreq2_p & v8ccbfa;
assign ad42ba = hbusreq1 & ad42b9 | !hbusreq1 & v845542;
assign d35659 = hgrant1_p & df54f3 | !hgrant1_p & d35658;
assign adea8c = hmaster0_p & v845542 | !hmaster0_p & !adea8b;
assign v8cc50a = hgrant2_p & v8cc472 | !hgrant2_p & v8cc509;
assign v9f77e6 = hbusreq2 & v9f77e4 | !hbusreq2 & v9f77e5;
assign ac148f = hmaster1_p & ac148c | !hmaster1_p & ac148e;
assign b1c4a4 = hbusreq4_p & b1c4a3 | !hbusreq4_p & !v84554a;
assign v9f7ce5 = hlock3 & v9f7cdd | !hlock3 & v9f7ce4;
assign d35712 = hbusreq2 & d356c7 | !hbusreq2 & v84554e;
assign d35742 = hgrant2_p & d3573f | !hgrant2_p & d35741;
assign v9f766c = hready & v9f766b | !hready & v9f7667;
assign v9e9e7b = hmaster1_p & v9e9e7a | !hmaster1_p & v9e9e77;
assign c5c93f = hmaster0_p & v845542 | !hmaster0_p & c5c930;
assign ad4894 = hbusreq1_p & ad4db7 | !hbusreq1_p & ad4dd4;
assign ad508e = hmaster1_p & c3d2d9 | !hmaster1_p & ad508d;
assign b1c55e = hmaster2_p & b1c858 | !hmaster2_p & b1c55d;
assign v9ea58d = hlock1 & v9ea586 | !hlock1 & v9ea58c;
assign d359e4 = hbusreq3 & d359e3 | !hbusreq3 & v845542;
assign ad4da0 = hbusreq1 & ad4d98 | !hbusreq1 & ad4d9c;
assign ad5026 = hready & ad4fbd | !hready & !v845542;
assign b579e6 = hbusreq3 & b579e4 | !hbusreq3 & b579e5;
assign ad4ecb = hbusreq4_p & v845542 | !hbusreq4_p & ad4e53;
assign ad3ccb = stateG10_4_p & c3cec2 | !stateG10_4_p & ad3cca;
assign c3cefd = hgrant2_p & v845551 | !hgrant2_p & c3d306;
assign ad4335 = hbusreq3 & ad4331 | !hbusreq3 & ad4334;
assign ad504b = hlock0_p & ad5049 | !hlock0_p & ad504a;
assign v8cc0c9 = hlock4 & v8ccbd8 | !hlock4 & v8cc0c5;
assign b05a98 = decide_p & b05a45 | !decide_p & !b05a97;
assign v9e9ef6 = decide_p & v9e9e75 | !decide_p & v9e9ef5;
assign bd5870 = hbusreq4_p & bd586d | !hbusreq4_p & bd586f;
assign v9f778a = hbusreq4 & v9f7788 | !hbusreq4 & v9f7789;
assign bd5bac = hgrant2_p & bd5bab | !hgrant2_p & !v845542;
assign v9e9f9a = hgrant1_p & v9e9ef0 | !hgrant1_p & v9e9f8e;
assign b059ce = hbusreq1_p & b058aa | !hbusreq1_p & b058a8;
assign b059ae = hgrant4_p & b058b6 | !hgrant4_p & b05953;
assign v9f7876 = hmaster0_p & v9f7730 | !hmaster0_p & v9f772c;
assign df511d = hready_p & v845542 | !hready_p & df511c;
assign ad4820 = hlock3_p & ad481b | !hlock3_p & ad481f;
assign bd58f7 = hbusreq1 & c3d685 | !hbusreq1 & !v845542;
assign b1c565 = hmaster2_p & b1c85e | !hmaster2_p & b1c564;
assign dc53c0 = hbusreq1_p & dc539f | !hbusreq1_p & v845564;
assign c3d6aa = hbusreq4_p & c3d6a7 | !hbusreq4_p & c3d6a9;
assign b1c769 = hmaster2_p & b1c755 | !hmaster2_p & ade4d9;
assign d35a1c = hmaster1_p & d359b3 | !hmaster1_p & d35a1b;
assign dc4fed = hbusreq0 & dc4fe7 | !hbusreq0 & dc4fec;
assign ad4898 = hmaster1_p & ad484d | !hmaster1_p & ad4897;
assign dc4f8a = hbusreq1 & dc4f68 | !hbusreq1 & dc4f89;
assign c3d66b = stateA1_p & v845542 | !stateA1_p & !v889629;
assign d35643 = hbusreq4_p & d35642 | !hbusreq4_p & !d35641;
assign c3d33c = hgrant4_p & v845542 | !hgrant4_p & !c3d33b;
assign d35492 = hbusreq2 & d35bed | !hbusreq2 & d35be8;
assign ade5b4 = hgrant1_p & ade5b3 | !hgrant1_p & !ade57c;
assign ba05ce = decide_p & ba05cd | !decide_p & v845550;
assign bd5851 = hbusreq4_p & bd584e | !hbusreq4_p & bd5850;
assign c3d51b = hbusreq1 & c3d512 | !hbusreq1 & c3d516;
assign ad4698 = hlock4_p & ad4e89 | !hlock4_p & b1cfcb;
assign dc504e = hburst1 & adea98 | !hburst1 & dc504d;
assign b0596e = hlock1_p & b058aa | !hlock1_p & b058ea;
assign ad4734 = hbusreq3 & ad4730 | !hbusreq3 & ad4733;
assign ad4f49 = hbusreq0_p & v845542 | !hbusreq0_p & v84556c;
assign v9f7d26 = hlock4 & v9f7d23 | !hlock4 & !v9f7d25;
assign b57aee = hgrant3_p & b57ae1 | !hgrant3_p & b57aed;
assign v8cc125 = hbusreq3 & v8cc0ee | !hbusreq3 & v8ccbd8;
assign bd589c = stateA1_p & bd589b | !stateA1_p & ade54b;
assign d35aa1 = hbusreq2_p & d35a97 | !hbusreq2_p & d35aa0;
assign v8da5a0 = stateG10_4_p & v84556e | !stateG10_4_p & !v8da59f;
assign ad45f3 = hbusreq4 & ad45ea | !hbusreq4 & ad45f2;
assign b1c72e = hmaster0_p & b1c719 | !hmaster0_p & b1c72d;
assign bd5929 = hmaster1_p & bd5928 | !hmaster1_p & v845542;
assign bd5ea7 = hlock2_p & bd5ea6 | !hlock2_p & !v845542;
assign c3d690 = hlock3_p & c3d680 | !hlock3_p & !c3d68f;
assign v8cc4a4 = hlock0 & v8cc494 | !hlock0 & v8cc4a1;
assign ad433c = hgrant1_p & ad4339 | !hgrant1_p & ad433b;
assign v9f7d81 = hgrant0_p & v9f7ca5 | !hgrant0_p & !v9f7d80;
assign c3ce73 = hready_p & c3ce5c | !hready_p & c3ce72;
assign bd5911 = hbusreq1 & bd5b82 | !hbusreq1 & v84556c;
assign d354da = hbusreq2 & d35c0b | !hbusreq2 & v84555a;
assign d3561b = stateG2_p & v845542 | !stateG2_p & d3561a;
assign d35a9c = hbusreq4_p & v845542 | !hbusreq4_p & v84554a;
assign d35650 = hmaster2_p & d35a5b | !hmaster2_p & d3564f;
assign df54dd = hmastlock_p & df54dc | !hmastlock_p & v845542;
assign d35499 = hbusreq2 & d35495 | !hbusreq2 & d35498;
assign ad4716 = hbusreq4_p & ad4715 | !hbusreq4_p & v845542;
assign c3d39a = hgrant4_p & v845542 | !hgrant4_p & c3d399;
assign d35804 = hready_p & d357f1 | !hready_p & d35803;
assign b57a8a = hmaster1_p & b57a89 | !hmaster1_p & v845542;
assign v8cc0e2 = hlock3 & v8cc4ad | !hlock3 & v8cc0e1;
assign v8cc7ba = hlock4_p & v8cc7b9 | !hlock4_p & v845542;
assign bd5b8f = hlock2_p & bd5b8e | !hlock2_p & !v845542;
assign bd5838 = locked_p & bd5837 | !locked_p & c3d674;
assign d357e8 = hgrant3_p & d357b3 | !hgrant3_p & d357e7;
assign ad46c9 = hmaster2_p & v845542 | !hmaster2_p & ad46c8;
assign v9f77fb = hlock3 & v9f77fa | !hlock3 & v9f77f9;
assign b1c071 = hbusreq4_p & b1c7c3 | !hbusreq4_p & !b1c070;
assign v9f7dba = hlock1 & v9f7db4 | !hlock1 & v9f7db9;
assign ad4f0f = hbusreq4_p & ad4f0e | !hbusreq4_p & ad4f00;
assign c3d2ec = stateG10_4_p & c3d2ea | !stateG10_4_p & c3d2eb;
assign df5136 = jx0_p & df5544 | !jx0_p & df5135;
assign cc36ec = decide_p & v845566 | !decide_p & cc36eb;
assign v9f77b0 = hmaster0_p & v9f77ab | !hmaster0_p & !v9f77af;
assign ad3d00 = hgrant4_p & ad3cde | !hgrant4_p & !ad3ceb;
assign ad46c1 = hready & ad46bb | !hready & ad46c0;
assign v9f775e = hbusreq4 & v9f775c | !hbusreq4 & v9f775d;
assign ad4f3f = hmaster2_p & v845542 | !hmaster2_p & ad4f3e;
assign v8ccbf4 = hmaster2_p & v8ccbee | !hmaster2_p & v8ccbf3;
assign v9f772a = stateA1_p & v845542 | !stateA1_p & v84557c;
assign df519d = hmaster1_p & df519c | !hmaster1_p & df5185;
assign bd58a1 = hburst0 & bd589d | !hburst0 & bd58a0;
assign d357ce = hgrant1_p & d357c0 | !hgrant1_p & d357cd;
assign bd5788 = stateA1_p & ade4b8 | !stateA1_p & !d3594a;
assign v9f7cbc = hready & v9f7cbb | !hready & v9f7cb7;
assign v9ea602 = hmaster1_p & v9ea580 | !hmaster1_p & v9ea405;
assign v9ea621 = hlock3 & v9ea3fa | !hlock3 & v9ea620;
assign v898970 = hmaster0_p & v845558 | !hmaster0_p & !v9041a4;
assign d359a4 = hbusreq0 & d3599d | !hbusreq0 & d359a3;
assign v9f7712 = hmaster1_p & v9f7711 | !hmaster1_p & v9f7ce9;
assign v9ea606 = hgrant1_p & v9ea605 | !hgrant1_p & v9ea45c;
assign ad426e = hlock1_p & ad426c | !hlock1_p & ad426d;
assign ad5054 = hbusreq4_p & ad5051 | !hbusreq4_p & ad5053;
assign v9f7673 = hlock2 & v9f7670 | !hlock2 & v9f7672;
assign b1cfcb = hlock0_p & v84556e | !hlock0_p & !v845542;
assign ad3d38 = hgrant2_p & ad3d35 | !hgrant2_p & ad3d37;
assign v9f7766 = hlock2 & v9f7763 | !hlock2 & v9f7765;
assign v9ea5a3 = hbusreq1 & v9ea5a1 | !hbusreq1 & v9ea5a2;
assign ad4fc8 = stateA1_p & ad4fc7 | !stateA1_p & ad4fab;
assign ad43b9 = hready & ad43a8 | !hready & ad43b8;
assign ade58d = hlock0_p & ade586 | !hlock0_p & ade58c;
assign b05a2c = hgrant3_p & b05949 | !hgrant3_p & b05a2b;
assign df50d2 = decide_p & df50d1 | !decide_p & d6ebca;
assign ad4f6a = stateG10_4_p & ad4f67 | !stateG10_4_p & !ad4f69;
assign cc36ba = hmaster1_p & cc36b9 | !hmaster1_p & v845542;
assign c3d667 = stateA1_p & v845578 | !stateA1_p & !v889629;
assign ad4f42 = hbusreq2 & ad4f3c | !hbusreq2 & ad4f41;
assign d356b2 = hlock1_p & v845542 | !hlock1_p & dc4fcb;
assign ad4432 = hready & ad4429 | !hready & ad4431;
assign d3564f = hbusreq4_p & d3564e | !hbusreq4_p & !d3564d;
assign dc4ff4 = hgrant4_p & v845542 | !hgrant4_p & !ade557;
assign ad4f82 = hgrant4_p & v845542 | !hgrant4_p & !ad4f80;
assign ac147d = hmaster1_p & ac145d | !hmaster1_p & ac147c;
assign bd5ba4 = hmaster1_p & bd5ba3 | !hmaster1_p & v845542;
assign c3d705 = hbusreq2_p & c3d6fe | !hbusreq2_p & c3d704;
assign bd58ff = hbusreq2_p & bd58fe | !hbusreq2_p & !v845542;
assign c3d2ad = stateA1_p & v845578 | !stateA1_p & !v84557c;
assign c3d31d = hbusreq0 & c3d31c | !hbusreq0 & c3d30a;
assign d354ba = hbusreq1 & d35c01 | !hbusreq1 & !d35c03;
assign v8cc506 = hbusreq2_p & v8ccbfb | !hbusreq2_p & v8cc504;
assign d356dd = hbusreq1_p & d356dc | !hbusreq1_p & v845542;
assign v9ea5bc = hmaster0_p & v9ea567 | !hmaster0_p & v9f20a1;
assign cc36e0 = hgrant1_p & v845566 | !hgrant1_p & cc36de;
assign v9ea5e2 = hgrant2_p & v9ea5df | !hgrant2_p & v9ea5e1;
assign ad4849 = hgrant1_p & ad4848 | !hgrant1_p & ad4845;
assign b1c772 = hmaster2_p & b1c771 | !hmaster2_p & !b1cf29;
assign ad47ef = hmaster0_p & ad47ee | !hmaster0_p & ad46e8;
assign b05932 = hmaster0_p & b0591e | !hmaster0_p & b05920;
assign v9f7d60 = hbusreq4_p & v9ea3fb | !hbusreq4_p & v9f7d5d;
assign ac1487 = hgrant4_p & v845542 | !hgrant4_p & ac1486;
assign v8cc625 = hgrant2_p & v8cc472 | !hgrant2_p & v8cc624;
assign ad4f1b = hbusreq2 & ad4e95 | !hbusreq2 & !ad4f1a;
assign ad4281 = hlock1_p & ad4e95 | !hlock1_p & v845542;
assign ad48cb = hbusreq3_p & ad5071 | !hbusreq3_p & ad48ca;
assign v857b36 = stateG3_0_p & v845542 | !stateG3_0_p & v845580;
assign v8cc7a6 = hmaster1_p & v8cc7a5 | !hmaster1_p & v845542;
assign d354c8 = hbusreq1 & d35c0b | !hbusreq1 & v84555a;
assign v9f7dc1 = hgrant1_p & v9f7dbf | !hgrant1_p & v9f7dc0;
assign df51bd = hmaster0_p & df519b | !hmaster0_p & df517c;
assign bd58da = hbusreq2_p & bd58d9 | !hbusreq2_p & !v845542;
assign d35497 = hbusreq4_p & d35496 | !hbusreq4_p & v845542;
assign b574fa = hbusreq2_p & b574d1 | !hbusreq2_p & b574f9;
assign ad40f4 = hmaster0_p & ad40f2 | !hmaster0_p & ad40f3;
assign b1c6ca = hmaster1_p & b1d00e | !hmaster1_p & b1c6c9;
assign v9f782e = hmaster2_p & v9f781d | !hmaster2_p & !v9f782d;
assign v9f7d31 = hlock3 & v9f7d12 | !hlock3 & v9f7d19;
assign b57a1c = hmaster2_p & b57a1b | !hmaster2_p & v845542;
assign v9ea3fb = locked_p & v845542 | !locked_p & v9ea3ec;
assign d35698 = decide_p & d35697 | !decide_p & v84556c;
assign v8ccb69 = hmastlock_p & v8ccb68 | !hmastlock_p & v845542;
assign d35436 = hmaster2_p & v84555a | !hmaster2_p & d35435;
assign ade4b7 = hburst0_p & c74a04 | !hburst0_p & !ade4b6;
assign b1c745 = hmaster0_p & b1c740 | !hmaster0_p & b1c744;
assign v9ea4e2 = hbusreq2_p & v9ea4dd | !hbusreq2_p & v9ea4e1;
assign v8ccbda = hmaster1_p & v8ccbd9 | !hmaster1_p & v845542;
assign ad4d9d = hbusreq3 & ad4d9c | !hbusreq3 & v845542;
assign d35905 = stateG2_p & v845542 | !stateG2_p & adea85;
assign v9f7719 = hmaster0_p & v9f76ab | !hmaster0_p & v9f7691;
assign v9e9f8c = stateG10_4_p & v9e9f8a | !stateG10_4_p & v9e9f8b;
assign hgrant1 = !df51e0;
assign ade57b = hmaster2_p & ade559 | !hmaster2_p & ade57a;
assign ac145b = hbusreq4_p & ac1459 | !hbusreq4_p & ac145a;
assign d354f0 = hmaster1_p & d354ef | !hmaster1_p & d35410;
assign ad445e = hmaster2_p & ad445d | !hmaster2_p & v845542;
assign ad4f22 = hmaster0_p & ad4f20 | !hmaster0_p & !ad4f21;
assign ad4dce = hlock0_p & ad4dc4 | !hlock0_p & v845542;
assign d35a30 = hbusreq1_p & d35a2f | !hbusreq1_p & !d35a2e;
assign b1c7dd = stateG10_4_p & b1c7bc | !stateG10_4_p & b1c7dc;
assign bd58a8 = stateG10_4_p & bd58a5 | !stateG10_4_p & !bd58a7;
assign d354e8 = hmaster1_p & d354e7 | !hmaster1_p & d354d3;
assign b06719 = stateG2_p & v845542 | !stateG2_p & c6d407;
assign v9ea5e9 = hready_p & v9ea436 | !hready_p & v9ea5e8;
assign bd5e9e = hbusreq4_p & bd5e9d | !hbusreq4_p & v845542;
assign d35a72 = hbusreq1_p & d35a71 | !hbusreq1_p & !v845542;
assign cc36c4 = hgrant1_p & df54f3 | !hgrant1_p & d35a49;
assign b574d6 = hbusreq2 & b574d5 | !hbusreq2 & b57942;
assign df51c7 = hmaster1_p & df51c3 | !hmaster1_p & df51c6;
assign ad4264 = hmaster2_p & v84556c | !hmaster2_p & ad4ef3;
assign v9f786b = hbusreq1_p & v9f7758 | !hbusreq1_p & v9f7864;
assign v9e9f59 = hlock4 & v9e9f57 | !hlock4 & v9e9f58;
assign dc5012 = hmaster2_p & dc4ff6 | !hmaster2_p & dc5011;
assign ad4845 = hready & ad4d96 | !hready & !ad4844;
assign v9f7d68 = hbusreq2_p & v9f7d65 | !hbusreq2_p & v9f7d67;
assign c3d328 = hmaster2_p & c3d327 | !hmaster2_p & c3d2fd;
assign c3d6c0 = hbusreq1_p & c3d67b | !hbusreq1_p & !c3d68a;
assign c3d32a = hbusreq4 & c3d311 | !hbusreq4 & !c3d329;
assign c3d51e = hmaster1_p & c3d51a | !hmaster1_p & c3d51d;
assign d35621 = hbusreq3 & d3560e | !hbusreq3 & d35620;
assign b1c086 = hbusreq0 & b1c085 | !hbusreq0 & b1c85e;
assign bd5e25 = hbusreq2_p & bd5e22 | !hbusreq2_p & v845542;
assign b1c78d = hmaster0_p & b1c78b | !hmaster0_p & b1c78c;
assign c3d5e1 = hgrant4_p & v845542 | !hgrant4_p & c3d5d9;
assign ad4e52 = hready & d35980 | !hready & v84556c;
assign v9f7698 = hmaster2_p & v9f768f | !hmaster2_p & !v9f7697;
assign v9e9e71 = hbusreq3_p & v9ea619 | !hbusreq3_p & v9e9e70;
assign ad434a = hready_p & ad432a | !hready_p & ad4349;
assign c3d355 = hmaster0_p & c3d351 | !hmaster0_p & c3d354;
assign b579eb = hgrant2_p & b579b0 | !hgrant2_p & b579ea;
assign v9f76b2 = hgrant3_p & v9f7d6a | !hgrant3_p & v9f76b1;
assign d35585 = hbusreq1 & d354f3 | !hbusreq1 & !d35a9b;
assign ad4fa6 = hmaster0_p & ad4f54 | !hmaster0_p & ad4fa5;
assign bd5772 = hbusreq3 & bd5771 | !hbusreq3 & !v845542;
assign ad4fc0 = hbusreq3 & ad4fbf | !hbusreq3 & v845542;
assign ad4471 = hbusreq1_p & ad4470 | !hbusreq1_p & ad40fe;
assign ad4377 = decide_p & ad42ce | !decide_p & ad4348;
assign v9f7cd0 = hbusreq1_p & v9f7cbe | !hbusreq1_p & v9f7ccf;
assign b05a75 = hlock3 & b05a74 | !hlock3 & b05a72;
assign d355af = hlock3_p & d355ae | !hlock3_p & v845552;
assign c3d342 = hmaster2_p & c3d341 | !hmaster2_p & v845576;
assign v9f7cbf = hlock3 & v9f7cb7 | !hlock3 & v9f7cbe;
assign d35800 = hmaster0_p & d357f8 | !hmaster0_p & d357ff;
assign d35909 = hburst0 & d35907 | !hburst0 & d35908;
assign d354b0 = hgrant0_p & v84556c | !hgrant0_p & !d354af;
assign df5191 = hbusreq1 & dc4fe0 | !hbusreq1 & v845542;
assign v9f76ee = hlock0_p & v9f7d81 | !hlock0_p & v9f76ed;
assign d35a3d = hmastlock_p & d35a3b | !hmastlock_p & v845542;
assign d359da = hmaster2_p & d359a2 | !hmaster2_p & d359d9;
assign c3d2c9 = hbusreq3 & c3d2c7 | !hbusreq3 & v845542;
assign bd5797 = hbusreq2 & bd5796 | !hbusreq2 & v845564;
assign df50d4 = hready_p & df50d2 | !hready_p & df50d3;
assign v9f7869 = hlock2 & v9f7866 | !hlock2 & v9f7868;
assign b1d012 = hmaster1_p & b1d00e | !hmaster1_p & b1d011;
assign d35a49 = hbusreq4_p & d35a48 | !hbusreq4_p & !dc500f;
assign v9e9f79 = hmaster2_p & v9e9f56 | !hmaster2_p & v9e9f77;
assign d3576b = jx1_p & d3575c | !jx1_p & d3576a;
assign v9ea583 = hmaster0_p & v9ea582 | !hmaster0_p & v9ea578;
assign v9ea3f6 = hmaster0_p & v9ea3f5 | !hmaster0_p & v9ea3e7;
assign ade590 = hgrant0_p & ade58f | !hgrant0_p & v84556c;
assign v8cc50f = hbusreq3_p & v8cc4df | !hbusreq3_p & v8cc50e;
assign v9f771b = hgrant2_p & v9f7718 | !hgrant2_p & v9f771a;
assign v8cc5ba = hmaster1_p & v8cc475 | !hmaster1_p & v8cc5b9;
assign b1c7e7 = hbusreq2 & b1c733 | !hbusreq2 & !b1c736;
assign ad41a8 = hmaster1_p & ad41a4 | !hmaster1_p & ad41a7;
assign ad4160 = hbusreq2 & ad415f | !hbusreq2 & v845542;
assign d357f1 = decide_p & d357f0 | !decide_p & v84556c;
assign c3d729 = hmaster1_p & c3d685 | !hmaster1_p & c3d68b;
assign v9ea5a0 = hbusreq4 & v9ea59f | !hbusreq4 & v9ea59b;
assign c3d6a4 = hbusreq1_p & c3d671 | !hbusreq1_p & !c3d683;
assign v9f7745 = hmaster2_p & v9f772a | !hmaster2_p & v84557a;
assign b059ff = hmaster1_p & b059fe | !hmaster1_p & b059f5;
assign b1c5eb = hmaster2_p & b1cfbf | !hmaster2_p & b1c5ea;
assign v9ea436 = decide_p & v9ea42b | !decide_p & v9ea435;
assign adeca1 = locked_p & v845542 | !locked_p & !adeca0;
assign bd5ea5 = hmaster1_p & bd5ea4 | !hmaster1_p & v84556c;
assign v8cc4ac = hgrant1_p & v845542 | !hgrant1_p & v8cc4ab;
assign ad433a = hbusreq1 & ad5021 | !hbusreq1 & ad5023;
assign v8cc4a6 = hlock4 & v8cc49d | !hlock4 & v8cc4a5;
assign ad4600 = hmaster0_p & ad45ff | !hmaster0_p & ad45c2;
assign d35689 = hbusreq2_p & v845552 | !hbusreq2_p & !v845542;
assign dc538d = hmaster2_p & v84556c | !hmaster2_p & !dc538c;
assign dc5000 = stateG10_4_p & adec89 | !stateG10_4_p & dc4fff;
assign b574f9 = hgrant2_p & b574d8 | !hgrant2_p & b574d0;
assign df54fd = hgrant2_p & v845542 | !hgrant2_p & !df54fc;
assign c5c894 = stateG2_p & v845542 | !stateG2_p & bb9bdd;
assign v8cc121 = hready_p & v8cc455 | !hready_p & v8cc120;
assign ad440f = hmaster2_p & b1c714 | !hmaster2_p & b1c70e;
assign dc5320 = hready_p & dc5315 | !hready_p & !dc531f;
assign v9f76fe = hlock3 & v9f76fd | !hlock3 & v9f76fb;
assign v8cc81f = decide_p & v845542 | !decide_p & v8cc81e;
assign ad4dec = hbusreq0 & ad4dde | !hbusreq0 & ad4deb;
assign c3ce90 = hmaster0_p & c3ce8f | !hmaster0_p & c3d2be;
assign v8cc4dc = decide_p & v8ccbd7 | !decide_p & v8cc4db;
assign ade56e = hbusreq4_p & ade56d | !hbusreq4_p & !v845542;
assign b57959 = hgrant2_p & b57948 | !hgrant2_p & b57958;
assign c3ceee = hlock0_p & c3d5b2 | !hlock0_p & c3ceed;
assign d35012 = hmaster2_p & d3580a | !hmaster2_p & d35011;
assign d354ab = hbusreq0 & d354a7 | !hbusreq0 & d354aa;
assign ad43d3 = hready & ad43c8 | !hready & !ad43d2;
assign c3d2b2 = hready & c3d2b1 | !hready & v845542;
assign v9f7cce = hlock1 & v9f7cc8 | !hlock1 & v9f7ccd;
assign b57423 = hready & b57422 | !hready & b57987;
assign ad46fd = hgrant4_p & v845542 | !hgrant4_p & cc36fc;
assign v9e9eef = hbusreq4_p & v9ea3fb | !hbusreq4_p & v9e9eec;
assign bd5790 = hburst0 & d3561d | !hburst0 & bd578f;
assign aa425d = jx0_p & v845542 | !jx0_p & aa425c;
assign d355a3 = hmaster2_p & v84556c | !hmaster2_p & d35a58;
assign b1c45e = hgrant3_p & b1cb00 | !hgrant3_p & b1c45d;
assign ad4f24 = hgrant2_p & ad4f23 | !hgrant2_p & !ad4f17;
assign b57983 = hgrant1_p & b578f1 | !hgrant1_p & b5794a;
assign d359b5 = hmastlock_p & v845542 | !hmastlock_p & d359b4;
assign b1c85a = hgrant1_p & b1d01a | !hgrant1_p & b1c859;
assign df54ea = hmaster0_p & df54e9 | !hmaster0_p & v845542;
assign ad4ee4 = hgrant4_p & ad4e5c | !hgrant4_p & ad4ee3;
assign c3d6d9 = hmaster0_p & c3d683 | !hmaster0_p & c3d6b5;
assign ad4814 = hmaster2_p & v845542 | !hmaster2_p & ad4f38;
assign c3cf21 = hmaster0_p & c3cf20 | !hmaster0_p & !c3d2be;
assign b059c3 = hmaster2_p & b058a3 | !hmaster2_p & b059c2;
assign d35762 = hgrant3_p & d3575e | !hgrant3_p & d35761;
assign v9ea463 = locked_p & v845542 | !locked_p & !v9ea3e9;
assign d356a1 = hbusreq1_p & d356a0 | !hbusreq1_p & v845542;
assign v8cc5fb = hbusreq2 & v8cc5f8 | !hbusreq2 & v8cc5f9;
assign v9f76e5 = hlock0_p & v9f7d70 | !hlock0_p & v9f76e4;
assign c3d585 = hbusreq2_p & c3d508 | !hbusreq2_p & c3d584;
assign ad4e46 = hmastlock_p & ad4e45 | !hmastlock_p & v845542;
assign d35706 = hgrant1_p & d35aa4 | !hgrant1_p & d35705;
assign d35770 = hmaster2_p & d3576e | !hmaster2_p & d3576f;
assign v9e9fbb = hmaster0_p & v9e9fb8 | !hmaster0_p & v9e9eed;
assign b57419 = hbusreq4_p & b5794f | !hbusreq4_p & b57418;
assign v9ea60d = hbusreq2 & v9ea60c | !hbusreq2 & v9ea486;
assign df516c = hbusreq2_p & df5164 | !hbusreq2_p & df516b;
assign d3579f = hbusreq0 & d3579e | !hbusreq0 & v845542;
assign v9e9ed6 = decide_p & v9ea4b2 | !decide_p & v9e9ed5;
assign ac146e = hgrant2_p & ac1456 | !hgrant2_p & ac146d;
assign ad4fd2 = hbusreq1_p & ad4fc2 | !hbusreq1_p & ad4fc1;
assign b1c6fe = decide_p & b1c6fd | !decide_p & b1c6cb;
assign v9f21c5 = locked_p & v9f21c4 | !locked_p & v845542;
assign v9e9edc = decide_p & v9e9e75 | !decide_p & v9e9edb;
assign ad4fd9 = hgrant0_p & ad4fae | !hgrant0_p & !v845542;
assign dc5088 = hgrant3_p & v84556a | !hgrant3_p & v845542;
assign c3d303 = hbusreq0 & v845542 | !hbusreq0 & adeaa5;
assign d35a4c = hbusreq3 & d35a4b | !hbusreq3 & v845542;
assign ad4efd = hgrant4_p & ad4ef3 | !hgrant4_p & v845542;
assign ad455f = hbusreq4 & ad455a | !hbusreq4 & ad455e;
assign ac1456 = hmaster1_p & ac1455 | !hmaster1_p & v845542;
assign v8da604 = hgrant3_p & v8da59e | !hgrant3_p & v8da603;
assign v9f7e0e = hmaster0_p & v9f7d9f | !hmaster0_p & v9f7e0d;
assign v9ea488 = hlock2 & v9ea486 | !hlock2 & v9ea487;
assign ad43a7 = hmaster2_p & b1c70e | !hmaster2_p & v845542;
assign v9f7cf1 = hbusreq2_p & v9f7cea | !hbusreq2_p & v9f7cf0;
assign ad4307 = hmaster1_p & ad4306 | !hmaster1_p & ad4300;
assign v9f7ce2 = hready & v9f7ce1 | !hready & v9f7cdd;
assign c3d381 = hmaster0_p & c3d380 | !hmaster0_p & !c3d2be;
assign bd5b97 = hmaster0_p & v84556c | !hmaster0_p & bd5b96;
assign c3d350 = hgrant1_p & v84554d | !hgrant1_p & c3d34f;
assign d35795 = hbusreq2 & d3578d | !hbusreq2 & d35794;
assign d35631 = hlock3_p & d3562d | !hlock3_p & d35630;
assign b1cf3a = hmaster2_p & v845542 | !hmaster2_p & d3591a;
assign v9ea47b = hmaster2_p & v9ea479 | !hmaster2_p & v9ea473;
assign ad41a1 = hbusreq3 & ad5027 | !hbusreq3 & ad502a;
assign c3d393 = decide_p & c3d392 | !decide_p & !c3d36c;
assign dc4f88 = hmaster0_p & dc4f67 | !hmaster0_p & dc4f87;
assign c3d71c = hmaster0_p & c3d6b5 | !hmaster0_p & c3d683;
assign ad4de5 = hbusreq2 & ad4de0 | !hbusreq2 & ad4de4;
assign d354b7 = hbusreq4 & d354ab | !hbusreq4 & d354b6;
assign ad3d10 = hready & ad3d0a | !hready & ad3d0f;
assign d35759 = decide_p & d35758 | !decide_p & v84556c;
assign v8cc76b = hbusreq2 & v8cc769 | !hbusreq2 & v8ccbd8;
assign c3d719 = decide_p & c3d695 | !decide_p & c3d718;
assign c3d703 = hmaster1_p & c3d702 | !hmaster1_p & c3d6fc;
assign b57403 = hready_p & b57a2e | !hready_p & b57402;
assign c3d72b = hmaster0_p & c3d685 | !hmaster0_p & c3d697;
assign d35021 = hbusreq2_p & d357e2 | !hbusreq2_p & d35020;
assign d357d3 = hgrant1_p & d357d1 | !hgrant1_p & d357cd;
assign v9f783b = hbusreq3 & v9f7837 | !hbusreq3 & v9f783a;
assign ad3cfa = hbusreq0 & ad3cf9 | !hbusreq0 & v845542;
assign d356db = hbusreq1 & d35910 | !hbusreq1 & v845542;
assign v9e9e73 = jx0_p & v9ea4e6 | !jx0_p & v9e9e72;
assign b57432 = hmaster0_p & v845542 | !hmaster0_p & b57431;
assign c3ce83 = hmaster0_p & c3ce82 | !hmaster0_p & c3ce4d;
assign ad5051 = hgrant4_p & ad5048 | !hgrant4_p & v84556c;
assign ad4314 = hbusreq1_p & ad4313 | !hbusreq1_p & v845542;
assign v84557a = stateA1_p & v845542 | !stateA1_p & !v845542;
assign ac1469 = hbusreq4_p & ac1467 | !hbusreq4_p & !ac1468;
assign ad431e = hgrant2_p & ad4312 | !hgrant2_p & ad431d;
assign ad4ff0 = hgrant2_p & ad4fb9 | !hgrant2_p & ad4fef;
assign d3597e = hready_p & d358e8 | !hready_p & d3597d;
assign ac144f = hmaster2_p & v845542 | !hmaster2_p & !ac144e;
assign c5c930 = hmaster2_p & v845542 | !hmaster2_p & c5c92f;
assign ad4f00 = hlock0_p & ad4e4c | !hlock0_p & !v845542;
assign v9f7838 = hbusreq1_p & v9f77c8 | !hbusreq1_p & v9f782f;
assign b1c084 = hbusreq4_p & b1c7db | !hbusreq4_p & !b1c083;
assign d35507 = decide_p & d35506 | !decide_p & !v84556c;
assign d35aab = hgrant4_p & v845542 | !hgrant4_p & !d35aaa;
assign ad4754 = hbusreq2_p & ad4750 | !hbusreq2_p & ad4753;
assign b5740d = hbusreq4 & b5740b | !hbusreq4 & b5740c;
assign b059e0 = stateG10_4_p & v9f7d42 | !stateG10_4_p & !b059df;
assign b579d3 = hmaster2_p & b579cb | !hmaster2_p & b579d2;
assign v9ea48d = hmaster2_p & v9ea439 | !hmaster2_p & v9ea44d;
assign ad4d9f = hmaster0_p & ad4d94 | !hmaster0_p & ad4d9e;
assign d354bf = hbusreq1_p & d354bb | !hbusreq1_p & !d354be;
assign ad43a2 = hmaster1_p & ad43a1 | !hmaster1_p & ad4f1a;
assign v9f7d11 = hmaster0_p & v9f7d03 | !hmaster0_p & v9f7d10;
assign v9e9fa2 = hbusreq1 & v9e9f6f | !hbusreq1 & v9e9f70;
assign v9f7dcb = hgrant4_p & v9f7cf5 | !hgrant4_p & v9f7c9f;
assign c3d57d = hbusreq0 & c3d57c | !hbusreq0 & v845542;
assign d359d1 = hlock4_p & d359cf | !hlock4_p & d359d0;
assign b57a73 = hbusreq2 & b57a71 | !hbusreq2 & b57a72;
assign v9ea577 = hbusreq4_p & v9ea403 | !hbusreq4_p & v9ea4bb;
assign ad4f76 = hbusreq4_p & ad4f75 | !hbusreq4_p & ad4f67;
assign v9ea5a6 = hlock3 & v9ea5a5 | !hlock3 & v9ea5a4;
assign v9f77e8 = hgrant4_p & d359c4 | !hgrant4_p & v9f772f;
assign c5c9b0 = hmaster1_p & c5c9af | !hmaster1_p & c5c8eb;
assign ad5039 = hbusreq3 & ad5037 | !hbusreq3 & ad5038;
assign ad481c = hbusreq2 & v845547 | !hbusreq2 & v845542;
assign d35a74 = hgrant1_p & d35a72 | !hgrant1_p & d35a73;
assign b1c052 = hgrant2_p & b1c04f | !hgrant2_p & b1c051;
assign v9ea3e9 = hmastlock_p & v845582 | !hmastlock_p & !v845542;
assign c3d6e8 = hgrant1_p & c3d671 | !hgrant1_p & c3d6e7;
assign v9f7652 = hgrant4_p & v9f7ca0 | !hgrant4_p & v9f7d78;
assign ad4404 = hmaster0_p & ad4403 | !hmaster0_p & ad43d7;
assign v9ea448 = hbusreq4_p & v9ea446 | !hbusreq4_p & v9ea447;
assign ad42f6 = hlock1_p & ad42f4 | !hlock1_p & ad42f5;
assign d355a0 = hready_p & d35596 | !hready_p & d3559f;
assign b57a82 = hmaster1_p & b579b4 | !hmaster1_p & b57a81;
assign d35a65 = hgrant4_p & v84556c | !hgrant4_p & !d35a64;
assign bd58b5 = hmaster0_p & bd58b0 | !hmaster0_p & bd58b4;
assign v8cc82a = hmaster1_p & v8cc500 | !hmaster1_p & v8cc829;
assign ad46d5 = hlock0_p & ad455b | !hlock0_p & !v845542;
assign ba7c6d = hmaster0_p & ba7c6b | !hmaster0_p & ba7c6c;
assign ad502d = hmaster0_p & ad5025 | !hmaster0_p & ad502c;
assign ad4e1f = hbusreq2_p & ad4df8 | !hbusreq2_p & ad4e0b;
assign d35ab8 = hgrant2_p & v845542 | !hgrant2_p & !d35ab7;
assign b1c7c8 = hbusreq0 & b1c7c7 | !hbusreq0 & b1cfcc;
assign c5c9ac = hmaster0_p & c5c8e9 | !hmaster0_p & c5c8e8;
assign v8cc768 = hbusreq3 & v8cc765 | !hbusreq3 & v8cc766;
assign ad4e7c = hgrant4_p & v845542 | !hgrant4_p & ad4e6f;
assign c3ce5d = hbusreq1 & c3d2d6 | !hbusreq1 & v845564;
assign adeab4 = hgrant2_p & v845542 | !hgrant2_p & adea95;
assign v9f7df8 = hmaster1_p & v9f7d9f | !hmaster1_p & v9f7df7;
assign v845576 = hgrant4_p & v845542 | !hgrant4_p & !v845542;
assign ad4332 = hbusreq1 & ad5029 | !hbusreq1 & ad5023;
assign v845570 = hgrant1_p & v845542 | !hgrant1_p & !v845542;
assign b1c7ac = hmaster2_p & b1c7a7 | !hmaster2_p & b1c7ab;
assign b574d8 = hmaster1_p & b574d7 | !hmaster1_p & v845542;
assign d35701 = hbusreq1_p & d35700 | !hbusreq1_p & v845542;
assign d35724 = hready_p & d35723 | !hready_p & d356f1;
assign ad4152 = hgrant4_p & v845542 | !hgrant4_p & ad4f38;
assign ad42d7 = hbusreq1 & ad501b | !hbusreq1 & v845542;
assign ad4f54 = hbusreq3 & ad4f53 | !hbusreq3 & v845542;
assign ad4ddd = hmaster2_p & v845542 | !hmaster2_p & !v9c81a4;
assign b8f74a = hmaster0_p & b8f6e1 | !hmaster0_p & b8f749;
assign c3d74e = hmaster1_p & c3d74d | !hmaster1_p & c3d6fc;
assign v9ea480 = hlock4 & v9ea46d | !hlock4 & v9ea476;
assign dc4fcb = hmaster2_p & v84556c | !hmaster2_p & v845542;
assign dc4f94 = hmaster1_p & dc4f88 | !hmaster1_p & dc4f93;
assign b574b9 = hbusreq1 & b574b8 | !hbusreq1 & b57942;
assign ad42d0 = hbusreq1 & ad5018 | !hbusreq1 & c3d2d9;
assign ad414c = hbusreq1 & ad4815 | !hbusreq1 & ad4f40;
assign d35441 = hlock2_p & d3543f | !hlock2_p & d35440;
assign v9e9f53 = hmaster2_p & v9e9f52 | !hmaster2_p & v9ea448;
assign b059ec = hready & b059eb | !hready & b059e7;
assign bd580e = hgrant4_p & adec89 | !hgrant4_p & bd580d;
assign bd593f = hgrant3_p & bd592d | !hgrant3_p & !bd593e;
assign ad4ea9 = hbusreq3 & ad4ea8 | !hbusreq3 & v845542;
assign b57ae6 = hbusreq3 & b579e4 | !hbusreq3 & b57ae5;
assign bd5bb0 = decide_p & bd5ba6 | !decide_p & !v845572;
assign bbb7c7 = hburst0_p & v845542 | !hburst0_p & bbb7c6;
assign v9e9ee7 = hlock0_p & v845542 | !hlock0_p & v9ea3e6;
assign v9f7843 = hbusreq4_p & v9f7841 | !hbusreq4_p & !v9f7842;
assign v9ea499 = hmaster1_p & v9ea498 | !hmaster1_p & v9ea43f;
assign b1c02f = hlock0_p & b1c754 | !hlock0_p & b1c02e;
assign d35a61 = hbusreq4_p & d35a60 | !hbusreq4_p & !d35a5f;
assign b059eb = hbusreq4 & b059e9 | !hbusreq4 & b059ea;
assign v9ea4bd = hmaster0_p & v9ea4b8 | !hmaster0_p & v9ea4bc;
assign c3d69a = hbusreq1_p & c3d697 | !hbusreq1_p & c3d699;
assign ad4db8 = hbusreq3 & ad4db7 | !hbusreq3 & v845542;
assign dc4fef = hgrant4_p & v845542 | !hgrant4_p & !ade553;
assign v9f788a = hbusreq4 & v9f7888 | !hbusreq4 & v9f7889;
assign v9f7889 = hlock4 & v9f77d8 | !hlock4 & v9f7888;
assign v9ea427 = hgrant2_p & v9ea40d | !hgrant2_p & v9ea426;
assign ad4356 = hbusreq2_p & ad4353 | !hbusreq2_p & ad4355;
assign dc5037 = locked_p & dc5036 | !locked_p & c3d66d;
assign d35628 = hmaster2_p & adea8a | !hmaster2_p & !d35627;
assign c3d5c2 = hbusreq4 & c3d5bc | !hbusreq4 & !c3d5c1;
assign c3d68b = hmaster0_p & c3d686 | !hmaster0_p & c3d68a;
assign b1c06a = hmaster2_p & b1c065 | !hmaster2_p & b1c069;
assign c3d34f = hready & c3d34e | !hready & c3d313;
assign d354ed = hgrant3_p & d35445 | !hgrant3_p & d354ec;
assign v9f7713 = hmaster1_p & v9f7683 | !hmaster1_p & v9f7675;
assign d358f9 = hburst0 & d358eb | !hburst0 & d358f8;
assign b1c044 = hmaster2_p & b1c043 | !hmaster2_p & !b1c844;
assign c3d723 = hmaster0_p & c3d6e9 | !hmaster0_p & c3d676;
assign dc5044 = stateG10_4_p & ade563 | !stateG10_4_p & !dc5043;
assign dc5066 = hbusreq3 & dc5065 | !hbusreq3 & v845542;
assign c3d4ff = hbusreq0 & c3d4fe | !hbusreq0 & v845542;
assign d35513 = hbusreq1 & d35421 | !hbusreq1 & d35512;
assign v9f7c9f = hmastlock_p & v9f7c9e | !hmastlock_p & !v845542;
assign d35656 = hbusreq4_p & d35655 | !hbusreq4_p & !d35654;
assign b57af0 = hlock3 & b57942 | !hlock3 & b579ec;
assign d35505 = hmaster1_p & d354fb | !hmaster1_p & d35504;
assign ad429b = hbusreq2_p & ad4298 | !hbusreq2_p & ad429a;
assign v9f7e25 = hlock1 & v9f7e1f | !hlock1 & v9f7e24;
assign v9ea5ca = hbusreq2_p & v9ea5bd | !hbusreq2_p & v9ea5be;
assign ade54c = stateA1_p & v845542 | !stateA1_p & !ade54b;
assign v9f765d = hgrant4_p & v9f7ca6 | !hgrant4_p & v9f7d89;
assign b1c055 = hmaster1_p & b1c054 | !hmaster1_p & b1c7eb;
assign ad4777 = hbusreq0 & ad45e5 | !hbusreq0 & ad4776;
assign v9f7d42 = hmastlock_p & v9f7d41 | !hmastlock_p & !v845542;
assign df5176 = hbusreq2 & df5146 | !hbusreq2 & df5148;
assign v9f767c = hmaster0_p & v9f7cc2 | !hmaster0_p & v9f767b;
assign v9ea45d = hgrant1_p & v9ea456 | !hgrant1_p & v9ea45c;
assign d3574a = hmaster0_p & d35748 | !hmaster0_p & d35749;
assign ad4f2b = hbusreq1 & ad4f1e | !hbusreq1 & !v845542;
assign ad4f96 = hgrant4_p & v845542 | !hgrant4_p & ad4f88;
assign c3d50a = hgrant1_p & v84554d | !hgrant1_p & c3d503;
assign ad42eb = hbusreq1 & ad4f57 | !hbusreq1 & v845542;
assign d35910 = hmaster2_p & d35909 | !hmaster2_p & !dc5318;
assign v9f7d06 = hlock0 & v9f7d05 | !hlock0 & v9f7d04;
assign d359e1 = hbusreq4 & d359db | !hbusreq4 & d359e0;
assign b1c7f2 = hbusreq1 & b1c722 | !hbusreq1 & b1c71d;
assign b579e8 = hbusreq2 & b579e6 | !hbusreq2 & b579e7;
assign b1d002 = hbusreq0 & b1cff7 | !hbusreq0 & b1d001;
assign v9f76f3 = hlock0 & v9f76f2 | !hlock0 & v9f76e9;
assign v8ccb88 = hbusreq2_p & v8ccb87 | !hbusreq2_p & v8ccb84;
assign v9e9ece = hmaster0_p & v9e9eba | !hmaster0_p & v9e9ea1;
assign v9f7697 = hbusreq4_p & v9f7695 | !hbusreq4_p & v9f7696;
assign v9f7723 = hgrant3_p & v9f76d2 | !hgrant3_p & v9f7722;
assign v9f76ae = hgrant2_p & v9f76aa | !hgrant2_p & v9f76ad;
assign cc370b = hbusreq3_p & cc36ee | !hbusreq3_p & !cc370a;
assign v9f21c4 = hmastlock_p & v9c81a4 | !hmastlock_p & v845542;
assign b059a0 = hmaster0_p & b05975 | !hmaster0_p & b0599f;
assign ad4488 = hgrant1_p & ad43ab | !hgrant1_p & ad4487;
assign v9f7cf7 = locked_p & v9f7cf2 | !locked_p & v9ea3ec;
assign dc4fc4 = hgrant2_p & dc4fc1 | !hgrant2_p & dc4fc3;
assign c3cef7 = hbusreq4 & c3cef3 | !hbusreq4 & !c3cef6;
assign bd588b = hlock4_p & bd5889 | !hlock4_p & !bd588a;
assign v9f769c = locked_p & v845542 | !locked_p & !v9f7d42;
assign b1cbf6 = hbusreq0 & b1cbf2 | !hbusreq0 & b1cbf5;
assign v9e9ef0 = hmaster2_p & v9e9eef | !hmaster2_p & v9ea4bb;
assign v9f7674 = hbusreq2 & v9f7672 | !hbusreq2 & v9f7673;
assign ad4559 = hbusreq4_p & ad4558 | !hbusreq4_p & v845542;
assign ad468f = hbusreq1 & ad4586 | !hbusreq1 & !v845542;
assign b1cfc8 = hbusreq0 & b1cfc3 | !hbusreq0 & b1cfc7;
assign v9f76a6 = hmaster0_p & v9f769a | !hmaster0_p & !v9f76a5;
assign v9ea5aa = hmaster0_p & v9ea599 | !hmaster0_p & v9ea5a9;
assign v845550 = hbusreq2_p & v845542 | !hbusreq2_p & !v845542;
assign v8cc7b0 = hlock1_p & v8cc79e | !hlock1_p & v845542;
assign b578ff = hlock0_p & b578f9 | !hlock0_p & v845542;
assign v8cc7bb = hbusreq4_p & v8cc7ba | !hbusreq4_p & v845542;
assign v8cc7ab = hmaster0_p & v845542 | !hmaster0_p & v8cc7a2;
assign v9f769f = stateG10_4_p & v9f769d | !stateG10_4_p & v9f769e;
assign adec9c = hmaster2_p & adec93 | !hmaster2_p & adec9b;
assign bd58e6 = hgrant3_p & bd57f0 | !hgrant3_p & !bd58e5;
assign ad41b6 = hmaster1_p & ad41b5 | !hmaster1_p & ad40f7;
assign v9f7773 = hmaster0_p & v9f774f | !hmaster0_p & v9f7772;
assign v9f781b = hgrant4_p & v9f7785 | !hgrant4_p & v9f781a;
assign b05a6c = hlock4 & b05a69 | !hlock4 & b05a6b;
assign c5c902 = hmaster1_p & c5c8f5 | !hmaster1_p & c5c901;
assign v9f7cfb = hlock4 & v9f7cf8 | !hlock4 & v9f7cfa;
assign c3d3a6 = hmaster0_p & c3d3a5 | !hmaster0_p & c3d395;
assign c3d479 = hready & c3d478 | !hready & v845542;
assign v9ea41e = hgrant0_p & v9ea41d | !hgrant0_p & v845542;
assign ade651 = hgrant3_p & ade63e | !hgrant3_p & ade650;
assign c3cf11 = hgrant2_p & c3d36c | !hgrant2_p & c3cf10;
assign c3d2f2 = hbusreq4_p & c3d2f0 | !hbusreq4_p & !c3d2f1;
assign d357da = hbusreq4_p & d357d7 | !hbusreq4_p & d357ca;
assign d35be8 = hbusreq4_p & d35be7 | !hbusreq4_p & v845542;
assign ade4c0 = hbusreq4_p & ade4bf | !hbusreq4_p & v845542;
assign b05a50 = hmaster1_p & b05a4f | !hmaster1_p & b059a0;
assign v8cc819 = decide_p & v8ccbd7 | !decide_p & v8cc50a;
assign ad4f68 = hgrant4_p & ad4f4a | !hgrant4_p & ad4f67;
assign b1c061 = hbusreq0_p & bd58a2 | !hbusreq0_p & v845542;
assign ad4481 = stateG10_4_p & c3cec2 | !stateG10_4_p & ad4480;
assign ade5c3 = hmaster1_p & ade5bf | !hmaster1_p & ade5c2;
assign ad442b = hbusreq4_p & ad442a | !hbusreq4_p & b1cfcd;
assign b1cf45 = hgrant2_p & b1cf43 | !hgrant2_p & b1cf3d;
assign ad4feb = hready & ad4fe0 | !hready & ad4fea;
assign d3569a = hgrant3_p & d3568d | !hgrant3_p & d35699;
assign dc53cf = hready_p & v845542 | !hready_p & dc53ce;
assign v9f7ddd = hgrant0_p & v9f7ca6 | !hgrant0_p & v9ea3ec;
assign ad46fc = hmaster1_p & ad46fb | !hmaster1_p & ad45a5;
assign ad46ba = hbusreq0 & ad46b9 | !hbusreq0 & ad4695;
assign b1c08a = hmaster0_p & b1c07a | !hmaster0_p & b1c089;
assign b05954 = hlock0_p & b05953 | !hlock0_p & v9f7d42;
assign df514c = hbusreq3 & df514b | !hbusreq3 & df5142;
assign ad4e9a = hgrant4_p & v845542 | !hgrant4_p & !ad4e98;
assign ad3cf1 = hready & ad3cf0 | !hready & !v845542;
assign dc531f = decide_p & dc531e | !decide_p & !v845542;
assign c3cecd = hmaster2_p & c3cecc | !hmaster2_p & v845542;
assign c5c96f = hgrant4_p & c5c8e7 | !hgrant4_p & c5c96e;
assign b1c7c6 = hbusreq4_p & b1c7c3 | !hbusreq4_p & !b1c7c5;
assign b1c7f9 = hbusreq2_p & b1c7ee | !hbusreq2_p & b1c7f8;
assign v8cc5c2 = hmaster0_p & v845542 | !hmaster0_p & v8cc5c1;
assign ad4343 = hbusreq1 & ad5034 | !hbusreq1 & c3d2d9;
assign ad4571 = hbusreq3 & ad4570 | !hbusreq3 & v845542;
assign b57b5b = jx1_p & b57abc | !jx1_p & b57b5a;
assign ad3d5c = hgrant3_p & ad3d32 | !hgrant3_p & ad3d5b;
assign ad4478 = hmaster1_p & ad4477 | !hmaster1_p & ad43ba;
assign ad4fbf = hgrant1_p & dc4fcb | !hgrant1_p & ad4fbe;
assign bd585e = hgrant4_p & bd5838 | !hgrant4_p & !bd574e;
assign b1c7d4 = hbusreq4_p & b1c7d1 | !hbusreq4_p & !b1c7d3;
assign c3cf26 = decide_p & c3cf23 | !decide_p & c3cf25;
assign ad3d45 = hgrant2_p & ad3d42 | !hgrant2_p & ad3d44;
assign ad4295 = hbusreq1 & ad4fb6 | !hbusreq1 & v845542;
assign bd5927 = hbusreq2 & dc5394 | !hbusreq2 & bd5926;
assign b1c6b9 = hlock1_p & b1c6b7 | !hlock1_p & b1c6b8;
assign ad45b5 = hbusreq4 & ad45b1 | !hbusreq4 & ad45b4;
assign b058a0 = stateG2_p & v845542 | !stateG2_p & !v845582;
assign ad4f07 = hgrant4_p & adea98 | !hgrant4_p & ad4e98;
assign d358e8 = decide_p & v845556 | !decide_p & v84556c;
assign cc36d8 = hmaster0_p & cc36be | !hmaster0_p & v845566;
assign ad476e = hbusreq1 & ad45b6 | !hbusreq1 & ad476b;
assign df5541 = decide_p & df552f | !decide_p & d6ebca;
assign ad4f48 = hbusreq4_p & v845542 | !hbusreq4_p & v84556c;
assign ad4770 = hbusreq1_p & ad476f | !hbusreq1_p & ad45ca;
assign b1c84f = hready_p & b1c82d | !hready_p & b1c84e;
assign v9f77a5 = hbusreq1 & v9f77a3 | !hbusreq1 & v9f77a4;
assign b1c030 = hbusreq4_p & b1c755 | !hbusreq4_p & b1c02f;
assign v9f7d18 = hlock1 & v9f7d12 | !hlock1 & v9f7d17;
assign bd56d8 = hmaster2_p & v845542 | !hmaster2_p & bd56d7;
assign dc5007 = hmaster2_p & dc4feb | !hmaster2_p & dc5006;
assign b058f9 = hlock4 & b058b8 | !hlock4 & b058f8;
assign ade667 = jx2_p & ade653 | !jx2_p & ade666;
assign c3d505 = hgrant1_p & v84554d | !hgrant1_p & c3d504;
assign c3cf2e = hmaster1_p & c3d5ec | !hmaster1_p & c3cf2d;
assign c3cdff = hmaster0_p & c3d306 | !hmaster0_p & c3cdfe;
assign c3ce44 = hbusreq1_p & c3ce43 | !hbusreq1_p & c3d305;
assign d35569 = hmaster1_p & d35568 | !hmaster1_p & d354d3;
assign ad4ee0 = hgrant4_p & ad4eae | !hgrant4_p & v845542;
assign b573e7 = hmaster0_p & v845542 | !hmaster0_p & b573e6;
assign v9f7c97 = stateA1_p & v845542 | !stateA1_p & !v9f7c96;
assign v9ea5df = hmaster1_p & v9ea5de | !hmaster1_p & v9ea583;
assign dc4f66 = hmaster2_p & ade4bf | !hmaster2_p & !v845566;
assign ad4e93 = hbusreq3 & ad4e92 | !hbusreq3 & v845542;
assign b05a18 = hgrant4_p & b058a7 | !hgrant4_p & v9f769d;
assign ad4325 = hgrant1_p & v845542 | !hgrant1_p & ad4324;
assign c3cea4 = hbusreq1 & c3ce9c | !hbusreq1 & c3ce9f;
assign df518d = hbusreq1 & dc501a | !hbusreq1 & !v845542;
assign ad4816 = hbusreq3 & ad4815 | !hbusreq3 & ad4f40;
assign dc5022 = hgrant4_p & adeca0 | !hgrant4_p & !ade563;
assign v9f770f = hmaster1_p & v9f770e | !hmaster1_p & v9f7675;
assign dc5079 = hbusreq1 & dc4fd4 | !hbusreq1 & v84556c;
assign b579bf = hbusreq4 & b579bd | !hbusreq4 & b579be;
assign ad5063 = hready & ad5058 | !hready & ad5062;
assign ad4fdf = hbusreq4_p & ad4fdd | !hbusreq4_p & ad4fde;
assign ad4f5f = hbusreq1_p & ad4f57 | !hbusreq1_p & ad4f5e;
assign ad5028 = hbusreq3 & ad5027 | !hbusreq3 & v845547;
assign c3cea7 = hmaster1_p & c3cea3 | !hmaster1_p & c3cea6;
assign v9f77d8 = hmaster2_p & v9f77c7 | !hmaster2_p & v9f772f;
assign c3d36f = busreq_p & c3d36e | !busreq_p & v845542;
assign d356c4 = hmaster0_p & d356c2 | !hmaster0_p & d356c3;
assign b1c068 = stateG10_4_p & b1c066 | !stateG10_4_p & b1c067;
assign d3558d = hbusreq4_p & d354ce | !hbusreq4_p & !d35aab;
assign ade5bb = hready_p & ade5b9 | !hready_p & ade5ba;
assign b579b7 = stateG2_p & v845542 | !stateG2_p & b579b6;
assign b058a9 = locked_p & b058a6 | !locked_p & !v9ea3e9;
assign ad4688 = hbusreq2 & ad4560 | !hbusreq2 & ad456b;
assign c3d73b = hmaster0_p & c3d685 | !hmaster0_p & c3d6b5;
assign v9f7789 = hlock4 & v9f772c | !hlock4 & v9f7788;
assign df50cd = hbusreq1_p & df50cc | !hbusreq1_p & !v845542;
assign dc4ffd = hbusreq1 & c3d66d | !hbusreq1 & !v845542;
assign df5188 = hbusreq1 & c3d66d | !hbusreq1 & v845542;
assign b1c4af = hmaster1_p & v845542 | !hmaster1_p & b1c4ae;
assign v9e9f9c = hbusreq3 & v9e9f99 | !hbusreq3 & v9e9f9b;
assign v9ea5f3 = hmaster0_p & v9f20a1 | !hmaster0_p & v9ea4a7;
assign v9f7d57 = stateA1_p & v845542 | !stateA1_p & !v9ea3e5;
assign v9f76a1 = hgrant4_p & v9f7d62 | !hgrant4_p & v9f7663;
assign v9e9fe5 = hgrant3_p & v9e9fdc | !hgrant3_p & v9e9fe4;
assign v8cc4f7 = hready_p & v8cc4e0 | !hready_p & v8cc4f6;
assign d354d4 = hmaster1_p & d354b8 | !hmaster1_p & d354d3;
assign d35416 = hlock3_p & d35bff | !hlock3_p & !d35415;
assign v845580 = stateG3_1_p & v845542 | !stateG3_1_p & !v845542;
assign d357ee = hmaster0_p & d357ea | !hmaster0_p & d357ed;
assign v8cc81e = hmaster1_p & v8cc81d | !hmaster1_p & v845542;
assign c3d677 = hbusreq1_p & c3d671 | !hbusreq1_p & c3d676;
assign dc5314 = hlock3_p & dc5311 | !hlock3_p & !v845542;
assign ad446c = hmaster0_p & ad481c | !hmaster0_p & v845547;
assign d35434 = hlock4_p & v845542 | !hlock4_p & !d3591a;
assign ad4edf = hmaster2_p & ad4ed6 | !hmaster2_p & ad4ede;
assign b1c75c = hbusreq0 & b1c75b | !hbusreq0 & !v845542;
assign b1c848 = hbusreq0 & b1c845 | !hbusreq0 & b1c847;
assign c3cee2 = hbusreq0 & c3cee1 | !hbusreq0 & v845542;
assign d357ac = hmaster0_p & d35799 | !hmaster0_p & d35795;
assign c3d6b6 = hbusreq1_p & c3d6b3 | !hbusreq1_p & !c3d6b5;
assign b1c708 = hready_p & b1c706 | !hready_p & b1c707;
assign ad4f4d = hbusreq3 & ad4f4c | !hbusreq3 & v845542;
assign b1c79e = hgrant4_p & b1c71a | !hgrant4_p & !b1c79d;
assign ad4e40 = decide_p & ad4e20 | !decide_p & ad4e24;
assign d35a45 = hgrant4_p & v845542 | !hgrant4_p & !d35a43;
assign v845566 = hmastlock_p & v845542 | !hmastlock_p & !v845542;
assign ad484b = hbusreq2 & ad484a | !hbusreq2 & v845542;
assign bd58ad = hmaster2_p & bd58a9 | !hmaster2_p & dc5011;
assign v9ea3e4 = start_p & v845542 | !start_p & !v845582;
assign v9f7831 = hbusreq0 & v9f782e | !hbusreq0 & v9f7830;
assign bd5936 = hbusreq2 & bd5931 | !hbusreq2 & bd5935;
assign b1c496 = hbusreq4_p & b1c495 | !hbusreq4_p & !v84554a;
assign ade58e = hgrant4_p & v84556c | !hgrant4_p & !ade58d;
assign c3d514 = hmaster2_p & c3d50f | !hmaster2_p & v845542;
assign b1c850 = hbusreq0 & b1cfb7 | !hbusreq0 & b1cfcc;
assign ad4fe6 = hlock0_p & v845542 | !hlock0_p & ad4fe5;
assign d35a08 = hbusreq4_p & d35a06 | !hbusreq4_p & d35a07;
assign b058c3 = hbusreq3 & b058c1 | !hbusreq3 & b058c2;
assign v8cc5ab = hready & v8cc5aa | !hready & v8cc494;
assign b1c610 = decide_p & b1c5fc | !decide_p & b1d013;
assign ad438a = hbusreq0 & ad4389 | !hbusreq0 & v845542;
assign b57a7e = hbusreq3 & b57a7c | !hbusreq3 & b57a7d;
assign dc4f9a = hbusreq3 & ade4bf | !hbusreq3 & v845542;
assign bd57ca = hgrant1_p & bd57c9 | !hgrant1_p & bd57c7;
assign b05a88 = hmaster0_p & b058c7 | !hmaster0_p & b059fb;
assign ad4721 = hmaster0_p & ad4706 | !hmaster0_p & ad4720;
assign b059d4 = hgrant4_p & b058a7 | !hgrant4_p & !b05953;
assign bd5804 = hgrant0_p & v84556c | !hgrant0_p & bd57fb;
assign b1c859 = hbusreq1_p & b1cfb7 | !hbusreq1_p & b1c858;
assign d35a03 = hlock0_p & v845542 | !hlock0_p & d35a02;
assign bd57c4 = hburst0 & bd57bf | !hburst0 & bd57c3;
assign ad4f1c = hmaster0_p & ad4f19 | !hmaster0_p & ad4f1b;
assign c3d2d7 = hbusreq3 & c3d2d6 | !hbusreq3 & v845542;
assign df5530 = decide_p & df552f | !decide_p & v845542;
assign v8cc600 = hready_p & v8cc4e0 | !hready_p & v8cc5ff;
assign ad416f = decide_p & ad4165 | !decide_p & ad416e;
assign ad458c = hbusreq1_p & ad4586 | !hbusreq1_p & ad458b;
assign b1c82e = hmaster0_p & v845542 | !hmaster0_p & b1cf2c;
assign v9f7cb5 = hmaster2_p & v9f7c9c | !hmaster2_p & !v9f7cb4;
assign ad4273 = hbusreq3 & ad4272 | !hbusreq3 & v845542;
assign ad45af = hlock4_p & dc4f78 | !hlock4_p & ad45ae;
assign d35565 = hbusreq2 & d35bf2 | !hbusreq2 & d35be8;
assign c3cf19 = hbusreq0 & c3cede | !hbusreq0 & v845564;
assign ad4766 = hmaster2_p & v845542 | !hmaster2_p & ad4765;
assign cc3703 = hgrant1_p & df54f3 | !hgrant1_p & cc3702;
assign b1c717 = hmaster2_p & b1c714 | !hmaster2_p & !b1c716;
assign ad4167 = hbusreq2 & ad4fbf | !hbusreq2 & v845542;
assign b058f0 = hlock1 & b058ea | !hlock1 & b058ef;
assign b1c71d = hbusreq0 & b1c714 | !hbusreq0 & v845542;
assign ad4ec0 = hmaster2_p & ad4e7c | !hmaster2_p & ad4ebf;
assign v9f7d8b = hgrant4_p & v9f7cb6 | !hgrant4_p & v9f7d8a;
assign v9ea5b8 = hbusreq2_p & v9ea5ac | !hbusreq2_p & v9ea5b7;
assign v9f7899 = hmaster0_p & v9f7898 | !hmaster0_p & !v9f77f3;
assign v9e9f88 = hbusreq2 & v9e9f86 | !hbusreq2 & v9e9f87;
assign b059e9 = hbusreq0 & b059de | !hbusreq0 & b059e8;
assign c3d376 = hgrant1_p & v845564 | !hgrant1_p & c3d375;
assign ad425e = decide_p & ad40f0 | !decide_p & ad41ab;
assign b57ab2 = hbusreq3 & b57a85 | !hbusreq3 & b57942;
assign bd5824 = hgrant1_p & bd57f3 | !hgrant1_p & bd5823;
assign d3562b = hmaster1_p & d35622 | !hmaster1_p & d3562a;
assign d35695 = hmaster1_p & d35aae | !hmaster1_p & d35694;
assign ad4fe1 = hgrant4_p & ad4fce | !hgrant4_p & !v84556c;
assign v9f7de9 = hbusreq0 & v9f7dd6 | !hbusreq0 & v9f7de8;
assign ade662 = jx1_p & ade661 | !jx1_p & adeab8;
assign df5157 = hbusreq1_p & df5156 | !hbusreq1_p & v845542;
assign dc5021 = hgrant4_p & adeca1 | !hgrant4_p & ade563;
assign b058de = hbusreq3 & b058dc | !hbusreq3 & b058dd;
assign ad4df6 = hmaster0_p & v845555 | !hmaster0_p & ad4df5;
assign ad47f6 = hgrant2_p & ad47f4 | !hgrant2_p & !ad47f5;
assign v9f7e08 = hbusreq1_p & v9f7e07 | !hbusreq1_p & v9f7d12;
assign bd591b = hgrant2_p & bd591a | !hgrant2_p & !v845542;
assign ad427a = hmaster0_p & ad4276 | !hmaster0_p & ad4279;
assign b8f6e5 = hgrant2_p & v845542 | !hgrant2_p & !b8f6e4;
assign d35a6d = hmaster1_p & d35a4c | !hmaster1_p & d35a6c;
assign b1c7b5 = hbusreq0 & b1c7b4 | !hbusreq0 & v845542;
assign ad4724 = hbusreq2_p & ad471d | !hbusreq2_p & ad4723;
assign c3ce99 = hmaster1_p & c3d35b | !hmaster1_p & c3ce98;
assign ad45e7 = hlock4_p & ad4daf | !hlock4_p & !ad45e6;
assign ad43f7 = hbusreq4_p & ad43f6 | !hbusreq4_p & v845542;
assign ad46b0 = hbusreq1 & ad4560 | !hbusreq1 & ad456b;
assign b1c0a6 = hbusreq1_p & b1cfd0 | !hbusreq1_p & b1c85f;
assign ade571 = hburst0 & v845542 | !hburst0 & ade570;
assign v9f7882 = hlock0_p & v9f77be | !hlock0_p & v9f7881;
assign b1c7b3 = hlock0_p & bd5838 | !hlock0_p & v845542;
assign c5c8e1 = hlock3_p & c5c8a4 | !hlock3_p & c5c8e0;
assign ad3cfc = hbusreq1 & ad3cf1 | !hbusreq1 & ad3cfb;
assign d3578f = hmaster2_p & d3578a | !hmaster2_p & d3578e;
assign b579d6 = hgrant4_p & b579ba | !hgrant4_p & v845542;
assign dc4f72 = hbusreq1_p & dc4f6e | !hbusreq1_p & dc4f71;
assign v8cc489 = hgrant1_p & v8ccbd8 | !hgrant1_p & v8cc474;
assign v9ea431 = hmaster2_p & v9ea42f | !hmaster2_p & v9ea430;
assign b05a8d = decide_p & b05a84 | !decide_p & b05a8c;
assign v8ccb66 = hburst1_p & bbbcd8 | !hburst1_p & !bb9c5a;
assign v8cc5a9 = hbusreq0 & v8cc5a8 | !hbusreq0 & v8cc494;
assign c3cdfa = hmaster0_p & c3d5ed | !hmaster0_p & c3d5cf;
assign d35714 = hmaster1_p & d35710 | !hmaster1_p & d35713;
assign b058d4 = hlock0_p & v9ea3e9 | !hlock0_p & b058d3;
assign v9f7753 = hbusreq0 & v9f7750 | !hbusreq0 & v9f7752;
assign dc53bf = hbusreq1_p & dc5394 | !hbusreq1_p & dc53a3;
assign c3d50b = hmaster0_p & c3d509 | !hmaster0_p & c3d50a;
assign ad4fb1 = hbusreq3 & ad4fb0 | !hbusreq3 & v845542;
assign ad45ef = hlock4_p & ad4daf | !hlock4_p & !v845542;
assign ad43e0 = hbusreq1_p & ad43df | !hbusreq1_p & ad43de;
assign c3d529 = hbusreq4 & c3d528 | !hbusreq4 & !v845542;
assign b573fa = hgrant3_p & b57946 | !hgrant3_p & b573f9;
assign bd5ba1 = hgrant3_p & bd5b7e | !hgrant3_p & !bd5ba0;
assign v9f7890 = hbusreq3 & v9f788e | !hbusreq3 & v9f788f;
assign b1c73d = hmaster2_p & b1c731 | !hmaster2_p & !b1c73c;
assign b058b1 = hbusreq1 & b058af | !hbusreq1 & b058b0;
assign ba7c7d = hready_p & ba7c7c | !hready_p & ba7c70;
assign v9f7d76 = stateG10_4_p & v9f7d72 | !stateG10_4_p & v9f7d74;
assign v9ea57b = hmaster0_p & v9ea571 | !hmaster0_p & v9ea575;
assign v9ea596 = hlock3 & v9ea595 | !hlock3 & v9ea593;
assign d356cb = hlock1_p & d35a21 | !hlock1_p & v845542;
assign v9f7dd5 = hbusreq4_p & v9f7dd3 | !hbusreq4_p & v9f7dd4;
assign df5116 = hbusreq1 & dc5394 | !hbusreq1 & dc539f;
assign b058cc = hlock2 & b058c9 | !hlock2 & b058cb;
assign ad4781 = hmaster0_p & ad4770 | !hmaster0_p & ad477d;
assign c3d6cf = hbusreq4_p & c3d6cc | !hbusreq4_p & !c3d6ce;
assign b578f8 = stateG2_p & v845542 | !stateG2_p & b578f7;
assign df507e = hready_p & v845542 | !hready_p & df507d;
assign c3d4f5 = hbusreq0 & v845542 | !hbusreq0 & c3d4f4;
assign c3d6c4 = hgrant4_p & c3d6b4 | !hgrant4_p & c3d6b8;
assign v9f7866 = hbusreq1_p & v9f775a | !hbusreq1_p & v9f785e;
assign bd579b = hmaster2_p & bd5786 | !hmaster2_p & !ade4e6;
assign d3598d = hbusreq2 & d3598c | !hbusreq2 & v845542;
assign ade653 = jx0_p & adeab9 | !jx0_p & ade652;
assign b05977 = hbusreq1_p & b05976 | !hbusreq1_p & b0590e;
assign ad4ed0 = hbusreq1 & ad4ecf | !hbusreq1 & v845542;
assign c3d5bc = hbusreq0 & c3d5b6 | !hbusreq0 & c3d5bb;
assign bd57d0 = hmaster2_p & bd57c4 | !hmaster2_p & v845542;
assign dc53c5 = decide_p & dc53c4 | !decide_p & !v845542;
assign v9f7822 = hbusreq4 & v9f7820 | !hbusreq4 & v9f7821;
assign v9f7851 = hgrant2_p & v9f7819 | !hgrant2_p & v9f7850;
assign b1c5e5 = hlock0_p & b1c5e4 | !hlock0_p & !v845542;
assign ad4320 = hbusreq1_p & ad431f | !hbusreq1_p & v845542;
assign ad46bd = hbusreq4_p & ad46bc | !hbusreq4_p & v845542;
assign d35a3a = stateG2_p & v845542 | !stateG2_p & adea96;
assign d35a4e = hburst0 & v8cc793 | !hburst0 & d35a4d;
assign ad4466 = hbusreq4 & ad445f | !hbusreq4 & ad4465;
assign ad4fef = hmaster1_p & ad4fc5 | !hmaster1_p & ad4fee;
assign ad4ff9 = hgrant2_p & ad4ff3 | !hgrant2_p & ad4ff8;
assign d35a7a = hlock3_p & d35a36 | !hlock3_p & d35a79;
assign d35bfc = hbusreq3 & d35bf2 | !hbusreq3 & d35be8;
assign c3d586 = decide_p & c3d585 | !decide_p & c3d50d;
assign c3ceac = hmaster2_p & d35a98 | !hmaster2_p & v845542;
assign ac1489 = hbusreq4_p & ac1459 | !hbusreq4_p & ac1488;
assign v9f7d24 = hlock0 & v9f7d23 | !hlock0 & !v9f7c9f;
assign c3d6d3 = hmaster1_p & c3d6b2 | !hmaster1_p & c3d6d2;
assign v9f789c = hbusreq2_p & v9f787e | !hbusreq2_p & v9f789b;
assign df54e3 = hbusreq1 & dc5394 | !hbusreq1 & df54e2;
assign ad45a5 = hmaster0_p & ad45a0 | !hmaster0_p & ad45a4;
assign ad4710 = hgrant1_p & ad470e | !hgrant1_p & ad470f;
assign ad3d0a = hbusreq4 & ad3d04 | !hbusreq4 & ad3d09;
assign bd5781 = hmastlock_p & ade4bc | !hmastlock_p & c3d668;
assign ad40ef = hlock2_p & ad40ed | !hlock2_p & !ad40ee;
assign ad4768 = hbusreq4_p & ad4767 | !hbusreq4_p & !v845542;
assign ad4dba = hmaster1_p & ad4d9f | !hmaster1_p & ad4db9;
assign b1c5d8 = hbusreq0 & b1c5d7 | !hbusreq0 & df54d6;
assign b1caf4 = hbusreq4_p & d35918 | !hbusreq4_p & b1cf29;
assign ad4e4b = hmaster2_p & v845542 | !hmaster2_p & ad4e47;
assign v91784a = hmaster0_p & v845542 | !hmaster0_p & v845564;
assign v8cc7e7 = hbusreq1_p & v8cc79e | !hbusreq1_p & v8cc7e6;
assign ad3cdd = hbusreq0_p & ad502f | !hbusreq0_p & !v845542;
assign ad46e1 = hbusreq4 & ad46d4 | !hbusreq4 & ad46e0;
assign b1c02e = hbusreq0_p & bd57c4 | !hbusreq0_p & v845542;
assign ad4fb5 = hbusreq3 & ad4fb4 | !hbusreq3 & v845542;
assign d35744 = hmaster0_p & d35743 | !hmaster0_p & d3570f;
assign ad45ff = hbusreq3 & ad45c6 | !hbusreq3 & ad45c9;
assign b1c808 = hbusreq1_p & b1c73e | !hbusreq1_p & b1c807;
assign v9f7dbc = hbusreq1_p & v9f7d97 | !hbusreq1_p & v9f7dbb;
assign c5c8fb = hbusreq4_p & c5c8fa | !hbusreq4_p & !v845542;
assign c3d396 = hmaster0_p & c3d306 | !hmaster0_p & c3d395;
assign v8cc508 = hmaster0_p & v8cc489 | !hmaster0_p & v8cc4ad;
assign d359f7 = hlock0_p & v845542 | !hlock0_p & d359f6;
assign v9e9e6a = hmaster0_p & v9e9e69 | !hmaster0_p & v9ea603;
assign c3d57c = hmaster2_p & c3d57b | !hmaster2_p & v845576;
assign b05a96 = hgrant2_p & b05a94 | !hgrant2_p & b05a95;
assign dc5038 = hgrant4_p & dc5037 | !hgrant4_p & adec89;
assign b059ba = hlock3 & b05964 | !hlock3 & b059b9;
assign c3ce9d = hgrant1_p & c3d2d6 | !hgrant1_p & c3ce9c;
assign d35657 = hmaster2_p & d35a5b | !hmaster2_p & d35656;
assign ad4429 = hbusreq0 & ad4103 | !hbusreq0 & v845542;
assign v9f77c4 = hgrant0_p & v9f772b | !hgrant0_p & v9f77c3;
assign ade4dd = hbusreq1_p & ade4d2 | !hbusreq1_p & ade4dc;
assign c3ce8b = hbusreq3_p & c3ce74 | !hbusreq3_p & c3ce8a;
assign c3d598 = hbusreq2 & c3d597 | !hbusreq2 & v84554d;
assign ad46e8 = hbusreq2 & ad4586 | !hbusreq2 & !v845547;
assign df54d8 = hlock1_p & df54d7 | !hlock1_p & v845542;
assign d35422 = hlock4_p & d358ef | !hlock4_p & !dc5318;
assign v9f7646 = hready & v9f7645 | !hready & v9f7e3f;
assign c3ce86 = hbusreq2_p & c3ce50 | !hbusreq2_p & c3ce85;
assign ad429e = hready & ad4ddd | !hready & !ad45ae;
assign ad46ef = hlock2_p & ad46e6 | !hlock2_p & !ad46ee;
assign d354a4 = hbusreq4_p & d354a3 | !hbusreq4_p & v845542;
assign d356ce = hmaster1_p & d356cd | !hmaster1_p & d356c9;
assign ad4f18 = hgrant2_p & ad4e62 | !hgrant2_p & ad4f17;
assign ad4392 = hbusreq0 & ad4380 | !hbusreq0 & v845542;
assign v9ea4c0 = hmaster1_p & v9ea4bf | !hmaster1_p & v9ea4bd;
assign c3d4f1 = hmaster2_p & c3d4f0 | !hmaster2_p & v845576;
assign c5c8a5 = hmaster0_p & c5c898 | !hmaster0_p & c5c897;
assign v9e9fc2 = hmaster0_p & v9e9fae | !hmaster0_p & v9e9f63;
assign ad3d5a = decide_p & ad4409 | !decide_p & ad3d59;
assign v9f7833 = hbusreq4 & v9f7831 | !hbusreq4 & v9f7832;
assign bd584e = hgrant4_p & v84556c | !hgrant4_p & bd5842;
assign ade4b0 = hmaster1_p & adec9f | !hmaster1_p & ade4af;
assign ad4fca = locked_p & ad4fc9 | !locked_p & v845542;
assign ad4d94 = hbusreq3 & ad4d93 | !hbusreq3 & v845542;
assign b1c723 = hbusreq1_p & b1c71c | !hbusreq1_p & b1c722;
assign bd5822 = hbusreq0 & bd5818 | !hbusreq0 & bd5821;
assign d354ef = hmaster0_p & d354ee | !hmaster0_p & d35c05;
assign v9f7e28 = hgrant1_p & v9f7cb7 | !hgrant1_p & v9f7e1f;
assign ade4e5 = hburst1 & v845542 | !hburst1 & ade4e4;
assign v9e9fd8 = hgrant3_p & v9e9fcf | !hgrant3_p & v9e9fd7;
assign ade57e = hgrant1_p & ade576 | !hgrant1_p & !ade57d;
assign ad473d = hready & ad4739 | !hready & !ad473c;
assign v8cc473 = hgrant4_p & v845542 | !hgrant4_p & v8d2b2e;
assign ad456c = hbusreq3 & ad4560 | !hbusreq3 & ad456b;
assign v9f77ff = hmaster0_p & v9f77d4 | !hmaster0_p & v9f77fe;
assign c3d523 = hbusreq4_p & c3d2b0 | !hbusreq4_p & !v845542;
assign v9ea4a0 = hready_p & v9ea436 | !hready_p & v9ea49f;
assign ad4f91 = hgrant4_p & v845542 | !hgrant4_p & ad4f80;
assign dc5051 = hgrant4_p & dc5050 | !hgrant4_p & adec89;
assign bd57f9 = stateA1_p & v845578 | !stateA1_p & !bd57f8;
assign v8ccbf6 = hgrant1_p & v845542 | !hgrant1_p & v8ccbf4;
assign v9ea4a3 = hmaster1_p & v9ea4a2 | !hmaster1_p & v845542;
assign b1d01a = hbusreq1_p & v845542 | !hbusreq1_p & d35a9c;
assign adea86 = stateG2_p & v845542 | !stateG2_p & !adea85;
assign v9f7701 = hbusreq2 & v9f76ff | !hbusreq2 & v9f7700;
assign df5169 = hbusreq2 & df5166 | !hbusreq2 & df5168;
assign b57b59 = hgrant3_p & b57af7 | !hgrant3_p & b57b58;
assign df51a5 = hbusreq3 & df5189 | !hbusreq3 & !v84554c;
assign ad4ec3 = hbusreq0 & ad4e83 | !hbusreq0 & ad4ea0;
assign b1c6bb = hgrant1_p & v845542 | !hgrant1_p & b1c6ba;
assign b57a1a = hbusreq0_p & b578f9 | !hbusreq0_p & v845542;
assign v8cc16a = hbusreq3_p & v8cc169 | !hbusreq3_p & v8cc50e;
assign v9ea444 = hbusreq4_p & v9ea442 | !hbusreq4_p & v9ea443;
assign ad5014 = stateA1_p & v9c81a4 | !stateA1_p & !adea96;
assign b058d0 = hlock0_p & b058b6 | !hlock0_p & b058cf;
assign b57401 = hready_p & b57a12 | !hready_p & b57400;
assign df5162 = hbusreq1_p & df5161 | !hbusreq1_p & v845542;
assign v9f7cd1 = hbusreq1_p & v9f7cb7 | !hbusreq1_p & v9f7cc8;
assign c3cf22 = hmaster1_p & c3cf1e | !hmaster1_p & c3cf21;
assign v9e9ee2 = decide_p & v9e9e75 | !decide_p & v9e9ee1;
assign bd56d0 = hburst1 & bd5b6a | !hburst1 & bd56cf;
assign ad44b5 = hbusreq0 & ad44b4 | !hbusreq0 & v845542;
assign b1c5f6 = decide_p & b1c5dd | !decide_p & b1d013;
assign ad4434 = hbusreq1 & ad4385 | !hbusreq1 & ad438b;
assign d35732 = hmaster0_p & d3572f | !hmaster0_p & !d35731;
assign bd5842 = hlock0_p & bd5840 | !hlock0_p & !bd5841;
assign c5c93c = hmaster0_p & c5c932 | !hmaster0_p & c5c93b;
assign ad4382 = hlock0_p & dc52fa | !hlock0_p & ad4381;
assign ad43f5 = hbusreq0 & ad43f4 | !hbusreq0 & v845542;
assign b1c755 = hbusreq0_p & b1c754 | !hbusreq0_p & !v845542;
assign ad4f36 = hmastlock_p & ad4f35 | !hmastlock_p & v845542;
assign d35abd = hbusreq3_p & d35a93 | !hbusreq3_p & !d35abc;
assign ad448c = hbusreq0_p & ad4fce | !hbusreq0_p & !v845542;
assign bd5767 = hbusreq2_p & bd5766 | !hbusreq2_p & v845542;
assign c5c973 = hgrant1_p & c5c8e9 | !hgrant1_p & c5c972;
assign ad4e74 = hmaster2_p & ad4e73 | !hmaster2_p & v845542;
assign ad4395 = hbusreq3 & ad4394 | !hbusreq3 & v845542;
assign v8ccb82 = hmaster1_p & v8d29fa | !hmaster1_p & v8ccb81;
assign ad46aa = hbusreq4_p & ad46a9 | !hbusreq4_p & v845542;
assign b1caeb = hlock4_p & b1cf26 | !hlock4_p & d3591a;
assign bd58b2 = hmaster2_p & bd58a9 | !hmaster2_p & v845542;
assign dc53ca = hbusreq3_p & dc53c9 | !hbusreq3_p & !dc5088;
assign ad4456 = hgrant4_p & ad437d | !hgrant4_p & v845542;
assign ad471f = hmaster1_p & ad471e | !hmaster1_p & ad45a5;
assign b57907 = hmaster0_p & b578fa | !hmaster0_p & b578f9;
assign df51dc = hready_p & df51da | !hready_p & df51db;
assign b57acb = hmaster0_p & b57aca | !hmaster0_p & b578f9;
assign v9ea56b = hmaster0_p & v9ea568 | !hmaster0_p & v9ea56a;
assign v8cc4fe = hbusreq1_p & v8ccbe3 | !hbusreq1_p & v8cc4fd;
assign df51c9 = hbusreq2_p & df51bf | !hbusreq2_p & df51c8;
assign b8f74d = hready_p & b8f74c | !hready_p & v845562;
assign v9f7e1b = hbusreq4_p & v9f7e19 | !hbusreq4_p & v9f7e1a;
assign bd5e20 = hmaster0_p & v845542 | !hmaster0_p & bd5e1f;
assign d357c0 = hbusreq1_p & d357bf | !hbusreq1_p & v84554a;
assign bd58ba = hgrant4_p & bd575d | !hgrant4_p & v84556c;
assign ade4eb = hbusreq0 & ade4e3 | !hbusreq0 & ade4ea;
assign b1c6df = decide_p & b1c6de | !decide_p & v845542;
assign v9f78a1 = hbusreq2_p & v9f789e | !hbusreq2_p & v9f78a0;
assign b57ab9 = decide_p & b57a21 | !decide_p & b57a8c;
assign dc53a9 = decide_p & dc53a8 | !decide_p & !v845542;
assign dc5058 = hbusreq4_p & dc5055 | !hbusreq4_p & dc5057;
assign ad4605 = hbusreq2_p & ad4604 | !hbusreq2_p & ad4603;
assign bd592c = decide_p & bd592b | !decide_p & v845542;
assign dc5031 = hbusreq1 & dc4fd9 | !hbusreq1 & v84556c;
assign v9f76eb = locked_p & v9f76ea | !locked_p & !v9f7ca4;
assign bd590b = hmaster0_p & v845542 | !hmaster0_p & bd590a;
assign v9041a4 = hmaster2_p & v845542 | !hmaster2_p & !v845558;
assign d359bc = hmastlock_p & d359b9 | !hmastlock_p & !v845542;
assign bd57ef = decide_p & bd57ee | !decide_p & v845542;
assign ad410d = hbusreq1 & ad4807 | !hbusreq1 & ad4809;
assign ad4747 = hbusreq0 & ad4743 | !hbusreq0 & ad4746;
assign b1c752 = hmastlock_p & b1c751 | !hmastlock_p & !b1c74e;
assign df51ad = hbusreq3 & df51ac | !hbusreq3 & !v84554c;
assign ac1490 = hgrant2_p & cc36d3 | !hgrant2_p & ac148f;
assign b1c759 = hbusreq0_p & ade4cc | !hbusreq0_p & !v845542;
assign v8a9702 = hmaster0_p & v845564 | !hmaster0_p & v845542;
assign c3d758 = hmaster0_p & c3d714 | !hmaster0_p & c3d70a;
assign c3d332 = hmaster1_p & c3d317 | !hmaster1_p & c3d331;
assign c3ce03 = hbusreq2 & c3d35d | !hbusreq2 & c3d306;
assign v8cc634 = hready_p & v8cc4e0 | !hready_p & v8cc633;
assign b1cae9 = hbusreq4_p & b1cf24 | !hbusreq4_p & b1cf29;
assign b1c866 = hgrant2_p & v845542 | !hgrant2_p & b1d00e;
assign d35a24 = hbusreq2 & d359e9 | !hbusreq2 & v845542;
assign c3d307 = hbusreq3 & c3d302 | !hbusreq3 & c3d306;
assign v9f773b = hmaster1_p & v9f772d | !hmaster1_p & v9f7736;
assign df54f6 = hmaster2_p & v84556c | !hmaster2_p & !dc5300;
assign v9ea41c = hgrant0_p & v9f21c5 | !hgrant0_p & v845542;
assign ade4e0 = hbusreq0_p & ade4df | !hbusreq0_p & !ade4d4;
assign ad4741 = hgrant4_p & v845542 | !hgrant4_p & ad5041;
assign d35022 = decide_p & d35021 | !decide_p & v84556c;
assign ad4fcd = hmastlock_p & ad4fcc | !hmastlock_p & !v845542;
assign d35a52 = hlock1_p & d35a51 | !hlock1_p & !v845542;
assign ad47fe = hmaster1_p & ad47fd | !hmaster1_p & ad45a5;
assign d354e3 = hbusreq1 & d35c08 | !hbusreq1 & !v84555a;
assign v9f7874 = decide_p & v9f7873 | !decide_p & v9f77b8;
assign v9f7757 = hbusreq1 & v9f7755 | !hbusreq1 & v9f7756;
assign v9f7845 = hgrant1_p & v9f77af | !hgrant1_p & !v9f7844;
assign ad505e = hlock0_p & v845542 | !hlock0_p & ad505d;
assign d354d9 = hbusreq2 & d35c09 | !hbusreq2 & !v84555a;
assign b0599e = hlock2 & b0599b | !hlock2 & b0599d;
assign v9f7e10 = hgrant2_p & v9f7e03 | !hgrant2_p & v9f7e0f;
assign dc539e = hmastlock_p & dc539d | !hmastlock_p & v845542;
assign ad42c4 = hmaster0_p & ad42a6 | !hmaster0_p & ad42c3;
assign b57942 = hmaster2_p & v845542 | !hmaster2_p & b57941;
assign ade4e1 = hlock0_p & ade4c5 | !hlock0_p & ade4e0;
assign c3ced0 = hready & c3cecf | !hready & c3d300;
assign v9e9e76 = hbusreq1_p & v9ea404 | !hbusreq1_p & v9ea4bc;
assign b57435 = hbusreq2_p & b5742d | !hbusreq2_p & b57434;
assign d3574c = hbusreq2 & d35730 | !hbusreq2 & d35aa4;
assign v8cc626 = hbusreq2_p & v8cc625 | !hbusreq2_p & v8cc50a;
assign v9f7d2c = hbusreq3 & v9f7d2a | !hbusreq3 & !v9f7d2b;
assign d357a1 = hlock4_p & d357a0 | !hlock4_p & v84554a;
assign b05913 = hmaster0_p & b05907 | !hmaster0_p & b05912;
assign bd58c0 = stateG10_4_p & bd58bd | !stateG10_4_p & !bd58bf;
assign v9f7d95 = hready & v9f7d94 | !hready & v9f7d90;
assign c3ce15 = hbusreq2 & c3d2d6 | !hbusreq2 & v845542;
assign v9e9f7b = hlock4 & v9e9f79 | !hlock4 & v9e9f7a;
assign d35438 = hmaster0_p & d35430 | !hmaster0_p & d35437;
assign ad4717 = hmaster2_p & v845542 | !hmaster2_p & ad4716;
assign bd5746 = hmaster2_p & v84556c | !hmaster2_p & !bd5744;
assign b1c07d = hgrant4_p & b1c7b3 | !hgrant4_p & b1c066;
assign b1c701 = hready_p & b1c6fe | !hready_p & b1c700;
assign v9f76c3 = hbusreq0_p & v9f7d3a | !hbusreq0_p & v9ea3e6;
assign cc36bd = locked_p & v845542 | !locked_p & !v845566;
assign d3559d = hmaster1_p & d35523 | !hmaster1_p & d3559c;
assign ad440d = hbusreq0 & ad440c | !hbusreq0 & v845542;
assign v9ea4c4 = hmaster0_p & v9ea4b7 | !hmaster0_p & v9ea3fa;
assign bd58ee = hbusreq3 & bd579e | !hbusreq3 & bd579f;
assign d3575f = hbusreq2_p & d35aa9 | !hbusreq2_p & d35aa7;
assign b05934 = hbusreq2_p & b05931 | !hbusreq2_p & b05933;
assign ade65c = hmaster1_p & adea95 | !hmaster1_p & ade65b;
assign v9ea60c = hbusreq3 & v9ea485 | !hbusreq3 & v9ea60b;
assign b1c57c = hmaster2_p & d35a9c | !hmaster2_p & b1c57b;
assign v9e9fc9 = hbusreq2_p & v9e9fc4 | !hbusreq2_p & v9e9fc8;
assign b1cfc5 = hlock0_p & b1cfc4 | !hlock0_p & !v845542;
assign b059a7 = hmaster0_p & b05901 | !hmaster0_p & b058e8;
assign ad4599 = hmaster2_p & adec93 | !hmaster2_p & ad4598;
assign v9f7d9b = hgrant1_p & v9f7d9a | !hgrant1_p & v9f7d90;
assign cc36bf = hmaster0_p & v845566 | !hmaster0_p & cc36be;
assign b058ab = hlock0 & b058aa | !hlock0 & b058a8;
assign bbb31e = hburst1_p & v845568 | !hburst1_p & v845542;
assign b058c9 = hbusreq1_p & b058b8 | !hbusreq1_p & b058c7;
assign ad4166 = hbusreq2 & ad4fc3 | !hbusreq2 & v845542;
assign bd5793 = hgrant1_p & bd5792 | !hgrant1_p & bd578c;
assign d35c06 = hmaster0_p & d35c04 | !hmaster0_p & d35c05;
assign b57448 = hmaster1_p & b57447 | !hmaster1_p & v845542;
assign b573e1 = hbusreq1 & b579c0 | !hbusreq1 & b57942;
assign c3d380 = hbusreq3 & c3d37f | !hbusreq3 & c3d2de;
assign b5743e = hmaster1_p & b5743d | !hmaster1_p & v845542;
assign ad4ec7 = hbusreq1_p & ad4ea7 | !hbusreq1_p & ad4ec6;
assign v8cc6b7 = jx1_p & v8cc604 | !jx1_p & v8cc6b6;
assign b05a57 = hmaster1_p & b05a56 | !hmaster1_p & b05913;
assign b1cf24 = hlock0_p & adea88 | !hlock0_p & !v845542;
assign ad4eab = hbusreq1 & ad4e49 | !hbusreq1 & ad4e4e;
assign bd5775 = hbusreq3 & c3d686 | !hbusreq3 & !v845542;
assign ad4dc9 = hbusreq1_p & ad4dc8 | !hbusreq1_p & ad4da1;
assign d359ac = hbusreq3 & d359ab | !hbusreq3 & v845542;
assign ad45e9 = hmaster2_p & v845542 | !hmaster2_p & !ad45e8;
assign v8cc603 = hgrant3_p & v8cc600 | !hgrant3_p & v8cc602;
assign v9e9fb6 = hbusreq3 & v9e9fa3 | !hbusreq3 & v9e9f68;
assign v9f7d33 = hlock2 & v9f7d12 | !hlock2 & v9f7d32;
assign ad413f = hlock4_p & ad413e | !hlock4_p & !v845576;
assign ad4e21 = hbusreq3 & v845542 | !hbusreq3 & c3d2d9;
assign ad4e5d = hmaster2_p & ad4e5a | !hmaster2_p & ad4e5c;
assign v8cc78f = hready_p & v8cc507 | !hready_p & v8cc78e;
assign ad4378 = hready_p & ad4376 | !hready_p & ad4377;
assign v9f7d85 = hgrant4_p & v9f7ca4 | !hgrant4_p & v9f7d83;
assign ad4809 = hready & ad4e4b | !hready & ad4808;
assign d356d6 = hmaster2_p & d35909 | !hmaster2_p & !d35617;
assign ad45c5 = hbusreq4 & ad4d92 | !hbusreq4 & v845542;
assign v9f7d6b = hmaster0_p & v9f7cc2 | !hmaster0_p & v9f7cb2;
assign v8cc76e = hmaster1_p & v8cc76c | !hmaster1_p & v845542;
assign v85746e = hmaster1_p & v845558 | !hmaster1_p & v898970;
assign ad4371 = hmaster0_p & df5142 | !hmaster0_p & ad4320;
assign ad4597 = hlock3_p & ad4584 | !hlock3_p & !ad4596;
assign b1cafe = hmaster1_p & v845542 | !hmaster1_p & b1cafd;
assign bd578e = hmastlock_p & bd578d | !hmastlock_p & v845542;
assign c3ce6b = hbusreq1_p & c3ce6a | !hbusreq1_p & c3d2de;
assign v9ea42d = hgrant1_p & v9ea3e1 | !hgrant1_p & v9ea40f;
assign bd5855 = hbusreq1_p & bd5823 | !hbusreq1_p & bd5854;
assign v9ea418 = hgrant4_p & v9f21c5 | !hgrant4_p & v845542;
assign bd5758 = hmaster2_p & bd5755 | !hmaster2_p & bd5757;
assign cc3701 = hmaster2_p & cc36fb | !hmaster2_p & cc3700;
assign c3d34b = hbusreq0 & c3d33a | !hbusreq0 & c3d34a;
assign c5c99b = decide_p & c5c8e1 | !decide_p & c5c99a;
assign ad45b3 = hbusreq4_p & ad45b2 | !hbusreq4_p & v845542;
assign b57ac4 = hlock1 & b578f9 | !hlock1 & b57ac3;
assign v9ea43e = hbusreq1_p & v9ea43a | !hbusreq1_p & v9ea43d;
assign ad46c3 = hgrant1_p & ad46b6 | !hgrant1_p & ad46c2;
assign cc36e2 = stateG10_4_p & cc36da | !stateG10_4_p & !cc36e1;
assign b0597f = hgrant0_p & b058e7 | !hgrant0_p & v9f7d42;
assign dc5072 = hbusreq3 & dc5071 | !hbusreq3 & v845542;
assign d35ab5 = hbusreq3 & d35aae | !hbusreq3 & d35ab4;
assign ac1485 = hbusreq0_p & ac1458 | !hbusreq0_p & ade562;
assign c3ce56 = hgrant1_p & v84554d | !hgrant1_p & c3ce55;
assign c3d6da = hmaster1_p & c3d6d9 | !hmaster1_p & c3d68b;
assign v9f7794 = hlock4 & v9f772d | !hlock4 & v9f7793;
assign ad4e88 = hbusreq0 & ad4e84 | !hbusreq0 & ad4e87;
assign cc36e9 = hmaster0_p & cc36e0 | !hmaster0_p & !cc36e8;
assign b0598b = hgrant0_p & b058a9 | !hgrant0_p & !v9ea3e9;
assign b058d9 = hbusreq4 & b058d7 | !hbusreq4 & b058d8;
assign b57534 = hgrant3_p & b57946 | !hgrant3_p & b57533;
assign v9ea5d3 = hlock3 & v9ea5cb | !hlock3 & v9ea5d2;
assign v9ea4d2 = hbusreq4_p & v9ea462 | !hbusreq4_p & v9ea4d1;
assign ba7c65 = hbusreq4_p & v845542 | !hbusreq4_p & !adeaa4;
assign df50dc = hmaster1_p & v845542 | !hmaster1_p & df50db;
assign adec95 = hburst0_p & v845542 | !hburst0_p & adec94;
assign ade5d3 = hbusreq1 & ade4c7 | !hbusreq1 & ade5d0;
assign b05a38 = hmaster0_p & b05920 | !hmaster0_p & b0591d;
assign d35710 = hmaster0_p & d3570e | !hmaster0_p & d3570f;
assign c3d6ac = hlock0_p & c3d6ab | !hlock0_p & !c3d66d;
assign v9f777a = hmaster0_p & v9f774f | !hmaster0_p & v9f7779;
assign v9f76d9 = hmaster1_p & v9f76d8 | !hmaster1_p & v9f7d2f;
assign bd58af = hgrant1_p & df5538 | !hgrant1_p & bd58ae;
assign dc52ff = hburst0 & dc52fd | !hburst0 & dc52fe;
assign v8cc7a1 = hlock2 & v8ccb6b | !hlock2 & v8cc7a0;
assign ad4dc1 = hmaster0_p & ad4d94 | !hmaster0_p & ad4dbc;
assign ade624 = hmaster1_p & ade5db | !hmaster1_p & ade4ec;
assign ad428b = hbusreq3 & ad4f1e | !hbusreq3 & !v845542;
assign ba7c74 = hready_p & ba7c73 | !hready_p & ba7c70;
assign ad4420 = hbusreq2 & ad438f | !hbusreq2 & v845542;
assign ade4c3 = hmastlock_p & v845542 | !hmastlock_p & v84557a;
assign ade555 = hgrant0_p & v84556c | !hgrant0_p & ade550;
assign c3d591 = hready & c3d590 | !hready & v845564;
assign ade5a2 = hbusreq0 & ade594 | !hbusreq0 & ade5a1;
assign v9f7806 = hbusreq3 & v9f7803 | !hbusreq3 & v9f7805;
assign dc4fb8 = hbusreq3 & dc4fb7 | !hbusreq3 & v845542;
assign ad4e62 = hmaster1_p & ad4e51 | !hmaster1_p & ad4e61;
assign c3d682 = hmaster2_p & c3d669 | !hmaster2_p & c3d681;
assign b1c790 = hmaster0_p & b1c78e | !hmaster0_p & b1c78f;
assign v8cc7d5 = hlock2_p & v8cc7d2 | !hlock2_p & v8cc7d3;
assign b1c826 = hmaster0_p & b1c825 | !hmaster0_p & b1c75e;
assign v9f7cdf = hbusreq0 & v9f7cd9 | !hbusreq0 & v9f7cde;
assign v9e9ec4 = hbusreq2 & v9e9ec2 | !hbusreq2 & v9e9ec3;
assign b1c7a1 = hbusreq4_p & b1c79e | !hbusreq4_p & !b1c7a0;
assign v9f773c = hmaster0_p & v9f772d | !hmaster0_p & v9f7730;
assign d3577e = hlock3_p & d3577d | !hlock3_p & v84554a;
assign ad45f0 = hbusreq4_p & ad45ef | !hbusreq4_p & !v845542;
assign b059fc = hmaster0_p & b058c5 | !hmaster0_p & b059fb;
assign v9ea593 = hgrant1_p & v9ea58f | !hgrant1_p & v9ea592;
assign b1c737 = hbusreq3 & b1c733 | !hbusreq3 & !b1c736;
assign cc36d1 = hgrant2_p & v84556c | !hgrant2_p & cc36d0;
assign v9f7710 = hgrant2_p & v9f76d4 | !hgrant2_p & v9f770f;
assign ad4564 = hbusreq4_p & ad4563 | !hbusreq4_p & v845542;
assign b1c5f4 = hbusreq2_p & b1d013 | !hbusreq2_p & b1c866;
assign df552e = hmaster0_p & df54e8 | !hmaster0_p & v845542;
assign c3cedc = jx1_p & c3ce8b | !jx1_p & c3cedb;
assign c3ce75 = hbusreq1_p & c3ce34 | !hbusreq1_p & !v845564;
assign bd5816 = stateG10_4_p & bd57fe | !stateG10_4_p & !bd5815;
assign bd5bae = hbusreq2_p & bd5bad | !hbusreq2_p & !v845542;
assign ad4eea = stateG10_4_p & ad4eb3 | !stateG10_4_p & ad4ebf;
assign b579c4 = hgrant1_p & b579c3 | !hgrant1_p & b579b3;
assign ad4283 = hbusreq3 & ad4281 | !hbusreq3 & !ad4282;
assign ad4e95 = hready & d359ad | !hready & v845542;
assign d3540f = hbusreq3 & d35c0b | !hbusreq3 & v84555a;
assign d35bf8 = hmaster2_p & v845542 | !hmaster2_p & d35be8;
assign ad42e4 = hbusreq2 & ad42e0 | !hbusreq2 & ad42e3;
assign b05908 = hlock0 & b058d5 | !hlock0 & v9f7d42;
assign b574ff = hlock2 & b57942 | !hlock2 & b574fe;
assign d35bf1 = hbusreq4_p & d35bf0 | !hbusreq4_p & v845542;
assign d357bb = hbusreq0 & d357ba | !hbusreq0 & v845542;
assign d35a32 = hbusreq3 & d35a31 | !hbusreq3 & v845542;
assign ad4f84 = hbusreq4_p & ad4f81 | !hbusreq4_p & ad4f83;
assign c3ce4a = hbusreq1 & c3d32a | !hbusreq1 & c3d32e;
assign d35958 = hbusreq0 & d35919 | !hbusreq0 & d35957;
assign b57af7 = hready_p & b57a12 | !hready_p & b57af6;
assign v9e9e9a = hmaster1_p & v9ea580 | !hmaster1_p & v9e9e77;
assign b1c784 = hlock2_p & b1c781 | !hlock2_p & b1c783;
assign bd589e = stateA1_p & bd589b | !stateA1_p & v84557c;
assign b1c718 = hbusreq0 & b1c717 | !hbusreq0 & v845542;
assign dc53b7 = jx0_p & dc5089 | !jx0_p & dc53b6;
assign v9f7717 = hmaster0_p & v9f7d5e | !hmaster0_p & v9f7d5a;
assign d358f0 = hmaster2_p & v845542 | !hmaster2_p & d358ef;
assign bd5733 = hburst0 & bd572f | !hburst0 & adec8e;
assign b1c711 = hlock0_p & bd5735 | !hlock0_p & b1c710;
assign v9f7752 = hlock0 & v9f7751 | !hlock0 & v9f7750;
assign ad3cd5 = hmaster2_p & ad3ccc | !hmaster2_p & ad4482;
assign ad13e2 = hgrant2_p & v84554c | !hgrant2_p & ad13df;
assign d3580a = hbusreq4_p & d357c4 | !hbusreq4_p & d35809;
assign v9f775c = hbusreq0 & v9f7759 | !hbusreq0 & v9f775b;
assign c3d2fe = hmaster2_p & c3d2fd | !hmaster2_p & v845542;
assign ade598 = locked_p & ade597 | !locked_p & v845542;
assign b1c073 = hbusreq0 & b1c072 | !hbusreq0 & b1c85e;
assign d354c6 = hgrant1_p & d354bf | !hgrant1_p & d354c5;
assign ad43c1 = hburst0_p & v9ea411 | !hburst0_p & !ad43c0;
assign ad47ec = hmaster1_p & ad47eb | !hmaster1_p & ad46e4;
assign d354bc = hlock4_p & d359c9 | !hlock4_p & !v845542;
assign v9ea465 = hgrant4_p & v9f20a1 | !hgrant4_p & v9ea457;
assign b05a8f = hmaster1_p & b05a8e | !hmaster1_p & b05943;
assign v8ccb74 = decide_p & v8ccb72 | !decide_p & v8ccb6e;
assign ad459f = hmaster0_p & ad459d | !hmaster0_p & ad459e;
assign bd57e6 = hbusreq2 & bd57e5 | !hbusreq2 & v845542;
assign ad4272 = hbusreq1_p & ad4271 | !hbusreq1_p & v845542;
assign v9f777d = hmaster0_p & v9f7772 | !hmaster0_p & v9f774f;
assign dc504c = stateA1_p & v845542 | !stateA1_p & bbbe36;
assign ad3d32 = hready_p & ad3d27 | !hready_p & ad3d31;
assign d3599a = hlock4_p & d35998 | !hlock4_p & !d35999;
assign ad44a3 = hgrant4_p & ad43a4 | !hgrant4_p & c3cec2;
assign b05a2a = decide_p & b05935 | !decide_p & !b05a29;
assign ad48c7 = hgrant2_p & ad508e | !hgrant2_p & ad48c6;
assign ad3d02 = hbusreq4_p & ad3cff | !hbusreq4_p & ad3d01;
assign ad4e4f = hbusreq3 & ad4e4e | !hbusreq3 & v845542;
assign b1c0a8 = hmaster0_p & b1c85a | !hmaster0_p & b1c0a7;
assign d357dd = hgrant1_p & d357d5 | !hgrant1_p & d357dc;
assign v9f7de3 = hgrant4_p & v9f7d22 | !hgrant4_p & v9f7de1;
assign v8ccbe6 = hlock1_p & v8ccb6b | !hlock1_p & v845542;
assign c3ce7b = hmaster1_p & c3ce78 | !hmaster1_p & c3ce7a;
assign v9f7d83 = hlock0_p & v9f7d81 | !hlock0_p & v9f7d82;
assign v9ea5dd = hready_p & v9ea4a4 | !hready_p & v9ea5dc;
assign ad501a = hmaster0_p & ad5013 | !hmaster0_p & ad5019;
assign ad4265 = hready & ad4e48 | !hready & ad4264;
assign ad3d31 = decide_p & ad4409 | !decide_p & ad3d30;
assign ad40f2 = hbusreq2 & ad5018 | !hbusreq2 & c3d2d9;
assign v9e9fbd = hbusreq2_p & v9e9fba | !hbusreq2_p & v9e9fbc;
assign v9ea623 = hbusreq2 & v9ea622 | !hbusreq2 & v9ea3fa;
assign c3d31b = hbusreq4_p & c3d319 | !hbusreq4_p & c3d31a;
assign bd58fd = hgrant2_p & bd5bab | !hgrant2_p & !bd58fc;
assign dc4f8f = hmaster2_p & dc4f7d | !hmaster2_p & !ade5d5;
assign ad46de = hbusreq4_p & ad46dd | !hbusreq4_p & v845542;
assign ade565 = hlock4_p & ade564 | !hlock4_p & !ade563;
assign b1c582 = hbusreq1_p & b1caf9 | !hbusreq1_p & b1c581;
assign ad43c4 = hmastlock_p & ad43c3 | !hmastlock_p & v845542;
assign c3d39c = hbusreq4_p & v845542 | !hbusreq4_p & c3d39b;
assign ade542 = hmaster0_p & ade540 | !hmaster0_p & ade541;
assign b05989 = hlock4_p & b05987 | !hlock4_p & !b05988;
assign b573ff = hmaster1_p & b573fe | !hmaster1_p & v845542;
assign v9f786d = hlock3 & v9f786c | !hlock3 & v9f786b;
assign ad4e57 = hbusreq1_p & ad4e52 | !hbusreq1_p & ad4e56;
assign v9e9fb0 = hmaster1_p & v9e9faf | !hmaster1_p & v9e9f9f;
assign b058ea = hmaster2_p & b058a3 | !hmaster2_p & b058e9;
assign d35802 = hbusreq2_p & d357af | !hbusreq2_p & d35801;
assign ad4e59 = hbusreq2 & ad4e58 | !hbusreq2 & v845542;
assign c3d32c = hgrant1_p & v84554d | !hgrant1_p & c3d32b;
assign c3d734 = hmaster0_p & c3d6dc | !hmaster0_p & c3d6b2;
assign b1c821 = hmaster0_p & b1c80e | !hmaster0_p & b1c820;
assign ad4e50 = hbusreq2 & ad4e4a | !hbusreq2 & ad4e4f;
assign bd58a7 = hgrant4_p & v845542 | !hgrant4_p & !bd58a5;
assign bd56cd = hgrant3_p & bd5e29 | !hgrant3_p & !bd56cc;
assign d3569d = jx0_p & d35abd | !jx0_p & d3569c;
assign ba7c6b = hgrant1_p & v845558 | !hgrant1_p & ba7c64;
assign d35a94 = decide_p & v845542 | !decide_p & !v84556c;
assign b57441 = decide_p & b57940 | !decide_p & b57440;
assign v9f76ca = hmaster1_p & v9f76c7 | !hmaster1_p & v9f76c9;
assign b05965 = hlock3 & b05964 | !hlock3 & b05963;
assign df51bf = hgrant2_p & df51bc | !hgrant2_p & !df51be;
assign b0592d = hbusreq2_p & b0592a | !hbusreq2_p & b0592c;
assign ad42a2 = hbusreq1 & ad4d9c | !hbusreq1 & v845542;
assign v9ea5e7 = hbusreq2_p & v9ea5e2 | !hbusreq2_p & v9ea5e6;
assign ad41a5 = hbusreq2 & ad5037 | !hbusreq2 & ad5038;
assign c3d37d = hmaster0_p & c3d377 | !hmaster0_p & c3d37c;
assign c5c979 = hgrant2_p & c5c96d | !hgrant2_p & c5c978;
assign bd5932 = hbusreq0_p & d355a8 | !hbusreq0_p & bd5b93;
assign bd57ea = hmaster0_p & bd57e9 | !hmaster0_p & bd57cd;
assign c3d2db = hbusreq2 & c3d2d8 | !hbusreq2 & c3d2da;
assign b1c77e = hbusreq2_p & b1c77a | !hbusreq2_p & b1c77d;
assign c74b29 = start_p & v845542 | !start_p & !c749e5;
assign ad3ccd = hmaster2_p & ad3ccc | !hmaster2_p & ad447b;
assign v9f7657 = hbusreq0_p & v9f7dce | !hbusreq0_p & v9f7656;
assign b1c095 = hgrant2_p & v845542 | !hgrant2_p & b1c094;
assign bd5866 = hgrant4_p & bd5757 | !hgrant4_p & bd5865;
assign v9ea4e4 = hready_p & v9ea436 | !hready_p & v9ea4e3;
assign bd5b88 = locked_p & bd5b87 | !locked_p & !v845542;
assign ad448a = hmaster2_p & b1c70e | !hmaster2_p & !ad4489;
assign d35571 = hbusreq2 & d354f4 | !hbusreq2 & !d354f5;
assign b1c743 = hbusreq0 & b1c742 | !hbusreq0 & v845542;
assign d35c0b = hlock4_p & d359e8 | !hlock4_p & !v845542;
assign ad4319 = hbusreq1 & ad4feb | !hbusreq1 & v845542;
assign bd5913 = hbusreq1_p & bd5912 | !hbusreq1_p & v84556c;
assign d354f2 = hbusreq4_p & d354bc | !hbusreq4_p & !v845542;
assign v9ea43f = hmaster0_p & v9ea43e | !hmaster0_p & v9ea404;
assign b1c774 = hbusreq4 & b1c76f | !hbusreq4 & b1c773;
assign v9f77bd = locked_p & v9f7743 | !locked_p & v9f772b;
assign b058e3 = hmaster0_p & b058b5 | !hmaster0_p & b058c7;
assign d354e0 = hmaster0_p & d354d6 | !hmaster0_p & d354df;
assign b059d5 = hgrant4_p & b059c2 | !hgrant4_p & v9f7d42;
assign d35a70 = hlock2_p & d35a6e | !hlock2_p & !d35a6f;
assign d3564d = hgrant4_p & v845542 | !hgrant4_p & !d3564b;
assign c3d6fa = hmaster2_p & c3d6f4 | !hmaster2_p & !c3d6f9;
assign adec8d = hmastlock_p & adec8c | !hmastlock_p & v845542;
assign d35a3f = hburst0 & d35a3c | !hburst0 & d35a3e;
assign ad4847 = hready & ad4d96 | !hready & !ad4846;
assign b1c764 = hbusreq0 & b1c763 | !hbusreq0 & !v845542;
assign d356e9 = hlock2_p & d356e6 | !hlock2_p & d356e8;
assign v9f7df3 = hlock3 & v9f7df2 | !hlock3 & v9f7def;
assign c3cee0 = hready & c3cedf | !hready & !v845542;
assign c3d5d3 = hmastlock_p & v84557c | !hmastlock_p & !v845542;
assign d35739 = hmaster1_p & d35736 | !hmaster1_p & d35738;
assign b574d4 = hbusreq3 & b574d2 | !hbusreq3 & b574d3;
assign bd5b81 = locked_p & bd5b80 | !locked_p & !v845542;
assign v9f7db2 = stateG10_4_p & v9f7dae | !stateG10_4_p & v9f7db0;
assign v8cc0e0 = hbusreq1 & v8cc0de | !hbusreq1 & v8cc0df;
assign bd57c1 = stateA1_p & bd57c0 | !stateA1_p & c5c88b;
assign b1c063 = hgrant4_p & b1c731 | !hgrant4_p & !b1c062;
assign b1c72c = hmaster1_p & b1c71f | !hmaster1_p & b1c72b;
assign b1c7ce = hbusreq1_p & b1c7cc | !hbusreq1_p & b1c7cd;
assign d357bc = hbusreq2 & d357b8 | !hbusreq2 & d357bb;
assign b1c0ac = decide_p & b1c0ab | !decide_p & b1d013;
assign b05a09 = hbusreq4_p & b05a07 | !hbusreq4_p & b05a08;
assign v8cc0e4 = hbusreq3 & v8cc0e1 | !hbusreq3 & v8cc0e2;
assign v9f7d01 = hbusreq3 & v9f7cff | !hbusreq3 & v9f7d00;
assign d35993 = hlock1_p & d35991 | !hlock1_p & !d35992;
assign v9e9fe9 = jx2_p & v9e9e73 | !jx2_p & v9e9fe8;
assign v8cc47f = hlock4 & v8ccbd8 | !hlock4 & v8cc47d;
assign d3565d = hbusreq2_p & d3565c | !hbusreq2_p & d35aa7;
assign v9f76d0 = hbusreq2_p & v9f76cd | !hbusreq2_p & v9f76cf;
assign c3d760 = decide_p & c3d72a | !decide_p & c3d75f;
assign d35a16 = hmaster2_p & d35a12 | !hmaster2_p & d35a15;
assign v9e9f71 = hbusreq1 & v9e9f70 | !hbusreq1 & v9e9f68;
assign ad436d = hmaster1_p & ad436c | !hmaster1_p & ad4297;
assign v8cc4e0 = decide_p & v845542 | !decide_p & v8ccb6e;
assign dc4fd7 = hbusreq2 & dc4fd6 | !hbusreq2 & dc4f61;
assign ade5d8 = hbusreq0 & ade4e3 | !hbusreq0 & ade5d7;
assign ad4693 = hmaster2_p & ad4692 | !hmaster2_p & v845542;
assign df5146 = hbusreq1_p & df5145 | !hbusreq1_p & v845542;
assign c3d6ed = hbusreq4_p & c3d6eb | !hbusreq4_p & c3d6ec;
assign c3cf34 = jx2_p & c3ce33 | !jx2_p & c3cf33;
assign dc4f81 = hbusreq4 & dc4f77 | !hbusreq4 & dc4f80;
assign v9f7d44 = hbusreq4_p & v9f7d40 | !hbusreq4_p & !v9f7d43;
assign ad3d27 = decide_p & ad43a2 | !decide_p & ad3d26;
assign ad4409 = hbusreq2_p & ad4408 | !hbusreq2_p & ad4407;
assign c3d2e2 = decide_p & c3d2d5 | !decide_p & !c3d2e1;
assign b579df = hlock4 & b579ce | !hlock4 & b579d5;
assign d3594e = hburst0 & dc5318 | !hburst0 & d3594d;
assign v9f7d66 = hmaster0_p & v9f7d5a | !hmaster0_p & v9f7d5e;
assign ba7c68 = hmaster1_p & ba7c64 | !hmaster1_p & ba7c67;
assign dc5010 = stateG10_4_p & ade563 | !stateG10_4_p & !dc500f;
assign c5c92e = hmastlock_p & c5c92d | !hmastlock_p & v845542;
assign b57a0d = hgrant2_p & b579f1 | !hgrant2_p & b579ea;
assign v9e9f92 = hmaster2_p & v9e9f91 | !hmaster2_p & v9ea4d8;
assign b1c847 = hmaster2_p & d35a9c | !hmaster2_p & !b1c846;
assign b05981 = hgrant4_p & b058d0 | !hgrant4_p & !b05980;
assign cc36fa = stateG10_4_p & cc36f2 | !stateG10_4_p & cc36f9;
assign bd5872 = hgrant0_p & bd576b | !hgrant0_p & !adec89;
assign ad4365 = hgrant2_p & ad4364 | !hgrant2_p & !ad4360;
assign bd58c9 = stateG10_4_p & bd58c6 | !stateG10_4_p & !bd58c8;
assign v8cc50c = decide_p & v8cc4f4 | !decide_p & v8cc50a;
assign ad441c = hmaster1_p & ad441b | !hmaster1_p & ad4419;
assign d356b9 = hmaster1_p & d356af | !hmaster1_p & d356b8;
assign b1c0b4 = jx0_p & b1c70d | !jx0_p & b1c0b3;
assign v84555a = hlock4_p & v845542 | !hlock4_p & !v845542;
assign v9f76e1 = stateA1_p & v845542 | !stateA1_p & !v9f76e0;
assign v9ea617 = decide_p & v9ea5f5 | !decide_p & v9ea616;
assign d35641 = hgrant4_p & v845542 | !hgrant4_p & !d3563f;
assign b1cf42 = hmaster0_p & v845542 | !hmaster0_p & b1cf41;
assign v8cc785 = hgrant3_p & v8ccbdc | !hgrant3_p & v8cc784;
assign ad4ff2 = hmaster0_p & dc4fcc | !hmaster0_p & ad4ff1;
assign v9f7deb = hbusreq4 & v9f7de9 | !hbusreq4 & v9f7dea;
assign v84556a = decide_p & v845542 | !decide_p & !v845542;
assign b059b1 = hmaster2_p & b05952 | !hmaster2_p & b059b0;
assign dc5386 = hready_p & v845542 | !hready_p & dc5385;
assign v8ccbee = hbusreq4_p & v8ccbec | !hbusreq4_p & v845542;
assign b1c739 = hbusreq0 & b1c738 | !hbusreq0 & v845542;
assign bd58f5 = hready_p & bd58ed | !hready_p & bd58f4;
assign c3d6de = hmaster1_p & c3d6dd | !hmaster1_p & c3d6d2;
assign bd56df = decide_p & bd56de | !decide_p & v845542;
assign ad4309 = hbusreq1 & ad4f5e | !hbusreq1 & v845542;
assign v9f7678 = hlock3 & v9f7e32 | !hlock3 & v9f7e39;
assign b57410 = hbusreq1 & b5740e | !hbusreq1 & b5740f;
assign c3cef9 = hgrant1_p & v84554d | !hgrant1_p & c3cef8;
assign ad42a0 = hlock1_p & ad429d | !hlock1_p & !ad429f;
assign v9f76f5 = hlock4 & v9f76f2 | !hlock4 & v9f76f4;
assign v8cc7de = hmaster2_p & v845542 | !hmaster2_p & v8cc7dd;
assign v9e9f95 = hbusreq4 & v9e9f94 | !hbusreq4 & v9e9f8e;
assign ad46a5 = hburst0 & ad46a4 | !hburst0 & ade54d;
assign v9f764a = hgrant1_p & v9f7e3a | !hgrant1_p & v9f7649;
assign b1c5b7 = hmaster2_p & v845542 | !hmaster2_p & b1c5b6;
assign v9f7ca1 = hmaster2_p & v9f7c9c | !hmaster2_p & !v9f7ca0;
assign v8cc483 = hlock1 & v8ccbd8 | !hlock1 & v8cc482;
assign v9ea609 = hbusreq3 & v9ea606 | !hbusreq3 & v9ea608;
assign b1c795 = hgrant0_p & v84556c | !hgrant0_p & !bd57fb;
assign v8cc7cf = hmaster0_p & v8cc7b8 | !hmaster0_p & v8cc7ce;
assign ad3d1a = hbusreq2 & ad3d18 | !hbusreq2 & ad3d19;
assign b57a0e = hbusreq2_p & b579eb | !hbusreq2_p & b57a0d;
assign c3cf0f = hmaster0_p & c3cf0e | !hmaster0_p & !c3d2be;
assign dc4f63 = hmaster1_p & dc4f62 | !hmaster1_p & v84556c;
assign df51d1 = hgrant3_p & df5531 | !hgrant3_p & df51d0;
assign ad42db = decide_p & ad42cf | !decide_p & ad42da;
assign d359a3 = hmaster2_p & d359a2 | !hmaster2_p & v845542;
assign v9e9f50 = hgrant4_p & v9e9ee7 | !hgrant4_p & v9e9f4f;
assign ad4158 = hbusreq0 & ad4154 | !hbusreq0 & ad4157;
assign ade4a9 = hbusreq0_p & adec89 | !hbusreq0_p & adeca1;
assign adea9c = hlock4_p & adea9b | !hlock4_p & !v845542;
assign c3ce27 = decide_p & c3ce26 | !decide_p & !c3d36c;
assign b1cfd1 = hgrant1_p & v845542 | !hgrant1_p & b1cfd0;
assign bd5925 = hmaster2_p & v845542 | !hmaster2_p & bd5924;
assign ad5062 = hmaster2_p & ad505b | !hmaster2_p & !ad5061;
assign v9f7783 = hbusreq2_p & v9f7780 | !hbusreq2_p & v9f7782;
assign ad3d56 = hmaster0_p & ad3d50 | !hmaster0_p & ad3d1a;
assign ad4556 = hmaster2_p & ad4554 | !hmaster2_p & ad4555;
assign v8cc502 = hmaster0_p & v8cc501 | !hmaster0_p & v8ccbf6;
assign b574b4 = hbusreq0 & b574b3 | !hbusreq0 & b57942;
assign c3d2be = hbusreq4 & c3d2bc | !hbusreq4 & !c3d2bd;
assign adeaa6 = hgrant1_p & v845542 | !hgrant1_p & !adeaa5;
assign c3ce20 = hmaster1_p & c3ce1d | !hmaster1_p & c3ce1f;
assign d356ee = hlock2_p & d356ec | !hlock2_p & d356ed;
assign v9ea61a = hmaster0_p & v9ea3e7 | !hmaster0_p & v9f20a1;
assign b1c6cc = decide_p & b1c6be | !decide_p & b1c6cb;
assign b1c0b2 = hbusreq3_p & b1c098 | !hbusreq3_p & b1c0b1;
assign d356f1 = decide_p & d356f0 | !decide_p & v84556c;
assign d3556d = hmaster1_p & d3556c | !hmaster1_p & d354db;
assign b1c4c8 = hbusreq4_p & d35918 | !hbusreq4_p & b1c843;
assign d3570f = hbusreq2 & d356c0 | !hbusreq2 & !d356c1;
assign ad48b4 = hmaster0_p & ad48b3 | !hmaster0_p & v845551;
assign ad470d = hready & ad4709 | !hready & ad470c;
assign bd5b74 = hlock2_p & bd5b73 | !hlock2_p & v845542;
assign c3d70e = hgrant1_p & c3d70b | !hgrant1_p & c3d70d;
assign c3d2d2 = hmaster1_p & c3d2ce | !hmaster1_p & c3d2d1;
assign d356ea = hbusreq2_p & d356e9 | !hbusreq2_p & d356e8;
assign ad4358 = hmaster0_p & ad4344 | !hmaster0_p & ad42d3;
assign ad4736 = hmaster0_p & ad4734 | !hmaster0_p & ad4735;
assign d356f7 = hbusreq1_p & d356f6 | !hbusreq1_p & v845542;
assign ad4ecd = hlock0_p & v845542 | !hlock0_p & ad4ecc;
assign b05929 = hmaster1_p & b05928 | !hmaster1_p & b05926;
assign ad4ed7 = hgrant0_p & ad4e47 | !hgrant0_p & v845542;
assign b574be = hlock2 & b579c5 | !hlock2 & b574bd;
assign ad4774 = hlock4_p & ad4dce | !hlock4_p & !ad45e6;
assign c3d5c6 = hmaster2_p & c3d5ba | !hmaster2_p & adeaa5;
assign c3cf06 = hbusreq0 & c3cf05 | !hbusreq0 & v845542;
assign c5c96a = hmaster2_p & c5c968 | !hmaster2_p & c5c88e;
assign b1c7f7 = hmaster1_p & b1c7f6 | !hmaster1_p & b1c7e3;
assign b8f749 = hgrant1_p & v845542 | !hgrant1_p & b8f748;
assign d35a39 = hmaster1_p & d35a38 | !hmaster1_p & v84556c;
assign d35915 = hlock1_p & d35914 | !hlock1_p & d3590a;
assign c3d4df = hbusreq4_p & c3d4de | !hbusreq4_p & !adeaa4;
assign v9f77b9 = decide_p & v9f7784 | !decide_p & v9f77b8;
assign b8f6e0 = hready_p & v845542 | !hready_p & v845562;
assign b1c81f = hbusreq1_p & v845542 | !hbusreq1_p & b1c81e;
assign bd581c = hbusreq4_p & bd5819 | !hbusreq4_p & bd581b;
assign d3542f = hlock1_p & d3542b | !hlock1_p & d3542e;
assign v8cc0cf = hlock1 & v8ccbd8 | !hlock1 & v8cc0ce;
assign ad4e72 = stateG10_4_p & ad4e6f | !stateG10_4_p & !ad4e71;
assign dc4fda = hbusreq3 & dc4fd9 | !hbusreq3 & v845542;
assign ad4756 = hready_p & ad4725 | !hready_p & ad4755;
assign b05907 = hbusreq2 & b05905 | !hbusreq2 & b05906;
assign v8cc455 = decide_p & v8cc434 | !decide_p & v8cc43f;
assign b1c4a6 = hbusreq0 & b1caf5 | !hbusreq0 & b1c4a5;
assign v9ea4ac = hbusreq0_p & v9ea3ec | !hbusreq0_p & v9ea4a6;
assign d35a76 = hmaster0_p & d35a75 | !hmaster0_p & d35a4c;
assign ad442f = hbusreq0 & ad442e | !hbusreq0 & v845542;
assign dc4feb = hbusreq4_p & dc4fe8 | !hbusreq4_p & dc4fea;
assign v9f77ce = hbusreq1 & v9f77cc | !hbusreq1 & v9f77cd;
assign v9f7d3b = hmaster2_p & v9f7d3a | !hmaster2_p & v9f7c9d;
assign v8ccbdd = hmaster0_p & v845542 | !hmaster0_p & v8ccb6b;
assign bd57f4 = hmastlock_p & bd5783 | !hmastlock_p & v845542;
assign d356bc = hbusreq3 & d356bb | !hbusreq3 & d356ad;
assign v845556 = hlock3_p & v845542 | !hlock3_p & !v845542;
assign ad4f7d = hbusreq4 & ad4f73 | !hbusreq4 & ad4f7c;
assign c5c88d = hmastlock_p & c5c88c | !hmastlock_p & !v845542;
assign ad42fb = hgrant2_p & ad42e9 | !hgrant2_p & ad42fa;
assign ade4ab = hbusreq4_p & ade4aa | !hbusreq4_p & v845542;
assign ad4f9f = hmaster1_p & ad4f5a | !hmaster1_p & ad4f9e;
assign b1c08e = decide_p & b1c08d | !decide_p & b1c866;
assign b57a86 = hbusreq3 & b57a84 | !hbusreq3 & b57a85;
assign v8ccb8c = hmaster1_p & v8ccb89 | !hmaster1_p & v8ccb81;
assign v8cc0c4 = hmaster2_p & v845542 | !hmaster2_p & v8cc0c3;
assign d356bf = hbusreq2_p & d356b9 | !hbusreq2_p & d356be;
assign d35a2a = hmaster0_p & d35a1e | !hmaster0_p & d35a29;
assign b1c079 = hbusreq1_p & b1c7ae | !hbusreq1_p & b1c074;
assign b05a5c = hbusreq0_p & b0594f | !hbusreq0_p & b05a5b;
assign c3d5c1 = hbusreq0 & c3d5be | !hbusreq0 & c3d5c0;
assign v8cc437 = hbusreq4_p & v8ccbeb | !hbusreq4_p & v8cc436;
assign b1c04f = hmaster1_p & b1c04e | !hmaster1_p & b1c790;
assign d35a1a = hbusreq3 & d35a19 | !hbusreq3 & v845542;
assign df512a = hgrant2_p & v845542 | !hgrant2_p & !df5129;
assign b579cb = hbusreq4_p & b579c9 | !hbusreq4_p & b579ca;
assign c3d5cd = hbusreq2 & c3d5cc | !hbusreq2 & c3d306;
assign v9f76b9 = hmaster1_p & v9f76b8 | !hmaster1_p & v9f7ce9;
assign c3d5d8 = hmaster2_p & c3d5d7 | !hmaster2_p & v845542;
assign ad4483 = hmaster2_p & ad447b | !hmaster2_p & ad4482;
assign d359cc = hbusreq1_p & d359c7 | !hbusreq1_p & !d359cb;
assign v9ea574 = hbusreq4_p & v9ea3fe | !hbusreq4_p & v9ea4b6;
assign b1cffb = hmaster2_p & b1cfbf | !hmaster2_p & b1cffa;
assign d3597c = hlock3_p & d35903 | !hlock3_p & d3597b;
assign ac1467 = hgrant4_p & v845542 | !hgrant4_p & !ac1466;
assign v9f767a = hlock2 & v9f7e32 | !hlock2 & v9f7679;
assign d35529 = hbusreq0 & d35526 | !hbusreq0 & d35528;
assign ad4f74 = hbusreq4_p & ad4f65 | !hbusreq4_p & ad4e98;
assign ade5c1 = hbusreq3 & ade583 | !hbusreq3 & v9041a4;
assign df515f = hlock1_p & df515d | !hlock1_p & df515e;
assign b57a71 = hbusreq3 & b57a6f | !hbusreq3 & b57a70;
assign c5c3b6 = hready_p & c5c953 | !hready_p & !c5c3b5;
assign v9f77bf = hgrant4_p & v9f772b | !hgrant4_p & v9f77be;
assign c5c932 = hgrant1_p & c5c931 | !hgrant1_p & c5c8f4;
assign ade64e = decide_p & ade64d | !decide_p & adeaa7;
assign ad45bb = hbusreq4_p & ad45ba | !hbusreq4_p & v845542;
assign b1c6b7 = hbusreq1 & b1cfc8 | !hbusreq1 & b1cfd0;
assign c3d516 = hready & c3d515 | !hready & !c3d47b;
assign d35511 = hmaster2_p & d35419 | !hmaster2_p & d35510;
assign c3d722 = hmaster1_p & c3d721 | !hmaster1_p & c3d67c;
assign b1c6fd = hbusreq2_p & b1c6be | !hbusreq2_p & b1c6fc;
assign df5174 = hbusreq2 & df5171 | !hbusreq2 & df5173;
assign v9e9faa = hgrant1_p & v9e9eed | !hgrant1_p & v9e9f79;
assign ad4150 = hgrant4_p & ad4f38 | !hgrant4_p & v845542;
assign b05a5e = hgrant4_p & b058a3 | !hgrant4_p & b05a5d;
assign ad46f9 = hgrant2_p & ad46f2 | !hgrant2_p & !ad46f8;
assign c3d70c = hmaster2_p & c3d669 | !hmaster2_p & !c3d6ed;
assign ad42e1 = hbusreq1 & ad4e4e | !hbusreq1 & v845542;
assign d3550a = hmaster2_p & d35419 | !hmaster2_p & d35509;
assign bd57af = hgrant1_p & bd57ae | !hgrant1_p & dc4f81;
assign ad4f46 = hbusreq3 & ad4f45 | !hbusreq3 & v845542;
assign ad431c = hmaster0_p & ad4318 | !hmaster0_p & ad431b;
assign v845572 = hgrant2_p & v845542 | !hgrant2_p & !v845542;
assign ad3cc8 = hmaster0_p & ad4411 | !hmaster0_p & ad440e;
assign d35a96 = hmaster0_p & v845542 | !hmaster0_p & d35a95;
assign v9f7cc4 = hmaster2_p & v9f7c9c | !hmaster2_p & v9f7c9f;
assign v9ea429 = hmaster1_p & v9ea428 | !hmaster1_p & v845542;
assign df5537 = hgrant2_p & v845542 | !hgrant2_p & !df5536;
assign b5740b = hbusreq0 & b57409 | !hbusreq0 & b5740a;
assign dc500e = hgrant4_p & v84556c | !hgrant4_p & ade563;
assign v8ccbfa = hgrant2_p & v845542 | !hgrant2_p & v8ccbf8;
assign d35a40 = locked_p & d35a3f | !locked_p & !v845542;
assign ad416d = hgrant2_p & v845542 | !hgrant2_p & ad416c;
assign ad4ee9 = hbusreq0 & ad4edf | !hbusreq0 & ad4ee8;
assign c3d518 = hbusreq3 & c3d513 | !hbusreq3 & c3d517;
assign c3d511 = hbusreq4 & c3d510 | !hbusreq4 & v845564;
assign d3597a = hgrant2_p & d3595b | !hgrant2_p & d35920;
assign adeab2 = decide_p & adeab1 | !decide_p & v845542;
assign ad481e = hmaster0_p & ad481c | !hmaster0_p & ad481d;
assign c5c937 = hbusreq0_p & c5c8fc | !hbusreq0_p & !c5c936;
assign ad439d = hbusreq3 & ad4393 | !hbusreq3 & v845542;
assign ad436b = hbusreq2_p & ad4366 | !hbusreq2_p & !ad436a;
assign d3572e = hbusreq1_p & d356c5 | !hbusreq1_p & v845542;
assign d356c7 = hlock1_p & d359e9 | !hlock1_p & !v845542;
assign dc4f7c = hburst0 & dc4f78 | !hburst0 & dc4f7b;
assign ad3cd8 = hready & ad3cd6 | !hready & !ad3cd7;
assign ad4e44 = hbusreq2 & ad4e43 | !hbusreq2 & v845542;
assign d355ae = hbusreq2_p & d355ad | !hbusreq2_p & v845542;
assign b1c082 = hgrant4_p & b1c7b6 | !hgrant4_p & b1c066;
assign d3541a = hlock4_p & v845542 | !hlock4_p & d3590d;
assign v9f7c99 = busreq_p & v9f7c95 | !busreq_p & v9f7c96;
assign bd58d9 = hlock2_p & bd589a | !hlock2_p & !bd58d8;
assign c3cf28 = decide_p & c3cf23 | !decide_p & c3cf15;
assign d356a8 = hbusreq1_p & d356a7 | !hbusreq1_p & v845542;
assign d359d3 = hbusreq4_p & d359d1 | !hbusreq4_p & d359d2;
assign ad426a = hmaster2_p & v845542 | !hmaster2_p & ad4566;
assign c5c971 = hbusreq4_p & c5c96f | !hbusreq4_p & c5c970;
assign bd5906 = jx0_p & bd5bb3 | !jx0_p & bd5905;
assign d35951 = hlock1_p & d35950 | !hlock1_p & d3590a;
assign b57508 = hgrant3_p & b57504 | !hgrant3_p & b57507;
assign bd575a = hbusreq2 & bd5759 | !hbusreq2 & v845542;
assign ad42ca = hmaster1_p & ad42c9 | !hmaster1_p & ad42bd;
assign b05a83 = hgrant2_p & b05a57 | !hgrant2_p & b05a82;
assign v9f7cb7 = hmaster2_p & v9f7ca5 | !hmaster2_p & !v9f7cb6;
assign ad42f3 = hgrant1_p & v845542 | !hgrant1_p & ad42f2;
assign bd581a = hgrant4_p & v845542 | !hgrant4_p & !bd5806;
assign ad4411 = hready & ad4410 | !hready & !v845542;
assign ad4daf = hlock0_p & ad4d9a | !hlock0_p & v845542;
assign b5742b = hmaster0_p & b57416 | !hmaster0_p & b5742a;
assign ad476c = hbusreq2 & ad45b6 | !hbusreq2 & ad476b;
assign b1c5e7 = hmaster2_p & b1cfbf | !hmaster2_p & b1c5e6;
assign c3d5ca = hbusreq4 & c3d5c7 | !hbusreq4 & !c3d5c9;
assign b1cc05 = decide_p & b1cc04 | !decide_p & b1c866;
assign c5c9ae = hgrant2_p & c5c9ad | !hgrant2_p & c5c978;
assign ad43cf = hbusreq0_p & ad4de2 | !hbusreq0_p & v845542;
assign c3d532 = hmaster1_p & c3d52e | !hmaster1_p & c3d531;
assign b1c50e = hready_p & b1c82d | !hready_p & b1c50d;
assign ad5044 = hbusreq4_p & ad5042 | !hbusreq4_p & ad5043;
assign ad3d4f = hmaster1_p & ad3d4e | !hmaster1_p & ad4419;
assign b05a46 = hmaster0_p & b05a0f | !hmaster0_p & b0593b;
assign dc5074 = hbusreq3 & dc5033 | !hbusreq3 & v845542;
assign d35010 = stateG10_4_p & d3580c | !stateG10_4_p & d3500f;
assign d359e8 = hlock0_p & v845542 | !hlock0_p & d359e7;
assign ad4f25 = hlock2_p & ad4f18 | !hlock2_p & !ad4f24;
assign c5c9a9 = hmaster1_p & c5c9a8 | !hmaster1_p & c5c8eb;
assign v9f76f0 = stateG10_4_p & v9f76ee | !stateG10_4_p & v9f76ef;
assign c3ce5b = hgrant2_p & v845551 | !hgrant2_p & c3ce5a;
assign c3d58e = hmaster2_p & c3d2ad | !hmaster2_p & v845542;
assign dc4f96 = hmaster1_p & dc4f88 | !hmaster1_p & dc4f83;
assign ad46bc = hlock4_p & ad4e89 | !hlock4_p & v845542;
assign df517e = hbusreq1_p & df517d | !hbusreq1_p & v845542;
assign d35626 = hbusreq1_p & d35625 | !hbusreq1_p & d35624;
assign v9f7829 = hbusreq2 & v9f7827 | !hbusreq2 & v9f7828;
assign ad4330 = hbusreq1_p & ad432f | !hbusreq1_p & v845547;
assign v8cc821 = hgrant1_p & v8cc7b1 | !hgrant1_p & v8cc4fe;
assign b1c03b = hbusreq3 & b1c035 | !hbusreq3 & b1c03a;
assign v889629 = hburst0_p & v845542 | !hburst0_p & v84555e;
assign ad42cf = hlock3_p & ad42c7 | !hlock3_p & ad42ce;
assign v9e9ebe = hbusreq2_p & v9e9eaf | !hbusreq2_p & v9e9ebd;
assign c3d2f1 = stateG10_4_p & c3d2ef | !stateG10_4_p & !c3d2f0;
assign c3d535 = hready_p & v845555 | !hready_p & c3d534;
assign v9ea497 = hbusreq2 & v9ea496 | !hbusreq2 & v9ea43b;
assign ad4f94 = hgrant4_p & ad4f3e | !hgrant4_p & v845542;
assign adec89 = locked_p & v845542 | !locked_p & c3d66d;
assign c3d746 = hgrant1_p & c3d6db | !hgrant1_p & c3d745;
assign ade61e = hmaster1_p & ade5b4 | !hmaster1_p & ade5a4;
assign c3d5b2 = hgrant0_p & v845542 | !hgrant0_p & c3d5b1;
assign v9e9ee5 = hbusreq3_p & v9e9ee4 | !hbusreq3_p & v9ea4e5;
assign b059e2 = hbusreq0_p & b0598b | !hbusreq0_p & b0597e;
assign b059c1 = hmastlock_p & b059c0 | !hmastlock_p & !v845542;
assign b57adf = hlock3_p & b57ad3 | !hlock3_p & b5793f;
assign df51cc = hready_p & df51ca | !hready_p & df51cb;
assign b1c78f = hbusreq2 & b1c727 | !hbusreq2 & b1c729;
assign ad504e = hbusreq4_p & ad504c | !hbusreq4_p & ad504d;
assign d35bfb = hmaster1_p & d35bef | !hmaster1_p & d35bfa;
assign bd5b6b = stateA1_p & d35905 | !stateA1_p & ade4b7;
assign ac148a = hmaster2_p & ac1489 | !hmaster2_p & v845542;
assign d3579c = hlock4_p & d3578b | !hlock4_p & v84554a;
assign d35654 = hgrant4_p & v845542 | !hgrant4_p & d35652;
assign dc501f = hbusreq4_p & adeca1 | !hbusreq4_p & dc501e;
assign ad4fbc = stateG10_4_p & cc36fc | !stateG10_4_p & ad4fbb;
assign bd5bb2 = hgrant3_p & bd5ba8 | !hgrant3_p & !bd5bb1;
assign df5183 = hbusreq1_p & df5182 | !hbusreq1_p & v845542;
assign c3d50d = hgrant2_p & v845551 | !hgrant2_p & c3d50c;
assign v8cc797 = hmaster2_p & v845542 | !hmaster2_p & v8cc796;
assign ad4db6 = hbusreq4 & ad4db1 | !hbusreq4 & !ad4db5;
assign v9f7725 = jx1_p & v857463 | !jx1_p & v9f7724;
assign dc5068 = hmaster1_p & dc5017 | !hmaster1_p & dc5067;
assign ad4f2d = hgrant1_p & ad4f2c | !hgrant1_p & ad4ec6;
assign ad45c0 = hready & ad45ad | !hready & !ad45bf;
assign v9f7e3c = hgrant4_p & v9f7cc7 | !hgrant4_p & v9f7dad;
assign ad4402 = hbusreq2_p & ad4401 | !hbusreq2_p & ad4400;
assign d35028 = jx2_p & d3569d | !jx2_p & d35027;
assign v9ea3ed = hbusreq0_p & v9ea3ec | !hbusreq0_p & v9ea3e6;
assign d356e4 = hbusreq1_p & d356e3 | !hbusreq1_p & d35a95;
assign ba7c6f = hgrant2_p & v845558 | !hgrant2_p & ba7c6e;
assign d35503 = hbusreq3 & d35500 | !hbusreq3 & d35502;
assign df51b3 = hmaster0_p & df51b2 | !hmaster0_p & df515b;
assign b059f9 = hbusreq3 & b059ca | !hbusreq3 & b059f8;
assign c3ce5f = hbusreq1 & c3d375 | !hbusreq1 & v845564;
assign v8cc5a7 = hmaster2_p & v8cc491 | !hmaster2_p & v8cc5a6;
assign ade54a = hbusreq1_p & ade547 | !hbusreq1_p & ade549;
assign b574b7 = hready & b574b6 | !hready & b57942;
assign v9f7d13 = hlock0 & v9f7d12 | !hlock0 & v9f7d04;
assign d3543a = hmaster0_p & d35426 | !hmaster0_p & d3542e;
assign v9f7e27 = hgrant1_p & v9f7cbe | !hgrant1_p & v9f7e26;
assign ad3d40 = hbusreq2_p & ad3d3a | !hbusreq2_p & ad3d3f;
assign ad4ddb = hbusreq2_p & ad4dc0 | !hbusreq2_p & ad4dda;
assign v8ccb6e = hmaster1_p & v8ccb6d | !hmaster1_p & v845542;
assign ad414e = hgrant1_p & ad414d | !hgrant1_p & ad4e8e;
assign df54eb = hmaster1_p & v845542 | !hmaster1_p & df54ea;
assign ad503e = hgrant0_p & ad5016 | !hgrant0_p & !v845542;
assign bd577e = hbusreq2_p & bd577b | !hbusreq2_p & v845542;
assign ade4d2 = hbusreq1 & ade4c7 | !hbusreq1 & ade4ce;
assign dc4fe7 = hmaster2_p & dc4fe6 | !hmaster2_p & v845542;
assign v9ea581 = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea574;
assign c3ce6e = hgrant1_p & c3ce6b | !hgrant1_p & c3ce6d;
assign c3d38b = hbusreq1_p & v845542 | !hbusreq1_p & !v845564;
assign df5193 = hbusreq2 & df5192 | !hbusreq2 & !v84554c;
assign ade5a8 = hbusreq2 & ade56f | !hbusreq2 & !ade574;
assign c3d383 = hgrant2_p & c3d36c | !hgrant2_p & c3d382;
assign d357ec = hbusreq0 & d357eb | !hbusreq0 & !v845542;
assign ad3d13 = hmaster1_p & ad3cdc | !hmaster1_p & ad3d12;
assign b57a31 = hgrant2_p & b579b0 | !hgrant2_p & b57a30;
assign dc53b9 = hbusreq1_p & dc538d | !hbusreq1_p & v845542;
assign bd588d = stateG10_4_p & bd5842 | !stateG10_4_p & !bd588c;
assign ad43a9 = hready & ad43a6 | !hready & ad43a8;
assign b1c7a6 = stateG10_4_p & b1c797 | !stateG10_4_p & b1c7a5;
assign c3d727 = hmaster0_p & c3d685 | !hmaster0_p & c3d683;
assign d35580 = hbusreq4_p & d354b4 | !hbusreq4_p & !d35aab;
assign d3568c = decide_p & d3568b | !decide_p & v84556c;
assign c3ce9a = hgrant2_p & v845551 | !hgrant2_p & c3ce99;
assign ad43db = hready & ad43da | !hready & !v845542;
assign adec9a = locked_p & adec99 | !locked_p & !v845542;
assign v8ccbf0 = hgrant0_p & v8ccb6a | !hgrant0_p & v845542;
assign v9f7d4b = hlock2_p & v9f7d48 | !hlock2_p & v9f7d4a;
assign b1c075 = hbusreq1_p & b1c7c9 | !hbusreq1_p & b1c074;
assign b57ac1 = hbusreq0 & b57abf | !hbusreq0 & b57ac0;
assign ad4fc2 = hready & ad4fc1 | !hready & ad4fbe;
assign b05a73 = hbusreq1_p & b0596b | !hbusreq1_p & b05a69;
assign b1c7e9 = hbusreq2 & b1c73f | !hbusreq2 & !v845542;
assign b574c8 = hlock1 & b579ce | !hlock1 & b574c7;
assign ad4dee = hbusreq0 & ad4ded | !hbusreq0 & ad4de2;
assign c3d318 = hgrant0_p & v845542 | !hgrant0_p & v84556c;
assign d35591 = hgrant1_p & d3558a | !hgrant1_p & d35590;
assign b57ae7 = hbusreq2 & b57ae6 | !hbusreq2 & b579e5;
assign ba7c7b = hmaster1_p & ba7c6b | !hmaster1_p & ba7c7a;
assign ad3d19 = hgrant1_p & ad4413 | !hgrant1_p & ad3cfb;
assign ad4ef1 = hbusreq0 & ad4eed | !hbusreq0 & ad4ef0;
assign v9ea60f = hmaster1_p & v9ea603 | !hmaster1_p & v9ea60e;
assign b57a23 = hready_p & b57a12 | !hready_p & b57a22;
assign d35746 = hgrant2_p & d35745 | !hgrant2_p & !d35741;
assign ad42b6 = hmaster2_p & ad42b4 | !hmaster2_p & ad45e6;
assign ad5058 = hbusreq4 & ad5050 | !hbusreq4 & ad5057;
assign v8cc0d0 = hbusreq1 & v8cc0cf | !hbusreq1 & v8ccbd8;
assign v9ea61f = hbusreq2_p & v9ea61e | !hbusreq2_p & v9ea4b1;
assign v9f7da8 = hready & v9f7da7 | !hready & v9f7da3;
assign v9ea58b = hbusreq4 & v9ea58a | !hbusreq4 & v9ea586;
assign ad4fd7 = stateG10_4_p & v84556c | !stateG10_4_p & !ad4fd6;
assign bd576a = hburst0 & v845542 | !hburst0 & bd5769;
assign v9ea4bb = hlock0_p & v9ea3fb | !hlock0_p & v9ea4ba;
assign b1c79b = hbusreq4_p & b1c798 | !hbusreq4_p & !b1c79a;
assign d359dc = hgrant4_p & v845542 | !hgrant4_p & d359ce;
assign v9e9e7e = hready_p & v9ea3e3 | !hready_p & v9e9e7d;
assign c3d362 = hgrant2_p & v845551 | !hgrant2_p & c3d361;
assign v9f7655 = hbusreq4_p & v9f7652 | !hbusreq4_p & !v9f7654;
assign bd5ea3 = hbusreq2 & bd5e9c | !hbusreq2 & bd5ea2;
assign v9f76fb = hgrant1_p & v9f7e05 | !hgrant1_p & v9f76fa;
assign d35985 = hbusreq1_p & d35980 | !hbusreq1_p & d35984;
assign ad4851 = hbusreq2 & ad4850 | !hbusreq2 & v845542;
assign c3d33e = hbusreq4_p & c3d33c | !hbusreq4_p & !c3d33d;
assign b57af6 = decide_p & b57a21 | !decide_p & b57af5;
assign b579c1 = hlock1 & b57942 | !hlock1 & b579c0;
assign b1c786 = hmaster1_p & b1c785 | !hmaster1_p & b1c775;
assign b059b6 = hready & b059b5 | !hready & b0595b;
assign bd5b98 = hmaster1_p & bd5b97 | !hmaster1_p & v84556c;
assign v9e9eda = hmaster1_p & v9ea3fd | !hmaster1_p & v9ea4bd;
assign cc3709 = hready_p & cc3708 | !hready_p & cc36ec;
assign v9ea5b6 = hmaster1_p & v9ea5b5 | !hmaster1_p & v9ea5aa;
assign c3d5a3 = hbusreq3 & c3d5a0 | !hbusreq3 & c3d5a2;
assign c3ceec = hready_p & v845555 | !hready_p & !c3ceeb;
assign ad4df8 = hlock2_p & ad4df3 | !hlock2_p & ad4df7;
assign v9f7818 = hmaster0_p & v9f779b | !hmaster0_p & v9f7790;
assign ad4ea0 = hmaster2_p & ad4e86 | !hmaster2_p & ad4e9f;
assign b1c86b = hbusreq3_p & b1d019 | !hbusreq3_p & b1c86a;
assign c3ceff = hbusreq0_p & c3d373 | !hbusreq0_p & v845542;
assign c3d2b4 = hbusreq3 & c3d2b2 | !hbusreq3 & v845542;
assign b05967 = hlock2 & b05964 | !hlock2 & b05966;
assign d3571c = hlock1_p & d3571b | !hlock1_p & d356ff;
assign dc5057 = stateG10_4_p & ade58d | !stateG10_4_p & !dc5056;
assign c3d71e = hmaster0_p & c3d6b5 | !hmaster0_p & c3d685;
assign ad4896 = hbusreq2 & ad4895 | !hbusreq2 & v845542;
assign d35587 = hbusreq1_p & d354b7 | !hbusreq1_p & d35582;
assign ad3d0d = hbusreq4_p & v845542 | !hbusreq4_p & !ad3d0c;
assign v8cc036 = hbusreq3_p & v8cc81c | !hbusreq3_p & v8cc035;
assign v9ea47d = hlock0 & v9ea46d | !hlock0 & v9ea47a;
assign v8cc5b1 = hgrant1_p & v845542 | !hgrant1_p & v8cc5b0;
assign v9e9eed = hmaster2_p & v9e9ee7 | !hmaster2_p & v9e9eec;
assign ad4fd0 = hready & ad4fcb | !hready & ad4fcf;
assign ad42d5 = hbusreq1 & ad5012 | !hbusreq1 & v845547;
assign ad475b = hmaster0_p & ad4758 | !hmaster0_p & ad4593;
assign dc504f = hburst0 & adea98 | !hburst0 & dc504e;
assign ade544 = hbusreq2 & ade4ac | !hbusreq2 & ade4ad;
assign v9f76df = hburst0_p & v9f7cf2 | !hburst0_p & !v9f76de;
assign ad43be = hbusreq2_p & ad43bb | !hbusreq2_p & ad43bd;
assign c5c896 = hmastlock_p & c5c895 | !hmastlock_p & !v845542;
assign c3d2cf = hbusreq1 & c3d2c7 | !hbusreq1 & c3d2cb;
assign v9ea401 = hbusreq4_p & v9ea3fb | !hbusreq4_p & v9ea3fe;
assign ad43d1 = hmaster2_p & v845542 | !hmaster2_p & ad43d0;
assign ad4602 = hmaster0_p & ad45ff | !hmaster0_p & ad45fa;
assign b059c5 = hbusreq0 & b059c3 | !hbusreq0 & b059c4;
assign b1cf40 = hbusreq0 & b1cf25 | !hbusreq0 & b1cf3f;
assign ad472c = hmaster0_p & ad460b | !hmaster0_p & ad460a;
assign b57426 = hgrant1_p & v845542 | !hgrant1_p & b57425;
assign b1cbff = hbusreq0 & b1cbfa | !hbusreq0 & b1cbfe;
assign b1c45c = decide_p & b1cafe | !decide_p & b1d013;
assign ad434e = hmaster1_p & ad434d | !hmaster1_p & ad4289;
assign bd5885 = hgrant4_p & v845542 | !hgrant4_p & !bd5865;
assign b1c5ed = hgrant1_p & v845542 | !hgrant1_p & b1c5ec;
assign ad4de7 = hbusreq1 & ad4ddf | !hbusreq1 & ad4de3;
assign d3591d = hmaster0_p & d35917 | !hmaster0_p & d3591c;
assign ad4423 = hbusreq2 & ad4394 | !hbusreq2 & v845542;
assign bd5b73 = hmaster1_p & bd5b72 | !hmaster1_p & v845542;
assign v9ea46c = hbusreq4_p & v9ea46a | !hbusreq4_p & v9ea46b;
assign v9f7775 = hlock2_p & v9f776e | !hlock2_p & v9f7774;
assign v9f7e31 = locked_p & v9f7c9d | !locked_p & !v9f7cc6;
assign d35754 = hgrant1_p & v84554c | !hgrant1_p & d35753;
assign v9ea5d0 = hready & v9ea5cf | !hready & v9ea5cb;
assign ad415f = hgrant1_p & v845542 | !hgrant1_p & ad415e;
assign b058c1 = hbusreq1 & b058bd | !hbusreq1 & b058be;
assign b1c7ec = hmaster1_p & b1c7e8 | !hmaster1_p & b1c7eb;
assign c3d6ca = hbusreq0_p & c3d6c8 | !hbusreq0_p & !c3d6c9;
assign v9f783d = hbusreq2 & v9f783b | !hbusreq2 & v9f783c;
assign c3ceda = hgrant3_p & c3ceba | !hgrant3_p & c3ced9;
assign df516e = hready_p & df5155 | !hready_p & df516d;
assign ad43a4 = hbusreq0_p & ad4fae | !hbusreq0_p & v845542;
assign ad4804 = hready_p & ad4802 | !hready_p & ad4803;
assign b05a21 = hmaster1_p & b05a0e | !hmaster1_p & b05a20;
assign b059d7 = hbusreq4_p & b059d4 | !hbusreq4_p & !b059d6;
assign ad3cce = hbusreq0 & ad3ccd | !hbusreq0 & v845542;
assign adec8e = hburst1 & adec8d | !hburst1 & v845542;
assign ac146c = hmaster0_p & ac1460 | !hmaster0_p & ac146b;
assign b57aea = hgrant2_p & b579b0 | !hgrant2_p & b57ae9;
assign c6d405 = stateG3_1_p & v845542 | !stateG3_1_p & !v845582;
assign ad47ea = hmaster1_p & ad47e9 | !hmaster1_p & ad468c;
assign v8cc470 = hmaster0_p & v845542 | !hmaster0_p & v8ccbd8;
assign b57409 = hmaster2_p & v845542 | !hmaster2_p & b57408;
assign d3571e = hgrant1_p & v845542 | !hgrant1_p & d3571d;
assign ad4efb = hbusreq4_p & ad4ef8 | !hbusreq4_p & ad4efa;
assign dc4f86 = hbusreq3 & dc4f70 | !hbusreq3 & v845542;
assign v8cc0d4 = hbusreq3 & v8cc0d2 | !hbusreq3 & v8cc0d3;
assign b1d010 = hgrant1_p & v845542 | !hgrant1_p & b1d00f;
assign d3590d = hmastlock_p & d3590c | !hmastlock_p & !v845542;
assign c3d368 = hbusreq3 & v845564 | !hbusreq3 & v845542;
assign d3579d = hbusreq4_p & d3579c | !hbusreq4_p & v84554a;
assign ad4da4 = hbusreq3 & ad4da3 | !hbusreq3 & v845542;
assign ade4bb = stateG2_p & v845542 | !stateG2_p & ade4ba;
assign c5c977 = hmaster0_p & c5c976 | !hmaster0_p & !c5c93b;
assign ad41a3 = hbusreq2 & ad5022 | !hbusreq2 & ad5024;
assign b1c85c = hgrant4_p & v84554a | !hgrant4_p & !b1c85b;
assign d3552e = decide_p & d3552d | !decide_p & v84556c;
assign d359b2 = hbusreq3 & d359b1 | !hbusreq3 & v845542;
assign b8f74b = hmaster1_p & b8f6e1 | !hmaster1_p & b8f74a;
assign v8cc4f0 = hbusreq1_p & v8ccb75 | !hbusreq1_p & v8cc4ee;
assign ad502f = locked_p & ad502e | !locked_p & v845542;
assign b573fd = hbusreq2 & b573fb | !hbusreq2 & b573fc;
assign bd58d2 = hbusreq0 & bd58cf | !hbusreq0 & bd58d1;
assign v9ea486 = hgrant1_p & v9ea404 | !hgrant1_p & v9ea46d;
assign ad4137 = hbusreq4_p & ad4136 | !hbusreq4_p & adeaa4;
assign d357a4 = hbusreq0 & d357a3 | !hbusreq0 & v845542;
assign c3d6b8 = hlock0_p & c3d6b7 | !hlock0_p & c3d674;
assign ac1465 = hgrant0_p & ac144e | !hgrant0_p & !v845542;
assign b058ba = hbusreq0 & b058b7 | !hbusreq0 & b058b9;
assign ad42c6 = hlock2_p & ad42be | !hlock2_p & ad42c5;
assign d35a47 = hbusreq4_p & d35a46 | !hbusreq4_p & !d35a45;
assign v9e9ef2 = hmaster1_p & v9e9eea | !hmaster1_p & v9e9ef1;
assign ad4783 = hmaster1_p & ad4602 | !hmaster1_p & ad4781;
assign b1c07f = hbusreq4_p & b1c7d1 | !hbusreq4_p & !b1c07e;
assign d3562e = hmaster1_p & d35624 | !hmaster1_p & d3562a;
assign v845568 = start_p & v845542 | !start_p & !v845542;
assign ad4822 = hmaster0_p & ad4821 | !hmaster0_p & bd5761;
assign v9f7dcd = hbusreq4_p & v9f7dca | !hbusreq4_p & !v9f7dcc;
assign b5741a = hgrant0_p & b57408 | !hgrant0_p & v845542;
assign v9f7801 = hgrant2_p & v9f77bc | !hgrant2_p & v9f7800;
assign d3557e = hmaster2_p & d3557c | !hmaster2_p & d3557d;
assign dc4f74 = hbusreq4_p & ade4c5 | !hbusreq4_p & !ade4d4;
assign dc5048 = stateG10_4_p & ade59c | !stateG10_4_p & dc5047;
assign c3cf0e = hgrant1_p & c3cf0c | !hgrant1_p & c3cf0d;
assign b1c776 = hmaster1_p & b1c75f | !hmaster1_p & b1c775;
assign b1c857 = stateG10_4_p & b1c855 | !stateG10_4_p & !b1c856;
assign b1c72b = hmaster0_p & b1c724 | !hmaster0_p & b1c72a;
assign ac1492 = decide_p & ac1491 | !decide_p & ac147e;
assign ac145d = hgrant1_p & v845542 | !hgrant1_p & ac145c;
assign dc4ffb = hbusreq3 & dc4ffa | !hbusreq3 & v845542;
assign bd5903 = hgrant3_p & bd58f5 | !hgrant3_p & !bd5902;
assign v8cc0f2 = hbusreq2 & v8cc0f1 | !hbusreq2 & v8ccbd8;
assign b1c7aa = stateG10_4_p & b1c79d | !stateG10_4_p & b1c7a9;
assign d35a01 = hgrant0_p & ade598 | !hgrant0_p & v845542;
assign df5532 = hgrant1_p & v84556c | !hgrant1_p & !v845542;
assign dc53a7 = hbusreq2_p & dc53a2 | !hbusreq2_p & dc53a6;
assign v9ea5a8 = hlock2 & v9ea5a5 | !hlock2 & v9ea5a7;
assign b0599c = hlock3 & b0599b | !hlock3 & b0599a;
assign ad4ea5 = hbusreq0 & ad4ea4 | !hbusreq0 & ad4e8e;
assign c3d2da = hbusreq3 & c3d2d9 | !hbusreq3 & v845542;
assign v9f77a3 = hbusreq4 & v9f77a1 | !hbusreq4 & v9f77a2;
assign ade4ce = hmaster2_p & ade4c0 | !hmaster2_p & !ade4cd;
assign v9f76e3 = hgrant0_p & v9f7c9b | !hgrant0_p & v9f76e2;
assign bd5924 = hlock0_p & dc539e | !hlock0_p & bd5923;
assign v9ea466 = stateG10_4_p & v9ea464 | !stateG10_4_p & v9ea465;
assign v9f787a = hgrant2_p & v9f7877 | !hgrant2_p & v9f7879;
assign b579d8 = hbusreq4_p & b579c9 | !hbusreq4_p & b579d7;
assign c3d6bd = hmaster2_p & c3d6aa | !hmaster2_p & c3d6bc;
assign d3594c = hmastlock_p & d3594b | !hmastlock_p & v845542;
assign c3d6e2 = stateG10_4_p & c3d6a5 | !stateG10_4_p & c3d6e1;
assign bd57fa = hmastlock_p & bd57f9 | !hmastlock_p & c3d668;
assign c3d344 = hmaster2_p & c3d343 | !hmaster2_p & v845542;
assign v9ea3e6 = hmastlock_p & v9ea3e5 | !hmastlock_p & v845542;
assign ad4f1e = hready & ad4f1d | !hready & v845542;
assign ad46b2 = hlock1_p & ad46b0 | !hlock1_p & !ad46b1;
assign v8da59f = hgrant4_p & v845542 | !hgrant4_p & !v84556e;
assign c3ce1a = hbusreq3 & c3d376 | !hbusreq3 & c3d37a;
assign v9ea3ea = stateG10_4_p & v9ea3e9 | !stateG10_4_p & !v9ea3e6;
assign ad46d7 = hlock4_p & ad46d6 | !hlock4_p & v845542;
assign b05a7f = hlock2 & b05a7c | !hlock2 & b05a7e;
assign ad4389 = hmaster2_p & v845542 | !hmaster2_p & !ad4388;
assign ad45ad = hbusreq4 & ad45ac | !hbusreq4 & v845542;
assign b05915 = hmaster0_p & b058f6 | !hmaster0_p & b058c7;
assign b1cbf9 = hbusreq4_p & b1cff6 | !hbusreq4_p & b1cfb7;
assign ac147b = hgrant1_p & v845542 | !hgrant1_p & !ac147a;
assign df51ba = hbusreq2 & df5150 | !hbusreq2 & df5142;
assign v8cc826 = hlock2 & v8cc501 | !hlock2 & v8cc825;
assign d35991 = hbusreq1 & d35980 | !hbusreq1 & v845542;
assign v9e9e67 = hmaster0_p & v9ea3ff | !hmaster0_p & v9ea3fa;
assign ad4316 = hbusreq1 & ad4fbe | !hbusreq1 & v845542;
assign b0590e = hbusreq1 & b0590c | !hbusreq1 & b0590d;
assign ad4573 = hbusreq4_p & ad4e54 | !hbusreq4_p & v845542;
assign bd583e = hbusreq4_p & bd574e | !hbusreq4_p & bd583d;
assign c3d6a2 = hmaster0_p & c3d671 | !hmaster0_p & c3d66f;
assign c3d3a0 = hbusreq4_p & v845576 | !hbusreq4_p & c3d39f;
assign d35c08 = hmaster2_p & d35c00 | !hmaster2_p & !d35c07;
assign ade55c = hlock4_p & ade55b | !hlock4_p & !v84556c;
assign ad4704 = hbusreq4 & ad4703 | !hbusreq4 & v845542;
assign v9f788c = hbusreq1 & v9f788a | !hbusreq1 & v9f788b;
assign b1c71f = hmaster0_p & b1c719 | !hmaster0_p & b1c71e;
assign d3575d = decide_p & d35a97 | !decide_p & v84556c;
assign dc502c = hbusreq0 & dc502b | !hbusreq0 & dc5012;
assign v9f7ca4 = hmastlock_p & v9f7ca3 | !hmastlock_p & !v845542;
assign ad3ce2 = hbusreq0_p & ad3ce1 | !hbusreq0_p & !v845542;
assign v9f7d0b = hlock1 & v9f7d05 | !hlock1 & v9f7d0a;
assign b1c619 = hmaster0_p & v845542 | !hmaster0_p & b1c618;
assign ade4db = hmaster2_p & ade4c0 | !hmaster2_p & !ade4da;
assign ad46b9 = hmaster2_p & ad4692 | !hmaster2_p & ad46b8;
assign c3cf17 = hready_p & c3cefe | !hready_p & !c3cf16;
assign bd5806 = hlock0_p & bd5804 | !hlock0_p & !bd5805;
assign dc4f6a = hmaster2_p & ade4bf | !hmaster2_p & !ade4cc;
assign v8cc81c = hgrant3_p & v8cc7aa | !hgrant3_p & v8cc81a;
assign v9e9f6b = hmaster2_p & v9e9ee7 | !hmaster2_p & v9e9f6a;
assign ad4144 = hready & ad4ef0 | !hready & ad4143;
assign v9ea4dd = hgrant2_p & v9ea4c5 | !hgrant2_p & v9ea4dc;
assign b574c3 = hmaster2_p & b574c2 | !hmaster2_p & b579cd;
assign v8cc79a = hlock4 & v8ccb6b | !hlock4 & v8cc799;
assign b059b0 = hbusreq4_p & b059ae | !hbusreq4_p & b059af;
assign ad45e0 = hmaster2_p & v845542 | !hmaster2_p & ad45df;
assign v9f7884 = stateG10_4_p & v9f7882 | !stateG10_4_p & v9f7883;
assign c3cdfd = hlock2_p & c3d5d2 | !hlock2_p & c3cdfc;
assign d35ab3 = hbusreq1_p & v845542 | !hbusreq1_p & d35ab2;
assign c3d680 = hbusreq2_p & c3d67d | !hbusreq2_p & c3d67f;
assign ad4fe4 = hgrant0_p & ad4fce | !hgrant0_p & v845542;
assign b058fb = hready & b058fa | !hready & b058b8;
assign v9f7d9d = hbusreq3 & v9f7d98 | !hbusreq3 & v9f7d9c;
assign v8cc59c = hbusreq1_p & v8ccbd8 | !hbusreq1_p & v8cc59b;
assign dc4fcd = hbusreq2 & dc4fca | !hbusreq2 & dc4fcc;
assign c3d321 = hbusreq4_p & c3d30d | !hbusreq4_p & c3d320;
assign d35a6f = hgrant2_p & v845542 | !hgrant2_p & !d35a6d;
assign v9f7dd7 = hgrant4_p & v9f7ca6 | !hgrant4_p & v9f7d8a;
assign b1c7b7 = hmaster2_p & v845542 | !hmaster2_p & b1c7b6;
assign d35443 = hlock3_p & d3543d | !hlock3_p & d35442;
assign dc4fa0 = hbusreq2 & dc4f9f | !hbusreq2 & dc4f6b;
assign adea96 = hburst0_p & bb9c5a | !hburst0_p & !bbbcd8;
assign v8cc79f = hlock3 & v8ccb6b | !hlock3 & v8cc79e;
assign v9f7689 = hmaster0_p & v9f7d5b | !hmaster0_p & v9f7d5a;
assign ad445d = hbusreq4_p & ad445c | !hbusreq4_p & adeaa4;
assign d35776 = hbusreq0 & d35775 | !hbusreq0 & v845542;
assign b57abf = hmaster2_p & b578f9 | !hmaster2_p & b57abe;
assign v9e9f73 = hgrant0_p & v9ea4b6 | !hgrant0_p & v9ea438;
assign b05a44 = hmaster1_p & b05a41 | !hmaster1_p & b05a43;
assign b579ef = hbusreq2 & b579ee | !hbusreq2 & b57942;
assign c3d4db = hlock4_p & c3d2eb | !hlock4_p & c3d337;
assign v9f7d46 = hmaster2_p & v9f7d44 | !hmaster2_p & v9f7d45;
assign b05a72 = hgrant1_p & b058c7 | !hgrant1_p & b05a71;
assign ad4faf = hmaster2_p & v84556c | !hmaster2_p & ad4fae;
assign d359ef = locked_p & d359ee | !locked_p & v845542;
assign ad4ed2 = hgrant4_p & ad4e47 | !hgrant4_p & v845542;
assign bd57e2 = hmaster1_p & bd57ce | !hmaster1_p & bd57e1;
assign v9e9fde = hmaster1_p & v9e9fdd | !hmaster1_p & v9e9fd0;
assign b05a1f = hgrant1_p & b05942 | !hgrant1_p & b05a1e;
assign v9ea458 = hgrant4_p & v9ea3fe | !hgrant4_p & v9ea457;
assign dc504a = hmaster2_p & dc5045 | !hmaster2_p & dc5049;
assign ad506e = hbusreq2_p & ad5068 | !hbusreq2_p & ad506d;
assign b058b8 = hmaster2_p & b058a3 | !hmaster2_p & v9ea3e9;
assign d357f8 = hbusreq1_p & d3579a | !hbusreq1_p & d357f6;
assign b1c801 = hmaster1_p & b1c800 | !hmaster1_p & b1c745;
assign v8cc783 = decide_p & v8ccbd7 | !decide_p & v8cc782;
assign ade4ed = hmaster1_p & ade4d1 | !hmaster1_p & ade4ec;
assign b05a86 = hmaster1_p & b05a85 | !hmaster1_p & b059f5;
assign ad43b6 = hbusreq4_p & v845542 | !hbusreq4_p & b1c70e;
assign b1c5b9 = hburst1 & d3561d | !hburst1 & bd56cf;
assign v8cc7dc = hmastlock_p & v8cc7db | !hmastlock_p & v845542;
assign ade5c9 = hbusreq3 & ade4d6 | !hbusreq3 & ade4db;
assign v9ea566 = hbusreq4_p & v9ea3e6 | !hbusreq4_p & v9ea4a6;
assign bd57bf = hmastlock_p & bd57be | !hmastlock_p & v845542;
assign ade4b1 = hbusreq3 & ade4a6 | !hbusreq3 & adec93;
assign v9f765f = stateG10_4_p & v9f7d42 | !stateG10_4_p & !v9f765e;
assign ad5041 = hlock0_p & ad503e | !hlock0_p & ad5040;
assign v9f7d74 = hgrant4_p & v9f7c9b | !hgrant4_p & v9f7d72;
assign ad4473 = hmaster0_p & ad4433 | !hmaster0_p & ad4472;
assign dc507e = hmaster0_p & dc4ffb | !hmaster0_p & dc507d;
assign b05a63 = hgrant0_p & b058a3 | !hgrant0_p & !b05a62;
assign c3ceb6 = hmaster0_p & c3ceb5 | !hmaster0_p & c3d2be;
assign d35903 = hbusreq2_p & d358f6 | !hbusreq2_p & d35902;
assign ad3d06 = hgrant4_p & ad3d05 | !hgrant4_p & c3cec2;
assign b1c73f = hbusreq1_p & b1c739 | !hbusreq1_p & b1c73e;
assign ad3d0c = stateG10_4_p & v845542 | !stateG10_4_p & ad3d0b;
assign v9f76bf = hmaster1_p & v9f76be | !hmaster1_p & v9f7d47;
assign ad4554 = hbusreq4_p & d3597f | !hbusreq4_p & v845542;
assign v9f769a = hgrant1_p & v9f7693 | !hgrant1_p & v9f7699;
assign b05944 = hmaster1_p & b0593c | !hmaster1_p & b05943;
assign d35beb = hmaster2_p & d35be8 | !hmaster2_p & !d35bea;
assign c3d2c7 = hready & c3d2c6 | !hready & v845542;
assign d35522 = hbusreq4 & d3551f | !hbusreq4 & d35521;
assign ad4fa4 = hgrant1_p & df553a | !hgrant1_p & ad4f5e;
assign b058f2 = hlock3 & b058ea | !hlock3 & b058f1;
assign v9f77f3 = hgrant1_p & v9f7735 | !hgrant1_p & !v9f77f2;
assign v9f77b7 = hmaster1_p & v9f77b6 | !hmaster1_p & v9f77b0;
assign b579e1 = hready & b579e0 | !hready & b579ce;
assign v9f77ef = hgrant4_p & v9f7734 | !hgrant4_p & !v9f77ee;
assign d3542d = hmaster2_p & d3541f | !hmaster2_p & v84555a;
assign d359f4 = hbusreq4_p & d359f1 | !hbusreq4_p & d359f3;
assign b05996 = hbusreq4 & b05994 | !hbusreq4 & b05995;
assign c5c8f7 = hbusreq1_p & c5c8f6 | !hbusreq1_p & v845542;
assign b57a12 = decide_p & v845542 | !decide_p & b578f3;
assign ba7c79 = hgrant1_p & v845558 | !hgrant1_p & ba7c78;
assign ad4e9c = hbusreq4_p & ad4e99 | !hbusreq4_p & ad4e9b;
assign d35418 = hlock4_p & v845542 | !hlock4_p & d35909;
assign c5c9b3 = decide_p & c5c8e0 | !decide_p & c5c9b2;
assign ad410a = hgrant1_p & ad4108 | !hgrant1_p & ad4109;
assign v9f769d = hgrant0_p & v9f769c | !hgrant0_p & !v9f7d42;
assign c3ce97 = hready_p & v845555 | !hready_p & c3ce96;
assign bd5864 = hbusreq0_p & bd5862 | !hbusreq0_p & !bd5863;
assign v9e9f68 = hmaster2_p & v9e9ee7 | !hmaster2_p & v9e9f67;
assign df519f = hbusreq2_p & df5187 | !hbusreq2_p & df519e;
assign c5c900 = hgrant1_p & v845542 | !hgrant1_p & !c5c8ff;
assign v9f7e01 = hbusreq2 & v9f7dff | !hbusreq2 & v9f7e00;
assign b05952 = hbusreq4_p & b05950 | !hbusreq4_p & b05951;
assign v9f781d = hbusreq4_p & v9f781b | !hbusreq4_p & v9f781c;
assign c3d6ff = hmaster0_p & c3d671 | !hmaster0_p & c3d6e9;
assign ad4744 = hgrant4_p & v845542 | !hgrant4_p & ad504b;
assign ad4779 = hbusreq4_p & ad4778 | !hbusreq4_p & !v845542;
assign ad45c7 = hmaster2_p & ad45bb | !hmaster2_p & !v845542;
assign ad4f66 = hbusreq4_p & ad4f65 | !hbusreq4_p & ad4e9b;
assign b059a2 = hgrant2_p & b0594b | !hgrant2_p & b059a1;
assign v9f7de0 = hbusreq0_p & v9f7dde | !hbusreq0_p & !v9f7ddf;
assign ad437a = hbusreq3_p & ad434b | !hbusreq3_p & !ad4379;
assign dc503e = hgrant4_p & ade581 | !hgrant4_p & ade58d;
assign b05a08 = stateG10_4_p & b05a06 | !stateG10_4_p & b05a07;
assign bd5801 = stateG10_4_p & bd57fe | !stateG10_4_p & bd5800;
assign adeab8 = hgrant3_p & adeab3 | !hgrant3_p & adeab7;
assign v9e9eb9 = hbusreq1_p & v9e9eb8 | !hbusreq1_p & v9ea4ca;
assign ad4345 = hmaster0_p & ad42d3 | !hmaster0_p & ad4344;
assign b579b1 = hgrant0_p & v845542 | !hgrant0_p & b57941;
assign b1c7d6 = hbusreq0 & b1c7d5 | !hbusreq0 & b1cfcc;
assign ad4ec1 = hbusreq0 & ad4ec0 | !hbusreq0 & ad4e7f;
assign v9ea470 = hlock0_p & v9f20a1 | !hlock0_p & v9ea46f;
assign v9ea479 = hbusreq4_p & v9ea462 | !hbusreq4_p & v9ea478;
assign b578fd = hlock4_p & b578f9 | !hlock4_p & v845542;
assign c5c8f0 = hmaster1_p & c5c8ef | !hmaster1_p & v845542;
assign ad442d = hbusreq4_p & ad442c | !hbusreq4_p & adeaa4;
assign ad4818 = hmaster0_p & ad4817 | !hmaster0_p & v845542;
assign b8f744 = hready_p & b8f743 | !hready_p & v845562;
assign ad468d = hmaster1_p & ad4689 | !hmaster1_p & ad468c;
assign dc538b = hburst0 & v8cc7d9 | !hburst0 & dc538a;
assign c3d3a8 = hgrant2_p & v845551 | !hgrant2_p & c3d3a7;
assign ade5b2 = hbusreq1 & ade5ab | !hbusreq1 & !v845558;
assign ad4eb3 = hlock0_p & ad4e54 | !hlock0_p & ad4e53;
assign df518f = hbusreq2 & df518c | !hbusreq2 & !df518e;
assign v8cc7e5 = hlock1 & v8ccb6b | !hlock1 & v8cc7e4;
assign d354ff = hmaster2_p & v845542 | !hmaster2_p & !d354fe;
assign d35720 = hmaster1_p & d3571f | !hmaster1_p & d3570b;
assign df553f = hbusreq2_p & df5537 | !hbusreq2_p & df553e;
assign d354cf = hbusreq4_p & d354ce | !hbusreq4_p & v845542;
assign ad4f01 = hgrant4_p & v84556c | !hgrant4_p & ad4f00;
assign adeab9 = hbusreq3_p & adeaad | !hbusreq3_p & adeab8;
assign df5155 = decide_p & df5154 | !decide_p & v845542;
assign b1c748 = hmaster0_p & b1c737 | !hmaster0_p & b1c747;
assign ad46ff = hgrant4_p & v845542 | !hgrant4_p & v84556c;
assign v9e9eca = decide_p & v9ea4b2 | !decide_p & v9e9ec9;
assign d35912 = hbusreq2 & d3590f | !hbusreq2 & d35911;
assign ad4363 = hmaster0_p & ad4362 | !hmaster0_p & ad42fd;
assign ad46d8 = hbusreq4_p & ad46d7 | !hbusreq4_p & v845542;
assign v9f7cf3 = hburst0_p & v9f7cf2 | !hburst0_p & !v9fa31b;
assign dc53d5 = hlock3_p & dc5390 | !hlock3_p & !v845542;
assign v9e9fe7 = jx1_p & v9e9fcd | !jx1_p & v9e9fe6;
assign ade5ae = hbusreq2 & ade583 | !hbusreq2 & v9041a4;
assign ad4323 = hbusreq1 & ad4fc1 | !hbusreq1 & v845542;
assign v9ea5ac = hgrant2_p & v9ea584 | !hgrant2_p & v9ea5ab;
assign v9ea44c = hmastlock_p & v9ea44b | !hmastlock_p & v845542;
assign b05983 = hlock4_p & b05981 | !hlock4_p & b05982;
assign v9f7ddf = hgrant0_p & v9f7da2 | !hgrant0_p & v9f7cc6;
assign c3cecb = hgrant4_p & v845542 | !hgrant4_p & c3cec2;
assign bd56d6 = hmaster2_p & v845542 | !hmaster2_p & bd56d5;
assign ad4566 = hburst0 & adea97 | !hburst0 & bd5b85;
assign d357d5 = hbusreq1_p & d357d4 | !hbusreq1_p & v84554a;
assign v9f77d6 = hbusreq1_p & v9f77d5 | !hbusreq1_p & v9f772c;
assign d35764 = hmaster1_p & d35aae | !hmaster1_p & d35763;
assign v9ea438 = hmastlock_p & v9ea437 | !hmastlock_p & v845542;
assign c5c93e = hgrant2_p & c5c8f0 | !hgrant2_p & c5c93d;
assign dc4f77 = hbusreq0 & dc4f75 | !hbusreq0 & dc4f76;
assign b1c863 = hmaster1_p & b1c85a | !hmaster1_p & b1c862;
assign v9e9eb2 = hlock3 & v9ea4cd | !hlock3 & v9e9eb1;
assign ad4583 = hmaster1_p & ad4582 | !hmaster1_p & ad457f;
assign b57a7d = hlock3 & b579e5 | !hlock3 & b57a7c;
assign d357b8 = hbusreq0 & d357b7 | !hbusreq0 & v845542;
assign adec94 = hburst1_p & v845542 | !hburst1_p & !bbbcd6;
assign v9f7e2d = stateA1_p & v845568 | !stateA1_p & c6d44d;
assign v8cc5c4 = hmaster1_p & v8cc5c2 | !hmaster1_p & v845542;
assign ad4749 = hbusreq4_p & ad505e | !hbusreq4_p & v845542;
assign c3d59f = hmaster2_p & c3d59e | !hmaster2_p & !v845542;
assign b1c5be = hbusreq1_p & b1c5b8 | !hbusreq1_p & b1c5bd;
assign d359c4 = locked_p & v84557a | !locked_p & !v845542;
assign c3d6d0 = hmaster2_p & c3d6c6 | !hmaster2_p & !c3d6cf;
assign v9f7dac = hmaster2_p & v9f7d77 | !hmaster2_p & v9f7c9f;
assign d354d2 = hgrant1_p & d354ca | !hgrant1_p & d354d1;
assign v8cc5a0 = hbusreq3 & v8cc59e | !hbusreq3 & v8cc59f;
assign ad41b8 = decide_p & ad40f0 | !decide_p & ad41b7;
assign c3cea2 = hbusreq2 & c3ce9d | !hbusreq2 & c3cea0;
assign v9f7748 = hlock4 & v9f7745 | !hlock4 & v9f7747;
assign v8ccbeb = hgrant4_p & v8ccb6a | !hgrant4_p & v845542;
assign ad4de9 = hbusreq1_p & ad4de8 | !hbusreq1_p & v845542;
assign v9f7d55 = hbusreq2_p & v9f7d52 | !hbusreq2_p & v9f7d54;
assign ad4305 = hbusreq2 & ad4304 | !hbusreq2 & !ad4282;
assign bd57c8 = hmaster2_p & bd57c4 | !hmaster2_p & ade5ce;
assign b1c7f0 = hmaster0_p & b1c7e6 | !hmaster0_p & b1c7ef;
assign c3ce49 = hbusreq1 & c3d32b | !hbusreq1 & c3d32e;
assign v8cc49a = hmaster2_p & v8cc491 | !hmaster2_p & v8cc499;
assign c3ce42 = hready_p & v845555 | !hready_p & c3ce41;
assign dc506b = hbusreq2 & dc506a | !hbusreq2 & !v845542;
assign bd5938 = hmaster1_p & bd5937 | !hmaster1_p & v84556c;
assign v9f778d = hlock3 & v9f772c | !hlock3 & v9f778c;
assign c3cea9 = decide_p & c3ce91 | !decide_p & !c3cea8;
assign d35411 = hmaster1_p & d35c06 | !hmaster1_p & d35410;
assign v9e9fa4 = hbusreq3 & v9e9fa2 | !hbusreq3 & v9e9fa3;
assign ad5037 = hgrant1_p & ad5035 | !hgrant1_p & ad5036;
assign v8cc4f9 = hbusreq0_p & v8ccbe1 | !hbusreq0_p & v845542;
assign v9e9ec6 = hmaster1_p & v9e9ec5 | !hmaster1_p & v9e9e77;
assign d35567 = hmaster1_p & d35566 | !hmaster1_p & d3549d;
assign b0591b = decide_p & b05918 | !decide_p & b058e5;
assign df5134 = hbusreq3_p & df512f | !hbusreq3_p & df5133;
assign dc4fbc = hmaster2_p & dc4fac | !hmaster2_p & !dc4fb9;
assign ad3d47 = hmaster1_p & ad3d46 | !hmaster1_p & ad43ba;
assign b1cf3c = hmaster0_p & v845542 | !hmaster0_p & b1cf3b;
assign ad4de2 = hburst0 & v845542 | !hburst0 & ade4c1;
assign ad4f5d = hbusreq1_p & ad4f5c | !hbusreq1_p & !v845542;
assign v9f76a4 = hmaster2_p & v9f76a0 | !hmaster2_p & v9f76a3;
assign v8ccb80 = hmaster2_p & v8ccb7b | !hmaster2_p & v8ccb7e;
assign b1cfcf = hmaster2_p & b1cfce | !hmaster2_p & b1cfcc;
assign adeaaf = hmaster2_p & adeaae | !hmaster2_p & !v845542;
assign c3cec6 = hmaster2_p & c3cec5 | !hmaster2_p & adeaa5;
assign bd58e4 = decide_p & bd57ee | !decide_p & !v845572;
assign ad42de = hbusreq1 & ad4e49 | !hbusreq1 & v845542;
assign v9e9f82 = hbusreq1_p & v9e9ee8 | !hbusreq1_p & v9e9f68;
assign dc4ff1 = hbusreq4_p & dc4fee | !hbusreq4_p & dc4ff0;
assign c3d5d5 = hgrant4_p & v845542 | !hgrant4_p & c3d5d4;
assign bd5748 = hbusreq2 & bd5747 | !hbusreq2 & v845542;
assign c3d69e = hmaster1_p & c3d69d | !hmaster1_p & c3d69b;
assign v9f779b = hbusreq2 & v9f7799 | !hbusreq2 & v9f779a;
assign b5794e = hgrant1_p & b5794d | !hgrant1_p & b5794a;
assign dc4fd5 = hbusreq1_p & adec89 | !hbusreq1_p & dc4fd4;
assign d359b3 = hmaster0_p & d359ac | !hmaster0_p & d359b2;
assign c3d2bb = hbusreq3 & c3d2ba | !hbusreq3 & v84554d;
assign ade5b8 = hbusreq2_p & ade5a6 | !hbusreq2_p & ade5b7;
assign v9f7cf4 = stateA1_p & v845542 | !stateA1_p & !v9f7cf3;
assign adea94 = hbusreq4_p & adea93 | !hbusreq4_p & !v845542;
assign v9e9ed3 = hmaster1_p & v9e9eba | !hmaster1_p & v9e9ead;
assign ad4258 = hmaster0_p & ad4257 | !hmaster0_p & ad4167;
assign c3d2c0 = hmaster1_p & c3d2b9 | !hmaster1_p & c3d2bf;
assign b059aa = hmaster0_p & b05968 | !hmaster0_p & b059a9;
assign ad4f7b = hmaster2_p & ad4f78 | !hmaster2_p & ad4f7a;
assign b57416 = hbusreq2 & b57414 | !hbusreq2 & b57415;
assign ad46a7 = hlock0_p & ad46a6 | !hlock0_p & ad46a5;
assign v8cc120 = decide_p & v8ccbd7 | !decide_p & v8cc11f;
assign dc53c8 = hready_p & v845542 | !hready_p & dc53c7;
assign d35a26 = hmaster1_p & d35a20 | !hmaster1_p & d35a25;
assign bd5874 = hbusreq0_p & bd5872 | !hbusreq0_p & bd5873;
assign b05901 = hbusreq2 & b058ff | !hbusreq2 & b05900;
assign df516f = hbusreq2 & df5141 | !hbusreq2 & df5142;
assign ad4743 = hmaster2_p & v845542 | !hmaster2_p & ad4742;
assign d359fd = hmaster2_p & d359f4 | !hmaster2_p & d359fc;
assign d35c02 = hlock4_p & d359c4 | !hlock4_p & v845542;
assign b5742c = hmaster1_p & b5794b | !hmaster1_p & b5742b;
assign bd5778 = hbusreq2 & bd5777 | !hbusreq2 & v845542;
assign dc53b8 = hbusreq1_p & dc5389 | !hbusreq1_p & v84556c;
assign c3d398 = hgrant2_p & v845551 | !hgrant2_p & c3d397;
assign ad4df0 = hready & v9c81a4 | !hready & ad4def;
assign c3d482 = hmaster1_p & c3d47f | !hmaster1_p & c3d481;
assign ad438c = hbusreq3 & ad4385 | !hbusreq3 & ad438b;
assign v9e9ea6 = hgrant1_p & v9ea4bc | !hgrant1_p & v9e9ea5;
assign ad4ff8 = hmaster1_p & ad4ff7 | !hmaster1_p & ad4fee;
assign b1cfc0 = hgrant0_p & bd5b81 | !hgrant0_p & !v845542;
assign v8cc0c5 = hbusreq0 & v8cc0c4 | !hbusreq0 & v8ccbd8;
assign c3d75f = hbusreq2_p & c3d75a | !hbusreq2_p & c3d75e;
assign d3580c = hlock0_p & v845542 | !hlock0_p & d3580b;
assign c3d2e1 = hmaster1_p & c3d2dc | !hmaster1_p & c3d2e0;
assign v9f7847 = hmaster1_p & v9f7829 | !hmaster1_p & v9f7846;
assign v8cc47d = hbusreq0 & v8cc47b | !hbusreq0 & v8cc47c;
assign d359ae = hbusreq1 & d359ad | !hbusreq1 & !v845542;
assign b05970 = hbusreq1_p & b0595b | !hbusreq1_p & b0596b;
assign c3d348 = hgrant1_p & v84554d | !hgrant1_p & c3d347;
assign c3d2d0 = hbusreq3 & c3d2cf | !hbusreq3 & v84554d;
assign b573fe = hmaster0_p & b573fd | !hmaster0_p & v845542;
assign d35bf0 = hlock4_p & d35983 | !hlock4_p & v84556c;
assign hmastlock = cc370b;
assign d35519 = hbusreq0 & d35433 | !hbusreq0 & d35518;
assign dc531a = hmaster2_p & v845542 | !hmaster2_p & dc5319;
assign v9f7dbd = hgrant1_p & v9f7dab | !hgrant1_p & v9f7dbc;
assign d357a5 = hbusreq4 & d3579f | !hbusreq4 & d357a4;
assign v9e9f90 = stateG10_4_p & v9e9f8a | !stateG10_4_p & v9e9f8f;
assign v9e9f8a = hlock0_p & v9e9f89 | !hlock0_p & v9ea464;
assign v8cc78d = hready_p & v8cc4e0 | !hready_p & v8cc78b;
assign b1c569 = hgrant1_p & b1d01a | !hgrant1_p & b1c568;
assign v8cc7cd = hlock2 & v8ccbf6 | !hlock2 & v8cc7cc;
assign b1c70e = hbusreq0_p & v84556c | !hbusreq0_p & v845542;
assign dc4fe5 = stateG10_4_p & ade553 | !stateG10_4_p & dc4fe4;
assign ade5a5 = hmaster1_p & ade569 | !hmaster1_p & ade5a4;
assign bd58ce = hbusreq4_p & bd58cd | !hbusreq4_p & bd58aa;
assign d35647 = hlock1_p & d35646 | !hlock1_p & !v845542;
assign ad4f4b = hmaster2_p & ad4f48 | !hmaster2_p & ad4f4a;
assign ad4f0a = hbusreq4_p & ad4f09 | !hbusreq4_p & ad4ef7;
assign v8cc796 = locked_p & v8cc793 | !locked_p & v845542;
assign ad45e2 = hlock0_p & ad45ae | !hlock0_p & !v845542;
assign v9e9f93 = hbusreq0 & v9e9f92 | !hbusreq0 & v9e9f8e;
assign ad413a = hgrant4_p & adea99 | !hgrant4_p & ad4e98;
assign ad4da3 = hbusreq1_p & ad4da2 | !hbusreq1_p & ad4da1;
assign b57a2f = hmaster0_p & b579c5 | !hmaster0_p & b579e5;
assign d359ca = hmaster2_p & v84557a | !hmaster2_p & !d359c9;
assign ad4e81 = hbusreq4 & ad4e7b | !hbusreq4 & ad4e80;
assign df5141 = hbusreq1_p & df5140 | !hbusreq1_p & v845542;
assign b1c6fc = hgrant2_p & b1d01a | !hgrant2_p & b1c6fb;
assign adeab0 = hmaster0_p & v845542 | !hmaster0_p & !adeaaf;
assign v9f76c1 = hmaster1_p & v9f76c0 | !hmaster1_p & v9f7d47;
assign df513c = hmaster2_p & v84556c | !hmaster2_p & df513b;
assign v9f77b4 = hlock2 & v9f779f | !hlock2 & v9f77b3;
assign ad4f85 = hmaster2_p & ad4f7f | !hmaster2_p & ad4f84;
assign c5c976 = hgrant1_p & c5c975 | !hgrant1_p & c5c972;
assign d354f7 = hbusreq4_p & d35c07 | !hbusreq4_p & !v845542;
assign c5c8f6 = hlock1_p & c5c88f | !hlock1_p & v845542;
assign d359f1 = hlock4_p & d359f0 | !hlock4_p & v845542;
assign v9f7d04 = hmaster2_p & v9f7c9b | !hmaster2_p & v9f7c9f;
assign c3d36b = hmaster0_p & c3d2de | !hmaster0_p & !c3d2be;
assign d356ec = hmaster1_p & d356eb | !hmaster1_p & d356e5;
assign v9e9fbf = hready_p & v9ea4a4 | !hready_p & v9e9fbe;
assign v9f7780 = hlock2_p & v9f777e | !hlock2_p & v9f777f;
assign v8ccb72 = hlock3_p & v8ccb6e | !hlock3_p & v845542;
assign v9f7d64 = hmaster0_p & v9f7d5f | !hmaster0_p & !v9f7d63;
assign v9f7d3d = hlock1_p & v9f7d3b | !hlock1_p & v9f7d3c;
assign ad4d90 = stateA1_p & v9ea412 | !stateA1_p & ad4d8f;
assign bd58f3 = hbusreq2_p & bd58f2 | !hbusreq2_p & v845542;
assign ad47fc = hgrant2_p & ad47f9 | !hgrant2_p & ad47fb;
assign v9f77cc = hbusreq4 & v9f77ca | !hbusreq4 & v9f77cb;
assign v9f7e40 = hlock0 & v9f7e3f | !hlock0 & v9f7e3b;
assign v9f7da9 = hlock1 & v9f7da3 | !hlock1 & v9f7da8;
assign c3d2e8 = hburst0 & c3d2e6 | !hburst0 & c3d2e7;
assign bd58cb = hmaster2_p & bd58c4 | !hmaster2_p & bd58ca;
assign d3570d = hgrant2_p & d356fd | !hgrant2_p & d3570c;
assign ad470b = hmaster2_p & adec93 | !hmaster2_p & !ad470a;
assign ad43cc = hbusreq0 & ad43cb | !hbusreq0 & !v845542;
assign d359e0 = hbusreq0 & d359df | !hbusreq0 & v845542;
assign dc53a3 = hmaster2_p & v845542 | !hmaster2_p & !v845566;
assign ad4730 = hgrant1_p & ad460b | !hgrant1_p & ad472f;
assign b579de = hlock4 & b579d5 | !hlock4 & b579dd;
assign bd5ea2 = hbusreq4 & bd5e9f | !hbusreq4 & bd5ea1;
assign ad4275 = hbusreq1_p & ad4e64 | !hbusreq1_p & v845542;
assign v9f7798 = hlock3 & v9f772d | !hlock3 & v9f7797;
assign v8cc7ee = hbusreq2 & v8cc7ea | !hbusreq2 & v8cc7eb;
assign b05990 = stateG10_4_p & b0598e | !stateG10_4_p & !b0598f;
assign ad430f = hgrant2_p & ad4307 | !hgrant2_p & !ad430e;
assign ad3d1c = hmaster1_p & ad3d1b | !hmaster1_p & ad3d12;
assign v9ea5da = hmaster1_p & v9ea5d9 | !hmaster1_p & v9ea579;
assign v9ea428 = hmaster0_p & v845542 | !hmaster0_p & v9ea415;
assign b1c0b0 = hready_p & b1c0ac | !hready_p & b1c868;
assign ad3cef = hmaster2_p & ad3ccc | !hmaster2_p & ad3cee;
assign v8cc7c2 = hbusreq0 & v8cc7c0 | !hbusreq0 & v8cc7c1;
assign d35a9f = hmaster0_p & d35a9a | !hmaster0_p & d35a9e;
assign ad3d52 = hmaster1_p & ad3d51 | !hmaster1_p & ad3d12;
assign ad443c = hready & ad4429 | !hready & ad443b;
assign v9f7df5 = hlock2 & v9f7df2 | !hlock2 & v9f7df4;
assign e0edf9 = stateG2_p & v845542 | !stateG2_p & c74a04;
assign c3d580 = hbusreq1_p & c3d4f7 | !hbusreq1_p & c3d57f;
assign v8cc59f = hlock3 & v8cc489 | !hlock3 & v8cc59e;
assign ad472d = hmaster1_p & ad472c | !hmaster1_p & ad460e;
assign b05979 = hgrant4_p & b058e7 | !hgrant4_p & b05954;
assign b1c841 = hmaster2_p & b1c840 | !hmaster2_p & d35a9c;
assign v84555e = hburst1_p & v845542 | !hburst1_p & !v845542;
assign d35432 = hbusreq4_p & d35431 | !hbusreq4_p & v845542;
assign bd5837 = hburst0 & c3d673 | !hburst0 & bd5836;
assign v9f76d2 = hready_p & v9f76bd | !hready_p & !v9f76d1;
assign v9f76ad = hmaster1_p & v9f76ac | !hmaster1_p & v9f76a6;
assign b1c588 = hgrant3_p & b1c50e | !hgrant3_p & b1c587;
assign c3d68d = hmaster0_p & c3d682 | !hmaster0_p & c3d685;
assign d357cb = hbusreq4_p & d357c9 | !hbusreq4_p & d357ca;
assign bd5819 = hgrant4_p & v84556c | !hgrant4_p & bd5806;
assign ade629 = hbusreq3_p & ade5bc | !hbusreq3_p & ade628;
assign ad441e = decide_p & ad440a | !decide_p & ad441d;
assign df512c = decide_p & df512b | !decide_p & d6ebca;
assign b578fc = hbusreq1_p & b578fb | !hbusreq1_p & b578fa;
assign c3d6ae = hgrant4_p & c3d66d | !hgrant4_p & !c3d6ac;
assign c3cec8 = hgrant4_p & v845542 | !hgrant4_p & !c3cebc;
assign d35917 = hbusreq3 & d35916 | !hbusreq3 & v845542;
assign d354de = hlock2_p & d354d5 | !hlock2_p & !d354dd;
assign b57a32 = decide_p & b57a21 | !decide_p & b57a31;
assign d35716 = hlock2_p & d3570d | !hlock2_p & !d35715;
assign v9f7755 = hbusreq4 & v9f7753 | !hbusreq4 & v9f7754;
assign df51c0 = hbusreq2 & df51ac | !hbusreq2 & !v84554c;
assign ad46a8 = hgrant4_p & v845542 | !hgrant4_p & ad46a7;
assign c3d6ee = hmaster2_p & c3d6e3 | !hmaster2_p & c3d6ed;
assign ad43ff = hmaster0_p & ad43d4 | !hmaster0_p & ad43fe;
assign c3d73f = hbusreq0_p & c3d669 | !hbusreq0_p & c3d73e;
assign c3d689 = hlock0_p & c3d66d | !hlock0_p & c3d688;
assign ad4581 = hbusreq3 & ad4576 | !hbusreq3 & v845542;
assign b059db = hgrant4_p & b058d0 | !hgrant4_p & !b059da;
assign b1c735 = hmaster2_p & v845542 | !hmaster2_p & b1c734;
assign ad41a7 = hmaster0_p & ad41a5 | !hmaster0_p & ad41a6;
assign b058e6 = stateA1_p & v845542 | !stateA1_p & v9fa31b;
assign c3d693 = hmaster0_p & c3d683 | !hmaster0_p & c3d685;
assign b579dd = hbusreq0 & b579db | !hbusreq0 & b579dc;
assign ad436a = hgrant2_p & ad4368 | !hgrant2_p & !ad4369;
assign ad4eec = hgrant4_p & v845542 | !hgrant4_p & ad4eda;
assign bd5ea9 = decide_p & bd5ea8 | !decide_p & v845572;
assign v8ccbd8 = hmaster2_p & v845542 | !hmaster2_p & v8d2b2b;
assign b05982 = hgrant4_p & v9f7d42 | !hgrant4_p & !b05980;
assign bd58a2 = locked_p & bd58a1 | !locked_p & v845542;
assign b1cf41 = hbusreq3 & b1cf40 | !hbusreq3 & b1cf2c;
assign b574ce = hbusreq2 & b574cc | !hbusreq2 & b574cd;
assign stateG10_2 = !ba05d0;
assign b059b4 = hlock4 & b0595b | !hlock4 & b059b3;
assign ad4364 = hmaster1_p & ad4363 | !hmaster1_p & ad4300;
assign b1c04d = hbusreq2 & b1c722 | !hbusreq2 & b1c71d;
assign v9f780b = hlock0_p & v9f77eb | !hlock0_p & v9f780a;
assign df54db = hmaster1_p & v845542 | !hmaster1_p & df54da;
assign b0589e = jx1_p & v85746e | !jx1_p & !v845542;
assign bd58fc = hmaster1_p & bd58fb | !hmaster1_p & bd5898;
assign b1c7a3 = hbusreq0 & b1c7a2 | !hbusreq0 & b1cfcc;
assign v8ccbe8 = hgrant1_p & v8ccbe7 | !hgrant1_p & v8ccbe3;
assign d35bf6 = hbusreq4_p & d35bf5 | !hbusreq4_p & v845542;
assign ad4edb = hgrant4_p & ad4e5c | !hgrant4_p & ad4eda;
assign v9e9e6c = hgrant2_p & v9e9e68 | !hgrant2_p & v9e9e6b;
assign v9f7695 = hgrant4_p & v9f7d5d | !hgrant4_p & v9f7694;
assign b1c6ce = hready_p & b1c6cc | !hready_p & b1c6cd;
assign d35a5a = hlock4_p & d35a59 | !hlock4_p & !dc500f;
assign ad447a = stateG10_4_p & c3cec2 | !stateG10_4_p & ad4479;
assign ad4ed1 = hbusreq1_p & ad4eca | !hbusreq1_p & ad4ed0;
assign bd58ac = hmaster2_p & bd58a9 | !hmaster2_p & bd58ab;
assign ad4339 = hbusreq1_p & ad4338 | !hbusreq1_p & c3d2d9;
assign ad501c = hbusreq3 & ad501b | !hbusreq3 & v845547;
assign bd5890 = hgrant4_p & v845542 | !hgrant4_p & !bd5875;
assign ad4269 = hbusreq1_p & ad4268 | !hbusreq1_p & v845542;
assign b058ed = hlock4 & b058ea | !hlock4 & b058ec;
assign ad40e8 = hmaster1_p & ad48b4 | !hmaster1_p & ad40e7;
assign b05966 = hbusreq3 & b05963 | !hbusreq3 & b05965;
assign b1c741 = hbusreq4_p & c3d66d | !hbusreq4_p & !b1c73c;
assign c3d32f = hgrant1_p & v84554d | !hgrant1_p & c3d32e;
assign v8cc815 = hgrant2_p & v8cc813 | !hgrant2_p & v8cc80a;
assign v8cc129 = hmaster1_p & v8cc128 | !hmaster1_p & v845542;
assign c3ce2a = hmaster1_p & c3d3a5 | !hmaster1_p & c3ce29;
assign v9f786f = hlock2 & v9f786c | !hlock2 & v9f786e;
assign ad4f26 = hbusreq2 & ad4eb0 | !hbusreq2 & !ad4f1a;
assign v9f772f = hmastlock_p & v84557a | !hmastlock_p & !v845542;
assign ade570 = hburst1 & v845542 | !hburst1 & !c3d673;
assign v8cc48d = hbusreq2 & v8cc48a | !hbusreq2 & v8cc48c;
assign d3561f = hbusreq1_p & d35618 | !hbusreq1_p & d3561e;
assign dc53c3 = hmaster1_p & dc53c2 | !hmaster1_p & v845542;
assign dc4ff3 = hgrant4_p & v84556c | !hgrant4_p & ade557;
assign dc4fbe = hbusreq4 & dc4fbb | !hbusreq4 & dc4fbd;
assign df5079 = hlock1_p & df5078 | !hlock1_p & v845542;
assign cc36ef = decide_p & cc36ba | !decide_p & !v84556c;
assign c5c97a = hmaster2_p & c5c968 | !hmaster2_p & !c5c92f;
assign v9f7676 = hmaster1_p & v9f7e2c | !hmaster1_p & v9f7675;
assign ad4737 = hbusreq4_p & ad502f | !hbusreq4_p & !v845542;
assign b574b2 = hlock0_p & b579ba | !hlock0_p & b574b1;
assign bd584c = hbusreq4_p & bd5849 | !hbusreq4_p & bd584b;
assign d35808 = hgrant4_p & v84554a | !hgrant4_p & d35807;
assign b058b7 = hmaster2_p & b058a3 | !hmaster2_p & b058b6;
assign c3ce4c = hbusreq1_p & c3ce4b | !hbusreq1_p & c3d305;
assign c5c88e = locked_p & c5c88d | !locked_p & !v845542;
assign d35956 = hlock0_p & d35955 | !hlock0_p & v845542;
assign b57abc = hbusreq3_p & b57a8f | !hbusreq3_p & b57abb;
assign ade5d6 = hbusreq4_p & ade5d5 | !hbusreq4_p & !v845542;
assign ad4570 = hready & ad456e | !hready & ad456f;
assign ad13e5 = hgrant3_p & ad13e1 | !hgrant3_p & ad13e4;
assign ad4824 = hbusreq2 & ad4fb6 | !hbusreq2 & v845542;
assign b059d8 = hgrant0_p & b059c2 | !hgrant0_p & v9f7d42;
assign ad4694 = hbusreq4_p & ad4e7e | !hbusreq4_p & v845542;
assign bd57a2 = hbusreq2 & bd57a1 | !hbusreq2 & v845542;
assign c3ceea = hmaster1_p & c3cee7 | !hmaster1_p & c3cee9;
assign c3d2fb = hmaster2_p & v8da5a1 | !hmaster2_p & adeaa5;
assign d357be = hmaster1_p & d357bd | !hmaster1_p & d3577c;
assign b574d2 = hbusreq1 & b574b7 | !hbusreq1 & b574b8;
assign dc4fdb = hbusreq2 & dc4fda | !hbusreq2 & dc4f61;
assign b573d7 = hbusreq1 & b579e1 | !hbusreq1 & b579ce;
assign d35424 = hmaster2_p & d35419 | !hmaster2_p & d35423;
assign d354f5 = hbusreq1_p & v84555a | !hbusreq1_p & d35a9b;
assign ad46ad = hbusreq4 & ad46a0 | !hbusreq4 & ad46ac;
assign b574c2 = hbusreq4_p & b579c9 | !hbusreq4_p & b574c1;
assign b1c5f2 = hlock2_p & b1c5e3 | !hlock2_p & b1c5f1;
assign dc4fce = hmaster2_p & adec89 | !hmaster2_p & adec90;
assign c5c96d = hmaster1_p & c5c96b | !hmaster1_p & c5c96c;
assign d35c0a = hbusreq3 & d35c09 | !hbusreq3 & !v84555a;
assign v9f777f = hmaster1_p & v9f7772 | !hmaster1_p & v9f776d;
assign df51c4 = hgrant1_p & df553a | !hgrant1_p & !df517e;
assign b574fe = hbusreq3 & b574d3 | !hbusreq3 & b57942;
assign v8cc621 = hbusreq2 & v8cc620 | !hbusreq2 & v8cc4ad;
assign c3d39f = hgrant4_p & v845542 | !hgrant4_p & !c3d399;
assign b1c074 = hbusreq4 & b1c06b | !hbusreq4 & b1c073;
assign v9e9fce = decide_p & v9ea3f4 | !decide_p & v9ea409;
assign ad4fad = hmastlock_p & ad4fac | !hmastlock_p & v845542;
assign v9f7ce8 = hbusreq2 & v9f7ce6 | !hbusreq2 & v9f7ce7;
assign v9e9f4c = locked_p & v9f20a1 | !locked_p & v9ea3e6;
assign ad45df = hbusreq4_p & ad4daa | !hbusreq4_p & v845542;
assign dc4ff8 = hbusreq0 & dc4ff2 | !hbusreq0 & dc4ff7;
assign b0592f = hmaster1_p & b0592e | !hmaster1_p & b05926;
assign v9ea56d = hmaster0_p & v9f20a1 | !hmaster0_p & v9ea567;
assign bd5820 = hbusreq4_p & bd581d | !hbusreq4_p & bd581f;
assign b57aeb = hbusreq2_p & b57aea | !hbusreq2_p & b57a31;
assign c6d44d = start_p & v845542 | !start_p & !v857440;
assign dc502b = hmaster2_p & dc4ff1 | !hmaster2_p & dc502a;
assign ad43c9 = hbusreq0_p & ad45ae | !hbusreq0_p & v845542;
assign v9f775a = hmaster2_p & v9f772a | !hmaster2_p & v9f772f;
assign dc4f8d = hmaster2_p & dc4f74 | !hmaster2_p & !ade5d5;
assign b1c7a8 = hgrant4_p & b1c714 | !hgrant4_p & !b1c79d;
assign dc505e = hgrant4_p & v84556c | !hgrant4_p & ade59c;
assign v9f7d8e = stateG10_4_p & v9f7d8a | !stateG10_4_p & v9f7d8c;
assign df51a9 = hmaster0_p & df51a7 | !hmaster0_p & df51a8;
assign ad419f = hmaster0_p & ad419e | !hmaster0_p & v845542;
assign df50d6 = hbusreq4_p & df54e1 | !hbusreq4_p & !v845542;
assign d3543d = hbusreq2_p & d3543c | !hbusreq2_p & d3543b;
assign ad4285 = hmaster0_p & ad4283 | !hmaster0_p & ad4284;
assign c5c3b5 = decide_p & c5c8e1 | !decide_p & c5c9b2;
assign dc4fa4 = hbusreq1_p & dc4fa2 | !hbusreq1_p & dc4fa3;
assign ad4e79 = hbusreq4_p & ad4e76 | !hbusreq4_p & ad4e78;
assign adea87 = stateA1_p & adea86 | !stateA1_p & !adea85;
assign d354a2 = hbusreq1_p & d354a1 | !hbusreq1_p & !d354a0;
assign v8cc504 = hgrant2_p & v845542 | !hgrant2_p & v8cc503;
assign ad4f9c = hgrant1_p & ad4f63 | !hgrant1_p & ad4f9b;
assign ad4dae = hmaster2_p & ad4dac | !hmaster2_p & ad4dad;
assign bd5b8b = hbusreq2 & bd5b83 | !hbusreq2 & bd5b8a;
assign ad43f3 = hbusreq4_p & ad43ca | !hbusreq4_p & !v845542;
assign c3d510 = hmaster2_p & c3d50f | !hmaster2_p & !v845542;
assign c3d6e9 = hmaster2_p & c3d66a | !hmaster2_p & c3d674;
assign adec9b = hbusreq4_p & adec9a | !hbusreq4_p & v845542;
assign v8cc5a5 = hbusreq2 & v8cc5a0 | !hbusreq2 & v8cc5a4;
assign d35747 = hlock2_p & d35742 | !hlock2_p & !d35746;
assign d354fc = hbusreq1_p & d35c01 | !hbusreq1_p & d354f8;
assign ad4f8f = hgrant4_p & ad4f3e | !hgrant4_p & ad4e98;
assign b05a1d = hbusreq4_p & b05a1b | !hbusreq4_p & b05a1c;
assign ad3ce3 = hmaster2_p & v845542 | !hmaster2_p & ad3ce2;
assign b1cf48 = decide_p & b1cf47 | !decide_p & v845542;
assign ad3d33 = hbusreq2 & ad4393 | !hbusreq2 & v845542;
assign ad426b = hready & ad4e4b | !hready & ad426a;
assign bd582e = hbusreq0 & bd582c | !hbusreq0 & bd582d;
assign v9f7666 = hbusreq4_p & v9f7664 | !hbusreq4_p & v9f7665;
assign dc5089 = hbusreq3_p & dc5087 | !hbusreq3_p & !dc5088;
assign ad4146 = hbusreq2 & ad4145 | !hbusreq2 & v845542;
assign v882b8e = hmaster1_p & v91784a | !hmaster1_p & v845542;
assign d355ad = hlock2_p & v845542 | !hlock2_p & d355ac;
assign ad4f77 = hmaster2_p & ad4f74 | !hmaster2_p & ad4f76;
assign v9ea48a = hmaster0_p & v9ea461 | !hmaster0_p & v9ea489;
assign ad430c = hgrant1_p & v845542 | !hgrant1_p & ad430b;
assign ad480b = hbusreq2 & ad480a | !hbusreq2 & v845542;
assign b1c757 = hmaster2_p & b1c755 | !hmaster2_p & !b1c756;
assign ad4705 = hready & ad4702 | !hready & ad4704;
assign v8cc80f = hlock2 & v8ccb6b | !hlock2 & v8cc80d;
assign ad43c2 = stateG2_p & v845542 | !stateG2_p & ad43c1;
assign df5148 = hbusreq1_p & df5147 | !hbusreq1_p & v845542;
assign d35573 = hbusreq2 & d354fc | !hbusreq2 & !d354f5;
assign v9f76b6 = hmaster1_p & v9f76b5 | !hmaster1_p & v9f7d2f;
assign v8cc498 = hlock0_p & v8cc492 | !hlock0_p & v8cc497;
assign bd58a5 = hlock0_p & bd58a3 | !hlock0_p & !bd58a4;
assign c3d5a2 = hready & c3d5a1 | !hready & !v845564;
assign v9ea434 = hmaster1_p & v9ea410 | !hmaster1_p & v9ea433;
assign d354c4 = hbusreq4 & d354c3 | !hbusreq4 & d354b6;
assign bd5b70 = hbusreq3 & bd5b6f | !hbusreq3 & v845564;
assign ad43f1 = hmaster2_p & ad43f0 | !hmaster2_p & v845542;
assign v9f77ea = hbusreq4_p & v9f77e7 | !hbusreq4_p & !v9f77e9;
assign ad4f30 = hmaster1_p & ad4f2f | !hmaster1_p & ad4f16;
assign b1c730 = hbusreq2_p & b1c72c | !hbusreq2_p & b1c72f;
assign df54f4 = hgrant1_p & df54f3 | !hgrant1_p & !v845542;
assign dc53de = jx1_p & dc53dd | !jx1_p & dc53d1;
assign dc539c = hburst1_p & v8f2540 | !hburst1_p & v857b36;
assign v9f7d2a = hbusreq1 & v9f7d28 | !hbusreq1 & !v9f7d29;
assign b1d019 = hgrant3_p & b1cf49 | !hgrant3_p & b1d018;
assign c3ce01 = hgrant2_p & v845551 | !hgrant2_p & c3ce00;
assign ad4fdd = hgrant4_p & v84556c | !hgrant4_p & ad4fdc;
assign b1c75f = hmaster0_p & b1c75d | !hmaster0_p & b1c75e;
assign ad455b = hburst0 & adec8c | !hburst0 & adec8d;
assign v9ea4e6 = hbusreq3_p & v9ea4a1 | !hbusreq3_p & v9ea4e5;
assign bd5784 = hmastlock_p & bd5783 | !hmastlock_p & c3d668;
assign cc36e8 = hgrant1_p & cc36bd | !hgrant1_p & !cc36e7;
assign d3549a = hmaster0_p & d35492 | !hmaster0_p & d35499;
assign b1cfc7 = hmaster2_p & b1cfbf | !hmaster2_p & b1cfc6;
assign c3d5ee = hmaster2_p & c3d5dc | !hmaster2_p & adeaa5;
assign b57442 = hready_p & b57436 | !hready_p & b57441;
assign ad4461 = hgrant4_p & ad4460 | !hgrant4_p & v845542;
assign v9f7d17 = hready & v9f7d16 | !hready & v9f7d12;
assign v9f7ded = hlock1 & v9f7de7 | !hlock1 & v9f7dec;
assign ad46ac = hbusreq0 & ad46a3 | !hbusreq0 & ad46ab;
assign c3ce18 = hmaster0_p & c3ce17 | !hmaster0_p & !c3d2be;
assign b1caf9 = hbusreq4 & b1caee | !hbusreq4 & b1caf8;
assign ad45c8 = hbusreq4 & v845542 | !hbusreq4 & !ad45c7;
assign v9ea403 = hlock0_p & v9ea3fb | !hlock0_p & v9ea402;
assign v9ea3ff = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea3fe;
assign b1c6be = hgrant2_p & v845542 | !hgrant2_p & b1c6bd;
assign v8cc4a9 = hready & v8cc4a8 | !hready & v8cc494;
assign v9f77c9 = hlock0 & v9f77c8 | !hlock0 & v9f77c2;
assign v9f7d6a = hready_p & v9f7d39 | !hready_p & !v9f7d69;
assign bd575d = locked_p & dc5036 | !locked_p & !v845542;
assign ade65e = decide_p & ade65d | !decide_p & adeaa7;
assign c3d6db = hbusreq1_p & c3d676 | !hbusreq1_p & !c3d685;
assign ad4416 = hmaster2_p & ad4415 | !hmaster2_p & v845542;
assign df50de = hready_p & v845542 | !hready_p & df50dd;
assign ad47f1 = hgrant2_p & ad47f0 | !hgrant2_p & !ad47ec;
assign dc5025 = hmaster2_p & dc4feb | !hmaster2_p & dc5024;
assign b57407 = hmastlock_p & b57406 | !hmastlock_p & v845542;
assign b05a55 = hlock2_p & b05a51 | !hlock2_p & b05a54;
assign v8cc7d2 = hgrant2_p & v8cc7ad | !hgrant2_p & v8cc7d0;
assign c3d35d = hgrant1_p & v84554d | !hgrant1_p & c3d313;
assign v9f77de = hbusreq1 & v9f77dc | !hbusreq1 & v9f77dd;
assign dc4fa1 = hmaster0_p & dc4f9a | !hmaster0_p & dc4fa0;
assign ad4719 = hready & ad4714 | !hready & ad4718;
assign bd58c6 = hlock0_p & bd58c5 | !hlock0_p & !ade562;
assign b57a84 = hbusreq1 & b57a6b | !hbusreq1 & b57a6c;
assign bd58eb = hlock2_p & bd58ea | !hlock2_p & !v845542;
assign ad4326 = hmaster0_p & ad4315 | !hmaster0_p & ad4325;
assign ad4d8e = hburst0_p & v9ea411 | !hburst0_p & !v84557e;
assign b1c791 = hmaster1_p & b1c78d | !hmaster1_p & b1c790;
assign ade63d = decide_p & ade63c | !decide_p & v845542;
assign cc36f7 = hgrant1_p & df54f3 | !hgrant1_p & cc36f6;
assign bd5735 = locked_p & bd5733 | !locked_p & c3d66d;
assign v9e9ec7 = hmaster0_p & v9e9ec4 | !hmaster0_p & v9e9e79;
assign ac1451 = hmaster1_p & ac1450 | !hmaster1_p & v845542;
assign b058a7 = locked_p & b058a6 | !locked_p & !v9f7d42;
assign ad4472 = hgrant1_p & ad4471 | !hgrant1_p & ad443c;
assign v9ea411 = start_p & v845542 | !start_p & !v84557e;
assign ad4424 = hbusreq2 & ad4399 | !hbusreq2 & v845542;
assign ad4803 = decide_p & ad4605 | !decide_p & ad4754;
assign v9f7d52 = hlock2_p & v9f7d50 | !hlock2_p & v9f7d51;
assign ade4ba = hburst0_p & c74a04 | !hburst0_p & !v8f96d9;
assign ade4d8 = hburst1 & v845542 | !hburst1 & !ade4d7;
assign v9ea59a = hbusreq4_p & v9ea46a | !hbusreq4_p & v9ea4d7;
assign v9f78a6 = hmaster1_p & v9f78a5 | !hmaster1_p & v9f7846;
assign bd58b7 = hbusreq1_p & bd58b6 | !hbusreq1_p & !v845542;
assign bd5898 = hmaster0_p & bd5857 | !hmaster0_p & bd5897;
assign df54e0 = hburst1 & df54dd | !hburst1 & df54df;
assign ad4435 = hlock1_p & ad4434 | !hlock1_p & v845547;
assign ade558 = hlock4_p & ade554 | !hlock4_p & !ade557;
assign ad3cdb = hbusreq2 & ad3cd0 | !hbusreq2 & ad3cd9;
assign v9ea5b0 = hlock2 & v9ea586 | !hlock2 & v9ea5af;
assign b574bc = hlock3 & b579c5 | !hlock3 & b574bb;
assign v8cc806 = hbusreq3 & v8cc803 | !hbusreq3 & v8cc805;
assign ad41ab = hbusreq2_p & ad41a9 | !hbusreq2_p & ad48c7;
assign v9f7c95 = hburst0_p & v9ea3e4 | !hburst0_p & !v845582;
assign v9e9e78 = hmaster1_p & v9ea3fd | !hmaster1_p & v9e9e77;
assign d35765 = hgrant2_p & v845542 | !hgrant2_p & !d35764;
assign b57439 = hgrant1_p & v845542 | !hgrant1_p & b579da;
assign v8cc800 = hready & v8cc7ff | !hready & v8cc439;
assign ad45b0 = hbusreq4_p & ad45af | !hbusreq4_p & v845542;
assign ad46f1 = hmaster0_p & ad46e7 | !hmaster0_p & ad46f0;
assign b1c86a = hgrant3_p & b1c84f | !hgrant3_p & b1c869;
assign d359bb = hmastlock_p & d359b9 | !hmastlock_p & !d359ba;
assign b1c864 = hgrant2_p & b1d01a | !hgrant2_p & b1c863;
assign ade4c6 = hbusreq4_p & ade4c5 | !hbusreq4_p & v845542;
assign d35410 = hmaster0_p & d35c0a | !hmaster0_p & !d3540f;
assign ad42b4 = hbusreq4_p & ad4de2 | !hbusreq4_p & !v845542;
assign ade4d9 = hburst0 & v845542 | !hburst0 & ade4d8;
assign dc5394 = hmaster2_p & v845542 | !hmaster2_p & !adea88;
assign ad4f11 = hbusreq0 & ad4f0b | !hbusreq0 & ad4f10;
assign c3d5db = stateG10_4_p & c3d5d9 | !stateG10_4_p & !c3d5da;
assign v8cc7d0 = hmaster1_p & v8ccbe5 | !hmaster1_p & v8cc7cf;
assign c3cecf = hbusreq4 & c3cec7 | !hbusreq4 & !c3cece;
assign b05a5a = locked_p & b05a59 | !locked_p & b058a3;
assign bd5923 = hbusreq0_p & d35617 | !hbusreq0_p & dc5318;
assign b059bc = hlock2 & b05964 | !hlock2 & b059bb;
assign b57a89 = hmaster0_p & v845542 | !hmaster0_p & b57a88;
assign bd5810 = stateG10_4_p & bd580d | !stateG10_4_p & bd580f;
assign bd5783 = stateA1_p & v845542 | !stateA1_p & bd5782;
assign ad4e70 = hgrant4_p & d3597f | !hgrant4_p & ad4e6f;
assign bd574a = hbusreq3 & bd5749 | !hbusreq3 & dc4fcb;
assign b1c79c = hgrant0_p & v84556c | !hgrant0_p & !adec89;
assign bd586b = hgrant4_p & bd5735 | !hgrant4_p & bd580d;
assign c3d51a = hmaster0_p & c3d518 | !hmaster0_p & c3d519;
assign v8cc791 = hbusreq3_p & v8cc785 | !hbusreq3_p & v8cc790;
assign d3559e = hbusreq2_p & d35441 | !hbusreq2_p & d3559d;
assign ad4712 = hbusreq4_p & ad4711 | !hbusreq4_p & v845542;
assign v9f7e11 = hbusreq2_p & v9f7dfd | !hbusreq2_p & v9f7e10;
assign v9f773a = hbusreq2_p & v9f7737 | !hbusreq2_p & v9f7739;
assign bd5827 = hbusreq1 & bd5771 | !hbusreq1 & !v845542;
assign b1c5da = hmaster0_p & v845542 | !hmaster0_p & b1c5d9;
assign b1c6c8 = hgrant1_p & v845542 | !hgrant1_p & b1c6c7;
assign ad468e = hbusreq1 & ad4570 | !hbusreq1 & v845542;
assign c3d4f8 = hgrant1_p & v84554d | !hgrant1_p & c3d4f7;
assign v9ea619 = hgrant3_p & v9ea5fa | !hgrant3_p & v9ea618;
assign c3cf0d = hbusreq1 & c3cf03 | !hbusreq1 & c3cf07;
assign v9ea56e = hmaster1_p & v9ea56d | !hmaster1_p & v9ea56b;
assign ad45bf = hbusreq4 & ad45b9 | !hbusreq4 & !ad45be;
assign b1c828 = hmaster0_p & b1c825 | !hmaster0_p & b1c777;
assign b57ab5 = hmaster0_p & b57ab4 | !hmaster0_p & v845542;
assign ad41b2 = hbusreq2_p & ad41b1 | !hbusreq2_p & v845542;
assign d3557f = hbusreq0 & d3557b | !hbusreq0 & d3557e;
assign bd5b82 = hmaster2_p & v84556c | !hmaster2_p & bd5b81;
assign cc36cc = hbusreq4_p & cc36cb | !hbusreq4_p & !cc36ca;
assign ad413d = hmaster2_p & ad413c | !hmaster2_p & ad4f0a;
assign d35617 = hmastlock_p & d35616 | !hmastlock_p & v845542;
assign b57a6a = hbusreq4 & b57a69 | !hbusreq4 & b57942;
assign df51cf = decide_p & df5537 | !decide_p & d6ebca;
assign d35027 = jx0_p & d3576b | !jx0_p & d35026;
assign v9f7651 = hbusreq2 & v9f764f | !hbusreq2 & v9f7650;
assign c3d5c4 = hgrant1_p & v84554d | !hgrant1_p & c3d5c3;
assign ad469e = hbusreq4_p & ad469d | !hbusreq4_p & v845542;
assign ad4e9b = stateG10_4_p & ad4e98 | !stateG10_4_p & !ad4e9a;
assign v8cc493 = hgrant4_p & v845542 | !hgrant4_p & v8cc492;
assign d35581 = hmaster2_p & d35580 | !hmaster2_p & d3557d;
assign c3d2f7 = hgrant4_p & v845542 | !hgrant4_p & c3d2ef;
assign b5b4ef = hgrant4_p & v845542 | !hgrant4_p & b5b40a;
assign ad4373 = hmaster1_p & ad4325 | !hmaster1_p & ad431c;
assign b05914 = hmaster1_p & b05902 | !hmaster1_p & b05913;
assign ad46c4 = hbusreq1 & ad457d | !hbusreq1 & v845542;
assign d3577c = hmaster0_p & d35778 | !hmaster0_p & d3577b;
assign d3552c = hmaster1_p & d35523 | !hmaster1_p & d3552b;
assign b1c7ea = hbusreq2 & b1c743 | !hbusreq2 & !v845542;
assign b1c5ef = hmaster0_p & b1cfb8 | !hmaster0_p & b1c5ee;
assign c3d597 = hbusreq1 & c3d58f | !hbusreq1 & c3d591;
assign c3d52c = hbusreq3 & c3d527 | !hbusreq3 & c3d52b;
assign dc52fa = locked_p & dc52f9 | !locked_p & !v845542;
assign ad4897 = hmaster0_p & ad4851 | !hmaster0_p & ad4896;
assign v9f7796 = hlock1 & v9f772d | !hlock1 & v9f7795;
assign b574c5 = hlock4 & b579ce | !hlock4 & b574c4;
assign d3568b = hbusreq2_p & d3562f | !hbusreq2_p & d35aa0;
assign ad457c = hbusreq4 & ade4ad | !hbusreq4 & v845542;
assign b1c6da = hbusreq1_p & b1c617 | !hbusreq1_p & b1c848;
assign d3551f = hmaster2_p & d3551e | !hmaster2_p & d35a9b;
assign ad473f = hbusreq1 & ad472f | !hbusreq1 & ad4732;
assign ad4e60 = hbusreq2 & ad4e5f | !hbusreq2 & v845542;
assign v9f7d35 = hmaster0_p & v9f7d03 | !hmaster0_p & v9f7d34;
assign ad4592 = hmaster1_p & ad4589 | !hmaster1_p & ad4591;
assign cc36ce = hgrant1_p & df54f3 | !hgrant1_p & cc36cd;
assign b0596c = hbusreq1_p & b05962 | !hbusreq1_p & b0596b;
assign ad4df7 = hmaster1_p & ad4df6 | !hmaster1_p & ad4df2;
assign bd5777 = hbusreq3 & c3d68a | !hbusreq3 & !v845542;
assign v8cc6b6 = hbusreq3_p & v8cc629 | !hbusreq3_p & v8cc6b5;
assign v9ea5d5 = hlock2 & v9ea5cb | !hlock2 & v9ea5d4;
assign v8ccb79 = hlock4_p & v8d29fa | !hlock4_p & v845542;
assign v9ea610 = hgrant2_p & v9ea602 | !hgrant2_p & v9ea60f;
assign v9f789e = hgrant2_p & v9f7877 | !hgrant2_p & v9f789d;
assign v9f7d1b = hbusreq1_p & v9f7d05 | !hbusreq1_p & v9f7d12;
assign ad4e0b = hmaster1_p & v845555 | !hmaster1_p & ad4df2;
assign c3ceae = hbusreq1_p & v845542 | !hbusreq1_p & c3cead;
assign d35ab4 = hgrant1_p & v84554c | !hgrant1_p & d35ab3;
assign v9f7dab = hbusreq1_p & v9f7da0 | !hbusreq1_p & v9f7daa;
assign v84554e = hlock1_p & v845542 | !hlock1_p & !v845542;
assign b57ad1 = hmaster1_p & b57ad0 | !hmaster1_p & b57901;
assign adec93 = hbusreq4_p & v84556c | !hbusreq4_p & v845542;
assign ad5071 = hgrant3_p & ad4e41 | !hgrant3_p & ad5070;
assign v8ccb81 = hmaster0_p & v8ccb78 | !hmaster0_p & v8ccb80;
assign ade540 = hbusreq2 & adec8a | !hbusreq2 & adec93;
assign cc36d3 = hmaster1_p & cc36d2 | !hmaster1_p & v845542;
assign c3d372 = locked_p & v845542 | !locked_p & !c3d371;
assign ad45c1 = hbusreq3 & ad45b6 | !hbusreq3 & ad45c0;
assign ad4dd5 = hbusreq3 & ad4dd4 | !hbusreq3 & v845542;
assign ad4e83 = hbusreq4_p & ad4e82 | !hbusreq4_p & b1cfbe;
assign b059bf = stateG2_p & v845542 | !stateG2_p & !b059be;
assign v9f776c = hmaster2_p & v9f776a | !hmaster2_p & v9f776b;
assign c3d4dd = hmaster2_p & c3d4dc | !hmaster2_p & v845542;
assign ad3d49 = hgrant2_p & ad3d47 | !hgrant2_p & ad3d48;
assign ad4759 = hmaster0_p & ad4758 | !hmaster0_p & ad4588;
assign df54d6 = hmaster2_p & v845542 | !hmaster2_p & dc5318;
assign b579af = hmaster0_p & v845542 | !hmaster0_p & b57942;
assign c3ce51 = hbusreq1 & c3d313 | !hbusreq1 & c3d305;
assign dc5073 = hbusreq2 & dc5072 | !hbusreq2 & !v845542;
assign bd5e22 = hlock2_p & bd5e21 | !hlock2_p & v845542;
assign b05a48 = hmaster0_p & b05a0f | !hmaster0_p & b0593d;
assign b57902 = hmaster1_p & b578f9 | !hmaster1_p & b57901;
assign c3d509 = hgrant1_p & v84554d | !hgrant1_p & c3d4f6;
assign v9e9eaa = hbusreq3 & v9e9ea6 | !hbusreq3 & v9e9ea9;
assign ad44b1 = hgrant4_p & ad448c | !hgrant4_p & !c3cec2;
assign v9f776b = hlock0_p & v84557a | !hlock0_p & !v9f7733;
assign ad46e3 = hgrant1_p & ad46c6 | !hgrant1_p & ad46e2;
assign df51db = decide_p & df511a | !decide_p & d6ebca;
assign c3cf30 = hready_p & c3cf2f | !hready_p & !c3d36c;
assign c3cede = hmaster2_p & c3cedd | !hmaster2_p & !v845542;
assign v9ea41b = hbusreq4_p & v9ea418 | !hbusreq4_p & v9ea41a;
assign d3598f = hmaster1_p & d35982 | !hmaster1_p & d3598e;
assign v9f7864 = hbusreq1 & v9f7862 | !hbusreq1 & v9f7863;
assign ad4590 = hbusreq3 & ad458f | !hbusreq3 & v845542;
assign b578f5 = decide_p & b578f4 | !decide_p & b578f3;
assign d3558e = hmaster2_p & d35aac | !hmaster2_p & d3558d;
assign b57af3 = hmaster0_p & b57af2 | !hmaster0_p & v845542;
assign v9f77c2 = hmaster2_p & v9f77c1 | !hmaster2_p & !v845542;
assign v9f7892 = hbusreq2 & v9f7890 | !hbusreq2 & v9f7891;
assign ad42e0 = hbusreq1_p & ad42df | !hbusreq1_p & v845542;
assign ad3ceb = hlock0_p & v84556e | !hlock0_p & c3cec2;
assign ad4e42 = hready & d35980 | !hready & dc4fcb;
assign bd591f = decide_p & bd590e | !decide_p & !v845572;
assign ad4f38 = hburst0 & dc504c | !hburst0 & adea98;
assign ad4388 = hlock0_p & d35a4e | !hlock0_p & !ad4387;
assign bd5795 = hbusreq2 & bd5794 | !hbusreq2 & v845542;
assign c3ce63 = hbusreq1_p & c3ce62 | !hbusreq1_p & v845542;
assign c3ce21 = hgrant2_p & c3ce19 | !hgrant2_p & c3ce20;
assign d3574f = hbusreq1_p & d3571c | !hbusreq1_p & d35aac;
assign v9f78b1 = jx2_p & v9f7c94 | !jx2_p & v9f78b0;
assign v9f785c = hlock0_p & v9f772a | !hlock0_p & v9f785b;
assign d357fe = hbusreq4 & d357fb | !hbusreq4 & d357fd;
assign ad4d96 = hmaster2_p & ad4d91 | !hmaster2_p & v9f21c4;
assign v9ea455 = hbusreq1 & v9ea454 | !hbusreq1 & v9ea3fa;
assign ad5016 = locked_p & ad5015 | !locked_p & !v845542;
assign b058bc = hbusreq4 & b058ba | !hbusreq4 & b058bb;
assign ade655 = hmaster0_p & v845542 | !hmaster0_p & !ade654;
assign ad4e69 = stateG2_p & v845542 | !stateG2_p & ad4e68;
assign v9e9fc8 = hgrant2_p & v9e9fc6 | !hgrant2_p & v9e9fc7;
assign v8cc5f8 = hbusreq3 & v8cc5be | !hbusreq3 & v8ccbd8;
assign adea9b = hgrant4_p & adea9a | !hgrant4_p & !v845542;
assign ba7c70 = decide_p & ba7c68 | !decide_p & ba7c6f;
assign d354ea = hbusreq2_p & d354de | !hbusreq2_p & !d354e9;
assign ad4464 = hmaster2_p & ad4463 | !hmaster2_p & v845542;
assign ad40ed = hmaster1_p & ad40ec | !hmaster1_p & ad4897;
assign d35bee = hbusreq3 & d35bed | !hbusreq3 & d35be8;
assign bd5761 = hbusreq2 & dc4fcb | !hbusreq2 & v845542;
assign d35a0f = stateG10_4_p & d359f7 | !stateG10_4_p & d35a0e;
assign b1c782 = hmaster0_p & b1c77f | !hmaster0_p & b1c777;
assign df5160 = hbusreq1_p & df515f | !hbusreq1_p & v845542;
assign df5129 = hmaster1_p & df54f4 | !hmaster1_p & df5128;
assign ad4ef4 = hgrant4_p & ad4ef3 | !hgrant4_p & ad4e98;
assign v8cc034 = hready_p & v8cc031 | !hready_p & v8cc50c;
assign c3cebe = stateG10_4_p & c3cebc | !stateG10_4_p & c3cebd;
assign df552c = hready_p & df54ff | !hready_p & df552b;
assign v9f7850 = hmaster1_p & v9f784f | !hmaster1_p & v9f7846;
assign v9f7d22 = hlock0_p & v9ea3ec | !hlock0_p & v9f7d21;
assign df5167 = hbusreq1 & dc4f70 | !hbusreq1 & v845542;
assign v9f7681 = hbusreq3 & v9f767e | !hbusreq3 & v9f7680;
assign v8cc75f = hbusreq2 & v8cc75c | !hbusreq2 & v8cc75e;
assign b1c76b = hbusreq1 & b1c768 | !hbusreq1 & b1c76a;
assign ad5069 = hbusreq3 & ad5034 | !hbusreq3 & c3d2d9;
assign ad4f5c = hlock1_p & ad4f5b | !hlock1_p & !v845542;
assign ad5017 = hmaster2_p & v84556c | !hmaster2_p & ad5016;
assign ad446b = hgrant2_p & ad4426 | !hgrant2_p & ad446a;
assign b57501 = hmaster0_p & b57500 | !hmaster0_p & v845542;
assign b57b57 = decide_p & b57a21 | !decide_p & b57aeb;
assign v9f7e1c = hgrant4_p & v9f7cb6 | !hgrant4_p & v9f7d89;
assign b1d003 = hgrant1_p & v845542 | !hgrant1_p & b1d002;
assign v9e9f6e = hbusreq4 & v9e9f6c | !hbusreq4 & v9e9f6d;
assign v9f78a2 = decide_p & v9f789c | !decide_p & v9f78a1;
assign ad4dc7 = hbusreq1 & ad4d98 | !hbusreq1 & ad4dc6;
assign v9f784a = hgrant1_p & v9f779f | !hgrant1_p & v9f782f;
assign v9ea4d1 = stateG10_4_p & v9ea464 | !stateG10_4_p & v9ea4d0;
assign c5c8a0 = hmaster1_p & c5c897 | !hmaster1_p & c5c89f;
assign bd5844 = hgrant4_p & c3d674 | !hgrant4_p & !bd5842;
assign v9f7e3a = hbusreq1_p & v9f7cae | !hbusreq1_p & v9f7e39;
assign v9f7cf9 = hlock0 & v9f7cf8 | !hlock0 & v9f7cf6;
assign c3d6c5 = stateG10_4_p & c3d6b8 | !stateG10_4_p & c3d6c4;
assign ade622 = hmaster0_p & ade5c9 | !hmaster0_p & ade4d0;
assign d6ebcb = hready_p & d6ebca | !hready_p & !v845560;
assign v9f7d7a = hgrant4_p & v9f7cb4 | !hgrant4_p & v9f7d79;
assign v9ea446 = hgrant4_p & v9ea3fb | !hgrant4_p & v9ea445;
assign v9f7743 = hmastlock_p & v9f7742 | !hmastlock_p & !v845542;
assign d357ea = hbusreq1_p & v84554a | !hbusreq1_p & d357e9;
assign v9f76ec = hgrant0_p & v9f7ca4 | !hgrant0_p & !v9f76eb;
assign d3569f = hbusreq1 & d3569e | !hbusreq1 & v845542;
assign v9ea4b2 = hbusreq2_p & v9ea4b0 | !hbusreq2_p & v9ea4b1;
assign v9e9ed4 = hgrant2_p & v9e9ed2 | !hgrant2_p & v9e9ed3;
assign dc507f = hmaster1_p & dc507e | !hmaster1_p & dc5067;
assign b1c7fa = decide_p & b1c7f9 | !decide_p & b1c866;
assign v8cc7b8 = hbusreq2 & v8cc7b5 | !hbusreq2 & v8cc7b6;
assign v9f7e07 = hlock1_p & v9f7cc8 | !hlock1_p & v9f7d12;
assign d3565a = hmaster0_p & d35649 | !hmaster0_p & d35659;
assign ad458d = hbusreq3 & ad458c | !hbusreq3 & !v845542;
assign adeaac = hready_p & adeaa8 | !hready_p & adeaab;
assign v9f7771 = hlock2 & v9f7751 | !hlock2 & v9f7770;
assign c3d6fe = hgrant2_p & c3d6a3 | !hgrant2_p & c3d6fd;
assign dc5061 = hbusreq4_p & dc505e | !hbusreq4_p & dc5060;
assign v9f7857 = hmaster1_p & v9f7856 | !hmaster1_p & v9f776d;
assign ad45a3 = hbusreq4 & ad45a2 | !hbusreq4 & v845542;
assign c5c8eb = hmaster0_p & c5c8e9 | !hmaster0_p & !v845542;
assign bd5ba7 = decide_p & bd5ba6 | !decide_p & v845542;
assign bd58d8 = hgrant2_p & v845542 | !hgrant2_p & bd58d7;
assign d356c9 = hmaster0_p & d356c6 | !hmaster0_p & !d356c8;
assign b05a0d = hmaster2_p & b05a09 | !hmaster2_p & !b05a0c;
assign v9f76f7 = hready & v9f76f6 | !hready & v9f76f2;
assign bd5b94 = hmaster2_p & v84556c | !hmaster2_p & !bd5b93;
assign dc5053 = stateG10_4_p & adeca1 | !stateG10_4_p & !dc5052;
assign v9f7e18 = hmaster2_p & v9f7e14 | !hmaster2_p & !v9f7e17;
assign v9f7873 = hbusreq2_p & v9f785a | !hbusreq2_p & v9f7872;
assign ad456e = hbusreq4 & ad456d | !hbusreq4 & v845542;
assign v8cc476 = stateA1_p & v8d29f9 | !stateA1_p & v8d29f8;
assign b57909 = hmaster1_p & b578fa | !hmaster1_p & b57901;
assign v8cc7e4 = hready & v8cc7e3 | !hready & v8ccb6b;
assign ad4e7a = hmaster2_p & ad4e79 | !hmaster2_p & v845542;
assign cc36c2 = decide_p & v845566 | !decide_p & cc36c1;
assign v9f7dc8 = hgrant4_p & v9f7ca0 | !hgrant4_p & v9f7d79;
assign v9ea4a9 = hbusreq1_p & v9f20a1 | !hbusreq1_p & v9ea4a7;
assign d356d1 = decide_p & d356d0 | !decide_p & v84556c;
assign v9f7826 = hlock3 & v9f77d0 | !hlock3 & v9f7825;
assign v9f774e = hlock2 & v9f7745 | !hlock2 & v9f774d;
assign b1c823 = hbusreq2_p & b1c801 | !hbusreq2_p & b1c822;
assign ad45b7 = hlock4_p & ad4d9a | !hlock4_p & !ad4de2;
assign bd5b9d = decide_p & bd5b9c | !decide_p & v845572;
assign c5c8e3 = stateG2_p & v845542 | !stateG2_p & !v845568;
assign ad5060 = stateG10_4_p & ad505e | !stateG10_4_p & !ad505f;
assign v9f7db0 = hgrant4_p & v9f7cc6 | !hgrant4_p & v9f7dae;
assign cc36d5 = hlock2_p & cc36d1 | !hlock2_p & !cc36d4;
assign b579d7 = stateG10_4_p & v845542 | !stateG10_4_p & b579d6;
assign ad4819 = hmaster1_p & ad4818 | !hmaster1_p & v845542;
assign d357fb = hbusreq0 & d357f9 | !hbusreq0 & d357fa;
assign ade57c = hbusreq0 & ade57b | !hbusreq0 & ade567;
assign c3d5e8 = hbusreq0 & c3d5e7 | !hbusreq0 & adeaa5;
assign d357c6 = hbusreq4_p & d357c4 | !hbusreq4_p & d357c5;
assign v9f7db9 = hready & v9f7db8 | !hready & v9f7db4;
assign b57430 = hlock2 & b578f1 | !hlock2 & b5742f;
assign c3d316 = hbusreq3 & c3d315 | !hbusreq3 & c3d306;
assign cc36da = hgrant0_p & cc36bd | !hgrant0_p & !v845566;
assign ad4ee2 = hbusreq4_p & ad4ed3 | !hbusreq4_p & ad4ee1;
assign b57956 = hgrant1_p & v845542 | !hgrant1_p & b57955;
assign v9f7840 = hbusreq4_p & d35a0b | !hbusreq4_p & !v9f783f;
assign bd58d7 = hmaster1_p & bd58b5 | !hmaster1_p & bd58d6;
assign c3d301 = hready & c3d2fa | !hready & c3d300;
assign ad4d9b = hmaster2_p & v845542 | !hmaster2_p & ad4d9a;
assign b1c6bd = hmaster1_p & b1cfb8 | !hmaster1_p & b1c6bc;
assign d356af = hmaster0_p & d356a9 | !hmaster0_p & d356ae;
assign b1cf30 = hlock0_p & bd56d1 | !hlock0_p & v845542;
assign ad410e = hlock1_p & ad410d | !hlock1_p & v845547;
assign b05a33 = hmaster1_p & b05a32 | !hmaster1_p & b058e1;
assign dc5029 = stateG10_4_p & adeca1 | !stateG10_4_p & !dc5028;
assign v9f788d = hbusreq1_p & v9f77de | !hbusreq1_p & v9f788c;
assign v9f7cda = hbusreq4_p & v9f7cb6 | !hbusreq4_p & !v9f7cc7;
assign bd588f = hgrant4_p & v84556c | !hgrant4_p & bd5875;
assign c3ce96 = decide_p & c3ce91 | !decide_p & !c3ce95;
assign c5c8e7 = locked_p & c5c8e6 | !locked_p & c5c896;
assign v9e9e7c = hbusreq2_p & v9e9e78 | !hbusreq2_p & v9e9e7b;
assign v9e9ecb = hready_p & v9ea4a4 | !hready_p & v9e9eca;
assign v9f7d48 = hmaster1_p & v9f7d3b | !hmaster1_p & v9f7d47;
assign b57aec = decide_p & b57adf | !decide_p & b57aeb;
assign b579ed = hbusreq3 & b579ec | !hbusreq3 & b57942;
assign bd57f6 = hburst0 & ade54d | !hburst0 & bd57f5;
assign bd5e9a = hbusreq4_p & bd5e99 | !hbusreq4_p & v84556c;
assign ad440e = hready & ad440d | !hready & !v845564;
assign ba05d0 = hgrant3_p & ba05cf | !hgrant3_p & ba05cd;
assign d3562c = hlock2_p & v845542 | !hlock2_p & !d3562b;
assign b059d9 = hbusreq0_p & b0597e | !hbusreq0_p & !b059d8;
assign bd5889 = hgrant4_p & bd587d | !hgrant4_p & bd580d;
assign ade59c = hlock0_p & ade595 | !hlock0_p & !ade59b;
assign dc5387 = hgrant3_p & dc5320 | !hgrant3_p & !dc5386;
assign c3cf14 = hgrant2_p & c3cf13 | !hgrant2_p & c3cf10;
assign v9ea49c = hmaster1_p & v9ea49b | !hmaster1_p & v9ea48a;
assign dc4fc9 = hmaster2_p & adec89 | !hmaster2_p & v845542;
assign d357de = hmaster0_p & d357d3 | !hmaster0_p & d357dd;
assign df5153 = hmaster1_p & df5152 | !hmaster1_p & df514d;
assign v9e9f57 = hmaster2_p & v9e9f56 | !hmaster2_p & v9ea448;
assign d35949 = hburst1_p & v845542 | !hburst1_p & !c74a04;
assign v8ccbd7 = hlock3_p & v8ccb88 | !hlock3_p & v8ccbd6;
assign c5c9a0 = decide_p & v845542 | !decide_p & c5c99f;
assign c3cf09 = hbusreq3 & c3cf04 | !hbusreq3 & c3cf08;
assign ad4555 = hbusreq4_p & ad4e47 | !hbusreq4_p & v845542;
assign v9e9f84 = hgrant1_p & v9e9f82 | !hgrant1_p & v9e9f83;
assign v8cc167 = hready_p & v8cc455 | !hready_p & v8cc819;
assign c3d669 = hmastlock_p & c3d667 | !hmastlock_p & c3d668;
assign bd5e99 = hlock4_p & bd5b81 | !hlock4_p & dc52fa;
assign b1c065 = hbusreq4_p & b1c798 | !hbusreq4_p & !b1c064;
assign c5c96b = hmaster0_p & c5c969 | !hmaster0_p & c5c96a;
assign d35a07 = stateG10_4_p & d35a03 | !stateG10_4_p & d35a05;
assign v9ea5f7 = hmaster1_p & v9ea5f6 | !hmaster1_p & v9ea4bd;
assign ad3ce0 = hbusreq0 & ad3cdf | !hbusreq0 & v845542;
assign ad4298 = hmaster1_p & ad4294 | !hmaster1_p & ad4297;
assign v9f7dd9 = hlock4_p & v9f7dd7 | !hlock4_p & v9f7dd8;
assign ad42ee = hgrant1_p & v845542 | !hgrant1_p & ad42ed;
assign c3d6d1 = hgrant1_p & c3d6c0 | !hgrant1_p & !c3d6d0;
assign c3d5c0 = hmaster2_p & c3d5bf | !hmaster2_p & c3d2fd;
assign b1c5bc = hmaster2_p & v845542 | !hmaster2_p & b1c5bb;
assign b573e3 = hlock3 & b57942 | !hlock3 & b573e2;
assign df54fc = hmaster1_p & df54f4 | !hmaster1_p & df54fb;
assign ac1462 = hlock4_p & ac1461 | !hlock4_p & adea92;
assign ad4eb1 = hbusreq1 & ad4eb0 | !hbusreq1 & !v845547;
assign b1cbf2 = hmaster2_p & b1cfb7 | !hmaster2_p & b1cbf1;
assign b574ca = hgrant1_p & v845542 | !hgrant1_p & b574c9;
assign v9e9eb0 = hbusreq1 & v9ea453 | !hbusreq1 & v9ea3fa;
assign v8cc6b8 = jx0_p & v8cc50f | !jx0_p & v8cc6b7;
assign ac1458 = hgrant0_p & v845542 | !hgrant0_p & !ac144e;
assign df5544 = hbusreq3_p & df552d | !hbusreq3_p & df5543;
assign d35760 = decide_p & d3575f | !decide_p & v84556c;
assign d354cd = hmaster2_p & v845542 | !hmaster2_p & d354cc;
assign b57a85 = hlock3 & b57942 | !hlock3 & b57a84;
assign c3d67e = hmaster0_p & c3d66f | !hmaster0_p & c3d676;
assign ad4eb7 = hbusreq4_p & ad4eb4 | !hbusreq4_p & ad4eb6;
assign df514f = hbusreq1 & dc4fd4 | !hbusreq1 & v845542;
assign bd590f = decide_p & bd590e | !decide_p & v845542;
assign ad4134 = hmaster2_p & ad4133 | !hmaster2_p & ad4efb;
assign b1c760 = hbusreq1 & b1c758 | !hbusreq1 & b1c75c;
assign v9e9fe1 = hgrant2_p & v9e9e68 | !hgrant2_p & v9e9fe0;
assign ad4788 = decide_p & ad4785 | !decide_p & ad4787;
assign ac1494 = hgrant3_p & ac1484 | !hgrant3_p & ac1493;
assign b1c80c = hmaster0_p & b1c806 | !hmaster0_p & b1c80b;
assign v9ea477 = hgrant4_p & v9ea44d | !hgrant4_p & v9ea457;
assign ad46be = hmaster2_p & ad4699 | !hmaster2_p & ad46bd;
assign ad4fa0 = hgrant2_p & ad4f50 | !hgrant2_p & ad4f9f;
assign c5c89a = hbusreq1_p & c5c899 | !hbusreq1_p & c5c898;
assign b059e4 = hgrant4_p & b058d4 | !hgrant4_p & !b059e3;
assign ad3d59 = hbusreq2_p & ad3d53 | !hbusreq2_p & ad3d58;
assign d35bec = hbusreq3 & d35be6 | !hbusreq3 & d35beb;
assign b058d8 = hlock4 & b058d5 | !hlock4 & b058d7;
assign b1cfd3 = hmaster0_p & b1cfb8 | !hmaster0_p & b1cfd2;
assign bd5803 = hmaster2_p & bd5802 | !hmaster2_p & dc5001;
assign v9f7803 = hgrant1_p & v9f772c | !hgrant1_p & v9f77df;
assign d357cc = hmaster2_p & d357c6 | !hmaster2_p & d357cb;
assign b1c7f4 = hbusreq1_p & b1c7f2 | !hbusreq1_p & b1c7f3;
assign b059f1 = hlock3 & b059f0 | !hlock3 & b059ef;
assign d35be4 = hlock4_p & d359b7 | !hlock4_p & dc52fa;
assign b1c7d0 = hgrant4_p & ade589 | !hgrant4_p & !b1c79d;
assign c3d3a3 = hbusreq4 & c3d39e | !hbusreq4 & !c3d3a2;
assign ad42cc = hmaster1_p & ad42cb | !hmaster1_p & ad42bd;
assign c3d6f3 = stateG10_4_p & c3d6b7 | !stateG10_4_p & c3d6f2;
assign c3ce6a = hbusreq1 & c3d2d6 | !hbusreq1 & v845542;
assign ad4eb0 = hready & ad4eaf | !hready & v845542;
assign b0591c = hmastlock_p & b058a4 | !hmastlock_p & v845542;
assign v9e9f66 = locked_p & v9f20a1 | !locked_p & v9e9f65;
assign ad4328 = hgrant2_p & ad4322 | !hgrant2_p & ad4327;
assign bd5b84 = stateA1_p & v845542 | !stateA1_p & !v8ccb67;
assign b5741c = hlock0_p & b57952 | !hlock0_p & b5741b;
assign d3590b = hbusreq3 & d3590a | !hbusreq3 & v845542;
assign dc53b3 = hready_p & v845542 | !hready_p & dc53b2;
assign v9f78ac = hready_p & v9f78a2 | !hready_p & v9f78ab;
assign d35ab1 = hbusreq4_p & v845542 | !hbusreq4_p & d35ab0;
assign b058cf = hbusreq0_p & b058b6 | !hbusreq0_p & v9f7d42;
assign ad43bc = hmaster0_p & ad43a9 | !hmaster0_p & ad43aa;
assign v9f7c93 = jx1_p & v845542 | !jx1_p & v857467;
assign ad432d = hbusreq1 & v845542 | !hbusreq1 & v845547;
assign v8cc4fd = hmaster2_p & v8cc4fc | !hmaster2_p & v845542;
assign v9f7dd0 = hlock0_p & v9f7dce | !hlock0_p & !v9f7dcf;
assign c74202 = start_p & v845542 | !start_p & c74198;
assign ad410c = hmaster0_p & ad4106 | !hmaster0_p & ad410b;
assign b579b4 = hgrant1_p & v845542 | !hgrant1_p & b579b3;
assign b05a14 = hmaster2_p & b05a09 | !hmaster2_p & !b05a13;
assign b1c798 = hgrant4_p & b1c70f | !hgrant4_p & !b1c797;
assign v9e9f5a = hbusreq4 & v9e9f58 | !hbusreq4 & v9e9f59;
assign b05920 = hmaster2_p & b0591c | !hmaster2_p & !v9f7d42;
assign c3d58f = hready & c3d58e | !hready & v845542;
assign bd5808 = hgrant4_p & c3d669 | !hgrant4_p & bd5806;
assign c5c9b5 = hgrant3_p & c5c9ab | !hgrant3_p & c5c9b4;
assign v9e9fe8 = jx0_p & v9e9ee6 | !jx0_p & v9e9fe7;
assign b1c704 = decide_p & b1c82f | !decide_p & v845542;
assign c3d761 = hready_p & c3d755 | !hready_p & !c3d760;
assign ba7c77 = jx0_p & ba7c72 | !jx0_p & ba7c76;
assign d35019 = hbusreq4_p & d357d7 | !hbusreq4_p & d35010;
assign d356f4 = hlock1_p & d35991 | !hlock1_p & df54f5;
assign v8cc82e = hbusreq2_p & v8cc7d5 | !hbusreq2_p & v8cc82c;
assign b0599d = hbusreq3 & b0599a | !hbusreq3 & b0599c;
assign dc503c = hbusreq4_p & dc5038 | !hbusreq4_p & dc503b;
assign v9f7d9a = hbusreq1_p & v9f7d99 | !hbusreq1_p & v9f7d05;
assign v9f7d15 = hlock4 & v9f7d12 | !hlock4 & v9f7d14;
assign c3d6cc = hgrant4_p & c3d67a | !hgrant4_p & !c3d6cb;
assign dc5317 = hmaster2_p & v845542 | !hmaster2_p & !dc5316;
assign bd585a = hbusreq1_p & bd5858 | !hbusreq1_p & bd5859;
assign c3ce48 = hgrant1_p & v84554d | !hgrant1_p & c3ce47;
assign b05a81 = hmaster0_p & b05a80 | !hmaster0_p & b0599f;
assign v9f788f = hlock3 & v9f77fa | !hlock3 & v9f788e;
assign b1c7c1 = hmaster2_p & b1c79b | !hmaster2_p & b1c7c0;
assign c3cea0 = hgrant1_p & c3d2d9 | !hgrant1_p & c3ce9f;
assign ade5ce = hburst0 & ade4c8 | !hburst0 & ade5cd;
assign v8cc4f4 = hbusreq2_p & v8ccb8f | !hbusreq2_p & v8cc4f3;
assign v9ea4ae = hmaster2_p & v9ea4ab | !hmaster2_p & v9ea4ad;
assign v8ccb7b = hbusreq4_p & v8ccb79 | !hbusreq4_p & v845542;
assign e199ba = hburst1_p & c76647 | !hburst1_p & v845542;
assign v9ea5ae = hlock3 & v9ea586 | !hlock3 & v9ea5ad;
assign v9e9ee1 = hbusreq2_p & v9e9ee0 | !hbusreq2_p & v9ea615;
assign bd572e = locked_p & v845542 | !locked_p & c3d669;
assign c3d673 = stateA1_p & v845542 | !stateA1_p & v889629;
assign v9f7704 = hbusreq1_p & v9f7d90 | !hbusreq1_p & v9f76f2;
assign ad4561 = hmaster2_p & v845542 | !hmaster2_p & ad4555;
assign bd56da = hbusreq2 & dc5317 | !hbusreq2 & bd56d9;
assign ad4485 = hmaster2_p & ad447b | !hmaster2_p & v845542;
assign ad4418 = hready & ad4417 | !hready & !v845542;
assign bd579d = hlock1_p & bd5799 | !hlock1_p & bd579c;
assign c5c92f = locked_p & c5c92e | !locked_p & v845542;
assign ad4347 = hgrant2_p & ad4346 | !hgrant2_p & ad4341;
assign ade54f = hburst0 & ade54c | !hburst0 & ade54e;
assign b574c0 = hgrant4_p & b574b2 | !hgrant4_p & v845542;
assign b57a66 = hbusreq4_p & b579ba | !hbusreq4_p & b57941;
assign d357c4 = hlock4_p & d357c2 | !hlock4_p & d357c3;
assign v9f7e33 = hlock0 & v9f7e32 | !hlock0 & v9f7e30;
assign v9e9f7a = hbusreq0 & v9e9f78 | !hbusreq0 & v9e9f79;
assign v8cc4ba = hmaster0_p & v845542 | !hmaster0_p & v8cc4b9;
assign v9e9fa5 = hlock2 & v9e9f68 | !hlock2 & v9e9fa4;
assign ad3cbc = hmaster1_p & ad4488 | !hmaster1_p & ad3cbb;
assign b1c7ba = hbusreq1_p & b1c7b2 | !hbusreq1_p & b1c7b9;
assign df553e = hgrant2_p & v845542 | !hgrant2_p & !df553d;
assign c3d5b0 = hready_p & v845555 | !hready_p & c3d5af;
assign v9ea569 = hbusreq4_p & v9ea3ee | !hbusreq4_p & v9ea4ad;
assign b05a3b = hmaster1_p & b05a3a | !hmaster1_p & b05926;
assign ad480f = hmaster0_p & ad480b | !hmaster0_p & ad480e;
assign v9ea4c6 = hgrant0_p & v9ea4b6 | !hgrant0_p & v9ea4a6;
assign b1c82f = hmaster1_p & v845542 | !hmaster1_p & b1c82e;
assign b05917 = hbusreq2_p & b05914 | !hbusreq2_p & b05916;
assign v9f7de5 = stateG10_4_p & v9f7de1 | !stateG10_4_p & v9f7de3;
assign d356f6 = hlock1_p & v845542 | !hlock1_p & df54f6;
assign ad4575 = hbusreq4 & ad4574 | !hbusreq4 & v845542;
assign b0593d = hmaster2_p & b05939 | !hmaster2_p & !v9f769c;
assign d356d7 = hbusreq1 & d356d6 | !hbusreq1 & v845542;
assign v8cc7f7 = hbusreq0_p & v8cc7bc | !hbusreq0_p & v8cc7f4;
assign ade55e = hmaster2_p & ade559 | !hmaster2_p & ade55d;
assign ad4725 = decide_p & ad46fa | !decide_p & ad4724;
assign bd57ce = hmaster0_p & bd57cc | !hmaster0_p & bd57cd;
assign b1c765 = hbusreq1 & b1c762 | !hbusreq1 & b1c764;
assign d3556f = hlock2_p & d3556a | !hlock2_p & !d3556e;
assign cc36f0 = hready_p & cc36ef | !hready_p & !cc36c2;
assign ad4de4 = hbusreq3 & ad4de3 | !hbusreq3 & !v845542;
assign v9ea573 = hmaster0_p & v9ea571 | !hmaster0_p & v9ea572;
assign c3d2ff = hbusreq0 & v845576 | !hbusreq0 & c3d2fe;
assign bd5757 = hlock0_p & adec89 | !hlock0_p & bd5756;
assign df5132 = hready_p & df5131 | !hready_p & df512d;
assign d35691 = hmaster1_p & d35690 | !hmaster1_p & d3565a;
assign d35775 = hmaster2_p & d3576e | !hmaster2_p & d35774;
assign ad476a = hbusreq4 & ad4766 | !hbusreq4 & !ad4769;
assign ad4ea7 = hready & ad4e81 | !hready & ad4ea6;
assign ad4df2 = hmaster0_p & ad4dea | !hmaster0_p & !ad4df1;
assign b57444 = hmaster0_p & b57431 | !hmaster0_p & v845542;
assign ac145f = hbusreq1_p & ac145e | !hbusreq1_p & cc36b8;
assign bd57fc = hgrant0_p & bd572e | !hgrant0_p & bd57fb;
assign v9f766d = hlock1 & v9f7667 | !hlock1 & v9f766c;
assign cc36fe = hlock0_p & v84556c | !hlock0_p & cc36fd;
assign v8cc12d = decide_p & v8cc4f4 | !decide_p & v8cc11f;
assign bd5829 = hmaster2_p & bd5802 | !hmaster2_p & v845542;
assign c3d70a = hgrant1_p & c3d697 | !hgrant1_p & c3d709;
assign v9f782b = hgrant4_p & v9f779d | !hgrant4_p & v9f782a;
assign ad4474 = hmaster1_p & ad4473 | !hmaster1_p & ad4469;
assign v9e9ec8 = hmaster1_p & v9e9ec7 | !hmaster1_p & v9e9e77;
assign v9ea417 = hgrant1_p & v9ea416 | !hgrant1_p & v9ea40f;
assign ad45ab = hbusreq4_p & v9f21c4 | !hbusreq4_p & v845542;
assign b05a60 = hbusreq4_p & b05950 | !hbusreq4_p & b05a5f;
assign b1c807 = hbusreq0 & b1c73d | !hbusreq0 & d35a9c;
assign b058b5 = hbusreq2 & b058b3 | !hbusreq2 & b058b4;
assign v9f7e1a = stateG10_4_p & v9f7d81 | !stateG10_4_p & v9f7e19;
assign bd5b8a = hbusreq3 & bd5b89 | !hbusreq3 & v845542;
assign ad4f6e = hgrant4_p & ad4f4a | !hgrant4_p & ad4f36;
assign ade5d2 = hmaster0_p & ade5c9 | !hmaster0_p & ade5d1;
assign b5b40a = hbusreq0_p & b5b409 | !hbusreq0_p & v845542;
assign ade4ea = hmaster2_p & adeaae | !hmaster2_p & ade4e9;
assign b1cf3e = hlock0_p & bd56d3 | !hlock0_p & v845542;
assign d354a9 = hbusreq4_p & d354a8 | !hbusreq4_p & v845542;
assign b1c7ff = hbusreq3 & b1c7b5 | !hbusreq3 & !b1c7b8;
assign ad4268 = hlock1_p & ad4266 | !hlock1_p & ad4267;
assign adec8c = stateA1_p & v845542 | !stateA1_p & !adec8b;
assign d35767 = decide_p & d35766 | !decide_p & v84556c;
assign v9f77d1 = hlock3 & v9f77d0 | !hlock3 & v9f77cf;
assign b1c05c = hbusreq2 & b1c81c | !hbusreq2 & !b1c81f;
assign v9e9ec1 = hgrant3_p & v9e9e7e | !hgrant3_p & v9e9ec0;
assign ad43d8 = hmaster0_p & ad43d4 | !hmaster0_p & ad43d7;
assign d357f6 = hbusreq0 & d357f5 | !hbusreq0 & d35a99;
assign b1c855 = hlock0_p & cc36fc | !hlock0_p & !v845548;
assign d3500f = hgrant4_p & v84554a | !hgrant4_p & d3580c;
assign b57a7b = hbusreq1 & b57a79 | !hbusreq1 & b57a7a;
assign ac148c = hgrant1_p & v845542 | !hgrant1_p & ac148b;
assign b0597d = hbusreq4_p & b0597a | !hbusreq4_p & !b0597c;
assign b058eb = hlock0 & b058ea | !hlock0 & b058e8;
assign c5c8f9 = hgrant4_p & c5c88e | !hgrant4_p & !v845542;
assign v9f7cb9 = hbusreq0 & v9f7cb5 | !hbusreq0 & v9f7cb8;
assign v9f7d9e = hlock2 & v9f7d9b | !hlock2 & v9f7d9d;
assign ad4f3b = hready & ad4f37 | !hready & ad4f3a;
assign v8cc79d = hlock1 & v8ccb6b | !hlock1 & v8cc79c;
assign cc36c9 = hbusreq4_p & dc500e | !hbusreq4_p & cc36c8;
assign b1c034 = hbusreq0 & b1c033 | !hbusreq0 & !b1c841;
assign v9f7dda = hgrant4_p & v9f7da2 | !hgrant4_p & v9f7dae;
assign bd573d = hmastlock_p & bd5739 | !hmastlock_p & !v845542;
assign dc507d = hbusreq3 & dc507c | !hbusreq3 & v845542;
assign d3572c = hbusreq3 & d3572b | !hbusreq3 & !d35aa4;
assign d357e2 = hlock2_p & d357e0 | !hlock2_p & d357e1;
assign dc5301 = hbusreq4_p & dc5300 | !hbusreq4_p & !v845542;
assign ade5c7 = hbusreq2_p & ade5c3 | !hbusreq2_p & ade5c6;
assign d35921 = hlock2_p & d3591e | !hlock2_p & d35920;
assign b5744c = decide_p & b57a21 | !decide_p & b57440;
assign ad4dbe = hmaster0_p & ad4d94 | !hmaster0_p & ad4dbd;
assign b1cf47 = hlock3_p & b1cf38 | !hlock3_p & b1cf46;
assign c3d757 = hmaster1_p & c3d756 | !hmaster1_p & c3d69b;
assign dc4fc7 = decide_p & dc4fc6 | !decide_p & !v845542;
assign b1c616 = hbusreq1 & b1cf28 | !hbusreq1 & b1cf2c;
assign v9ea5e5 = hmaster1_p & v9ea5b4 | !hmaster1_p & v9ea5aa;
assign ad4e96 = hbusreq1 & ad4e95 | !hbusreq1 & !v845542;
assign d356c0 = hlock1_p & d359ad | !hlock1_p & v845542;
assign v8cc628 = hready_p & v8cc455 | !hready_p & v8cc627;
assign v8cc4b3 = hgrant2_p & v8cc472 | !hgrant2_p & v8cc4b2;
assign b058fd = hbusreq1 & b058fb | !hbusreq1 & b058fc;
assign ad4fb4 = hbusreq1_p & ad4fb3 | !hbusreq1_p & v84556c;
assign v9f77a1 = hbusreq0 & v9f779e | !hbusreq0 & v9f77a0;
assign v8cc765 = hbusreq1_p & v8cc763 | !hbusreq1_p & v8ccbd8;
assign b05958 = stateG10_4_p & b05954 | !stateG10_4_p & b05956;
assign ad4109 = hready & ad4103 | !hready & ad4e90;
assign ad46b3 = hbusreq4 & ad4eaf | !hbusreq4 & !v845542;
assign ad4321 = hmaster0_p & ad4293 | !hmaster0_p & ad4320;
assign v8d29f8 = start_p & v845542 | !start_p & !v845580;
assign ac1491 = hbusreq2_p & ac1470 | !hbusreq2_p & ac1490;
assign v9f787f = locked_p & v9f7742 | !locked_p & v9f772b;
assign c3ced6 = hbusreq2_p & c3ce9a | !hbusreq2_p & c3ced5;
assign ad46cb = hmaster2_p & v845542 | !hmaster2_p & ad46ca;
assign v9f7670 = hgrant1_p & v9f7cdd | !hgrant1_p & v9f7667;
assign dc53a8 = hlock3_p & dc53a7 | !hlock3_p & v845542;
assign d35525 = hbusreq4_p & d35431 | !hbusreq4_p & v84554a;
assign d359e6 = hbusreq4_p & v845542 | !hbusreq4_p & adeca0;
assign ad4fe9 = hbusreq4_p & ad4fe7 | !hbusreq4_p & ad4fe8;
assign b5793f = hbusreq2_p & b5790a | !hbusreq2_p & b57909;
assign c3d2ca = hmaster2_p & c3d2c5 | !hmaster2_p & !v845542;
assign df54e9 = hbusreq3 & df54e5 | !hbusreq3 & df54e8;
assign hmaster1 = b8ef53;
assign v9f77b2 = hlock3 & v9f779f | !hlock3 & v9f77a5;
assign d35430 = hbusreq1_p & d3542f | !hbusreq1_p & d3542e;
assign df51ab = hbusreq1 & dc5070 | !hbusreq1 & v845542;
assign ad4102 = hgrant4_p & v845542 | !hgrant4_p & ad4101;
assign v9f771f = hgrant2_p & v9f771d | !hgrant2_p & v9f771e;
assign v9e9ebb = hmaster0_p & v9e9ea1 | !hmaster0_p & v9e9eba;
assign b058c7 = hmaster2_p & b058a3 | !hmaster2_p & v9f7d42;
assign c3cf00 = hgrant4_p & v845542 | !hgrant4_p & c3ceff;
assign v9f7e0b = hbusreq3 & v9f7e06 | !hbusreq3 & v9f7e0a;
assign b57ac8 = hlock3 & b578f9 | !hlock3 & b57ac7;
assign b05a61 = hmaster2_p & b05a60 | !hmaster2_p & v9f7d42;
assign v9ea5ea = hgrant3_p & v9ea5dd | !hgrant3_p & v9ea5e9;
assign d35c07 = hlock4_p & adeca0 | !hlock4_p & !v845542;
assign bd56d4 = hlock4_p & bd56d1 | !hlock4_p & bd56d3;
assign bd5921 = hgrant3_p & bd5910 | !hgrant3_p & !bd5920;
assign ad42a9 = hbusreq1 & ad4d93 | !hbusreq1 & v845542;
assign v9ea3eb = hbusreq4_p & v9f20a1 | !hbusreq4_p & !v9ea3ea;
assign ad4304 = hlock1_p & ad4eb0 | !hlock1_p & v845542;
assign ad4762 = hbusreq2_p & ad475f | !hbusreq2_p & ad4761;
assign v9f7778 = hlock2 & v9f775a | !hlock2 & v9f7777;
assign ad438e = hbusreq0 & ad438d | !hbusreq0 & v845542;
assign ad3d09 = hbusreq0 & ad3d08 | !hbusreq0 & v845542;
assign c3cef3 = hbusreq0 & c3cef2 | !hbusreq0 & adeaa5;
assign d356fc = hmaster0_p & d356fa | !hmaster0_p & d356fb;
assign b573d8 = hbusreq1_p & b573d7 | !hbusreq1_p & b579ce;
assign dc53bb = hmaster0_p & dc53ba | !hmaster0_p & v84556c;
assign ad46df = hmaster2_p & v845542 | !hmaster2_p & ad46de;
assign b059f0 = hgrant1_p & b058d5 | !hgrant1_p & !b059e7;
assign v9f76ba = hmaster0_p & v9f767b | !hmaster0_p & v9f7cee;
assign b1c0a9 = hmaster1_p & b1c85a | !hmaster1_p & b1c0a8;
assign v9f77a9 = hbusreq3 & v9f77a6 | !hbusreq3 & v9f77a8;
assign v8cc75e = hlock2 & v8cc4ad | !hlock2 & v8cc75c;
assign v9f7df1 = hbusreq1_p & v9f7df0 | !hbusreq1_p & v9f7d23;
assign d3564a = hgrant0_p & adea9a | !hgrant0_p & v84556c;
assign ad46d0 = hmaster2_p & v845542 | !hmaster2_p & ad46cf;
assign ad46b4 = hready & ad46b3 | !hready & v845542;
assign b05a01 = hbusreq2_p & b059f7 | !hbusreq2_p & b05a00;
assign d357d0 = hlock1_p & d357cf | !hlock1_p & v84554a;
assign ad3d42 = hmaster1_p & ad3d41 | !hmaster1_p & ad43ba;
assign c3d6b9 = hgrant4_p & c3d675 | !hgrant4_p & c3d6b8;
assign v9e9fdc = hready_p & v9ea3e3 | !hready_p & v9e9fdb;
assign b05a9d = jx0_p & b05a9c | !jx0_p & v867d75;
assign ad427c = hbusreq1_p & ad4f2a | !hbusreq1_p & v845542;
assign ad13e0 = decide_p & ad13df | !decide_p & v84554c;
assign v9ea568 = hbusreq1_p & v9f20a1 | !hbusreq1_p & v9ea567;
assign adea98 = hmastlock_p & adea97 | !hmastlock_p & v845542;
assign b05a11 = hgrant4_p & v9f769c | !hgrant4_p & v9f769d;
assign ad4fc4 = hbusreq3 & ad4fc3 | !hbusreq3 & v845542;
assign bd5918 = hbusreq2 & bd5913 | !hbusreq2 & bd5917;
assign v9f7808 = hbusreq2 & v9f7806 | !hbusreq2 & v9f7807;
assign dc4fdd = hmaster1_p & dc4fd3 | !hmaster1_p & dc4fdc;
assign d35749 = hbusreq2 & d35729 | !hbusreq2 & !d35aa4;
assign df515d = hbusreq1 & dc4f66 | !hbusreq1 & v845564;
assign ad4ec6 = hready & ad4ec2 | !hready & ad4ec5;
assign v8cc5ff = decide_p & v8cc4f4 | !decide_p & v8cc5fe;
assign ad3d2b = hbusreq3 & ad3ce5 | !hbusreq3 & ad3ce7;
assign v8cc5b2 = hlock3 & v8cc4ad | !hlock3 & v8cc5b1;
assign ad5049 = hgrant0_p & ad5048 | !hgrant0_p & !v845542;
assign dc5033 = hmaster2_p & dc5032 | !hmaster2_p & ade581;
assign b1c600 = decide_p & b1c5ff | !decide_p & b1c5f4;
assign c5c897 = hmaster2_p & c5c896 | !hmaster2_p & c5c88d;
assign ad4f79 = hgrant4_p & v845542 | !hgrant4_p & ad4f36;
assign b1c7e0 = hbusreq0 & b1c7df | !hbusreq0 & b1cfcc;
assign df5127 = hgrant1_p & df5126 | !hgrant1_p & !v845542;
assign v9f7d4f = hmaster0_p & v9f7d3c | !hmaster0_p & v9f7d3b;
assign bd5794 = hbusreq3 & bd5787 | !hbusreq3 & bd5793;
assign ade5a3 = hgrant1_p & ade585 | !hgrant1_p & !ade5a2;
assign v9e9ede = hmaster1_p & v9ea580 | !hmaster1_p & v9ea4bd;
assign dc5004 = hgrant4_p & c3d66d | !hgrant4_p & ade563;
assign v9ea5ce = hbusreq0 & v9ea5cc | !hbusreq0 & v9ea5cd;
assign v8cc61c = hbusreq2 & v8cc61a | !hbusreq2 & v8cc489;
assign ade5ac = hbusreq1_p & ade548 | !hbusreq1_p & ade5ab;
assign ad4397 = hmaster2_p & ad4396 | !hmaster2_p & v845542;
assign bbbcd6 = stateG3_0_p & v845580 | !stateG3_0_p & !v845580;
assign b57954 = hgrant4_p & v845542 | !hgrant4_p & b57953;
assign b57944 = hmaster1_p & b57943 | !hmaster1_p & v845542;
assign bd581b = stateG10_4_p & bd5806 | !stateG10_4_p & !bd581a;
assign b57a70 = hlock3 & b579c5 | !hlock3 & b57a6f;
assign c3d4fe = hmaster2_p & v845576 | !hmaster2_p & c3d4f0;
assign ad3d15 = hbusreq2 & ad3ce5 | !hbusreq2 & ad3ce7;
assign v8cc593 = hbusreq0 & v8cc590 | !hbusreq0 & v8cc592;
assign d354e5 = hbusreq1_p & d354e4 | !hbusreq1_p & !d354e3;
assign v9f7cd5 = hbusreq2 & v9f7cd3 | !hbusreq2 & v9f7cd4;
assign b57a26 = hmaster2_p & b57a25 | !hmaster2_p & v845542;
assign c3ce8c = hbusreq3 & v845542 | !hbusreq3 & v845564;
assign v8cc4a2 = hmaster2_p & v8cc4a0 | !hmaster2_p & v8cc499;
assign c3d687 = hbusreq4_p & c3d66d | !hbusreq4_p & !c3d674;
assign c3d72e = hmaster1_p & c3d72d | !hmaster1_p & c3d69b;
assign v9f7d4d = hmaster1_p & v9f7d4c | !hmaster1_p & v9f7d47;
assign v9ea46f = hbusreq0_p & v9f20a1 | !hbusreq0_p & v9ea46e;
assign bd57e3 = hlock2_p & bd57b2 | !hlock2_p & !bd57e2;
assign d35649 = hgrant1_p & d35648 | !hgrant1_p & d35644;
assign ad3d0f = hbusreq0 & ad3d0e | !hbusreq0 & v845542;
assign c3d752 = hmaster1_p & c3d701 | !hmaster1_p & c3d6fc;
assign v9e9ee8 = hmaster2_p & v9e9ee7 | !hmaster2_p & v9f20a1;
assign ad415d = hbusreq4 & ad4158 | !hbusreq4 & ad415c;
assign d35711 = hbusreq2 & d356c5 | !hbusreq2 & !v84554e;
assign ad4fa2 = hlock2_p & ad4fa0 | !hlock2_p & !ad4fa1;
assign ad43dc = hbusreq0 & ad43da | !hbusreq0 & v845542;
assign b059c8 = hready & b059c7 | !hready & b058a8;
assign v9f77e3 = hlock3 & v9f77e2 | !hlock3 & v9f77e0;
assign v9ea432 = hgrant1_p & v845542 | !hgrant1_p & v9ea431;
assign d35740 = hmaster0_p & d3571e | !hmaster0_p & d35702;
assign c3d351 = hbusreq3 & c3d350 | !hbusreq3 & c3d306;
assign v9ea46e = hgrant0_p & v9ea44d | !hgrant0_p & v9ea3e6;
assign d35793 = hmaster2_p & d3578a | !hmaster2_p & d35792;
assign c3d2fd = hgrant4_p & v845542 | !hgrant4_p & v84556e;
assign dc4f84 = hmaster1_p & dc4f6d | !hmaster1_p & dc4f83;
assign ad42b3 = hbusreq0 & ad42b1 | !hbusreq0 & ad42b2;
assign b1c703 = hbusreq3_p & b1c6cf | !hbusreq3_p & b1c702;
assign bb9bdc = hburst1_p & v845542 | !hburst1_p & !v845568;
assign v9f7814 = hmaster1_p & v9f77ff | !hmaster1_p & v9f7811;
assign ad4769 = hmaster2_p & ad45bb | !hmaster2_p & !ad4768;
assign b059ca = hbusreq1 & b059c8 | !hbusreq1 & b059c9;
assign b1c7cc = hbusreq1 & b1c727 | !hbusreq1 & b1c729;
assign c5c890 = hmaster0_p & c5c88f | !hmaster0_p & v845542;
assign ad3cbb = hmaster0_p & ad449a | !hmaster0_p & ad44b7;
assign ad5035 = hbusreq1_p & ad5018 | !hbusreq1_p & ad5034;
assign v9f7df7 = hmaster0_p & v9f7dc5 | !hmaster0_p & !v9f7df6;
assign v8cc0ce = hready & v8cc0ca | !hready & v8ccbd8;
assign v9ea587 = hbusreq4_p & v9ea44d | !hbusreq4_p & v9ea4b3;
assign b1c059 = hbusreq2 & b1c803 | !hbusreq2 & !b1c805;
assign c3d2cd = hbusreq2 & c3d2c9 | !hbusreq2 & c3d2cc;
assign d35a7b = decide_p & d35a7a | !decide_p & v84556c;
assign ad3cc3 = hgrant2_p & ad3cbf | !hgrant2_p & ad3cc2;
assign c3d716 = hmaster1_p & c3d715 | !hmaster1_p & c3d70f;
assign v9e9eb6 = hmaster0_p & v9ea3fc | !hmaster0_p & v9e9eb5;
assign c3cf2f = hgrant2_p & v845551 | !hgrant2_p & c3cf2e;
assign ad4131 = hgrant4_p & dc52fa | !hgrant4_p & ad4e98;
assign ad481f = hmaster1_p & ad481e | !hmaster1_p & ad481d;
assign b05a5d = hlock0_p & b0594f | !hlock0_p & b05a5c;
assign v9f7c9b = hmastlock_p & v9f7c9a | !hmastlock_p & !v845542;
assign v8cc0d2 = hgrant1_p & v8cc0d1 | !hgrant1_p & v8cc474;
assign d3572a = hbusreq3 & d35729 | !hbusreq3 & !d35aa4;
assign v9ea3f8 = hbusreq2_p & v9ea3f1 | !hbusreq2_p & v9ea3f7;
assign d35a1d = hgrant2_p & d3598f | !hgrant2_p & d35a1c;
assign d35729 = hbusreq1_p & d35717 | !hbusreq1_p & v845542;
assign d35a3b = stateA1_p & v845542 | !stateA1_p & !d35a3a;
assign c3d6a8 = hgrant4_p & c3d669 | !hgrant4_p & !c3d6a6;
assign bbbe35 = hburst1_p & v845542 | !hburst1_p & bbbcd8;
assign b059a9 = hgrant1_p & b058c7 | !hgrant1_p & b0596b;
assign v9f77f6 = hgrant2_p & v9f77bc | !hgrant2_p & v9f77f5;
assign b058db = hlock1 & b058d5 | !hlock1 & b058da;
assign ad4da1 = hready & ad4d92 | !hready & !v845542;
assign ad4801 = hbusreq2_p & ad47fc | !hbusreq2_p & ad4800;
assign v8cc5b9 = hmaster0_p & v8cc5a5 | !hmaster0_p & v8cc5b5;
assign v9ea4d4 = hbusreq0_p & v9f20a1 | !hbusreq0_p & v9ea4d3;
assign d35aa5 = hgrant1_p & d35aa4 | !hgrant1_p & v845542;
assign bd5880 = hlock4_p & bd587e | !hlock4_p & !bd587f;
assign bd5815 = hgrant4_p & v845542 | !hgrant4_p & !bd57fe;
assign dc4f6b = hbusreq3 & dc4f6a | !hbusreq3 & v845542;
assign v9e9ea0 = hbusreq1_p & v9e9e9f | !hbusreq1_p & v9ea449;
assign b059b7 = hlock1 & b0595b | !hlock1 & b059b6;
assign c3d38a = hmaster1_p & c3d388 | !hmaster1_p & c3d389;
assign d3595b = hmaster1_p & d3590b | !hmaster1_p & d3595a;
assign ad42e9 = hmaster1_p & ad42e5 | !hmaster1_p & ad42e8;
assign dc4ffa = hgrant1_p & dc4fe2 | !hgrant1_p & dc4ff9;
assign ade665 = jx1_p & adeaad | !jx1_p & adeab8;
assign v8cc62d = hbusreq2 & v8cc62c | !hbusreq2 & v8ccbd8;
assign c3d2b6 = hready & c3d2b5 | !hready & v845564;
assign ad4f4e = hbusreq2 & ad4f4d | !hbusreq2 & v845542;
assign d35aaf = hgrant1_p & d35aa4 | !hgrant1_p & d35aad;
assign v8cc4f2 = hmaster0_p & v8cc4f1 | !hmaster0_p & v8ccb80;
assign d35510 = hbusreq4_p & d3550f | !hbusreq4_p & v845542;
assign v9f7758 = hlock1_p & v9f774b | !hlock1_p & v9f7757;
assign d35520 = hbusreq4_p & d3541e | !hbusreq4_p & v845548;
assign v9e9fac = hbusreq3 & v9e9fa9 | !hbusreq3 & v9e9fab;
assign ad43a3 = hlock3_p & ad43a0 | !hlock3_p & ad43a2;
assign dc4f79 = stateA1_p & adea86 | !stateA1_p & bbb7c7;
assign df511a = hmaster1_p & v845542 | !hmaster1_p & df5119;
assign d3501e = hmaster0_p & d35017 | !hmaster0_p & d3501d;
assign ad4eff = hbusreq4_p & ad4efe | !hbusreq4_p & adeaa4;
assign c3d5ec = hgrant1_p & v84554d | !hgrant1_p & c3d5eb;
assign bd5769 = hburst1 & v845542 | !hburst1 & c3d66b;
assign v8cc784 = hready_p & v8cc455 | !hready_p & v8cc783;
assign d35687 = hready_p & d3565e | !hready_p & d35632;
assign c3d2bd = hbusreq0 & v845564 | !hbusreq0 & v845542;
assign c3d2c5 = hburst0 & c3d2ad | !hburst0 & c3d2c4;
assign bd5876 = hgrant4_p & bd5757 | !hgrant4_p & bd5875;
assign ad45ea = hbusreq0 & ad45e5 | !hbusreq0 & ad45e9;
assign c3d399 = hlock0_p & v845542 | !hlock0_p & v84556e;
assign c3d708 = hmaster1_p & c3d707 | !hmaster1_p & c3d69b;
assign d354b4 = hlock4_p & v845542 | !hlock4_p & !d354b3;
assign v8cc5c0 = hlock2 & v8ccbd8 | !hlock2 & v8cc5bf;
assign v9e9ead = hmaster0_p & v9e9ea3 | !hmaster0_p & v9e9eac;
assign ad4ead = hlock1_p & ad4eab | !hlock1_p & !ad4eac;
assign d354bd = hmaster2_p & d35c00 | !hmaster2_p & !d354bc;
assign c3d5dd = hmaster2_p & c3d5dc | !hmaster2_p & v8da5a1;
assign b57ab8 = hready_p & b57a12 | !hready_p & b57ab7;
assign cc3707 = hbusreq2_p & cc36d5 | !hbusreq2_p & !cc3706;
assign cc36b9 = hmaster0_p & cc36b8 | !hmaster0_p & v845542;
assign v9ea40d = hmaster1_p & v9ea40c | !hmaster1_p & v845542;
assign d35756 = hmaster1_p & d35750 | !hmaster1_p & d35755;
assign b058ff = hbusreq3 & b058fd | !hbusreq3 & b058fe;
assign v9f77bb = hmaster0_p & v9f772d | !hmaster0_p & v9f772c;
assign bd5887 = hbusreq4_p & bd5884 | !hbusreq4_p & bd5886;
assign ade4d4 = hburst0 & c3d674 | !hburst0 & ade4d3;
assign bd576d = hbusreq3 & bd5768 | !hbusreq3 & !bd576c;
assign b57532 = decide_p & b57940 | !decide_p & b57a31;
assign b1cfc2 = hgrant4_p & v845542 | !hgrant4_p & !b1cfc1;
assign c3d5ba = hbusreq4_p & c3d5b8 | !hbusreq4_p & !c3d5b9;
assign d356df = hmaster0_p & d356da | !hmaster0_p & d356de;
assign d354d6 = hbusreq2 & d35c01 | !hbusreq2 & !v84555a;
assign ad4f59 = hbusreq3 & ad4f58 | !hbusreq3 & v845542;
assign b1cc00 = hbusreq4 & b1cbf6 | !hbusreq4 & b1cbff;
assign d35439 = hmaster1_p & d3542a | !hmaster1_p & d35438;
assign df5195 = hbusreq1_p & df5194 | !hbusreq1_p & v845542;
assign df51ca = decide_p & df51c9 | !decide_p & d6ebca;
assign b57436 = decide_p & b57982 | !decide_p & b57435;
assign c3d385 = decide_p & c3d2d5 | !decide_p & !c3d383;
assign v9ea484 = hbusreq1 & v9ea482 | !hbusreq1 & v9ea483;
assign c3d369 = hbusreq2 & v845564 | !hbusreq2 & v845542;
assign b579bc = hlock0 & b57942 | !hlock0 & b579bb;
assign ac146b = hgrant1_p & v845542 | !hgrant1_p & !ac146a;
assign v9ea5a9 = hbusreq2 & v9ea5a7 | !hbusreq2 & v9ea5a8;
assign v8cc0d6 = hbusreq2 & v8cc0d4 | !hbusreq2 & v8cc0d5;
assign c3ce1f = hmaster0_p & c3ce1e | !hmaster0_p & !c3d2be;
assign d358f6 = hmaster1_p & v845542 | !hmaster1_p & d358f5;
assign b579c6 = hbusreq3 & b579c4 | !hbusreq3 & b579c5;
assign c3d47d = hbusreq3 & c3d479 | !hbusreq3 & c3d47c;
assign c3d588 = hready_p & c3d586 | !hready_p & c3d587;
assign d35624 = hmaster2_p & dc5318 | !hmaster2_p & v845542;
assign d357b1 = hlock3_p & d357ab | !hlock3_p & d357b0;
assign d3599b = stateG10_4_p & d35997 | !stateG10_4_p & !d35999;
assign ad42c8 = hbusreq3 & ad42bf | !hbusreq3 & ad42c2;
assign c3d346 = hbusreq4 & c3d340 | !hbusreq4 & !c3d345;
assign dc4f93 = hmaster0_p & dc4f8c | !hmaster0_p & dc4f92;
assign ad439f = hmaster1_p & ad439e | !hmaster1_p & ad439b;
assign c5c934 = stateG10_4_p & v845542 | !stateG10_4_p & c5c933;
assign ade61c = hmaster0_p & ade61b | !hmaster0_p & ade5a8;
assign v9ea5a2 = hlock1 & v9ea59b | !hlock1 & v9ea5a1;
assign c5c966 = stateA1_p & c5c88b | !stateA1_p & v845542;
assign df5539 = hgrant1_p & df5538 | !hgrant1_p & !v845542;
assign ad42f1 = hlock1_p & ad42ef | !hlock1_p & ad42f0;
assign df54ee = hbusreq2_p & df54db | !hbusreq2_p & df54ed;
assign c3d748 = hgrant1_p & c3d6b6 | !hgrant1_p & c3d747;
assign v9ea616 = hbusreq2_p & v9ea610 | !hbusreq2_p & v9ea615;
assign d3543b = hmaster1_p & d3543a | !hmaster1_p & d35438;
assign v8cc4b1 = hmaster0_p & v8cc48d | !hmaster0_p & v8cc4b0;
assign c3d6e4 = hgrant4_p & c3d670 | !hgrant4_p & c3d6ab;
assign d35496 = hlock4_p & v845542 | !hlock4_p & !dc5300;
assign ad4611 = hready_p & ad45aa | !hready_p & ad4610;
assign dc500c = hbusreq4_p & dc5009 | !hbusreq4_p & dc500b;
assign ad460d = hready & ad457c | !hready & !v845542;
assign c5c89d = hlock0_p & c5c88d | !hlock0_p & !v845542;
assign ad5021 = hready & ad4fbe | !hready & !v845542;
assign c3d718 = hbusreq2_p & c3d711 | !hbusreq2_p & c3d717;
assign ad48c5 = hmaster0_p & ad5038 | !hmaster0_p & v845542;
assign b1c4c6 = hmaster2_p & d35a9c | !hmaster2_p & b1c4c5;
assign c5c939 = hgrant4_p & v845542 | !hgrant4_p & !c5c938;
assign b05a0e = hgrant1_p & b0593b | !hgrant1_p & b05a0d;
assign c3ce77 = hbusreq2 & c3ce75 | !hbusreq2 & c3ce37;
assign dc4fd1 = hbusreq3 & dc4fd0 | !hbusreq3 & v845542;
assign ad4400 = hmaster1_p & ad43ff | !hmaster1_p & ad43fc;
assign ad4156 = hbusreq4_p & ad4155 | !hbusreq4_p & ad4f3e;
assign ad480d = hbusreq3 & ad480c | !hbusreq3 & v845542;
assign ad4e7f = hmaster2_p & ad4e7e | !hmaster2_p & v845542;
assign bd58b1 = hbusreq1_p & dc4fcb | !hbusreq1_p & !v845542;
assign df51a4 = hbusreq3 & df518c | !hbusreq3 & !df518e;
assign v9f783e = hgrant4_p & d359c4 | !hgrant4_p & !v9f782a;
assign dc4f7e = hmaster2_p & dc4f7d | !hmaster2_p & ade4e1;
assign ad4f3c = hbusreq3 & ad4f3b | !hbusreq3 & v845542;
assign v9f7d0e = hbusreq3 & v9f7d0c | !hbusreq3 & v9f7d0d;
assign d356b7 = hbusreq3 & d356b6 | !hbusreq3 & d356ad;
assign ad4f90 = hbusreq4_p & ad4f8f | !hbusreq4_p & b1cfbe;
assign d35751 = hbusreq1_p & d35704 | !hbusreq1_p & d35aac;
assign b05a94 = hmaster1_p & b05a93 | !hmaster1_p & b05943;
assign d35982 = hbusreq2 & d35981 | !hbusreq2 & v845542;
assign ad4318 = hgrant1_p & v845542 | !hgrant1_p & ad4317;
assign d35596 = decide_p & d35595 | !decide_p & v84556c;
assign v9f7cee = hbusreq2 & v9f7cec | !hbusreq2 & v9f7ced;
assign v9f7cd4 = hlock2 & v9f7cd1 | !hlock2 & v9f7cd3;
assign ad42f0 = hbusreq1 & ad4e90 | !hbusreq1 & v845542;
assign ade4ee = hbusreq2 & ade4d6 | !hbusreq2 & ade4db;
assign ade56a = hbusreq1 & adec92 | !hbusreq1 & adec9c;
assign df517c = hgrant1_p & v84556c | !hgrant1_p & !df517b;
assign b5741d = hgrant4_p & v845542 | !hgrant4_p & b5741c;
assign d35980 = hmaster2_p & d3597f | !hmaster2_p & v845542;
assign bd592b = hbusreq2_p & bd592a | !hbusreq2_p & v845542;
assign c3d740 = hlock0_p & c3d6a5 | !hlock0_p & !c3d73f;
assign v9e9f80 = hbusreq1_p & v9e9f5d | !hbusreq1_p & v9e9f7f;
assign d3579a = hlock1_p & d35797 | !hlock1_p & d35799;
assign b05961 = hlock1 & b0595b | !hlock1 & b05960;
assign ad4606 = hlock3_p & ad45fe | !hlock3_p & ad4605;
assign v8cc759 = hgrant1_p & v845542 | !hgrant1_p & v8cc758;
assign d35a99 = hmaster2_p & d35a98 | !hmaster2_p & !v845542;
assign ad4ee8 = hmaster2_p & ad4ee2 | !hmaster2_p & ad4ee7;
assign df5172 = hbusreq1 & dc4fd0 | !hbusreq1 & v845542;
assign dc4fac = hbusreq4_p & dc4f7c | !hbusreq4_p & !v845542;
assign b05a9b = hbusreq3_p & b05a2c | !hbusreq3_p & b05a9a;
assign ade619 = hmaster1_p & ade618 | !hmaster1_p & ade5a4;
assign b57428 = hbusreq3 & b57426 | !hbusreq3 & b57427;
assign c5c3b7 = hgrant3_p & c5c8ee | !hgrant3_p & c5c3b6;
assign ad4f72 = hmaster2_p & ad4f6d | !hmaster2_p & ad4f71;
assign v9f7da7 = hbusreq4 & v9f7da5 | !hbusreq4 & v9f7da6;
assign b1c048 = hmaster0_p & b1c03f | !hmaster0_p & !b1c047;
assign c3d323 = hbusreq0 & c3d31f | !hbusreq0 & c3d322;
assign ac1479 = hbusreq4_p & ac1477 | !hbusreq4_p & !ac1478;
assign c3d5f1 = hbusreq0 & c3d5e0 | !hbusreq0 & c3d5f0;
assign v9f7684 = hmaster0_p & v9f7e2c | !hmaster0_p & v9f7683;
assign ad43cb = hmaster2_p & v845542 | !hmaster2_p & !ad43ca;
assign b57988 = hgrant1_p & v845542 | !hgrant1_p & b57987;
assign bd593b = hbusreq2_p & bd593a | !hbusreq2_p & !v845542;
assign c3d33b = hgrant0_p & v845542 | !hgrant0_p & !c3d2e8;
assign v9f7e22 = hlock4 & v9f7e1f | !hlock4 & v9f7e21;
assign ad4f87 = hbusreq4_p & ad4f86 | !hbusreq4_p & adeaa4;
assign b1cffd = hgrant1_p & v845542 | !hgrant1_p & b1cffc;
assign b1c71c = hbusreq0 & b1c71b | !hbusreq0 & v845542;
assign ad4f97 = hbusreq4_p & ad4f96 | !hbusreq4_p & ad4f88;
assign bd576c = hmaster2_p & v845542 | !hmaster2_p & bd576b;
assign d35987 = hbusreq2 & d35986 | !hbusreq2 & v845542;
assign c3cefc = hgrant2_p & v845551 | !hgrant2_p & c3cefb;
assign d35445 = hready_p & d35417 | !hready_p & d35444;
assign ad4806 = hbusreq3_p & ad4757 | !hbusreq3_p & !ad4805;
assign ad44b2 = stateG10_4_p & c3cec2 | !stateG10_4_p & !ad44b1;
assign c3d530 = hbusreq1_p & c3d480 | !hbusreq1_p & c3d52f;
assign c3d5ae = hbusreq2_p & c3d5ad | !hbusreq2_p & c3d38a;
assign b059b2 = hlock0 & b0595b | !hlock0 & b059b1;
assign v8cc5be = hlock3 & v8ccbd8 | !hlock3 & v8cc5bd;
assign dc4f98 = hbusreq2_p & dc4f84 | !hbusreq2_p & dc4f97;
assign ad4412 = hmaster0_p & ad440e | !hmaster0_p & ad4411;
assign v9e9f72 = hbusreq1_p & v9e9ee8 | !hbusreq1_p & v9e9f71;
assign c3d66e = locked_p & c3d66c | !locked_p & c3d66d;
assign d35501 = hmaster2_p & v845542 | !hmaster2_p & !d35a9b;
assign ad4708 = hmaster2_p & adec93 | !hmaster2_p & !ad4707;
assign d35a50 = hmaster2_p & v84556c | !hmaster2_p & !d35a4f;
assign d355a8 = locked_p & d355a7 | !locked_p & v845542;
assign c3cedb = hbusreq3_p & c3ceab | !hbusreq3_p & c3ceda;
assign ad3cdc = hmaster0_p & ad3cda | !hmaster0_p & ad3cdb;
assign ad5055 = hmaster2_p & ad5054 | !hmaster2_p & ad5044;
assign b5790a = hlock2_p & b57908 | !hlock2_p & b57909;
assign d35016 = hbusreq1_p & d357d0 | !hbusreq1_p & d357e9;
assign bd577b = hlock2_p & bd577a | !hlock2_p & !v845542;
assign c3d500 = hbusreq4 & c3d4fd | !hbusreq4 & !c3d4ff;
assign v8cc763 = hbusreq1 & v8cc482 | !hbusreq1 & v8ccbd8;
assign ade597 = hburst0 & v845542 | !hburst0 & ade596;
assign bd5908 = hlock1_p & bd5907 | !hlock1_p & df54d6;
assign v8cc7c0 = hmaster2_p & v8cc7bb | !hmaster2_p & v8cc7bf;
assign b1c563 = hmaster2_p & b1c858 | !hmaster2_p & b1c562;
assign ad3cd6 = hbusreq0 & ad3cd5 | !hbusreq0 & v845542;
assign v9f76fd = hgrant1_p & v9f7e08 | !hgrant1_p & v9f76fc;
assign d359f6 = hbusreq0_p & v845542 | !hbusreq0_p & d359f5;
assign v8cc5c7 = decide_p & v8ccbd7 | !decide_p & v8cc5c6;
assign ad42d4 = hmaster0_p & ad42d1 | !hmaster0_p & ad42d3;
assign v9ea494 = hbusreq1 & v9ea492 | !hbusreq1 & v9ea493;
assign df5179 = hmaster1_p & df5175 | !hmaster1_p & df5178;
assign ad4ef5 = hlock4_p & ad4ef4 | !hlock4_p & !ad4e9a;
assign v86cea1 = hmaster0_p & v8587b7 | !hmaster0_p & v84554c;
assign ad4f2f = hmaster0_p & ad4e93 | !hmaster0_p & ad4f2e;
assign c3d364 = decide_p & c3d359 | !decide_p & c3d362;
assign bd5b6d = hburst1 & bd5b6a | !hburst1 & bd5b6c;
assign v9ea410 = hgrant1_p & v845542 | !hgrant1_p & v9ea40f;
assign d359d6 = hgrant4_p & adeca0 | !hgrant4_p & v845542;
assign d35a20 = hmaster0_p & d35a1e | !hmaster0_p & d35a1f;
assign v9ea5dc = decide_p & v9ea5ca | !decide_p & v9ea5db;
assign d35527 = hbusreq4_p & d35516 | !hbusreq4_p & v84554a;
assign c3cee9 = hmaster0_p & c3cee8 | !hmaster0_p & !c3d2be;
assign b05a70 = hbusreq1 & b05a6e | !hbusreq1 & b05a6f;
assign df51b1 = decide_p & df51b0 | !decide_p & v845542;
assign ba7c80 = jx0_p & ba7c7f | !jx0_p & ba7c75;
assign ad435f = hmaster0_p & ad430c | !hmaster0_p & ad42ee;
assign ad4fec = hgrant1_p & ad4fb6 | !hgrant1_p & ad4feb;
assign ad43b8 = hbusreq0 & ad43b7 | !hbusreq0 & v845542;
assign ad460c = hmaster0_p & ad460a | !hmaster0_p & ad460b;
assign ad5046 = stateA1_p & c74b29 | !stateA1_p & !adea96;
assign bd589f = hmastlock_p & bd589e | !hmastlock_p & !v845542;
assign df51b5 = hmaster0_p & df51b2 | !hmaster0_p & df5169;
assign ad4ebd = hmaster2_p & ad4e79 | !hmaster2_p & ad4ebc;
assign b1c06d = stateG10_4_p & b1c062 | !stateG10_4_p & b1c06c;
assign v9f7e42 = hlock4 & v9f7e3f | !hlock4 & v9f7e41;
assign ad506b = hmaster1_p & ad506a | !hmaster1_p & ad501e;
assign v857440 = stateG3_0_p & v845542 | !stateG3_0_p & v93a916;
assign b57a77 = hbusreq0 & b57a76 | !hbusreq0 & b579ce;
assign d358f5 = hmaster0_p & d358f4 | !hmaster0_p & v845542;
assign c3d30c = hbusreq0 & c3d2ee | !hbusreq0 & c3d30b;
assign d35a42 = hgrant0_p & v845542 | !hgrant0_p & !d35a40;
assign b57958 = hmaster1_p & b5794b | !hmaster1_p & b57957;
assign ad13e3 = decide_p & ad13df | !decide_p & ad13e2;
assign b1c613 = hbusreq3_p & b1c5f8 | !hbusreq3_p & b1c612;
assign c3d738 = hmaster1_p & c3d737 | !hmaster1_p & c3d68b;
assign dc5316 = hbusreq4_p & adea88 | !hbusreq4_p & v845566;
assign c3d756 = hmaster0_p & c3d699 | !hmaster0_p & c3d696;
assign ad3d36 = hmaster0_p & ad4472 | !hmaster0_p & ad4433;
assign c3ce23 = decide_p & c3d5ae | !decide_p & !c3ce22;
assign ad4ea1 = hbusreq0 & ad4e9d | !hbusreq0 & ad4ea0;
assign d35954 = hburst1 & df54dd | !hburst1 & d3594c;
assign ad4f80 = hlock0_p & ad4f39 | !hlock0_p & !v845542;
assign b058dd = hlock3 & b058d5 | !hlock3 & b058dc;
assign v9ea604 = hbusreq1 & v9ea493 | !hbusreq1 & v9ea43b;
assign d3561d = hmastlock_p & d3561c | !hmastlock_p & v845542;
assign b05939 = locked_p & b05937 | !locked_p & !b05938;
assign dc53ba = hbusreq3 & dc53b8 | !hbusreq3 & dc53b9;
assign b1c4c4 = hmaster2_p & d35a9c | !hmaster2_p & !b1c4c3;
assign v9f7764 = hlock3 & v9f7763 | !hlock3 & v9f7761;
assign ad4ed3 = hlock4_p & ad4ed2 | !hlock4_p & v845542;
assign b574d0 = hmaster1_p & b579b4 | !hmaster1_p & b574cf;
assign ad4440 = hbusreq1_p & ad443f | !hbusreq1_p & ad40fe;
assign ad4287 = hlock1_p & ad4ecf | !hlock1_p & !v845542;
assign df51c6 = hmaster0_p & df51c4 | !hmaster0_p & df51c5;
assign df512e = hready_p & df512c | !hready_p & df512d;
assign d35694 = hmaster0_p & d35aaf | !hmaster0_p & d35693;
assign ad501e = hmaster0_p & ad501c | !hmaster0_p & ad501d;
assign bd58aa = stateG10_4_p & v84556c | !stateG10_4_p & !cc36ca;
assign bd57e7 = hmaster0_p & bd57e6 | !hmaster0_p & bd5797;
assign d35bf4 = hbusreq3 & d35bf3 | !hbusreq3 & d35be8;
assign b05a06 = hgrant0_p & b05939 | !hgrant0_p & !b05a05;
assign ad475f = hmaster1_p & ad475e | !hmaster1_p & ad45a5;
assign ade594 = hmaster2_p & adea94 | !hmaster2_p & ade593;
assign v9f770b = hmaster1_p & v9f7701 | !hmaster1_p & v9f770a;
assign c3ce79 = hbusreq1_p & c3ce3d | !hbusreq1_p & !c3d2de;
assign d35806 = hbusreq0_p & d3563c | !hbusreq0_p & v845542;
assign bd5b8d = hmaster1_p & bd5b8c | !hmaster1_p & v84556c;
assign bd580b = hgrant0_p & v84556c | !hgrant0_p & adec89;
assign c3ce7c = hbusreq2_p & c3ce40 | !hbusreq2_p & c3ce7b;
assign ade572 = locked_p & ade571 | !locked_p & v845542;
assign c3d319 = hgrant4_p & v845542 | !hgrant4_p & c3d318;
assign v9e9fc6 = hmaster1_p & v9e9fc5 | !hmaster1_p & v9e9ef1;
assign v8da5a1 = hbusreq4_p & v8da59f | !hbusreq4_p & !v8da5a0;
assign v8ccbf8 = hmaster1_p & v8ccbe5 | !hmaster1_p & v8ccbf7;
assign b05931 = hlock2_p & b0592f | !hlock2_p & b05930;
assign bd5b96 = hbusreq2 & df54f5 | !hbusreq2 & bd5b95;
assign v9f7714 = hgrant2_p & v9f7712 | !hgrant2_p & v9f7713;
assign b1c74e = stateA1_p & b1c74d | !stateA1_p & !v845542;
assign v9f7e34 = hbusreq0 & v9f7e30 | !hbusreq0 & v9f7e33;
assign bd5893 = hmaster2_p & bd588e | !hmaster2_p & bd5892;
assign b1c4cf = hmaster0_p & b1c842 | !hmaster0_p & b1c4ce;
assign v8cc127 = hbusreq2 & v8cc125 | !hbusreq2 & v8cc126;
assign ad43c7 = hmaster2_p & ad43c4 | !hmaster2_p & ad43c6;
assign c3d68f = hbusreq2_p & c3d68c | !hbusreq2_p & c3d68e;
assign bd5862 = hgrant0_p & ade589 | !hgrant0_p & adec89;
assign v9ea422 = hgrant4_p & v845542 | !hgrant4_p & v9ea421;
assign c3d5ac = hmaster1_p & c3d5a8 | !hmaster1_p & c3d5ab;
assign b574fc = hready_p & b5799c | !hready_p & b574fb;
assign dc5018 = hbusreq1 & dc4fce | !hbusreq1 & dc4fd0;
assign cc36ea = hmaster1_p & cc36df | !hmaster1_p & cc36e9;
assign c3d31e = hgrant4_p & v845542 | !hgrant4_p & !c3d318;
assign ad474e = hmaster0_p & ad4740 | !hmaster0_p & ad474d;
assign v9f77f1 = hbusreq4_p & v9f77ef | !hbusreq4_p & !v9f77f0;
assign b1cf2b = hmaster2_p & v845542 | !hmaster2_p & !v84554a;
assign b57a28 = hgrant1_p & v845542 | !hgrant1_p & b57a27;
assign ad4764 = hlock4_p & ad4dc4 | !hlock4_p & !ad4de2;
assign ad4568 = hbusreq4_p & ad4567 | !hbusreq4_p & v845542;
assign ade4f2 = decide_p & ade4f1 | !decide_p & v845542;
assign b57a8f = hgrant3_p & b57946 | !hgrant3_p & b57a8e;
assign b058ef = hready & b058ee | !hready & b058ea;
assign c3d66c = hmastlock_p & c3d66b | !hmastlock_p & !v845542;
assign ad42a5 = hbusreq1_p & ad42a4 | !hbusreq1_p & v845542;
assign ade5d4 = hbusreq1_p & ade5d3 | !hbusreq1_p & ade4dc;
assign b05a52 = hmaster0_p & b058c7 | !hmaster0_p & b058f6;
assign c3d2d9 = hready & v845542 | !hready & !v845564;
assign ad4e54 = locked_p & v845542 | !locked_p & ad4e53;
assign ad425c = decide_p & ad4165 | !decide_p & ad425b;
assign cc36e5 = stateG10_4_p & v845566 | !stateG10_4_p & !cc36e4;
assign d354fe = hbusreq4_p & d35c0b | !hbusreq4_p & !v845542;
assign d35575 = hmaster0_p & d35573 | !hmaster0_p & !d35574;
assign bd57a0 = hbusreq1 & bd579e | !hbusreq1 & bd579f;
assign dc4ff6 = hbusreq4_p & dc4ff3 | !hbusreq4_p & dc4ff5;
assign bd585c = hgrant4_p & ade589 | !hgrant4_p & adec89;
assign ade4f0 = hmaster1_p & ade4ef | !hmaster1_p & ade4ec;
assign dc5002 = hmaster2_p & dc4fe6 | !hmaster2_p & dc5001;
assign bd5935 = hbusreq0 & bd5934 | !hbusreq0 & v845542;
assign ade4b5 = decide_p & ade4b4 | !decide_p & v845542;
assign ad46af = hgrant1_p & ad4690 | !hgrant1_p & ad46ae;
assign bd574c = hmaster0_p & bd5748 | !hmaster0_p & bd574b;
assign c3d314 = hready & c3d310 | !hready & c3d313;
assign b1c78b = hbusreq2 & b1c71c | !hbusreq2 & b1c71d;
assign d357e3 = hbusreq2_p & d357e2 | !hbusreq2_p & d357e1;
assign v9f7cd7 = hbusreq0_p & v9f7cb4 | !hbusreq0_p & !v9f7c9f;
assign c3d512 = hready & c3d511 | !hready & !v845542;
assign c5c969 = hmaster2_p & c5c968 | !hmaster2_p & !v845542;
assign b1c076 = hgrant1_p & b1c060 | !hgrant1_p & b1c075;
assign dc4f8b = hbusreq1_p & dc4f8a | !hbusreq1_p & dc4f71;
assign ade620 = hbusreq2_p & ade61a | !hbusreq2_p & ade61f;
assign ad43c0 = hburst1_p & v84557e | !hburst1_p & !v845542;
assign b058ca = hlock3 & b058c9 | !hlock3 & b058c8;
assign v8cc132 = hbusreq3_p & v8cc122 | !hbusreq3_p & v8cc130;
assign v9f772d = hmaster2_p & v9f772b | !hmaster2_p & !v845542;
assign d354c2 = hmaster2_p & d354a4 | !hmaster2_p & d354c1;
assign v9ea4ce = hbusreq1_p & v9ea449 | !hbusreq1_p & v9ea4ca;
assign adea89 = hlock4_p & adea88 | !hlock4_p & !v845542;
assign b5798b = hgrant2_p & b57948 | !hgrant2_p & b5798a;
assign v9ea4a7 = hmaster2_p & v9f20a1 | !hmaster2_p & v9ea4a6;
assign v9e9f4e = hbusreq0_p & v9e9f4d | !hbusreq0_p & v9ea441;
assign df51a7 = hbusreq3 & df5192 | !hbusreq3 & !v84554c;
assign v9f771a = hmaster1_p & v9f7719 | !hmaster1_p & v9f76a6;
assign v9f7664 = hgrant4_p & v9f7cdc | !hgrant4_p & v9f7663;
assign dc507a = hbusreq1 & dc5070 | !hbusreq1 & !v845542;
assign b05a2e = hmaster1_p & b05a2d | !hmaster1_p & b05913;
assign dc53d2 = jx1_p & dc53ca | !jx1_p & dc53d1;
assign d3594a = hburst0_p & v845542 | !hburst0_p & d35949;
assign v9ea40b = hready_p & v9ea3e3 | !hready_p & v9ea40a;
assign v9f7dc6 = hlock1_p & v9f7ce4 | !hlock1_p & !v9f7d2a;
assign v9ea61e = hlock2_p & v9ea61b | !hlock2_p & v9ea61d;
assign df515b = hbusreq2 & df5157 | !hbusreq2 & df5159;
assign d3542b = hbusreq1 & d35421 | !hbusreq1 & d35425;
assign v8cc810 = hbusreq2 & v8cc80d | !hbusreq2 & v8cc80f;
assign d358ed = hmastlock_p & d358ec | !hmastlock_p & v845542;
assign c3cf03 = hready & c3cf02 | !hready & !v845542;
assign d359a9 = hbusreq0 & d359a8 | !hbusreq0 & v845542;
assign ad4dad = hlock0_p & dc4f78 | !hlock0_p & !v845542;
assign b0592b = hmaster0_p & b0591d | !hmaster0_p & b05920;
assign v9f768e = stateG10_4_p & v9f768c | !stateG10_4_p & v9f768d;
assign ad3d4a = hbusreq2_p & ad3d45 | !hbusreq2_p & ad3d49;
assign c3ce71 = hgrant2_p & c3d36c | !hgrant2_p & c3ce70;
assign b1c05f = hbusreq1 & b1c807 | !hbusreq1 & !b1c809;
assign b1c73a = hbusreq3 & b1c739 | !hbusreq3 & !v845542;
assign bd5916 = hlock1_p & bd5914 | !hlock1_p & bd5915;
assign bd5892 = hbusreq4_p & bd588f | !hbusreq4_p & bd5891;
assign bd5e29 = hready_p & v845542 | !hready_p & bd5e26;
assign ad40e6 = hbusreq2 & ad4df0 | !hbusreq2 & v845542;
assign v9f77fd = hlock2 & v9f77fa | !hlock2 & v9f77fc;
assign ad4490 = hbusreq1_p & ad43a9 | !hbusreq1_p & ad448f;
assign c3ce3a = hmaster0_p & c3ce38 | !hmaster0_p & c3ce39;
assign ad4e98 = hlock0_p & v84556c | !hlock0_p & !v845542;
assign v9f7d7c = hlock4_p & v9f7d7a | !hlock4_p & !v9f7d7b;
assign v8cc4af = hlock2 & v8cc4ad | !hlock2 & v8cc4ae;
assign ad426d = hbusreq1 & ad4f40 | !hbusreq1 & v845542;
assign bd58d5 = hbusreq2 & bd58d4 | !hbusreq2 & v845542;
assign ade4b9 = busreq_p & v845542 | !busreq_p & !ade4b8;
assign ad4810 = hready & v845542 | !hready & v84556c;
assign ade5a7 = hbusreq2 & ade548 | !hbusreq2 & !v845558;
assign v9f7668 = hlock0 & v9f7667 | !hlock0 & v9f765c;
assign bd5869 = hbusreq4_p & bd5866 | !hbusreq4_p & bd5868;
assign v9e9f56 = hbusreq4_p & v9e9f54 | !hbusreq4_p & v9e9f55;
assign v9f77ca = hbusreq0 & v9f77c2 | !hbusreq0 & v9f77c9;
assign df51a0 = decide_p & df519f | !decide_p & d6ebca;
assign v9f7cff = hbusreq1 & v9f7cfd | !hbusreq1 & v9f7cfe;
assign b5794c = hlock1_p & b578f1 | !hlock1_p & v845542;
assign d35a12 = hbusreq4_p & d35a0c | !hbusreq4_p & v845542;
assign b05984 = stateG10_4_p & b05980 | !stateG10_4_p & !b05982;
assign ac147e = hgrant2_p & ac1456 | !hgrant2_p & ac147d;
assign b1cfb7 = hgrant4_p & v845542 | !hgrant4_p & !b1cfb6;
assign b57414 = hbusreq3 & b57412 | !hbusreq3 & b57413;
assign c3ce26 = hbusreq2_p & c3d5ad | !hbusreq2_p & c3d391;
assign b1c586 = decide_p & b1c585 | !decide_p & b1d013;
assign b1c04b = decide_p & b1c04a | !decide_p & !v845542;
assign ad5066 = hmaster0_p & ad5039 | !hmaster0_p & ad5065;
assign bd57bb = hburst1_p & v8f2540 | !hburst1_p & !v845568;
assign v9e9f7d = hready & v9e9f7c | !hready & v9e9f79;
assign b57abb = hgrant3_p & b57ab8 | !hgrant3_p & b57aba;
assign dc4f64 = decide_p & dc4f63 | !decide_p & v845542;
assign v9e9ed8 = hgrant3_p & v9e9ecb | !hgrant3_p & v9e9ed7;
assign v8cc0da = hmaster2_p & v8cc0d9 | !hmaster2_p & v8cc493;
assign d3590e = hmaster2_p & d35909 | !hmaster2_p & d3590d;
assign c3d6bb = stateG10_4_p & c3d6b8 | !stateG10_4_p & c3d6ba;
assign c3d484 = hready_p & v845555 | !hready_p & c3d483;
assign ad3ce6 = hbusreq0 & ad3ce3 | !hbusreq0 & v845564;
assign v9ea58f = hbusreq1_p & v9ea3fa | !hbusreq1_p & v9ea58e;
assign v9f7e2a = hbusreq3 & v9f7e27 | !hbusreq3 & v9f7e29;
assign b1c803 = hbusreq1_p & b1c7b5 | !hbusreq1_p & b1c802;
assign c3d75d = hmaster1_p & c3d714 | !hmaster1_p & c3d70f;
assign v8d2b2e = hgrant0_p & v845542 | !hgrant0_p & v8d2b2b;
assign v9f76c8 = hbusreq1_p & v9f7d3d | !hbusreq1_p & v9f76c6;
assign v9f7ccb = hlock4 & v9f7cc8 | !hlock4 & v9f7cca;
assign b1c869 = hready_p & b1c867 | !hready_p & b1c868;
assign b1cfcd = stateG10_4_p & b1cfcb | !stateG10_4_p & !b1cfcc;
assign d359b8 = hmaster2_p & d3597f | !hmaster2_p & d359b7;
assign b578fa = hmaster2_p & b578f9 | !hmaster2_p & v845542;
assign ad3d35 = hmaster1_p & ad3d34 | !hmaster1_p & ad4425;
assign ad4ff6 = hbusreq3 & ad4ff5 | !hbusreq3 & v845542;
assign b1c4a3 = hlock0_p & d3594e | !hlock0_p & v845542;
assign v9f7782 = hmaster1_p & v9f7781 | !hmaster1_p & v9f776d;
assign d3563f = hlock0_p & d3563d | !hlock0_p & !d3563e;
assign dc53c1 = hbusreq3 & dc53bf | !hbusreq3 & dc53c0;
assign d355a6 = hmastlock_p & v8cc792 | !hmastlock_p & d355a5;
assign v9f76cd = hmaster1_p & v9f76cc | !hmaster1_p & v9f7d64;
assign ad419d = hbusreq2 & v845542 | !hbusreq2 & c3d2d9;
assign b059cc = hbusreq1_p & b059b8 | !hbusreq1_p & b0596b;
assign v9e9ed1 = hmaster0_p & v9e9e79 | !hmaster0_p & v9e9eb5;
assign b05a20 = hmaster0_p & b05a16 | !hmaster0_p & !b05a1f;
assign d35919 = hmaster2_p & adea8a | !hmaster2_p & d35918;
assign c5c9b6 = hbusreq3_p & c5c99d | !hbusreq3_p & c5c9b5;
assign ad4e5c = hlock0_p & v845542 | !hlock0_p & ad4e5b;
assign ade4bc = stateA1_p & ade4b9 | !stateA1_p & !ade4bb;
assign d359fb = stateG10_4_p & d359f7 | !stateG10_4_p & d359f9;
assign ad40f1 = hlock3_p & ad40ea | !hlock3_p & ad40f0;
assign ad4778 = hlock4_p & ad4dce | !hlock4_p & !v845542;
assign dc4fd3 = hmaster0_p & dc4fcd | !hmaster0_p & dc4fd2;
assign ad42ff = hbusreq2 & ad4287 | !hbusreq2 & v845542;
assign df5143 = hbusreq3 & df5141 | !hbusreq3 & df5142;
assign v8cc47b = hmaster2_p & v845542 | !hmaster2_p & v8cc47a;
assign ad458f = hready & ad458e | !hready & !v845542;
assign ade56c = hburst0 & v889629 | !hburst0 & ade56b;
assign b05903 = hbusreq1_p & b058fd | !hbusreq1_p & b058c7;
assign v9f77ae = hlock0_p & v845542 | !hlock0_p & v9f77ad;
assign v9f7c9d = hmastlock_p & c6d44d | !hmastlock_p & v845542;
assign v8cc798 = hlock0 & v8ccb6b | !hlock0 & v8cc797;
assign b1c778 = hmaster0_p & b1c75d | !hmaster0_p & b1c777;
assign v9f7d62 = hlock0_p & v9ea3fb | !hlock0_p & v9f7d61;
assign d357ef = hmaster1_p & d357ea | !hmaster1_p & d357ee;
assign ad3d54 = hmaster0_p & ad4413 | !hmaster0_p & ad3d15;
assign dc53c6 = hready_p & dc53be | !hready_p & !dc53c5;
assign bd591d = hbusreq2_p & bd591c | !hbusreq2_p & !v845542;
assign d35a35 = hgrant2_p & d35a2b | !hgrant2_p & !d35a34;
assign ad4e4a = hbusreq3 & ad4e49 | !hbusreq3 & v845542;
assign df51c2 = hmaster1_p & df51c1 | !hmaster1_p & df5197;
assign v9f76f2 = hmaster2_p & v9f76f1 | !hmaster2_p & v9f7db3;
assign c5c8f4 = hmaster2_p & c5c8f3 | !hmaster2_p & v845542;
assign dc5082 = decide_p & dc5081 | !decide_p & v845542;
assign b57b5c = jx0_p & b57a35 | !jx0_p & b57b5b;
assign b579db = hlock0 & b579d9 | !hlock0 & b579da;
assign d3570b = hmaster0_p & d35706 | !hmaster0_p & d3570a;
assign v9f7ce1 = hbusreq4 & v9f7cdf | !hbusreq4 & v9f7ce0;
assign c3d2c8 = hbusreq3 & c3d2c7 | !hbusreq3 & !v845542;
assign b579cc = hgrant0_p & b57941 | !hgrant0_p & v845542;
assign ad4fa7 = hmaster1_p & ad4fa6 | !hmaster1_p & ad4f9e;
assign b1c80f = hmaster2_p & b1c741 | !hmaster2_p & d35a9c;
assign ad472f = hready & ad472e | !hready & !v845542;
assign d3557d = hbusreq4_p & d354a5 | !hbusreq4_p & !d35aab;
assign adea8a = hbusreq4_p & adea89 | !hbusreq4_p & !v845542;
assign dc5017 = hmaster0_p & dc4ffb | !hmaster0_p & dc5016;
assign v8f2540 = start_p & v845542 | !start_p & v857b36;
assign v9f76d4 = hmaster1_p & v9f76d3 | !hmaster1_p & v9f7ce9;
assign d35aad = hbusreq1_p & v845542 | !hbusreq1_p & d35aac;
assign v9f784c = hbusreq3 & v9f7849 | !hbusreq3 & v9f784b;
assign d35a59 = hgrant4_p & d35a58 | !hgrant4_p & ade563;
assign dc531d = hmaster1_p & dc531c | !hmaster1_p & v845542;
assign b1cff5 = hlock0_p & b1cff4 | !hlock0_p & !v845542;
assign df51d5 = hready_p & v845542 | !hready_p & df51d4;
assign ad4430 = hbusreq0 & ad4e8e | !hbusreq0 & v845542;
assign ad4696 = hbusreq0 & ad4693 | !hbusreq0 & ad4695;
assign c3cf0b = hmaster0_p & c3cf09 | !hmaster0_p & c3cf0a;
assign b05a4d = hmaster0_p & b058c7 | !hmaster0_p & b058b5;
assign b05a3d = hbusreq0_p & b0591c | !hbusreq0_p & b05938;
assign b1cfc9 = hgrant1_p & v845542 | !hgrant1_p & b1cfc8;
assign c3d5a8 = hmaster0_p & c3d5a6 | !hmaster0_p & c3d5a7;
assign d35645 = hgrant1_p & df54f3 | !hgrant1_p & d35644;
assign ad4487 = hready & ad4484 | !hready & ad4486;
assign v8cc491 = hbusreq4_p & v8cc48e | !hbusreq4_p & v8cc48f;
assign b1c780 = hmaster0_p & b1c77f | !hmaster0_p & b1c75e;
assign bd5858 = hbusreq1 & bd5758 | !hbusreq1 & v84556c;
assign c3d2e6 = hmastlock_p & c3d2e5 | !hmastlock_p & v845542;
assign ad46eb = hbusreq2 & ad458f | !hbusreq2 & v845542;
assign b1c843 = hlock0_p & v845566 | !hlock0_p & v845542;
assign ad4dd3 = hbusreq4 & ad4dd0 | !hbusreq4 & !ad4dd2;
assign d354a0 = hbusreq1 & d35c01 | !hbusreq1 & !v84555a;
assign ade58b = hgrant0_p & ade56d | !hgrant0_p & !v84556c;
assign v9f76af = hbusreq2_p & v9f76a8 | !hbusreq2_p & v9f76ae;
assign ad40f7 = hmaster0_p & ad40f5 | !hmaster0_p & ad40f6;
assign d354ee = hbusreq3 & d354bd | !hbusreq3 & !v84555a;
assign ade4af = hmaster0_p & ade4a8 | !hmaster0_p & ade4ae;
assign b1c715 = hbusreq0_p & df513b | !hbusreq0_p & v845542;
assign ad46a1 = hlock4_p & ad4e8c | !hlock4_p & v845542;
assign c3d691 = decide_p & c3d690 | !decide_p & c3d680;
assign ad4d92 = hmaster2_p & ad4d91 | !hmaster2_p & v845542;
assign v9ea5e0 = hmaster0_p & v9ea5b4 | !hmaster0_p & v9ea44a;
assign c3cf10 = hmaster1_p & c3cf0b | !hmaster1_p & c3cf0f;
assign v9ea437 = stateA1_p & v9ea3e5 | !stateA1_p & v845542;
assign ad433e = hbusreq1_p & ad433d | !hbusreq1_p & v845542;
assign c3d50f = hbusreq4_p & c3d374 | !hbusreq4_p & v845542;
assign d3575b = hgrant3_p & d3573c | !hgrant3_p & !d3575a;
assign ad4732 = hready & ad4702 | !hready & !ad4731;
assign bd5ea0 = hbusreq4_p & bd5b93 | !hbusreq4_p & !v845542;
assign ad45fb = hmaster0_p & ad45c1 | !hmaster0_p & ad45fa;
assign ade4a8 = hbusreq3 & ade4a7 | !hbusreq3 & adec93;
assign b058f7 = hlock0 & b058b8 | !hlock0 & b058c7;
assign b1c093 = hmaster0_p & b1cfb8 | !hmaster0_p & b1cfd1;
assign b57a1f = hmaster0_p & b57a1e | !hmaster0_p & b57900;
assign v9f7653 = hgrant4_p & v9f7e2f | !hgrant4_p & !v9f7c9f;
assign d35494 = hbusreq4_p & d35493 | !hbusreq4_p & v845542;
assign ad4336 = hbusreq2 & ad4331 | !hbusreq2 & ad4334;
assign ad3d1e = hbusreq2_p & ad3d14 | !hbusreq2_p & ad3d1d;
assign cc36dd = hbusreq4_p & cc36db | !hbusreq4_p & cc36dc;
assign ad4362 = hbusreq2 & ad4f1e | !hbusreq2 & !v845542;
assign b57a34 = hgrant3_p & b57a23 | !hgrant3_p & b57a33;
assign ad41a9 = hgrant2_p & ad41a0 | !hgrant2_p & ad41a8;
assign bd5910 = hready_p & v845542 | !hready_p & bd590f;
assign df5139 = hbusreq1_p & df5138 | !hbusreq1_p & v845542;
assign v9ea626 = hbusreq2_p & v9ea625 | !hbusreq2_p & v9ea4c0;
assign ad4f9b = hready & ad4f7d | !hready & ad4f9a;
assign df5534 = hgrant1_p & df5533 | !hgrant1_p & !v845542;
assign ad432f = hbusreq1 & ad5026 | !hbusreq1 & v845547;
assign b1c567 = hbusreq4 & b1c561 | !hbusreq4 & b1c566;
assign v9f7787 = hlock0 & v9f772c | !hlock0 & v9f7786;
assign c3d704 = hgrant2_p & c3d700 | !hgrant2_p & c3d703;
assign v9ea5b4 = hgrant1_p & v9ea581 | !hgrant1_p & v9ea591;
assign v8cc7bd = hlock0_p & v8cc7bc | !hlock0_p & v845542;
assign b05a7d = hlock3 & b05a7c | !hlock3 & b05a7a;
assign b1c76f = hbusreq0 & b1c76e | !hbusreq0 & b1cf2b;
assign ade4b4 = hbusreq2_p & ade4b0 | !hbusreq2_p & ade4b3;
assign d35640 = hgrant4_p & v84556c | !hgrant4_p & d3563f;
assign ad4369 = hmaster1_p & ad430c | !hmaster1_p & ad42f9;
assign ad45f1 = hmaster2_p & v845542 | !hmaster2_p & !ad45f0;
assign c3d595 = hbusreq2 & c3d58f | !hbusreq2 & !v845542;
assign v8cc813 = hmaster1_p & v8cc812 | !hmaster1_p & v845542;
assign ad3d3e = hmaster1_p & ad4472 | !hmaster1_p & ad4469;
assign v9f7761 = hbusreq1_p & v9f7758 | !hbusreq1_p & v9f7760;
assign c3d4e0 = hlock4_p & c3d308 | !hlock4_p & v8da59f;
assign b57900 = hmaster2_p & b578fe | !hmaster2_p & b578ff;
assign ad44b6 = hready & ad44a8 | !hready & ad44b5;
assign ad4262 = jx1_p & ad4806 | !jx1_p & ad4261;
assign b5742e = hlock3 & b578f1 | !hlock3 & b57410;
assign dc4fb3 = hmaster1_p & dc4fa1 | !hmaster1_p & dc4fb2;
assign b1c5e0 = hbusreq2 & b1cfc9 | !hbusreq2 & b1cfd1;
assign b578f3 = hmaster1_p & b578f2 | !hmaster1_p & v845542;
assign d35426 = hbusreq3 & d35421 | !hbusreq3 & d35425;
assign v8ccbf2 = hlock0_p & v8ccbf0 | !hlock0_p & v845542;
assign v9f7d37 = hbusreq2_p & v9f7d30 | !hbusreq2_p & v9f7d36;
assign ad443e = hgrant1_p & ad4436 | !hgrant1_p & ad443d;
assign c3ceb4 = hbusreq1 & c3cead | !hbusreq1 & c3ceaf;
assign ad3ced = stateG10_4_p & ad3ceb | !stateG10_4_p & ad3cec;
assign v9ea421 = hlock0_p & v9ea41c | !hlock0_p & v9ea420;
assign b05a35 = hmaster1_p & b05a34 | !hmaster1_p & b058e1;
assign ad45a8 = hmaster1_p & ad45a7 | !hmaster1_p & ad45a5;
assign v9f776e = hmaster1_p & v9f774f | !hmaster1_p & v9f776d;
assign v9f7683 = hbusreq2 & v9f7681 | !hbusreq2 & v9f7682;
assign v8cc7a8 = decide_p & v8cc7a7 | !decide_p & v8cc7a6;
assign v8cc48f = stateG10_4_p & v845542 | !stateG10_4_p & v8cc48e;
assign dc5075 = hbusreq2 & dc5074 | !hbusreq2 & !v845542;
assign ad448f = hready & ad448b | !hready & ad448e;
assign cc36ed = hready_p & cc36d7 | !hready_p & cc36ec;
assign ad40eb = hbusreq2 & ad4da1 | !hbusreq2 & v845542;
assign v9e9eac = hbusreq2 & v9e9eaa | !hbusreq2 & v9e9eab;
assign b57a8c = hbusreq2_p & b57a83 | !hbusreq2_p & b57a8b;
assign adec91 = hbusreq4_p & adec90 | !hbusreq4_p & v845542;
assign d359b1 = hgrant1_p & d359b0 | !hgrant1_p & d359aa;
assign c5c8ed = decide_p & c5c8e1 | !decide_p & c5c8ec;
assign v9f7871 = hmaster0_p & v9f7870 | !hmaster0_p & v9f776c;
assign v9ea4b8 = hbusreq1_p & v9ea3fc | !hbusreq1_p & v9ea4b7;
assign v9ea612 = hmaster1_p & v9ea611 | !hmaster1_p & v9ea4bd;
assign v9f7dad = hgrant0_p & v9f7cc7 | !hgrant0_p & v9f7cc6;
assign d35a19 = hgrant1_p & d359ec | !hgrant1_p & d35a18;
assign ad4294 = hmaster0_p & ad4291 | !hmaster0_p & ad4293;
assign d356e6 = hmaster1_p & d356df | !hmaster1_p & d356e5;
assign b0593b = hmaster2_p & b05939 | !hmaster2_p & !v9ea463;
assign c3ce91 = hmaster1_p & c3ce8e | !hmaster1_p & c3ce90;
assign d35a9a = hbusreq1_p & v845542 | !hbusreq1_p & d35a99;
assign d357b6 = hlock0_p & v845542 | !hlock0_p & adea9a;
assign ad4f0c = hgrant4_p & adea98 | !hgrant4_p & v845542;
assign bd584a = hgrant4_p & v845542 | !hgrant4_p & !bd574e;
assign d356c3 = hbusreq3 & d356c0 | !hbusreq3 & !v84554e;
assign v9f7894 = hgrant1_p & v9f77d6 | !hgrant1_p & v9f7893;
assign df513e = hbusreq1_p & df513d | !hbusreq1_p & v845542;
assign v9f7855 = hgrant3_p & v9f77ba | !hgrant3_p & v9f7854;
assign ade657 = decide_p & ade656 | !decide_p & v845542;
assign ad42af = hbusreq1 & ad4db7 | !hbusreq1 & v845542;
assign v9f7728 = hmaster1_p & d35aaa | !hmaster1_p & v9f7727;
assign dc501e = stateG10_4_p & adeca1 | !stateG10_4_p & !dc501d;
assign df5165 = hbusreq1 & dc4f6f | !hbusreq1 & v845542;
assign c3cee7 = hmaster0_p & c3cee5 | !hmaster0_p & c3cee6;
assign c5c8ff = hmaster2_p & c5c8fb | !hmaster2_p & !c5c8fe;
assign d3558c = hmaster2_p & d35aac | !hmaster2_p & d3558b;
assign ad47fa = hmaster0_p & ad4720 | !hmaster0_p & ad4706;
assign c3ce2c = hbusreq2_p & c3cdfd | !hbusreq2_p & c3ce2b;
assign cc36bc = decide_p & cc36bb | !decide_p & v84556c;
assign b57904 = hmaster1_p & b57903 | !hmaster1_p & b57901;
assign d359a6 = stateG10_4_p & d35997 | !stateG10_4_p & d359a5;
assign d354dc = hmaster1_p & d354d8 | !hmaster1_p & d354db;
assign d356ca = hmaster1_p & d356c4 | !hmaster1_p & d356c9;
assign ad4105 = hgrant1_p & ad40ff | !hgrant1_p & ad4104;
assign df51b8 = decide_p & df51b7 | !decide_p & v845542;
assign bd5ba9 = hbusreq2 & v84556c | !hbusreq2 & v845542;
assign d35578 = hbusreq1_p & d354e4 | !hbusreq1_p & !d35577;
assign bd588a = hgrant4_p & bd576b | !hgrant4_p & !bd580d;
assign b1c57f = hmaster2_p & d35a9c | !hmaster2_p & b1c57e;
assign v9f7862 = hbusreq4 & v9f7860 | !hbusreq4 & v9f7861;
assign ade586 = hgrant0_p & adec90 | !hgrant0_p & v84556c;
assign c3d30e = hmaster2_p & c3d2f7 | !hmaster2_p & c3d30d;
assign c3d744 = hmaster2_p & c3d743 | !hmaster2_p & c3d6bc;
assign df50d8 = hbusreq1 & dc5317 | !hbusreq1 & df50d7;
assign df54e7 = hlock1_p & df54e6 | !hlock1_p & v845542;
assign jx2 = aa4260;
assign ad471b = hmaster0_p & ad4710 | !hmaster0_p & ad471a;
assign df518b = hbusreq1 & dc5019 | !hbusreq1 & v845542;
assign d359eb = hlock1_p & d359e5 | !hlock1_p & d359ea;
assign d355ab = hmaster0_p & d355aa | !hmaster0_p & dc4fcb;
assign v9f7707 = hbusreq3 & v9f7703 | !hbusreq3 & v9f7706;
assign b1c762 = hbusreq0 & b1c761 | !hbusreq0 & !v845542;
assign ad4d97 = hmaster2_p & v845542 | !hmaster2_p & !dc4f78;
assign d359d0 = hgrant4_p & adeca0 | !hgrant4_p & d359ce;
assign ad428e = hbusreq2_p & ad428a | !hbusreq2_p & ad428d;
assign ac1453 = decide_p & ac1452 | !decide_p & ac1451;
assign c3d698 = hmaster0_p & c3d696 | !hmaster0_p & c3d697;
assign ad4459 = hmaster2_p & ad4458 | !hmaster2_p & v845542;
assign b1d00d = hlock3_p & b1cfd5 | !hlock3_p & b1d007;
assign c5c8e5 = stateA1_p & c5c88b | !stateA1_p & c5c8e4;
assign b1d005 = hmaster0_p & b1cfb8 | !hmaster0_p & b1d004;
assign v9e9f6c = hbusreq0 & v9e9f6b | !hbusreq0 & v9e9f68;
assign c3ce61 = hgrant1_p & c3ce5e | !hgrant1_p & c3ce60;
assign ad4dc5 = hmaster2_p & v845542 | !hmaster2_p & ad4dc4;
assign ad4fce = locked_p & ad4fcd | !locked_p & v845542;
assign v9f78a4 = hmaster1_p & v9f78a3 | !hmaster1_p & v9f77b0;
assign ade5db = hmaster0_p & ade5c9 | !hmaster0_p & ade4ee;
assign c3d392 = hbusreq2_p & c3d38a | !hbusreq2_p & c3d391;
assign c3d3aa = decide_p & c3d3a9 | !decide_p & c3d398;
assign d35a29 = hbusreq2 & d359ca | !hbusreq2 & !v845542;
assign v9ea5ba = hready_p & v9ea436 | !hready_p & v9ea5b9;
assign ad5019 = hbusreq3 & ad5018 | !hbusreq3 & c3d2d9;
assign v9fa31b = stateG3_0_p & v845542 | !stateG3_0_p & v845582;
assign b57a79 = hready & b57a78 | !hready & b579ce;
assign b1c6fa = hmaster0_p & b1c85a | !hmaster0_p & b1c6f9;
assign v9f7d20 = hbusreq4_p & v9ea3ec | !hbusreq4_p & !v9f7cc6;
assign v9f774c = hlock3 & v9f7745 | !hlock3 & v9f774b;
assign d358fd = hbusreq1_p & d358fc | !hbusreq1_p & v845542;
assign v9f7dbf = hbusreq1_p & v9f7dbe | !hbusreq1_p & v9f7da3;
assign b1c498 = hbusreq0 & b1caea | !hbusreq0 & b1c497;
assign dc5087 = hgrant3_p & dc4fc8 | !hgrant3_p & !dc5086;
assign c3d57f = hready & c3d57e | !hready & c3d4f6;
assign b1c80a = hbusreq1_p & v845542 | !hbusreq1_p & b1c809;
assign c3d763 = hbusreq3_p & c3d71b | !hbusreq3_p & !c3d762;
assign bd5b9f = decide_p & bd5b7c | !decide_p & !v845572;
assign v8cc825 = hbusreq3 & v8cc821 | !hbusreq3 & v8cc822;
assign dc502d = hbusreq4 & dc5026 | !hbusreq4 & dc502c;
assign v9f7721 = decide_p & v9f76cb | !decide_p & !v9f7720;
assign ad4e85 = hgrant4_p & v84556c | !hgrant4_p & b1cfcb;
assign ad4e49 = hready & ad4e48 | !hready & df54f5;
assign b1cf32 = hbusreq0 & b1cf25 | !hbusreq0 & b1cf31;
assign df507a = hbusreq1_p & df5079 | !hbusreq1_p & v845542;
assign ad4739 = hbusreq4 & ad4738 | !hbusreq4 & v845542;
assign bd5b79 = hmaster1_p & bd5b78 | !hmaster1_p & v845542;
assign c3d582 = hmaster0_p & c3d581 | !hmaster0_p & c3d505;
assign c3ced4 = hmaster1_p & c3ced2 | !hmaster1_p & c3ced3;
assign cc36ff = hgrant4_p & v845542 | !hgrant4_p & !cc36fe;
assign v9f7e1e = hbusreq4_p & v9f7e1c | !hbusreq4_p & v9f7e1d;
assign d3573b = decide_p & d3573a | !decide_p & v84556c;
assign b57503 = decide_p & b57a21 | !decide_p & b57502;
assign v9e9f8e = hmaster2_p & v9e9f8d | !hmaster2_p & v9ea4d8;
assign ad4757 = hgrant3_p & ad4611 | !hgrant3_p & ad4756;
assign bd5848 = hbusreq0 & bd583f | !hbusreq0 & bd5847;
assign v9f76b4 = hmaster1_p & v9f76b3 | !hmaster1_p & v9f7d2f;
assign v9ea4a4 = decide_p & v9ea4a3 | !decide_p & v9ea3e3;
assign ad505b = hbusreq4_p & v845542 | !hbusreq4_p & !ad505a;
assign b1cf28 = hbusreq0 & b1cf25 | !hbusreq0 & b1cf27;
assign b05956 = hgrant4_p & v9f7d42 | !hgrant4_p & b05954;
assign b1c4c3 = hbusreq4_p & b1cf24 | !hbusreq4_p & b1c843;
assign ade650 = hready_p & ade64e | !hready_p & ade64f;
assign d356d3 = hlock1_p & v845542 | !hlock1_p & d356d2;
assign v9f7da4 = hlock0 & v9f7da3 | !hlock0 & v9f7cf6;
assign b1caf7 = hmaster2_p & v845542 | !hmaster2_p & b1caf6;
assign v8cc633 = decide_p & v8cc4f4 | !decide_p & v8cc630;
assign v8cc7b6 = hlock2 & v8ccbe8 | !hlock2 & v8cc7b5;
assign b1c721 = hmaster2_p & b1c70f | !hmaster2_p & b1c720;
assign v9f7693 = hbusreq1_p & v9f7d5a | !hbusreq1_p & v9f7692;
assign b1c709 = hgrant3_p & b1c705 | !hgrant3_p & b1c708;
assign b1c5ff = hbusreq2_p & b1c5f2 | !hbusreq2_p & b1c864;
assign c3d5e6 = hgrant1_p & v84554d | !hgrant1_p & c3d5e5;
assign d359de = hbusreq4_p & d359dc | !hbusreq4_p & d359dd;
assign c3d6c7 = hgrant0_p & c3d66e | !hgrant0_p & c3d66d;
assign d35a0d = hbusreq4_p & d35a0c | !hbusreq4_p & d359dd;
assign v9f7cb2 = hbusreq2 & v9f7cb0 | !hbusreq2 & v9f7cb1;
assign d356ad = hbusreq1_p & d356ac | !hbusreq1_p & v845542;
assign cc36c0 = hmaster0_p & cc36be | !hmaster0_p & !cc36bd;
assign ad4f8d = hmaster2_p & ad4f87 | !hmaster2_p & ad4f8c;
assign ade617 = hmaster1_p & ade616 | !hmaster1_p & ade545;
assign df5151 = hbusreq3 & df5150 | !hbusreq3 & df5142;
assign ad4f28 = hmaster1_p & ad4f27 | !hmaster1_p & ad4f22;
assign v8cc6b4 = hready_p & v8cc507 | !hready_p & v8cc6b3;
assign bd5846 = hbusreq4_p & bd5843 | !hbusreq4_p & bd5845;
assign c3d6c9 = hgrant0_p & c3d6b4 | !hgrant0_p & c3d674;
assign c5c8e9 = hmaster2_p & c5c8e7 | !hmaster2_p & !v845542;
assign v8cc7eb = hlock2 & v8cc435 | !hlock2 & v8cc7ea;
assign v9e9f77 = hbusreq4_p & v9e9f75 | !hbusreq4_p & v9e9f76;
assign b57a35 = hbusreq3_p & b57a11 | !hbusreq3_p & b57a34;
assign d356fe = hbusreq1 & d359aa | !hbusreq1 & v845542;
assign c3cf20 = hbusreq1_p & c3cee8 | !hbusreq1_p & c3cf1f;
assign bd587d = locked_p & bd587c | !locked_p & !v845542;
assign c3d35f = hmaster0_p & c3d35c | !hmaster0_p & c3d35e;
assign c6d407 = start_p & v845542 | !start_p & c6d406;
assign ad4110 = hgrant1_p & ad410f | !hgrant1_p & ad4104;
assign v9f76e6 = hgrant4_p & v9f7c9b | !hgrant4_p & v9f76e5;
assign v9f764f = hbusreq3 & v9f764a | !hbusreq3 & v9f764e;
assign v8cc7c9 = hbusreq1 & v8cc7c5 | !hbusreq1 & v8cc7c8;
assign ad4594 = hmaster0_p & ad4587 | !hmaster0_p & ad4593;
assign v9c81a4 = stateG2_p & v845542 | !stateG2_p & c74b29;
assign ad457d = hready & ad457b | !hready & ad457c;
assign b1c862 = hmaster0_p & b1c85a | !hmaster0_p & b1c861;
assign b57422 = hbusreq4 & b57420 | !hbusreq4 & b57421;
assign d35632 = decide_p & d35631 | !decide_p & v84556c;
assign v9ea4e1 = hgrant2_p & v9ea4df | !hgrant2_p & v9ea4e0;
assign b57951 = hbusreq4_p & b57950 | !hbusreq4_p & v845542;
assign v9f77ec = hgrant0_p & d359c4 | !hgrant0_p & v9f772f;
assign v8cc808 = hbusreq2 & v8cc806 | !hbusreq2 & v8cc807;
assign v9ea3fd = hmaster0_p & v9ea3fa | !hmaster0_p & v9ea3fc;
assign v9f7d29 = hlock1 & v9f7d23 | !hlock1 & !v9f7d28;
assign v9f7e05 = hbusreq1_p & v9f7e04 | !hbusreq1_p & v9f7d19;
assign bd5b9b = hbusreq2_p & bd5b9a | !hbusreq2_p & !v845542;
assign ad484e = hbusreq1 & ad4d98 | !hbusreq1 & ad4845;
assign ad46c6 = hbusreq1_p & ad46c4 | !hbusreq1_p & ad46c5;
assign v9e9f86 = hbusreq3 & v9e9f81 | !hbusreq3 & v9e9f85;
assign bd5786 = hburst0 & bd5781 | !hburst0 & bd5785;
assign dc53dc = hgrant3_p & dc53d9 | !hgrant3_p & !dc53db;
assign v9f77dc = hbusreq4 & v9f77da | !hbusreq4 & v9f77db;
assign df54f2 = hlock1_p & v84556c | !hlock1_p & !v845542;
assign c3d52e = hmaster0_p & c3d52c | !hmaster0_p & c3d52d;
assign v9f78a8 = hmaster1_p & v9f784e | !hmaster1_p & v9f7846;
assign d3501b = hbusreq0 & d3501a | !hbusreq0 & d35aac;
assign v9f7d19 = hbusreq1 & v9f7d17 | !hbusreq1 & v9f7d18;
assign bd5e9c = hbusreq4 & bd5e9b | !hbusreq4 & dc52fc;
assign v9e9faf = hmaster0_p & v9e9f63 | !hmaster0_p & v9e9fae;
assign ad46f3 = hbusreq1 & ad4576 | !hbusreq1 & v845542;
assign v9f7e17 = hbusreq4_p & v9f7e15 | !hbusreq4_p & v9f7e16;
assign ad45e4 = hbusreq4_p & ad45e3 | !hbusreq4_p & v845542;
assign v9f7e0d = hbusreq2 & v9f7e0b | !hbusreq2 & v9f7e0c;
assign b57af2 = hbusreq2 & b57af1 | !hbusreq2 & b57942;
assign ade4c8 = hmastlock_p & adea85 | !hmastlock_p & v845542;
assign v8cc7d9 = hburst0_p & bb9c5a | !hburst0_p & !v8cc7d8;
assign v9f7658 = hlock0_p & v9f7dce | !hlock0_p & v9f7657;
assign v9e9fda = hbusreq2_p & v9ea61b | !hbusreq2_p & v9e9fd9;
assign d354b9 = hbusreq1 & d35be6 | !hbusreq1 & d35beb;
assign v9f7663 = hlock0_p & v9f7ddd | !hlock0_p & v9f7662;
assign c3d6fc = hmaster0_p & c3d6f0 | !hmaster0_p & c3d6fb;
assign b05a53 = hmaster1_p & b05a52 | !hmaster1_p & b05913;
assign b1c793 = hbusreq1 & b1c739 | !hbusreq1 & !v845542;
assign d35412 = hbusreq3 & d35c08 | !hbusreq3 & !v84555a;
assign v9ea4c8 = stateG10_4_p & v9ea4c6 | !stateG10_4_p & v9ea4c7;
assign d359d9 = hbusreq4_p & d359d7 | !hbusreq4_p & d359d8;
assign b05a4f = hmaster0_p & b059a9 | !hmaster0_p & b05968;
assign ad4fdb = hbusreq0_p & ad4fd9 | !hbusreq0_p & !ad4fda;
assign v9f7816 = hbusreq2_p & v9f7813 | !hbusreq2_p & v9f7815;
assign d354ae = hburst0 & d354ac | !hburst0 & d354ad;
assign b1c789 = decide_p & b1c788 | !decide_p & !v845542;
assign b1c5e9 = hlock0_p & b1c5e8 | !hlock0_p & v845542;
assign b1d017 = decide_p & b1cf47 | !decide_p & b1d013;
assign v9f7649 = hbusreq1_p & v9f7e26 | !hbusreq1_p & v9f7648;
assign ad4308 = hbusreq1 & ad4ec6 | !hbusreq1 & v845542;
assign v8cc7df = hlock0 & v8ccb6b | !hlock0 & v8cc7de;
assign c5c8a2 = hmaster1_p & c5c8a1 | !hmaster1_p & c5c89f;
assign ad5031 = stateA1_p & d35905 | !stateA1_p & !v845542;
assign d359ff = stateG10_4_p & v845542 | !stateG10_4_p & d359fe;
assign c3d2b3 = hbusreq3 & c3d2b2 | !hbusreq3 & !v845542;
assign c3d5b9 = stateG10_4_p & c3d5b7 | !stateG10_4_p & !c3d5b8;
assign bd5737 = hburst1_p & v845542 | !hburst1_p & !bb9c5a;
assign c3ce57 = hbusreq1_p & c3ce4a | !hbusreq1_p & c3d305;
assign dc4fe3 = hgrant4_p & adec89 | !hgrant4_p & ade553;
assign v8cc170 = jx2_p & v8cc6b8 | !jx2_p & v8cc16f;
assign bd58c4 = hbusreq4_p & bd58c3 | !hbusreq4_p & dc5010;
assign ade579 = hlock4_p & ade578 | !hlock4_p & !v84556c;
assign b0590a = hlock4 & b058d5 | !hlock4 & b05909;
assign v9ea413 = stateA1_p & v9ea412 | !stateA1_p & v9ea411;
assign d35a5c = hgrant0_p & dc52fa | !hgrant0_p & v84556c;
assign ad440a = hlock3_p & ad4402 | !hlock3_p & ad4409;
assign v9f7d5a = hmaster2_p & v9f7d59 | !hmaster2_p & !v9f7ca6;
assign bd5882 = stateG10_4_p & bd574e | !stateG10_4_p & !bd5881;
assign v9ea440 = hmaster1_p & v9ea43c | !hmaster1_p & v9ea43f;
assign ad46db = hlock0_p & ad46da | !hlock0_p & !v84556e;
assign ad469c = hmaster2_p & ad4699 | !hmaster2_p & ad469b;
assign v9f7774 = hmaster1_p & v9f7773 | !hmaster1_p & v9f776d;
assign v8cc0e7 = hbusreq2 & v8cc0e4 | !hbusreq2 & v8cc0e6;
assign dc5303 = hbusreq3 & dc52fc | !hbusreq3 & dc5302;
assign b05922 = hlock4_p & b058a6 | !hlock4_p & !v9ea3e9;
assign dc53df = jx0_p & dc53d2 | !jx0_p & dc53de;
assign ad504c = hgrant4_p & v84556c | !hgrant4_p & ad504b;
assign ad45bd = hbusreq4_p & ad45bc | !hbusreq4_p & !v845542;
assign ad468c = hmaster0_p & ad468a | !hmaster0_p & ad468b;
assign bd5825 = hbusreq2 & bd5824 | !hbusreq2 & v845542;
assign v9e9e9e = hbusreq4_p & v9e9e9c | !hbusreq4_p & v9e9e9d;
assign v9f768b = locked_p & v9f7d3a | !locked_p & v9ea3e6;
assign v8cc50e = hgrant3_p & v8cc4f7 | !hgrant3_p & v8cc50d;
assign v9ea3ef = hmaster2_p & v9ea3eb | !hmaster2_p & v9ea3ee;
assign ad4351 = hbusreq2_p & ad434e | !hbusreq2_p & ad4350;
assign bd5833 = hbusreq1 & bd5736 | !hbusreq1 & bd5746;
assign v9f7736 = hmaster0_p & v9f7731 | !hmaster0_p & !v9f7735;
assign v9f7d94 = hbusreq4 & v9f7d92 | !hbusreq4 & v9f7d93;
assign d359bd = stateA1_p & v8ccb68 | !stateA1_p & !v845542;
assign ad4437 = hgrant4_p & ad4380 | !hgrant4_p & v845542;
assign v9f7d6f = locked_p & v9f7d3a | !locked_p & !v9f7c9b;
assign b0594f = hgrant0_p & b058a3 | !hgrant0_p & !b0594e;
assign bd586d = hlock4_p & bd586b | !hlock4_p & bd586c;
assign v9f7d88 = hbusreq4_p & v9f7d86 | !hbusreq4_p & v9f7d87;
assign ad4e9d = hmaster2_p & ad4e83 | !hmaster2_p & ad4e9c;
assign v9f7ccc = hbusreq4 & v9f7cca | !hbusreq4 & v9f7ccb;
assign df507d = decide_p & df507c | !decide_p & v845542;
assign d354f9 = hbusreq1_p & d35c08 | !hbusreq1_p & d354f8;
assign c3ce8f = hbusreq1 & v845542 | !hbusreq1 & v845564;
assign ad4deb = hmaster2_p & ad4dde | !hmaster2_p & ad4de2;
assign v9f7878 = hmaster0_p & v9f77fe | !hmaster0_p & v9f77d4;
assign b57acf = hbusreq3 & b578f9 | !hbusreq3 & b57ace;
assign v9e9fb3 = decide_p & v9e9e75 | !decide_p & v9e9fb2;
assign b57ab3 = hlock2 & b57942 | !hlock2 & b57ab2;
assign b1c81b = hbusreq0 & b1c80f | !hbusreq0 & d35a9c;
assign d35583 = hbusreq1_p & d354c4 | !hbusreq1_p & d35582;
assign v9e9e6e = decide_p & v9ea61f | !decide_p & v9e9e6d;
assign b57a6c = hlock1 & b57942 | !hlock1 & b57a6b;
assign bd58fa = hbusreq2 & bd58f9 | !hbusreq2 & v845542;
assign d3577a = hmaster2_p & d3576e | !hmaster2_p & v845542;
assign v9e9fd4 = hgrant2_p & v9ea602 | !hgrant2_p & v9e9fd3;
assign ade583 = hmaster2_p & v845542 | !hmaster2_p & ade582;
assign b1c5dc = hlock2_p & b1c5b5 | !hlock2_p & b1c5db;
assign ade564 = hgrant4_p & v84556c | !hgrant4_p & !ade563;
assign bd587b = hbusreq0 & bd586a | !hbusreq0 & bd587a;
assign d3551d = hlock2_p & d3551b | !hlock2_p & d3551c;
assign d35801 = hmaster1_p & d357f7 | !hmaster1_p & d35800;
assign ad43ac = hmaster0_p & ad43a9 | !hmaster0_p & ad43ab;
assign v9f780d = stateG10_4_p & v9f780b | !stateG10_4_p & !v9f780c;
assign dc52fc = hmaster2_p & v84556c | !hmaster2_p & dc52fb;
assign ad4edd = stateG10_4_p & ad4eda | !stateG10_4_p & ad4edc;
assign v9f7ca8 = hlock0 & v9f7ca7 | !hlock0 & v9f7ca1;
assign c3ce08 = hgrant2_p & v845551 | !hgrant2_p & c3ce07;
assign dc53a5 = hmaster0_p & dc53a4 | !hmaster0_p & v845542;
assign b1c7c3 = hgrant4_p & b1c714 | !hgrant4_p & !b1c7bc;
assign b058e8 = hmaster2_p & b058a3 | !hmaster2_p & b058e7;
assign b1c858 = hbusreq4_p & b1cfb7 | !hbusreq4_p & !b1c857;
assign ad4609 = hbusreq4 & ad4608 | !hbusreq4 & v845542;
assign b1c767 = hmaster2_p & b1c755 | !hmaster2_p & ade4d4;
assign v9f7d99 = hlock1_p & v9f7cb7 | !hlock1_p & v9f7d05;
assign v9f766a = hlock4 & v9f7667 | !hlock4 & v9f7669;
assign ad4745 = hbusreq4_p & ad4744 | !hbusreq4_p & v845542;
assign b1c6dc = hmaster1_p & b1c842 | !hmaster1_p & b1c6db;
assign v9ea3f3 = hmaster1_p & v9ea3f2 | !hmaster1_p & v9ea3f0;
assign bd5812 = hmaster2_p & bd580a | !hmaster2_p & bd5811;
assign b058a5 = stateA1_p & b058a4 | !stateA1_p & !v857440;
assign b5742a = hbusreq2 & b57428 | !hbusreq2 & b57429;
assign v8cc49d = hbusreq0 & v8cc49c | !hbusreq0 & v8cc494;
assign v9ea48b = hmaster1_p & v9ea44a | !hmaster1_p & v9ea48a;
assign bd57fe = hlock0_p & bd57fc | !hlock0_p & bd57fd;
assign c3d524 = hmaster2_p & c3d523 | !hmaster2_p & v845542;
assign ade4ca = hmastlock_p & ade4c9 | !hmastlock_p & v845542;
assign d357f4 = hbusreq4_p & d3578a | !hbusreq4_p & d357f3;
assign cc36f2 = hlock0_p & v84556c | !hlock0_p & !cc36f1;
assign ad4291 = hbusreq1_p & ad4290 | !hbusreq1_p & v845542;
assign v9ea570 = hbusreq4_p & v9ea439 | !hbusreq4_p & v9ea3e6;
assign bd57cc = hbusreq2 & bd57cb | !hbusreq2 & !v845542;
assign dc505c = stateG10_4_p & ade563 | !stateG10_4_p & !dc505b;
assign v9f7cbb = hbusreq4 & v9f7cb9 | !hbusreq4 & v9f7cba;
assign b05a67 = stateG10_4_p & b05a65 | !stateG10_4_p & b05a66;
assign d354a7 = hmaster2_p & d354a4 | !hmaster2_p & d354a6;
assign ad4f56 = hbusreq1_p & ad4f55 | !hbusreq1_p & !v845542;
assign ad44a7 = hmaster2_p & ad44a6 | !hmaster2_p & v845542;
assign bd5841 = hgrant0_p & v845542 | !hgrant0_p & !bd574e;
assign bd5ba3 = hmaster0_p & v845542 | !hmaster0_p & bd5ba2;
assign v9f77da = hbusreq0 & v9f77d7 | !hbusreq0 & v9f77d9;
assign df5158 = hbusreq1 & dc4f6a | !hbusreq1 & v845542;
assign d356a5 = hmaster2_p & v845542 | !hmaster2_p & !d356a4;
assign v9ea571 = hmaster2_p & v9ea570 | !hmaster2_p & v9f20a1;
assign c3d6b4 = locked_p & c3d673 | !locked_p & c3d674;
assign v9f7880 = hgrant0_p & v9f772b | !hgrant0_p & v9f787f;
assign v9ea5d7 = hmaster0_p & v9ea5d6 | !hmaster0_p & v9ea572;
assign v9e9eaf = hgrant2_p & v9e9e9a | !hgrant2_p & v9e9eae;
assign ad503b = hgrant4_p & ad502f | !hgrant4_p & !cc36fc;
assign v8cc0f4 = hmaster0_p & v845542 | !hmaster0_p & v8cc0f2;
assign c3d5e4 = hbusreq4 & c3d5de | !hbusreq4 & !c3d5e3;
assign v9ea5e3 = hmaster0_p & v9ea581 | !hmaster0_p & v9ea5b1;
assign v9f7d78 = hgrant0_p & v9f7cb4 | !hgrant0_p & !v9f7c9f;
assign bd5902 = hready_p & bd5900 | !hready_p & !bd5901;
assign b1c080 = hmaster2_p & b1c07f | !hmaster2_p & b1c858;
assign ad4f63 = hbusreq1_p & ad4f62 | !hbusreq1_p & !v845542;
assign b05951 = stateG10_4_p & b0594f | !stateG10_4_p & b05950;
assign v9e9ea9 = hlock3 & v9e9ea8 | !hlock3 & v9e9ea6;
assign v9ea3e2 = hmaster0_p & v9ea3e1 | !hmaster0_p & v845542;
assign ad43a0 = hbusreq2_p & ad439c | !hbusreq2_p & ad439f;
assign c3d2dd = hbusreq1 & c3d2d6 | !hbusreq1 & c3d2d9;
assign bd5884 = hgrant4_p & v84556c | !hgrant4_p & bd5865;
assign c3d378 = hbusreq3 & c3d376 | !hbusreq3 & v845564;
assign ade5af = hmaster0_p & ade5ad | !hmaster0_p & ade5ae;
assign b1c7ae = hbusreq4 & b1c7a3 | !hbusreq4 & b1c7ad;
assign cc36c7 = hgrant1_p & cc36c6 | !hgrant1_p & d35a49;
assign bd5b7e = hready_p & v845542 | !hready_p & bd5b7d;
assign d357c1 = hlock0_p & v845542 | !hlock0_p & !d3563c;
assign b05a7a = hgrant1_p & b0596a | !hgrant1_p & b05a79;
assign d35769 = hgrant3_p & d35aa3 | !hgrant3_p & !d35768;
assign dc4f71 = hbusreq1 & dc4f6f | !hbusreq1 & dc4f70;
assign bd5934 = hmaster2_p & v84556c | !hmaster2_p & !bd5933;
assign v9f76bc = hbusreq2_p & v9f76b9 | !hbusreq2_p & v9f76bb;
assign ade569 = hgrant1_p & ade54a | !hgrant1_p & !ade568;
assign b1c089 = hgrant1_p & b1c07c | !hgrant1_p & b1c088;
assign ad42ec = hlock1_p & ad42ea | !hlock1_p & ad42eb;
assign v9f7ddc = hbusreq4_p & v9f7dd9 | !hbusreq4_p & !v9f7ddb;
assign bd578a = hburst1 & d35617 | !hburst1 & bd5789;
assign v8cc761 = hmaster1_p & v8cc475 | !hmaster1_p & v8cc760;
assign c3d379 = hmaster2_p & c3d374 | !hmaster2_p & v845542;
assign ade4bf = hburst0 & ade4bd | !hburst0 & ade4be;
assign v9f7dfb = hmaster1_p & v9f7dfa | !hmaster1_p & v9f7d2f;
assign b1c036 = hlock0_p & ade4d9 | !hlock0_p & v845542;
assign b1c77b = hbusreq2 & b1c768 | !hbusreq2 & b1c76a;
assign d35414 = hmaster1_p & d35413 | !hmaster1_p & d35410;
assign ad40fd = hbusreq1 & ad4810 | !hbusreq1 & v845542;
assign v8cc7da = stateG2_p & v845542 | !stateG2_p & v8cc7d9;
assign v9f7dca = hlock4_p & v9f7dc8 | !hlock4_p & !v9f7dc9;
assign bd58b8 = hgrant1_p & bd58b7 | !hgrant1_p & bd58ae;
assign v9ea4e3 = decide_p & v9ea4b2 | !decide_p & v9ea4e2;
assign v8cc7fe = hlock4 & v8cc439 | !hlock4 & v8cc7fd;
assign b05910 = hbusreq3 & b0590e | !hbusreq3 & b0590f;
assign v9ea61c = hmaster0_p & v9ea3e7 | !hmaster0_p & v9ea3f5;
assign d35622 = hmaster0_p & d35621 | !hmaster0_p & dc5318;
assign b1c7fd = hready_p & b1c7fa | !hready_p & !b1c7fc;
assign b0597b = hgrant4_p & b058e7 | !hgrant4_p & v9f7d42;
assign d356b4 = hbusreq3 & d356b1 | !hbusreq3 & d356b3;
assign v9e9fe3 = decide_p & v9e9fda | !decide_p & v9e9fe2;
assign d35aa2 = decide_p & d35aa1 | !decide_p & v84556c;
assign b1c614 = jx1_p & b1c589 | !jx1_p & b1c613;
assign v9f76e8 = hbusreq4_p & v9f7d75 | !hbusreq4_p & v9f76e7;
assign v8cc595 = hbusreq4 & v8cc593 | !hbusreq4 & v8ccbd8;
assign ad46d2 = hbusreq4_p & ad46d1 | !hbusreq4_p & v845542;
assign b1c08c = hgrant2_p & b1c05e | !hgrant2_p & b1c08b;
assign ade5d0 = hmaster2_p & ade4c0 | !hmaster2_p & !ade5cf;
assign v8cc75c = hbusreq3 & v8cc759 | !hbusreq3 & v8cc75b;
assign v9f7672 = hbusreq3 & v9f766f | !hbusreq3 & v9f7671;
assign b1c5b5 = hmaster1_p & v845542 | !hmaster1_p & b1c5b4;
assign ade5c5 = hmaster0_p & ade5bd | !hmaster0_p & ade5c4;
assign b1c706 = decide_p & b1c854 | !decide_p & b1c866;
assign bd581d = hgrant4_p & v84556c | !hgrant4_p & bd580d;
assign bd56d2 = hburst1 & dc5318 | !hburst1 & df54df;
assign b1c7b1 = hbusreq1 & b1c733 | !hbusreq1 & !b1c736;
assign v9f7dd2 = hgrant4_p & v9f7c9f | !hgrant4_p & !v9f7dd0;
assign d356fa = hbusreq2 & d356b1 | !hbusreq2 & d356b3;
assign ad4ed5 = stateG10_4_p & ad4eb3 | !stateG10_4_p & ad4ed4;
assign b05972 = hlock3 & b05971 | !hlock3 & b0596d;
assign d35c00 = hlock4_p & v84557a | !hlock4_p & v845542;
assign d35421 = hbusreq4 & d3541c | !hbusreq4 & d35420;
assign ad4103 = hmaster2_p & ad4102 | !hmaster2_p & v845542;
assign b57ae4 = hbusreq2 & b57ae3 | !hbusreq2 & b579c5;
assign d35a57 = hburst0 & d35a56 | !hburst0 & adea98;
assign b5744e = hgrant3_p & b5744a | !hgrant3_p & b5744d;
assign v9e9ec3 = hlock2 & v9ea4cd | !hlock2 & v9e9ec2;
assign b1c805 = hbusreq1_p & b1c7b8 | !hbusreq1_p & b1c804;
assign b1c7df = hmaster2_p & b1c7de | !hmaster2_p & b1cfb7;
assign d3557b = hmaster2_p & d35579 | !hmaster2_p & d3557a;
assign c3ceb9 = decide_p & c3ceb8 | !decide_p & !c3ce95;
assign ad4776 = hmaster2_p & v845542 | !hmaster2_p & !ad4775;
assign d3543f = hmaster1_p & d3543e | !hmaster1_p & d35438;
assign d35727 = hmaster0_p & d35726 | !hmaster0_p & d356c3;
assign c3d2fa = hbusreq4 & c3d2f4 | !hbusreq4 & !c3d2f9;
assign b05a03 = hmaster0_p & b0593b | !hmaster0_p & b0593a;
assign v9f77a7 = hbusreq1_p & v9f772d | !hbusreq1_p & v9f779f;
assign v9e9f70 = hlock1 & v9e9f68 | !hlock1 & v9e9f6f;
assign df519a = hbusreq1_p & df5199 | !hbusreq1_p & v845542;
assign d35598 = hbusreq4_p & d35434 | !hbusreq4_p & v84554a;
assign ad439b = hmaster0_p & ad4395 | !hmaster0_p & ad439a;
assign ad46b6 = hbusreq1_p & ad46b2 | !hbusreq1_p & !ad46b5;
assign ad5067 = hmaster1_p & ad502d | !hmaster1_p & ad5066;
assign df54f9 = hbusreq1_p & df54f8 | !hbusreq1_p & !v845542;
assign v9f7cfd = hready & v9f7cfc | !hready & v9f7cf8;
assign v9ea45b = hmaster2_p & v9ea444 | !hmaster2_p & v9ea45a;
assign ad4169 = hbusreq2 & ad4fd3 | !hbusreq2 & v845542;
assign b57a2c = hgrant2_p & v845542 | !hgrant2_p & b57a2b;
assign v8cc79b = hbusreq4 & v8cc799 | !hbusreq4 & v8cc79a;
assign b1c07b = hbusreq1 & b1c81b | !hbusreq1 & !b1c81e;
assign ad459a = hbusreq4 & ad4599 | !hbusreq4 & v845542;
assign v84554d = hbusreq1 & v845542 | !hbusreq1 & !v845542;
assign v9f765b = hbusreq4_p & v9f7659 | !hbusreq4_p & v9f765a;
assign b059e7 = hmaster2_p & b059e1 | !hmaster2_p & !b059e6;
assign b058c5 = hbusreq2 & b058c3 | !hbusreq2 & b058c4;
assign b05968 = hbusreq2 & b05966 | !hbusreq2 & b05967;
assign c3ce94 = hmaster0_p & c3d2dd | !hmaster0_p & !c3d2be;
assign v8cc81a = hready_p & v8cc818 | !hready_p & v8cc819;
assign d3549c = hbusreq2 & d35bf7 | !hbusreq2 & d35bf8;
assign v9f7d59 = locked_p & v9f7d58 | !locked_p & !v9ea3e6;
assign c3d69c = hmaster1_p & c3d698 | !hmaster1_p & c3d69b;
assign dc4fba = hmaster2_p & dc4fa6 | !hmaster2_p & !dc4fb9;
assign d35a22 = hbusreq1_p & d359ad | !hbusreq1_p & d35a21;
assign d35523 = hbusreq1_p & d3542e | !hbusreq1_p & d35522;
assign d3568f = hgrant1_p & d35a72 | !hgrant1_p & d3568e;
assign ad4577 = hbusreq1_p & ad4570 | !hbusreq1_p & ad4576;
assign b1c042 = hbusreq0 & b1c041 | !hbusreq0 & b1c847;
assign b1c75b = hmaster2_p & b1c755 | !hmaster2_p & b1c75a;
assign ad4fb6 = hready & v84556c | !hready & ad4f4b;
assign hmaster0 = d6ebcc;
assign ad4fe7 = hgrant4_p & ad4f4a | !hgrant4_p & ad4fe6;
assign d35a02 = hbusreq0_p & d35a01 | !hbusreq0_p & v845542;
assign v8cc5c9 = hgrant3_p & v8ccbdc | !hgrant3_p & v8cc5c8;
assign ad4302 = hgrant2_p & ad4301 | !hgrant2_p & !ad42fa;
assign v8cc4a7 = hlock4 & v8cc494 | !hlock4 & v8cc49d;
assign d35651 = hgrant0_p & dc538c | !hgrant0_p & !v84556c;
assign b05a1b = hgrant4_p & b05941 | !hgrant4_p & b059e3;
assign ad5053 = stateG10_4_p & v84556c | !stateG10_4_p & !ad5052;
assign v9f7d08 = hlock4 & v9f7d05 | !hlock4 & v9f7d07;
assign v9ea598 = hlock2 & v9ea595 | !hlock2 & v9ea597;
assign dc53bd = hlock3_p & dc53bc | !hlock3_p & !v845542;
assign c5c905 = hlock2_p & c5c903 | !hlock2_p & c5c904;
assign d359c3 = hbusreq1 & d359b8 | !hbusreq1 & d359c2;
assign ad4340 = hmaster0_p & ad433c | !hmaster0_p & ad433f;
assign df553a = hbusreq1_p & df5533 | !hbusreq1_p & !v845542;
assign v9e9fcd = hbusreq3_p & v9e9fb5 | !hbusreq3_p & v9e9fcc;
assign b059f3 = hlock2 & b059f0 | !hlock2 & b059f2;
assign b579b5 = hburst1_p & v8b08c1 | !hburst1_p & v84557e;
assign df54fa = hgrant1_p & df54f9 | !hgrant1_p & !v845542;
assign ad3cfe = hgrant1_p & ad3ce9 | !hgrant1_p & ad3cfd;
assign b058d6 = hlock0 & b058d5 | !hlock0 & b058d1;
assign b1c7d2 = hgrant4_p & b1c7b3 | !hgrant4_p & b1c7bc;
assign ad4ffa = hbusreq2_p & ad4ff0 | !hbusreq2_p & ad4ff9;
assign b1c5ba = hburst0 & d3561d | !hburst0 & b1c5b9;
assign bd5909 = hbusreq1_p & bd5908 | !hbusreq1_p & v845564;
assign v9f77f8 = hlock2_p & v9f77f6 | !hlock2_p & v9f77f7;
assign bd58e8 = hbusreq2 & bd58e7 | !hbusreq2 & v845542;
assign c3d67c = hmaster0_p & c3d677 | !hmaster0_p & c3d67b;
assign bd56db = hmaster0_p & v845542 | !hmaster0_p & bd56da;
assign ad4fab = hburst0_p & c73a9a | !hburst0_p & !e199ba;
assign c3d527 = hbusreq1_p & c3d479 | !hbusreq1_p & c3d526;
assign ad4349 = decide_p & ad42cf | !decide_p & ad4348;
assign ac1460 = hgrant1_p & ac145f | !hgrant1_p & ac145c;
assign b579b0 = hmaster1_p & b579af | !hmaster1_p & v845542;
assign dc52f8 = hmastlock_p & adea97 | !hmastlock_p & !v845542;
assign d35a05 = hgrant4_p & d359e8 | !hgrant4_p & d35a03;
assign v9f7d41 = stateA1_p & v845542 | !stateA1_p & v845582;
assign b05993 = hlock0 & b05992 | !hlock0 & b05986;
assign ad4e23 = hmaster0_p & ad4e22 | !hmaster0_p & v845542;
assign b05949 = hready_p & b0591b | !hready_p & !b05948;
assign dc53aa = hready_p & dc5393 | !hready_p & !dc53a9;
assign v9f771d = hmaster1_p & v9f771c | !hmaster1_p & v9f7d64;
assign v845551 = hbusreq2 & v845542 | !hbusreq2 & !v845542;
assign b05940 = hbusreq0_p & v9ea463 | !hbusreq0_p & v9f769c;
assign v9f7805 = hlock3 & v9f7804 | !hlock3 & v9f7803;
assign bd5805 = hgrant0_p & v845542 | !hgrant0_p & !bd57fb;
assign bd5b87 = hburst0 & d35a56 | !hburst0 & bd5b86;
assign adeab5 = decide_p & adeab4 | !decide_p & adeaa7;
assign ba7c75 = hgrant3_p & ba7c6a | !hgrant3_p & ba7c74;
assign c3ce46 = hbusreq1 & c3d301 | !hbusreq1 & c3d305;
assign dc4f68 = hmaster2_p & ade4bf | !hmaster2_p & ade4c5;
assign ade5aa = hbusreq4_p & adeca0 | !hbusreq4_p & !v845542;
assign d35be6 = hmaster2_p & d35be3 | !hmaster2_p & d35be5;
assign ad468a = hbusreq2 & ad4577 | !hbusreq2 & v845542;
assign ad505d = hbusreq0_p & v845542 | !hbusreq0_p & !ad5032;
assign b57537 = jx0_p & b57450 | !jx0_p & b57536;
assign ad4e9f = hbusreq4_p & ad4e9e | !hbusreq4_p & adeaa4;
assign d354cb = hlock4_p & d35a0e | !hlock4_p & !d35a5f;
assign d359f0 = hgrant4_p & d359ef | !hgrant4_p & v845542;
assign bd5e1e = hbusreq4 & bd5e1d | !hbusreq4 & dc531a;
assign b1cbf4 = hbusreq4_p & b1cbf3 | !hbusreq4_p & b1cfcc;
assign ad474b = hbusreq4 & ad474a | !hbusreq4 & v845542;
assign c3cec3 = hgrant4_p & v845542 | !hgrant4_p & !c3cec2;
assign c3cea5 = hgrant1_p & c3d2dd | !hgrant1_p & c3cea4;
assign v9f7d71 = hgrant0_p & v9f7c9b | !hgrant0_p & !v9f7d6f;
assign b05a0b = stateG10_4_p & v9ea464 | !stateG10_4_p & b05a0a;
assign b1c7b8 = hbusreq0 & b1c7b7 | !hbusreq0 & !v845542;
assign ade5b6 = hmaster1_p & ade5b5 | !hmaster1_p & ade5a4;
assign ad414b = hbusreq2 & ad414a | !hbusreq2 & v845542;
assign df514a = hbusreq1 & dc4fd9 | !hbusreq1 & v845542;
assign c3cdfc = hgrant2_p & v845551 | !hgrant2_p & c3cdfb;
assign v9f76a8 = hgrant2_p & v9f768a | !hgrant2_p & v9f76a7;
assign c3d349 = hbusreq3 & c3d348 | !hbusreq3 & c3d306;
assign v8ccb84 = hmaster1_p & v8ccb83 | !hmaster1_p & v8ccb81;
assign ad42bb = hlock1_p & ad42af | !hlock1_p & ad42ba;
assign v9ea5f5 = hbusreq2_p & v9ea3f1 | !hbusreq2_p & v9ea5f4;
assign adec9f = hmaster0_p & adec9d | !hmaster0_p & adec9e;
assign v9f7cdc = hlock0_p & v9f7cb6 | !hlock0_p & v9f7cdb;
assign ad4278 = hbusreq1_p & ad4277 | !hbusreq1_p & v845542;
assign v9ea405 = hmaster0_p & v9ea400 | !hmaster0_p & v9ea404;
assign ad4136 = hlock4_p & ad4135 | !hlock4_p & !v845576;
assign c3cf1d = hbusreq2 & c3cf1b | !hbusreq2 & c3cee4;
assign ad4f05 = hmaster2_p & ad4eff | !hmaster2_p & ad4f04;
assign c3d357 = hgrant2_p & v845551 | !hgrant2_p & c3d356;
assign v9e9ef4 = hmaster1_p & v9e9ef3 | !hmaster1_p & v9e9ef1;
assign ad4f5b = hbusreq1 & ad4f3b | !hbusreq1 & ad4f40;
assign dc503a = hgrant4_p & ade56d | !hgrant4_p & !adeca1;
assign v8cc16f = jx0_p & v8cc038 | !jx0_p & v8cc16c;
assign b573f9 = hready_p & b5799c | !hready_p & b573f8;
assign ad3cbe = hmaster0_p & ad43ab | !hmaster0_p & ad448f;
assign b1cbf0 = hlock4_p & b1cfc2 | !hlock4_p & b1cff6;
assign v9f770c = hgrant2_p & v9f76dd | !hgrant2_p & v9f770b;
assign dc4fae = hmaster2_p & dc4fac | !hmaster2_p & !dc4fa9;
assign ad4746 = hmaster2_p & v845542 | !hmaster2_p & ad4745;
assign bd583b = hbusreq1_p & bd5835 | !hbusreq1_p & bd583a;
assign c3d33d = stateG10_4_p & c3d33b | !stateG10_4_p & !c3d33c;
assign b574cc = hbusreq3 & b574ca | !hbusreq3 & b574cb;
assign b1c85d = stateG10_4_p & b1c85b | !stateG10_4_p & !b1c85c;
assign d357e9 = hbusreq0 & v84554a | !hbusreq0 & !v845542;
assign d357ab = hbusreq2_p & d357aa | !hbusreq2_p & d357a9;
assign d355a5 = hburst0_p & v845542 | !hburst0_p & !d355a4;
assign b05a78 = hbusreq2 & b05a76 | !hbusreq2 & b05a77;
assign v9f78ae = hbusreq3_p & v9f7855 | !hbusreq3_p & v9f78ad;
assign b5741f = hlock0 & b57987 | !hlock0 & b5741e;
assign ad4eb5 = hgrant4_p & ad4e53 | !hgrant4_p & ad4eb3;
assign b1c7bc = hlock0_p & b1c7bb | !hlock0_p & !b1c70e;
assign v9f7e39 = hbusreq1 & v9f7e37 | !hbusreq1 & v9f7e38;
assign v9f7747 = hbusreq0 & v9f7744 | !hbusreq0 & v9f7746;
assign bd5860 = hbusreq4_p & bd585d | !hbusreq4_p & bd585f;
assign c3d6f8 = stateG10_4_p & c3d6f6 | !stateG10_4_p & !c3d6f7;
assign b579e3 = hbusreq1 & b579e1 | !hbusreq1 & b579e2;
assign ade59b = hbusreq0_p & ade599 | !hbusreq0_p & ade59a;
assign b0591e = hmaster2_p & b0591c | !hmaster2_p & !v9ea3e9;
assign ade59e = hlock0_p & ade595 | !hlock0_p & !ade562;
assign ade5cc = hmastlock_p & ade5cb | !hmastlock_p & v845542;
assign c3d701 = hgrant1_p & c3d676 | !hgrant1_p & c3d6ee;
assign c3d333 = hgrant2_p & v845551 | !hgrant2_p & c3d332;
assign ad42da = hmaster1_p & ad42d4 | !hmaster1_p & ad42d9;
assign b05925 = hmaster2_p & b05923 | !hmaster2_p & b05924;
assign v9f7706 = hlock3 & v9f7705 | !hlock3 & v9f7703;
assign v8cc487 = hbusreq1_p & v8ccbd8 | !hbusreq1_p & v8cc484;
assign ad42ce = hbusreq2_p & ad42cd | !hbusreq2_p & ad42cc;
assign v8cc0dc = hlock4 & v8cc494 | !hlock4 & v8cc0db;
assign v9ea57d = hbusreq2_p & v9ea57a | !hbusreq2_p & v9ea57c;
assign ad477c = hbusreq4 & ad4777 | !hbusreq4 & ad477b;
assign b1cf34 = hmaster0_p & v845542 | !hmaster0_p & b1cf33;
assign b058be = hlock1 & b058b8 | !hlock1 & b058bd;
assign df553c = hmaster0_p & df553b | !hmaster0_p & df5539;
assign b573e5 = hlock2 & b57942 | !hlock2 & b573e4;
assign c3d6f5 = hbusreq0_p & c3d6c7 | !hbusreq0_p & !c3d674;
assign b1cfd4 = hmaster1_p & b1cfb8 | !hmaster1_p & b1cfd3;
assign bd5867 = hgrant4_p & c3d689 | !hgrant4_p & bd5865;
assign ad42be = hmaster1_p & ad42a8 | !hmaster1_p & ad42bd;
assign b05a16 = hgrant1_p & b05a10 | !hgrant1_p & b05a15;
assign ad4557 = hbusreq4 & ad4556 | !hbusreq4 & v845542;
assign v8cc789 = hmaster0_p & v8cc788 | !hmaster0_p & v845542;
assign c3d2ed = hbusreq4_p & c3d2eb | !hbusreq4_p & c3d2ec;
assign b059d2 = hlock2 & b059cf | !hlock2 & b059d1;
assign v8cc169 = hgrant3_p & v8ccbdc | !hgrant3_p & v8cc167;
assign bd57f0 = hready_p & bd5780 | !hready_p & bd57ef;
assign d35998 = hgrant4_p & d3597f | !hgrant4_p & d35997;
assign bd579f = hmaster2_p & bd5786 | !hmaster2_p & !ade4d9;
assign dc53d7 = hlock3_p & dc53a2 | !hlock3_p & v845542;
assign b8f6e4 = hmaster1_p & b8f6e1 | !hmaster1_p & b8f6e3;
assign d357fc = hmaster2_p & d357a2 | !hmaster2_p & d35a9c;
assign bd58bd = hlock0_p & bd58bc | !hlock0_p & !ade562;
assign v9f7691 = hgrant1_p & v9f7d5b | !hgrant1_p & v9f7690;
assign v9f7e36 = hbusreq4 & v9f7e34 | !hbusreq4 & v9f7e35;
assign v9e9fa7 = hmaster0_p & v9e9ee9 | !hmaster0_p & v9e9fa6;
assign v9e9eeb = locked_p & v845542 | !locked_p & v9ea438;
assign v8cc4f6 = decide_p & v8cc4f4 | !decide_p & v8ccbda;
assign d35778 = hbusreq0 & d3576e | !hbusreq0 & v845542;
assign dc5062 = hmaster2_p & dc505d | !hmaster2_p & dc5061;
assign c3ce6c = hbusreq1 & c3d375 | !hbusreq1 & v845542;
assign b5740f = hlock1 & b578f1 | !hlock1 & b5740e;
assign v9f7d50 = hmaster1_p & v9f7d4f | !hmaster1_p & v9f7d47;
assign v8cc7e9 = hlock3 & v8cc435 | !hlock3 & v8cc7e8;
assign v9f786a = hbusreq2 & v9f7868 | !hbusreq2 & v9f7869;
assign b0595d = hbusreq0 & b0595a | !hbusreq0 & b0595c;
assign ad4e7d = hmaster2_p & ad4e7c | !hmaster2_p & v845542;
assign d354ec = hready_p & d354eb | !hready_p & d35444;
assign d357e0 = hgrant2_p & d357be | !hgrant2_p & d357df;
assign c3cef5 = hmaster2_p & c3cef4 | !hmaster2_p & v845576;
assign df50d1 = hgrant2_p & v845542 | !hgrant2_p & !df50d0;
assign v9f7836 = hbusreq1_p & v9f7824 | !hbusreq1_p & v9f7835;
assign v84556e = hgrant0_p & v845542 | !hgrant0_p & !v845542;
assign c3ce35 = hbusreq1_p & c3ce34 | !hbusreq1_p & v845542;
assign d35a67 = hlock4_p & d35a65 | !hlock4_p & !d35a66;
assign d35736 = hbusreq1_p & d356e1 | !hbusreq1_p & d35a99;
assign b1c56d = hbusreq2_p & b1cc04 | !hbusreq2_p & b1c56c;
assign ad5023 = hready & v845542 | !hready & !c3d327;
assign d35a92 = hready_p & d35a7b | !hready_p & d3597d;
assign ad3d22 = hmaster0_p & ad448f | !hmaster0_p & ad43ab;
assign b5740a = hlock0 & b578f1 | !hlock0 & b57409;
assign c5c89f = hmaster0_p & c5c89a | !hmaster0_p & c5c89e;
assign ad4f3e = hburst0 & v845542 | !hburst0 & adec8d;
assign b0591f = hlock1_p & b0591d | !hlock1_p & b0591e;
assign d3541f = hbusreq4_p & d3541e | !hbusreq4_p & v845542;
assign c3d47b = hbusreq4 & v845564 | !hbusreq4 & !v845542;
assign v9ea3e7 = hmaster2_p & v9f20a1 | !hmaster2_p & v9ea3e6;
assign df51a2 = hready_p & df51a0 | !hready_p & df51a1;
assign b1c03e = hbusreq1 & b1c034 | !hbusreq1 & b1c039;
assign c3d742 = stateG10_4_p & c3d740 | !stateG10_4_p & !c3d741;
assign d35024 = hgrant3_p & d35804 | !hgrant3_p & d35023;
assign bd5835 = hlock1_p & bd5833 | !hlock1_p & bd5834;
assign v8cc82c = hgrant2_p & v845542 | !hgrant2_p & v8cc82a;
assign bd58f1 = hmaster1_p & bd58f0 | !hmaster1_p & bd57b1;
assign dc4f91 = hbusreq4 & dc4f8e | !hbusreq4 & dc4f90;
assign d356aa = hlock1_p & d35991 | !hlock1_p & v84556c;
assign v9f7716 = decide_p & v9f770d | !decide_p & v9f7715;
assign c3d6b2 = hgrant1_p & c3d6a4 | !hgrant1_p & c3d6b1;
assign df517a = hbusreq1 & dc5014 | !hbusreq1 & v845542;
assign d3573d = hbusreq2 & d356bb | !hbusreq2 & d356ad;
assign c3d3ac = hgrant3_p & c3d394 | !hgrant3_p & c3d3ab;
assign ade55b = hgrant4_p & v84556c | !hgrant4_p & !adec89;
assign ac145a = stateG10_4_p & ac1458 | !stateG10_4_p & ac1459;
assign d35703 = hbusreq1 & d35a73 | !hbusreq1 & v845542;
assign bd573f = hburst1 & d35a4d | !hburst1 & bd573d;
assign c3d5b6 = hmaster2_p & c3d5b5 | !hmaster2_p & v845542;
assign d356d0 = hlock3_p & d356bf | !hlock3_p & !d356cf;
assign ade61a = hgrant2_p & ade617 | !hgrant2_p & ade619;
assign b579d1 = hlock0_p & b579cc | !hlock0_p & b579d0;
assign c5c931 = hbusreq1_p & c5c88f | !hbusreq1_p & c5c930;
assign ade57a = hbusreq4_p & ade579 | !hbusreq4_p & !v845542;
assign c3ce38 = hbusreq3 & c3ce35 | !hbusreq3 & c3ce37;
assign d3576e = hlock0_p & v845542 | !hlock0_p & v84556c;
assign ad460f = hmaster1_p & ad460c | !hmaster1_p & ad460e;
assign ad4ee6 = stateG10_4_p & ad4ee3 | !stateG10_4_p & ad4ee5;
assign d356c2 = hbusreq3 & d356c0 | !hbusreq3 & !d356c1;
assign ad504a = hbusreq0_p & ad5049 | !hbusreq0_p & !ad503f;
assign v9f7cc8 = hmaster2_p & v9f7ca5 | !hmaster2_p & v9f7cc7;
assign df5177 = hbusreq2 & df514b | !hbusreq2 & df5142;
assign b05963 = hgrant1_p & b0594d | !hgrant1_p & b05962;
assign ad41b4 = hbusreq2 & ad5034 | !hbusreq2 & c3d2d9;
assign v9e9eb4 = hlock2 & v9ea4cd | !hlock2 & v9e9eb3;
assign v9f7cea = hmaster1_p & v9f7cc3 | !hmaster1_p & v9f7ce9;
assign v9e9f61 = hbusreq3 & v9e9f5e | !hbusreq3 & v9e9f60;
assign dc4f9b = hmastlock_p & ade4c1 | !hmastlock_p & !v845542;
assign ad4fb8 = hmaster0_p & ad4fb5 | !hmaster0_p & ad4fb7;
assign c3ce67 = hbusreq3 & c3ce61 | !hbusreq3 & c3ce66;
assign ac147c = hmaster0_p & ac1474 | !hmaster0_p & ac147b;
assign c3ce81 = hbusreq1_p & c3ce46 | !hbusreq1_p & c3d3a3;
assign v8cc757 = hbusreq1 & v8cc4a9 | !hbusreq1 & v8cc494;
assign v9f77c7 = hbusreq4_p & v9f77c5 | !hbusreq4_p & v9f77c6;
assign bd5942 = jx2_p & bd5906 | !jx2_p & bd5941;
assign bd593d = decide_p & bd592b | !decide_p & !v845572;
assign d356b5 = hlock1_p & d359e5 | !hlock1_p & v84556c;
assign v9f7cf0 = hmaster1_p & v9f7cef | !hmaster1_p & v9f7ce9;
assign c3d6d7 = hgrant2_p & c3d6d6 | !hgrant2_p & !c3d6d3;
assign b1c561 = hbusreq0 & b1c55e | !hbusreq0 & b1c560;
assign ad4ebb = stateG10_4_p & v845542 | !stateG10_4_p & ad4eba;
assign v9f7887 = hlock0 & v9f77d8 | !hlock0 & v9f7886;
assign b57a75 = hmaster2_p & b579cb | !hmaster2_p & b57a74;
assign ad46e4 = hmaster0_p & ad46c3 | !hmaster0_p & ad46e3;
assign ad4699 = hbusreq4_p & ad4698 | !hbusreq4_p & v845542;
assign b1c06b = hbusreq0 & b1c06a | !hbusreq0 & b1c85e;
assign b573df = hmaster1_p & b579b4 | !hmaster1_p & b573de;
assign c5c952 = hbusreq2_p & c5c93e | !hbusreq2_p & c5c951;
assign df5170 = hbusreq1 & dc4fce | !hbusreq1 & v845542;
assign d356e8 = hmaster1_p & d356e7 | !hmaster1_p & d356e5;
assign v9f7caf = hlock3 & v9f7ca7 | !hlock3 & v9f7cae;
assign d358f3 = hbusreq1_p & d358f2 | !hbusreq1_p & v845542;
assign ad4ddf = hready & ad4ddd | !hready & !ad4dde;
assign v9f77c0 = stateG10_4_p & v9f77be | !stateG10_4_p & v9f77bf;
assign ad42d2 = hbusreq1 & ad501b | !hbusreq1 & v845547;
assign c3d731 = hready_p & c3d726 | !hready_p & c3d730;
assign b059e6 = hbusreq4_p & b059e4 | !hbusreq4_p & !b059e5;
assign c3d759 = hmaster1_p & c3d758 | !hmaster1_p & c3d70f;
assign c3d5a6 = hbusreq2 & c3d5a3 | !hbusreq2 & c3d368;
assign c3d503 = hbusreq4 & c3d502 | !hbusreq4 & !c3d304;
assign b1c040 = hbusreq4_p & b1c756 | !hbusreq4_p & !b1c031;
assign d35a63 = hgrant0_p & dc5300 | !hgrant0_p & !v84556c;
assign ad42d9 = hmaster0_p & ad42d6 | !hmaster0_p & ad42d8;
assign b1c039 = hbusreq0 & b1c038 | !hbusreq0 & !b1c841;
assign d3599e = hgrant4_p & d3597f | !hgrant4_p & v845542;
assign ad4414 = hbusreq1_p & ad4411 | !hbusreq1_p & ad4413;
assign d35014 = hbusreq1_p & d357cd | !hbusreq1_p & d35013;
assign c5c9ab = hready_p & c5c9a0 | !hready_p & !c5c9aa;
assign c3d37e = hbusreq1 & c3d375 | !hbusreq1 & c3d379;
assign ad4ece = hmaster2_p & ad4ecb | !hmaster2_p & ad4ecd;
assign d35517 = hbusreq4_p & d35516 | !hbusreq4_p & v845542;
assign b1cfff = hlock0_p & b1cffe | !hlock0_p & v845542;
assign v9ea3f1 = hmaster1_p & v9f20a1 | !hmaster1_p & v9ea3f0;
assign c3d359 = hlock3_p & c3d333 | !hlock3_p & c3d357;
assign df54de = stateA1_p & e0edf9 | !stateA1_p & ade4b7;
assign b57986 = hgrant4_p & v845542 | !hgrant4_p & b57952;
assign c5c8f2 = hgrant0_p & v845542 | !hgrant0_p & !c5c8f1;
assign dc5077 = hmaster1_p & dc506f | !hmaster1_p & dc5076;
assign d35984 = hmaster2_p & d3597f | !hmaster2_p & d35983;
assign b574ba = hbusreq1_p & b57942 | !hbusreq1_p & b574b9;
assign v9e9e7a = hmaster0_p & v9ea3fa | !hmaster0_p & v9e9e79;
assign ad47f8 = hmaster0_p & ad456f | !hmaster0_p & ad459d;
assign b059de = hmaster2_p & b059d7 | !hmaster2_p & !b059dd;
assign v9f77ac = hbusreq4_p & v845542 | !hbusreq4_p & v9f779d;
assign b1c5b3 = hbusreq2 & b1c58b | !hbusreq2 & b1cf2c;
assign ad42f7 = hbusreq1_p & ad42f6 | !hbusreq1_p & v845542;
assign v9f76b0 = decide_p & v9f7d56 | !decide_p & !v9f76af;
assign v9ea424 = hgrant1_p & v845542 | !hgrant1_p & v9ea423;
assign v8cc12f = hready_p & v8cc507 | !hready_p & v8cc12d;
assign ad4fa9 = hbusreq2_p & ad4fa2 | !hbusreq2_p & !ad4fa8;
assign c3ceef = hgrant4_p & v845542 | !hgrant4_p & c3ceee;
assign ad4154 = hmaster2_p & ad4151 | !hmaster2_p & ad4153;
assign v9ea492 = hready & v9ea491 | !hready & v9ea43b;
assign df5137 = hmaster2_p & adec89 | !hmaster2_p & dc5037;
assign v9ea5b2 = hmaster0_p & v9ea3fc | !hmaster0_p & v9ea5b1;
assign v9f7d1d = hbusreq3 & v9f7d1a | !hbusreq3 & v9f7d1c;
assign ad4dd1 = hmaster2_p & ad4db2 | !hmaster2_p & ad4dce;
assign ad4ef7 = hlock0_p & dc52fa | !hlock0_p & !v845542;
assign b059ee = hbusreq1 & b059ec | !hbusreq1 & b059ed;
assign d356e1 = hlock1_p & v845542 | !hlock1_p & d356e0;
assign ad481a = hlock2_p & ad4813 | !hlock2_p & ad4819;
assign v9ea491 = hbusreq4 & v9ea48f | !hbusreq4 & v9ea490;
assign d35515 = hbusreq1_p & d35514 | !hbusreq1_p & d3542e;
assign ad4140 = hbusreq4_p & ad413f | !hbusreq4_p & adeaa4;
assign v9f7742 = stateA1_p & v9f7741 | !stateA1_p & v84557c;
assign v9ea624 = hmaster0_p & v9ea623 | !hmaster0_p & v9ea3fc;
assign v9ea57e = decide_p & v9ea56f | !decide_p & v9ea57d;
assign ad433b = hbusreq1_p & ad433a | !hbusreq1_p & ad5023;
assign dc5042 = hgrant4_p & dc5037 | !hgrant4_p & ade563;
assign ad427e = hmaster0_p & ad4270 | !hmaster0_p & ad427d;
assign bd582c = hmaster2_p & bd5817 | !hmaster2_p & v845542;
assign c3d74c = hbusreq2_p & c3d73a | !hbusreq2_p & !c3d74b;
assign adec97 = hmastlock_p & adec96 | !hmastlock_p & v845542;
assign ad4f70 = stateG10_4_p & ad4f36 | !stateG10_4_p & !ad4f6f;
assign b059dd = hbusreq4_p & b059db | !hbusreq4_p & !b059dc;
assign c3d725 = hbusreq2_p & c3d722 | !hbusreq2_p & c3d724;
assign v9f767e = hgrant1_p & v9f7ccf | !hgrant1_p & v9f7648;
assign v8cc599 = hlock1 & v8ccbd8 | !hlock1 & v8cc598;
assign b5743a = hmaster0_p & b57438 | !hmaster0_p & b57439;
assign ac1477 = hgrant4_p & v845542 | !hgrant4_p & !ac1465;
assign ad435d = hmaster0_p & ad435c | !hmaster0_p & ad42e4;
assign b1c581 = hbusreq4 & b1c57d | !hbusreq4 & b1c580;
assign v9f7686 = hgrant2_p & v9f767d | !hgrant2_p & v9f7685;
assign v9f7d39 = decide_p & v9f7d38 | !decide_p & v9f7cf1;
assign dc5070 = hmaster2_p & c3d66d | !hmaster2_p & !adeca0;
assign b05a6e = hready & b05a6d | !hready & b05a69;
assign v8cc496 = hgrant0_p & v8cc47a | !hgrant0_p & v845542;
assign v9ea482 = hready & v9ea481 | !hready & v9ea46d;
assign ad43de = hbusreq1 & ad43db | !hbusreq1 & ad43dd;
assign b1c7ca = hbusreq1_p & b1c7ae | !hbusreq1_p & b1c7c9;
assign v9f7d30 = hmaster1_p & v9f7d11 | !hmaster1_p & v9f7d2f;
assign c3cf12 = hmaster0_p & c3d368 | !hmaster0_p & c3ce15;
assign ad4fc6 = hburst0_p & c73a9a | !hburst0_p & !c76647;
assign cc3705 = hmaster1_p & cc36f7 | !hmaster1_p & cc3704;
assign ad42fc = hbusreq2 & ad4281 | !hbusreq2 & !v845542;
assign ad48b6 = hlock1_p & ad48b5 | !hlock1_p & v845542;
assign v8cc5b5 = hbusreq2 & v8cc5b3 | !hbusreq2 & v8cc5b4;
assign df54ef = decide_p & df54ee | !decide_p & v845542;
assign c3d578 = hbusreq4_p & c3d4db | !hbusreq4_p & c3d39b;
assign ad4701 = hmaster2_p & ad46fe | !hmaster2_p & ad4700;
assign b573fc = hlock2 & b57942 | !hlock2 & b573fb;
assign v8cc61a = hbusreq3 & v8cc488 | !hbusreq3 & v8cc619;
assign c3d6a6 = hlock0_p & c3d6a5 | !hlock0_p & !c3d669;
assign d354b2 = hlock0_p & d354b0 | !hlock0_p & !d354b1;
assign d35797 = hbusreq1 & d3578d | !hbusreq1 & d35790;
assign c5c899 = hlock1_p & c5c897 | !hlock1_p & c5c898;
assign v8cc7e2 = hlock4 & v8ccb6b | !hlock4 & v8cc7e1;
assign c3d2cb = hready & c3d2ca | !hready & v845564;
assign b1c61b = decide_p & b1c61a | !decide_p & v845542;
assign v9ea585 = hbusreq4_p & v9f20a1 | !hbusreq4_p & v9ea4b3;
assign v8cc12a = decide_p & v8cc4f4 | !decide_p & v8cc129;
assign d35aa8 = hgrant2_p & v845542 | !hgrant2_p & d35aa7;
assign v9ea47a = hmaster2_p & v9ea479 | !hmaster2_p & v9ea46c;
assign d35791 = hbusreq3 & d3578d | !hbusreq3 & d35790;
assign v85746a = hbusreq3_p & v92e9d9 | !hbusreq3_p & !v845542;
assign dc501b = hbusreq1 & dc5019 | !hbusreq1 & !dc501a;
assign ad431b = hgrant1_p & v845542 | !hgrant1_p & ad431a;
assign b57947 = hmaster0_p & v845542 | !hmaster0_p & b578f1;
assign ad45a1 = hbusreq4_p & ad4f4a | !hbusreq4_p & v845542;
assign c3d754 = hbusreq2_p & c3d74f | !hbusreq2_p & c3d753;
assign v8cc7f1 = hbusreq4_p & v8cc7b9 | !hbusreq4_p & v8cc7f0;
assign dc4f6d = hmaster0_p & dc4f67 | !hmaster0_p & dc4f6c;
assign ba7c7e = hgrant3_p & ba7c6a | !hgrant3_p & ba7c7d;
assign d3591e = hmaster1_p & d35913 | !hmaster1_p & d3591d;
assign v8cc4a0 = hbusreq4_p & v8cc48e | !hbusreq4_p & v8cc49f;
assign b059a3 = hmaster0_p & b05901 | !hmaster0_p & b058f6;
assign bd575e = hmaster2_p & v84556c | !hmaster2_p & bd575d;
assign b05933 = hmaster1_p & b05932 | !hmaster1_p & b05926;
assign bd5b69 = stateA1_p & d35905 | !stateA1_p & adea85;
assign v9ea5b9 = decide_p & v9ea56f | !decide_p & v9ea5b8;
assign c3d72c = hmaster1_p & c3d72b | !hmaster1_p & c3d69b;
assign b57a29 = hgrant1_p & b5794d | !hgrant1_p & b57a27;
assign v845547 = hready & v845542 | !hready & !v845542;
assign ade4ac = hmaster2_p & v845542 | !hmaster2_p & ade4ab;
assign dc4f82 = hbusreq3 & dc4f81 | !hbusreq3 & v845542;
assign dc5391 = hbusreq2_p & dc5390 | !hbusreq2_p & dc4f63;
assign bd57e9 = hbusreq2 & bd57d0 | !hbusreq2 & !v845542;
assign ad4db3 = hmaster2_p & ad4db2 | !hmaster2_p & !ad4dad;
assign v9f7dff = hbusreq3 & v9f7daa | !hbusreq3 & v9f7dfe;
assign c3d2f4 = hbusreq0 & c3d2ee | !hbusreq0 & c3d2f3;
assign v9e9e72 = jx1_p & v9ea5eb | !jx1_p & v9e9e71;
assign c3d5d7 = hbusreq4_p & c3d5d5 | !hbusreq4_p & c3d5d6;
assign ad42e6 = hbusreq2 & ad4275 | !hbusreq2 & v845542;
assign ad4313 = hbusreq1 & ad4fc2 | !hbusreq1 & v845542;
assign ade547 = hbusreq1 & adec8a | !hbusreq1 & adec93;
assign ad3d16 = hmaster0_p & ad4411 | !hmaster0_p & ad3d15;
assign bd5e1c = hbusreq4_p & bd5e1b | !hbusreq4_p & !v845542;
assign v8cc4da = hgrant2_p & v8cc4bb | !hgrant2_p & v8cc4b2;
assign hmaster2 = !v8da604;
assign b1c7be = hgrant4_p & b1c73c | !hgrant4_p & b1c7bc;
assign v9f76ff = hbusreq3 & v9f76fb | !hbusreq3 & v9f76fe;
assign v9ea4d7 = stateG10_4_p & v9ea4d5 | !stateG10_4_p & v9ea4d6;
assign b1c7e2 = hgrant1_p & b1c7ce | !hgrant1_p & b1c7e1;
assign ad42e7 = hbusreq2 & ad4278 | !hbusreq2 & v845542;
assign c3d685 = hmaster2_p & c3d669 | !hmaster2_p & !c3d674;
assign b05a92 = hgrant2_p & b05a8f | !hgrant2_p & b05a91;
assign v8d29fa = hmastlock_p & v8d29f9 | !hmastlock_p & v845542;
assign v9f77e1 = hbusreq1_p & v9f77c8 | !hbusreq1_p & v9f77d8;
assign c5c975 = hbusreq1_p & c5c8e8 | !hbusreq1_p & c5c974;
assign v9ea460 = hlock2 & v9ea45e | !hlock2 & v9ea45f;
assign ad42c1 = hlock1_p & ad42c0 | !hlock1_p & !v84554d;
assign ad42b1 = hmaster2_p & ad42b0 | !hmaster2_p & ad45e2;
assign v9f7699 = hbusreq1_p & v9f7690 | !hbusreq1_p & v9f7698;
assign ad4e91 = hready & ad4e81 | !hready & ad4e90;
assign b1c050 = hmaster0_p & b1c7f5 | !hmaster0_p & b1c7af;
assign d354e7 = hmaster0_p & d354b8 | !hmaster0_p & d354e6;
assign d3578d = hbusreq0 & d3578c | !hbusreq0 & v845542;
assign c3d38c = hbusreq3 & c3d38b | !hbusreq3 & !v845542;
assign b1cc02 = hmaster0_p & b1cfb8 | !hmaster0_p & b1cc01;
assign v9e9ea2 = hbusreq1_p & v9e9e9f | !hbusreq1_p & v9ea4ca;
assign d35798 = hmaster2_p & d3578a | !hmaster2_p & v84554a;
assign ad4fbd = hbusreq4_p & ad4fbb | !hbusreq4_p & ad4fbc;
assign ade596 = hburst1 & v845542 | !hburst1 & !v889629;
assign v9f76c6 = hmaster2_p & v9f76c5 | !hmaster2_p & !v9f7cc6;
assign d35a79 = hbusreq2_p & d35a70 | !hbusreq2_p & !d35a78;
assign c3d2b1 = hmaster2_p & c3d2b0 | !hmaster2_p & v845542;
assign df511c = decide_p & df511b | !decide_p & v845542;
assign v9ea45a = hbusreq4_p & v9ea458 | !hbusreq4_p & v9ea459;
assign c3d714 = hgrant1_p & c3d699 | !hgrant1_p & c3d70c;
assign ad3cf8 = hbusreq4_p & ad3cf6 | !hbusreq4_p & ad3cf7;
assign ad3d5f = jx0_p & ad437b | !jx0_p & ad3d5e;
assign cc36fc = hgrant0_p & v84556c | !hgrant0_p & !v845542;
assign c3d5ea = hbusreq0 & c3d5e9 | !hbusreq0 & v845542;
assign v9ea408 = hmaster1_p & v9ea407 | !hmaster1_p & v9ea405;
assign b059fb = hbusreq2 & b059f9 | !hbusreq2 & b059fa;
assign b05a25 = hgrant1_p & b0593d | !hgrant1_p & b05a14;
assign c5c892 = hlock3_p & c5c891 | !hlock3_p & v845542;
assign ad415a = hmaster2_p & ad4159 | !hmaster2_p & ad4153;
assign ad455e = hmaster2_p & v845542 | !hmaster2_p & ad455d;
assign ad4fd4 = hbusreq3 & ad4fd3 | !hbusreq3 & v845542;
assign ad4dab = hmaster2_p & ad4da9 | !hmaster2_p & ad4daa;
assign ade554 = hgrant4_p & v84556c | !hgrant4_p & !ade553;
assign d3552a = hbusreq1_p & d35519 | !hbusreq1_p & d35529;
assign v9e9f64 = stateA1_p & v9ea3e4 | !stateA1_p & v845542;
assign ad4427 = hbusreq1 & ad438f | !hbusreq1 & v845542;
assign b1c7d9 = hgrant4_p & b1c7d8 | !hgrant4_p & !b1c79d;
assign ad4f57 = hready & ad4e90 | !hready & ad4ea6;
assign ad4687 = hbusreq2 & ad4570 | !hbusreq2 & v845542;
assign c3d387 = hgrant3_p & c3d2e3 | !hgrant3_p & c3d386;
assign v9f7d3f = hbusreq1_p & v9f7d3d | !hbusreq1_p & v9f7d3e;
assign c5c893 = decide_p & c5c892 | !decide_p & c5c891;
assign dc4fff = hgrant4_p & c3d66d | !hgrant4_p & adec89;
assign ad436f = hmaster1_p & ad436e | !hmaster1_p & ad431c;
assign c3d71b = hgrant3_p & c3d6a1 | !hgrant3_p & c3d71a;
assign d358eb = hmastlock_p & d358ea | !hmastlock_p & v845542;
assign v8cc11e = hgrant2_p & v8cc0f5 | !hgrant2_p & v8cc0e9;
assign df5190 = hmaster0_p & df518a | !hmaster0_p & df518f;
assign c3d5df = hgrant4_p & v845542 | !hgrant4_p & !c3d5d4;
assign dc4fa6 = hbusreq4_p & dc4f9d | !hbusreq4_p & !v845542;
assign ad47ee = hbusreq2 & ad458b | !hbusreq2 & !v845542;
assign ade591 = hlock0_p & ade590 | !hlock0_p & !ade562;
assign v9f76dc = hmaster0_p & v9f7d34 | !hmaster0_p & v9f7e01;
assign v9f7d2f = hmaster0_p & v9f7d1f | !hmaster0_p & v9f7d2e;
assign ad4fd6 = hgrant4_p & ad4fca | !hgrant4_p & !v84556c;
assign c3d671 = hmaster2_p & c3d66a | !hmaster2_p & c3d670;
assign ad5033 = hmaster2_p & v845542 | !hmaster2_p & ad5032;
assign d3549f = hbusreq1 & d35bed | !hbusreq1 & d35be8;
assign dc53d0 = hgrant3_p & dc53cd | !hgrant3_p & !dc53cf;
assign c3d2b8 = hbusreq2 & c3d2b4 | !hbusreq2 & c3d2b7;
assign b573f6 = hgrant2_p & b573e8 | !hgrant2_p & b573df;
assign ad43fd = hmaster1_p & ad43d8 | !hmaster1_p & ad43fc;
assign df5197 = hmaster0_p & df5193 | !hmaster0_p & df5196;
assign v9f7e2c = hbusreq2 & v9f7e2a | !hbusreq2 & v9f7e2b;
assign dc4fb1 = hbusreq3 & dc4fb0 | !hbusreq3 & v845542;
assign adec8a = hbusreq4_p & adec89 | !hbusreq4_p & v845542;
assign v9f7cc1 = hlock2 & v9f7cb7 | !hlock2 & v9f7cc0;
assign v9f785e = hmaster2_p & v9f785d | !hmaster2_p & v9f772f;
assign c3cf24 = hmaster0_p & c3d2d7 | !hmaster0_p & c3d369;
assign dc53cd = hready_p & dc4f64 | !hready_p & !dc53cc;
assign ad43a5 = hmaster2_p & b1c70e | !hmaster2_p & ad43a4;
assign dc53b5 = hbusreq3_p & dc53b4 | !hbusreq3_p & !dc5088;
assign ad4162 = hmaster1_p & ad414b | !hmaster1_p & ad4161;
assign ad502a = hgrant1_p & ad501b | !hgrant1_p & ad5029;
assign d35908 = hburst1 & d35907 | !hburst1 & v845566;
assign df516a = hmaster0_p & df515a | !hmaster0_p & df5169;
assign b57a68 = hlock0 & b57942 | !hlock0 & b57a67;
assign c3d38f = hbusreq1_p & v84554d | !hbusreq1_p & !c3d2de;
assign df5186 = hmaster1_p & df517c | !hmaster1_p & df5185;
assign b57ae1 = hready_p & b578f5 | !hready_p & b57ae0;
assign ade5bd = hbusreq3 & ade56f | !hbusreq3 & !ade574;
assign d35708 = hlock1_p & d35707 | !hlock1_p & d35a6a;
assign v8cc786 = hbusreq3 & v8cc766 | !hbusreq3 & v8ccbd8;
assign v9f7858 = hmaster0_p & v9f7779 | !hmaster0_p & v9f7772;
assign bd5738 = hburst0_p & v845542 | !hburst0_p & bd5737;
assign d3549e = hmaster1_p & d3549a | !hmaster1_p & d3549d;
assign v9ea5a4 = hgrant1_p & v9ea578 | !hgrant1_p & v9ea5a3;
assign v9ea5b7 = hgrant2_p & v9ea5b3 | !hgrant2_p & v9ea5b6;
assign aa425e = jx1_p & v857463 | !jx1_p & v845542;
assign c5c970 = stateG10_4_p & c5c96e | !stateG10_4_p & c5c96f;
assign d35a4b = hgrant1_p & df54f3 | !hgrant1_p & d35a4a;
assign ad4f23 = hmaster1_p & ad4f1c | !hmaster1_p & ad4f22;
assign b1c051 = hmaster1_p & b1c050 | !hmaster1_p & b1c7e3;
assign b05a76 = hbusreq3 & b05a72 | !hbusreq3 & b05a75;
assign d3564e = hlock4_p & d3564c | !hlock4_p & !d3564d;
assign v9ea5cb = hmaster2_p & v9ea570 | !hmaster2_p & v9ea585;
assign c3ceed = hbusreq0_p & c3d5d4 | !hbusreq0_p & v84556e;
assign b1c7ee = hlock2_p & b1c7e5 | !hlock2_p & b1c7ed;
assign ad4fc7 = stateG2_p & v845542 | !stateG2_p & ad4fc6;
assign v9f7d0a = hready & v9f7d09 | !hready & v9f7d05;
assign decide = !ad3d60;
assign d3591c = hbusreq0 & d35919 | !hbusreq0 & d3591b;
assign c3d711 = hgrant2_p & c3d708 | !hgrant2_p & c3d710;
assign ad3cf7 = stateG10_4_p & ad3ceb | !stateG10_4_p & ad3cf6;
assign d354ac = hmastlock_p & ade54b | !hmastlock_p & v845542;
assign ad484c = hbusreq2 & ad4d93 | !hbusreq2 & v845542;
assign c3d71d = hmaster1_p & c3d71c | !hmaster1_p & c3d68b;
assign ad48b3 = hbusreq2 & ad48b2 | !hbusreq2 & !v845542;
assign v9ea42f = hbusreq4_p & v9ea418 | !hbusreq4_p & v9ea42e;
assign v8cc4b8 = hlock2 & v8ccbd8 | !hlock2 & v8cc4b6;
assign b57a22 = decide_p & b57a21 | !decide_p & b57944;
assign v9ea462 = hgrant4_p & v9f20a1 | !hgrant4_p & v9ea445;
assign d359b4 = hburst0_p & v845542 | !hburst0_p & !bbb31e;
assign c3cdf9 = hmaster0_p & c3d5ed | !hmaster0_p & c3d5f5;
assign v8cc820 = hready_p & v8cc81f | !hready_p & v8cc4f6;
assign v9ea3ec = hmastlock_p & v9ea3e4 | !hmastlock_p & v845542;
assign ad4ecc = hbusreq0_p & v845542 | !hbusreq0_p & ad4e53;
assign ad4de6 = hmaster0_p & v845555 | !hmaster0_p & ad4de5;
assign ade561 = hbusreq4_p & ade560 | !hbusreq4_p & !v845542;
assign d3590c = stateA1_p & v845542 | !stateA1_p & !adea85;
assign v9ea474 = hmaster2_p & v9ea467 | !hmaster2_p & v9ea473;
assign d355a4 = hburst1_p & v845568 | !hburst1_p & !v845542;
assign b57a10 = hready_p & b5799c | !hready_p & b57a0f;
assign ad4715 = hgrant4_p & v845542 | !hgrant4_p & ad4fe6;
assign v9f7ccf = hbusreq1 & v9f7ccd | !hbusreq1 & v9f7cce;
assign b57418 = stateG10_4_p & v845542 | !stateG10_4_p & b57417;
assign d35753 = hbusreq1_p & d35708 | !hbusreq1_p & d35aac;
assign b1d011 = hmaster0_p & b1d00e | !hmaster0_p & b1d010;
assign b1c054 = hmaster0_p & b1c053 | !hmaster0_p & b1c7e7;
assign b059c4 = hlock0 & b058a8 | !hlock0 & b059c3;
assign v8cc5a8 = hlock0 & v8cc494 | !hlock0 & v8cc5a7;
assign v9f7e0f = hmaster1_p & v9f7e0e | !hmaster1_p & v9f7df7;
assign b05a22 = hgrant2_p & b05a04 | !hgrant2_p & b05a21;
assign v8ccbe1 = hgrant0_p & v845542 | !hgrant0_p & v8ccb6a;
assign adec8f = hburst0 & adec8c | !hburst0 & adec8e;
assign v8cc76c = hmaster0_p & v845542 | !hmaster0_p & v8cc76b;
assign v9e9e74 = hmaster1_p & v9f20a1 | !hmaster1_p & v9ea4af;
assign d357ed = hbusreq1_p & v84554a | !hbusreq1_p & d357ec;
assign d35521 = hmaster2_p & d35520 | !hmaster2_p & d35a9b;
assign b058f3 = hbusreq3 & b058f1 | !hbusreq3 & b058f2;
assign c3d721 = hmaster0_p & c3d6e9 | !hmaster0_p & c3d671;
assign b1c7e4 = hmaster1_p & b1c7af | !hmaster1_p & b1c7e3;
assign b579c7 = hlock2 & b579c5 | !hlock2 & b579c6;
assign df5117 = hlock1_p & df5116 | !hlock1_p & v845542;
assign v9f78aa = hbusreq2_p & v9f78a7 | !hbusreq2_p & v9f78a9;
assign ad443f = hbusreq1 & ad4399 | !hbusreq1 & v845542;
assign ad3d12 = hmaster0_p & ad3cfe | !hmaster0_p & ad3d11;
assign b05918 = hlock3_p & b058e5 | !hlock3_p & b05917;
assign v84554c = hbusreq1_p & v845542 | !hbusreq1_p & !v845542;
assign c6d406 = stateG3_0_p & v845542 | !stateG3_0_p & c6d405;
assign d35630 = hbusreq2_p & d3562f | !hbusreq2_p & d35a97;
assign b57a69 = hbusreq0 & b57a67 | !hbusreq0 & b57a68;
assign v9ea489 = hbusreq2 & v9ea487 | !hbusreq2 & v9ea488;
assign d3568e = hmaster2_p & d35643 | !hmaster2_p & v845542;
assign bd5749 = hmaster2_p & bd572e | !hmaster2_p & v845542;
assign v9f783c = hlock2 & v9f7839 | !hlock2 & v9f783b;
assign v9f77c5 = hgrant4_p & v9f772b | !hgrant4_p & v9f77c4;
assign ad42fa = hmaster1_p & ad42ee | !hmaster1_p & ad42f9;
assign ad3d11 = hgrant1_p & ad4418 | !hgrant1_p & ad3d10;
assign d35758 = hbusreq2_p & d35747 | !hbusreq2_p & !d35757;
assign v9f7cbe = hbusreq1 & v9f7cbc | !hbusreq1 & v9f7cbd;
assign ad469a = hlock4_p & ad4ea2 | !hlock4_p & v845542;
assign ad5059 = hgrant4_p & ad5032 | !hgrant4_p & v845542;
assign ad4ded = hmaster2_p & ad4de2 | !hmaster2_p & ad4dde;
assign v9f7791 = hmaster2_p & v9f7785 | !hmaster2_p & !v845542;
assign b5740e = hready & b5740d | !hready & b578f1;
assign c3d2c6 = hmaster2_p & c3d2c5 | !hmaster2_p & v845542;
assign ade5c2 = hmaster0_p & ade5c0 | !hmaster0_p & ade5c1;
assign bd5798 = hmaster0_p & bd5795 | !hmaster0_p & bd5797;
assign b1cffa = hgrant4_p & v845542 | !hgrant4_p & b1cff9;
assign c3d341 = hgrant4_p & v845542 | !hgrant4_p & !c3d336;
assign ba7c7c = hgrant2_p & v845558 | !hgrant2_p & ba7c7b;
assign v8cc43b = hmaster0_p & v8cc435 | !hmaster0_p & v8cc43a;
assign v9f76be = hmaster0_p & v9f7d3e | !hmaster0_p & v9f7d3b;
assign v9f77e0 = hgrant1_p & v9f77d6 | !hgrant1_p & v9f77df;
assign ad431f = hbusreq1 & ad4fd0 | !hbusreq1 & v845542;
assign bd5912 = hlock1_p & bd5911 | !hlock1_p & df54f5;
assign b1c78c = hbusreq2 & b1c713 | !hbusreq2 & b1c718;
assign v8cc12b = hready_p & v8cc4e0 | !hready_p & v8cc12a;
assign b1c7cf = hgrant4_p & b1c711 | !hgrant4_p & !b1c79d;
assign ad4376 = decide_p & ad436b | !decide_p & ad4375;
assign b57a11 = hgrant3_p & b57946 | !hgrant3_p & b57a10;
assign d356f0 = hlock3_p & d356ea | !hlock3_p & d356ef;
assign c3d331 = hmaster0_p & c3d316 | !hmaster0_p & c3d330;
assign b1c849 = hbusreq1_p & b1cf2c | !hbusreq1_p & b1c848;
assign ad4efc = hmaster2_p & ad4ef6 | !hmaster2_p & ad4efb;
assign c3d6a3 = hmaster1_p & c3d6a2 | !hmaster1_p & c3d67c;
assign df5189 = hbusreq1_p & df5188 | !hbusreq1_p & v845542;
assign ad47e9 = hmaster0_p & ad47e8 | !hmaster0_p & ad4688;
assign v9f77db = hlock4 & v9f77d8 | !hlock4 & v9f77da;
assign ad45ba = hlock4_p & ade4bc | !hlock4_p & v845542;
assign v9ea584 = hmaster1_p & v9ea580 | !hmaster1_p & v9ea583;
assign b1c72f = hmaster1_p & b1c72e | !hmaster1_p & b1c72b;
assign c3d670 = locked_p & v845542 | !locked_p & !c3d66d;
assign ad3d5d = hbusreq3_p & ad3d21 | !hbusreq3_p & ad3d5c;
assign ad416e = hbusreq2_p & ad416d | !hbusreq2_p & v845542;
assign d35a3e = hburst1 & d35a3d | !hburst1 & v845542;
assign d357f9 = hmaster2_p & d3579d | !hmaster2_p & d35a9c;
assign v9ea3f5 = hmaster2_p & v9f20a1 | !hmaster2_p & v9ea3ec;
assign v9f7d2d = hlock2 & v9f7d23 | !hlock2 & !v9f7d2c;
assign ad481b = hbusreq2_p & ad481a | !hbusreq2_p & v845542;
assign c3d515 = hbusreq4 & c3d514 | !hbusreq4 & v845542;
assign ad3d18 = hgrant1_p & ad4413 | !hgrant1_p & ad3cf1;
assign ba7c67 = hmaster0_p & ba7c64 | !hmaster0_p & ba7c66;
assign d35ab0 = stateG10_4_p & d35aaa | !stateG10_4_p & !d35aab;
assign bd5e1d = hmaster2_p & v845542 | !hmaster2_p & bd5e1c;
assign b05a2d = hmaster0_p & b058e8 | !hmaster0_p & b05901;
assign d3572f = hbusreq3 & d3572e | !hbusreq3 & !d35aa4;
assign b579c0 = hready & b579bf | !hready & b57942;
assign ad4e22 = hbusreq3 & v845542 | !hbusreq3 & v845547;
assign ad46e6 = hgrant2_p & ad468d | !hgrant2_p & ad46e5;
assign c3d706 = decide_p & c3d6e0 | !decide_p & c3d705;
assign adeab3 = hready_p & v845542 | !hready_p & adeab2;
assign b1c7bf = stateG10_4_p & b1c7bc | !stateG10_4_p & b1c7be;
assign ad42e5 = hmaster0_p & ad42dd | !hmaster0_p & ad42e4;
assign v9ea407 = hmaster0_p & v9ea3fa | !hmaster0_p & v9ea3ff;
assign v9ea439 = locked_p & v9ea438 | !locked_p & v9ea3e6;
assign d35ab7 = hmaster1_p & d35aae | !hmaster1_p & d35ab6;
assign v8cc4ee = hmaster2_p & v8cc4ed | !hmaster2_p & v845542;
assign v9ea4be = hmaster1_p & v9ea4b5 | !hmaster1_p & v9ea4bd;
assign bd580d = hlock0_p & bd580b | !hlock0_p & !bd580c;
assign v9f7c98 = hmastlock_p & v9f7c97 | !hmastlock_p & !v845542;
assign v8cc590 = hmaster2_p & v845542 | !hmaster2_p & v8cc58f;
assign ade56f = hmaster2_p & ade548 | !hmaster2_p & !ade56e;
assign ad5032 = hmastlock_p & ad5031 | !hmastlock_p & v845542;
assign v8cc4dd = hready_p & v8cc455 | !hready_p & v8cc4dc;
assign v867d75 = jx1_p & v845542 | !jx1_p & !v845542;
assign v9f7817 = decide_p & v9f7802 | !decide_p & v9f7816;
assign ad42c2 = hbusreq1_p & ad42c1 | !hbusreq1_p & v845542;
assign ad4850 = hbusreq1_p & ad484f | !hbusreq1_p & ad4da1;
assign v9ea400 = hbusreq1_p & v9ea3fc | !hbusreq1_p & v9ea3ff;
assign dc5001 = hbusreq4_p & adec89 | !hbusreq4_p & dc5000;
assign ade551 = hgrant0_p & adec89 | !hgrant0_p & ade550;
assign b058a3 = hmastlock_p & b058a2 | !hmastlock_p & !v845542;
assign d35725 = hgrant3_p & d356f2 | !hgrant3_p & d35724;
assign ad47f5 = hmaster1_p & ad46f6 | !hmaster1_p & ad46e4;
assign ad42ed = hbusreq1_p & ad42ec | !hbusreq1_p & v845542;
assign df50d3 = decide_p & df507c | !decide_p & d6ebca;
assign ad4fa5 = hbusreq3 & ad4fa4 | !hbusreq3 & v845542;
assign d359f9 = hgrant4_p & d359e8 | !hgrant4_p & d359f7;
assign b059c0 = stateA1_p & b059bf | !stateA1_p & v857440;
assign c3cf0a = hbusreq2 & c3cf04 | !hbusreq2 & c3cf08;
assign bd5bb1 = hready_p & bd5baf | !hready_p & !bd5bb0;
assign ad4ee3 = hlock0_p & ad4ed7 | !hlock0_p & v845542;
assign d35a95 = hmaster2_p & v84555a | !hmaster2_p & v845542;
assign dc538c = locked_p & dc538b | !locked_p & v845542;
assign d35506 = hbusreq2_p & d354f0 | !hbusreq2_p & d35505;
assign ad4f2a = hbusreq1 & ad4e56 | !hbusreq1 & v845542;
assign v9ea498 = hmaster0_p & v9ea43a | !hmaster0_p & v9ea497;
assign ad4f95 = hbusreq4_p & ad4f94 | !hbusreq4_p & adeaa4;
assign c3cefe = decide_p & c3cefc | !decide_p & c3cefd;
assign d35514 = hlock1_p & d35513 | !hlock1_p & d3542e;
assign d358f2 = hlock1_p & d358f1 | !hlock1_p & v845542;
assign c3ce7e = hready_p & v845555 | !hready_p & c3ce7d;
assign c3d5be = hmaster2_p & c3d5bd | !hmaster2_p & v845576;
assign c3ce84 = hmaster1_p & c3ce80 | !hmaster1_p & c3ce83;
assign d358ea = stateA1_p & c5c894 | !stateA1_p & bb9bdd;
assign c3cf27 = hready_p & v845555 | !hready_p & !c3cf26;
assign b1c562 = hbusreq4_p & b1cff6 | !hbusreq4_p & !b1c857;
assign ade54d = hmastlock_p & ade54c | !hmastlock_p & v845542;
assign v9ea481 = hbusreq4 & v9ea47f | !hbusreq4 & v9ea480;
assign v8cc782 = hbusreq2_p & v8cc762 | !hbusreq2_p & v8cc781;
assign dc5067 = hmaster0_p & dc5030 | !hmaster0_p & dc5066;
assign d358f1 = hbusreq1 & v845542 | !hbusreq1 & d358f0;
assign ad435b = hready_p & ad4357 | !hready_p & !ad435a;
assign ad414d = hlock1_p & ad414c | !hlock1_p & !v845542;
assign ba7c6e = hmaster1_p & ba7c6b | !hmaster1_p & ba7c6d;
assign ad4e47 = locked_p & ad4e46 | !locked_p & v845542;
assign dc5008 = hbusreq0 & dc5002 | !hbusreq0 & dc5007;
assign v9f786c = hbusreq1_p & v9f7762 | !hbusreq1_p & v9f785e;
assign v9ea57c = hmaster1_p & v9ea57b | !hmaster1_p & v9ea579;
assign c3d584 = hgrant2_p & v845551 | !hgrant2_p & c3d583;
assign bd5e26 = decide_p & bd5e25 | !decide_p & v845542;
assign ac148d = hgrant1_p & ac145f | !hgrant1_p & ac148b;
assign v8da5a4 = hgrant1_p & v845542 | !hgrant1_p & !v8da5a1;
assign v8cc7e1 = hbusreq0 & v8cc7de | !hbusreq0 & v8cc7df;
assign c3d68a = hmaster2_p & c3d687 | !hmaster2_p & c3d689;
assign d35644 = hmaster2_p & d35643 | !hmaster2_p & d35a49;
assign b059e8 = hlock0 & b059e7 | !hlock0 & b059de;
assign ad41a0 = hmaster1_p & ad419d | !hmaster1_p & ad419f;
assign d356d4 = hbusreq1_p & d356d3 | !hbusreq1_p & v845542;
assign b059ed = hlock1 & b059e7 | !hlock1 & b059ec;
assign bd588c = hgrant4_p & ade572 | !hgrant4_p & !bd5842;
assign c3d47c = hready & c3d47a | !hready & c3d47b;
assign b1c07c = hbusreq1_p & b1c7cc | !hbusreq1_p & b1c07b;
assign v9f21c6 = hgrant0_p & v845542 | !hgrant0_p & v9f21c5;
assign d35794 = hbusreq0 & d35793 | !hbusreq0 & v845542;
assign ad4fde = stateG10_4_p & ad4fdc | !stateG10_4_p & ad4fdd;
assign d35620 = hgrant1_p & d3561f | !hgrant1_p & d35618;
assign ac1466 = hlock0_p & ac1465 | !hlock0_p & cc36fc;
assign v9e9f74 = hlock0_p & v9e9f73 | !hlock0_p & v9ea4c6;
assign b05a17 = hgrant4_p & b058a9 | !hgrant4_p & v9ea464;
assign ad4ffb = decide_p & ad4faa | !decide_p & ad4ffa;
assign df5182 = hbusreq1 & dc5064 | !hbusreq1 & v845542;
assign d35a60 = hlock4_p & d35a5e | !hlock4_p & !d35a5f;
assign b1c043 = hbusreq4_p & b1c770 | !hbusreq4_p & !b1c036;
assign ad4e7b = hbusreq0 & ad4e74 | !hbusreq0 & ad4e7a;
assign ade4a6 = hmaster2_p & adec8a | !hmaster2_p & adeca2;
assign v9f7df2 = hgrant1_p & v9f7df1 | !hgrant1_p & v9f7de7;
assign c5c904 = hgrant2_p & v845542 | !hgrant2_p & c5c902;
assign v8cc5b0 = hbusreq1 & v8cc5ab | !hbusreq1 & v8cc5ac;
assign c3d74f = hgrant2_p & c3d733 | !hgrant2_p & c3d74e;
assign c3d390 = hmaster0_p & c3d38f | !hmaster0_p & c3d2be;
assign c3ce98 = hmaster0_p & c3d35b | !hmaster0_p & c3d306;
assign b1c067 = hgrant4_p & b1c73c | !hgrant4_p & b1c066;
assign ad503f = hgrant0_p & ad502f | !hgrant0_p & v845542;
assign b1c5e2 = hmaster1_p & b1cfb8 | !hmaster1_p & b1c5e1;
assign ade4d1 = hmaster0_p & ade4cf | !hmaster0_p & ade4d0;
assign b579ea = hmaster1_p & b579b4 | !hmaster1_p & b579e9;
assign v9f76f9 = hbusreq1 & v9f76f7 | !hbusreq1 & v9f76f8;
assign c3d724 = hmaster1_p & c3d723 | !hmaster1_p & c3d67c;
assign d35417 = decide_p & d35416 | !decide_p & v84556c;
assign b059df = hgrant4_p & b058a7 | !hgrant4_p & !v9f7d42;
assign d35a75 = hbusreq3 & d35a74 | !hbusreq3 & v845542;
assign ade4d0 = hbusreq2 & ade4c7 | !hbusreq2 & ade4ce;
assign ad429a = hmaster1_p & ad4299 | !hmaster1_p & ad4297;
assign b0595a = hmaster2_p & b05952 | !hmaster2_p & b05959;
assign ad4151 = hbusreq4_p & ad4150 | !hbusreq4_p & v845542;
assign v8ccbfb = hlock2_p & v8ccbf9 | !hlock2_p & v8ccbfa;
assign v8cc769 = hlock2 & v8ccbd8 | !hlock2 & v8cc768;
assign b57a74 = hbusreq4_p & b579d2 | !hbusreq4_p & b579cd;
assign v9e9fa0 = hmaster1_p & v9e9f63 | !hmaster1_p & v9e9f9f;
assign b05a90 = hmaster0_p & b05a25 | !hmaster0_p & b05a0e;
assign ad4368 = hmaster1_p & ad4367 | !hmaster1_p & ad4300;
assign c3d2e5 = stateA1_p & v845542 | !stateA1_p & !v84557c;
assign c3d394 = hready_p & v845555 | !hready_p & c3d393;
assign b1c7ab = hbusreq4_p & b1c7a8 | !hbusreq4_p & !b1c7aa;
assign d35999 = hgrant4_p & v84557a | !hgrant4_p & !d35997;
assign c3d312 = hbusreq0 & v845576 | !hbusreq0 & c3d2fd;
assign d3597f = locked_p & v845542 | !locked_p & !v84557a;
assign ad4f75 = hgrant4_p & v845542 | !hgrant4_p & ad4f67;
assign dc5049 = hbusreq4_p & dc5046 | !hbusreq4_p & dc5048;
assign ad4ea6 = hbusreq4 & ad4ea1 | !hbusreq4 & ad4ea5;
assign ad4406 = hmaster0_p & ad4403 | !hmaster0_p & ad43fe;
assign v8cc7fa = hmaster2_p & v8cc7f1 | !hmaster2_p & v8cc7f9;
assign ad4db0 = hmaster2_p & ad4dac | !hmaster2_p & !ad4daf;
assign bd58e7 = hbusreq3 & bd5839 | !hbusreq3 & !dc501a;
assign d356da = hbusreq3 & d356d4 | !hbusreq3 & d356d9;
assign d359d2 = stateG10_4_p & d359ce | !stateG10_4_p & d359d0;
assign b579d4 = hlock0 & b579ce | !hlock0 & b579d3;
assign v9f781c = stateG10_4_p & v9f781a | !stateG10_4_p & v9f781b;
assign b1c58b = hgrant1_p & b1c58a | !hgrant1_p & b1cf28;
assign ad4751 = hmaster0_p & ad460b | !hmaster0_p & ad473d;
assign v8cc7e8 = hgrant1_p & v8cc7e7 | !hgrant1_p & v8ccbe3;
assign c3d360 = hmaster0_p & c3d35e | !hmaster0_p & c3d354;
assign v9e9fa1 = hgrant2_p & v9e9f4a | !hgrant2_p & v9e9fa0;
assign d3565e = decide_p & d3565d | !decide_p & v84556c;
assign d35aaa = hlock0_p & v845542 | !hlock0_p & v845548;
assign v8ccb8f = hlock2_p & v8ccb8c | !hlock2_p & v8ccb8d;
assign v9ea60e = hmaster0_p & v9ea60a | !hmaster0_p & v9ea60d;
assign c3cece = hbusreq0 & c3ceca | !hbusreq0 & c3cecd;
assign df5130 = hbusreq2_p & df512a | !hbusreq2_p & df553e;
assign d35992 = hbusreq1 & v84557a | !hbusreq1 & !v845542;
assign b574d7 = hmaster0_p & v845542 | !hmaster0_p & b574d6;
assign v9f7688 = decide_p & v9f7e11 | !decide_p & v9f7687;
assign ad42f5 = hbusreq1 & ad4f9b | !hbusreq1 & v845542;
assign dc4f69 = hbusreq3 & dc4f68 | !hbusreq3 & v845542;
assign ad42b7 = hbusreq0 & ad42b5 | !hbusreq0 & ad42b6;
assign b57a81 = hmaster0_p & b57a73 | !hmaster0_p & b57a80;
assign bd58b4 = hbusreq2 & bd58b3 | !hbusreq2 & v845542;
assign c5c9ad = hmaster1_p & c5c9ac | !hmaster1_p & c5c8eb;
assign d35986 = hbusreq3 & d35985 | !hbusreq3 & v845542;
assign ad4317 = hbusreq1_p & ad4316 | !hbusreq1_p & v845542;
assign c3d2b5 = hmaster2_p & c3d2b0 | !hmaster2_p & !v845542;
assign v8cc75b = hlock3 & v8cc4ad | !hlock3 & v8cc759;
assign bd58db = decide_p & bd58da | !decide_p & v845572;
assign v9f7e3e = hbusreq4_p & v9f7e3c | !hbusreq4_p & v9f7e3d;
assign d35508 = hlock4_p & v845542 | !hlock4_p & !d35955;
assign d356a2 = hmastlock_p & d359b9 | !hmastlock_p & d355a5;
assign ad4296 = hbusreq1_p & ad4295 | !hbusreq1_p & v845542;
assign v9f7dde = hgrant0_p & v9f7cf7 | !hgrant0_p & v9ea3ec;
assign b059b5 = hbusreq4 & b059b3 | !hbusreq4 & b059b4;
assign v8cc766 = hlock3 & v8ccbd8 | !hlock3 & v8cc765;
assign d35a64 = hlock0_p & d35a63 | !hlock0_p & ade562;
assign ad42f4 = hbusreq1 & ad4f13 | !hbusreq1 & v845542;
assign b1cc04 = hgrant2_p & v845542 | !hgrant2_p & b1cc03;
assign c5c8ef = hmaster0_p & v845542 | !hmaster0_p & c5c88f;
assign dc4f97 = hgrant2_p & dc4f94 | !hgrant2_p & dc4f96;
assign ac144e = locked_p & v845566 | !locked_p & !v845542;
assign d356b3 = hbusreq1_p & d356b2 | !hbusreq1_p & v845542;
assign ac1468 = stateG10_4_p & ac1466 | !stateG10_4_p & !ac1467;
assign c3d743 = hbusreq4_p & c3d6a7 | !hbusreq4_p & c3d742;
assign ad4f43 = hmaster0_p & ad4f33 | !hmaster0_p & ad4f42;
assign ad44b7 = hgrant1_p & ad43b9 | !hgrant1_p & ad44b6;
assign d357f2 = hbusreq0_p & dc5318 | !hbusreq0_p & v845542;
assign v8cc4a5 = hbusreq0 & v8cc4a3 | !hbusreq0 & v8cc4a4;
assign ad4565 = hmaster2_p & v845542 | !hmaster2_p & ad4564;
assign d357d6 = hgrant4_p & d3576f | !hgrant4_p & d3576e;
assign v845582 = stateG3_2_p & v845542 | !stateG3_2_p & !v845542;
assign v9e9f54 = hgrant4_p & v9e9ee7 | !hgrant4_p & v9ea441;
assign c3cec0 = hmaster2_p & c3cebf | !hmaster2_p & v845542;
assign df5540 = decide_p & df553f | !decide_p & d6ebca;
assign v9e9fe4 = hready_p & v9ea435 | !hready_p & v9e9fe3;
assign v9f7ca3 = stateA1_p & v845542 | !stateA1_p & !v9f7ca2;
assign d35aa6 = hmaster0_p & d35aa5 | !hmaster0_p & v845542;
assign bd57be = stateA1_p & bd57ba | !stateA1_p & bd57bd;
assign c3d2ea = hgrant0_p & v845542 | !hgrant0_p & c3d2e9;
assign c3d67a = hlock0_p & c3d670 | !hlock0_p & c3d679;
assign v9f7df9 = hgrant2_p & v9f7d6c | !hgrant2_p & v9f7df8;
assign v9ea5f4 = hmaster1_p & v9ea5f3 | !hmaster1_p & v9ea4af;
assign ac146d = hmaster1_p & ac145d | !hmaster1_p & ac146c;
assign v9e9ea3 = hgrant1_p & v9ea4cd | !hgrant1_p & v9e9ea2;
assign v9f7cb6 = locked_p & v9f7cb3 | !locked_p & v9ea3ec;
assign ad471c = hmaster1_p & ad4706 | !hmaster1_p & ad471b;
assign c3d36e = stateG2_p & v845542 | !stateG2_p & !d359ba;
assign b1c732 = hmaster2_p & b1c731 | !hmaster2_p & ade589;
assign b57404 = hgrant3_p & b57401 | !hgrant3_p & b57403;
assign b1c7d8 = hlock0_p & bd587d | !hlock0_p & b1c7d7;
assign v9ea5de = hmaster0_p & v9ea581 | !hmaster0_p & v9ea3fa;
assign ad476f = hlock1_p & ad476e | !hlock1_p & ad45ca;
assign ad45e6 = hlock0_p & ad4de2 | !hlock0_p & !v845542;
assign dc53b4 = hgrant3_p & dc53aa | !hgrant3_p & !dc53b3;
assign c3d4fa = hbusreq4_p & c3d4f9 | !hbusreq4_p & v845542;
assign ad4702 = hbusreq4 & ad4701 | !hbusreq4 & v845542;
assign b5743d = hmaster0_p & v845542 | !hmaster0_p & b579bb;
assign v9ea4d3 = hgrant0_p & v9ea4b3 | !hgrant0_p & v9ea4a6;
assign v9f770e = hmaster0_p & v9f7683 | !hmaster0_p & v9f7e2c;
assign ac1476 = hbusreq4_p & ac1461 | !hbusreq4_p & !ac1475;
assign ad4dd2 = hbusreq0 & ad4db3 | !hbusreq0 & ad4dd1;
assign b8f743 = hgrant2_p & v845542 | !hgrant2_p & !b8f6e1;
assign b57a7c = hgrant1_p & v845542 | !hgrant1_p & b57a7b;
assign ad3d44 = hmaster1_p & ad3d43 | !hmaster1_p & ad3cbb;
assign v9e9fcb = hready_p & v9ea436 | !hready_p & v9e9fca;
assign v9e9fdf = hgrant2_p & v9e9e68 | !hgrant2_p & v9e9fde;
assign df513a = hburst0 & adea98 | !hburst0 & adec98;
assign dc4fbb = hbusreq0 & dc4fa8 | !hbusreq0 & dc4fba;
assign c3cf04 = hgrant1_p & v845564 | !hgrant1_p & c3cf03;
assign d35777 = hbusreq3 & d35771 | !hbusreq3 & d35776;
assign b573f8 = decide_p & b57940 | !decide_p & b573f7;
assign b579be = hlock4 & b57942 | !hlock4 & b579bd;
assign b1c73c = hlock0_p & c3d674 | !hlock0_p & v845542;
assign ad475a = hmaster1_p & ad4759 | !hmaster1_p & ad4591;
assign c3d3a5 = hgrant1_p & v84554d | !hgrant1_p & c3d3a4;
assign c3d528 = hmaster2_p & c3d523 | !hmaster2_p & !v845542;
assign v8cc7dd = locked_p & v8cc7dc | !locked_p & v845542;
assign b1c865 = hbusreq2_p & b1c854 | !hbusreq2_p & b1c864;
assign b1cbf5 = hmaster2_p & b1cfcc | !hmaster2_p & b1cbf4;
assign dc5080 = hgrant2_p & dc5077 | !hgrant2_p & dc507f;
assign c3d375 = hmaster2_p & c3d374 | !hmaster2_p & !v845542;
assign v9f7e2b = hlock2 & v9f7e28 | !hlock2 & v9f7e2a;
assign b058a8 = hmaster2_p & b058a3 | !hmaster2_p & !b058a7;
assign b05945 = hmaster0_p & b0593a | !hmaster0_p & b0593d;
assign v8cc7f9 = hgrant4_p & v845542 | !hgrant4_p & v8cc7f8;
assign v9f77d7 = hmaster2_p & v9f77c1 | !hmaster2_p & v9f772f;
assign d354d5 = hgrant2_p & d3549e | !hgrant2_p & d354d4;
assign b05a64 = hbusreq0_p & b0594f | !hbusreq0_p & b05a63;
assign d3550f = hlock4_p & d358f9 | !hlock4_p & !d3594e;
assign ade5ad = hbusreq2 & ade5ac | !hbusreq2 & !v845558;
assign dc4faf = hbusreq0 & dc4fad | !hbusreq0 & dc4fae;
assign c3d5f5 = hbusreq2 & c3d5f4 | !hbusreq2 & c3d5ec;
assign ad5064 = hgrant1_p & ad501b | !hgrant1_p & ad5063;
assign v9f7cf6 = hmaster2_p & v9f7c9b | !hmaster2_p & v9f7cf5;
assign ad4341 = hmaster1_p & ad4337 | !hmaster1_p & ad4340;
assign ad4eb4 = hgrant4_p & ad4e54 | !hgrant4_p & ad4eb3;
assign v9e9f9f = hmaster0_p & v9e9f88 | !hmaster0_p & v9e9f9e;
assign v9f787d = hgrant2_p & v9f787c | !hgrant2_p & v9f7879;
assign ad46b8 = hbusreq4_p & ad46b7 | !hbusreq4_p & v845542;
assign ad432e = hbusreq1_p & ad432d | !hbusreq1_p & v845547;
assign v9e9ecd = hmaster1_p & v9e9ecc | !hmaster1_p & v9e9e77;
assign b1c7c5 = stateG10_4_p & b1c7bc | !stateG10_4_p & b1c7c4;
assign c3d6b7 = hgrant0_p & c3d675 | !hgrant0_p & c3d674;
assign ad4353 = hmaster1_p & ad4352 | !hmaster1_p & ad4297;
assign df518c = hbusreq1_p & df518b | !hbusreq1_p & v845542;
assign ad4479 = hgrant4_p & b1c70e | !hgrant4_p & c3cec2;
assign c3d6f7 = hgrant4_p & c3d67a | !hgrant4_p & !c3d6f6;
assign v9e9ef3 = hmaster0_p & v9e9ee8 | !hmaster0_p & v9e9eed;
assign v9f76e4 = hbusreq0_p & v9f7d71 | !hbusreq0_p & v9f76e3;
assign df50ce = hgrant1_p & df50cd | !hgrant1_p & !v845542;
assign ade625 = hbusreq2_p & ade623 | !hbusreq2_p & ade624;
assign b05a6d = hbusreq4 & b05a6b | !hbusreq4 & b05a6c;
assign v9f77f9 = hgrant1_p & v9f7730 | !hgrant1_p & v9f77de;
assign b1d001 = hmaster2_p & b1cfbf | !hmaster2_p & b1d000;
assign c3cec7 = hbusreq0 & c3cec0 | !hbusreq0 & c3cec6;
assign b05a10 = hbusreq1_p & b0593a | !hbusreq1_p & b05a0f;
assign ad4306 = hmaster0_p & ad42fc | !hmaster0_p & ad4305;
assign v8cc7b1 = hbusreq1_p & v8cc7b0 | !hbusreq1_p & v845542;
assign bd579a = hmaster2_p & bd5786 | !hmaster2_p & ade4df;
assign v9f7724 = hbusreq3_p & v9f76b2 | !hbusreq3_p & v9f7723;
assign ad436e = hmaster0_p & ad4325 | !hmaster0_p & ad4315;
assign v9f76f4 = hbusreq0 & v9f76e9 | !hbusreq0 & v9f76f3;
assign v9f785f = hlock0 & v9f785e | !hlock0 & v9f7759;
assign d35a53 = hbusreq1_p & d35a52 | !hbusreq1_p & !v845542;
assign v9f7d05 = hmaster2_p & v9f7ca4 | !hmaster2_p & !v9ea3ec;
assign ad4748 = hbusreq4 & ad4747 | !hbusreq4 & v845542;
assign b57b5a = hbusreq3_p & b57aee | !hbusreq3_p & b57b59;
assign v9f7776 = hlock3 & v9f775a | !hlock3 & v9f7760;
assign b0590c = hready & b0590b | !hready & b058d5;
assign ad410b = hbusreq2 & ad410a | !hbusreq2 & v845542;
assign v9f76a5 = hgrant1_p & v9f7d63 | !hgrant1_p & v9f76a4;
assign b573e6 = hbusreq2 & b573e5 | !hbusreq2 & b57942;
assign v9f7cfa = hbusreq0 & v9f7cf6 | !hbusreq0 & v9f7cf9;
assign v9f7832 = hlock4 & v9f782f | !hlock4 & v9f7831;
assign b1c56c = hgrant2_p & b1d01a | !hgrant2_p & b1c56b;
assign ad5047 = hmastlock_p & ad5046 | !hmastlock_p & v845542;
assign b1c060 = hbusreq1_p & b1c7f2 | !hbusreq1_p & b1c05f;
assign v845558 = hbusreq4_p & v845542 | !hbusreq4_p & !v845542;
assign d359c7 = hlock1_p & d359c3 | !hlock1_p & !d359c6;
assign b57943 = hmaster0_p & b57942 | !hmaster0_p & v845542;
assign ad4f09 = hgrant4_p & v845542 | !hgrant4_p & ad4ef7;
assign v9f7781 = hmaster0_p & v9f7772 | !hmaster0_p & v9f7779;
assign ad42c3 = hbusreq2 & ad42bf | !hbusreq2 & ad42c2;
assign v9ea41f = hgrant0_p & v9ea414 | !hgrant0_p & v845542;
assign d35700 = hlock1_p & d356fe | !hlock1_p & d356ff;
assign bd58f9 = hgrant1_p & bd58f8 | !hgrant1_p & bd5854;
assign b1c618 = hbusreq1_p & b1c617 | !hbusreq1_p & b1cf2c;
assign dc505f = hgrant4_p & v845542 | !hgrant4_p & !ade59c;
assign b05955 = hgrant4_p & b058b6 | !hgrant4_p & b05954;
assign b1c71e = hbusreq3 & b1c71c | !hbusreq3 & b1c71d;
assign b1c5bf = hgrant1_p & b1c5be | !hgrant1_p & b1c5b8;
assign v9e9f98 = hbusreq1 & v9e9f96 | !hbusreq1 & v9e9f97;
assign ad46b1 = hbusreq1 & ad4586 | !hbusreq1 & !v845547;
assign v857463 = hmaster1_p & v84554c | !hmaster1_p & v86cea1;
assign b579e0 = hbusreq4 & b579de | !hbusreq4 & b579df;
assign ad3d55 = hmaster1_p & ad3d54 | !hmaster1_p & ad4419;
assign dc53d9 = hready_p & dc53d6 | !hready_p & !dc53d8;
assign c3ce6f = hmaster0_p & c3ce6e | !hmaster0_p & !c3d2be;
assign b05a80 = hbusreq2 & b05a7e | !hbusreq2 & b05a7f;
assign ade5b3 = hbusreq1_p & ade5b1 | !hbusreq1_p & ade5b2;
assign b1c7d5 = hmaster2_p & b1c7d4 | !hmaster2_p & b1cfb7;
assign d359e9 = hmaster2_p & d359e6 | !hmaster2_p & d359e8;
assign d357ad = hmaster1_p & d357ac | !hmaster1_p & d357a6;
assign cc370a = hgrant3_p & cc36f0 | !hgrant3_p & !cc3709;
assign b57424 = hlock1 & b57987 | !hlock1 & b57423;
assign c3d337 = hgrant4_p & v845542 | !hgrant4_p & c3d336;
assign b1c041 = hmaster2_p & b1c040 | !hmaster2_p & !b1c844;
assign b059f5 = hmaster0_p & b059d3 | !hmaster0_p & b059f4;
assign b8f6e2 = hgrant1_p & v845542 | !hgrant1_p & c3d328;
assign df514b = hbusreq1_p & df514a | !hbusreq1_p & v845542;
assign v9f7e09 = hgrant1_p & v9f7e08 | !hgrant1_p & v9f7db4;
assign ad46fb = hmaster0_p & ad459e | !hmaster0_p & ad459d;
assign ad4342 = hgrant2_p & ad432c | !hgrant2_p & ad4341;
assign v9e9f62 = hlock2 & v9e9f5f | !hlock2 & v9e9f61;
assign d357a9 = hmaster1_p & d357a8 | !hmaster1_p & d357a6;
assign d357aa = hlock2_p & d357a7 | !hlock2_p & d357a9;
assign d35588 = hgrant1_p & d35586 | !hgrant1_p & d35587;
assign b05937 = hmastlock_p & b05936 | !hmastlock_p & !v845542;
assign v9ea5ab = hmaster1_p & v9ea44a | !hmaster1_p & v9ea5aa;
assign v9f77a4 = hlock1 & v9f779f | !hlock1 & v9f77a3;
assign b1c7b2 = hlock1_p & b1c7b0 | !hlock1_p & b1c7b1;
assign ad46bb = hbusreq4 & ad46ba | !hbusreq4 & v845542;
assign bd56d9 = hbusreq4 & bd56d6 | !hbusreq4 & bd56d8;
assign ad4fe3 = hbusreq4_p & v845542 | !hbusreq4_p & ad4fe2;
assign df5156 = hbusreq1 & dc4f68 | !hbusreq1 & v845542;
assign c3ce2e = decide_p & c3ce26 | !decide_p & !c3ce22;
assign ad4dd9 = hmaster1_p & ad4dc1 | !hmaster1_p & ad4db9;
assign c3d389 = hmaster0_p & v84554d | !hmaster0_p & c3d2be;
assign ad4322 = hmaster1_p & ad4321 | !hmaster1_p & ad4297;
assign ad459c = hbusreq4 & ad459b | !hbusreq4 & v845542;
assign c3ce59 = hmaster0_p & c3ce56 | !hmaster0_p & c3ce58;
assign v9ea595 = hgrant1_p & v9ea594 | !hgrant1_p & v9ea592;
assign d3562a = hmaster0_p & d35626 | !hmaster0_p & !d35629;
assign ad4e4e = hready & ad4e4b | !hready & ad4e4d;
assign b1c7b4 = hmaster2_p & b1c731 | !hmaster2_p & !b1c7b3;
assign v8cc4ad = hgrant1_p & v845542 | !hgrant1_p & v8cc494;
assign dc5034 = hbusreq1 & dc5033 | !hbusreq1 & !v845542;
assign d35a48 = hlock4_p & dc500e | !hlock4_p & !dc500f;
assign b8f6e6 = hready_p & b8f6e5 | !hready_p & v845562;
assign ad45ae = hburst0 & dc4f7a | !hburst0 & dc4f78;
assign v9ea45c = hbusreq1_p & v9ea449 | !hbusreq1_p & v9ea45b;
assign ad3cf6 = hlock0_p & c3d318 | !hlock0_p & ad4480;
assign ad4f55 = hbusreq1 & ad4f44 | !hbusreq1 & v845542;
assign d35696 = hgrant2_p & v845542 | !hgrant2_p & !d35695;
assign b57ae3 = hbusreq3 & b579c4 | !hbusreq3 & b57ae2;
assign ad4138 = hmaster2_p & ad4137 | !hmaster2_p & ad4f04;
assign v9e9f87 = hlock2 & v9e9f84 | !hlock2 & v9e9f86;
assign v9e9e68 = hmaster1_p & v9e9e67 | !hmaster1_p & v9ea405;
assign v9ea419 = hgrant4_p & v9ea414 | !hgrant4_p & v845542;
assign b57a6f = hgrant1_p & b57a6e | !hgrant1_p & b579b3;
assign ad3d2e = hmaster0_p & ad3d2b | !hmaster0_p & ad4413;
assign v9f7749 = hbusreq4 & v9f7747 | !hbusreq4 & v9f7748;
assign bd5904 = hbusreq3_p & bd58e6 | !hbusreq3_p & bd5903;
assign b1c4d0 = hmaster1_p & b1c842 | !hmaster1_p & b1c4cf;
assign d35a44 = hgrant4_p & v84556c | !hgrant4_p & d35a43;
assign c3d50c = hmaster1_p & c3d509 | !hmaster1_p & c3d50b;
assign bd57c9 = hbusreq1_p & bd57c7 | !hbusreq1_p & bd57c8;
assign v9f7d75 = hlock4_p & v9f7d73 | !hlock4_p & v9f7d74;
assign b5744f = hbusreq3_p & b57443 | !hbusreq3_p & b5744e;
assign v9ea430 = hgrant4_p & v845542 | !hgrant4_p & v9ea41c;
assign v9ea5f9 = decide_p & v9ea5f5 | !decide_p & v9ea5f8;
assign b1c77d = hmaster1_p & b1c77c | !hmaster1_p & b1c775;
assign ad45ee = hmaster2_p & v845542 | !hmaster2_p & ad45ed;
assign b57acd = hbusreq1_p & b578f9 | !hbusreq1_p & b57abf;
assign dc5020 = hmaster2_p & dc4fe6 | !hmaster2_p & dc501f;
assign d3571f = hmaster0_p & d35702 | !hmaster0_p & d3571e;
assign d35a6a = hbusreq0 & d35a62 | !hbusreq0 & d35a69;
assign b05a43 = hmaster0_p & b05a42 | !hmaster0_p & b05925;
assign df516b = hmaster1_p & df516a | !hmaster1_p & df5163;
assign v9f7dd4 = stateG10_4_p & v9f7dd0 | !stateG10_4_p & !v9f7dd2;
assign ad43a8 = hbusreq0 & ad43a7 | !hbusreq0 & v845542;
assign dc4fb5 = hmaster0_p & dc4f9a | !hmaster0_p & dc4fb4;
assign v9f7de6 = hbusreq4_p & v9f7de4 | !hbusreq4_p & v9f7de5;
assign ad4daa = hlock0_p & v9f21c4 | !hlock0_p & v845542;
assign c3d382 = hmaster1_p & c3d37d | !hmaster1_p & c3d381;
assign v9f7891 = hlock2 & v9f77fa | !hlock2 & v9f7890;
assign b05a1e = hmaster2_p & b05a1a | !hmaster2_p & b05a1d;
assign bd57cb = hbusreq3 & bd57c5 | !hbusreq3 & bd57ca;
assign v9ea457 = hgrant0_p & v9ea3fe | !hgrant0_p & v9ea3e6;
assign bd581f = stateG10_4_p & bd580d | !stateG10_4_p & !bd581e;
assign b57a7f = hlock2 & b579e5 | !hlock2 & b57a7e;
assign d35428 = hbusreq4 & d35427 | !hbusreq4 & d3541f;
assign ad3d05 = hbusreq0_p & ad5048 | !hbusreq0_p & v845542;
assign ade5bc = hgrant3_p & ade4f3 | !hgrant3_p & ade5bb;
assign b058fc = hlock1 & b058b8 | !hlock1 & b058fb;
assign v8cc4fa = hgrant4_p & v845542 | !hgrant4_p & v8cc4f9;
assign b1c802 = hbusreq0 & b1c7b4 | !hbusreq0 & d35a9c;
assign c3d6ce = stateG10_4_p & c3d6cb | !stateG10_4_p & c3d6cd;
assign c5c93b = hgrant1_p & v845542 | !hgrant1_p & !c5c93a;
assign d35a6e = hgrant2_p & d35a39 | !hgrant2_p & d35a6d;
assign b1c031 = hlock0_p & ade4d4 | !hlock0_p & v845542;
assign ad5040 = hbusreq0_p & ad503e | !hbusreq0_p & !ad503f;
assign cc36d9 = hmaster1_p & cc36d8 | !hmaster1_p & cc36c0;
assign c3ce85 = hgrant2_p & v845551 | !hgrant2_p & c3ce84;
assign ad4168 = hmaster0_p & ad4166 | !hmaster0_p & ad4167;
assign c3d678 = hbusreq4_p & c3d670 | !hbusreq4_p & c3d675;
assign b05997 = hready & b05996 | !hready & b05992;
assign ad4489 = hbusreq0_p & ad4fca | !hbusreq0_p & !v845542;
assign dc4fdf = hbusreq1 & dc4fc9 | !hbusreq1 & dc4fcb;
assign c3ce36 = hbusreq1 & c3d2b6 | !hbusreq1 & !v845542;
assign bd56e0 = hready_p & v845542 | !hready_p & bd56df;
assign c3cee3 = hbusreq0 & v845564 | !hbusreq0 & !v845542;
assign v9f7709 = hbusreq2 & v9f7707 | !hbusreq2 & v9f7708;
assign b1c611 = hready_p & b1c600 | !hready_p & b1c610;
assign ad4f1d = hmaster2_p & v84557a | !hmaster2_p & !ad4e53;
assign ad4689 = hmaster0_p & ad4687 | !hmaster0_p & ad4688;
assign v9e9eea = hmaster0_p & v9e9ee8 | !hmaster0_p & v9e9ee9;
assign v9f77f4 = hmaster0_p & v9f77e6 | !hmaster0_p & !v9f77f3;
assign ad42a7 = hbusreq2 & ad42a1 | !hbusreq2 & ad42a5;
assign v9f7dce = hgrant0_p & v9f7ca0 | !hgrant0_p & !v9f7c9f;
assign dc4fc3 = hmaster1_p & dc4fb5 | !hmaster1_p & dc4fb2;
assign b05a87 = hgrant2_p & b05a4e | !hgrant2_p & b05a86;
assign dc503f = stateG10_4_p & ade58d | !stateG10_4_p & dc503e;
assign b1c853 = hmaster1_p & b1cfb8 | !hmaster1_p & b1c852;
assign dc4f9f = hbusreq3 & dc4f9e | !hbusreq3 & v845542;
assign ad4784 = hlock2_p & ad4782 | !hlock2_p & ad4783;
assign ad4e75 = hgrant0_p & v845542 | !hgrant0_p & !ad4e6c;
assign bd5807 = hgrant4_p & bd572e | !hgrant4_p & bd5806;
assign v9f7d58 = hmastlock_p & v9f7d57 | !hmastlock_p & !v845542;
assign ad43bb = hmaster1_p & ad43ac | !hmaster1_p & ad43ba;
assign b57a2a = hmaster0_p & b57a29 | !hmaster0_p & b57956;
assign c3d478 = hbusreq4 & c3d2b1 | !hbusreq4 & !v845564;
assign b1caec = hbusreq4_p & b1caeb | !hbusreq4_p & !v84554a;
assign b05a8a = hmaster1_p & b059a9 | !hmaster1_p & b059f5;
assign ad40fb = decide_p & ad40f1 | !decide_p & ad40fa;
assign c3ceb7 = hmaster1_p & c3ceb3 | !hmaster1_p & c3ceb6;
assign v9ea3e3 = hmaster1_p & v9ea3e2 | !hmaster1_p & v845542;
assign ac1455 = hmaster0_p & v845542 | !hmaster0_p & ac144f;
assign bd5ba0 = hready_p & bd5b9d | !hready_p & !bd5b9f;
assign b1c75d = hbusreq3 & b1c758 | !hbusreq3 & b1c75c;
assign b058c2 = hlock3 & b058b8 | !hlock3 & b058c1;
assign ad4723 = hgrant2_p & ad471f | !hgrant2_p & ad4722;
assign c3d6e5 = stateG10_4_p & c3d6ab | !stateG10_4_p & c3d6e4;
assign dc5315 = decide_p & dc5314 | !decide_p & v845542;
assign v9e9f5e = hgrant1_p & v9e9ee9 | !hgrant1_p & v9e9f5d;
assign ad4f8b = stateG10_4_p & ad4f88 | !stateG10_4_p & !ad4f8a;
assign ad4e4c = hburst0 & dc52f8 | !hburst0 & bd5b85;
assign v8cc5ac = hlock1 & v8cc494 | !hlock1 & v8cc5ab;
assign v8cc829 = hmaster0_p & v8cc827 | !hmaster0_p & v8cc7ce;
assign ad40e7 = hmaster0_p & ad40ba | !hmaster0_p & !ad40e6;
assign v8cc81d = hmaster0_p & v8cc810 | !hmaster0_p & v845542;
assign b05a07 = hgrant4_p & b05939 | !hgrant4_p & b05a06;
assign b579b2 = hgrant4_p & v845542 | !hgrant4_p & b579b1;
assign c3d502 = hbusreq0 & v845542 | !hbusreq0 & c3d501;
assign v9f7839 = hgrant1_p & v9f772c | !hgrant1_p & v9f7838;
assign b0597a = hlock4_p & b05978 | !hlock4_p & !b05979;
assign v9f7ceb = hlock3 & v9f7cc8 | !hlock3 & v9f7ccf;
assign c5c8f1 = locked_p & c5c896 | !locked_p & !v845542;
assign ad4f67 = hlock0_p & ad4f36 | !hlock0_p & !v845542;
assign ad4fb0 = hready & ad4faf | !hready & dc4fcb;
assign b1c82d = decide_p & b1c82c | !decide_p & v845542;
assign bd5843 = hgrant4_p & bd574e | !hgrant4_p & bd5842;
assign v8cc0d8 = stateG10_4_p & v845542 | !stateG10_4_p & v8cc0d7;
assign b05962 = hbusreq1 & b05960 | !hbusreq1 & b05961;
assign ad4572 = hmaster0_p & ad456c | !hmaster0_p & ad4571;
assign c3cf18 = hgrant3_p & c3ceec | !hgrant3_p & c3cf17;
assign b059d3 = hbusreq2 & b059d1 | !hbusreq2 & b059d2;
assign v8cc43a = hgrant1_p & v845542 | !hgrant1_p & v8cc439;
assign v845548 = hbusreq0_p & v845542 | !hbusreq0_p & !v845542;
assign d35566 = hmaster0_p & d35565 | !hmaster0_p & d35499;
assign ad3ce7 = hready & ad3ce0 | !hready & !ad3ce6;
assign bd583f = hmaster2_p & bd5802 | !hmaster2_p & bd583e;
assign v8cc601 = decide_p & v8cc4f4 | !decide_p & v8cc5c6;
assign bd5937 = hmaster0_p & v84556c | !hmaster0_p & bd5936;
assign bd57c3 = hburst1 & bd57bf | !hburst1 & bd57c2;
assign cc3704 = hmaster0_p & cc36f8 | !hmaster0_p & cc3703;
assign bd5e1b = hlock4_p & bd5b6e | !hlock4_p & dc5318;
assign ad46d6 = hgrant4_p & v845542 | !hgrant4_p & ad46d5;
assign b05a65 = hlock0_p & b0594f | !hlock0_p & b05a64;
assign v9ea48c = hgrant2_p & v9ea440 | !hgrant2_p & v9ea48b;
assign v8cc0e8 = hmaster0_p & v8cc0d6 | !hmaster0_p & v8cc0e7;
assign v9ea43b = hmaster2_p & v9ea439 | !hmaster2_p & v9f20a1;
assign ac1486 = hlock0_p & ac1458 | !hlock0_p & ac1485;
assign v9f7cd9 = hmaster2_p & v9f7cd6 | !hmaster2_p & v9f7cd8;
assign d35616 = stateA1_p & ade4b8 | !stateA1_p & ade4b7;
assign cc36ca = hgrant4_p & v845542 | !hgrant4_p & !v84556c;
assign v9f773d = hmaster1_p & v9f773c | !hmaster1_p & v9f7736;
assign ad4dc4 = hburst0 & ad4dc3 | !hburst0 & d3561c;
assign v9e9fd7 = hready_p & v9ea435 | !hready_p & v9e9fd6;
assign ad4596 = hbusreq2_p & ad4592 | !hbusreq2_p & ad4595;
assign ade661 = hgrant3_p & ade658 | !hgrant3_p & ade660;
assign v9f7cbd = hlock1 & v9f7cb7 | !hlock1 & v9f7cbc;
assign b5743c = hgrant2_p & b579b0 | !hgrant2_p & b5743b;
assign v9f7d32 = hbusreq3 & v9f7d19 | !hbusreq3 & v9f7d31;
assign ad3ccc = hbusreq4_p & ad3cca | !hbusreq4_p & ad3ccb;
assign d354fd = hbusreq3 & d354fc | !hbusreq3 & !d354f5;
assign ac1482 = hgrant3_p & ac1454 | !hgrant3_p & ac1481;
assign b57940 = hlock3_p & b57906 | !hlock3_p & b5793f;
assign ad4142 = hbusreq0 & ad413d | !hbusreq0 & ad4141;
assign c3ce09 = hbusreq2_p & c3ce08 | !hbusreq2_p & c3ce01;
assign bd57c5 = hmaster2_p & bd57c4 | !hmaster2_p & !dc4f9d;
assign d35a09 = hmaster2_p & d35a00 | !hmaster2_p & d35a08;
assign v9f7647 = hlock1 & v9f7e3f | !hlock1 & v9f7646;
assign b574bf = hbusreq2 & b574bd | !hbusreq2 & b574be;
assign v9f7ca5 = locked_p & v9f7c98 | !locked_p & v9f7ca4;
assign v9f7d93 = hlock4 & v9f7d90 | !hlock4 & v9f7d92;
assign ad45e8 = hbusreq4_p & ad45e7 | !hbusreq4_p & !v845542;
assign bd5854 = hbusreq4 & bd5848 | !hbusreq4 & bd5853;
assign ade5dd = hbusreq2_p & ade5da | !hbusreq2_p & ade5dc;
assign ad4147 = hmaster0_p & ad4111 | !hmaster0_p & ad4146;
assign bd5830 = hgrant1_p & bd5828 | !hgrant1_p & bd582f;
assign b05a39 = hmaster1_p & b05a38 | !hmaster1_p & b05926;
assign ad4eee = hbusreq4_p & ad4ed3 | !hbusreq4_p & v845542;
assign bbb7c6 = hburst1_p & v845542 | !hburst1_p & v8f2540;
assign v9f774b = hbusreq1 & v9f7749 | !hbusreq1 & v9f774a;
assign d35423 = hbusreq4_p & d35422 | !hbusreq4_p & v845542;
assign ad4383 = hmaster2_p & ad4380 | !hmaster2_p & ad4382;
assign v9f7dc5 = hbusreq2 & v9f7dc3 | !hbusreq2 & v9f7dc4;
assign ad4e6e = hgrant0_p & v84557a | !hgrant0_p & ad4e6c;
assign cc36de = hmaster2_p & v845566 | !hmaster2_p & !cc36dd;
assign v9f76a3 = hbusreq4_p & v9f76a1 | !hbusreq4_p & v9f76a2;
assign b1c779 = hmaster1_p & b1c778 | !hmaster1_p & b1c775;
assign c3d306 = hgrant1_p & v84554d | !hgrant1_p & c3d305;
assign d3577f = decide_p & d3577e | !decide_p & v84556c;
assign c3ce9e = hmaster2_p & c3d30d | !hmaster2_p & v845542;
assign ad4fcc = stateA1_p & d35a3a | !stateA1_p & !v845542;
assign c3ce3d = hlock1_p & c3ce3b | !hlock1_p & c3ce3c;
assign v9f76db = hlock2_p & v9f76d7 | !hlock2_p & v9f76da;
assign d35715 = hgrant2_p & d35714 | !hgrant2_p & !d3570c;
assign dc4fb7 = hbusreq1_p & dc4fb6 | !hbusreq1_p & dc4fa3;
assign b57aba = hready_p & b57a2e | !hready_p & b57ab9;
assign v845555 = hbusreq3 & v845542 | !hbusreq3 & !v845542;
assign b1c825 = hbusreq3 & b1c768 | !hbusreq3 & b1c76a;
assign ade4aa = hlock0_p & adec89 | !hlock0_p & ade4a9;
assign ade627 = hready_p & ade621 | !hready_p & ade626;
assign v9e9fd0 = hmaster0_p & v9ea45e | !hmaster0_p & v9ea486;
assign b059cd = hgrant1_p & b059cb | !hgrant1_p & b059cc;
assign b57aca = hbusreq2 & b57ac9 | !hbusreq2 & b578f9;
assign ad45c4 = hbusreq1 & ad45b6 | !hbusreq1 & ad45c0;
assign c3ce4e = hmaster0_p & c3ce48 | !hmaster0_p & c3ce4d;
assign b059fd = hmaster1_p & b059fc | !hmaster1_p & b058e1;
assign v9f768d = hgrant4_p & v9f7d59 | !hgrant4_p & v9f768c;
assign v9f7d5d = locked_p & v845542 | !locked_p & !v9f7cc6;
assign c5c99e = hmaster0_p & c5c930 | !hmaster0_p & v845542;
assign v9ea49a = hgrant1_p & v9ea3ff | !hgrant1_p & v9ea45b;
assign b1c495 = hlock4_p & b1cf30 | !hlock4_p & b1cf3e;
assign ade4e4 = hmastlock_p & c3d66b | !hmastlock_p & v845542;
assign c3d5aa = hbusreq2 & c3d5a9 | !hbusreq2 & c3d2de;
assign b058f6 = hbusreq2 & b058f3 | !hbusreq2 & b058f5;
assign v9e9f7c = hbusreq4 & v9e9f7a | !hbusreq4 & v9e9f7b;
assign v8cc802 = hbusreq1 & v8cc800 | !hbusreq1 & v8cc801;
assign d35a2d = hbusreq1 & d35984 | !hbusreq1 & v845542;
assign v8ccbec = hlock4_p & v8ccbeb | !hlock4_p & v845542;
assign bd590c = hmaster1_p & bd590b | !hmaster1_p & v845542;
assign cc36f9 = hgrant4_p & v84556c | !hgrant4_p & cc36f2;
assign c3cee5 = hbusreq3 & c3cee0 | !hbusreq3 & c3cee4;
assign c3d51d = hmaster0_p & c3d51c | !hmaster0_p & !c3d2be;
assign d35023 = hready_p & d35022 | !hready_p & d35803;
assign v8cc031 = decide_p & v8cc82e | !decide_p & v8cc816;
assign ad45ec = hlock4_p & ad45eb | !hlock4_p & v845542;
assign bd586f = stateG10_4_p & bd5842 | !stateG10_4_p & !bd586e;
assign v8ccbf7 = hmaster0_p & v8ccbe8 | !hmaster0_p & v8ccbf6;
assign v8cc482 = hready & v8cc481 | !hready & v8ccbd8;
assign c3d592 = hbusreq3 & c3d58f | !hbusreq3 & c3d591;
assign v9f7867 = hlock3 & v9f7866 | !hlock3 & v9f7865;
assign c3d5ce = hmaster0_p & c3d5c5 | !hmaster0_p & c3d5cd;
assign d357a0 = hlock0_p & v845542 | !hlock0_p & adea88;
assign b05927 = hmaster1_p & b0591d | !hmaster1_p & b05926;
assign ade573 = hbusreq4_p & ade572 | !hbusreq4_p & !v845542;
assign d354e9 = hgrant2_p & d354e1 | !hgrant2_p & !d354e8;
assign d3574b = hbusreq2 & d3572e | !hbusreq2 & !d35aa4;
assign ad4f1a = hbusreq3 & v845547 | !hbusreq3 & v845542;
assign v9f7875 = hready_p & v9f773a | !hready_p & v9f7874;
assign ad438b = hready & ad437f | !hready & ad438a;
assign ad46f4 = hbusreq1 & ad458b | !hbusreq1 & !v845542;
assign ad4e67 = hbusreq1_p & ad4e64 | !hbusreq1_p & !ad4e66;
assign adec96 = stateA1_p & v845542 | !stateA1_p & adec95;
assign c3d370 = stateA1_p & c3d36f | !stateA1_p & c5c8e4;
assign ad429d = hbusreq1 & ad4d98 | !hbusreq1 & v845542;
assign ad4465 = hbusreq0 & ad4464 | !hbusreq0 & v845542;
assign ad4e65 = hready & v84557a | !hready & v845542;
assign dc53cb = hlock3_p & dc53a6 | !hlock3_p & v845542;
assign c3d755 = decide_p & c3d74c | !decide_p & c3d754;
assign v9f7d27 = hbusreq4 & v9f7d25 | !hbusreq4 & !v9f7d26;
assign bd58ef = hbusreq2 & bd58ee | !hbusreq2 & v845542;
assign c3cf2b = hbusreq3_p & c3cf18 | !hbusreq3_p & c3cf2a;
assign v9e9f5c = hlock1 & v9e9f57 | !hlock1 & v9e9f5b;
assign d359c8 = stateA1_p & v889629 | !stateA1_p & v845542;
assign b1c753 = hburst1 & b1c74f | !hburst1 & b1c752;
assign bd574f = hmaster2_p & bd572e | !hmaster2_p & bd574e;
assign c74620 = hburst1_p & v845542 | !hburst1_p & v857b36;
assign v9ea5d2 = hbusreq1 & v9ea5d0 | !hbusreq1 & v9ea5d1;
assign v9f7754 = hlock4 & v9f7751 | !hlock4 & v9f7753;
assign bd5b7c = hlock3_p & bd5b75 | !hlock3_p & bd5b7b;
assign bd58c3 = hgrant4_p & bd575d | !hgrant4_p & ade563;
assign c3d6c3 = hlock4_p & c3d6c1 | !hlock4_p & c3d6c2;
assign v9ea4dc = hmaster1_p & v9ea4cc | !hmaster1_p & v9ea4db;
assign ad505f = hgrant4_p & v845542 | !hgrant4_p & !ad505e;
assign ad4e8b = hmaster2_p & ad4e8a | !hmaster2_p & v845542;
assign ad41ad = hready_p & ad416f | !hready_p & ad41ac;
assign ad46ce = hlock4_p & ad4f09 | !hlock4_p & ad4f38;
assign v9f7e14 = hbusreq4_p & v9f7e12 | !hbusreq4_p & v9f7e13;
assign b0593a = hmaster2_p & b05939 | !hmaster2_p & !b058a9;
assign ade65b = hmaster0_p & adea95 | !hmaster0_p & ade65a;
assign ad41b5 = hmaster0_p & ad41b4 | !hmaster0_p & ad40f3;
assign df5124 = hbusreq1 & dc5389 | !hbusreq1 & dc538d;
assign df51ae = hmaster0_p & df51a4 | !hmaster0_p & df51ad;
assign b57421 = hlock4 & b57987 | !hlock4 & b57420;
assign ad4ede = hbusreq4_p & ad4edb | !hbusreq4_p & ad4edd;
assign c3d2eb = hgrant4_p & v845542 | !hgrant4_p & c3d2ea;
assign b058ae = hbusreq4 & b058ac | !hbusreq4 & b058ad;
assign d356a3 = hburst0 & d356a2 | !hburst0 & d359bf;
assign d35658 = hbusreq0 & d35650 | !hbusreq0 & d35657;
assign bd584f = hgrant4_p & v845542 | !hgrant4_p & !bd5842;
assign c3ce16 = hmaster0_p & c3ce14 | !hmaster0_p & c3ce15;
assign b57447 = hmaster0_p & b579bb | !hmaster0_p & v845542;
assign v8cc62c = hbusreq3 & v8cc62b | !hbusreq3 & v8ccbd8;
assign v9f7d86 = hlock4_p & v9f7d84 | !hlock4_p & v9f7d85;
assign d35435 = hbusreq4_p & d35434 | !hbusreq4_p & v845542;
assign ad44a4 = hgrant4_p & ad4489 | !hgrant4_p & !c3cec2;
assign c3d480 = hbusreq1 & c3d479 | !hbusreq1 & c3d47c;
assign bd5926 = hbusreq0 & bd5925 | !hbusreq0 & v845564;
assign c3ced3 = hmaster0_p & c3ced2 | !hmaster0_p & c3d306;
assign b059d0 = hlock3 & b059cf | !hlock3 & b059cd;
assign df54f0 = hready_p & v845542 | !hready_p & df54ef;
assign d3578b = hlock0_p & v845542 | !hlock0_p & d3590d;
assign v9f768c = hgrant0_p & v9f7d59 | !hgrant0_p & !v9f768b;
assign d357b7 = hmaster2_p & d3576e | !hmaster2_p & d357b6;
assign b058d3 = hbusreq0_p & v9ea3e9 | !hbusreq0_p & v9f7d42;
assign b058e0 = hbusreq2 & b058de | !hbusreq2 & b058df;
assign v9f7db7 = hlock4 & v9f7db4 | !hlock4 & v9f7db6;
assign b05a3c = hlock2_p & b05a39 | !hlock2_p & b05a3b;
assign b1c734 = hlock0_p & bd576b | !hlock0_p & v845542;
assign c3d4fc = hmaster2_p & adeaa5 | !hmaster2_p & c3d4e1;
assign bd5b91 = hmastlock_p & v8ccb68 | !hmastlock_p & !v845542;
assign b1c720 = hlock0_p & bd574e | !hlock0_p & b1c70e;
assign bd578c = hmaster2_p & bd5786 | !hmaster2_p & !bd578b;
assign b1cf27 = hmaster2_p & v845542 | !hmaster2_p & b1cf26;
assign d357db = hmaster2_p & d357da | !hmaster2_p & v845542;
assign ad4f32 = hbusreq2_p & ad4f25 | !hbusreq2_p & !ad4f31;
assign bd57e8 = hmaster1_p & bd57e7 | !hmaster1_p & bd57b1;
assign v9f7daf = hgrant4_p & v9f7cc7 | !hgrant4_p & v9f7dae;
assign df51df = jx0_p & df51d3 | !jx0_p & df51de;
assign c3ce65 = hbusreq1_p & c3ce64 | !hbusreq1_p & v845542;
assign v8cc7b2 = hgrant1_p & v8cc7b1 | !hgrant1_p & v8ccbe3;
assign b1c726 = hmaster2_p & b1c725 | !hmaster2_p & v845542;
assign d3550d = hbusreq2 & d35421 | !hbusreq2 & d3550c;
assign v9ea5d9 = hmaster0_p & v9ea5d6 | !hmaster0_p & v9ea575;
assign df5163 = hmaster0_p & df5160 | !hmaster0_p & df5162;
assign c3d5ab = hmaster0_p & c3d5aa | !hmaster0_p & !c3d2be;
assign v9f7d6c = hmaster1_p & v9f7d6b | !hmaster1_p & v9f7ce9;
assign dc5064 = hbusreq4 & dc504b | !hbusreq4 & dc5063;
assign ad46f7 = hmaster0_p & ad46af | !hmaster0_p & ad46f6;
assign v9f7d8c = hgrant4_p & v9ea3ec | !hgrant4_p & v9f7d8a;
assign c3ceba = hready_p & v845555 | !hready_p & c3ceb9;
assign ad45b6 = hready & ad45ad | !hready & !ad45b5;
assign v9f7700 = hlock2 & v9f76fd | !hlock2 & v9f76ff;
assign ad4f33 = hbusreq2 & dc4fcc | !hbusreq2 & v845542;
assign b1c74f = hmastlock_p & bd57be | !hmastlock_p & !b1c74e;
assign adeaa1 = hmaster1_p & adea95 | !hmaster1_p & adeaa0;
assign dc4f9d = hburst0 & dc4f9b | !hburst0 & dc4f9c;
assign d355aa = hbusreq3 & d355a3 | !hbusreq3 & d355a9;
assign ad456b = hready & ad4562 | !hready & ad456a;
assign ad448d = hmaster2_p & b1c70e | !hmaster2_p & !ad448c;
assign ad4f6d = hbusreq4_p & ad4f65 | !hbusreq4_p & adeaa4;
assign dc4ffc = hbusreq1 & adec89 | !hbusreq1 & v84556c;
assign v9f7da3 = hmaster2_p & v9f7ca4 | !hmaster2_p & v9f7da2;
assign c3cea6 = hmaster0_p & c3cea5 | !hmaster0_p & !c3d2be;
assign b1c0ab = hbusreq2_p & b1c095 | !hbusreq2_p & b1c0aa;
assign ad473c = hbusreq4 & ad473b | !hbusreq4 & v845564;
assign dc502a = hbusreq4_p & dc5027 | !hbusreq4_p & dc5029;
assign b1c6de = hbusreq2_p & b1c61a | !hbusreq2_p & b1c6dc;
assign c3ce34 = hbusreq1 & c3d2b2 | !hbusreq1 & v845542;
assign v8cc818 = decide_p & v8cc7d7 | !decide_p & v8cc816;
assign ad445c = hlock4_p & ad445b | !hlock4_p & !v845576;
assign b57a80 = hbusreq2 & b57a7e | !hbusreq2 & b57a7f;
assign c3d6fb = hgrant1_p & c3d67b | !hgrant1_p & !c3d6fa;
assign v9f789b = hgrant2_p & v9f7877 | !hgrant2_p & v9f789a;
assign d3573f = hmaster1_p & d3573e | !hmaster1_p & d356fc;
assign b1caee = hbusreq0 & b1caea | !hbusreq0 & b1caed;
assign v8cc038 = jx1_p & v8cc791 | !jx1_p & v8cc036;
assign d3598a = hlock0_p & v845542 | !hlock0_p & d35989;
assign d6ebca = hgrant2_p & v845542 | !hgrant2_p & !v845570;
assign d356c5 = hlock1_p & v84557a | !hlock1_p & v845542;
assign dc501c = hbusreq1_p & dc5018 | !hbusreq1_p & dc501b;
assign ad3ce5 = hready & ad3ce0 | !hready & !ad3ce4;
assign bd575f = hbusreq3 & bd575e | !hbusreq3 & df513c;
assign ad4e77 = hgrant4_p & v84557a | !hgrant4_p & !ad4e75;
assign ad4d99 = hbusreq3 & ad4d98 | !hbusreq3 & v845542;
assign v9f7e02 = hmaster0_p & v9f7d10 | !hmaster0_p & v9f7e01;
assign c3ce43 = hbusreq1 & c3d314 | !hbusreq1 & c3d305;
assign ad425a = hgrant2_p & v845542 | !hgrant2_p & ad4259;
assign ade556 = hgrant0_p & v845542 | !hgrant0_p & !ade550;
assign ad40ea = hbusreq2_p & ad40e9 | !hbusreq2_p & v845542;
assign b1c749 = hmaster1_p & b1c748 | !hmaster1_p & b1c745;
assign c5c8e0 = hbusreq2_p & c5c8a8 | !hbusreq2_p & c5c8a7;
assign ade5da = hmaster1_p & ade5d2 | !hmaster1_p & ade5d9;
assign d35a0c = hlock4_p & d359f0 | !hlock4_p & !d35a0b;
assign d3576a = hbusreq3_p & d35762 | !hbusreq3_p & !d35769;
assign b0595b = hmaster2_p & b05952 | !hmaster2_p & v9ea3e9;
assign b05a85 = hmaster0_p & b059a9 | !hmaster0_p & b059bd;
assign ad4ec9 = hbusreq3 & ad4ec8 | !hbusreq3 & v845542;
assign v9ea56a = hmaster2_p & v9ea4ab | !hmaster2_p & v9ea569;
assign v8cc5fe = hmaster1_p & v8cc5fd | !hmaster1_p & v845542;
assign c3d5a0 = hready & c3d59f | !hready & !v845542;
assign b5795b = hlock2_p & b57959 | !hlock2_p & b5795a;
assign d3558a = hbusreq1_p & d354c9 | !hbusreq1_p & !d35589;
assign v9ea443 = stateG10_4_p & v9ea441 | !stateG10_4_p & v9ea442;
assign v9e9f60 = hlock3 & v9e9f5f | !hlock3 & v9e9f5e;
assign df5531 = hready_p & v845542 | !hready_p & df5530;
assign v9f7860 = hbusreq0 & v9f7759 | !hbusreq0 & v9f785f;
assign bd582a = hmaster2_p & bd580a | !hmaster2_p & v845542;
assign c5c903 = hgrant2_p & c5c8f0 | !hgrant2_p & c5c902;
assign ad45a6 = hmaster1_p & ad459f | !hmaster1_p & ad45a5;
assign c5c8a4 = hbusreq2_p & c5c8a3 | !hbusreq2_p & c5c8a2;
assign b059ad = hbusreq2_p & b059a6 | !hbusreq2_p & b059ac;
assign b578f9 = hmastlock_p & b578f8 | !hmastlock_p & v845542;
assign c3d4f6 = hbusreq4 & c3d4f5 | !hbusreq4 & !c3d304;
assign v9ea4b9 = hbusreq4_p & v9ea3fb | !hbusreq4_p & v9ea4b6;
assign bd57de = hbusreq1_p & dc4fb0 | !hbusreq1_p & dc4fbe;
assign v9ea4d9 = hmaster2_p & v9ea4d2 | !hmaster2_p & v9ea4d8;
assign af7f59 = hburst1_p & c74202 | !hburst1_p & v845542;
assign ad5042 = hgrant4_p & v84556c | !hgrant4_p & ad5041;
assign v9f7810 = hgrant1_p & v9f7735 | !hgrant1_p & !v9f780f;
assign b1c5e4 = hgrant0_p & d35a58 | !hgrant0_p & !v845542;
assign ad45f8 = hmaster0_p & ad45cc | !hmaster0_p & ad45f4;
assign c3ceb0 = hbusreq1_p & v845564 | !hbusreq1_p & c3ceaf;
assign df54e4 = hlock1_p & df54e3 | !hlock1_p & v845542;
assign v9f7740 = decide_p & v9f773f | !decide_p & v9f773a;
assign b05909 = hbusreq0 & v9f7d42 | !hbusreq0 & b05908;
assign d35bff = hbusreq2_p & d35bfb | !hbusreq2_p & d35bfe;
assign ad4457 = hlock4_p & ad4456 | !hlock4_p & v845542;
assign v9f7d5f = hbusreq1_p & v9f7d5b | !hbusreq1_p & v9f7d5e;
assign c3ceb5 = hbusreq1_p & c3ce8f | !hbusreq1_p & c3ceb4;
assign d35a55 = hbusreq3 & d35a54 | !hbusreq3 & v845542;
assign ad5048 = locked_p & ad5047 | !locked_p & !v845542;
assign v9f7825 = hgrant1_p & v9f7797 | !hgrant1_p & v9f7824;
assign c3d2f3 = hmaster2_p & c3d2f2 | !hmaster2_p & adeaa5;
assign d35a46 = hlock4_p & d35a44 | !hlock4_p & !d35a45;
assign b57a8d = decide_p & b57940 | !decide_p & b57a8c;
assign c3d320 = stateG10_4_p & ade562 | !stateG10_4_p & c3d30d;
assign b059a5 = hgrant2_p & b059a4 | !hgrant2_p & b059a1;
assign dc538f = hmaster0_p & dc538e | !hmaster0_p & v84556c;
assign b1c56a = hmaster0_p & b1c85a | !hmaster0_p & b1c569;
assign ad4742 = hbusreq4_p & ad4741 | !hbusreq4_p & v845542;
assign d3551a = hmaster0_p & d35515 | !hmaster0_p & d35519;
assign b05a41 = hbusreq1_p & b05920 | !hbusreq1_p & b05a40;
assign ad4f7e = hgrant4_p & ad4f39 | !hgrant4_p & ad4e98;
assign c3d5b4 = stateG10_4_p & c3d5b2 | !stateG10_4_p & c3d5b3;
assign ade593 = hbusreq4_p & ade592 | !hbusreq4_p & !v845542;
assign ad42ea = hbusreq1 & ad4ea7 | !hbusreq1 & v845542;
assign adeaa7 = hgrant2_p & v845542 | !hgrant2_p & adeaa6;
assign v9f7d98 = hgrant1_p & v9f7d6e | !hgrant1_p & v9f7d97;
assign c3d2d5 = hlock3_p & c3d2c0 | !hlock3_p & c3d2d2;
assign v9e9fc3 = hmaster1_p & v9e9fc2 | !hmaster1_p & v9e9f9f;
assign ad4db1 = hbusreq0 & ad4dae | !hbusreq0 & ad4db0;
assign v9f7854 = hready_p & v9f7817 | !hready_p & v9f7853;
assign c3d4f2 = hbusreq0 & c3d4f1 | !hbusreq0 & v845542;
assign b1c50c = hbusreq2_p & b1c4af | !hbusreq2_p & b1c4d0;
assign df54d9 = hbusreq1_p & df54d8 | !hbusreq1_p & v845542;
assign c5c8fc = hgrant0_p & c5c88e | !hgrant0_p & !v845542;
assign b57949 = hgrant4_p & v845542 | !hgrant4_p & b5b409;
assign ad428c = hmaster0_p & ad4283 | !hmaster0_p & ad428b;
assign b059f7 = hgrant2_p & b0594b | !hgrant2_p & b059f6;
assign ad4428 = hbusreq1_p & ad4427 | !hbusreq1_p & ad40fe;
assign bd5baa = hmaster0_p & v84556c | !hmaster0_p & bd5ba9;
assign c3d599 = hmaster0_p & c3d598 | !hmaster0_p & c3d2be;
assign b57ac5 = hbusreq1 & b57ac3 | !hbusreq1 & b57ac4;
assign ad4468 = hgrant1_p & ad4440 | !hgrant1_p & ad4467;
assign c3d34c = hmaster2_p & c3d343 | !hmaster2_p & c3d2fd;
assign v9e9ed7 = hready_p & v9ea436 | !hready_p & v9e9ed6;
assign d35a4d = hmastlock_p & v8cc792 | !hmastlock_p & !v845542;
assign ade615 = hbusreq2 & ade4a6 | !hbusreq2 & adec93;
assign c3cedf = hbusreq0 & c3cede | !hbusreq0 & !v845542;
assign v9f776f = hlock3 & v9f7751 | !hlock3 & v9f7757;
assign v9f7896 = hbusreq3 & v9f7894 | !hbusreq3 & v9f7895;
assign ade4de = hburst1 & c3d66d | !hburst1 & ade4c3;
assign v8cc7c5 = hready & v8cc7c4 | !hready & v8ccbf4;
assign b05a28 = hgrant2_p & b05a24 | !hgrant2_p & b05a27;
assign ad4f14 = hgrant1_p & ad4ed1 | !hgrant1_p & ad4f13;
assign v9ea4c3 = hready_p & v9ea4a4 | !hready_p & v9ea4c2;
assign v9f7cad = hlock1 & v9f7ca7 | !hlock1 & v9f7cac;
assign ade4e8 = hlock0_p & ade4cc | !hlock0_p & ade4e7;
assign b05a51 = hgrant2_p & b05a4e | !hgrant2_p & b05a50;
assign c76645 = stateG3_0_p & v845580 | !stateG3_0_p & v845542;
assign c3d733 = hmaster1_p & c3d732 | !hmaster1_p & c3d67c;
assign d3559c = hmaster0_p & d35597 | !hmaster0_p & d3559b;
assign ad4dbd = hbusreq2 & ad4da1 | !hbusreq2 & ad4dbc;
assign ade4da = hbusreq4_p & ade4d9 | !hbusreq4_p & !v845542;
assign v9f7d1f = hbusreq2 & v9f7d1d | !hbusreq2 & v9f7d1e;
assign c3d4e3 = hbusreq0 & c3d4dd | !hbusreq0 & c3d4e2;
assign v9f7763 = hbusreq1_p & v9f7762 | !hbusreq1_p & v9f775a;
assign adeaa0 = hmaster0_p & adea95 | !hmaster0_p & adea9f;
assign ad5025 = hbusreq3 & ad5022 | !hbusreq3 & ad5024;
assign c3d5c9 = hbusreq0 & c3d5be | !hbusreq0 & c3d5c8;
assign c3d6bc = hbusreq4_p & c3d6b9 | !hbusreq4_p & c3d6bb;
assign bd5b77 = hbusreq2 & dc5394 | !hbusreq2 & df54d6;
assign v9f7d3a = hmastlock_p & b06735 | !hmastlock_p & v845542;
assign b05988 = hgrant4_p & b058e9 | !hgrant4_p & v9ea3e9;
assign b1cf2f = hmaster1_p & v845542 | !hmaster1_p & b1cf2e;
assign d357cf = hbusreq1 & d35771 | !hbusreq1 & d35776;
assign bd5b89 = hmaster2_p & v84556c | !hmaster2_p & bd5b88;
assign bd5744 = locked_p & bd5740 | !locked_p & v845542;
assign v9ea44a = hgrant1_p & v9ea3fc | !hgrant1_p & v9ea449;
assign bd5789 = hmastlock_p & bd5788 | !hmastlock_p & v845542;
assign c3d66a = locked_p & v845542 | !locked_p & !c3d669;
assign v8cc7cc = hbusreq3 & v8cc7ca | !hbusreq3 & v8cc7cb;
assign b57a0f = decide_p & b57940 | !decide_p & b57a0e;
assign v9f77b8 = hbusreq2_p & v9f77b1 | !hbusreq2_p & v9f77b7;
assign b1c785 = hmaster0_p & b1c77f | !hmaster0_p & b1c77b;
assign v9ea608 = hlock3 & v9ea607 | !hlock3 & v9ea606;
assign v9f77e5 = hlock2 & v9f77e2 | !hlock2 & v9f77e4;
assign d354c9 = hlock1_p & d354c7 | !hlock1_p & d354c8;
assign dc53a4 = hbusreq3 & dc53a3 | !hbusreq3 & v845564;
assign b1c6cb = hgrant2_p & v845542 | !hgrant2_p & b1c6ca;
assign c3d697 = hmaster2_p & c3d669 | !hmaster2_p & !c3d670;
assign c3ce60 = hbusreq1_p & c3ce5f | !hbusreq1_p & v845564;
assign ad46dc = hgrant4_p & v845542 | !hgrant4_p & ad46db;
assign v9ea402 = hbusreq0_p & v9ea3fb | !hbusreq0_p & v9ea3fe;
assign v9e9fb5 = hgrant3_p & v9e9ef7 | !hgrant3_p & v9e9fb4;
assign d3591a = hlock0_p & dc5318 | !hlock0_p & v845542;
assign d35570 = hbusreq2 & d354f9 | !hbusreq2 & !d354f5;
assign ad42cd = hlock2_p & ad42ca | !hlock2_p & ad42cc;
assign v9ea5bd = hmaster1_p & v9ea5bc | !hmaster1_p & v9ea56b;
assign d35743 = hbusreq2 & d356cb | !hbusreq2 & !v84554e;
assign ad4782 = hmaster1_p & ad476d | !hmaster1_p & ad4781;
assign v9f7662 = hbusreq0_p & v9f7ddd | !hbusreq0_p & v9f7661;
assign d356bd = hmaster0_p & d356a9 | !hmaster0_p & d356bc;
assign ad4391 = hmaster0_p & ad438c | !hmaster0_p & ad4390;
assign b574b5 = hlock4 & b57942 | !hlock4 & b574b4;
assign bd57d1 = hbusreq1_p & bd57cf | !hbusreq1_p & bd57d0;
assign v9f7ce4 = hbusreq1 & v9f7ce2 | !hbusreq1 & v9f7ce3;
assign b579e5 = hgrant1_p & v845542 | !hgrant1_p & b579ce;
assign b0598f = hgrant4_p & b058d4 | !hgrant4_p & !b0598e;
assign b05a99 = hready_p & b05a8d | !hready_p & !b05a98;
assign v9f7dfd = hlock2_p & v9f7df9 | !hlock2_p & v9f7dfc;
assign ad4334 = hgrant1_p & ad432e | !hgrant1_p & ad4333;
assign c3d69b = hmaster0_p & c3d69a | !hmaster0_p & !c3d67b;
assign ad508f = decide_p & v845542 | !decide_p & ad508e;
assign ad437f = hbusreq0 & ad437e | !hbusreq0 & v845542;
assign ad4f5a = hmaster0_p & ad4f54 | !hmaster0_p & ad4f59;
assign d3570a = hgrant1_p & v845542 | !hgrant1_p & d35709;
assign b8f746 = jx1_p & b8f745 | !jx1_p & b8f6e7;
assign d35a9b = hbusreq4_p & v84555a | !hbusreq4_p & !v845542;
assign ad449a = hgrant1_p & ad4490 | !hgrant1_p & ad4499;
assign b57af1 = hbusreq3 & b57af0 | !hbusreq3 & b57942;
assign ad4374 = hgrant2_p & ad4372 | !hgrant2_p & ad4373;
assign v8cc435 = hgrant1_p & v8ccb6b | !hgrant1_p & v8ccbe3;
assign bd5771 = hmaster2_p & c3d669 | !hmaster2_p & v845542;
assign v8cc0e1 = hgrant1_p & v845542 | !hgrant1_p & v8cc0e0;
assign b1c05e = hmaster1_p & b1c05a | !hmaster1_p & b1c05d;
assign v8cc792 = stateA1_p & v8ccb68 | !stateA1_p & v8ccb67;
assign v8cc436 = stateG10_4_p & v845542 | !stateG10_4_p & v8ccbeb;
assign v8cc494 = hmaster2_p & v8cc491 | !hmaster2_p & v8cc493;
assign ade5b5 = hmaster0_p & ade569 | !hmaster0_p & ade5b4;
assign dc4fee = hgrant4_p & v84556c | !hgrant4_p & ade553;
assign v9f778b = hlock1 & v9f772c | !hlock1 & v9f778a;
assign ad4733 = hgrant1_p & ad460b | !hgrant1_p & ad4732;
assign dc4fd8 = hbusreq4_p & adec89 | !hbusreq4_p & adeca1;
assign v9f780f = hmaster2_p & v9f7809 | !hmaster2_p & !v9f780e;
assign b1c585 = hbusreq2_p & b1cafe | !hbusreq2_p & b1c584;
assign c3d5d9 = hgrant0_p & v845542 | !hgrant0_p & c3d5d3;
assign v9f76d6 = hmaster1_p & v9f76d5 | !hmaster1_p & v9f7df7;
assign ad5090 = hready_p & v845542 | !hready_p & ad508f;
assign c3d2bf = hmaster0_p & c3d2bb | !hmaster0_p & c3d2be;
assign d3579e = hmaster2_p & d3579d | !hmaster2_p & v845542;
assign c3ce28 = hready_p & v845555 | !hready_p & c3ce27;
assign b1c568 = hbusreq1_p & b1cc00 | !hbusreq1_p & b1c567;
assign ba05cd = hbusreq2_p & v845542 | !hbusreq2_p & v845572;
assign v9ea4ca = hmaster2_p & v9ea444 | !hmaster2_p & v9ea4c9;
assign d35914 = hbusreq1 & d3590e | !hbusreq1 & d35910;
assign c3cec5 = hbusreq4_p & v8da59f | !hbusreq4_p & !c3cec4;
assign ad445f = hbusreq0 & ad445e | !hbusreq0 & v845542;
assign v9f7cb3 = hmastlock_p & v9f7c95 | !hmastlock_p & v845542;
assign b059af = stateG10_4_p & b05953 | !stateG10_4_p & b059ae;
assign c3ce74 = hgrant3_p & c3ce42 | !hgrant3_p & c3ce73;
assign v9ea576 = hbusreq1_p & v9ea572 | !hbusreq1_p & v9ea575;
assign bd58f6 = hbusreq1 & bd574f | !hbusreq1 & v84556c;
assign ad3d1f = decide_p & ad440a | !decide_p & ad3d1e;
assign b05935 = hlock3_p & b0592d | !hlock3_p & b05934;
assign b579ce = hmaster2_p & b579cb | !hmaster2_p & b579cd;
assign b1c7eb = hmaster0_p & b1c7e9 | !hmaster0_p & b1c7ea;
assign dc506e = hbusreq2 & dc506c | !hbusreq2 & !dc506d;
assign bd5877 = hgrant4_p & c3d689 | !hgrant4_p & bd5875;
assign ad4f9e = hmaster0_p & ad4f61 | !hmaster0_p & ad4f9d;
assign d3594f = hmaster2_p & d35909 | !hmaster2_p & !d3594e;
assign ad4753 = hgrant2_p & ad4752 | !hgrant2_p & ad474f;
assign ade4e9 = hbusreq4_p & ade4e8 | !hbusreq4_p & !v845542;
assign b058e9 = locked_p & v9fa31b | !locked_p & v9ea3e9;
assign b05974 = hlock2 & b05971 | !hlock2 & b05973;
assign b1c045 = hbusreq0 & b1c044 | !hbusreq0 & b1c847;
assign v9e9f51 = stateG10_4_p & v9e9f4f | !stateG10_4_p & v9e9f50;
assign b1c55f = hbusreq4_p & b1cbf3 | !hbusreq4_p & !b1c85d;
assign v9f77fa = hgrant1_p & v9f7730 | !hgrant1_p & v9f77d8;
assign jx1 = !b05a9e;
assign v9f76c4 = hlock0_p & v9f7d3a | !hlock0_p & v9f76c3;
assign v9ea4cb = hgrant1_p & v9ea4b7 | !hgrant1_p & v9ea4ca;
assign v8ccbdc = hready_p & v8ccb74 | !hready_p & v8ccbdb;
assign d35697 = hbusreq2_p & d35692 | !hbusreq2_p & !d35696;
assign ad4df3 = hmaster1_p & ad4de6 | !hmaster1_p & ad4df2;
assign cc36ee = hgrant3_p & cc36c3 | !hgrant3_p & cc36ed;
assign d357e7 = hready_p & d357e4 | !hready_p & d357b2;
assign b05904 = hlock3 & b058c9 | !hlock3 & b05903;
assign b5794a = hmaster2_p & b57949 | !hmaster2_p & v845542;
assign b058b2 = hlock3 & b058aa | !hlock3 & b058b1;
assign ad46ee = hgrant2_p & ad46ed | !hgrant2_p & !ad46e5;
assign ad4588 = hbusreq3 & ad4586 | !hbusreq3 & !v845542;
assign bd5852 = hmaster2_p & bd581c | !hmaster2_p & bd5851;
assign v8cc0de = hready & v8cc0dd | !hready & v8cc494;
assign ad4333 = hbusreq1_p & ad4332 | !hbusreq1_p & ad5023;
assign v9e9e79 = hbusreq1_p & v9ea3ff | !hbusreq1_p & v9ea4b7;
assign v9f7784 = hlock3_p & v9f777c | !hlock3_p & v9f7783;
assign ad4f61 = hbusreq3 & ad4f60 | !hbusreq3 & v845542;
assign c3d6ea = hbusreq1_p & c3d66f | !hbusreq1_p & c3d6e9;
assign bd57f2 = hbusreq1 & c3d683 | !hbusreq1 & !v845542;
assign b8ef51 = jx1_p & b8ef50 | !jx1_p & b8f745;
assign df51bc = hmaster1_p & df51bb | !hmaster1_p & df5178;
assign v9f779f = hmaster2_p & v9f772b | !hmaster2_p & !v9f779d;
assign v9f7da0 = hlock1_p & v9f7cae | !hlock1_p & v9f7cff;
assign stateG10_3 = !bcd5a7;
assign c5c8a8 = hlock2_p & c5c8a6 | !hlock2_p & c5c8a7;
assign c3d6f2 = hgrant4_p & c3d674 | !hgrant4_p & c3d6b7;
assign c5c9b1 = hgrant2_p & c5c9b0 | !hgrant2_p & c5c978;
assign v9ea472 = stateG10_4_p & v9ea470 | !stateG10_4_p & v9ea471;
assign ade566 = hbusreq4_p & ade565 | !hbusreq4_p & !v845542;
assign ad473b = hmaster2_p & v845542 | !hmaster2_p & ad473a;
assign ad3d24 = hmaster0_p & ad448f | !hmaster0_p & ad43aa;
assign ad430a = hlock1_p & ad4308 | !hlock1_p & ad4309;
assign ad4159 = hbusreq4_p & ad4f94 | !hbusreq4_p & v845542;
assign df513f = hbusreq3 & df5139 | !hbusreq3 & df513e;
assign ad475d = hbusreq2_p & ad475a | !hbusreq2_p & ad475c;
assign df5536 = hmaster1_p & df5532 | !hmaster1_p & df5535;
assign b05a4a = hbusreq2_p & b05a47 | !hbusreq2_p & b05a49;
assign cc36e1 = hgrant4_p & v845566 | !hgrant4_p & !cc36da;
assign b1c844 = hbusreq4_p & b1cf29 | !hbusreq4_p & b1c843;
assign ad3d30 = hbusreq2_p & ad3d2d | !hbusreq2_p & ad3d2f;
assign ad46a3 = hmaster2_p & ad46a2 | !hmaster2_p & v845542;
assign b05943 = hmaster0_p & b0593e | !hmaster0_p & !b05942;
assign ad48c8 = decide_p & v845542 | !decide_p & ad48c7;
assign ad4ff3 = hmaster1_p & ad4ff2 | !hmaster1_p & ad4fb8;
assign v9f76ab = hgrant1_p & v9f7d5e | !hgrant1_p & v9f7698;
assign d359a5 = hgrant4_p & v845542 | !hgrant4_p & d35997;
assign d355a1 = hgrant3_p & d3552f | !hgrant3_p & !d355a0;
assign ad46a4 = hmastlock_p & ade54c | !hmastlock_p & !v845542;
assign dc4fe1 = hbusreq1 & dc4fe0 | !hbusreq1 & !v845542;
assign ad43fb = hready & ad43f2 | !hready & ad43fa;
assign ad4813 = hmaster1_p & ad480f | !hmaster1_p & ad4812;
assign c3d5d0 = hmaster0_p & c3d5c5 | !hmaster0_p & c3d5cf;
assign df51d2 = hbusreq3_p & df51d1 | !hbusreq3_p & df5543;
assign ad441a = hmaster1_p & ad4412 | !hmaster1_p & ad4419;
assign ad45cc = hbusreq1_p & ad45cb | !hbusreq1_p & ad45ca;
assign ade543 = hbusreq2 & ade4a7 | !hbusreq2 & adec93;
assign ad42dc = hready_p & ad429c | !hready_p & ad42db;
assign v8cc48a = hbusreq3 & v8cc488 | !hbusreq3 & v8cc489;
assign c3ce5c = decide_p & c3ce50 | !decide_p & c3ce5b;
assign d35013 = hbusreq0 & d35012 | !hbusreq0 & d35aac;
assign v9f7d67 = hmaster1_p & v9f7d66 | !hmaster1_p & v9f7d64;
assign ad470e = hbusreq1_p & ad459d | !hbusreq1_p & ad470d;
assign df51d3 = jx1_p & df51ce | !jx1_p & df51d2;
assign ba7c69 = decide_p & ba7c68 | !decide_p & v845558;
assign bd56dd = hlock2_p & bd56dc | !hlock2_p & v845542;
assign df5145 = hbusreq1 & dc4fc9 | !hbusreq1 & v845542;
assign v9f775f = hlock1 & v9f775a | !hlock1 & v9f775e;
assign ad40fa = hbusreq2_p & ad40f8 | !hbusreq2_p & ad508e;
assign adea8d = hmaster1_p & v845542 | !hmaster1_p & adea8c;
assign ad4f41 = hbusreq3 & ad4f40 | !hbusreq3 & v845542;
assign d3599c = hbusreq4_p & d3599a | !hbusreq4_p & d3599b;
assign b57433 = hmaster1_p & b57432 | !hmaster1_p & v845542;
assign b1c087 = hbusreq4 & b1c081 | !hbusreq4 & b1c086;
assign ad4ed8 = hgrant0_p & ad4eae | !hgrant0_p & v845542;
assign d358fe = hbusreq3 & d358fd | !hbusreq3 & v845542;
assign ad48b1 = hready & ad4de1 | !hready & ad48b0;
assign c3d31c = hmaster2_p & v845542 | !hmaster2_p & c3d31b;
assign c5c9a8 = hmaster0_p & c5c974 | !hmaster0_p & c5c8e9;
assign d356b1 = hbusreq1_p & d356b0 | !hbusreq1_p & v845542;
assign d354f8 = hmaster2_p & d354f1 | !hmaster2_p & !d354f7;
assign c3d32b = hready & c3d324 | !hready & c3d32a;
assign b1c771 = hbusreq4_p & b1c770 | !hbusreq4_p & !ade4d9;
assign v9ea4e5 = hgrant3_p & v9ea4c3 | !hgrant3_p & v9ea4e4;
assign ad43c3 = stateA1_p & v845542 | !stateA1_p & ad43c2;
assign c3d5e9 = hmaster2_p & v8da59f | !hmaster2_p & v845576;
assign ad4e51 = hmaster0_p & ad4e44 | !hmaster0_p & ad4e50;
assign dc4ff7 = hmaster2_p & dc4ff6 | !hmaster2_p & v845542;
assign v9f7d69 = decide_p & v9f7d56 | !decide_p & !v9f7d68;
assign v9ea3fa = hmaster2_p & v9ea3e6 | !hmaster2_p & v9f20a1;
assign c3d2dc = hmaster0_p & c3d2d7 | !hmaster0_p & c3d2db;
assign ad4826 = hmaster1_p & ad4822 | !hmaster1_p & ad4825;
assign ad3cd7 = hbusreq0 & v845542 | !hbusreq0 & c3d327;
assign ade4cc = hburst0 & ade4c8 | !hburst0 & ade4cb;
assign v8ccbdb = decide_p & v8ccbd7 | !decide_p & v8ccbda;
assign dc5054 = hbusreq4_p & dc5051 | !hbusreq4_p & dc5053;
assign bd5865 = hlock0_p & bd5861 | !hlock0_p & bd5864;
assign ade4b8 = stateG2_p & v845542 | !stateG2_p & ade4b7;
assign c3d2ae = hmastlock_p & c3d2ad | !hmastlock_p & !v845542;
assign v9e9fba = hmaster1_p & v9e9fb9 | !hmaster1_p & v9e9ef1;
assign ad42a1 = hbusreq1_p & ad42a0 | !hbusreq1_p & v845542;
assign v9e9e9d = stateG10_4_p & v9e9e9b | !stateG10_4_p & v9e9e9c;
assign v9e9edb = hbusreq2_p & v9e9eda | !hbusreq2_p & v9ea5f7;
assign ad40f5 = hbusreq2 & ad501b | !hbusreq2 & v845547;
assign v9f7ccd = hready & v9f7ccc | !hready & v9f7cc8;
assign ad4eca = hbusreq1 & ad4e5e | !hbusreq1 & v845542;
assign v9ea58c = hready & v9ea58b | !hready & v9ea586;
assign adea85 = hburst0_p & c74a04 | !hburst0_p & !v8f2540;
assign b1c85f = hbusreq0 & b1c858 | !hbusreq0 & b1c85e;
assign ad4f81 = hgrant4_p & v84556c | !hgrant4_p & ad4f80;
assign d35906 = stateA1_p & ade4b9 | !stateA1_p & !d35905;
assign cc36c5 = hlock1_p & v84556c | !hlock1_p & !cc36b8;
assign bd5ba5 = hlock2_p & bd5ba4 | !hlock2_p & v845542;
assign v9f7d7d = stateG10_4_p & v9f7d79 | !stateG10_4_p & !v9f7d7b;
assign d3563d = hgrant0_p & v84556c | !hgrant0_p & !d3563c;
assign v9f7842 = stateG10_4_p & v9f780b | !stateG10_4_p & !v9f7841;
assign b1c746 = hmaster1_p & b1c73b | !hmaster1_p & b1c745;
assign ad4d9c = hready & ad4d96 | !hready & !ad4d9b;
assign ad4895 = hgrant1_p & ad4894 | !hgrant1_p & ad4db7;
assign b57a1b = hbusreq4_p & b578f9 | !hbusreq4_p & b57a1a;
assign c3cf1b = hbusreq1_p & c3cee0 | !hbusreq1_p & c3cf1a;
assign ad4398 = hbusreq0 & ad4397 | !hbusreq0 & v845542;
assign ad4844 = hmaster2_p & v845542 | !hmaster2_p & d35616;
assign b1c7de = hbusreq4_p & b1c7db | !hbusreq4_p & !b1c7dd;
assign ad4282 = hlock1_p & ad40fe | !hlock1_p & !v845542;
assign dc504b = hbusreq0 & dc5041 | !hbusreq0 & dc504a;
assign c3d5e2 = hmaster2_p & c3d5e1 | !hmaster2_p & c3d2fd;
assign v8ccbe5 = hgrant1_p & v845542 | !hgrant1_p & v8ccbe3;
assign v9f782f = hmaster2_p & v9f77c7 | !hmaster2_p & !v9f782d;
assign d354f1 = hbusreq4_p & d35c00 | !hbusreq4_p & v845542;
assign v8cc16c = jx1_p & v8cc132 | !jx1_p & v8cc16a;
assign ad4848 = hbusreq1_p & ad4845 | !hbusreq1_p & ad4847;
assign v8ccb8d = hmaster1_p & v8ccb75 | !hmaster1_p & v8ccb81;
assign v9f7d02 = hlock2 & v9f7cf8 | !hlock2 & v9f7d01;
assign d359c1 = locked_p & d359c0 | !locked_p & !v845542;
assign b1c5d7 = hmaster2_p & v845542 | !hmaster2_p & !d3590d;
assign dc5013 = hbusreq0 & dc500d | !hbusreq0 & dc5012;
assign c3d325 = hmaster2_p & adeaa5 | !hmaster2_p & v845576;
assign b1c078 = hbusreq1_p & b1c7b2 | !hbusreq1_p & b1c077;
assign d35a73 = hmaster2_p & d35a47 | !hmaster2_p & v845542;
assign d35733 = hmaster1_p & d3572d | !hmaster1_p & d35732;
assign ad43f8 = hmaster2_p & ad43f7 | !hmaster2_p & !v845542;
assign d35629 = hbusreq0 & d35919 | !hbusreq0 & d35628;
assign bd5891 = stateG10_4_p & bd5875 | !stateG10_4_p & !bd5890;
assign b574d5 = hlock2 & b57942 | !hlock2 & b574d4;
assign b1c7a5 = hgrant4_p & v845542 | !hgrant4_p & b1c797;
assign b1c062 = hlock0_p & b1c795 | !hlock0_p & b1c061;
assign v9f76f6 = hbusreq4 & v9f76f4 | !hbusreq4 & v9f76f5;
assign ade5ca = hburst0_p & c74a04 | !hburst0_p & !v857b36;
assign b1c06f = hgrant4_p & v845542 | !hgrant4_p & b1c066;
assign b0596d = hgrant1_p & b0596a | !hgrant1_p & b0596c;
assign v9ea607 = hgrant1_p & v9ea43b | !hgrant1_p & v9ea45c;
assign b1c5df = hready_p & v845542 | !hready_p & b1c5de;
assign v8cc126 = hlock2 & v8ccbd8 | !hlock2 & v8cc125;
assign v9e9f9b = hlock3 & v9e9f9a | !hlock3 & v9e9f99;
assign ad3d39 = hgrant2_p & ad446d | !hgrant2_p & ad3d37;
assign b1cf2a = hmaster2_p & v845542 | !hmaster2_p & !b1cf29;
assign b1c710 = hbusreq0_p & bd575d | !hbusreq0_p & v845542;
assign d3561a = hburst0_p & c74a04 | !hburst0_p & !d35619;
assign ad443d = hbusreq1_p & ad4432 | !hbusreq1_p & ad443c;
assign bd5bab = hmaster1_p & bd5baa | !hmaster1_p & v84556c;
assign b57908 = hmaster1_p & b57907 | !hmaster1_p & b57901;
assign v9f7dfc = hgrant2_p & v9f7dfb | !hgrant2_p & v9f7df8;
assign d35a17 = hbusreq0 & d35a11 | !hbusreq0 & d35a16;
assign bd56ce = stateA1_p & c74a04 | !stateA1_p & ade4b7;
assign ad4713 = hmaster2_p & v845542 | !hmaster2_p & ad4712;
assign ad13e1 = hready_p & v84554c | !hready_p & ad13e0;
assign ad46c8 = hbusreq4_p & ad46c7 | !hbusreq4_p & v845542;
assign v9f76b3 = hmaster0_p & v9f7e01 | !hmaster0_p & v9f7d10;
assign b0599a = hgrant1_p & b05977 | !hgrant1_p & !b05999;
assign d35577 = hbusreq1 & d354f8 | !hbusreq1 & !d35a9b;
assign d35bf2 = hmaster2_p & d35be3 | !hmaster2_p & d35bf1;
assign bd5780 = decide_p & bd577f | !decide_p & v845542;
assign dc4f89 = hmaster2_p & ade4bf | !hmaster2_p & !ade5ce;
assign adeca0 = hmastlock_p & v889629 | !hmastlock_p & v845542;
assign d35aa0 = hmaster1_p & d35a9a | !hmaster1_p & d35a9f;
assign b1c070 = stateG10_4_p & b1c066 | !stateG10_4_p & b1c06f;
assign c3ceab = hgrant3_p & c3ce97 | !hgrant3_p & c3ceaa;
assign bd5ea6 = hgrant2_p & bd5ea5 | !hgrant2_p & !v845542;
assign v9f76ef = hgrant4_p & v9f7ca4 | !hgrant4_p & v9f76ee;
assign ad4ebf = hgrant4_p & v845542 | !hgrant4_p & ad4eb3;
assign v9f7d80 = locked_p & v9f7d3a | !locked_p & !v9f7ca4;
assign v9f7849 = hgrant1_p & v9f77a5 | !hgrant1_p & v9f7835;
assign v9ea5e1 = hmaster1_p & v9ea5e0 | !hmaster1_p & v9ea5aa;
assign d35805 = hbusreq1_p & d357bf | !hbusreq1_p & d357e9;
assign ad42b8 = hbusreq4 & ad42b3 | !hbusreq4 & ad42b7;
assign df519c = hmaster0_p & df517c | !hmaster0_p & df519b;
assign bd5894 = hbusreq0 & bd5888 | !hbusreq0 & bd5893;
assign ad4690 = hbusreq1_p & ad468e | !hbusreq1_p & !ad468f;
assign ad3d01 = stateG10_4_p & ad3ceb | !stateG10_4_p & !ad3d00;
assign ad42ab = hbusreq1_p & ad42aa | !hbusreq1_p & v845542;
assign d354a5 = hlock4_p & v845542 | !hlock4_p & !dc500f;
assign b1c094 = hmaster1_p & b1cfb8 | !hmaster1_p & b1c093;
assign ad45ca = hbusreq1 & ad45c6 | !hbusreq1 & ad45c9;
assign b058df = hlock2 & b058d5 | !hlock2 & b058de;
assign dc505a = hgrant4_p & dc5050 | !hgrant4_p & ade563;
assign ad4eae = locked_p & d359c8 | !locked_p & ad4e53;
assign ad43aa = hbusreq0 & b1c70e | !hbusreq0 & v845542;
assign b1c4a5 = hmaster2_p & v845542 | !hmaster2_p & b1c4a4;
assign cc36e4 = hgrant4_p & cc36bd | !hgrant4_p & !v845566;
assign v9e9fe2 = hbusreq2_p & v9e9fdf | !hbusreq2_p & v9e9fe1;
assign v9f7dd3 = hlock4_p & v9f7dd1 | !hlock4_p & !v9f7dd2;
assign v9f77b1 = hmaster1_p & v9f779c | !hmaster1_p & v9f77b0;
assign ad4271 = hlock1_p & ad4e94 | !hlock1_p & ad4f55;
assign c3d683 = hmaster2_p & c3d669 | !hmaster2_p & c3d66d;
assign b57413 = hlock3 & b57983 | !hlock3 & b57412;
assign ad426f = hbusreq1_p & ad426e | !hbusreq1_p & v845542;
assign c3d30f = hbusreq0 & c3d2f6 | !hbusreq0 & c3d30e;
assign ad4ea3 = hbusreq4_p & ad4ea2 | !hbusreq4_p & ad4e98;
assign v8cc78a = hmaster1_p & v8cc789 | !hmaster1_p & v845542;
assign bd58a0 = hburst1 & bd589d | !hburst1 & bd589f;
assign v8f96d9 = hburst1_p & v8f2540 | !hburst1_p & v845542;
assign b1cfcc = hgrant4_p & v845542 | !hgrant4_p & !b1cfcb;
assign ad46e9 = hmaster0_p & ad46e7 | !hmaster0_p & ad46e8;
assign c3d668 = stateA1_p & v845578 | !stateA1_p & !v845542;
assign df552f = hmaster1_p & v845542 | !hmaster1_p & df552e;
assign c3d6dd = hmaster0_p & c3d6b2 | !hmaster0_p & c3d6dc;
assign ad4601 = hmaster1_p & ad4600 | !hmaster1_p & ad45f8;
assign dc4fe8 = hgrant4_p & adec89 | !hgrant4_p & ade557;
assign v9ea603 = hgrant1_p & v9ea43a | !hgrant1_p & v9ea449;
assign ade4be = hburst1 & ade4bd | !hburst1 & v845566;
assign v93a916 = stateG3_1_p & v845542 | !stateG3_1_p & v845582;
assign d359a2 = hbusreq4_p & d359a0 | !hbusreq4_p & d359a1;
assign c3cebf = hbusreq4_p & v845542 | !hbusreq4_p & c3cebe;
assign ad4f53 = hgrant1_p & ad4f52 | !hgrant1_p & ad4e90;
assign v9ea599 = hbusreq2 & v9ea597 | !hbusreq2 & v9ea598;
assign df517f = hgrant1_p & df5533 | !hgrant1_p & !df517e;
assign b1c705 = hready_p & v845542 | !hready_p & b1c704;
assign d35011 = hbusreq4_p & d357c9 | !hbusreq4_p & d35010;
assign v8ccb6d = hmaster0_p & v8ccb6b | !hmaster0_p & v845542;
assign ad4f93 = hmaster2_p & ad4f90 | !hmaster2_p & ad4f92;
assign ad4ee1 = stateG10_4_p & v845542 | !stateG10_4_p & ad4ee0;
assign v9f7828 = hlock2 & v9f77d0 | !hlock2 & v9f7827;
assign d35bfa = hmaster0_p & d35bf4 | !hmaster0_p & d35bf9;
assign dc4fcc = hbusreq3 & dc4fcb | !hbusreq3 & v845542;
assign v9f7821 = hlock4 & v9f77c8 | !hlock4 & v9f7820;
assign b574b8 = hlock1 & b57942 | !hlock1 & b574b7;
assign ad415e = hready & ad4f7b | !hready & ad415d;
assign b1c5b8 = hbusreq0 & b1cf25 | !hbusreq0 & b1c5b7;
assign b1c7c9 = hbusreq4 & b1c7c2 | !hbusreq4 & b1c7c8;
assign b059c2 = locked_p & b059c1 | !locked_p & v9f7d42;
assign ad4331 = hgrant1_p & ad432e | !hgrant1_p & ad4330;
assign df51b4 = hmaster1_p & df51b3 | !hmaster1_p & df5163;
assign b05a45 = hbusreq2_p & b05a3c | !hbusreq2_p & b05a44;
assign b57ae5 = hlock3 & b579e5 | !hlock3 & b579e4;
assign dc5069 = hgrant2_p & dc4fdd | !hgrant2_p & dc5068;
assign v8cc5c6 = hbusreq2_p & v8cc5bb | !hbusreq2_p & v8cc5c5;
assign ad434f = hmaster0_p & ad434c | !hmaster0_p & ad428b;
assign ad4735 = hbusreq2 & ad4730 | !hbusreq2 & ad4733;
assign d35a38 = hmaster0_p & dc4fcb | !hmaster0_p & d35a37;
assign ad4fbb = hgrant4_p & v84556c | !hgrant4_p & cc36fc;
assign df51b0 = hbusreq2_p & df51aa | !hbusreq2_p & df51af;
assign c3d5af = decide_p & c3d5ae | !decide_p & !c3d36c;
assign v9ea589 = hlock0 & v9ea586 | !hlock0 & v9ea588;
assign d35512 = hbusreq4 & d35511 | !hbusreq4 & d3550b;
assign ad469f = hmaster2_p & ad469e | !hmaster2_p & v845542;
assign bd5b6c = hmastlock_p & bd5b6b | !hmastlock_p & v845542;
assign v9ea46a = hgrant4_p & v9ea403 | !hgrant4_p & v9f20a1;
assign c3d745 = hbusreq1_p & c3d6bd | !hbusreq1_p & c3d744;
assign b57427 = hlock3 & b57988 | !hlock3 & b57426;
assign v9ea5ad = hbusreq1 & v9ea58c | !hbusreq1 & v9ea58d;
assign b05928 = hmaster0_p & b0591d | !hmaster0_p & b0591e;
assign b1c03a = hbusreq1_p & b1c76a | !hbusreq1_p & b1c039;
assign bd5bb3 = hbusreq3_p & bd5ba1 | !hbusreq3_p & bd5bb2;
assign df5184 = hgrant1_p & v84556c | !hgrant1_p & !df5183;
assign v9ea495 = hbusreq3 & v9ea494 | !hbusreq3 & v9ea43b;
assign d35959 = hbusreq3 & d35958 | !hbusreq3 & v845542;
assign v9f7e3b = hmaster2_p & v9f7e14 | !hmaster2_p & v9f7c9f;
assign c5c936 = hgrant0_p & c5c92f | !hgrant0_p & v845542;
assign ad414f = hbusreq2 & ad414e | !hbusreq2 & v845542;
assign v9f7d12 = hmaster2_p & v9f7ca4 | !hmaster2_p & v9f7cc6;
assign v9ea57a = hmaster1_p & v9ea573 | !hmaster1_p & v9ea579;
assign v9ea46b = stateG10_4_p & v9f20a1 | !stateG10_4_p & v9ea46a;
assign c3d67f = hmaster1_p & c3d67e | !hmaster1_p & c3d67c;
assign b05a34 = hmaster0_p & b059fb | !hmaster0_p & b058c7;
assign ad45b9 = hmaster2_p & v845542 | !hmaster2_p & ad45b8;
assign ad5038 = hgrant1_p & c3d2d9 | !hgrant1_p & ad5023;
assign c3ce5e = hbusreq1_p & c3ce5d | !hbusreq1_p & v845564;
assign c5c88c = stateA1_p & c5c88b | !stateA1_p & !bb9bdd;
assign ad4db7 = hready & ad4dab | !hready & ad4db6;
assign d35996 = hgrant0_p & v84557a | !hgrant0_p & !v845542;
assign v8ccb7e = hlock0_p & v8d29fa | !hlock0_p & v845542;
assign ad5052 = hgrant4_p & ad502f | !hgrant4_p & !v84556c;
assign dc5036 = hburst0 & adec8d | !hburst0 & adec8e;
assign d354b6 = hmaster2_p & d354b5 | !hmaster2_p & d354a6;
assign ad42bf = hlock1_p & ad4da1 | !hlock1_p & !v845542;
assign ad4f2c = hbusreq1_p & ad4f2a | !hbusreq1_p & !ad4f2b;
assign v9ea496 = hlock2 & v9ea43b | !hlock2 & v9ea495;
assign v9ea45e = hgrant1_p & v9ea3fa | !hgrant1_p & v9ea45c;
assign ade54b = stateG2_p & v845542 | !stateG2_p & adec8b;
assign d35a77 = hmaster1_p & d35a76 | !hmaster1_p & d35a6c;
assign v9f7df0 = hlock1_p & v9f7cdd | !hlock1_p & v9f7d23;
assign c3ce5a = hmaster1_p & c3ce53 | !hmaster1_p & c3ce59;
assign v9f7e26 = hbusreq1 & v9f7e24 | !hbusreq1 & v9f7e25;
assign v8b08c2 = hburst1_p & v8b08c1 | !hburst1_p & v845542;
assign v9f7d1a = hbusreq1_p & v9f7d0c | !hbusreq1_p & v9f7d19;
assign b059e1 = hbusreq4_p & b05987 | !hbusreq4_p & !b059e0;
assign d356dc = hlock1_p & v845542 | !hlock1_p & d356db;
assign ad460a = hready & ad4609 | !hready & !v845564;
assign b1cf31 = hmaster2_p & v845542 | !hmaster2_p & b1cf30;
assign d35504 = hmaster0_p & d354fd | !hmaster0_p & !d35503;
assign c3d2f9 = hbusreq0 & c3d2f6 | !hbusreq0 & c3d2f8;
assign v9f7d43 = stateG10_4_p & v9f7d42 | !stateG10_4_p & v9f7cc6;
assign b05906 = hlock2 & b058c9 | !hlock2 & b05905;
assign ad4311 = hmaster0_p & ad4293 | !hmaster0_p & ad4291;
assign ad4dda = hgrant2_p & ad4dd7 | !hgrant2_p & ad4dd9;
assign d3571d = hbusreq1_p & d3571c | !hbusreq1_p & v845542;
assign d35988 = hbusreq4_p & v845542 | !hbusreq4_p & d35983;
assign v9ea582 = hbusreq1_p & v9ea3fc | !hbusreq1_p & v9ea581;
assign c5c99f = hmaster1_p & c5c99e | !hmaster1_p & v845542;
assign ad503d = hbusreq4_p & ad503a | !hbusreq4_p & ad503c;
assign v9ea48e = hlock0 & v9ea43b | !hlock0 & v9ea48d;
assign ade64f = decide_p & ade63c | !decide_p & adeaa7;
assign d3597d = decide_p & d3597c | !decide_p & v84556c;
assign ad4dd0 = hbusreq0 & ad4dae | !hbusreq0 & ad4dcf;
assign d3597b = hbusreq2_p & d35921 | !hbusreq2_p & d3597a;
assign df515e = hbusreq1 & ade4bf | !hbusreq1 & v845542;
assign v8cc0d3 = hlock3 & v8cc489 | !hlock3 & v8cc0d2;
assign b1c7fc = decide_p & b1c788 | !decide_p & !b1d013;
assign b05999 = hbusreq1 & b05997 | !hbusreq1 & b05998;
assign ad42f2 = hbusreq1_p & ad42f1 | !hbusreq1_p & v845542;
assign c3d6e7 = hmaster2_p & c3d6e3 | !hmaster2_p & c3d6e6;
assign c5c933 = hgrant4_p & c5c92f | !hgrant4_p & v845542;
assign b1c6b8 = hbusreq1 & b1cffc | !hbusreq1 & b1d002;
assign v8cc49c = hlock0 & v8cc494 | !hlock0 & v8cc49a;
assign bd57ae = hbusreq1_p & dc4f81 | !hbusreq1_p & dc4f91;
assign c3cf1f = hbusreq1 & c3cf1a | !hbusreq1 & c3cee4;
assign dc500d = hmaster2_p & dc4ff1 | !hmaster2_p & dc500c;
assign v9e9fa3 = hlock3 & v9e9f68 | !hlock3 & v9e9fa2;
assign v9f76e2 = locked_p & v9f76e1 | !locked_p & v9f7c9b;
assign v8cc4a3 = hlock0 & v8cc4a1 | !hlock0 & v8cc4a2;
assign b05a5f = stateG10_4_p & b05a5d | !stateG10_4_p & b05a5e;
assign ad4dcf = hmaster2_p & ad4dac | !hmaster2_p & !ad4dce;
assign ad439e = hmaster0_p & ad438c | !hmaster0_p & ad439d;
assign v9f7cc5 = stateA1_p & v845542 | !stateA1_p & !v9ea3e4;
assign ad45b2 = hlock4_p & ade4c1 | !hlock4_p & v845542;
assign b1c560 = hmaster2_p & b1c85e | !hmaster2_p & b1c55f;
assign d35bed = hmaster2_p & d35be3 | !hmaster2_p & d35be8;
assign d35a97 = hmaster1_p & v845542 | !hmaster1_p & d35a96;
assign v8ccb6b = hmaster2_p & v845542 | !hmaster2_p & v8ccb6a;
assign v9f771e = hmaster1_p & v9f76ab | !hmaster1_p & v9f76a6;
assign ad43a1 = hmaster0_p & v845547 | !hmaster0_p & ad4f1a;
assign v9e9eb3 = hbusreq3 & v9e9eb1 | !hbusreq3 & v9e9eb2;
assign d35a31 = hgrant1_p & d35a30 | !hgrant1_p & d359e1;
assign d35a69 = hmaster2_p & d35a5b | !hmaster2_p & d35a68;
assign ad3d20 = hready_p & ad3cc5 | !hready_p & ad3d1f;
assign b57af5 = hbusreq2_p & b57af4 | !hbusreq2_p & b57944;
assign ad4fa1 = hgrant2_p & v845542 | !hgrant2_p & !ad4f9f;
assign v8cc43d = hmaster1_p & v8ccbe5 | !hmaster1_p & v8cc43b;
assign df50cf = hmaster0_p & df50ce | !hmaster0_p & df54f4;
assign v9e9ecf = hmaster1_p & v9e9ece | !hmaster1_p & v9e9ead;
assign ade61f = hgrant2_p & ade61d | !hgrant2_p & ade61e;
assign v9f76b8 = hmaster0_p & v9f767b | !hmaster0_p & v9f7cc2;
assign bd5905 = jx1_p & bd572c | !jx1_p & bd5904;
assign b5743f = hgrant2_p & b5743e | !hgrant2_p & b5743b;
assign ad4ef2 = hbusreq4 & ad4ee9 | !hbusreq4 & ad4ef1;
assign b1cbfd = hbusreq4_p & b1d000 | !hbusreq4_p & b1cfcc;
assign ad4ea8 = hgrant1_p & ad4e97 | !hgrant1_p & ad4ea7;
assign ad4786 = hmaster0_p & ad473d | !hmaster0_p & ad460b;
assign b57509 = hbusreq3_p & b574fd | !hbusreq3_p & b57508;
assign d35952 = hbusreq1_p & d35951 | !hbusreq1_p & d3590a;
assign c3cf29 = hready_p & c3cefe | !hready_p & !c3cf28;
assign ad4e45 = stateA1_p & v845542 | !stateA1_p & af7f5a;
assign v9ea5a5 = hgrant1_p & v9ea578 | !hgrant1_p & v9ea59b;
assign b1c6cd = decide_p & b1c61a | !decide_p & b1d013;
assign v9ea59c = hbusreq4_p & v9ea471 | !hbusreq4_p & v9ea4d7;
assign bd575b = hmaster0_p & bd5754 | !hmaster0_p & bd575a;
assign d359db = hbusreq0 & d359d4 | !hbusreq0 & d359da;
assign d35bf9 = hbusreq3 & d35bf7 | !hbusreq3 & d35bf8;
assign dc538a = hmastlock_p & v8cc7d9 | !hmastlock_p & !v845542;
assign c5c895 = busreq_p & c5c88b | !busreq_p & !c5c894;
assign c3d2f0 = hgrant4_p & v845542 | !hgrant4_p & !c3d2ef;
assign b57a7a = hlock1 & b579ce | !hlock1 & b57a79;
assign d358f8 = hburst1 & d358eb | !hburst1 & v845542;
assign c5c9af = hmaster0_p & c5c8e9 | !hmaster0_p & c5c974;
assign ad4410 = hbusreq0 & ad440f | !hbusreq0 & v845542;
assign d35705 = hbusreq1_p & d35704 | !hbusreq1_p & v845542;
assign c3ceeb = decide_p & c3ceea | !decide_p & c3d36c;
assign c3d30a = hbusreq4_p & c3d308 | !hbusreq4_p & !c3d309;
assign v8cc0eb = hgrant2_p & v8cc472 | !hgrant2_p & v8cc0e9;
assign d35592 = hmaster0_p & d35588 | !hmaster0_p & d35591;
assign ad4de8 = hlock1_p & ad4de7 | !hlock1_p & v845542;
assign b059c7 = hbusreq4 & b059c5 | !hbusreq4 & b059c6;
assign bd58d3 = hbusreq4 & bd58cc | !hbusreq4 & bd58d2;
assign aa425c = jx1_p & v85746e | !jx1_p & v845542;
assign ad43d4 = hbusreq3 & ad43cd | !hbusreq3 & ad43d3;
assign v9f7819 = hmaster1_p & v9f7818 | !hmaster1_p & v9f77b0;
assign b1c85b = hlock0_p & v84556e | !hlock0_p & !v845548;
assign ad4297 = hmaster0_p & df5148 | !hmaster0_p & ad4296;
assign d35718 = hbusreq2 & d35717 | !hbusreq2 & !v84554e;
assign v9ea47c = hlock0 & v9ea47a | !hlock0 & v9ea47b;
assign v9f7746 = hlock0 & v9f7745 | !hlock0 & v9f7744;
assign c3d353 = hgrant1_p & v84554d | !hgrant1_p & c3d32a;
assign c3d59e = stateA1_p & c3d59d | !stateA1_p & c5c8e2;
assign b1cbfe = hmaster2_p & b1cfcc | !hmaster2_p & b1cbfd;
assign c3cf15 = hbusreq2_p & c3cf11 | !hbusreq2_p & c3cf14;
assign v8cc4b6 = hbusreq3 & v8cc4b4 | !hbusreq3 & v8ccbd8;
assign d35803 = decide_p & d35802 | !decide_p & v84556c;
assign v9f7812 = hmaster1_p & v9f77d4 | !hmaster1_p & v9f7811;
assign b1c056 = hgrant2_p & b1c055 | !hgrant2_p & b1c051;
assign ad46fe = hbusreq4_p & ad46fd | !hbusreq4_p & v845542;
assign ad4603 = hmaster1_p & ad4602 | !hmaster1_p & ad45f8;
assign v9e9eee = hbusreq1_p & v9e9ee9 | !hbusreq1_p & v9e9eed;
assign ad416b = hmaster0_p & ad4169 | !hmaster0_p & ad416a;
assign ade578 = hgrant4_p & v84556c | !hgrant4_p & !adeca1;
assign v9f78ab = decide_p & v9f7873 | !decide_p & v9f78aa;
assign dc5056 = hgrant4_p & v845542 | !hgrant4_p & !ade58d;
assign b0594b = hmaster1_p & b0594a | !hmaster1_p & b058e1;
assign ad4403 = hbusreq3 & ad43db | !hbusreq3 & ad43dd;
assign d35723 = decide_p & d35722 | !decide_p & v84556c;
assign v9f7d4a = hmaster1_p & v9f7d49 | !hmaster1_p & v9f7d47;
assign bd5886 = stateG10_4_p & bd5865 | !stateG10_4_p & !bd5885;
assign bd580f = hgrant4_p & c3d66d | !hgrant4_p & bd580d;
assign b059c6 = hlock4 & b058a8 | !hlock4 & b059c5;
assign v8cc592 = hlock0 & v8ccbd8 | !hlock0 & v8cc590;
assign v9e9ee4 = hgrant3_p & v9e9edd | !hgrant3_p & v9e9ee3;
assign c3d71f = hmaster1_p & c3d71e | !hmaster1_p & c3d68b;
assign b5b407 = hmastlock_p & b0ed8b | !hmastlock_p & v845542;
assign b05a29 = hbusreq2_p & b05a22 | !hbusreq2_p & b05a28;
assign v9f76de = hburst1_p & v9fa31b | !hburst1_p & !v9f7cf2;
assign ad4817 = hbusreq2 & ad4816 | !hbusreq2 & v845542;
assign ad477b = hbusreq0 & ad45ee | !hbusreq0 & ad477a;
assign ad4fd8 = hbusreq4_p & ad4fd5 | !hbusreq4_p & ad4fd7;
assign ad4ef9 = hgrant4_p & v845542 | !hgrant4_p & !ad4ef7;
assign v9ea567 = hmaster2_p & v9f20a1 | !hmaster2_p & v9ea566;
assign ad416c = hmaster1_p & ad4168 | !hmaster1_p & ad416b;
assign c3d5f3 = hready & c3d5f2 | !hready & c3d300;
assign dc4f87 = hbusreq2 & dc4f85 | !hbusreq2 & dc4f86;
assign b1c45d = hready_p & b1cc05 | !hready_p & b1c45c;
assign b1c78e = hbusreq2 & b1c723 | !hbusreq2 & b1c71d;
assign c3d519 = hbusreq2 & c3d513 | !hbusreq2 & c3d517;
assign b058f5 = hlock2 & b058ea | !hlock2 & b058f3;
assign c3d517 = hgrant1_p & v845542 | !hgrant1_p & c3d516;
assign df5175 = hmaster0_p & df516f | !hmaster0_p & df5174;
assign c3d504 = hready & c3d500 | !hready & c3d503;
assign b1c7e6 = hbusreq2 & b1c739 | !hbusreq2 & !v845542;
assign c3d317 = hmaster0_p & c3d307 | !hmaster0_p & c3d316;
assign v9ea487 = hbusreq3 & v9ea485 | !hbusreq3 & v9ea486;
assign v9f76a2 = stateG10_4_p & v9f7663 | !stateG10_4_p & v9f76a1;
assign b57984 = stateG10_4_p & v845542 | !stateG10_4_p & b5794f;
assign d3571b = hbusreq1 & d359e1 | !hbusreq1 & v845542;
assign b1c5d9 = hbusreq2 & b1c5bf | !hbusreq2 & b1c5d8;
assign v9e9f9d = hlock2 & v9e9f9a | !hlock2 & v9e9f9c;
assign ad4efa = stateG10_4_p & ad4ef7 | !stateG10_4_p & !ad4ef9;
assign v9ea45f = hbusreq3 & v9ea45d | !hbusreq3 & v9ea45e;
assign d35020 = hgrant2_p & d357ef | !hgrant2_p & d3501f;
assign bd577f = hlock3_p & bd5767 | !hlock3_p & bd577e;
assign bd57bc = hburst0_p & c74a04 | !hburst0_p & !bd57bb;
assign v9f7cf2 = start_p & v845542 | !start_p & !v9fa31b;
assign v9f7d34 = hbusreq2 & v9f7d32 | !hbusreq2 & v9f7d33;
assign b05a62 = locked_p & b05a58 | !locked_p & !b058a3;
assign ad4422 = hmaster0_p & ad4420 | !hmaster0_p & ad4421;
assign ad4805 = hgrant3_p & ad4789 | !hgrant3_p & !ad4804;
assign b8f74c = hgrant2_p & v845542 | !hgrant2_p & !b8f74b;
assign v9e9fdd = hmaster0_p & v9ea49a | !hmaster0_p & v9ea44a;
assign c3d6b0 = hbusreq4_p & c3d6ad | !hbusreq4_p & c3d6af;
assign v9ea5cd = hlock0 & v9ea5cb | !hlock0 & v9ea5cc;
assign bd5b72 = hmaster0_p & v845542 | !hmaster0_p & bd5b71;
assign ad4355 = hmaster1_p & ad4354 | !hmaster1_p & ad4297;
assign b1c72a = hbusreq3 & b1c727 | !hbusreq3 & b1c729;
assign v9f7739 = hmaster1_p & v9f7738 | !hmaster1_p & v9f7736;
assign ad3d0e = hmaster2_p & ad3d0d | !hmaster2_p & v845542;
assign b1c053 = hbusreq2 & b1c73e | !hbusreq2 & !v845542;
assign b574c7 = hready & b574c6 | !hready & b579ce;
assign ad3d5b = hready_p & ad3d4b | !hready_p & ad3d5a;
assign ade5a9 = hmaster0_p & ade5a7 | !hmaster0_p & ade5a8;
assign c3ce9b = hmaster2_p & c3d30d | !hmaster2_p & !v845542;
assign bd588e = hbusreq4_p & bd588b | !hbusreq4_p & bd588d;
assign ad443a = hbusreq0 & ad4439 | !hbusreq0 & v845542;
assign c3ce50 = hgrant2_p & v845551 | !hgrant2_p & c3ce4f;
assign d3568d = hready_p & d3568a | !hready_p & d3568c;
assign c3d5ef = hbusreq0 & c3d5d8 | !hbusreq0 & c3d5ee;
assign v9f775d = hlock4 & v9f775a | !hlock4 & v9f775c;
assign ad42e2 = hlock1_p & ad42e1 | !hlock1_p & ad426d;
assign b1c79a = stateG10_4_p & b1c797 | !stateG10_4_p & !b1c799;
assign v8cc5a6 = hbusreq4_p & v8cc499 | !hbusreq4_p & v8cc493;
assign b57a25 = hbusreq4_p & b57949 | !hbusreq4_p & b5b4ef;
assign bd57f5 = hburst1 & ade54d | !hburst1 & bd57f4;
assign v9ea48f = hbusreq0 & v9ea48d | !hbusreq0 & v9ea48e;
assign c3d343 = hgrant4_p & v845542 | !hgrant4_p & c3d33b;
assign bd5817 = hbusreq4_p & bd5814 | !hbusreq4_p & bd5816;
assign ad3cc0 = hgrant1_p & ad43aa | !hgrant1_p & ad4484;
assign c3ce76 = hbusreq3 & c3ce75 | !hbusreq3 & c3ce37;
assign v9f764b = hbusreq1_p & v9f7ca7 | !hbusreq1_p & v9f7e32;
assign af7f5a = hburst0_p & c74202 | !hburst0_p & af7f59;
assign ad5030 = hmaster2_p & v84556c | !hmaster2_p & !ad502f;
assign b05a74 = hgrant1_p & b058c7 | !hgrant1_p & b05a73;
assign v9e9edf = hmaster1_p & v9ea44a | !hmaster1_p & v9ea4db;
assign c3d35b = hgrant1_p & v84554d | !hgrant1_p & c3d300;
assign ad4fc1 = hmaster2_p & ad4fbd | !hmaster2_p & v84556c;
assign ad506f = decide_p & ad4e20 | !decide_p & ad506e;
assign ade5ab = hmaster2_p & ade548 | !hmaster2_p & !ade5aa;
assign v9ea459 = stateG10_4_p & v9ea457 | !stateG10_4_p & v9ea458;
assign b059d6 = stateG10_4_p & v9f7d42 | !stateG10_4_p & b059d5;
assign v9e9fab = hlock3 & v9e9faa | !hlock3 & v9e9fa9;
assign bd5940 = jx1_p & bd593f | !jx1_p & bd5bb2;
assign b058e4 = hmaster1_p & b058e3 | !hmaster1_p & b058e1;
assign df5538 = hbusreq1_p & v84556c | !hbusreq1_p & !v845542;
assign b1c7cd = hbusreq1 & b1c743 | !hbusreq1 & !v845542;
assign ba7c7a = hmaster0_p & ba7c6b | !hmaster0_p & ba7c79;
assign v8ccbe3 = hmaster2_p & v8ccbe2 | !hmaster2_p & v845542;
assign v9ea592 = hbusreq1_p & v9ea449 | !hbusreq1_p & v9ea591;
assign c3d37a = hgrant1_p & v845542 | !hgrant1_p & c3d379;
assign cc36e3 = hbusreq4_p & cc36e1 | !hbusreq4_p & !cc36e2;
assign v9f7770 = hbusreq3 & v9f7757 | !hbusreq3 & v9f776f;
assign c3d50e = decide_p & c3d508 | !decide_p & c3d50d;
assign d35be7 = hlock4_p & v845542 | !hlock4_p & v84556c;
assign v9ea5b5 = hmaster0_p & v9ea44a | !hmaster0_p & v9ea5b4;
assign c749e5 = stateG3_0_p & v845580 | !stateG3_0_p & !v845542;
assign d35599 = hmaster2_p & d35a9b | !hmaster2_p & d35598;
assign dc5307 = hmaster0_p & dc5303 | !hmaster0_p & v84556c;
assign ad4def = hbusreq4 & ad4dec | !hbusreq4 & ad4dee;
assign c3d534 = decide_p & c3d533 | !decide_p & !c3d36c;
assign d3572d = hmaster0_p & d3572a | !hmaster0_p & d3572c;
assign ad5057 = hbusreq0 & ad5055 | !hbusreq0 & ad5056;
assign c3d728 = hmaster1_p & c3d727 | !hmaster1_p & c3d68b;
assign v8cc4df = hgrant3_p & v8ccbdc | !hgrant3_p & v8cc4dd;
assign v845578 = busreq_p & v845542 | !busreq_p & !v845542;
assign v8cc5bb = hgrant2_p & v8cc472 | !hgrant2_p & v8cc5ba;
assign c3d6a1 = hready_p & c3d691 | !hready_p & !c3d6a0;
assign c3d31a = stateG10_4_p & c3d318 | !stateG10_4_p & c3d319;
assign bd58fe = hlock2_p & bd58fd | !hlock2_p & !bd58d8;
assign v9f7d0c = hbusreq1 & v9f7d0a | !hbusreq1 & v9f7d0b;
assign v9ea464 = hgrant0_p & v9ea463 | !hgrant0_p & !v9ea3e9;
assign c3d361 = hmaster1_p & c3d35f | !hmaster1_p & c3d360;
assign b059fe = hmaster0_p & b059bd | !hmaster0_p & b059a9;
assign b1c7c7 = hmaster2_p & b1c7a7 | !hmaster2_p & b1c7c6;
assign bd5b99 = hgrant2_p & bd5b98 | !hgrant2_p & !v845542;
assign v9f7732 = hbusreq4_p & v845542 | !hbusreq4_p & !v9f772f;
assign v9ea4bc = hmaster2_p & v9ea4b9 | !hmaster2_p & v9ea4bb;
assign ad45fc = hmaster1_p & ad45fb | !hmaster1_p & ad45f8;
assign d354c7 = hbusreq1 & d35bf7 | !hbusreq1 & d35bf8;
assign b579c2 = hbusreq1 & b579c1 | !hbusreq1 & b57942;
assign b0599f = hbusreq2 & b0599d | !hbusreq2 & b0599e;
assign b0596a = hbusreq1_p & b05969 | !hbusreq1_p & b058e8;
assign b1c809 = hbusreq0 & v845542 | !hbusreq0 & !d35a9c;
assign ad4fae = locked_p & ad4fad | !locked_p & !v845542;
assign v9f7d9c = hlock3 & v9f7d9b | !hlock3 & v9f7d98;
assign ad4143 = hbusreq4 & ad4139 | !hbusreq4 & ad4142;
assign v9f7dd6 = hmaster2_p & v9f7dcd | !hmaster2_p & v9f7dd5;
assign v8cc762 = hgrant2_p & v8cc472 | !hgrant2_p & v8cc761;
assign c3cdfe = hbusreq2 & c3d306 | !hbusreq2 & c3d32f;
assign b573e0 = hgrant2_p & b579b0 | !hgrant2_p & b573df;
assign b57abe = hmastlock_p & b57abd | !hmastlock_p & v845542;
assign c3d3a1 = hmaster2_p & c3d3a0 | !hmaster2_p & v845576;
assign v9f7768 = hlock4_p & v84557a | !hlock4_p & !v845542;
assign ad4f47 = hbusreq2 & ad4f46 | !hbusreq2 & v845542;
assign v9f7d45 = hlock0_p & v9f7c9d | !hlock0_p & v9f7d21;
assign ad457a = hmaster2_p & v845542 | !hmaster2_p & ad4579;
assign b05a8c = hbusreq2_p & b05a87 | !hbusreq2_p & b05a8b;
assign ad4765 = hbusreq4_p & ad4764 | !hbusreq4_p & !v845542;
assign d35a51 = hbusreq1 & df54f5 | !hbusreq1 & d35a50;
assign d35abb = hready_p & d35aba | !hready_p & d35aa2;
assign c3d700 = hmaster1_p & c3d6ff | !hmaster1_p & c3d67c;
assign ade4d3 = hburst1 & c3d674 | !hburst1 & !v845566;
assign b579d0 = hbusreq0_p & b579cc | !hbusreq0_p & b579cf;
assign b573de = hmaster0_p & b579c5 | !hmaster0_p & b573dd;
assign b059cb = hbusreq1_p & b058b1 | !hbusreq1_p & b059ca;
assign b05a7e = hbusreq3 & b05a7a | !hbusreq3 & b05a7d;
assign d356cd = hmaster0_p & d356c2 | !hmaster0_p & d356cc;
assign ade5ba = decide_p & ade4f1 | !decide_p & adeaa7;
assign b1c7d7 = hbusreq0_p & dc5050 | !hbusreq0_p & v845542;
assign c3d324 = hbusreq4 & c3d31d | !hbusreq4 & !c3d323;
assign v9e9ebf = decide_p & v9e9e75 | !decide_p & v9e9ebe;
assign b1cf25 = hmaster2_p & v845542 | !hmaster2_p & !b1cf24;
assign ba7c71 = hready_p & ba7c6f | !hready_p & ba7c70;
assign b058a1 = busreq_p & v845582 | !busreq_p & !b058a0;
assign c3cea8 = hgrant2_p & c3ce95 | !hgrant2_p & c3cea7;
assign bd578f = hburst1 & d3561d | !hburst1 & bd578e;
assign b1c7b6 = hlock0_p & ade572 | !hlock0_p & v845542;
assign c3d521 = hready_p & c3d50e | !hready_p & c3d520;
assign b058fe = hlock3 & b058b8 | !hlock3 & b058fd;
assign b57ac2 = hlock4 & b578f9 | !hlock4 & b57ac1;
assign v9f765e = hgrant4_p & v9f7e31 | !hgrant4_p & !v9f7dad;
assign v845560 = hmaster0_p & v845542 | !hmaster0_p & !v845542;
assign ad3d07 = hbusreq4_p & ad3d06 | !hbusreq4_p & ad3d01;
assign v9ea426 = hmaster1_p & v9ea410 | !hmaster1_p & v9ea425;
assign c5c9b2 = hbusreq2_p & c5c9ae | !hbusreq2_p & c5c9b1;
assign b058b9 = hlock0 & b058b8 | !hlock0 & b058b7;
assign v9f7d73 = hgrant4_p & v9f7c9c | !hgrant4_p & v9f7d72;
assign c3d374 = hgrant4_p & v845542 | !hgrant4_p & c3d373;
assign adea95 = hgrant1_p & v845542 | !hgrant1_p & !adea94;
assign c3d2c4 = hburst1 & c3d2ad | !hburst1 & v845542;
assign b058b0 = hlock1 & b058aa | !hlock1 & b058af;
assign d35ab6 = hmaster0_p & d35aaf | !hmaster0_p & d35ab5;
assign ad4e6a = stateA1_p & v845542 | !stateA1_p & !ad4e69;
assign v9ea433 = hmaster0_p & v9ea42d | !hmaster0_p & v9ea432;
assign c5c99a = hbusreq2_p & c5c979 | !hbusreq2_p & c5c999;
assign d357f7 = hbusreq1_p & d35799 | !hbusreq1_p & d357f6;
assign v9f769e = hgrant4_p & v9f7e31 | !hgrant4_p & v9f7694;
assign d35440 = hmaster1_p & d3542e | !hmaster1_p & d35438;
assign c3ce41 = decide_p & c3ce40 | !decide_p & !c3d36c;
assign b05a00 = hgrant2_p & b059fd | !hgrant2_p & b059ff;
assign ad3d08 = hmaster2_p & ad3d07 | !hmaster2_p & v845542;
assign ad4ebc = hbusreq4_p & ad4eb9 | !hbusreq4_p & ad4ebb;
assign d35619 = hburst1_p & v857b36 | !hburst1_p & !c74a04;
assign dc5041 = hmaster2_p & dc503c | !hmaster2_p & dc5040;
assign v9f7726 = hmaster2_p & d35aaa | !hmaster2_p & !v845542;
assign b1c033 = hmaster2_p & b1c030 | !hmaster2_p & b1c032;
assign c3d73a = hlock2_p & c3d736 | !hlock2_p & !c3d739;
assign ad42d8 = hbusreq1_p & ad42d7 | !hbusreq1_p & v845542;
assign c3cea3 = hmaster0_p & c3cea1 | !hmaster0_p & c3cea2;
assign v9e9f76 = stateG10_4_p & v9e9f74 | !stateG10_4_p & v9e9f75;
assign cc36d7 = decide_p & cc36d6 | !decide_p & v84556c;
assign v9f7de8 = hlock0 & v9f7de7 | !hlock0 & v9f7dd6;
assign bd57e1 = hmaster0_p & bd57d2 | !hmaster0_p & !bd57e0;
assign d359ee = hburst0 & d359ed | !hburst0 & v845542;
assign c3d74a = hmaster1_p & c3d746 | !hmaster1_p & c3d749;
assign d3594d = hburst1 & dc5318 | !hburst1 & d3594c;
assign d35be2 = hlock4_p & d3597f | !hlock4_p & v84556c;
assign bd583d = stateG10_4_p & bd574e | !stateG10_4_p & !bd583c;
assign ac145c = hmaster2_p & ac145b | !hmaster2_p & v845542;
assign ad4f4c = hready & ad4f4b | !hready & v84556c;
assign b1cf3b = hbusreq0 & b1cf25 | !hbusreq0 & b1cf3a;
assign v9f7696 = stateG10_4_p & v9f7694 | !stateG10_4_p & v9f7695;
assign bd58e5 = hready_p & bd58db | !hready_p & !bd58e4;
assign c3cf16 = decide_p & c3ceea | !decide_p & c3cf15;
assign v9f7e30 = hmaster2_p & v9f7c9c | !hmaster2_p & !v9f7e2f;
assign c5c93d = hmaster1_p & c5c8f5 | !hmaster1_p & c5c93c;
assign ad4823 = hbusreq2 & ad4fb4 | !hbusreq2 & v845542;
assign df51bb = hmaster0_p & df51ba | !hmaster0_p & df5174;
assign bd57fb = locked_p & bd57f6 | !locked_p & bd57fa;
assign ad4f1f = hbusreq1_p & ad4e95 | !hbusreq1_p & ad4f1e;
assign b1c851 = hgrant1_p & v845542 | !hgrant1_p & b1c850;
assign ad41b9 = hready_p & ad41b3 | !hready_p & ad41b8;
assign ad4f5e = hready & ad4ea6 | !hready & ad4ec5;
assign b1c856 = hgrant4_p & v84554a | !hgrant4_p & !b1c855;
assign b8ef53 = jx2_p & b8f747 | !jx2_p & b8ef52;
assign ad4fb2 = hmaster0_p & dc4fcc | !hmaster0_p & ad4fb1;
assign v9ea3f0 = hmaster0_p & v9ea3e8 | !hmaster0_p & v9ea3ef;
assign v8cc0f1 = hlock2 & v8ccbd8 | !hlock2 & v8cc0f0;
assign v9e9f67 = hlock0_p & v9e9f66 | !hlock0_p & v9ea4b3;
assign c3cef6 = hbusreq0 & c3cef5 | !hbusreq0 & v845542;
assign ad3ce1 = locked_p & ad5032 | !locked_p & v845542;
assign d35a6c = hmaster0_p & d35a55 | !hmaster0_p & d35a6b;
assign b1c069 = hbusreq4_p & b1c7bd | !hbusreq4_p & !b1c068;
assign c5c901 = hmaster0_p & c5c8f8 | !hmaster0_p & c5c900;
assign b1c4cb = hmaster2_p & d35a9c | !hmaster2_p & b1c4ca;
assign dc5300 = locked_p & dc52ff | !locked_p & v845542;
assign ad4574 = hmaster2_p & ad4554 | !hmaster2_p & ad4573;
assign c74a04 = start_p & v845542 | !start_p & !v857b36;
assign v9ea3e5 = stateG2_p & v845542 | !stateG2_p & v9ea3e4;
assign ad502c = hbusreq2 & ad5028 | !hbusreq2 & ad502b;
assign dc53a6 = hmaster1_p & dc53a5 | !hmaster1_p & v845542;
assign v9f77a2 = hlock4 & v9f779f | !hlock4 & v9f77a1;
assign dc4fc5 = hbusreq2_p & dc4fb3 | !hbusreq2_p & dc4fc4;
assign dc5023 = stateG10_4_p & ade563 | !stateG10_4_p & !dc5022;
assign c3ce87 = decide_p & c3ce86 | !decide_p & c3ce5b;
assign ad3d14 = hgrant2_p & ad3cc9 | !hgrant2_p & ad3d13;
assign dc4f73 = hbusreq3 & dc4f72 | !hbusreq3 & v845542;
assign ad4f40 = hready & ad4f3d | !hready & ad4f3f;
assign c3d676 = hmaster2_p & c3d66a | !hmaster2_p & c3d675;
assign v8cc827 = hbusreq2 & v8cc825 | !hbusreq2 & v8cc826;
assign b1c84a = hmaster0_p & b1c842 | !hmaster0_p & b1c849;
assign bd589b = busreq_p & v84557c | !busreq_p & !v845542;
assign v8cc5c5 = hgrant2_p & v8cc5c4 | !hgrant2_p & v8cc5ba;
assign v9f788b = hlock1 & v9f77d8 | !hlock1 & v9f788a;
assign v9f7d96 = hlock1 & v9f7d90 | !hlock1 & v9f7d95;
assign ad3d4e = hmaster0_p & ad4413 | !hmaster0_p & ad440e;
assign cc3702 = hbusreq1_p & cc36cd | !hbusreq1_p & cc3701;
assign bd5930 = hmaster2_p & v84556c | !hmaster2_p & bd592f;
assign d35728 = hmaster1_p & d35727 | !hmaster1_p & d356c9;
assign c3ce1b = hbusreq2 & c3ce1a | !hbusreq2 & c3d368;
assign ad4703 = hmaster2_p & ad46fe | !hmaster2_p & v845542;
assign b574c4 = hbusreq0 & b574c3 | !hbusreq0 & b579ce;
assign d357d7 = hlock4_p & d357d6 | !hlock4_p & d357c8;
assign b0590d = hlock1 & b058d5 | !hlock1 & b0590c;
assign ac147a = hmaster2_p & ac1476 | !hmaster2_p & !ac1479;
assign dc5006 = hbusreq4_p & dc5003 | !hbusreq4_p & dc5005;
assign d35c09 = hbusreq1_p & d35c01 | !hbusreq1_p & d35c08;
assign ad45ac = hmaster2_p & ad4d91 | !hmaster2_p & ad45ab;
assign ade55d = hbusreq4_p & ade55c | !hbusreq4_p & !v845542;
assign b058c8 = hbusreq1_p & b058c1 | !hbusreq1_p & b058c7;
assign ac1493 = hready_p & ac1492 | !hready_p & !v845542;
assign v8cc62e = hmaster0_p & v8cc62d | !hmaster0_p & v845542;
assign ad4e41 = hready_p & v845542 | !hready_p & ad4e40;
assign v9f7675 = hmaster0_p & v9f7651 | !hmaster0_p & !v9f7674;
assign ac1474 = hgrant1_p & ac144f | !hgrant1_p & ac145c;
assign v9e9f6a = hlock0_p & v9ea44c | !hlock0_p & v9e9f69;
assign c3cecc = hbusreq4_p & c3d2fd | !hbusreq4_p & c3cecb;
assign ad4274 = hmaster0_p & ad4270 | !hmaster0_p & ad4273;
assign v9e9f89 = hgrant0_p & v9ea463 | !hgrant0_p & v845542;
assign adec9d = hbusreq3 & adec92 | !hbusreq3 & adec9c;
assign ad43d9 = hbusreq1 & ad43cd | !hbusreq1 & ad43d3;
assign v9f77d5 = hlock1_p & v9f772c | !hlock1_p & v9f772d;
assign d35763 = hmaster0_p & d35aaf | !hmaster0_p & d35aae;
assign v9ea5fa = hready_p & v9ea3e3 | !hready_p & v9ea5f9;
assign d35abc = hgrant3_p & d35aa3 | !hgrant3_p & !d35abb;
assign b05947 = hbusreq2_p & b05944 | !hbusreq2_p & b05946;
assign v9ea4d5 = hlock0_p & v9f20a1 | !hlock0_p & v9ea4d4;
assign df5115 = hbusreq3_p & df50d5 | !hbusreq3_p & df5114;
assign v9f7e2e = hmastlock_p & v9f7e2d | !hmastlock_p & v845542;
assign df5542 = hready_p & df5540 | !hready_p & df5541;
assign ad4f73 = hbusreq0 & ad4f6c | !hbusreq0 & ad4f72;
assign df514d = hmaster0_p & df5149 | !hmaster0_p & df514c;
assign adeaae = hbusreq4_p & v845566 | !hbusreq4_p & !v845542;
assign b1c5bd = hbusreq0 & b1cf25 | !hbusreq0 & b1c5bc;
assign d359c5 = hmaster2_p & v845542 | !hmaster2_p & !d359c4;
assign b0598e = hlock0_p & b0598b | !hlock0_p & !b0598d;
assign df5199 = hbusreq1 & dc502d | !hbusreq1 & v845542;
assign d35c04 = hbusreq3 & d35c01 | !hbusreq3 & !d35c03;
assign b57402 = decide_p & b57a21 | !decide_p & b573f7;
assign bd5809 = stateG10_4_p & bd5806 | !stateG10_4_p & bd5808;
assign v9e9fe6 = hbusreq3_p & v9e9fd8 | !hbusreq3_p & v9e9fe5;
assign df50db = hmaster0_p & df50da | !hmaster0_p & v845542;
assign v9ea44b = stateA1_p & b06719 | !stateA1_p & c6d407;
assign ad46d9 = hmaster2_p & v845542 | !hmaster2_p & ad46d8;
assign b05a24 = hmaster1_p & b05a23 | !hmaster1_p & b05943;
assign v8cc629 = hgrant3_p & v8ccbdc | !hgrant3_p & v8cc628;
assign ade4e6 = hburst0 & v845542 | !hburst0 & ade4e5;
assign d35018 = hbusreq1_p & d357d4 | !hbusreq1_p & d357ec;
assign v9f7df6 = hbusreq2 & v9f7df4 | !hbusreq2 & v9f7df5;
assign v9f7885 = hbusreq4_p & v9f77bf | !hbusreq4_p & v9f7884;
assign v9f7d56 = hlock3_p & v9f7d4e | !hlock3_p & v9f7d55;
assign ad4579 = hbusreq4_p & ad4e5c | !hbusreq4_p & v845542;
assign dc506c = hbusreq3 & dc5019 | !hbusreq3 & v845542;
assign d35911 = hbusreq3 & d35910 | !hbusreq3 & v845542;
assign dc4f67 = hbusreq3 & dc4f66 | !hbusreq3 & v845564;
assign d355a2 = hbusreq3_p & d354ed | !hbusreq3_p & !d355a1;
assign b573e8 = hmaster1_p & b573e7 | !hmaster1_p & v845542;
assign ad4163 = hgrant2_p & v845542 | !hgrant2_p & ad4162;
assign bd582f = hbusreq4 & bd582b | !hbusreq4 & bd582e;
assign ad4e92 = hgrant1_p & ad4e67 | !hgrant1_p & ad4e91;
assign v9ea409 = hbusreq2_p & v9ea406 | !hbusreq2_p & v9ea408;
assign d35989 = hbusreq0_p & v845542 | !hbusreq0_p & d35983;
assign v8cc7fc = hlock0 & v8cc439 | !hlock0 & v8cc7fa;
assign v8cc7aa = hready_p & v8cc7a8 | !hready_p & v8ccbdb;
assign b57a72 = hlock2 & b579c5 | !hlock2 & b57a71;
assign d354d3 = hmaster0_p & d354c6 | !hmaster0_p & d354d2;
assign ad4f04 = hbusreq4_p & ad4f01 | !hbusreq4_p & ad4f03;
assign c3d6f9 = hbusreq4_p & c3d6f7 | !hbusreq4_p & !c3d6f8;
assign d35568 = hmaster0_p & d354e6 | !hmaster0_p & d354b8;
assign ad4f60 = hgrant1_p & ad4f5d | !hgrant1_p & ad4f5f;
assign df5135 = jx1_p & df5115 | !jx1_p & df5134;
assign df5192 = hbusreq1_p & df5191 | !hbusreq1_p & v845542;
assign c3ce80 = hgrant1_p & v84554d | !hgrant1_p & c3ce7f;
assign b1c7f1 = hmaster1_p & b1c7f0 | !hmaster1_p & b1c7eb;
assign ad3d46 = hmaster0_p & ad43aa | !hmaster0_p & ad448f;
assign b579c9 = hgrant4_p & b57941 | !hgrant4_p & v845542;
assign v9ea49e = hbusreq2_p & v9ea48c | !hbusreq2_p & v9ea49d;
assign c3d522 = hgrant3_p & c3d484 | !hgrant3_p & c3d521;
assign ac1464 = hbusreq4_p & ac1462 | !hbusreq4_p & !ac1463;
assign stateG3_1 = !v8cc170;
assign v9f779a = hlock2 & v9f772d | !hlock2 & v9f7799;
assign d3590a = hmaster2_p & d35909 | !hmaster2_p & !v845542;
assign ad4381 = hbusreq0_p & ad4f38 | !hbusreq0_p & v845542;
assign b57533 = hready_p & b5799c | !hready_p & b57532;
assign b579e2 = hlock1 & b579ce | !hlock1 & b579e1;
assign c3d339 = hbusreq4_p & c3d337 | !hbusreq4_p & c3d338;
assign v9f77aa = hlock2 & v9f77a7 | !hlock2 & v9f77a9;
assign ad42c5 = hmaster1_p & ad42c4 | !hmaster1_p & ad42bd;
assign b059a1 = hmaster1_p & b05968 | !hmaster1_p & b059a0;
assign ad4470 = hbusreq1 & ad4393 | !hbusreq1 & v845542;
assign v9f7de1 = hlock0_p & v9f7ddd | !hlock0_p & v9f7de0;
assign ade4ec = hmaster0_p & ade4dd | !hmaster0_p & !ade4eb;
assign b05976 = hlock1_p & b058dc | !hlock1_p & b0590e;
assign ad4eb8 = hmaster2_p & ad4e73 | !hmaster2_p & ad4eb7;
assign ad3cf0 = hbusreq0 & ad3cef | !hbusreq0 & v845542;
assign v9f7809 = hbusreq4_p & d35a0b | !hbusreq4_p & !v9f77e9;
assign v9f7dcf = hgrant0_p & v9f7cf5 | !hgrant0_p & v9f7c9f;
assign v9f778c = hbusreq1 & v9f778a | !hbusreq1 & v9f778b;
assign v9ea41d = locked_p & v9ea411 | !locked_p & v845542;
assign d35419 = hbusreq4_p & d35418 | !hbusreq4_p & v845542;
assign ade5b1 = hbusreq1 & ade4a6 | !hbusreq1 & adec93;
assign d35aa9 = hlock2_p & d35aa8 | !hlock2_p & d35aa7;
assign b1c74a = hbusreq2_p & b1c746 | !hbusreq2_p & b1c749;
assign d35a1f = hbusreq2 & d359ad | !hbusreq2 & !d359c5;
assign v9f781e = hmaster2_p & v9f781d | !hmaster2_p & !v845542;
assign b05a19 = stateG10_4_p & v9f769d | !stateG10_4_p & b05a18;
assign b05a6b = hbusreq0 & b05a61 | !hbusreq0 & b05a6a;
assign ad3d0b = hgrant4_p & ad3ce2 | !hgrant4_p & v845542;
assign b05a12 = stateG10_4_p & v9f769d | !stateG10_4_p & b05a11;
assign hgrant4 = !ade667;
assign ad5027 = hgrant1_p & ad501b | !hgrant1_p & ad5026;
assign v9ea471 = hgrant4_p & v9ea403 | !hgrant4_p & v9ea470;
assign v84554a = hlock0_p & v845542 | !hlock0_p & !v845542;
assign bd5863 = hgrant0_p & bd5838 | !hgrant0_p & !bd574e;
assign d357a3 = hmaster2_p & d357a2 | !hmaster2_p & v845542;
assign v8cc61e = hlock3 & v8cc4ad | !hlock3 & v8cc4ac;
assign d357af = hlock2_p & d357ad | !hlock2_p & d357ae;
assign c3d6d6 = hmaster1_p & c3d6d5 | !hmaster1_p & c3d68b;
assign b578fe = hbusreq4_p & b578fd | !hbusreq4_p & v845542;
assign b5740c = hlock4 & b578f1 | !hlock4 & b5740b;
assign v8ccb89 = hmaster0_p & v8ccb75 | !hmaster0_p & v8d29fa;
assign d35a00 = hbusreq4_p & d359f1 | !hbusreq4_p & d359ff;
assign b579e7 = hlock2 & b579e5 | !hlock2 & b579e6;
assign d359f3 = stateG10_4_p & d359ce | !stateG10_4_p & d359f2;
assign v9f77b6 = hmaster0_p & v9f7790 | !hmaster0_p & v9f77b5;
assign ad4dd7 = hmaster1_p & ad4dc1 | !hmaster1_p & ad4dd6;
assign d35bea = hbusreq4_p & d35be9 | !hbusreq4_p & !v845542;
assign v9f787b = hmaster0_p & v9f7730 | !hmaster0_p & v9f772d;
assign v9f769b = hgrant4_p & v9f7ca6 | !hgrant4_p & v9ea445;
assign bd585f = stateG10_4_p & bd574e | !stateG10_4_p & !bd585e;
assign v9f7834 = hlock1 & v9f782f | !hlock1 & v9f7833;
assign v9ea4c1 = hbusreq2_p & v9ea4be | !hbusreq2_p & v9ea4c0;
assign d35721 = hgrant2_p & d3571a | !hgrant2_p & !d35720;
assign df51cd = hgrant3_p & df51b9 | !hgrant3_p & df51cc;
assign df5078 = hbusreq1 & dc5317 | !hbusreq1 & dc531a;
assign d359e7 = hbusreq0_p & v845542 | !hbusreq0_p & adeca0;
assign c5c8f8 = hgrant1_p & c5c8f7 | !hgrant1_p & c5c8f4;
assign df518e = hbusreq1_p & df518d | !hbusreq1_p & !v845542;
assign ad4344 = hbusreq1_p & ad4343 | !hbusreq1_p & c3d2d9;
assign ad476d = hmaster0_p & ad45ff | !hmaster0_p & ad476c;
assign d3575e = hready_p & d358e8 | !hready_p & d3575d;
assign c3d356 = hmaster1_p & c3d352 | !hmaster1_p & c3d355;
assign c3d3a7 = hmaster1_p & c3d3a5 | !hmaster1_p & c3d3a6;
assign c5c8e2 = stateG2_p & v845542 | !stateG2_p & v845568;
assign b1c7f8 = hgrant2_p & b1c7f1 | !hgrant2_p & b1c7f7;
assign adeab7 = hready_p & adeab5 | !hready_p & adeab6;
assign b05953 = hgrant0_p & b058b6 | !hgrant0_p & v9f7d42;
assign b57945 = decide_p & b57940 | !decide_p & b57944;
assign ad41b0 = hmaster0_p & ad41af | !hmaster0_p & bd5761;
assign ad4df5 = hbusreq2 & v845542 | !hbusreq2 & v845555;
assign bd579c = hbusreq1 & bd579a | !hbusreq1 & bd579b;
assign b579ee = hlock2 & b57942 | !hlock2 & b579ed;
assign v9f7800 = hmaster1_p & v9f77ff | !hmaster1_p & v9f77f4;
assign b1c5ea = hgrant4_p & v845542 | !hgrant4_p & b1c5e9;
assign v9f77ee = hlock0_p & v9f77eb | !hlock0_p & !v9f77ed;
assign b1cff9 = hlock0_p & b1cff8 | !hlock0_p & v845542;
assign ad4480 = hbusreq0_p & c3d318 | !hbusreq0_p & v845542;
assign ad4eb9 = hgrant4_p & ad4e54 | !hgrant4_p & v845542;
assign b1c08f = decide_p & b1c04a | !decide_p & !b1d013;
assign v8cc122 = hgrant3_p & v8ccbdc | !hgrant3_p & v8cc121;
assign v9f7cb8 = hlock0 & v9f7cb7 | !hlock0 & v9f7cb5;
assign c3d395 = hbusreq3 & c3d306 | !hbusreq3 & c3d32f;
assign b8f745 = hgrant3_p & b8f6e0 | !hgrant3_p & b8f744;
assign b1c82c = hbusreq2_p & v845542 | !hbusreq2_p & b1d01a;
assign ad442e = hmaster2_p & ad442b | !hmaster2_p & ad442d;
assign v8cc7f4 = hgrant0_p & v8cc7dd | !hgrant0_p & v845542;
assign bd5800 = hgrant4_p & c3d669 | !hgrant4_p & bd57fe;
assign b1c702 = hgrant3_p & b1c6e0 | !hgrant3_p & b1c701;
assign ad4eb2 = hbusreq1_p & ad4ead | !hbusreq1_p & !ad4eb1;
assign d359e2 = hbusreq1_p & d359aa | !hbusreq1_p & d359e1;
assign ad427b = hmaster1_p & ad4274 | !hmaster1_p & ad427a;
assign df5154 = hbusreq2_p & df514e | !hbusreq2_p & df5153;
assign v9f7e41 = hbusreq0 & v9f7e3b | !hbusreq0 & v9f7e40;
assign ade57f = hbusreq1 & ade4ac | !hbusreq1 & ade4ad;
assign b579ba = locked_p & b579b9 | !locked_p & v845542;
assign ad4f02 = hgrant4_p & v845542 | !hgrant4_p & !ad4f00;
assign c3ce06 = hmaster0_p & c3ce03 | !hmaster0_p & c3d5cf;
assign b05a31 = hbusreq2_p & b05a2e | !hbusreq2_p & b05a30;
assign c3ce1d = hmaster0_p & c3ce1b | !hmaster0_p & c3ce1c;
assign v9f77fe = hbusreq2 & v9f77fc | !hbusreq2 & v9f77fd;
assign b0598c = hgrant0_p & b058e9 | !hgrant0_p & v9ea3e9;
assign ad4fcb = hmaster2_p & v84556c | !hmaster2_p & !ad4fca;
assign v9ea60b = hlock3 & v9ea486 | !hlock3 & v9ea485;
assign ad4431 = hbusreq4 & ad442f | !hbusreq4 & ad4430;
assign ad4f86 = hgrant4_p & ad4f39 | !hgrant4_p & v845542;
assign c3d6be = hbusreq1_p & c3d6b1 | !hbusreq1_p & c3d6bd;
assign v9f7702 = hbusreq1_p & v9f7d97 | !hbusreq1_p & v9f76f9;
assign b579d5 = hbusreq0 & b579d4 | !hbusreq0 & b579ce;
assign adeaa5 = hbusreq4_p & v845576 | !hbusreq4_p & !adeaa4;
assign bd58b3 = hgrant1_p & bd58b1 | !hgrant1_p & bd58b2;
assign d356d5 = hbusreq1 & d358f0 | !hbusreq1 & v845542;
assign d357c8 = hgrant4_p & v84554a | !hgrant4_p & d3576e;
assign v8cc7a7 = hlock3_p & v8cc7a6 | !hlock3_p & v845542;
assign dc5385 = decide_p & dc531e | !decide_p & v845542;
assign c3cef1 = hbusreq4_p & c3ceef | !hbusreq4_p & c3cef0;
assign ad4f35 = stateA1_p & v845542 | !stateA1_p & ad4f34;
assign df5168 = hbusreq1_p & df5167 | !hbusreq1_p & v845542;
assign c5c8a6 = hmaster1_p & c5c8a5 | !hmaster1_p & c5c89f;
assign ad4ec2 = hbusreq4 & ad4ebe | !hbusreq4 & ad4ec1;
assign b058d1 = hmaster2_p & b058ce | !hmaster2_p & b058d0;
assign c5bed6 = jx2_p & c5c3bf | !jx2_p & c5c3be;
assign v9f7e29 = hlock3 & v9f7e28 | !hlock3 & v9f7e27;
assign v9f7703 = hgrant1_p & v9f7dab | !hgrant1_p & v9f7702;
assign df50d5 = hgrant3_p & df507e | !hgrant3_p & df50d4;
assign b57507 = hready_p & b57a2e | !hready_p & b57506;
assign v9ea445 = hgrant0_p & v9ea3fb | !hgrant0_p & v9ea3ec;
assign v9f782d = hbusreq4_p & v9f782b | !hbusreq4_p & v9f782c;
assign v8ccb83 = hmaster0_p & v8d29fa | !hmaster0_p & v8ccb75;
assign b1c6ba = hbusreq1_p & b1c6b9 | !hbusreq1_p & b1c850;
assign bd5766 = hlock2_p & bd575c | !hlock2_p & bd5765;
assign ade546 = hmaster1_p & ade542 | !hmaster1_p & ade545;
assign v9f7cd2 = hlock3 & v9f7cd1 | !hlock3 & v9f7cd0;
assign ad5013 = hbusreq3 & ad5012 | !hbusreq3 & v845547;
assign bd58bf = hgrant4_p & v845542 | !hgrant4_p & !bd58bd;
assign v9f7d8a = hlock0_p & v9f7d89 | !hlock0_p & v9ea3ec;
assign v9ea44d = locked_p & v9ea44c | !locked_p & v9ea3ec;
assign ade4e2 = hbusreq4_p & ade4e1 | !hbusreq4_p & v845542;
assign b579ca = stateG10_4_p & v845542 | !stateG10_4_p & b579c9;
assign v9f784e = hbusreq2 & v9f784c | !hbusreq2 & v9f784d;
assign dc4fa9 = hlock0_p & ade4cc | !hlock0_p & v845542;
assign v9f7883 = hgrant4_p & v9f772b | !hgrant4_p & v9f7882;
assign d354d1 = hbusreq0 & d354cd | !hbusreq0 & d354d0;
assign df50dd = decide_p & df50dc | !decide_p & v845542;
assign v857467 = hbusreq2_p & v882b8e | !hbusreq2_p & !v845542;
assign v9f7dec = hready & v9f7deb | !hready & v9f7de7;
assign d356ae = hbusreq3 & d356ab | !hbusreq3 & d356ad;
assign v9f785a = hlock2_p & v9f7857 | !hlock2_p & v9f7859;
assign v8cc816 = hbusreq2_p & v8cc80b | !hbusreq2_p & v8cc815;
assign v9f77d3 = hlock2 & v9f77d0 | !hlock2 & v9f77d2;
assign b573db = hbusreq3 & b573d9 | !hbusreq3 & b573da;
assign ad448b = hbusreq0 & ad448a | !hbusreq0 & v845542;
assign c3ceb2 = hbusreq2 & c3ceae | !hbusreq2 & c3ceb0;
assign d35a0a = hbusreq0 & d359fd | !hbusreq0 & d35a09;
assign ad446d = hmaster1_p & ad446c | !hmaster1_p & ad481c;
assign c3ce31 = hbusreq3_p & c3ce25 | !hbusreq3_p & c3ce30;
assign b1c724 = hbusreq3 & b1c723 | !hbusreq3 & b1c71d;
assign c5c972 = hmaster2_p & c5c971 | !hmaster2_p & !v845542;
assign bd56d7 = hbusreq4_p & d3594e | !hbusreq4_p & !v845542;
assign v8da59e = hready_p & v845542 | !hready_p & !v845564;
assign ad456d = hmaster2_p & ad4554 | !hmaster2_p & v845542;
assign c3d327 = hbusreq4_p & c3d2fd | !hbusreq4_p & c3d326;
assign v9f7d7f = hmaster2_p & v9f7d77 | !hmaster2_p & !v9f7d7e;
assign d3501f = hmaster1_p & d35015 | !hmaster1_p & d3501e;
assign v9ea59f = hbusreq0 & v9ea59e | !hbusreq0 & v9ea59b;
assign v9f7caa = hlock4 & v9f7ca7 | !hlock4 & v9f7ca9;
assign ad4f99 = hbusreq0 & ad4f93 | !hbusreq0 & ad4f98;
assign c3ce22 = hbusreq2_p & c3ce21 | !hbusreq2_p & c3d36c;
assign v8ccb78 = hbusreq1_p & v8ccb76 | !hbusreq1_p & v8ccb75;
assign b578f7 = hburst0_p & v9ea411 | !hburst0_p & !b578f6;
assign ade652 = jx1_p & ade629 | !jx1_p & ade651;
assign ad3cc1 = hmaster0_p & ad4488 | !hmaster0_p & ad3cc0;
assign ad4fee = hmaster0_p & ad4fd4 | !hmaster0_p & ad4fed;
assign v9f789d = hmaster1_p & v9f7878 | !hmaster1_p & v9f7811;
assign d35a25 = hmaster0_p & d35a23 | !hmaster0_p & !d35a24;
assign df54e2 = hmaster2_p & v845542 | !hmaster2_p & df54e1;
assign bd589d = hmastlock_p & bd589c | !hmastlock_p & !v845542;
assign dc4fd6 = hbusreq3 & dc4fd5 | !hbusreq3 & v845542;
assign ad432b = hmaster0_p & ad42d3 | !hmaster0_p & ad42d1;
assign v9e9fc1 = hmaster1_p & v9e9fc0 | !hmaster1_p & v9e9ef1;
assign d35bfd = hmaster0_p & d35bec | !hmaster0_p & d35bfc;
assign v9f7865 = hbusreq1_p & v9f7760 | !hbusreq1_p & v9f7864;
assign b1c71a = hbusreq0_p & adec89 | !hbusreq0_p & v845542;
assign v9f7e00 = hlock2 & v9f7da3 | !hlock2 & v9f7dff;
assign v9f7765 = hbusreq3 & v9f7761 | !hbusreq3 & v9f7764;
assign ac1488 = stateG10_4_p & ac1486 | !stateG10_4_p & ac1487;
assign c3d57b = hbusreq4_p & v8da59f | !hbusreq4_p & c3d39f;
assign v9ea4b1 = hmaster1_p & v9ea4a7 | !hmaster1_p & v9ea4af;
assign c3ced8 = decide_p & c3ceb8 | !decide_p & !c3cea8;
assign v9f7e20 = hlock0 & v9f7e1f | !hlock0 & v9f7e18;
assign ad3d50 = hbusreq3 & ad3d18 | !hbusreq3 & ad3d19;
assign dc5071 = hbusreq1_p & c3d66d | !hbusreq1_p & dc5070;
assign c3d5bb = hmaster2_p & c3d5ba | !hmaster2_p & v8da5a1;
assign c3d6d4 = hgrant2_p & c3d6a3 | !hgrant2_p & c3d6d3;
assign v8cc7e6 = hbusreq1 & v8cc7e4 | !hbusreq1 & v8cc7e5;
assign b1c5e6 = hgrant4_p & v845542 | !hgrant4_p & !b1c5e5;
assign ad428a = hmaster1_p & ad4285 | !hmaster1_p & ad4289;
assign ad45a4 = hready & ad457c | !hready & ad45a3;
assign d359f8 = hgrant4_p & d3598a | !hgrant4_p & d359f7;
assign c3d4f0 = hbusreq4_p & v8da59f | !hbusreq4_p & v845576;
assign d35a5f = hgrant4_p & v845542 | !hgrant4_p & !d35a5d;
assign v9f7852 = hbusreq2_p & v9f7848 | !hbusreq2_p & v9f7851;
assign b1c0a7 = hgrant1_p & b1d01a | !hgrant1_p & b1c0a6;
assign df51e0 = jx2_p & df5136 | !jx2_p & df51df;
assign df51dd = hgrant3_p & df51d5 | !hgrant3_p & df51dc;
assign df51a6 = hmaster0_p & df51a4 | !hmaster0_p & df51a5;
assign ad458b = hready & ad458a | !hready & v845542;
assign b574c9 = hbusreq1 & b574c7 | !hbusreq1 & b574c8;
assign d3565b = hmaster1_p & d35645 | !hmaster1_p & d3565a;
assign d357b0 = hbusreq2_p & d357af | !hbusreq2_p & d357ae;
assign ade4dc = hbusreq1 & ade4d6 | !hbusreq1 & ade4db;
assign dc503d = hgrant4_p & ade4aa | !hgrant4_p & ade58d;
assign c3d5c7 = hbusreq0 & c3d5b6 | !hbusreq0 & c3d5c6;
assign c5c8fa = hlock4_p & c5c8f9 | !hlock4_p & !v845542;
assign b1c5fd = decide_p & b1c5fc | !decide_p & v845542;
assign ad4f17 = hmaster1_p & ad4eaa | !hmaster1_p & ad4f16;
assign b1cb00 = hready_p & v845542 | !hready_p & b1caff;
assign c5c940 = hmaster1_p & c5c93f | !hmaster1_p & v845542;
assign v9ea4b7 = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea4b6;
assign ad47ff = hmaster1_p & ad4720 | !hmaster1_p & ad471b;
assign ad4738 = hmaster2_p & adec93 | !hmaster2_p & !ad4737;
assign d3560e = hmaster2_p & dc5318 | !hmaster2_p & !d3590d;
assign b1c02d = hlock2_p & b1c827 | !hlock2_p & b1c829;
assign d3542e = hbusreq4 & d3542c | !hbusreq4 & d3542d;
assign bd5782 = stateG2_p & v889629 | !stateG2_p & v845542;
assign ad45fe = hbusreq2_p & ad45fd | !hbusreq2_p & ad45fc;
assign ad45b4 = hmaster2_p & v845542 | !hmaster2_p & !ad45b3;
assign df552d = hgrant3_p & df54f0 | !hgrant3_p & df552c;
assign ad4695 = hmaster2_p & ad4694 | !hmaster2_p & v845542;
assign c3d4f4 = hbusreq4_p & v8da59f | !hbusreq4_p & !adeaa4;
assign d3541b = hbusreq4_p & d3541a | !hbusreq4_p & v845542;
assign ad4260 = hgrant3_p & ad41b9 | !hgrant3_p & ad425f;
assign d359a0 = hlock4_p & d3599e | !hlock4_p & !d3599f;
assign ad46c0 = hbusreq4 & ad46bf | !hbusreq4 & ad46ac;
assign ad4f16 = hmaster0_p & ad4ec9 | !hmaster0_p & ad4f15;
assign d354a3 = hlock4_p & d359a5 | !hlock4_p & !d35a45;
assign ad3cde = hlock0_p & ad502f | !hlock0_p & ad3cdd;
assign ad440c = hmaster2_p & b1c714 | !hmaster2_p & ad440b;
assign v9ea620 = hbusreq1 & v9ea453 | !hbusreq1 & v9ea454;
assign cc36eb = hgrant2_p & cc36d9 | !hgrant2_p & cc36ea;
assign ad441f = hready_p & ad43bf | !hready_p & ad441e;
assign v9ea450 = hbusreq0 & v9ea44e | !hbusreq0 & v9ea44f;
assign v9ea4c5 = hmaster1_p & v9ea4c4 | !hmaster1_p & v9ea4bd;
assign c5c88f = hmaster2_p & v845542 | !hmaster2_p & !c5c88e;
assign v9f77c3 = locked_p & v9f772a | !locked_p & v9f772b;
assign ad46e0 = hbusreq0 & ad46d9 | !hbusreq0 & ad46df;
assign df54d7 = hbusreq1 & dc5394 | !hbusreq1 & df54d6;
assign v9f7898 = hbusreq2 & v9f7896 | !hbusreq2 & v9f7897;
assign b1c4ce = hbusreq1_p & b1c4a7 | !hbusreq1_p & b1c4cd;
assign v9ea4b4 = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea4b3;
assign v9e9fd5 = hbusreq2_p & v9e9fd2 | !hbusreq2_p & v9e9fd4;
assign dc501a = hmaster2_p & v845542 | !hmaster2_p & ade572;
assign b1c747 = hbusreq3 & b1c73e | !hbusreq3 & !v845542;
assign v9f7711 = hmaster0_p & v9f7cee | !hmaster0_p & v9f767b;
assign b1c80e = hbusreq3 & b1c80d | !hbusreq3 & !b1c80a;
assign c3ce53 = hgrant1_p & v84554d | !hgrant1_p & c3ce52;
assign v9f7ce6 = hbusreq3 & v9f7ce4 | !hbusreq3 & v9f7ce5;
assign ad45c6 = hready & ad45c5 | !hready & !v845542;
assign ade580 = hbusreq0_p & c3d66d | !hbusreq0_p & !adeca0;
assign c3d34a = hmaster2_p & c3d33e | !hmaster2_p & v8da5a1;
assign c3d2b7 = hbusreq3 & c3d2b6 | !hbusreq3 & !v845542;
assign ad4379 = hgrant3_p & ad435b | !hgrant3_p & !ad4378;
assign ba7c73 = hgrant2_p & v845558 | !hgrant2_p & ba7c6b;
assign ad4ec8 = hgrant1_p & ad4eb2 | !hgrant1_p & ad4ec7;
assign ad4e87 = hmaster2_p & ad4e86 | !hmaster2_p & v845542;
assign ad4dc2 = stateG2_p & v845542 | !stateG2_p & ade5ca;
assign ade4cf = hbusreq3 & ade4c7 | !hbusreq3 & ade4ce;
assign ad4e20 = hlock3_p & ad4ddb | !hlock3_p & !ad4e1f;
assign d35572 = hmaster0_p & d35570 | !hmaster0_p & d35571;
assign ad4d93 = hready & ad4d92 | !hready & !v845564;
assign v9ea4de = hmaster0_p & v9ea4b7 | !hmaster0_p & v9ea4b4;
assign v9f778e = hbusreq3 & v9f778c | !hbusreq3 & v9f778d;
assign b0589f = jx0_p & v85746a | !jx0_p & !b0589e;
assign c3ce3f = hmaster0_p & c3ce3e | !hmaster0_p & c3d2be;
assign c3d330 = hbusreq3 & c3d32c | !hbusreq3 & c3d32f;
assign ad4808 = hmaster2_p & v845542 | !hmaster2_p & !d35a4e;
assign dc52fe = hmastlock_p & v8ccb67 | !hmastlock_p & !v845542;
assign b1c827 = hmaster1_p & b1c826 | !hmaster1_p & b1c775;
assign b1c73e = hbusreq0 & b1c73d | !hbusreq0 & v845542;
assign ad471e = hmaster0_p & ad459e | !hmaster0_p & ad470d;
assign bd5774 = hmaster0_p & bd576e | !hmaster0_p & bd5773;
assign v9f777b = hmaster1_p & v9f777a | !hmaster1_p & v9f776d;
assign ad413e = hgrant4_p & adea99 | !hgrant4_p & v845542;
assign v9f7dc3 = hbusreq3 & v9f7dbd | !hbusreq3 & v9f7dc2;
assign ad5012 = hready & dc4fcb | !hready & !v845542;
assign d359d5 = hgrant4_p & d35983 | !hgrant4_p & v845542;
assign bd578d = stateA1_p & d3561b | !stateA1_p & !d3594a;
assign ade581 = hlock0_p & c3d66d | !hlock0_p & ade580;
assign cc36e6 = hbusreq4_p & cc36e4 | !hbusreq4_p & !cc36e5;
assign c3ce9c = hready & c3ce9b | !hready & !v845542;
assign b1c700 = decide_p & b1c6de | !decide_p & b1d013;
assign cc36cf = hmaster0_p & cc36c7 | !hmaster0_p & cc36ce;
assign stateA1 = !c3d763;
assign ad4598 = hbusreq4_p & ad4fae | !hbusreq4_p & v845542;
assign b1caff = decide_p & b1cafe | !decide_p & v845542;
assign b57ac3 = hbusreq4 & b57ac1 | !hbusreq4 & b57ac2;
assign d354c0 = hlock4_p & d359dc | !hlock4_p & !dc500f;
assign ade568 = hbusreq0 & ade55e | !hbusreq0 & ade567;
assign b57a87 = hlock2 & b57942 | !hlock2 & b57a86;
assign v9ea42e = stateG10_4_p & v845542 | !stateG10_4_p & v9ea418;
assign c3d750 = hmaster0_p & c3d676 | !hmaster0_p & c3d6e9;
assign v9ea5d4 = hbusreq3 & v9ea5d3 | !hbusreq3 & v9ea5cb;
assign v9ea49f = decide_p & v9ea3f9 | !decide_p & v9ea49e;
assign dc53a1 = hmaster0_p & dc53a0 | !hmaster0_p & v845542;
assign b058f8 = hbusreq0 & b058c7 | !hbusreq0 & b058f7;
assign ad4421 = hbusreq2 & ad4385 | !hbusreq2 & ad438b;
assign dc4fa2 = hbusreq1 & dc4f9e | !hbusreq1 & dc4f6a;
assign cc36f4 = hbusreq4_p & d35a48 | !hbusreq4_p & !cc36f3;
assign c3d590 = hmaster2_p & c3d2ad | !hmaster2_p & !v845542;
assign v8cc7db = stateA1_p & v8cc7da | !stateA1_p & v8ccb67;
assign bd5856 = hgrant1_p & bd583b | !hgrant1_p & bd5855;
assign v8cc492 = hgrant0_p & v8d2b2b | !hgrant0_p & v845542;
assign dc4fb9 = hlock0_p & ade5ce | !hlock0_p & v845542;
assign b059ea = hlock4 & b059e7 | !hlock4 & b059e9;
assign d3577d = hmaster1_p & d35779 | !hmaster1_p & d3577c;
assign v9ea43d = hmaster2_p & v9ea439 | !hmaster2_p & v9ea3fe;
assign bd572c = hbusreq3_p & bd56cd | !hbusreq3_p & bd5728;
assign ad4f8e = hbusreq0 & ad4f85 | !hbusreq0 & ad4f8d;
assign b1c6c9 = hmaster0_p & b1d00e | !hmaster0_p & b1c6c8;
assign v9e9e70 = hgrant3_p & v9ea628 | !hgrant3_p & v9e9e6f;
assign bd57f8 = busreq_p & v889629 | !busreq_p & bd57f7;
assign ad47f3 = hmaster0_p & ad47ee | !hmaster0_p & ad46f0;
assign v9f7793 = hbusreq0 & v9f7791 | !hbusreq0 & v9f7792;
assign b05a58 = stateG2_p & v845542 | !stateG2_p & !v9fa31b;
assign ad4591 = hmaster0_p & ad458d | !hmaster0_p & !ad4590;
assign b05a37 = decide_p & b05a31 | !decide_p & b05a36;
assign ad44b4 = hmaster2_p & ad44b3 | !hmaster2_p & v845542;
assign ad445a = hbusreq0 & ad4459 | !hbusreq0 & v845542;
assign ad4586 = hready & ad4585 | !hready & v845542;
assign v9e9fb7 = hlock2 & v9e9f68 | !hlock2 & v9e9fb6;
assign ad433f = hgrant1_p & v845542 | !hgrant1_p & ad433e;
assign d359ab = hgrant1_p & d35994 | !hgrant1_p & d359aa;
assign c3d300 = hbusreq4 & c3d2fc | !hbusreq4 & !c3d2ff;
assign v9f7807 = hlock2 & v9f7804 | !hlock2 & v9f7806;
assign bd5799 = hbusreq1 & bd5787 | !hbusreq1 & bd578c;
assign v9e9ec5 = hmaster0_p & v9e9ec4 | !hmaster0_p & v9ea3fc;
assign bd5e21 = hmaster1_p & bd5e20 | !hmaster1_p & v845542;
assign v9f7823 = hlock1 & v9f77c8 | !hlock1 & v9f7822;
assign v9f7cde = hlock0 & v9f7cdd | !hlock0 & v9f7cd9;
assign bd5896 = hgrant1_p & bd585a | !hgrant1_p & bd5895;
assign c3d681 = locked_p & c3d66b | !locked_p & c3d66d;
assign b57535 = hbusreq3_p & b57534 | !hbusreq3_p & b57a34;
assign v9f7d54 = hmaster1_p & v9f7d53 | !hmaster1_p & v9f7d47;
assign v9e9f7e = hlock1 & v9e9f79 | !hlock1 & v9e9f7d;
assign c5c99c = hready_p & c5c953 | !hready_p & !c5c99b;
assign d35a2f = hlock1_p & d35a2d | !hlock1_p & !d35a2e;
assign ade599 = hgrant0_p & ade598 | !hgrant0_p & !v84556c;
assign ac1484 = hready_p & ac1483 | !hready_p & !v845542;
assign b579c3 = hbusreq1_p & b57942 | !hbusreq1_p & b579c2;
assign ade4b2 = hmaster0_p & adec9d | !hmaster0_p & ade4b1;
assign ad46f6 = hgrant1_p & ad46f5 | !hgrant1_p & ad46c1;
assign cc36d0 = hmaster1_p & cc36c4 | !hmaster1_p & cc36cf;
assign bd58ae = hbusreq0 & bd58ac | !hbusreq0 & bd58ad;
assign b1c756 = hbusreq0_p & ade4c5 | !hbusreq0_p & v845542;
assign df51ac = hbusreq1_p & df51ab | !hbusreq1_p & v845542;
assign ade575 = hbusreq1 & ade56f | !hbusreq1 & !ade574;
assign ad41b7 = hbusreq2_p & ad41b6 | !hbusreq2_p & ad508e;
assign b57953 = hlock0_p & b57952 | !hlock0_p & v845542;
assign v9f7e13 = stateG10_4_p & v9f7d70 | !stateG10_4_p & v9f7e12;
assign b059cf = hgrant1_p & b059ce | !hgrant1_p & b05970;
assign c3d75b = hmaster0_p & c3d699 | !hmaster0_p & c3d685;
assign df54dc = stateG2_p & v845542 | !stateG2_p & dc539d;
assign b5741b = hbusreq0_p & b57952 | !hbusreq0_p & b5741a;
assign b05912 = hbusreq2 & b05910 | !hbusreq2 & b05911;
assign ad4604 = hlock2_p & ad4601 | !hlock2_p & ad4603;
assign v9e9e6b = hmaster1_p & v9e9e6a | !hmaster1_p & v9ea60e;
assign v9f7d8f = hbusreq4_p & v9f7d8d | !hbusreq4_p & v9f7d8e;
assign b0590f = hlock3 & b058d5 | !hlock3 & b0590e;
assign ade659 = hbusreq1_p & adea9e | !hbusreq1_p & adea94;
assign dc4fca = hbusreq3 & dc4fc9 | !hbusreq3 & v845542;
assign b1cfbe = stateG10_4_p & b1cfb6 | !stateG10_4_p & !b1cfb7;
assign b1c07e = stateG10_4_p & b1c066 | !stateG10_4_p & b1c07d;
assign dc5059 = hmaster2_p & dc5054 | !hmaster2_p & dc5058;
assign b0599b = hgrant1_p & b058d5 | !hgrant1_p & !b05992;
assign c3d6e1 = hgrant4_p & c3d66a | !hgrant4_p & c3d6a5;
assign adea9f = hgrant1_p & v845542 | !hgrant1_p & !adea9e;
assign dc5030 = hbusreq3 & dc502f | !hbusreq3 & v845542;
assign c3d5cc = hgrant1_p & v84554d | !hgrant1_p & c3d5cb;
assign b1d013 = hgrant2_p & v845542 | !hgrant2_p & b1d012;
assign ad4132 = hlock4_p & ad4131 | !hlock4_p & !ad4e9a;
assign b05a97 = hbusreq2_p & b05a92 | !hbusreq2_p & b05a96;
assign ad4f83 = stateG10_4_p & ad4f80 | !stateG10_4_p & !ad4f82;
assign bd592d = hready_p & v845542 | !hready_p & bd592c;
assign b058e2 = hmaster1_p & b058c6 | !hmaster1_p & b058e1;
assign v9e9e75 = hbusreq2_p & v9e9e74 | !hbusreq2_p & v9ea5f4;
assign bbbcd9 = hburst1_p & bbbcd8 | !hburst1_p & v845542;
assign df5126 = hbusreq1_p & df5125 | !hbusreq1_p & !v845542;
assign d354d8 = hmaster0_p & d354d6 | !hmaster0_p & d354d7;
assign v8ccbde = hmaster1_p & v8ccbdd | !hmaster1_p & v845542;
assign b5b409 = hgrant0_p & v845542 | !hgrant0_p & b5b408;
assign v9f7d25 = hbusreq0 & v9f7c9f | !hbusreq0 & !v9f7d24;
assign ade4d6 = hmaster2_p & ade4c0 | !hmaster2_p & !ade4d5;
assign v9f7db5 = hlock0 & v9f7db4 | !hlock0 & v9f7dac;
assign v9f7cf8 = hmaster2_p & v9f7ca4 | !hmaster2_p & !v9f7cf7;
assign v9f786e = hbusreq3 & v9f786b | !hbusreq3 & v9f786d;
assign ad4e5e = hready & ad4e5d | !hready & v84556c;
assign c5c97c = hmaster1_p & c5c97b | !hmaster1_p & c5c96c;
assign b57449 = decide_p & b57a21 | !decide_p & b57448;
assign v8cc619 = hlock3 & v8cc489 | !hlock3 & v8cc488;
assign c3cf33 = jx0_p & c3cedc | !jx0_p & c3cf32;
assign bd58c1 = hbusreq4_p & bd58be | !hbusreq4_p & bd58c0;
assign bd56d1 = hburst0 & bd5b6a | !hburst0 & bd56d0;
assign b05a3e = hlock0_p & b0591c | !hlock0_p & b05a3d;
assign v9f7d2b = hlock3 & v9f7d23 | !hlock3 & !v9f7d2a;
assign ad4718 = hbusreq4 & ad4717 | !hbusreq4 & v845542;
assign bd5792 = hbusreq1_p & bd578c | !hbusreq1_p & bd5791;
assign v9ea453 = hready & v9ea452 | !hready & v9ea3fa;
assign b1caf5 = hmaster2_p & v845542 | !hmaster2_p & !b1caf4;
assign v9ea4a2 = hmaster0_p & v9ea415 | !hmaster0_p & v845542;
assign df5140 = hbusreq1 & adec89 | !hbusreq1 & v845542;
assign c3d322 = hmaster2_p & c3d321 | !hmaster2_p & c3d30d;
assign v9f7d91 = hlock0 & v9f7d90 | !hlock0 & v9f7d7f;
assign bd5b7a = hlock2_p & bd5b79 | !hlock2_p & v845542;
assign ad455a = hmaster2_p & adec93 | !hmaster2_p & ad4559;
assign v9ea614 = hmaster1_p & v9ea613 | !hmaster1_p & v9ea4db;
assign ad484a = hbusreq3 & ad4d98 | !hbusreq3 & ad4849;
assign ade560 = hlock4_p & ade55f | !hlock4_p & !ade557;
assign b059a8 = hmaster1_p & b059a7 | !hmaster1_p & b05913;
assign df54f7 = hbusreq1 & df54f5 | !hbusreq1 & df54f6;
assign v8cc627 = decide_p & v8ccbd7 | !decide_p & v8cc626;
assign d357b9 = hlock0_p & v845542 | !hlock0_p & !dc538c;
assign v9f76c2 = hlock2_p & v9f76bf | !hlock2_p & v9f76c1;
assign ad4165 = hbusreq2_p & ad4164 | !hbusreq2_p & v845542;
assign ade65d = hgrant2_p & v845542 | !hgrant2_p & ade65c;
assign b1c750 = stateG2_p & v889629 | !stateG2_p & bb9bdd;
assign c3d4dc = hbusreq4_p & c3d4db | !hbusreq4_p & v845542;
assign ad434c = hbusreq3 & ad4304 | !hbusreq3 & !ad4282;
assign d3569b = hbusreq3_p & d35688 | !hbusreq3_p & d3569a;
assign cc36be = hmaster2_p & v845566 | !hmaster2_p & !cc36bd;
assign bd5823 = hbusreq4 & bd5813 | !hbusreq4 & bd5822;
assign b57434 = hgrant2_p & b57433 | !hgrant2_p & b5742c;
assign b058ac = hbusreq0 & b058a8 | !hbusreq0 & b058ab;
assign dc539f = hmaster2_p & v845542 | !hmaster2_p & dc539e;
assign c3ced1 = hbusreq1_p & c3d300 | !hbusreq1_p & c3ced0;
assign bd58ed = decide_p & bd58ec | !decide_p & v845542;
assign d359ec = hbusreq1_p & d359eb | !hbusreq1_p & d359ea;
assign v9ea4da = hgrant1_p & v9ea4bc | !hgrant1_p & v9ea4d9;
assign df51be = hmaster1_p & df51bd | !hmaster1_p & df5185;
assign c3d507 = hmaster1_p & c3d4f8 | !hmaster1_p & c3d506;
assign bd584d = hmaster2_p & bd5817 | !hmaster2_p & bd584c;
assign d357a2 = hbusreq4_p & d357a1 | !hbusreq4_p & v84554a;
assign bbbe36 = hburst0_p & v845542 | !hburst0_p & bbbe35;
assign cc36df = hgrant1_p & cc36be | !hgrant1_p & cc36de;
assign c3d308 = hgrant4_p & v845542 | !hgrant4_p & !ade562;
assign b1c57d = hbusreq0 & b1c4c4 | !hbusreq0 & b1c57c;
assign bd5740 = hburst0 & d355a6 | !hburst0 & bd573f;
assign v8cc472 = hmaster1_p & v8cc470 | !hmaster1_p & v845542;
assign ad45e1 = hbusreq4 & ad45e0 | !hbusreq4 & v845542;
assign b1c751 = stateA1_p & bd57c0 | !stateA1_p & !b1c750;
assign c3ceca = hmaster2_p & c3cec9 | !hmaster2_p & v845576;
assign ad42a8 = hmaster0_p & ad42a6 | !hmaster0_p & ad42a7;
assign d3563b = hburst0 & ade54b | !hburst0 & d354ad;
assign d358fc = hlock1_p & d358fb | !hlock1_p & v845542;
assign b1c5f7 = hready_p & b1c5f5 | !hready_p & b1c5f6;
assign v8cc80a = hmaster1_p & v8ccbe5 | !hmaster1_p & v8cc809;
assign d357eb = hmaster2_p & v84554a | !hmaster2_p & !v845542;
assign ad4846 = hmaster2_p & v845542 | !hmaster2_p & d3561c;
assign dc5319 = hbusreq4_p & dc5318 | !hbusreq4_p & !v845542;
assign bd57eb = hmaster1_p & bd57ea | !hmaster1_p & bd57e1;
assign v9f7cec = hbusreq3 & v9f7ccf | !hbusreq3 & v9f7ceb;
assign b1c085 = hmaster2_p & b1c084 | !hmaster2_p & b1c858;
assign b05964 = hgrant1_p & b058b8 | !hgrant1_p & b0595b;
assign ad446a = hmaster1_p & ad4433 | !hmaster1_p & ad4469;
assign ad4100 = locked_p & ad4e6a | !locked_p & !v845542;
assign v9f76cb = hbusreq2_p & v9f76c2 | !hbusreq2_p & v9f76ca;
assign bd5750 = hbusreq1_p & bd574d | !hbusreq1_p & bd574f;
assign b1c05a = hmaster0_p & b1c058 | !hmaster0_p & b1c059;
assign d35655 = hlock4_p & d35653 | !hlock4_p & !d35654;
assign ad46dd = hlock4_p & ad46dc | !hlock4_p & v845542;
assign c3d32d = hbusreq0 & c3d325 | !hbusreq0 & v845542;
assign dc4ff5 = stateG10_4_p & ade557 | !stateG10_4_p & !dc4ff4;
assign v8ccb68 = stateG2_p & v845542 | !stateG2_p & v8ccb67;
assign d356f2 = hready_p & d356d1 | !hready_p & d356f1;
assign b574d3 = hlock3 & b57942 | !hlock3 & b574d2;
assign ad42a3 = hbusreq1 & ad4de3 | !hbusreq1 & !v845542;
assign ad480a = hbusreq3 & ad4807 | !hbusreq3 & ad4809;
assign c3d37c = hbusreq2 & c3d378 | !hbusreq2 & c3d37b;
assign bd58a6 = hgrant4_p & v84556c | !hgrant4_p & bd58a5;
assign ad4e58 = hbusreq3 & ad4e57 | !hbusreq3 & v845542;
assign d35a71 = hlock1_p & dc4fcb | !hlock1_p & !v845542;
assign ad4266 = hbusreq1 & ad4265 | !hbusreq1 & v845542;
assign v9ea56c = hmaster1_p & v9f20a1 | !hmaster1_p & v9ea56b;
assign ad4e56 = hready & ad4e55 | !hready & v84556c;
assign b1c744 = hbusreq3 & b1c743 | !hbusreq3 & !v845542;
assign c3cebc = hlock0_p & v845542 | !hlock0_p & c3cebb;
assign d35498 = hmaster2_p & d35be8 | !hmaster2_p & d35497;
assign bd57c2 = hmastlock_p & bd57c1 | !hmastlock_p & v845542;
assign bd593e = hready_p & bd593c | !hready_p & !bd593d;
assign bd58a9 = hbusreq4_p & bd58a6 | !hbusreq4_p & bd58a8;
assign c3d5d2 = hgrant2_p & v845551 | !hgrant2_p & c3d5d1;
assign v9f78af = jx1_p & v9f7728 | !jx1_p & v9f78ae;
assign d35627 = hlock0_p & dc539e | !hlock0_p & v845542;
assign bd5bad = hlock2_p & bd5bac | !hlock2_p & !v845542;
assign v9f77be = hgrant0_p & v9f772b | !hgrant0_p & v9f77bd;
assign ad41a2 = hbusreq2 & ad41a1 | !hbusreq2 & ad5024;
assign c3d315 = hgrant1_p & v84554d | !hgrant1_p & c3d314;
assign c3d5e7 = hmaster2_p & c3d327 | !hmaster2_p & v845542;
assign d35738 = hmaster0_p & d35736 | !hmaster0_p & d35737;
assign dc5011 = hbusreq4_p & dc500e | !hbusreq4_p & dc5010;
assign b1c773 = hbusreq0 & b1c772 | !hbusreq0 & b1cf2b;
assign b0592e = hmaster0_p & b0591e | !hmaster0_p & b0591d;
assign ad4d9e = hbusreq2 & ad4d99 | !hbusreq2 & ad4d9d;
assign b5794f = hgrant4_p & b5b408 | !hgrant4_p & v845542;
assign df51da = decide_p & df512a | !decide_p & d6ebca;
assign v9f767b = hbusreq2 & v9f7679 | !hbusreq2 & v9f767a;
assign d35731 = hbusreq3 & d35730 | !hbusreq3 & d35aa4;
assign ad473e = hbusreq1_p & ad460a | !hbusreq1_p & ad473d;
assign c5c978 = hmaster1_p & c5c973 | !hmaster1_p & c5c977;
assign v9f7d3c = hmaster2_p & v9f7d3a | !hmaster2_p & v9ea3ec;
assign d354f3 = hmaster2_p & d354f1 | !hmaster2_p & !d354f2;
assign bd56cf = hmastlock_p & bd56ce | !hmastlock_p & v845542;
assign v9f7844 = hmaster2_p & v9f7840 | !hmaster2_p & !v9f7843;
assign bd57b0 = hbusreq2 & bd57af | !hbusreq2 & v845542;
assign bd58d1 = hmaster2_p & bd58d0 | !hmaster2_p & bd58ca;
assign b1c763 = hmaster2_p & b1c755 | !hmaster2_p & ade4e6;
assign d357c5 = stateG10_4_p & d357c1 | !stateG10_4_p & d357c3;
assign bd5b80 = hburst0 & bd5b7f | !hburst0 & adea98;
assign ad3ccf = hready & ad3cce | !hready & !v845542;
assign v8cc624 = hmaster1_p & v8cc475 | !hmaster1_p & v8cc623;
assign bd5845 = stateG10_4_p & bd5842 | !stateG10_4_p & !bd5844;
assign b1c7a7 = hbusreq4_p & b1c7a4 | !hbusreq4_p & !b1c7a6;
assign d356b0 = hlock1_p & d35991 | !hlock1_p & dc4fcb;
assign bd5914 = hbusreq1 & bd5b89 | !hbusreq1 & v845542;
assign d35699 = hready_p & d35698 | !hready_p & d3568c;
assign ade64d = hbusreq2_p & adeaa2 | !hbusreq2_p & adeab4;
assign v9e9f8d = hbusreq4_p & v9ea462 | !hbusreq4_p & v9e9f8c;
assign v9f7751 = hmaster2_p & v9f772a | !hmaster2_p & !v845542;
assign v9f768f = hbusreq4_p & v9f768d | !hbusreq4_p & v9f768e;
assign d354fa = hbusreq3 & d354f9 | !hbusreq3 & !d354f5;
assign v8cc4ab = hbusreq1 & v8cc4a9 | !hbusreq1 & v8cc4aa;
assign d357f0 = hbusreq2_p & v84554a | !hbusreq2_p & d357ef;
assign ad4e94 = hbusreq1 & ad4e52 | !hbusreq1 & v845542;
assign v8ccbe7 = hbusreq1_p & v8ccbe6 | !hbusreq1_p & v845542;
assign c3d33f = hmaster2_p & c3d33e | !hmaster2_p & adeaa5;
assign ad41af = hbusreq2 & ad4fd0 | !hbusreq2 & v845542;
assign d35594 = hgrant2_p & d35576 | !hgrant2_p & !d35593;
assign c3d5e0 = hmaster2_p & c3d5df | !hmaster2_p & v845576;
assign v9f7654 = stateG10_4_p & v9f7d42 | !stateG10_4_p & !v9f7653;
assign d35579 = hbusreq4_p & d354a3 | !hbusreq4_p & !d35aab;
assign bd590a = hbusreq2 & dc53bf | !hbusreq2 & bd5909;
assign v9f7d10 = hbusreq2 & v9f7d0e | !hbusreq2 & v9f7d0f;
assign v9e9e9b = hgrant0_p & v9ea439 | !hgrant0_p & v9f20a1;
assign c5c92d = stateA1_p & v845542 | !stateA1_p & bb9bdd;
assign v9f7d82 = hgrant0_p & v9f7ca4 | !hgrant0_p & !v9f7d80;
assign v9f7718 = hmaster1_p & v9f7717 | !hmaster1_p & v9f7d64;
assign b0596f = hbusreq1_p & b0596e | !hbusreq1_p & b058e8;
assign adeca2 = hbusreq4_p & adeca1 | !hbusreq4_p & v845542;
assign b1c77f = hbusreq3 & b1c762 | !hbusreq3 & b1c764;
assign b05994 = hbusreq0 & b05986 | !hbusreq0 & b05993;
assign ad42e3 = hbusreq1_p & ad42e2 | !hbusreq1_p & v845542;
assign dc4fe6 = hbusreq4_p & dc4fe3 | !hbusreq4_p & dc4fe5;
assign v9ea5eb = hbusreq3_p & v9ea5bb | !hbusreq3_p & v9ea5ea;
assign v9f76ea = stateG2_p & v845542 | !stateG2_p & v9f7cf2;
assign c3cead = hready & c3ceac | !hready & v845542;
assign dc53b6 = jx1_p & dc5388 | !jx1_p & dc53b5;
assign d356a9 = hbusreq3 & d356a1 | !hbusreq3 & d356a8;
assign b57a8b = hgrant2_p & b57a8a | !hgrant2_p & b57a82;
assign c5c951 = hgrant2_p & c5c940 | !hgrant2_p & c5c93d;
assign v9f7645 = hbusreq4 & v9f7e41 | !hbusreq4 & v9f7e42;
assign v9ea594 = hbusreq1_p & v9ea3fa | !hbusreq1_p & v9ea586;
assign b57ae8 = hmaster0_p & b57ae4 | !hmaster0_p & b57ae7;
assign b05986 = hmaster2_p & b0597d | !hmaster2_p & !b05985;
assign ad4408 = hlock2_p & ad4405 | !hlock2_p & ad4407;
assign bd5839 = hmaster2_p & c3d669 | !hmaster2_p & !bd5838;
assign ad4e73 = hbusreq4_p & ad4e70 | !hbusreq4_p & ad4e72;
assign bd586a = hmaster2_p & bd5860 | !hmaster2_p & bd5869;
assign b1c712 = hmaster2_p & b1c70f | !hmaster2_p & b1c711;
assign b1c072 = hmaster2_p & b1c06e | !hmaster2_p & b1c071;
assign ad4563 = hlock4_p & ad4e4c | !hlock4_p & ad4f3e;
assign c3d2e3 = hready_p & v845555 | !hready_p & c3d2e2;
assign d35957 = hmaster2_p & adea8a | !hmaster2_p & !d35956;
assign bd5ba6 = hbusreq2_p & bd5ba5 | !hbusreq2_p & v845542;
assign ad4499 = hbusreq1_p & ad4487 | !hbusreq1_p & ad4484;
assign v9f7737 = hmaster1_p & v9f772e | !hmaster1_p & v9f7736;
assign c3d735 = hmaster1_p & c3d734 | !hmaster1_p & c3d6d2;
assign v9f7660 = hbusreq4_p & v9f765d | !hbusreq4_p & !v9f765f;
assign bd5931 = hbusreq0 & bd5930 | !hbusreq0 & v84556c;
assign v9f7730 = hmaster2_p & v9f772b | !hmaster2_p & v9f772f;
assign b1c74d = busreq_p & bb9bdd | !busreq_p & !v845542;
assign ad3d03 = hmaster2_p & ad3d02 | !hmaster2_p & v845542;
assign b579d9 = hmaster2_p & b579d8 | !hmaster2_p & b579cd;
assign d356f8 = hbusreq2 & d356f5 | !hbusreq2 & d356f7;
assign v9e9fbc = hmaster1_p & v9e9fbb | !hmaster1_p & v9e9ef1;
assign b1c046 = hbusreq4 & b1c042 | !hbusreq4 & b1c045;
assign ad47ed = hgrant2_p & ad47ea | !hgrant2_p & ad47ec;
assign v9f7de2 = hgrant4_p & v9f7cdc | !hgrant4_p & v9f7de1;
assign d35425 = hbusreq4 & d35424 | !hbusreq4 & d3541f;
assign c3ce2b = hgrant2_p & v845551 | !hgrant2_p & c3ce2a;
assign b058cd = hbusreq2 & b058cb | !hbusreq2 & b058cc;
assign ad459e = hready & ad456f | !hready & ad459c;
assign c3d58a = hbusreq3_p & c3d522 | !hbusreq3_p & c3d589;
assign c3d39b = stateG10_4_p & c3d399 | !stateG10_4_p & c3d39a;
assign ad4107 = hbusreq1 & ad480c | !hbusreq1 & v845542;
assign ad501b = hready & v84556c | !hready & !v845542;
assign v9f7893 = hbusreq1_p & v9f77ce | !hbusreq1_p & v9f788c;
assign b1c583 = hmaster0_p & b1c842 | !hmaster0_p & b1c582;
assign d356a0 = hlock1_p & d3569f | !hlock1_p & d355a3;
assign ad4fc9 = hmastlock_p & ad4fc8 | !hmastlock_p & !v845542;
assign ad4828 = decide_p & ad4820 | !decide_p & ad4827;
assign v9f77cf = hgrant1_p & v9f772d | !hgrant1_p & v9f77ce;
assign c3ce7a = hmaster0_p & c3ce79 | !hmaster0_p & c3d2be;
assign v8cc7ca = hgrant1_p & v845542 | !hgrant1_p & v8cc7c9;
assign c3d6df = hgrant2_p & c3d6da | !hgrant2_p & !c3d6de;
assign df516d = decide_p & df516c | !decide_p & v845542;
assign d356ef = hbusreq2_p & d356ee | !hbusreq2_p & d356ed;
assign ad4f7c = hbusreq0 & ad4f77 | !hbusreq0 & ad4f7b;
assign ad4767 = hlock4_p & ad4dc4 | !hlock4_p & !v845542;
assign ad4393 = hready & v845542 | !hready & ad4392;
assign ad441b = hmaster0_p & ad440e | !hmaster0_p & ad4413;
assign ad4815 = hready & ad4f3d | !hready & ad4814;
assign d357cd = hbusreq0 & d357cc | !hbusreq0 & v845542;
assign bd5b83 = hbusreq3 & bd5b82 | !hbusreq3 & v84556c;
assign c3d695 = hbusreq2_p & c3d692 | !hbusreq2_p & c3d694;
assign v8cc438 = hgrant4_p & v845542 | !hgrant4_p & v8ccbf0;
assign d3565c = hlock2_p & v845542 | !hlock2_p & d3565b;
assign b574b3 = hmaster2_p & v845542 | !hmaster2_p & b574b2;
assign c3ce8a = hgrant3_p & c3ce7e | !hgrant3_p & c3ce89;
assign c3d70f = hmaster0_p & c3d70e | !hmaster0_p & !c3d6fb;
assign b57411 = hbusreq1_p & b578f1 | !hbusreq1_p & b57410;
assign ade4c2 = hmastlock_p & ade4c1 | !hmastlock_p & v84557a;
assign d357dc = hbusreq0 & d357db | !hbusreq0 & v845542;
assign ad48a6 = hready & ad4ddd | !hready & ad48a5;
assign v9f76d8 = hmaster0_p & v9f7d34 | !hmaster0_p & v9f7d03;
assign ad4821 = hbusreq2 & ad4fb0 | !hbusreq2 & v845542;
assign c3cf07 = hready & c3cf06 | !hready & !c3cee3;
assign b1c55d = hbusreq4_p & b1cbf0 | !hbusreq4_p & !b1c857;
assign v9f7786 = hmaster2_p & v9f7785 | !hmaster2_p & d359c4;
assign v9f780a = hbusreq0_p & v9f77eb | !hbusreq0_p & v9f77ec;
assign d35437 = hbusreq0 & d35433 | !hbusreq0 & d35436;
assign b8f748 = hbusreq1_p & c3d328 | !hbusreq1_p & c3d2fd;
assign v8cc0c3 = hlock0_p & v8cc47a | !hlock0_p & v8cc0c2;
assign b1cf2d = hbusreq3 & b1cf28 | !hbusreq3 & b1cf2c;
assign b1c4a7 = hbusreq4 & b1c498 | !hbusreq4 & b1c4a6;
assign d3569c = jx1_p & d355a2 | !jx1_p & d3569b;
assign cc36dc = stateG10_4_p & cc36da | !stateG10_4_p & cc36db;
assign b1c7f6 = hmaster0_p & b1c7af | !hmaster0_p & b1c7f5;
assign v8da603 = hready_p & v8da5a6 | !hready_p & !v845564;
assign ad3d57 = hmaster1_p & ad3d56 | !hmaster1_p & ad3d12;
assign ad458e = hbusreq4 & ad4ecd | !hbusreq4 & v845542;
assign ad4760 = hmaster0_p & ad470d | !hmaster0_p & ad456f;
assign d356eb = hmaster0_p & d356e2 | !hmaster0_p & d356de;
assign b1c7db = hlock4_p & b1c7d9 | !hlock4_p & !b1c7da;
assign bd57e5 = hbusreq3 & bd579a | !hbusreq3 & bd579b;
assign v8ccb75 = hmaster2_p & v8d29fa | !hmaster2_p & v845542;
assign ade5a1 = hmaster2_p & adea94 | !hmaster2_p & ade5a0;
assign bd5755 = hbusreq4_p & adec89 | !hbusreq4_p & bd574e;
assign c3cefa = hmaster0_p & c3cef9 | !hmaster0_p & c3d306;
assign b579f0 = hmaster0_p & v845542 | !hmaster0_p & b579ef;
assign ad48c6 = hmaster1_p & ad5024 | !hmaster1_p & ad48c5;
assign bd5b75 = hbusreq2_p & bd5b74 | !hbusreq2_p & v845542;
assign ad4755 = decide_p & ad4606 | !decide_p & ad4754;
assign d356be = hmaster1_p & d356bd | !hmaster1_p & d356b8;
assign c3d5b3 = hgrant4_p & v845542 | !hgrant4_p & c3d5b2;
assign b1c4c9 = hmaster2_p & d35a9c | !hmaster2_p & !b1c4c8;
assign d3556a = hgrant2_p & d35567 | !hgrant2_p & d35569;
assign d35916 = hbusreq1_p & d35915 | !hbusreq1_p & d3590a;
assign d35690 = hmaster0_p & d35645 | !hmaster0_p & d3568f;
assign d357ba = hmaster2_p & d3576e | !hmaster2_p & d357b9;
assign b1c566 = hbusreq0 & b1c563 | !hbusreq0 & b1c565;
assign c3d51c = hgrant1_p & c3d2de | !hgrant1_p & c3d51b;
assign d359ce = hlock0_p & d35983 | !hlock0_p & d359cd;
assign d3564c = hgrant4_p & v84556c | !hgrant4_p & d3564b;
assign hgrant0 = !b1c0b5;
assign ad4eeb = hbusreq4_p & ad4ed3 | !hbusreq4_p & ad4eea;
assign dc4fec = hmaster2_p & dc4feb | !hmaster2_p & v845542;
assign ad4149 = hgrant2_p & v845542 | !hgrant2_p & ad4148;
assign bd5773 = hbusreq2 & bd5772 | !hbusreq2 & v845542;
assign c3ce29 = hmaster0_p & c3d3a5 | !hmaster0_p & c3cdfe;
assign v8cc80b = hgrant2_p & v8cc7ad | !hgrant2_p & v8cc80a;
assign c3d6ab = hgrant0_p & c3d670 | !hgrant0_p & !c3d66d;
assign bd57f3 = hbusreq1_p & bd57f1 | !hbusreq1_p & bd57f2;
assign v9e9f91 = hbusreq4_p & v9ea462 | !hbusreq4_p & v9e9f90;
assign b1c796 = hbusreq0_p & bd58a2 | !hbusreq0_p & !v845542;
assign bd58c8 = hgrant4_p & v845542 | !hgrant4_p & !bd58c6;
assign df5147 = hbusreq1 & dc4fcb | !hbusreq1 & v845542;
assign ad4157 = hmaster2_p & ad4151 | !hmaster2_p & ad4156;
assign ad4284 = hbusreq3 & ad4281 | !hbusreq3 & !v845542;
assign d35bf7 = hmaster2_p & v845542 | !hmaster2_p & d35bf6;
assign ad4f92 = hbusreq4_p & ad4f91 | !hbusreq4_p & ad4f80;
assign bd5b93 = locked_p & bd5b92 | !locked_p & v845542;
assign c3d6ec = stateG10_4_p & c3d6b7 | !stateG10_4_p & c3d6eb;
assign d35a9d = hmaster2_p & d35a9b | !hmaster2_p & d35a9c;
assign c3ce4b = hlock1_p & c3ce49 | !hlock1_p & c3ce4a;
assign ad4463 = hbusreq4_p & ad4462 | !hbusreq4_p & adeaa4;
assign ad4366 = hlock2_p & ad4361 | !hlock2_p & !ad4365;
assign ad46ab = hmaster2_p & ad46aa | !hmaster2_p & v845542;
assign dc4f62 = hmaster0_p & dc4f61 | !hmaster0_p & v84556c;
assign adeab1 = hmaster1_p & v845542 | !hmaster1_p & adeab0;
assign v8ccbd6 = hbusreq2_p & v8ccb8f | !hbusreq2_p & v8ccb8d;
assign v9e9f96 = hready & v9e9f95 | !hready & v9e9f8e;
assign b0594e = locked_p & b0591c | !locked_p & !b058a3;
assign ad4e8d = hbusreq4_p & ad4e8c | !hbusreq4_p & b1cfcb;
assign ad46a6 = hgrant0_p & v845542 | !hgrant0_p & ad46a5;
assign ade5d9 = hmaster0_p & ade5d4 | !hmaster0_p & !ade5d8;
assign ad3d26 = hbusreq2_p & ad3d23 | !hbusreq2_p & ad3d25;
assign d35950 = hbusreq1 & d3590e | !hbusreq1 & d3594f;
assign ade5cf = hbusreq4_p & ade5ce | !hbusreq4_p & !v845542;
assign v8cc48c = hlock2 & v8cc489 | !hlock2 & v8cc48a;
assign df552b = decide_p & df54ee | !decide_p & d6ebca;
assign ad4ff1 = hbusreq3 & ad4fd0 | !hbusreq3 & v845542;
assign d3598c = hbusreq3 & d3598b | !hbusreq3 & v845542;
assign b1c72d = hbusreq3 & b1c722 | !hbusreq3 & b1c71d;
assign v9e9fc0 = hmaster0_p & v9e9eed | !hmaster0_p & v9e9ee8;
assign c3d6ef = hbusreq1_p & c3d6e7 | !hbusreq1_p & c3d6ee;
assign ad436c = hmaster0_p & df5142 | !hmaster0_p & ad4291;
assign stateG10_4 = !ba7c81;
assign ad3cd0 = hgrant1_p & ad4411 | !hgrant1_p & ad3ccf;
assign ad43f6 = hlock0_p & adea85 | !hlock0_p & !ad43cf;
assign v8d2b2b = locked_p & v8d29fa | !locked_p & v845542;
assign v9f7d65 = hmaster1_p & v9f7d5c | !hmaster1_p & v9f7d64;
assign ad3d41 = hmaster0_p & ad43aa | !hmaster0_p & ad43a9;
assign adea99 = hburst0 & adea97 | !hburst0 & adea98;
assign v8cc7ad = hmaster1_p & v8cc7ab | !hmaster1_p & v845542;
assign bd58ec = hbusreq2_p & bd58eb | !hbusreq2_p & v845542;
assign bd5871 = hgrant0_p & adec9a | !hgrant0_p & adec89;
assign v9f7cc3 = hmaster0_p & v9f7cb2 | !hmaster0_p & v9f7cc2;
assign ad508d = hmaster0_p & v845547 | !hmaster0_p & v845542;
assign c3d6e0 = hbusreq2_p & c3d6d8 | !hbusreq2_p & !c3d6df;
assign d35a33 = hmaster0_p & d359ac | !hmaster0_p & d35a32;
assign ad437d = hbusreq0_p & ad4e47 | !hbusreq0_p & v845542;
assign d3574d = hmaster0_p & d3574b | !hmaster0_p & !d3574c;
assign c3d2e0 = hmaster0_p & c3d2df | !hmaster0_p & !c3d2be;
assign d6ebc9 = hready_p & v845542 | !hready_p & v845560;
assign d35994 = hbusreq1_p & d35993 | !hbusreq1_p & !d35992;
assign d35a15 = hbusreq4_p & d35a13 | !hbusreq4_p & d35a14;
assign b1c719 = hbusreq3 & b1c713 | !hbusreq3 & b1c718;
assign b1cffc = hbusreq0 & b1cff7 | !hbusreq0 & b1cffb;
assign d35713 = hmaster0_p & d35711 | !hmaster0_p & !d35712;
assign ad481d = hbusreq2 & ad4f1a | !hbusreq2 & v845542;
assign v9e9ea4 = hbusreq1 & v9ea482 | !hbusreq1 & v9ea46d;
assign bd5ea4 = hmaster0_p & v84556c | !hmaster0_p & bd5ea3;
assign b1c846 = hbusreq4_p & v84554a | !hbusreq4_p & v845542;
assign b1cf43 = hmaster1_p & v845542 | !hmaster1_p & b1cf42;
assign v9e9ee3 = hready_p & v9ea436 | !hready_p & v9e9ee2;
assign df5161 = hbusreq1 & dc4f81 | !hbusreq1 & v845542;
assign d35642 = hlock4_p & d35640 | !hlock4_p & !d35641;
assign bd58cf = hmaster2_p & bd58ce | !hmaster2_p & bd58c1;
assign c3d6f0 = hgrant1_p & c3d6ea | !hgrant1_p & c3d6ef;
assign d35745 = hmaster1_p & d35744 | !hmaster1_p & d35713;
assign ad4e43 = hbusreq3 & ad4e42 | !hbusreq3 & v845542;
assign d359cb = hbusreq1 & d359ca | !hbusreq1 & !v845542;
assign v9f772b = hmastlock_p & v9f772a | !hmastlock_p & !v845542;
assign b05a2b = hready_p & b05a02 | !hready_p & !b05a2a;
assign b05980 = hlock0_p & b0597e | !hlock0_p & !b0597f;
assign v9f7679 = hbusreq3 & v9f7e39 | !hbusreq3 & v9f7678;
assign c3cef8 = hready & c3cef7 | !hready & c3d305;
assign bd58f4 = decide_p & bd58f3 | !decide_p & v845542;
assign c3d73d = locked_p & c3d667 | !locked_p & c3d669;
assign v9ea415 = hmaster2_p & v845542 | !hmaster2_p & v9ea414;
assign dc5086 = hready_p & dc5082 | !hready_p & dc5085;
assign b1c783 = hmaster1_p & b1c782 | !hmaster1_p & b1c775;
assign ad4692 = hbusreq4_p & ad4691 | !hbusreq4_p & v845542;
assign v9ea40f = hmaster2_p & v9ea40e | !hmaster2_p & v845542;
assign dc5026 = hbusreq0 & dc5020 | !hbusreq0 & dc5025;
assign df51d0 = hready_p & df51cf | !hready_p & df5541;
assign bd57ec = hlock2_p & bd57e8 | !hlock2_p & !bd57eb;
assign b1cfb8 = hgrant1_p & v845542 | !hgrant1_p & b1cfb7;
assign dc4f80 = hbusreq0 & dc4f7e | !hbusreq0 & dc4f7f;
assign b1c800 = hmaster0_p & b1c7ff | !hmaster0_p & b1c73a;
assign d354bb = hlock1_p & d354b9 | !hlock1_p & !d354ba;
assign b1c788 = hlock3_p & b1c77e | !hlock3_p & b1c787;
assign b574bd = hbusreq3 & b574bb | !hbusreq3 & b574bc;
assign ad470c = hbusreq4 & ad470b | !hbusreq4 & v845542;
assign bd5879 = hbusreq4_p & bd5876 | !hbusreq4_p & bd5878;
assign b57440 = hbusreq2_p & b5743c | !hbusreq2_p & b5743f;
assign ad4e6c = locked_p & ad4e6b | !locked_p & !v845542;
assign ad4f6b = hbusreq4_p & ad4f68 | !hbusreq4_p & ad4f6a;
assign ade541 = hbusreq2 & adec92 | !hbusreq2 & adec9c;
assign ade5c0 = hbusreq3 & ade5ac | !hbusreq3 & !v845558;
assign v9f779d = locked_p & v845542 | !locked_p & !v9f772f;
assign ad432a = decide_p & ad4310 | !decide_p & ad4329;
assign ad4357 = decide_p & ad4351 | !decide_p & !ad4356;
assign dc4fab = hbusreq0 & dc4fa8 | !hbusreq0 & dc4faa;
assign v9f7d53 = hmaster0_p & v9f7d3c | !hmaster0_p & v9f7d3e;
assign v9ea4d0 = hgrant4_p & v9ea4b3 | !hgrant4_p & v9ea4c6;
assign v9f7777 = hbusreq3 & v9f7760 | !hbusreq3 & v9f7776;
assign b1cfd0 = hbusreq0 & b1cfca | !hbusreq0 & b1cfcf;
assign d359ed = hmastlock_p & v845542 | !hmastlock_p & !d359ba;
assign d357ae = hmaster1_p & d35799 | !hmaster1_p & d357a6;
assign c3d6d2 = hmaster0_p & c3d6bf | !hmaster0_p & c3d6d1;
assign ad47eb = hmaster0_p & ad46f6 | !hmaster0_p & ad46af;
assign v9f7720 = hbusreq2_p & v9f771b | !hbusreq2_p & v9f771f;
assign d359e5 = hbusreq1 & d3598b | !hbusreq1 & v845542;
assign dc4fbf = hbusreq3 & dc4fbe | !hbusreq3 & v845542;
assign b1c7b9 = hbusreq1 & b1c7b5 | !hbusreq1 & !b1c7b8;
assign v9e9ebd = hgrant2_p & v9e9eb7 | !hgrant2_p & v9e9ebc;
assign bd593a = hlock2_p & bd5939 | !hlock2_p & !v845542;
assign ad4f06 = hbusreq0 & ad4efc | !hbusreq0 & ad4f05;
assign bd579e = hmaster2_p & bd5786 | !hmaster2_p & !ade4d4;
assign ad4fbe = hmaster2_p & ad4fbd | !hmaster2_p & v845542;
assign bd58ea = hmaster1_p & bd58e9 | !hmaster1_p & bd5779;
assign ad4101 = hgrant0_p & v845542 | !hgrant0_p & !ad4100;
assign d3563e = hgrant0_p & v845542 | !hgrant0_p & d3563c;
assign dc503b = stateG10_4_p & adeca1 | !stateG10_4_p & !dc503a;
assign v9e9ef5 = hbusreq2_p & v9e9ef2 | !hbusreq2_p & v9e9ef4;
assign ad4e9e = hgrant4_p & v84556c | !hgrant4_p & v845542;
assign c3ced9 = hready_p & c3ced7 | !hready_p & c3ced8;
assign bd58b9 = hbusreq2 & bd58b8 | !hbusreq2 & v845542;
assign v8cc481 = hbusreq4 & v8cc47d | !hbusreq4 & v8cc47f;
assign ad3cc2 = hmaster1_p & ad3cc1 | !hmaster1_p & ad3cbb;
assign b57982 = hbusreq2_p & b5795b | !hbusreq2_p & b5795a;
assign v9f7d14 = hbusreq0 & v9f7d04 | !hbusreq0 & v9f7d13;
assign v9f7d72 = hlock0_p & v9f7d70 | !hlock0_p & v9f7d71;
assign v9e9ed5 = hbusreq2_p & v9e9ed0 | !hbusreq2_p & v9e9ed4;
assign dc53d6 = decide_p & dc53d5 | !decide_p & v845542;
assign ad4329 = hbusreq2_p & ad431e | !hbusreq2_p & ad4328;
assign d354d0 = hmaster2_p & v845542 | !hmaster2_p & d354cf;
assign dc4f76 = hmaster2_p & dc4f74 | !hmaster2_p & !ade4e8;
assign v9f76f8 = hlock1 & v9f76f2 | !hlock1 & v9f76f7;
assign v9e9f5b = hready & v9e9f5a | !hready & v9e9f57;
assign c3d3a2 = hbusreq0 & c3d3a1 | !hbusreq0 & v845542;
assign ad468b = hbusreq2 & ad457d | !hbusreq2 & v845542;
assign b57538 = jx2_p & b57b5c | !jx2_p & b57537;
assign ad4569 = hmaster2_p & v845542 | !hmaster2_p & ad4568;
assign b1c08d = hbusreq2_p & b1c057 | !hbusreq2_p & b1c08c;
assign v9ea44e = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea44d;
assign v9e9ee0 = hgrant2_p & v9e9ede | !hgrant2_p & v9e9edf;
assign b1cfca = hmaster2_p & b1cfbf | !hmaster2_p & b1cfb7;
assign ade5cd = hburst1 & ade4c8 | !hburst1 & ade5cc;
assign c3d70d = hbusreq1_p & c3d709 | !hbusreq1_p & c3d70c;
assign b059a4 = hmaster1_p & b059a3 | !hmaster1_p & b05913;
assign b1c797 = hlock0_p & b1c795 | !hlock0_p & b1c796;
assign v9e9ebc = hmaster1_p & v9e9ebb | !hmaster1_p & v9e9ead;
assign v8cc79e = hbusreq1 & v8cc79c | !hbusreq1 & v8cc79d;
assign d3574e = hmaster1_p & d3574a | !hmaster1_p & d3574d;
assign v9f7d09 = hbusreq4 & v9f7d07 | !hbusreq4 & v9f7d08;
assign b579b3 = hmaster2_p & b579b2 | !hmaster2_p & v845542;
assign ade54e = hburst1 & ade54d | !hburst1 & v845542;
assign v8cc0dd = hbusreq4 & v8cc0dc | !hbusreq4 & v8cc494;
assign v9f77e9 = stateG10_4_p & v845542 | !stateG10_4_p & !v9f77e8;
assign df553d = hmaster1_p & df5539 | !hmaster1_p & df553c;
assign d357c3 = hgrant4_p & v84554a | !hgrant4_p & d357c1;
assign c3d506 = hmaster0_p & c3d4f8 | !hmaster0_p & c3d505;
assign df5114 = hgrant3_p & df50de | !hgrant3_p & df50d4;
assign d35779 = hmaster0_p & d35777 | !hmaster0_p & d35778;
assign ad457b = hbusreq4 & ad457a | !hbusreq4 & v845542;
assign adea8f = decide_p & adea8d | !decide_p & v845542;
assign v84556c = locked_p & v845542 | !locked_p & !v845542;
assign c3d310 = hbusreq4 & c3d30c | !hbusreq4 & !c3d30f;
assign v9e9fa6 = hbusreq2 & v9e9fa5 | !hbusreq2 & v9e9f68;
assign bd581e = hgrant4_p & v845542 | !hgrant4_p & !bd580d;
assign c3d6f4 = hbusreq4_p & c3d6f1 | !hbusreq4_p & !c3d6f3;
assign ad4161 = hmaster0_p & ad414f | !hmaster0_p & ad4160;
assign cc36d4 = hgrant2_p & cc36d3 | !hgrant2_p & !cc36d0;
assign dc4f7b = hburst1 & dc4f78 | !hburst1 & dc4f7a;
assign d356f3 = hbusreq2 & d356ab | !hbusreq2 & d356ad;
assign bd572f = hmastlock_p & adec8c | !hmastlock_p & !d359ba;
assign bd5b85 = hmastlock_p & bd5b84 | !hmastlock_p & v845542;
assign v9f7872 = hmaster1_p & v9f786a | !hmaster1_p & v9f7871;
assign ad410f = hbusreq1_p & ad410e | !hbusreq1_p & v845547;
assign b1cf38 = hbusreq2_p & b1cf2f | !hbusreq2_p & b1cf37;
assign b05959 = hbusreq4_p & b05957 | !hbusreq4_p & b05958;
assign b57408 = locked_p & b57407 | !locked_p & v845542;
assign b05a79 = hbusreq1_p & b05962 | !hbusreq1_p & b05a70;
assign c3d6b3 = hlock1_p & c3d66f | !hlock1_p & !c3d682;
assign c5c9b4 = hready_p & c5c953 | !hready_p & !c5c9b3;
assign v9f767f = hgrant1_p & v9f7cc8 | !hgrant1_p & v9f7e3f;
assign v9e9f58 = hbusreq0 & v9e9f53 | !hbusreq0 & v9e9f57;
assign ad42f9 = hmaster0_p & ad42f3 | !hmaster0_p & ad42f8;
assign ad4558 = hlock4_p & dc52fa | !hlock4_p & ad4f39;
assign c3cf08 = hgrant1_p & v845542 | !hgrant1_p & c3cf07;
assign b579ec = hbusreq1 & b579c0 | !hbusreq1 & b579c1;
assign v9f7ddb = stateG10_4_p & v9f7d42 | !stateG10_4_p & v9f7dda;
assign ad434b = hgrant3_p & ad42dc | !hgrant3_p & ad434a;
assign v9f782c = stateG10_4_p & v9f782a | !stateG10_4_p & v9f782b;
assign v8cc6b5 = hgrant3_p & v8cc634 | !hgrant3_p & v8cc6b4;
assign ade567 = hmaster2_p & ade561 | !hmaster2_p & ade566;
assign d35a06 = hlock4_p & d35a04 | !hlock4_p & d35a05;
assign df514e = hmaster1_p & df5144 | !hmaster1_p & df514d;
assign ac1461 = hgrant4_p & ac144e | !hgrant4_p & !v845542;
assign df553b = hgrant1_p & df553a | !hgrant1_p & !v845542;
assign ad4475 = hgrant2_p & ad446d | !hgrant2_p & ad4474;
assign b579bb = hmaster2_p & v845542 | !hmaster2_p & b579ba;
assign ad4e82 = hgrant4_p & v84556c | !hgrant4_p & b1cfb6;
assign v9f7785 = locked_p & v9f772b | !locked_p & v9f7743;
assign b579b6 = hburst0_p & v9ea411 | !hburst0_p & !b579b5;
assign ad3cff = hgrant4_p & ad440b | !hgrant4_p & c3cec2;
assign ad42c7 = hbusreq2_p & ad42c6 | !hbusreq2_p & ad42c5;
assign df5133 = hgrant3_p & df511d | !hgrant3_p & df5132;
assign v9f7cdb = hbusreq0_p & v9f7cb6 | !hbusreq0_p & !v9f7cc7;
assign c3d762 = hgrant3_p & c3d731 | !hgrant3_p & !c3d761;
assign ad4482 = hbusreq4_p & ad4480 | !hbusreq4_p & ad4481;
assign b57a67 = hmaster2_p & v845542 | !hmaster2_p & b57a66;
assign b05a13 = hbusreq4_p & b05a11 | !hbusreq4_p & b05a12;
assign ad4290 = hbusreq1 & ad4fb0 | !hbusreq1 & v845542;
assign ad4401 = hlock2_p & ad43fd | !hlock2_p & ad4400;
assign c3d4de = hlock4_p & c3d2f0 | !hlock4_p & c3d33c;
assign adeab6 = decide_p & adeab1 | !decide_p & adeaa7;
assign c5c96c = hmaster0_p & c5c969 | !hmaster0_p & !v845542;
assign b1caea = hmaster2_p & v845542 | !hmaster2_p & !b1cae9;
assign ad506d = hgrant2_p & ad506b | !hgrant2_p & ad5067;
assign v84557c = stateG2_p & v845542 | !stateG2_p & !v845542;
assign df54fb = hmaster0_p & df54fa | !hmaster0_p & df54f4;
assign c3cf13 = hmaster1_p & c3cf12 | !hmaster1_p & c3d36b;
assign v9f778f = hlock2 & v9f772c | !hlock2 & v9f778e;
assign d35aa7 = hmaster1_p & v845542 | !hmaster1_p & d35aa6;
assign b06735 = stateG2_p & v845542 | !stateG2_p & c6d44d;
assign b1c064 = stateG10_4_p & b1c062 | !stateG10_4_p & !b1c063;
assign ad48a5 = hmaster2_p & v845542 | !hmaster2_p & !ad4dde;
assign v9ea49b = hmaster0_p & v9ea44a | !hmaster0_p & v9ea49a;
assign b1cbf1 = hbusreq4_p & b1cbf0 | !hbusreq4_p & b1cfb7;
assign b1c5bb = hlock0_p & b1c5ba | !hlock0_p & v845542;
assign df5152 = hmaster0_p & df513f | !hmaster0_p & df5151;
assign ad43da = hmaster2_p & ad43c4 | !hmaster2_p & v845542;
assign c3d67d = hmaster1_p & c3d672 | !hmaster1_p & c3d67c;
assign dc4fa3 = hmaster2_p & ade4bf | !hmaster2_p & !v845542;
assign ad4299 = hmaster0_p & ad4291 | !hmaster0_p & df5142;
assign bd5802 = hbusreq4_p & bd57ff | !hbusreq4_p & bd5801;
assign d35413 = hmaster0_p & d35c04 | !hmaster0_p & d35412;
assign d35726 = hbusreq3 & d35717 | !hbusreq3 & !v84554e;
assign b058bb = hlock4 & b058b8 | !hlock4 & b058ba;
assign d355b0 = decide_p & d355af | !decide_p & v84556c;
assign v9f7802 = hbusreq2_p & v9f77f8 | !hbusreq2_p & v9f7801;
assign ad4eb6 = stateG10_4_p & ad4eb3 | !stateG10_4_p & ad4eb5;
assign v9ea41a = stateG10_4_p & v845542 | !stateG10_4_p & v9ea419;
assign v9f783f = stateG10_4_p & v845542 | !stateG10_4_p & !v9f783e;
assign ad47f4 = hmaster1_p & ad47f3 | !hmaster1_p & ad46ec;
assign ad476b = hready & ad45ad | !hready & !ad476a;
assign ad3d48 = hmaster1_p & ad3cc0 | !hmaster1_p & ad3cbb;
assign ad3d58 = hgrant2_p & ad3d55 | !hgrant2_p & ad3d57;
assign b05a3a = hmaster0_p & b05920 | !hmaster0_p & b0591e;
assign v9f78b0 = jx0_p & v9f7725 | !jx0_p & !v9f78af;
assign b1c5ec = hbusreq0 & b1c5e7 | !hbusreq0 & b1c5eb;
assign v9e9eb8 = hmaster2_p & v9e9e9e | !hmaster2_p & v9ea45a;
assign v8cc488 = hgrant1_p & v8cc487 | !hgrant1_p & v8cc474;
assign ad4f03 = stateG10_4_p & ad4f00 | !stateG10_4_p & !ad4f02;
assign dc5388 = hbusreq3_p & dc5387 | !hbusreq3_p & !dc5088;
assign v9e9fe0 = hmaster1_p & v9ea49a | !hmaster1_p & v9e9fd0;
assign ad4787 = hmaster1_p & ad4786 | !hmaster1_p & ad460e;
assign ac1495 = hbusreq3_p & ac1482 | !hbusreq3_p & ac1494;
assign bd590e = hbusreq2_p & bd590d | !hbusreq2_p & v845542;
assign ad4f64 = hgrant4_p & ad4f36 | !hgrant4_p & v845542;
assign v9f7dfa = hmaster0_p & v9f7d10 | !hmaster0_p & v9f7d03;
assign ad4e97 = hbusreq1_p & ad4e94 | !hbusreq1_p & !ad4e96;
assign v9e9fb8 = hbusreq2 & v9e9fb6 | !hbusreq2 & v9e9fb7;
assign b1c7f5 = hgrant1_p & b1c7f4 | !hgrant1_p & b1c7c9;
assign dc4fc8 = hready_p & dc4f64 | !hready_p & !dc4fc7;
assign v9ea58a = hbusreq0 & v9ea588 | !hbusreq0 & v9ea589;
assign b059e3 = hlock0_p & b0598b | !hlock0_p & b059e2;
assign df5543 = hgrant3_p & df5531 | !hgrant3_p & df5542;
assign c5c8ea = hmaster0_p & c5c8e8 | !hmaster0_p & c5c8e9;
assign v8cc760 = hmaster0_p & v8cc489 | !hmaster0_p & v8cc75f;
assign ad4133 = hbusreq4_p & ad4132 | !hbusreq4_p & ad4e9b;
assign v8cc7fd = hbusreq0 & v8cc7fa | !hbusreq0 & v8cc7fc;
assign bd580c = hgrant0_p & v845542 | !hgrant0_p & !adec89;
assign d35aba = decide_p & d35ab9 | !decide_p & v84556c;
assign ad4562 = hbusreq4 & ad4561 | !hbusreq4 & v845542;
assign d356c1 = hlock1_p & d359c5 | !hlock1_p & !v845542;
assign c3d702 = hmaster0_p & c3d6e8 | !hmaster0_p & c3d701;
assign b05a69 = hmaster2_p & b05a68 | !hmaster2_p & v9f7d42;
assign b05a1a = hbusreq4_p & b05a17 | !hbusreq4_p & b05a19;
assign b05a02 = decide_p & b059ad | !decide_p & b05a01;
assign d35593 = hmaster1_p & d35584 | !hmaster1_p & d35592;
assign ad4eba = hgrant4_p & ad4e53 | !hgrant4_p & v845542;
assign d35625 = hlock1_p & d35623 | !hlock1_p & d35624;
assign c5c97b = hmaster0_p & c5c969 | !hmaster0_p & c5c97a;
assign b05973 = hbusreq3 & b0596d | !hbusreq3 & b05972;
assign c3d5cb = hready & c3d5ca | !hready & c3d300;
assign b1cf3d = hmaster1_p & v845542 | !hmaster1_p & b1cf3c;
assign ad438f = hready & v845542 | !hready & ad438e;
assign ad5043 = stateG10_4_p & ad5041 | !stateG10_4_p & ad5042;
assign d3599f = hgrant4_p & v84557a | !hgrant4_p & !v845542;
assign d35a41 = hgrant0_p & v84556c | !hgrant0_p & d35a40;
assign v9e9f65 = hmastlock_p & v9e9f64 | !hmastlock_p & v845542;
assign v9e9e69 = hgrant1_p & v9ea43d | !hgrant1_p & v9ea45b;
assign d35526 = hmaster2_p & d35a9b | !hmaster2_p & d35525;
assign v9f77a0 = hlock0 & v9f779f | !hlock0 & v9f779e;
assign v9f77f5 = hmaster1_p & v9f77d4 | !hmaster1_p & v9f77f4;
assign b058ec = hbusreq0 & b058e8 | !hbusreq0 & b058eb;
assign ad415c = hbusreq0 & ad415a | !hbusreq0 & ad415b;
assign b05a8e = hmaster0_p & b0593d | !hmaster0_p & b0593a;
assign b1cf46 = hbusreq2_p & b1cf3d | !hbusreq2_p & b1cf45;
assign ad439a = hbusreq3 & ad4399 | !hbusreq3 & v845542;
assign v9f7762 = hlock1_p & v9f7745 | !hlock1_p & v9f7751;
assign v9f7dd8 = hgrant4_p & v9f7cf7 | !hgrant4_p & v9f7d8a;
assign d35431 = hlock4_p & v845542 | !hlock4_p & d35918;
assign ad5061 = hbusreq4_p & ad505f | !hbusreq4_p & !ad5060;
assign d356fd = hmaster1_p & d356f9 | !hmaster1_p & d356fc;
assign b1c5b6 = hlock0_p & d35617 | !hlock0_p & v845542;
assign ad46b5 = hbusreq1 & ad46b4 | !hbusreq1 & !v845547;
assign v9ea5af = hbusreq3 & v9ea5ad | !hbusreq3 & v9ea5ae;
assign b05950 = hgrant4_p & b058a3 | !hgrant4_p & b0594f;
assign d3579b = hbusreq1_p & d3579a | !hbusreq1_p & d35799;
assign dc4fc6 = hlock3_p & dc4f98 | !hlock3_p & dc4fc5;
assign d359c2 = hmaster2_p & v845542 | !hmaster2_p & !d359c1;
assign ad4303 = hlock2_p & ad42fb | !hlock2_p & !ad4302;
assign d354b5 = hbusreq4_p & d354b4 | !hbusreq4_p & v845542;
assign v9f7750 = hmaster2_p & v9f7743 | !hmaster2_p & !v845542;
assign ad43b5 = hbusreq1_p & ad43ab | !hbusreq1_p & ad43aa;
assign b1c713 = hbusreq0 & b1c712 | !hbusreq0 & v845542;
assign c3d674 = hmastlock_p & c3d673 | !hmastlock_p & v845542;
assign d3549b = hbusreq2 & d35bf3 | !hbusreq2 & d35be8;
assign b573dc = hlock2 & b579e5 | !hlock2 & b573db;
assign v9f7d47 = hmaster0_p & v9f7d3f | !hmaster0_p & v9f7d46;
assign c3cf2a = hgrant3_p & c3cf27 | !hgrant3_p & c3cf29;
assign ad46cc = hbusreq0 & ad46c9 | !hbusreq0 & ad46cb;
assign b05a9c = jx1_p & v857463 | !jx1_p & !b05a9b;
assign v9f7769 = stateG10_4_p & v845542 | !stateG10_4_p & !v9f772f;
assign v9f77d9 = hlock0 & v9f77d8 | !hlock0 & v9f77d7;
assign v9f76a9 = hmaster0_p & v9f7d5b | !hmaster0_p & v9f7692;
assign ad42d6 = hbusreq1_p & ad42d5 | !hbusreq1_p & v845547;
assign ad469d = hlock4_p & ad4e8c | !hlock4_p & b1cfcb;
assign ad42bd = hmaster0_p & ad42ab | !hmaster0_p & ad42bc;
assign ade4cb = hburst1 & ade4c8 | !hburst1 & ade4ca;
assign ad4720 = hgrant1_p & ad456f | !hgrant1_p & ad4702;
assign v9f7e32 = hmaster2_p & v9f7ca5 | !hmaster2_p & !v9f7e31;
assign bd57e4 = hbusreq2_p & bd57e3 | !hbusreq2_p & v845542;
assign b1c617 = hlock1_p & b1c616 | !hlock1_p & b1cf3b;
assign b058c6 = hmaster0_p & b058b5 | !hmaster0_p & b058c5;
assign b1c7e8 = hmaster0_p & b1c7e6 | !hmaster0_p & b1c7e7;
assign dc5024 = hbusreq4_p & dc5021 | !hbusreq4_p & dc5023;
assign bd5e9b = hmaster2_p & v84556c | !hmaster2_p & bd5e9a;
assign b573d9 = hgrant1_p & v845542 | !hgrant1_p & b573d8;
assign bd5768 = hmaster2_p & c3d669 | !hmaster2_p & ade589;
assign ad4350 = hmaster1_p & ad434f | !hmaster1_p & ad4289;
assign v8cc5c8 = hready_p & v8cc455 | !hready_p & v8cc5c7;
assign c5c3bf = jx0_p & c5c9b6 | !jx0_p & c5c3be;
assign v8cc4bb = hmaster1_p & v8cc4ba | !hmaster1_p & v845542;
assign bd5922 = jx1_p & bd5921 | !jx1_p & bd5bb2;
assign v9f77a8 = hlock3 & v9f77a7 | !hlock3 & v9f77a6;
assign v845562 = hmaster1_p & v845542 | !hmaster1_p & !v845542;
assign v9f766f = hgrant1_p & v9f7ce4 | !hgrant1_p & v9f766e;
assign bd56d5 = hbusreq4_p & bd56d4 | !hbusreq4_p & !v845542;
assign ad46c5 = hbusreq1 & ad458f | !hbusreq1 & v845542;
assign ad46d1 = hlock4_p & ad4f0e | !hlock4_p & ad4f3e;
assign d3564b = hlock0_p & d3564a | !hlock0_p & !ade562;
assign cc3700 = hbusreq4_p & cc36cb | !hbusreq4_p & !cc36ff;
assign bd56dc = hmaster1_p & bd56db | !hmaster1_p & v845542;
assign v9f7cb1 = hlock2 & v9f7ca7 | !hlock2 & v9f7cb0;
assign ade55f = hgrant4_p & v84556c | !hgrant4_p & !ade557;
assign dc5318 = hmastlock_p & ade4b8 | !hmastlock_p & v845542;
assign c3ce1c = hbusreq2 & c3d376 | !hbusreq2 & v845542;
assign ad4fac = stateA1_p & v845542 | !stateA1_p & !ad4fab;
assign ad45aa = decide_p & ad4597 | !decide_p & ad45a9;
assign v9e9f49 = hmaster0_p & v9e9ee9 | !hmaster0_p & v9e9ee8;
assign v9ea572 = hmaster2_p & v9ea570 | !hmaster2_p & v9ea3fb;
assign b05a84 = hbusreq2_p & b05a55 | !hbusreq2_p & b05a83;
assign d3562f = hlock2_p & v845542 | !hlock2_p & !d3562e;
assign b05a68 = hbusreq4_p & b05950 | !hbusreq4_p & b05a67;
assign b05941 = hlock0_p & v9ea463 | !hlock0_p & b05940;
assign ad4346 = hmaster1_p & ad4345 | !hmaster1_p & ad42d9;
assign v8cc0f5 = hmaster1_p & v8cc0f4 | !hmaster1_p & v845542;
assign c3d525 = hbusreq4 & c3d524 | !hbusreq4 & !v845564;
assign c3d6bf = hgrant1_p & c3d6b6 | !hgrant1_p & c3d6be;
assign v9ea404 = hmaster2_p & v9ea401 | !hmaster2_p & v9ea403;
assign df5194 = hbusreq1 & dc5033 | !hbusreq1 & v845542;
assign d3556e = hgrant2_p & d3556d | !hgrant2_p & !d35569;
assign c3ce95 = hmaster1_p & c3ce93 | !hmaster1_p & c3ce94;
assign ad4267 = hbusreq1 & ad4f3b | !hbusreq1 & v845542;
assign dc4f75 = hmaster2_p & dc4f74 | !hmaster2_p & ade4e1;
assign df5159 = hbusreq1_p & df5158 | !hbusreq1_p & v845542;
assign v9f7cc0 = hbusreq3 & v9f7cbe | !hbusreq3 & v9f7cbf;
assign d3550b = hmaster2_p & d3541f | !hmaster2_p & d35509;
assign d354be = hbusreq1 & d354bd | !hbusreq1 & !v84555a;
assign ad4576 = hready & ad4575 | !hready & ad456f;
assign b05a71 = hbusreq1_p & b0596b | !hbusreq1_p & b05a70;
assign bd5b6f = hmaster2_p & v845542 | !hmaster2_p & bd5b6e;
assign v9e9eae = hmaster1_p & v9e9ea1 | !hmaster1_p & v9e9ead;
assign v9f7d70 = hgrant0_p & v9f7c9c | !hgrant0_p & !v9f7d6f;
assign cc36f1 = hbusreq0_p & ade562 | !hbusreq0_p & v845542;
assign v9ea3e8 = hbusreq1_p & v9f20a1 | !hbusreq1_p & v9ea3e7;
assign v8cc49e = hgrant4_p & v8cc47a | !hgrant4_p & v845542;
assign c3d5e5 = hready & c3d5e4 | !hready & c3d313;
assign v9f7835 = hbusreq1 & v9f7833 | !hbusreq1 & v9f7834;
assign v9f771c = hmaster0_p & v9f7d5e | !hmaster0_p & v9f7692;
assign d35653 = hgrant4_p & v84556c | !hgrant4_p & !d35652;
assign v9ea5a7 = hbusreq3 & v9ea5a4 | !hbusreq3 & v9ea5a6;
assign v9f76e0 = stateG2_p & v845542 | !stateG2_p & v9f76df;
assign v9f785b = hbusreq0_p & v9f772a | !hbusreq0_p & v9f772b;
assign b57ab6 = hmaster1_p & b57ab5 | !hmaster1_p & v845542;
assign dc505b = hgrant4_p & ade572 | !hgrant4_p & !ade563;
assign b058a6 = hmastlock_p & b058a5 | !hmastlock_p & v845542;
assign d358ef = hburst0 & d358eb | !hburst0 & d358ee;
assign ac1450 = hmaster0_p & ac144f | !hmaster0_p & v845542;
assign v9e9f83 = hbusreq1_p & v9e9f57 | !hbusreq1_p & v9e9f79;
assign b1c7c0 = hbusreq4_p & b1c7bd | !hbusreq4_p & !b1c7bf;
assign b1c035 = hbusreq1_p & b1c768 | !hbusreq1_p & b1c034;
assign b1c854 = hgrant2_p & v845542 | !hgrant2_p & b1c853;
assign ad4dca = hbusreq3 & ad4dc9 | !hbusreq3 & v845542;
assign bd5933 = hlock0_p & dc538c | !hlock0_p & bd5932;
assign bd5b7f = hmastlock_p & adea97 | !hmastlock_p & !d359b4;
assign c3d715 = hmaster0_p & c3d70a | !hmaster0_p & c3d714;
assign bd57fd = hgrant0_p & c3d669 | !hgrant0_p & bd57fb;
assign ad4fe0 = hmaster2_p & ad4fd8 | !hmaster2_p & ad4fdf;
assign bd57cf = hbusreq1 & bd57c5 | !hbusreq1 & bd57c7;
assign d354aa = hmaster2_p & d354a9 | !hmaster2_p & d354a6;
assign ac145e = hlock1_p & ac144f | !hlock1_p & cc36b8;
assign ad4436 = hbusreq1_p & ad4435 | !hbusreq1_p & v845547;
assign ad4f3a = hmaster2_p & v84556c | !hmaster2_p & ad4f39;
assign v9f76bb = hmaster1_p & v9f76ba | !hmaster1_p & v9f7ce9;
assign b1c083 = stateG10_4_p & b1c066 | !stateG10_4_p & b1c082;
assign v9f77f0 = stateG10_4_p & v9f77ee | !stateG10_4_p & !v9f77ef;
assign bd5ba8 = hready_p & v845542 | !hready_p & bd5ba7;
assign ad4f45 = hbusreq1_p & ad4f44 | !hbusreq1_p & v84556c;
assign v9ea5e6 = hgrant2_p & v9ea5e4 | !hgrant2_p & v9ea5e5;
assign dc507c = hgrant1_p & dc507b | !hgrant1_p & dc502d;
assign c3d520 = decide_p & c3d482 | !decide_p & !c3d51f;
assign ad502e = hmastlock_p & d35a3a | !hmastlock_p & !v845542;
assign v9f7cc7 = locked_p & v9f7c9f | !locked_p & v9f7cc6;
assign b1c05b = hbusreq2 & b1c80d | !hbusreq2 & !b1c80a;
assign v9f7d9f = hbusreq2 & v9f7d9d | !hbusreq2 & v9f7d9e;
assign c5c89b = hlock4_p & c5c88d | !hlock4_p & !v845542;
assign c3cdfb = hmaster1_p & c3cdf9 | !hmaster1_p & c3cdfa;
assign b1c766 = hlock1_p & b1c760 | !hlock1_p & b1c765;
assign ad46f8 = hmaster1_p & ad46f7 | !hmaster1_p & ad46e4;
assign ade5b7 = hgrant2_p & ade5b0 | !hgrant2_p & ade5b6;
assign dc4f85 = hbusreq3 & dc4f6f | !hbusreq3 & v845542;
assign ad445b = hgrant4_p & ad4382 | !hgrant4_p & v845542;
assign ade5c6 = hmaster1_p & ade5c5 | !hmaster1_p & ade5c2;
assign bd5900 = decide_p & bd58ff | !decide_p & v845572;
assign ad43d7 = hbusreq2 & ad43cd | !hbusreq2 & ad43d3;
assign dc5302 = hmaster2_p & adec93 | !hmaster2_p & !dc5301;
assign v9e9eb1 = hbusreq1_p & v9e9eb0 | !hbusreq1_p & v9ea4b4;
assign v9ea412 = stateG2_p & v845542 | !stateG2_p & v9ea411;
assign d356a7 = hlock1_p & d356a6 | !hlock1_p & d355a9;
assign c3d69d = hmaster0_p & c3d696 | !hmaster0_p & c3d699;
assign v9f766e = hbusreq1 & v9f766c | !hbusreq1 & v9f766d;
assign ad40f3 = hbusreq2 & ad5012 | !hbusreq2 & v845547;
assign c3ce32 = jx1_p & c3d58a | !jx1_p & c3ce31;
assign v8cc4b4 = hbusreq1 & v8cc482 | !hbusreq1 & v8cc483;
assign b57a78 = hbusreq4 & b57a77 | !hbusreq4 & b579ce;
assign c3d747 = hbusreq1_p & c3d6b1 | !hbusreq1_p & c3d744;
assign v9f76d3 = hmaster0_p & v9f7cee | !hmaster0_p & v9f7cb2;
assign d3595a = hmaster0_p & d35953 | !hmaster0_p & d35959;
assign ad48b0 = hmaster2_p & v845542 | !hmaster2_p & !ad4de2;
assign ad4de0 = hbusreq3 & ad4ddf | !hbusreq3 & !v845542;
assign v9e9fad = hlock2 & v9e9faa | !hlock2 & v9e9fac;
assign b57a33 = hready_p & b57a2e | !hready_p & b57a32;
assign v9e9eb7 = hmaster1_p & v9e9eb6 | !hmaster1_p & v9e9e77;
assign v9f7886 = hmaster2_p & v9f7885 | !hmaster2_p & v9f772f;
assign dc4f6c = hbusreq2 & dc4f69 | !hbusreq2 & dc4f6b;
assign bd5814 = hgrant4_p & v84556c | !hgrant4_p & bd57fe;
assign v8cc4f1 = hbusreq1_p & v8ccb76 | !hbusreq1_p & v8cc4ee;
assign dc4fcf = hbusreq3 & dc4fce | !hbusreq3 & v845542;
assign c74198 = stateG3_0_p & v845542 | !stateG3_0_p & !v845580;
assign b0594a = hmaster0_p & b058c5 | !hmaster0_p & b058b5;
assign ad4610 = decide_p & ad4606 | !decide_p & ad460f;
assign ade59a = hgrant0_p & ade572 | !hgrant0_p & !v84556c;
assign v8cc5a4 = hlock2 & v8cc489 | !hlock2 & v8cc5a0;
assign v8cc602 = hready_p & v8cc507 | !hready_p & v8cc601;
assign d35750 = hgrant1_p & v84554c | !hgrant1_p & d3574f;
assign v8cc5bd = hbusreq1 & v8cc598 | !hbusreq1 & v8cc599;
assign b5b408 = locked_p & b5b407 | !locked_p & v845542;
assign d35709 = hbusreq1_p & d35708 | !hbusreq1_p & v845542;
assign v9ea3f2 = hmaster0_p & v9f20a1 | !hmaster0_p & v9ea3e7;
assign c3d5ed = hbusreq2 & c3d5e6 | !hbusreq2 & c3d5ec;
assign ad43bf = decide_p & ad43a3 | !decide_p & ad43be;
assign v9ea47e = hbusreq0 & v9ea47c | !hbusreq0 & v9ea47d;
assign c5c9aa = decide_p & c5c8e0 | !decide_p & c5c9a9;
assign v8cc5b3 = hbusreq3 & v8cc5b1 | !hbusreq3 & v8cc5b2;
assign cc36b8 = hmaster2_p & v845542 | !hmaster2_p & !v84556c;
assign d3572b = hbusreq1_p & d356cb | !hbusreq1_p & v845542;
assign v9f7815 = hgrant2_p & v9f77bc | !hgrant2_p & v9f7814;
assign b058ce = hbusreq4_p & b058b6 | !hbusreq4_p & v9f7d42;
assign ade666 = jx0_p & ade662 | !jx0_p & ade665;
assign bd5907 = hbusreq1 & bd5b6f | !hbusreq1 & v845564;
assign b05a26 = hmaster0_p & b05a0e | !hmaster0_p & b05a25;
assign c3d710 = hmaster1_p & c3d70a | !hmaster1_p & c3d70f;
assign v9ea47f = hlock4 & v9ea476 | !hlock4 & v9ea47e;
assign ad45eb = hlock0_p & ade4c1 | !hlock0_p & !v845542;
assign ad4fed = hbusreq3 & ad4fec | !hbusreq3 & v845542;
assign dc53bc = hmaster1_p & dc53bb | !hmaster1_p & v84556c;
assign b57ae0 = decide_p & b57adf | !decide_p & b57944;
assign b1c7dc = hgrant4_p & b1c7b6 | !hgrant4_p & b1c7bc;
assign c3d692 = hmaster1_p & c3d683 | !hmaster1_p & c3d68b;
assign ad42f8 = hgrant1_p & v845542 | !hgrant1_p & ad42f7;
assign c3d707 = hmaster0_p & c3d697 | !hmaster0_p & c3d696;
assign b059b8 = hbusreq1 & b059b6 | !hbusreq1 & b059b7;
assign d35755 = hmaster0_p & d35752 | !hmaster0_p & d35754;
assign df51cb = decide_p & df51b7 | !decide_p & d6ebca;
assign ad4eac = hbusreq1 & ad4e95 | !hbusreq1 & !v845547;
assign ac146a = hmaster2_p & ac1464 | !hmaster2_p & !ac1469;
assign b1cc01 = hgrant1_p & v845542 | !hgrant1_p & b1cc00;
assign ad477d = hready & ad45e1 | !hready & ad477c;
assign bd5888 = hmaster2_p & bd5883 | !hmaster2_p & bd5887;
assign c3d38d = hbusreq2 & c3d38b | !hbusreq2 & !v845542;
assign locked = d35028;
assign c3d2b9 = hmaster0_p & c3d2b3 | !hmaster0_p & c3d2b8;
assign d354d7 = hbusreq2 & d35c01 | !hbusreq2 & !d35c03;
assign c3d6cb = hlock0_p & c3d6c7 | !hlock0_p & c3d6ca;
assign c3ce55 = hbusreq1_p & c3ce54 | !hbusreq1_p & c3d305;
assign b57437 = hbusreq1_p & b57942 | !hbusreq1_p & b579bb;
assign ad4fd5 = hgrant4_p & ad4fae | !hgrant4_p & v84556c;
assign ad43d2 = hbusreq0 & ad43d1 | !hbusreq0 & !v845542;
assign d35748 = hbusreq2 & d3572b | !hbusreq2 & !d35aa4;
assign df5185 = hmaster0_p & df517f | !hmaster0_p & df5184;
assign b1cfc3 = hmaster2_p & b1cfbf | !hmaster2_p & b1cfc2;
assign ad4f71 = hbusreq4_p & ad4f6e | !hbusreq4_p & ad4f70;
assign v8cc4a1 = hmaster2_p & v8cc4a0 | !hmaster2_p & v8cc493;
assign v9f7d4c = hmaster0_p & v9f7d3b | !hmaster0_p & v9f7d3e;
assign c3d2ef = hgrant0_p & v845542 | !hgrant0_p & !c3d2e9;
assign v9ea588 = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea587;
assign d356f5 = hbusreq1_p & d356f4 | !hbusreq1_p & v845542;
assign d3571a = hmaster1_p & d35719 | !hmaster1_p & d35713;
assign v8cc0d1 = hbusreq1_p & v8ccbd8 | !hbusreq1_p & v8cc0d0;
assign c3d688 = hbusreq0_p & c3d66d | !hbusreq0_p & !c3d674;
assign c3d397 = hmaster1_p & c3d306 | !hmaster1_p & c3d396;
assign v9f76dd = hmaster1_p & v9f76dc | !hmaster1_p & v9f7d2f;
assign ad447b = hbusreq4_p & ad4479 | !hbusreq4_p & ad447a;
assign b058d7 = hbusreq0 & b058d1 | !hbusreq0 & b058d6;
assign df515c = hmaster0_p & df515a | !hmaster0_p & df515b;
assign dc5043 = hgrant4_p & ade56d | !hgrant4_p & !ade563;
assign ad431a = hbusreq1_p & ad4319 | !hbusreq1_p & v845542;
assign b1cf2e = hmaster0_p & v845542 | !hmaster0_p & b1cf2d;
assign df54da = hmaster0_p & df54d9 | !hmaster0_p & v845542;
assign v9ea5b3 = hmaster1_p & v9ea5b2 | !hmaster1_p & v9ea583;
assign v9e9edd = hready_p & v9ea3e3 | !hready_p & v9e9edc;
assign b1c742 = hmaster2_p & b1c741 | !hmaster2_p & v845542;
assign dc5005 = stateG10_4_p & ade563 | !stateG10_4_p & dc5004;
assign v9f7d4e = hbusreq2_p & v9f7d4b | !hbusreq2_p & v9f7d4d;
assign cc36fd = hbusreq0_p & v84556c | !hbusreq0_p & cc36fc;
assign ad4396 = hbusreq4_p & b1c714 | !hbusreq4_p & ad4380;
assign d35a4f = locked_p & d35a4e | !locked_p & v845542;
assign ad416a = hbusreq2 & ad4fec | !hbusreq2 & v845542;
assign ad4fc3 = hgrant1_p & ad4fb3 | !hgrant1_p & ad4fc2;
assign b1c70d = jx1_p & b1c703 | !jx1_p & b1c70c;
assign c3d32e = hbusreq4 & c3d303 | !hbusreq4 & !c3d32d;
assign v9ea5cf = hbusreq4 & v9ea5ce | !hbusreq4 & v9ea5cb;
assign c3ce6d = hbusreq1_p & c3ce6c | !hbusreq1_p & c3d2de;
assign d35be9 = hlock4_p & d359c1 | !hlock4_p & d35a4f;
assign c3cf1e = hmaster0_p & c3cf1c | !hmaster0_p & c3cf1d;
assign ad4ec5 = hbusreq4 & ad4ec3 | !hbusreq4 & ad4ec4;
assign c3d354 = hbusreq3 & c3d353 | !hbusreq3 & c3d32f;
assign b1c7e1 = hbusreq4 & b1c7d6 | !hbusreq4 & b1c7e0;
assign c3d345 = hbusreq0 & c3d342 | !hbusreq0 & c3d344;
assign b57ab7 = decide_p & b57a21 | !decide_p & b57ab6;
assign b57955 = hmaster2_p & b57951 | !hmaster2_p & b57954;
assign d35528 = hmaster2_p & d35a9b | !hmaster2_p & d35527;
assign v8cc5b4 = hlock2 & v8cc4ad | !hlock2 & v8cc5b3;
assign dc4fdc = hmaster0_p & dc4fd7 | !hmaster0_p & dc4fdb;
assign c3d751 = hmaster1_p & c3d750 | !hmaster1_p & c3d67c;
assign ade4ae = hbusreq3 & ade4ac | !hbusreq3 & ade4ad;
assign v8cc4b2 = hmaster1_p & v8cc475 | !hmaster1_p & v8cc4b1;
assign ba7c7f = jx1_p & ba7c7e | !jx1_p & ba7c75;
assign v9e9ea5 = hbusreq1_p & v9e9ea4 | !hbusreq1_p & v9ea4d9;
assign c3d5a9 = hbusreq1 & c3d5a0 | !hbusreq1 & c3d5a2;
assign b1c85e = hbusreq4_p & b1cfcc | !hbusreq4_p & !b1c85d;
assign v9ea46d = hmaster2_p & v9ea467 | !hmaster2_p & v9ea46c;
assign b058dc = hbusreq1 & b058da | !hbusreq1 & b058db;
assign ad4fd3 = hgrant1_p & ad4fd1 | !hgrant1_p & ad4fd2;
assign ad48b7 = hbusreq1_p & ad48b6 | !hbusreq1_p & v845542;
assign ade5d7 = hmaster2_p & adeaae | !hmaster2_p & ade5d6;
assign v9e9ec0 = hready_p & v9ea436 | !hready_p & v9e9ebf;
assign v9f20a1 = hmastlock_p & b06719 | !hmastlock_p & v845542;
assign b1c7cb = hgrant1_p & b1c7ba | !hgrant1_p & b1c7ca;
assign ad5036 = hbusreq1 & ad5026 | !hbusreq1 & ad5029;
assign bd592a = hlock2_p & bd5929 | !hlock2_p & v845542;
assign ad42b2 = hmaster2_p & ad42b0 | !hmaster2_p & ad45e6;
assign b1c61a = hmaster1_p & v845542 | !hmaster1_p & b1c619;
assign c3d2f5 = hgrant4_p & v845542 | !hgrant4_p & !c3d2ea;
assign dc5390 = hmaster1_p & dc538f | !hmaster1_p & v84556c;
assign c3d72f = hbusreq2_p & c3d72c | !hbusreq2_p & c3d72e;
assign c3ce39 = hbusreq2 & c3ce35 | !hbusreq2 & c3ce37;
assign b1c058 = hbusreq2 & b1c808 | !hbusreq2 & !b1c80a;
assign ad4807 = hready & ad4e4b | !hready & df54f5;
assign v9f77e4 = hbusreq3 & v9f77e0 | !hbusreq3 & v9f77e3;
assign b1c057 = hlock2_p & b1c052 | !hlock2_p & b1c056;
assign v9f76fa = hbusreq1_p & v9f7dbb | !hbusreq1_p & v9f76f9;
assign d35799 = hbusreq0 & d35798 | !hbusreq0 & v845542;
assign ad43dd = hready & ad43dc | !hready & !v845549;
assign d35792 = hlock0_p & v845542 | !hlock0_p & !dc539e;
assign c3d6d8 = hlock2_p & c3d6d4 | !hlock2_p & !c3d6d7;
assign bd58d0 = hbusreq4_p & dc505a | !hbusreq4_p & dc5010;
assign v8d29fb = hbusreq0_p & v8d29fa | !hbusreq0_p & v845542;
assign v9ea42b = hbusreq2_p & v9ea427 | !hbusreq2_p & v9ea42a;
assign c3d6a7 = hgrant4_p & c3d66a | !hgrant4_p & c3d6a6;
assign ad4607 = hbusreq4_p & ad5016 | !hbusreq4_p & v845542;
assign d35017 = hgrant1_p & d35016 | !hgrant1_p & d35014;
assign v9f7859 = hmaster1_p & v9f7858 | !hmaster1_p & v9f776d;
assign v8cc4fc = hbusreq4_p & v8ccbe2 | !hbusreq4_p & v8cc4fa;
assign b1cffe = hgrant0_p & bd5b93 | !hgrant0_p & v845542;
assign b578f6 = hburst1_p & v8b08c1 | !hburst1_p & !v9ea411;
assign c3d5ad = hlock2_p & c3d59a | !hlock2_p & !c3d5ac;
assign d3575a = hready_p & d35759 | !hready_p & d3573b;
assign bd5b6e = hburst0 & bd5b6a | !hburst0 & bd5b6d;
assign b1c806 = hbusreq3 & b1c803 | !hbusreq3 & !b1c805;
assign df51b2 = hbusreq3 & df5166 | !hbusreq3 & df5168;
assign ad44b3 = hbusreq4_p & v845542 | !hbusreq4_p & ad44b2;
assign v9f7e21 = hbusreq0 & v9f7e18 | !hbusreq0 & v9f7e20;
assign ad4da2 = hlock1_p & ad4da0 | !hlock1_p & ad4da1;
assign c3d533 = hbusreq2_p & c3d482 | !hbusreq2_p & c3d532;
assign c3d5f2 = hbusreq4 & c3d5ef | !hbusreq4 & !c3d5f1;
assign d35a78 = hgrant2_p & v845542 | !hgrant2_p & !d35a77;
assign c3d57a = hbusreq0 & c3d579 | !hbusreq0 & c3d4e2;
assign d35a3c = hmastlock_p & d35a3b | !hmastlock_p & !v845542;
assign c3d73c = hmaster1_p & c3d73b | !hmaster1_p & c3d68b;
assign b1c06e = hbusreq4_p & b1c7a4 | !hbusreq4_p & !b1c06d;
assign v8cc598 = hready & v8cc595 | !hready & v8ccbd8;
assign ba7c78 = hbusreq1_p & ba7c66 | !hbusreq1_p & ba7c64;
assign v9f77d4 = hbusreq2 & v9f77d2 | !hbusreq2 & v9f77d3;
assign v9f76c0 = hmaster0_p & v9f7d3e | !hmaster0_p & v9f7d3c;
assign c5c935 = hbusreq4_p & c5c8f9 | !hbusreq4_p & !c5c934;
assign v9f7685 = hmaster1_p & v9f7684 | !hmaster1_p & v9f7675;
assign b57989 = hmaster0_p & b57983 | !hmaster0_p & b57988;
assign v8cc43f = hgrant2_p & v8ccbde | !hgrant2_p & v8cc43d;
assign v9ea5db = hbusreq2_p & v9ea5d8 | !hbusreq2_p & v9ea5da;
assign v9ea467 = hbusreq4_p & v9ea462 | !hbusreq4_p & v9ea466;
assign c3ce8d = hbusreq2 & v845542 | !hbusreq2 & v845564;
assign d358ee = hburst1 & d358eb | !hburst1 & d358ed;
assign d356b8 = hmaster0_p & d356b4 | !hmaster0_p & d356b7;
assign b1c7d1 = hlock4_p & b1c7cf | !hlock4_p & b1c7d0;
assign ade5d1 = hbusreq2 & ade4c7 | !hbusreq2 & ade5d0;
assign c3ce47 = hbusreq1_p & c3ce46 | !hbusreq1_p & c3d305;
assign d355a9 = hmaster2_p & v84556c | !hmaster2_p & !d355a8;
assign b57987 = hmaster2_p & b57985 | !hmaster2_p & b57986;
assign v9f76a0 = hbusreq4_p & v9f769b | !hbusreq4_p & v9f769f;
assign v9e9ed2 = hmaster1_p & v9e9ed1 | !hmaster1_p & v9e9e77;
assign d357df = hmaster1_p & d357ce | !hmaster1_p & d357de;
assign c3d6b1 = hmaster2_p & c3d6aa | !hmaster2_p & c3d6b0;
assign df51b6 = hmaster1_p & df51b5 | !hmaster1_p & df5163;
assign d35900 = hmaster1_p & v845542 | !hmaster1_p & d358ff;
assign ade592 = hlock4_p & ade58e | !hlock4_p & !ade591;
assign ad4ef6 = hbusreq4_p & ad4ef5 | !hbusreq4_p & b1cfbe;
assign v9ea493 = hlock1 & v9ea43b | !hlock1 & v9ea492;
assign ad3d3a = hlock2_p & ad3d38 | !hlock2_p & ad3d39;
assign d35aae = hgrant1_p & v84554c | !hgrant1_p & d35aad;
assign c3cea1 = hbusreq3 & c3ce9d | !hbusreq3 & c3cea0;
assign ad4707 = hbusreq4_p & ad4fca | !hbusreq4_p & !v845542;
assign ad460b = hready & ad456f | !hready & !v845542;
assign d359f5 = hgrant0_p & d359c9 | !hgrant0_p & v845542;
assign v9f7738 = hmaster0_p & v9f772c | !hmaster0_p & v9f7730;
assign d35981 = hbusreq3 & d35980 | !hbusreq3 & v845542;
assign c5c974 = hmaster2_p & c5c8e7 | !hmaster2_p & !c5c92f;
assign c3d730 = decide_p & c3d72a | !decide_p & c3d72f;
assign bd582d = hmaster2_p & bd581c | !hmaster2_p & v845542;
assign v8cc5c1 = hbusreq2 & v8cc5c0 | !hbusreq2 & v8ccbd8;
assign v9f76b1 = hready_p & v9f7688 | !hready_p & !v9f76b0;
assign d3541c = hmaster2_p & d35419 | !hmaster2_p & d3541b;
assign ad4fb7 = hbusreq3 & ad4fb6 | !hbusreq3 & v845542;
assign d35502 = hbusreq1_p & v84555a | !hbusreq1_p & !d35501;
assign ad4f88 = hlock0_p & ad4f3e | !hlock0_p & !v845542;
assign ad4f2e = hbusreq3 & ad4f2d | !hbusreq3 & v845542;
assign d35576 = hmaster1_p & d35572 | !hmaster1_p & d35575;
assign ad435e = hmaster1_p & ad435d | !hmaster1_p & ad42e8;
assign d356e0 = hbusreq1 & d3590a | !hbusreq1 & v845542;
assign d356d8 = hlock1_p & d356d5 | !hlock1_p & d356d7;
assign bd576b = locked_p & bd576a | !locked_p & v845542;
assign c3d3a9 = hbusreq2_p & c3d398 | !hbusreq2_p & c3d3a8;
assign b1c047 = hbusreq1_p & b1c774 | !hbusreq1_p & b1c046;
assign ad3cc9 = hmaster1_p & ad3cc8 | !hmaster1_p & ad4419;
assign c3cef0 = stateG10_4_p & c3ceee | !stateG10_4_p & c3ceef;
assign ade4ef = hmaster0_p & ade4cf | !hmaster0_p & ade4ee;
assign ad4ea2 = hgrant4_p & v845542 | !hgrant4_p & ad4e98;
assign adec8b = hburst0_p & bb9c5a | !hburst0_p & !bbbcd9;
assign d3543c = hlock2_p & d35439 | !hlock2_p & d3543b;
assign df51a3 = hgrant3_p & df516e | !hgrant3_p & df51a2;
assign dc4f92 = hbusreq3 & dc4f91 | !hbusreq3 & v845542;
assign v9ea485 = hgrant1_p & v9ea404 | !hgrant1_p & v9ea484;
assign c3d47a = hbusreq4 & c3d2b5 | !hbusreq4 & !v845542;
assign v9f7cd3 = hbusreq3 & v9f7cd0 | !hbusreq3 & v9f7cd2;
assign df5173 = hbusreq1_p & df5172 | !hbusreq1_p & v845542;
assign ad3d21 = hgrant3_p & ad441f | !hgrant3_p & ad3d20;
assign c5c898 = hmaster2_p & c5c896 | !hmaster2_p & !v845542;
assign b05a0f = hmaster2_p & b05939 | !hmaster2_p & !b058a7;
assign bd58b0 = hbusreq2 & bd58af | !hbusreq2 & v845542;
assign b059da = hlock0_p & b0597e | !hlock0_p & b059d9;
assign ad4155 = hgrant4_p & v845542 | !hgrant4_p & ad4f3e;
assign c5c967 = hmastlock_p & c5c966 | !hmastlock_p & !v845542;
assign d35a68 = hbusreq4_p & d35a67 | !hbusreq4_p & !d35a66;
assign v8cc0d5 = hlock2 & v8cc489 | !hlock2 & v8cc0d4;
assign v9f7ced = hlock2 & v9f7cc8 | !hlock2 & v9f7cec;
assign d358ff = hmaster0_p & d358fe | !hmaster0_p & v845542;
assign ad415b = hmaster2_p & ad4159 | !hmaster2_p & ad4156;
assign d356de = hbusreq2 & d356d4 | !hbusreq2 & d356dd;
assign ad3d51 = hmaster0_p & ad3d50 | !hmaster0_p & ad3cdb;
assign ad4f4a = hlock0_p & v845542 | !hlock0_p & ad4f49;
assign d35442 = hbusreq2_p & d35441 | !hbusreq2_p & d35440;
assign c3d587 = decide_p & c3d533 | !decide_p & !c3d51f;
assign d357b2 = decide_p & d357b1 | !decide_p & v84556c;
assign b57429 = hlock2 & b57988 | !hlock2 & b57428;
assign b1c56e = decide_p & b1c56d | !decide_p & b1c866;
assign ad4de1 = hmaster2_p & v845542 | !hmaster2_p & !c74b29;
assign d354ce = hlock4_p & d35a13 | !hlock4_p & !d35a66;
assign dc500b = stateG10_4_p & adec89 | !stateG10_4_p & !dc500a;
assign v9ea478 = stateG10_4_p & v9ea464 | !stateG10_4_p & v9ea477;
assign c3cf23 = hbusreq2_p & c3ceea | !hbusreq2_p & c3cf22;
assign c3d47f = hmaster0_p & c3d47d | !hmaster0_p & c3d47e;
assign v9f7c9c = locked_p & v9f7c98 | !locked_p & v9f7c9b;
assign ad4da9 = hbusreq4_p & ad4da8 | !hbusreq4_p & v845542;
assign ac1472 = hbusreq2_p & ac1470 | !hbusreq2_p & ac146f;
assign ad4310 = hbusreq2_p & ad4303 | !hbusreq2_p & !ad430f;
assign ad4efe = hlock4_p & ad4efd | !hlock4_p & !v845576;
assign v8cc5aa = hbusreq4 & v8cc5a9 | !hbusreq4 & v8cc494;
assign b059b9 = hgrant1_p & b058c1 | !hgrant1_p & b059b8;
assign d35730 = hbusreq1_p & d356c7 | !hbusreq1_p & !v845542;
assign ade56b = hburst1 & v889629 | !hburst1 & !v845542;
assign c5c938 = hlock0_p & c5c8fc | !hlock0_p & c5c937;
assign v9f77bc = hmaster1_p & v9f77bb | !hmaster1_p & v9f7736;
assign ad429f = hbusreq1 & ad429e | !hbusreq1 & !v845542;
assign c3d2d8 = hbusreq3 & c3d2d6 | !hbusreq3 & v845564;
assign v8cc758 = hbusreq1_p & v8cc757 | !hbusreq1_p & v8cc494;
assign c76647 = start_p & v845542 | !start_p & !c76645;
assign ad4ee7 = hbusreq4_p & ad4ee4 | !hbusreq4_p & ad4ee6;
assign c3d679 = hbusreq0_p & c3d670 | !hbusreq0_p & c3d675;
assign c3ce68 = hbusreq2 & c3ce61 | !hbusreq2 & c3ce66;
assign v9f7d0d = hlock3 & v9f7d05 | !hlock3 & v9f7d0c;
assign b05a9a = hgrant3_p & b05a4c | !hgrant3_p & b05a99;
assign b059c9 = hlock1 & b058a8 | !hlock1 & b059c8;
assign v9ea423 = hmaster2_p & v9ea41b | !hmaster2_p & v9ea422;
assign v8cc7bf = hgrant4_p & v845542 | !hgrant4_p & v8cc7bd;
assign dc53e0 = jx2_p & dc53b7 | !jx2_p & dc53df;
assign c3d6fd = hmaster1_p & c3d6e8 | !hmaster1_p & c3d6fc;
assign b058e5 = hbusreq2_p & b058e2 | !hbusreq2_p & b058e4;
assign ad43cd = hready & ad43c8 | !hready & !ad43cc;
assign d35a9e = hbusreq1_p & d35a95 | !hbusreq1_p & d35a9d;
assign v9f7788 = hbusreq0 & v9f7786 | !hbusreq0 & v9f7787;
assign v8cc59e = hgrant1_p & v8cc59c | !hgrant1_p & v8cc474;
assign d3570e = hbusreq2 & d356c0 | !hbusreq2 & !v84554e;
assign ade4c4 = hburst1 & ade4c2 | !hburst1 & ade4c3;
assign v9f7790 = hbusreq2 & v9f778e | !hbusreq2 & v9f778f;
assign d359f2 = hgrant4_p & d359c9 | !hgrant4_p & d359ce;
assign ad3d60 = jx2_p & ad4263 | !jx2_p & ad3d5f;
assign bd58f2 = hlock2_p & bd58f1 | !hlock2_p & !bd57eb;
assign ade4a7 = hbusreq1_p & adec8a | !hbusreq1_p & ade4a6;
assign d35574 = hbusreq2 & d35500 | !hbusreq2 & d35502;
assign ad437b = jx1_p & ad437a | !jx1_p & v845542;
assign v9f7797 = hbusreq1 & v9f7795 | !hbusreq1 & v9f7796;
assign ad4f10 = hmaster2_p & ad4f0d | !hmaster2_p & ad4f0f;
assign c3d66f = hmaster2_p & c3d66a | !hmaster2_p & !c3d66e;
assign c5c8f5 = hgrant1_p & v845542 | !hgrant1_p & c5c8f4;
assign b05991 = hbusreq4_p & b0598f | !hbusreq4_p & !b05990;
assign adea88 = hmastlock_p & adea87 | !hmastlock_p & !v845542;
assign b1c6cf = hgrant3_p & b1c61c | !hgrant3_p & b1c6ce;
assign ad46ea = hbusreq2 & ad458c | !hbusreq2 & !v845542;
assign c3d5f4 = hgrant1_p & v84554d | !hgrant1_p & c3d5f3;
assign v9f7df4 = hbusreq3 & v9f7def | !hbusreq3 & v9f7df3;
assign d35a14 = stateG10_4_p & d35a03 | !stateG10_4_p & d35a13;
assign df513b = locked_p & df513a | !locked_p & !v845542;
assign df512b = hbusreq2_p & df512a | !hbusreq2_p & df5537;
assign ade5b0 = hmaster1_p & ade5a9 | !hmaster1_p & ade5af;
assign b1cafd = hmaster0_p & v845542 | !hmaster0_p & b1caf9;
assign b1c0b3 = jx1_p & b1c092 | !jx1_p & b1c0b2;
assign v9e9fbe = decide_p & v9ea4b2 | !decide_p & v9e9fbd;
assign ade4bd = hmastlock_p & ade4bc | !hmastlock_p & !v845542;
assign b1c077 = hbusreq1 & b1c802 | !hbusreq1 & !b1c804;
assign v9e9fcf = hready_p & v9ea3e3 | !hready_p & v9e9fce;
assign bd57c7 = hmaster2_p & bd57c4 | !hmaster2_p & ade4cc;
assign b05998 = hlock1 & b05992 | !hlock1 & b05997;
assign v9f7d03 = hbusreq2 & v9f7d01 | !hbusreq2 & v9f7d02;
assign v9f77cd = hlock1 & v9f77c8 | !hlock1 & v9f77cc;
assign d354df = hbusreq2 & d354bd | !hbusreq2 & !v84555a;
assign b1c092 = hbusreq3_p & b1c7fe | !hbusreq3_p & b1c091;
assign ad4f37 = hmaster2_p & v84556c | !hmaster2_p & ad4f36;
assign ba7c66 = hmaster2_p & ba7c65 | !hmaster2_p & ba7c64;
assign v8cc48e = hgrant4_p & v8d2b2b | !hgrant4_p & v845542;
assign ad4e89 = hgrant4_p & v845542 | !hgrant4_p & b1cfb6;
assign b05987 = hgrant4_p & b058a9 | !hgrant4_p & !v9ea3e9;
assign ad430e = hmaster1_p & ad430d | !hmaster1_p & ad42f9;
assign ad42d3 = hbusreq1_p & ad42d2 | !hbusreq1_p & v845547;
assign b1c7a0 = stateG10_4_p & b1c79d | !stateG10_4_p & !b1c79f;
assign b1c714 = hlock0_p & v84556c | !hlock0_p & b1c70e;
assign df519e = hgrant2_p & df5198 | !hgrant2_p & !df519d;
assign ad46a9 = hlock4_p & ad46a8 | !hlock4_p & v845542;
assign c3d37b = hbusreq3 & c3d37a | !hbusreq3 & v845542;
assign ad3d1b = hmaster0_p & ad3cda | !hmaster0_p & ad3d1a;
assign ad477a = hmaster2_p & v845542 | !hmaster2_p & !ad4779;
assign d359d7 = hlock4_p & d359d5 | !hlock4_p & d359d6;
assign d359a1 = stateG10_4_p & v845542 | !stateG10_4_p & !d3599f;
assign dc5027 = hgrant4_p & v84556c | !hgrant4_p & adeca1;
assign v9ea4cf = hgrant1_p & v9ea4cd | !hgrant1_p & v9ea4ce;
assign d354dd = hgrant2_p & d354dc | !hgrant2_p & !d354d4;
assign b57af4 = hmaster1_p & b57af3 | !hmaster1_p & v845542;
assign ad4276 = hbusreq3 & ad4275 | !hbusreq3 & v845542;
assign v9f7e2f = locked_p & v9f7e2e | !locked_p & !v9f7c9f;
assign c3d73e = hgrant0_p & c3d669 | !hgrant0_p & c3d73d;
assign ad43f4 = hmaster2_p & ad43f3 | !hmaster2_p & v845542;
assign ad40f8 = hmaster1_p & ad40f4 | !hmaster1_p & ad40f7;
assign b579dc = hlock0 & b579ce | !hlock0 & b579d9;
assign v9f7735 = hmaster2_p & v9f7732 | !hmaster2_p & v9f7734;
assign ad4337 = hmaster0_p & ad4335 | !hmaster0_p & ad4336;
assign b1c04a = hbusreq2_p & b1c02d | !hbusreq2_p & b1c049;
assign v9ea61d = hmaster1_p & v9ea61c | !hmaster1_p & v9ea3f0;
assign ad4584 = hbusreq2_p & ad4580 | !hbusreq2_p & ad4583;
assign d35918 = hlock0_p & d3590d | !hlock0_p & !v845542;
assign c3cec9 = hbusreq4_p & v845576 | !hbusreq4_p & c3cec8;
assign ad41b1 = hmaster1_p & ad41b0 | !hmaster1_p & ad4825;
assign bd591e = decide_p & bd591d | !decide_p & v845572;
assign b1c57b = hbusreq4_p & b1caeb | !hbusreq4_p & !v845542;
assign ad441d = hbusreq2_p & ad441a | !hbusreq2_p & ad441c;
assign ad45c9 = hready & ad45c5 | !hready & !ad45c8;
assign b57417 = hgrant4_p & b57408 | !hgrant4_p & v845542;
assign d356ed = hmaster1_p & d356e2 | !hmaster1_p & d356e5;
assign v9f77b5 = hbusreq2 & v9f77b3 | !hbusreq2 & v9f77b4;
assign ad4f7a = hbusreq4_p & ad4f79 | !hbusreq4_p & ad4f36;
assign bd58d6 = hmaster0_p & bd58b9 | !hmaster0_p & bd58d5;
assign b578fb = hlock1_p & b578f9 | !hlock1_p & b578fa;
assign ad4eed = hmaster2_p & ad4eeb | !hmaster2_p & ad4eec;
assign b1c589 = hbusreq3_p & b1c45e | !hbusreq3_p & b1c588;
assign c3d340 = hbusreq0 & c3d33a | !hbusreq0 & c3d33f;
assign b579e9 = hmaster0_p & b579c8 | !hmaster0_p & b579e8;
assign bd58a4 = hgrant0_p & v845542 | !hgrant0_p & bd58a2;
assign v9f7da6 = hlock4 & v9f7da3 | !hlock4 & v9f7da5;
assign b059b3 = hbusreq0 & b059b1 | !hbusreq0 & b059b2;
assign bd5836 = hburst1 & c3d673 | !hburst1 & !v845542;
assign c3d69f = hbusreq2_p & c3d69c | !hbusreq2_p & c3d69e;
assign bd5873 = hgrant0_p & ade572 | !hgrant0_p & !bd574e;
assign ad42dd = hbusreq2 & ad4272 | !hbusreq2 & v845542;
assign ad474f = hmaster1_p & ad4736 | !hmaster1_p & ad474e;
assign dc53c4 = hlock3_p & dc53c3 | !hlock3_p & v845542;
assign c3d2f8 = hmaster2_p & c3d2f7 | !hmaster2_p & v845542;
assign d35704 = hlock1_p & d356fe | !hlock1_p & d35703;
assign v8cc439 = hmaster2_p & v8cc437 | !hmaster2_p & v8cc438;
assign v9ea5be = hmaster1_p & v9ea567 | !hmaster1_p & v9ea56b;
assign ad419e = hbusreq2 & v845542 | !hbusreq2 & v845547;
assign ad4f0b = hmaster2_p & ad4f08 | !hmaster2_p & ad4f0a;
assign ad4361 = hgrant2_p & ad435e | !hgrant2_p & ad4360;
assign b1c7ef = hbusreq2 & b1c7b5 | !hbusreq2 & !b1c7b8;
assign b0594c = hlock1_p & b058c1 | !hlock1_p & b058fd;
assign d35719 = hmaster0_p & d3570e | !hmaster0_p & d35718;
assign c3d481 = hmaster0_p & c3d480 | !hmaster0_p & c3d2be;
assign b05946 = hmaster1_p & b05945 | !hmaster1_p & b05943;
assign df517d = hbusreq1 & dc4ff9 | !hbusreq1 & v845542;
assign v8cc787 = hlock2 & v8ccbd8 | !hlock2 & v8cc786;
assign d35a13 = hgrant4_p & v845542 | !hgrant4_p & d35a03;
assign c3d6ba = hgrant4_p & c3d674 | !hgrant4_p & c3d6b8;
assign b1c4c7 = hbusreq0 & b1c4c4 | !hbusreq0 & b1c4c6;
assign ad4dd6 = hmaster0_p & ad4dca | !hmaster0_p & ad4dd5;
assign v9f7813 = hgrant2_p & v9f77bc | !hgrant2_p & v9f7812;
assign c3cee8 = hbusreq1 & c3cee0 | !hbusreq1 & c3cee4;
assign ade61d = hmaster1_p & ade61c | !hmaster1_p & ade5af;
assign c3d59d = busreq_p & c5c88b | !busreq_p & v845542;
assign v9f78a0 = hgrant2_p & v9f7877 | !hgrant2_p & v9f789f;
assign b1c861 = hgrant1_p & b1d01a | !hgrant1_p & b1c860;
assign ad4706 = hgrant1_p & ad459e | !hgrant1_p & ad4705;
assign ad5022 = hgrant1_p & ad5012 | !hgrant1_p & ad5021;
assign b05900 = hlock2 & b058b8 | !hlock2 & b058ff;
assign c3d2bc = hbusreq0 & v845542 | !hbusreq0 & v845564;
assign c3d75e = hgrant2_p & c3d75c | !hgrant2_p & c3d75d;
assign v9f7cef = hmaster0_p & v9f7cb2 | !hmaster0_p & v9f7cee;
assign ad5029 = hready & ad4fc1 | !hready & !v845542;
assign v9f7c9a = stateA1_p & v845542 | !stateA1_p & !v9f7c99;
assign b05938 = hmastlock_p & b058a0 | !hmastlock_p & v845542;
assign c3d736 = hgrant2_p & c3d733 | !hgrant2_p & c3d735;
assign d35495 = hmaster2_p & d35be3 | !hmaster2_p & d35494;
assign c3ce78 = hmaster0_p & c3ce76 | !hmaster0_p & c3ce77;
assign b574d1 = hgrant2_p & b579b0 | !hgrant2_p & b574d0;
assign b5794d = hbusreq1_p & b5794c | !hbusreq1_p & v845542;
assign b1c0b5 = jx2_p & b1c615 | !jx2_p & b1c0b4;
assign c3d579 = hmaster2_p & c3d578 | !hmaster2_p & v845542;
assign b574b1 = hbusreq0_p & b579ba | !hbusreq0_p & b57941;
assign d359fc = hbusreq4_p & d359fa | !hbusreq4_p & d359fb;
assign v9e9fc7 = hmaster1_p & v9e9fae | !hmaster1_p & v9e9f9f;
assign b05971 = hgrant1_p & b0596f | !hgrant1_p & b05970;
assign v9f775b = hlock0 & v9f775a | !hlock0 & v9f7759;
assign d3569e = hmaster2_p & d3597f | !hmaster2_p & d359ef;
assign bd58cd = hgrant4_p & dc5050 | !hgrant4_p & v84556c;
assign b1cfc4 = hgrant0_p & bd5b88 | !hgrant0_p & !v845542;
assign b05a95 = hmaster1_p & b05a25 | !hmaster1_p & b05a20;
assign ad4370 = hgrant2_p & ad436d | !hgrant2_p & ad436f;
assign v8cc479 = hmastlock_p & v8cc476 | !hmastlock_p & v845542;
assign ad3d34 = hmaster0_p & ad3d33 | !hmaster0_p & ad4421;
assign d354e2 = hbusreq1 & d35bf2 | !hbusreq1 & d35be8;
assign b1c84b = hmaster1_p & b1c842 | !hmaster1_p & b1c84a;
assign bcd5a7 = hbusreq3_p & v845542 | !hbusreq3_p & v845574;
assign v9e9f94 = hlock4 & v9e9f8e | !hlock4 & v9e9f93;
assign c3d720 = hbusreq2_p & c3d71d | !hbusreq2_p & c3d71f;
assign bb9c5a = start_p & v845542 | !start_p & bbbcd6;
assign b05a23 = hmaster0_p & b0593b | !hmaster0_p & b05a0f;
assign bd57bd = stateG2_p & v845542 | !stateG2_p & bd57bc;
assign v8cc501 = hgrant1_p & v8ccbe7 | !hgrant1_p & v8cc4fe;
assign d35444 = decide_p & d35443 | !decide_p & v84556c;
assign ad45e3 = hlock4_p & ad4dad | !hlock4_p & ad45e2;
assign ad43ca = hlock0_p & dc4f78 | !hlock0_p & ad43c9;
assign b1c781 = hmaster1_p & b1c780 | !hmaster1_p & b1c775;
assign ad4f65 = hlock4_p & ad4f64 | !hlock4_p & v845542;
assign c3d694 = hmaster1_p & c3d693 | !hmaster1_p & c3d68b;
assign ad4e71 = hgrant4_p & v84557a | !hgrant4_p & !ad4e6f;
assign b1c840 = hbusreq4_p & v845542 | !hbusreq4_p & d35aaa;
assign dc4f8e = hbusreq0 & dc4f75 | !hbusreq0 & dc4f8d;
assign ade58a = hgrant0_p & ade589 | !hgrant0_p & v84556c;
assign v9ea3f7 = hmaster1_p & v9ea3f6 | !hmaster1_p & v9ea3f0;
assign v9f772e = hmaster0_p & v9f772c | !hmaster0_p & v9f772d;
assign ad4e99 = hgrant4_p & v84556c | !hgrant4_p & ad4e98;
assign bd5861 = hgrant0_p & adec90 | !hgrant0_p & adec89;
assign v9f7db3 = hbusreq4_p & v9f7db1 | !hbusreq4_p & v9f7db2;
assign v9e9f4d = hgrant0_p & v9ea3e6 | !hgrant0_p & v9e9f4c;
assign b1c7a9 = hgrant4_p & v845542 | !hgrant4_p & b1c79d;
assign b05a7c = hgrant1_p & b0596f | !hgrant1_p & b05a7b;
assign dc4ff2 = hmaster2_p & dc4ff1 | !hmaster2_p & v845542;
assign v8cc62f = hmaster1_p & v8cc62e | !hmaster1_p & v845542;
assign v9f76b7 = hbusreq2_p & v9f76b4 | !hbusreq2_p & v9f76b6;
assign b1c820 = hbusreq3 & b1c81c | !hbusreq3 & !b1c81f;
assign v9f7e3f = hmaster2_p & v9f7e1b | !hmaster2_p & v9f7e3e;
assign d358fa = hmaster2_p & v845542 | !hmaster2_p & d358f9;
assign b1c4cc = hbusreq0 & b1c4c9 | !hbusreq0 & b1c4cb;
assign ad43fe = hbusreq2 & ad43db | !hbusreq2 & ad43dd;
assign dc4fe4 = hgrant4_p & c3d66d | !hgrant4_p & ade553;
assign c3ce04 = hbusreq2 & c3d35b | !hbusreq2 & c3d306;
assign c3ce4d = hgrant1_p & v84554d | !hgrant1_p & c3ce4c;
assign b0592a = hlock2_p & b05927 | !hlock2_p & b05929;
assign v9ea40c = hmaster0_p & v845542 | !hmaster0_p & v9ea3e1;
assign ad4697 = hbusreq4 & ad4696 | !hbusreq4 & v845542;
assign d354c5 = hbusreq1_p & d354b7 | !hbusreq1_p & d354c4;
assign bd57a1 = hbusreq1_p & bd579d | !hbusreq1_p & bd57a0;
assign ad470a = hbusreq4_p & ad4fce | !hbusreq4_p & !v845542;
assign ade5bf = hmaster0_p & ade5bd | !hmaster0_p & ade5be;
assign c3cf0c = hbusreq1_p & c3d2de | !hbusreq1_p & c3ce6a;
assign b1c775 = hmaster0_p & b1c76c | !hmaster0_p & !b1c774;
assign b57b58 = hready_p & b57a2e | !hready_p & b57b57;
assign v9f7dae = hlock0_p & v9f7dad | !hlock0_p & v9f7cc6;
assign d359ad = hmaster2_p & v84557a | !hmaster2_p & !v845542;
assign dc5050 = locked_p & dc504f | !locked_p & !v845542;
assign df5119 = hmaster0_p & df5118 | !hmaster0_p & v845542;
assign v9ea625 = hmaster1_p & v9ea624 | !hmaster1_p & v9ea405;
assign ad4ec4 = hbusreq0 & ad4e8a | !hbusreq0 & ad4e8e;
assign d357e4 = decide_p & d357e3 | !decide_p & v84556c;
assign v9f7cc6 = hmastlock_p & v9f7cc5 | !hmastlock_p & !v845542;
assign b57400 = decide_p & b57a21 | !decide_p & b573ff;
assign ad46c2 = hbusreq1_p & ad46ae | !hbusreq1_p & ad46c1;
assign v8cc7a5 = hmaster0_p & v8cc7a2 | !hmaster0_p & v845542;
assign ad4f9d = hbusreq3 & ad4f9c | !hbusreq3 & v845542;
assign ad42a4 = hlock1_p & ad42a2 | !hlock1_p & !ad42a3;
assign ad433d = hbusreq1 & ad5063 | !hbusreq1 & v845542;
assign v9ea435 = hgrant2_p & v9ea40d | !hgrant2_p & v9ea434;
assign bd57c0 = busreq_p & c5c88b | !busreq_p & !v845542;
assign c3d68c = hmaster1_p & c3d684 | !hmaster1_p & c3d68b;
assign ad4394 = hbusreq1_p & ad438f | !hbusreq1_p & ad4393;
assign bd5baf = decide_p & bd5bae | !decide_p & v845572;
assign v8cc499 = hgrant4_p & v845542 | !hgrant4_p & v8cc498;
assign d3594b = stateA1_p & e0edf9 | !stateA1_p & !d3594a;
assign d35902 = hgrant2_p & d35900 | !hgrant2_p & d358f6;
assign c3d6ad = hgrant4_p & c3d670 | !hgrant4_p & c3d6ac;
assign ad4433 = hgrant1_p & ad4428 | !hgrant1_p & ad4432;
assign c3d6a9 = stateG10_4_p & c3d6a6 | !stateG10_4_p & !c3d6a8;
assign cc3708 = decide_p & cc3707 | !decide_p & v84556c;
assign d359b0 = hbusreq1_p & d359af | !hbusreq1_p & !d359ae;
assign b579cd = hgrant4_p & v845542 | !hgrant4_p & b579cc;
assign c3ce2f = hready_p & c3ce2d | !hready_p & c3ce2e;
assign c3cf02 = hbusreq0 & c3cf01 | !hbusreq0 & v845564;
assign ad4eaa = hmaster0_p & ad4e93 | !hmaster0_p & ad4ea9;
assign b1c76e = hmaster2_p & b1c76d | !hmaster2_p & !b1cf29;
assign bd5917 = hbusreq1_p & bd5916 | !hbusreq1_p & v845542;
assign d35737 = hbusreq1_p & d356e3 | !hbusreq1_p & d35a9d;
assign d35aa4 = hbusreq1_p & v84554e | !hbusreq1_p & !v845542;
assign v9f7def = hgrant1_p & v9f7dc7 | !hgrant1_p & v9f7dee;
assign b1c770 = hbusreq0_p & dc4f7c | !hbusreq0_p & v845542;
assign ade5c8 = decide_p & ade5c7 | !decide_p & v845542;
assign ad4f78 = hbusreq4_p & ad4f65 | !hbusreq4_p & v845542;
assign v9ea44f = hlock0 & v9ea3fa | !hlock0 & v9ea44e;
assign b1c70c = hbusreq3_p & b1c709 | !hbusreq3_p & b1c86a;
assign v9f7667 = hmaster2_p & v9f7660 | !hmaster2_p & v9f7666;
assign ade5a4 = hmaster0_p & ade57e | !hmaster0_p & ade5a3;
assign ad40ff = hbusreq1_p & ad40fd | !hbusreq1_p & ad40fe;
assign dc505d = hbusreq4_p & dc505a | !hbusreq4_p & dc505c;
assign c3ce70 = hmaster1_p & c3ce69 | !hmaster1_p & c3ce6f;
assign ad503c = stateG10_4_p & cc36fc | !stateG10_4_p & !ad503b;
assign v9ea591 = hmaster2_p & v9ea444 | !hmaster2_p & v9ea590;
assign v9f7d3e = hmaster2_p & v9f7d3a | !hmaster2_p & !v9f7cc6;
assign ad480c = hready & v845542 | !hready & dc4fcb;
assign ad46a0 = hbusreq0 & ad469c | !hbusreq0 & ad469f;
assign c3d5d4 = hgrant0_p & v845542 | !hgrant0_p & !c3d5d3;
assign d355ac = hmaster1_p & d355ab | !hmaster1_p & v84556c;
assign dc4ff0 = stateG10_4_p & ade553 | !stateG10_4_p & !dc4fef;
assign v9f76d1 = decide_p & v9f76cb | !decide_p & !v9f76d0;
assign ad3ce4 = hbusreq0 & ad3ce3 | !hbusreq0 & !v845542;
assign ad4e55 = hmaster2_p & d3597f | !hmaster2_p & ad4e54;
assign b574c1 = stateG10_4_p & v845542 | !stateG10_4_p & b574c0;
assign bd5ea8 = hbusreq2_p & bd5ea7 | !hbusreq2_p & !v845542;
assign b57ad3 = hbusreq2_p & b57ad2 | !hbusreq2_p & b57904;
assign b1c098 = hgrant3_p & b1c705 | !hgrant3_p & b1c097;
assign dc53c9 = hgrant3_p & dc53c6 | !hgrant3_p & !dc53c8;
assign b57abd = stateA1_p & v9ea412 | !stateA1_p & b578f7;
assign c3ce24 = hready_p & c3ce0a | !hready_p & c3ce23;
assign ad4261 = hbusreq3_p & ad41ae | !hbusreq3_p & ad4260;
assign v9ea452 = hbusreq4 & v9ea450 | !hbusreq4 & v9ea451;
assign bd580a = hbusreq4_p & bd5807 | !hbusreq4_p & bd5809;
assign ad4ed4 = hgrant4_p & ad4eae | !hgrant4_p & ad4eb3;
assign v8cc58f = hbusreq4_p & v8cc47a | !hbusreq4_p & v8d2b2b;
assign bd5b8c = hmaster0_p & v84556c | !hmaster0_p & bd5b8b;
assign v8cc781 = hgrant2_p & v8cc76e | !hgrant2_p & v8cc761;
assign ad4338 = hbusreq1 & v845542 | !hbusreq1 & c3d2d9;
assign v9f7846 = hmaster0_p & v9f783d | !hmaster0_p & !v9f7845;
assign c3d30b = hmaster2_p & c3d2f2 | !hmaster2_p & c3d30a;
assign ade5b9 = decide_p & ade5b8 | !decide_p & adeaa7;
assign d3580b = hbusreq0_p & v84556c | !hbusreq0_p & !v845542;
assign d35a2b = hmaster1_p & d35a2a | !hmaster1_p & d35a25;
assign b05985 = hbusreq4_p & b05983 | !hbusreq4_p & !b05984;
assign ad4fb9 = hmaster1_p & ad4fb2 | !hmaster1_p & ad4fb8;
assign d3561e = hmaster2_p & dc5318 | !hmaster2_p & d3561d;
assign b5742d = hgrant2_p & b57948 | !hgrant2_p & b5742c;
assign bd57e0 = hbusreq2 & bd57df | !hbusreq2 & v845542;
assign v9f77eb = hgrant0_p & d359c4 | !hgrant0_p & !v845542;
assign v9f76c9 = hmaster0_p & v9f76c8 | !hmaster0_p & v9f7d46;
assign v9f780c = hgrant4_p & v9f7734 | !hgrant4_p & !v9f780b;
assign ad4f9a = hbusreq4 & ad4f8e | !hbusreq4 & ad4f99;
assign d35955 = hburst0 & df54dd | !hburst0 & d35954;
assign dc4fbd = hbusreq0 & dc4fad | !hbusreq0 & dc4fbc;
assign ad501d = hbusreq3 & ad501b | !hbusreq3 & v845542;
assign bd58ab = hbusreq4_p & v84556c | !hbusreq4_p & bd58aa;
assign v8cc7c3 = hlock4 & v8ccbf4 | !hlock4 & v8cc7c2;
assign d35995 = hgrant0_p & d3597f | !hgrant0_p & v845542;
assign c3d39e = hbusreq0 & c3d39d | !hbusreq0 & adeaa5;
assign b058b6 = locked_p & v9ea3e9 | !locked_p & v9f7d42;
assign ad3d53 = hgrant2_p & ad3d4f | !hgrant2_p & ad3d52;
assign d35809 = stateG10_4_p & d35807 | !stateG10_4_p & d35808;
assign v9f7cd6 = hbusreq4_p & v9f7cb4 | !hbusreq4_p & !v9f7c9f;
assign ad4ff7 = hmaster0_p & ad4fc0 | !hmaster0_p & ad4ff6;
assign b1c038 = hmaster2_p & b1c030 | !hmaster2_p & b1c037;
assign v8cc78b = decide_p & v8cc4f4 | !decide_p & v8cc78a;
assign b1c5f5 = decide_p & b1c5f3 | !decide_p & b1c5f4;
assign d357bd = hmaster0_p & d35778 | !hmaster0_p & d357bc;
assign df51c3 = hgrant1_p & df5538 | !hgrant1_p & !df519a;
assign bd5b78 = hmaster0_p & v845542 | !hmaster0_p & bd5b77;
assign v9f7677 = hgrant2_p & v9f7d6c | !hgrant2_p & v9f7676;
assign b05a1c = stateG10_4_p & b059e3 | !stateG10_4_p & b05a1b;
assign dc4fd4 = hmaster2_p & adec89 | !hmaster2_p & adeca1;
assign c3d39d = hmaster2_p & c3d39c | !hmaster2_p & v845542;
assign v9f7d84 = hgrant4_p & v9f7ca5 | !hgrant4_p & v9f7d83;
assign d356cf = hbusreq2_p & d356ca | !hbusreq2_p & d356ce;
assign v9f7ce7 = hlock2 & v9f7cdd | !hlock2 & v9f7ce6;
assign ad4ed9 = hbusreq0_p & v845542 | !hbusreq0_p & ad4ed8;
assign b57a2e = decide_p & b57a2d | !decide_p & b5798b;
assign bd5747 = hbusreq3 & bd5736 | !hbusreq3 & bd5746;
assign c3d329 = hbusreq0 & c3d325 | !hbusreq0 & c3d328;
assign ade4f1 = hbusreq2_p & ade4ed | !hbusreq2_p & ade4f0;
assign v9f7694 = hgrant0_p & v9f7d5d | !hgrant0_p & !v9f7cc6;
assign c3d2fc = hbusreq0 & v845542 | !hbusreq0 & c3d2fb;
assign ad4139 = hbusreq0 & ad4134 | !hbusreq0 & ad4138;
assign d3542c = hmaster2_p & d35419 | !hmaster2_p & v84555a;
assign v8ccbf9 = hgrant2_p & v8ccbde | !hgrant2_p & v8ccbf8;
assign b574fd = hgrant3_p & b57946 | !hgrant3_p & b574fc;
assign ad40f0 = hbusreq2_p & ad40ef | !hbusreq2_p & v845542;
assign d359a8 = hmaster2_p & d359a7 | !hmaster2_p & v845542;
assign ad4e80 = hbusreq0 & ad4e7d | !hbusreq0 & ad4e7f;
assign d3557c = hbusreq4_p & d354a8 | !hbusreq4_p & !d35aab;
assign v8cc7ce = hbusreq2 & v8cc7cc | !hbusreq2 & v8cc7cd;
assign v9f7895 = hlock3 & v9f77e2 | !hlock3 & v9f7894;
assign b57438 = hgrant1_p & b57437 | !hgrant1_p & b579b3;
assign ad472e = hbusreq4 & ad46fe | !hbusreq4 & v845542;
assign bd5811 = hbusreq4_p & bd580e | !hbusreq4_p & bd5810;
assign b0597e = hgrant0_p & b058a7 | !hgrant0_p & !v9f7d42;
assign ad42fe = hmaster0_p & ad42fc | !hmaster0_p & ad42fd;
assign ad46e5 = hmaster1_p & ad46af | !hmaster1_p & ad46e4;
assign ad44a8 = hbusreq0 & ad44a7 | !hbusreq0 & v845542;
assign ade549 = hbusreq1 & ade548 | !hbusreq1 & !v845558;
assign v8d29f9 = stateG2_p & v845542 | !stateG2_p & v8d29f8;
assign b0593e = hbusreq1_p & b0593b | !hbusreq1_p & b0593d;
assign df54e8 = hbusreq1_p & df54e7 | !hbusreq1_p & v845542;
assign ade623 = hmaster1_p & ade622 | !hmaster1_p & ade4ec;
assign ad428f = hlock3_p & ad4280 | !hlock3_p & !ad428e;
assign dc5393 = decide_p & dc5392 | !decide_p & v845542;
assign dc5016 = hbusreq3 & dc5015 | !hbusreq3 & v845542;
assign c3d35c = hbusreq3 & c3d35b | !hbusreq3 & c3d306;
assign ad45be = hmaster2_p & ad45bb | !hmaster2_p & !ad45bd;
assign d35a34 = hmaster1_p & d35a33 | !hmaster1_p & d35a1b;
assign bd5857 = hbusreq2 & bd5856 | !hbusreq2 & v845542;
assign v9f7d90 = hmaster2_p & v9f7d88 | !hmaster2_p & !v9f7d8f;
assign c5c8a1 = hmaster0_p & c5c897 | !hmaster0_p & c5c898;
assign v8ccbe2 = hgrant4_p & v845542 | !hgrant4_p & v8ccbe1;
assign d3556c = hmaster0_p & d3556b | !hmaster0_p & d354d7;
assign b059e5 = stateG10_4_p & b059e3 | !stateG10_4_p & !b059e4;
assign b1c5ee = hbusreq2 & b1c5ed | !hbusreq2 & b1d003;
assign cc36cd = hmaster2_p & cc36c9 | !hmaster2_p & cc36cc;
assign v9ea56f = hbusreq2_p & v9ea56c | !hbusreq2_p & v9ea56e;
assign ad45f9 = hmaster1_p & ad45c3 | !hmaster1_p & ad45f8;
assign ba7c6a = hready_p & v845558 | !hready_p & ba7c69;
assign df51aa = hmaster1_p & df51a6 | !hmaster1_p & df51a9;
assign d3559f = decide_p & d3559e | !decide_p & v84556c;
assign ad434d = hmaster0_p & ad434c | !hmaster0_p & ad4284;
assign bd5776 = hbusreq2 & bd5775 | !hbusreq2 & v845542;
assign b1c81c = hbusreq1_p & b1c743 | !hbusreq1_p & b1c81b;
assign c3d336 = hgrant0_p & v845542 | !hgrant0_p & c3d2e8;
assign v9f7e0a = hlock3 & v9f7e09 | !hlock3 & v9f7e06;
assign v8cc7d3 = hgrant2_p & v845542 | !hgrant2_p & v8cc7d0;
assign v9ea49d = hgrant2_p & v9ea499 | !hgrant2_p & v9ea49c;
assign bd5ea1 = hmaster2_p & adec93 | !hmaster2_p & !bd5ea0;
assign v9f7827 = hbusreq3 & v9f7825 | !hbusreq3 & v9f7826;
assign v9f77c1 = hbusreq4_p & v9f77bf | !hbusreq4_p & v9f77c0;
assign d3576f = hlock0_p & v845542 | !hlock0_p & d35a58;
assign b57a6b = hready & b57a6a | !hready & b57942;
assign b1c6c7 = hbusreq1_p & b1d00f | !hbusreq1_p & v8da59f;
assign v9f7ca9 = hbusreq0 & v9f7ca1 | !hbusreq0 & v9f7ca8;
assign b574c6 = hbusreq4 & b574c5 | !hbusreq4 & b579ce;
assign ade582 = hbusreq4_p & ade581 | !hbusreq4_p & v845542;
assign v8cc80d = hbusreq3 & v8cc7e6 | !hbusreq3 & v8cc80c;
assign v9f7db8 = hbusreq4 & v9f7db6 | !hbusreq4 & v9f7db7;
assign v9e9fd3 = hmaster1_p & v9ea49b | !hmaster1_p & v9e9fd0;
assign b1cff4 = hgrant0_p & dc52fa | !hgrant0_p & !v845542;
assign ad4593 = hbusreq3 & ad458b | !hbusreq3 & !v845542;
assign c3d302 = hgrant1_p & v84554d | !hgrant1_p & c3d301;
assign d3551e = hbusreq4_p & d35418 | !hbusreq4_p & v845548;
assign v9ea4ab = hbusreq4_p & v9f20a1 | !hbusreq4_p & !v9ea4aa;
assign v9f774f = hbusreq2 & v9f774d | !hbusreq2 & v9f774e;
assign d35774 = hlock0_p & v845542 | !hlock0_p & !d355a8;
assign v9f7d36 = hmaster1_p & v9f7d35 | !hmaster1_p & v9f7d2f;
assign c3d5b1 = hburst0 & c3d2e5 | !hburst0 & c3d2e6;
assign d356ac = hlock1_p & v845542 | !hlock1_p & v84556c;
assign d35c05 = hbusreq3 & d35c01 | !hbusreq3 & !v84555a;
assign d3568a = decide_p & d35689 | !decide_p & v84556c;
assign ad413c = hbusreq4_p & ad413b | !hbusreq4_p & ad4e9b;
assign b57ace = hgrant1_p & b57acd | !hgrant1_p & b578f9;
assign b1c6db = hmaster0_p & b1c842 | !hmaster0_p & b1c6da;
assign b0596b = hmaster2_p & b05952 | !hmaster2_p & v9f7d42;
assign adea97 = stateA1_p & v845542 | !stateA1_p & !adea96;
assign v9f7795 = hbusreq4 & v9f7793 | !hbusreq4 & v9f7794;
assign ad46ca = hbusreq4_p & ad4eef | !hbusreq4_p & v845542;
assign v8cc799 = hbusreq0 & v8cc797 | !hbusreq0 & v8cc798;
assign d35692 = hlock2_p & v845542 | !hlock2_p & d35691;
assign cc36d2 = hmaster0_p & v845542 | !hmaster0_p & cc36b8;
assign ad4f27 = hmaster0_p & ad4f19 | !hmaster0_p & ad4f26;
assign d35582 = hbusreq4 & d3557f | !hbusreq4 & d35581;
assign ad457e = hbusreq3 & ad457d | !hbusreq3 & v845542;
assign v8cc50d = hready_p & v8cc507 | !hready_p & v8cc50c;
assign ad40ba = hbusreq2 & ad48b7 | !hbusreq2 & !v845542;
assign v9ea4a8 = hmaster0_p & v9ea4a7 | !hmaster0_p & v9f20a1;
assign v9e9e77 = hmaster0_p & v9ea4b8 | !hmaster0_p & v9e9e76;
assign ad455c = hlock4_p & ad455b | !hlock4_p & v845542;
assign ba7c72 = hgrant3_p & ba7c6a | !hgrant3_p & ba7c71;
assign b058aa = hmaster2_p & b058a3 | !hmaster2_p & !b058a9;
assign bd5b71 = hbusreq2 & dc5394 | !hbusreq2 & bd5b70;
assign ad4dc0 = hlock2_p & ad4dba | !hlock2_p & ad4dbf;
assign b57406 = stateA1_p & b0ed8b | !stateA1_p & c74202;
assign ad4417 = hbusreq0 & ad4416 | !hbusreq0 & v845542;
assign ad4111 = hbusreq2 & ad4110 | !hbusreq2 & v845542;
assign d3578a = hlock0_p & v845542 | !hlock0_p & !dc5318;
assign adec92 = hmaster2_p & adec8a | !hmaster2_p & adec91;
assign c3ce3e = hbusreq1_p & c3ce3d | !hbusreq1_p & v84554d;
assign ad4802 = decide_p & ad47f7 | !decide_p & ad4801;
assign v9ea5d6 = hbusreq2 & v9ea5d4 | !hbusreq2 & v9ea5d5;
assign c5c8ec = hmaster1_p & c5c8ea | !hmaster1_p & c5c8eb;
assign b058af = hready & b058ae | !hready & b058aa;
assign ad4750 = hgrant2_p & ad472d | !hgrant2_p & ad474f;
assign ad4fdc = hlock0_p & ad4fd9 | !hlock0_p & ad4fdb;
assign c3ce17 = hbusreq2 & c3d2dd | !hbusreq2 & c3d2de;
assign ad4d8f = stateG2_p & v845542 | !stateG2_p & ad4d8e;
assign v9f7c94 = jx0_p & v85746a | !jx0_p & !v9f7c93;
assign dc506f = hmaster0_p & dc506b | !hmaster0_p & dc506e;
assign df54f5 = hmaster2_p & v84556c | !hmaster2_p & dc52fa;
assign b1cf49 = hready_p & v845542 | !hready_p & b1cf48;
assign ad4164 = hlock2_p & ad4149 | !hlock2_p & ad4163;
assign v9f77df = hbusreq1_p & v9f77ce | !hbusreq1_p & v9f77de;
assign b05a56 = hmaster0_p & b058c7 | !hmaster0_p & b058e8;
assign df5142 = hbusreq1_p & df5533 | !hbusreq1_p & v845542;
assign v9e9e6d = hbusreq2_p & v9e9e6c | !hbusreq2_p & v9ea4e1;
assign d3552f = hready_p & d35507 | !hready_p & !d3552e;
assign cc36cb = hlock4_p & v84556c | !hlock4_p & !cc36ca;
assign v8cc7a0 = hbusreq3 & v8cc79e | !hbusreq3 & v8cc79f;
assign v9ea580 = hmaster0_p & v9ea3fc | !hmaster0_p & v9ea3fa;
assign ad4eda = hlock0_p & ad4ed7 | !hlock0_p & ad4ed9;
assign dc53dd = hbusreq3_p & dc53dc | !hbusreq3_p & !dc5088;
assign bd5897 = hbusreq2 & bd5896 | !hbusreq2 & v845542;
assign ade63e = hready_p & v845542 | !hready_p & ade63d;
assign c3d596 = hmaster0_p & c3d594 | !hmaster0_p & c3d595;
assign ade550 = locked_p & ade54f | !locked_p & !v845542;
assign ad47f9 = hmaster1_p & ad47f8 | !hmaster1_p & ad45a5;
assign ad43f2 = hbusreq0 & ad43f1 | !hbusreq0 & v845542;
assign ade4c5 = hburst0 & ade4c2 | !hburst0 & ade4c4;
assign bd58c7 = hgrant4_p & v84556c | !hgrant4_p & bd58c6;
assign ad4e8f = hbusreq0 & ad4e8b | !hbusreq0 & ad4e8e;
assign v9f7dc9 = hgrant4_p & v9f7cf5 | !hgrant4_p & !v9f7d79;
assign v9ea3fe = locked_p & v845542 | !locked_p & v9ea3e6;
assign d35bf5 = hlock4_p & d3598a | !hlock4_p & v84556c;
assign bd5785 = hburst1 & bd5781 | !hburst1 & bd5784;
assign ade65f = decide_p & ade656 | !decide_p & adeaa7;
assign ad5050 = hbusreq0 & ad5045 | !hbusreq0 & ad504f;
assign bd587a = hmaster2_p & bd5870 | !hmaster2_p & bd5879;
assign b0598a = hbusreq4_p & b05989 | !hbusreq4_p & !b0597c;
assign bd5847 = hmaster2_p & bd580a | !hmaster2_p & bd5846;
assign v9f7ca2 = busreq_p & v9ea3e4 | !busreq_p & v9ea3e5;
assign d3598e = hmaster0_p & d35987 | !hmaster0_p & d3598d;
assign c3d5da = hgrant4_p & v845542 | !hgrant4_p & !c3d5d9;
assign v8cc0f0 = hbusreq3 & v8cc0ec | !hbusreq3 & v8cc0ee;
assign ad42b5 = hmaster2_p & ad42b4 | !hmaster2_p & ad45e2;
assign dc4f6f = hmaster2_p & ade4bf | !hmaster2_p & !ade4d4;
assign ade557 = hlock0_p & ade555 | !hlock0_p & !ade556;
assign bd57ee = hlock3_p & bd57e4 | !hlock3_p & bd57ed;
assign bd584b = stateG10_4_p & bd574e | !stateG10_4_p & !bd584a;
assign b57ac0 = hlock0 & b578f9 | !hlock0 & b57abf;
assign ad4425 = hmaster0_p & ad4423 | !hmaster0_p & ad4424;
assign c3ced7 = decide_p & c3ced6 | !decide_p & c3ce9a;
assign bd5752 = hbusreq3 & bd5750 | !hbusreq3 & v84556c;
assign v9f7d89 = hgrant0_p & v9f7cb6 | !hgrant0_p & v9ea3ec;
assign d359be = hmastlock_p & d359bd | !hmastlock_p & !v845542;
assign d35766 = hbusreq2_p & d35aa9 | !hbusreq2_p & !d35765;
assign df50d7 = hmaster2_p & v845542 | !hmaster2_p & df50d6;
assign bd5760 = hbusreq2 & bd575f | !hbusreq2 & v845542;
assign v8ccbf3 = hgrant4_p & v845542 | !hgrant4_p & v8ccbf2;
assign v9f76cc = hmaster0_p & v9f7692 | !hmaster0_p & v9f7d5b;
assign d3501c = hbusreq1_p & d357dc | !hbusreq1_p & d3501b;
assign bd574b = hbusreq2 & bd574a | !hbusreq2 & v845542;
assign ad45f2 = hbusreq0 & ad45ee | !hbusreq0 & ad45f1;
assign dc539d = hburst0_p & c74a04 | !hburst0_p & !dc539c;
assign v8cc790 = hgrant3_p & v8cc78d | !hgrant3_p & v8cc78f;
assign b5744b = decide_p & b57a2d | !decide_p & b57435;
assign bd5736 = hmaster2_p & bd572e | !hmaster2_p & bd5735;
assign v9f76e9 = hmaster2_p & v9f76e8 | !hmaster2_p & v9f7c9f;
assign d359ea = hbusreq1 & d359e9 | !hbusreq1 & v845542;
assign ad46f0 = hbusreq2 & ad46b4 | !hbusreq2 & !v845547;
assign ade4d7 = hmastlock_p & c3d673 | !hmastlock_p & !v845542;
assign ad4e5b = hbusreq0_p & v845542 | !hbusreq0_p & ad4e54;
assign df5166 = hbusreq1_p & df5165 | !hbusreq1_p & v845542;
assign bd5821 = hmaster2_p & bd581c | !hmaster2_p & bd5820;
assign b1c792 = hbusreq1 & b1c71c | !hbusreq1 & b1c71d;
assign ac1452 = hlock3_p & ac1451 | !hlock3_p & cc36ba;
assign df5128 = hmaster0_p & df5127 | !hmaster0_p & df54f4;
assign v9f78ad = hgrant3_p & v9f7875 | !hgrant3_p & v9f78ac;
assign b1c758 = hbusreq0 & b1c757 | !hbusreq0 & !v845542;
assign v8cc807 = hlock2 & v8cc43a | !hlock2 & v8cc806;
assign v9f7d51 = hmaster1_p & v9f7d3c | !hmaster1_p & v9f7d47;
assign ad41ac = decide_p & ad40f1 | !decide_p & ad41ab;
assign v9f78a7 = hgrant2_p & v9f78a4 | !hgrant2_p & v9f78a6;
assign v9ea5e8 = decide_p & v9ea5ca | !decide_p & v9ea5e7;
assign df507b = hmaster0_p & df507a | !hmaster0_p & v845542;
assign b05921 = hbusreq1_p & b0591f | !hbusreq1_p & b05920;
assign ad4e61 = hmaster0_p & ad4e59 | !hmaster0_p & ad4e60;
assign c3d6c6 = hbusreq4_p & c3d6c3 | !hbusreq4_p & !c3d6c5;
assign b57500 = hbusreq2 & b574fe | !hbusreq2 & b574ff;
assign v9e9f6f = hready & v9e9f6e | !hready & v9e9f68;
assign v9ea59d = hmaster2_p & v9ea4d2 | !hmaster2_p & v9ea59c;
assign v8cc507 = decide_p & v8cc506 | !decide_p & v8cc43f;
assign adea9a = locked_p & adea99 | !locked_p & !v845542;
assign v9f78a3 = hmaster0_p & v9f77b5 | !hmaster0_p & v9f7790;
assign ad47fd = hmaster0_p & ad456f | !hmaster0_p & ad470d;
assign c3ce88 = decide_p & c3ce7c | !decide_p & !c3ce71;
assign adeaad = hgrant3_p & adea90 | !hgrant3_p & adeaac;
assign ad40fe = hbusreq1 & v845547 | !hbusreq1 & v845542;
assign v9f7e06 = hgrant1_p & v9f7e05 | !hgrant1_p & v9f7dbb;
assign b1c6fb = hmaster1_p & b1c85a | !hmaster1_p & b1c6fa;
assign d35648 = hbusreq1_p & d35647 | !hbusreq1_p & !v845542;
assign dc502e = hbusreq1_p & dc5014 | !hbusreq1_p & dc502d;
assign ad46bf = hbusreq0 & ad46be | !hbusreq0 & ad469f;
assign bd5b9a = hlock2_p & bd5b99 | !hlock2_p & !v845542;
assign ac1463 = stateG10_4_p & v845542 | !stateG10_4_p & !adea92;
assign c5c8e4 = busreq_p & c5c8e2 | !busreq_p & !c5c8e3;
assign c3d581 = hgrant1_p & v84554d | !hgrant1_p & c3d580;
assign v9f784b = hlock3 & v9f784a | !hlock3 & v9f7849;
assign b1c6f9 = hgrant1_p & b1d01a | !hgrant1_p & b1c6f8;
assign d356d9 = hbusreq1_p & d356d8 | !hbusreq1_p & v845542;
assign bd586c = hgrant4_p & ade589 | !hgrant4_p & bd580d;
assign b1cf33 = hbusreq3 & b1cf32 | !hbusreq3 & b1cf2c;
assign d357b3 = hready_p & d3577f | !hready_p & d357b2;
assign ad4104 = hready & ad4103 | !hready & ad4ea6;
assign d357ff = hbusreq1_p & d357a5 | !hbusreq1_p & d357fe;
assign v8cc630 = hbusreq2_p & v8cc62f | !hbusreq2_p & v8ccbda;
assign v9ea447 = stateG10_4_p & v9ea445 | !stateG10_4_p & v9ea446;
assign ad4d98 = hready & ad4d96 | !hready & !ad4d97;
assign c3d5c5 = hbusreq2 & c3d5c4 | !hbusreq2 & c3d306;
assign dc5060 = stateG10_4_p & ade59c | !stateG10_4_p & !dc505f;
assign v8cc7d8 = hburst1_p & bbbcd8 | !hburst1_p & !bbbcd6;
assign v9f7772 = hbusreq2 & v9f7770 | !hbusreq2 & v9f7771;
assign v9f7e1d = stateG10_4_p & v9f7d89 | !stateG10_4_p & v9f7e1c;
assign ad41a4 = hmaster0_p & ad41a2 | !hmaster0_p & ad41a3;
assign b1c74b = hlock3_p & b1c730 | !hlock3_p & b1c74a;
assign d356c8 = hbusreq3 & d356c7 | !hbusreq3 & v84554e;
assign v9ea4c7 = hgrant4_p & v9ea4b6 | !hgrant4_p & v9ea4c6;
assign b1d004 = hbusreq3 & b1cffd | !hbusreq3 & b1d003;
assign ad4d9a = hburst0 & bd5b69 | !hburst0 & bd5b6b;
assign c3ce7d = decide_p & c3ce7c | !decide_p & !c3d36c;
assign d3573a = hbusreq2_p & d356ee | !hbusreq2_p & d35739;
assign v9f7dc2 = hlock3 & v9f7dc1 | !hlock3 & v9f7dbd;
assign d357a6 = hmaster0_p & d3579b | !hmaster0_p & d357a5;
assign d354e1 = hmaster1_p & d354e0 | !hmaster1_p & d354db;
assign d35026 = jx1_p & d35025 | !jx1_p & d3576a;
assign d356e3 = hlock1_p & v845542 | !hlock1_p & d3591c;
assign b57a2d = hbusreq2_p & b5795b | !hbusreq2_p & b57a2c;
assign v8cc4f3 = hmaster1_p & v8cc4f0 | !hmaster1_p & v8cc4f2;
assign b05a0c = hbusreq4_p & b05a0a | !hbusreq4_p & b05a0b;
assign v9f7dee = hbusreq1 & v9f7dec | !hbusreq1 & v9f7ded;
assign b1c79d = hlock0_p & b1c79c | !hlock0_p & !b1c70e;
assign c3cee1 = hmaster2_p & c3cedd | !hmaster2_p & v845542;
assign v8cc7b9 = hgrant4_p & v8cc796 | !hgrant4_p & v845542;
assign v9f7879 = hmaster1_p & v9f7878 | !hmaster1_p & v9f77f4;
assign b1c04e = hmaster0_p & b1c04d | !hmaster0_p & b1c78c;
assign ad456f = hbusreq4 & adec93 | !hbusreq4 & v845542;
assign cc36c3 = hready_p & cc36bc | !hready_p & cc36c2;
assign c3ce69 = hmaster0_p & c3ce67 | !hmaster0_p & c3ce68;
assign b0595f = hbusreq4 & b0595d | !hbusreq4 & b0595e;
assign v9f788e = hgrant1_p & v9f7730 | !hgrant1_p & v9f788d;
assign ad426c = hbusreq1 & ad426b | !hbusreq1 & v845542;
assign ad504f = hmaster2_p & ad503d | !hmaster2_p & ad504e;
assign c3d6d5 = hmaster0_p & c3d683 | !hmaster0_p & c3d682;
assign d35a28 = hlock2_p & d35a1d | !hlock2_p & !d35a27;
assign ade57d = hbusreq1_p & ade568 | !hbusreq1_p & ade57c;
assign c5c8e8 = hmaster2_p & c5c8e7 | !hmaster2_p & c5c88e;
assign b1c6bc = hmaster0_p & b1cfb8 | !hmaster0_p & b1c6bb;
assign d35a27 = hgrant2_p & d35a26 | !hgrant2_p & !d35a1c;
assign ad4785 = hbusreq2_p & ad4784 | !hbusreq2_p & ad4783;
assign d35589 = hbusreq1 & d354ff | !hbusreq1 & d35501;
assign v9f7680 = hlock3 & v9f767f | !hlock3 & v9f767e;
assign ad45b8 = hbusreq4_p & ad45b7 | !hbusreq4_p & !v845542;
assign ad4db5 = hbusreq0 & ad4db3 | !hbusreq0 & ad4db4;
assign c3d313 = hbusreq4 & c3d311 | !hbusreq4 & !c3d312;
assign b1c5fc = hbusreq2_p & b1c5dc | !hbusreq2_p & b1c84b;
assign d359df = hmaster2_p & d359a7 | !hmaster2_p & d359de;
assign v9ea4a1 = hgrant3_p & v9ea40b | !hgrant3_p & v9ea4a0;
assign ad3cea = hbusreq1 & ad3ccf | !hbusreq1 & ad3cd8;
assign c3ce2d = decide_p & c3ce2c | !decide_p & c3ce09;
assign v84557e = stateG3_0_p & v845542 | !stateG3_0_p & !v845542;
assign b578f4 = hlock3_p & b578f3 | !hlock3_p & v845542;
assign b57ac9 = hbusreq3 & b578f9 | !hbusreq3 & b57ac8;
assign b059be = hburst0_p & v845568 | !hburst0_p & d355a4;
assign bd575c = hmaster1_p & bd574c | !hmaster1_p & bd575b;
assign v8cc7c8 = hlock1 & v8ccbf4 | !hlock1 & v8cc7c5;
assign c3d508 = hgrant2_p & v845551 | !hgrant2_p & c3d507;
assign v9f770a = hmaster0_p & v9f7709 | !hmaster0_p & !v9f7df6;
assign v9f7767 = hbusreq2 & v9f7765 | !hbusreq2 & v9f7766;
assign d3577b = hbusreq0 & d3577a | !hbusreq0 & v845542;
assign adeaa4 = stateG10_4_p & v845542 | !stateG10_4_p & !v845576;
assign b57ad2 = hlock2_p & b57acc | !hlock2_p & b57ad1;
assign ad4462 = hlock4_p & ad4461 | !hlock4_p & !v845576;
assign bd587c = hburst0 & adea97 | !hburst0 & dc504e;
assign c3d52b = hbusreq1_p & c3d47c | !hbusreq1_p & c3d52a;
assign v9e9f75 = hgrant4_p & v9e9eec | !hgrant4_p & v9e9f74;
assign ade4c9 = stateA1_p & adea85 | !stateA1_p & !c74621;
assign ad48ca = hgrant3_p & ad5090 | !hgrant3_p & ad48c9;
assign v9ea4b5 = hmaster0_p & v9ea4b4 | !hmaster0_p & v9ea3fc;
assign v9f7759 = hmaster2_p & v9f7743 | !hmaster2_p & v9f772f;
assign v9f7760 = hbusreq1 & v9f775e | !hbusreq1 & v9f775f;
assign ad4dc8 = hlock1_p & ad4dc7 | !hlock1_p & ad4da1;
assign b1c75e = hbusreq2 & b1c758 | !hbusreq2 & b1c75c;
assign v9e9fd6 = decide_p & v9ea3f4 | !decide_p & v9e9fd5;
assign v9f789f = hmaster1_p & v9f77fe | !hmaster1_p & v9f7811;
assign ad4469 = hmaster0_p & ad443e | !hmaster0_p & ad4468;
assign ad431d = hmaster1_p & ad4315 | !hmaster1_p & ad431c;
assign ad46e2 = hready & ad46cd | !hready & ad46e1;
assign v9ea5f8 = hbusreq2_p & v9ea406 | !hbusreq2_p & v9ea5f7;
assign b1c729 = hbusreq0 & b1c728 | !hbusreq0 & v845542;
assign v9f777c = hbusreq2_p & v9f7775 | !hbusreq2_p & v9f777b;
assign ad3ce9 = hbusreq1_p & ad440e | !hbusreq1_p & ad3ce8;
assign ad45a9 = hbusreq2_p & ad45a6 | !hbusreq2_p & ad45a8;
assign ade4b3 = hmaster1_p & ade4b2 | !hmaster1_p & ade4af;
assign v8cc7ea = hbusreq3 & v8cc7e8 | !hbusreq3 & v8cc7e9;
assign df51ce = hbusreq3_p & df51a3 | !hbusreq3_p & df51cd;
assign ad4ef3 = locked_p & adea98 | !locked_p & !v845542;
assign v9f7dbe = hlock1_p & v9f7ca7 | !hlock1_p & v9f7cf8;
assign b1c738 = hmaster2_p & b1c731 | !hmaster2_p & c3d66d;
assign b1c5f3 = hbusreq2_p & b1c5f2 | !hbusreq2_p & b1c854;
assign c3ceb3 = hmaster0_p & c3ceb1 | !hmaster0_p & c3ceb2;
assign v9f7cb0 = hbusreq3 & v9f7cae | !hbusreq3 & v9f7caf;
assign ad40ee = hmaster1_p & v845551 | !hmaster1_p & ad40e7;
assign v9f7dbb = hbusreq1 & v9f7db9 | !hbusreq1 & v9f7dba;
assign v9f7863 = hlock1 & v9f785e | !hlock1 & v9f7862;
assign b1c80b = hbusreq3 & b1c808 | !hbusreq3 & !b1c80a;
assign v8cc5f9 = hlock2 & v8ccbd8 | !hlock2 & v8cc5f8;
assign ade585 = hbusreq1_p & ade57f | !hbusreq1_p & ade584;
assign v9ea622 = hbusreq3 & v9ea621 | !hbusreq3 & v9ea3fa;
assign v9f7656 = hgrant0_p & v9f7e2f | !hgrant0_p & !v9f7c9f;
assign v9f7744 = hmaster2_p & v9f7743 | !hmaster2_p & v84557a;
assign dc4fb2 = hmaster0_p & dc4fa5 | !hmaster0_p & dc4fb1;
assign ade654 = hbusreq1_p & adea8b | !hbusreq1_p & adeaaf;
assign v9f7820 = hbusreq0 & v9f781e | !hbusreq0 & v9f781f;
assign v8587b7 = hbusreq1_p & v845564 | !hbusreq1_p & !v845542;
assign dc506a = hbusreq3 & dc4fe0 | !hbusreq3 & v845542;
assign d35427 = hmaster2_p & d35419 | !hmaster2_p & d3541f;
assign adea9d = hbusreq4_p & adea9c | !hbusreq4_p & !v845542;
assign b059bb = hbusreq3 & b059b9 | !hbusreq3 & b059ba;
assign ad5015 = hmastlock_p & ad5014 | !hmastlock_p & v845542;
assign b1c829 = hmaster1_p & b1c828 | !hmaster1_p & b1c775;
assign ad45c2 = hbusreq2 & ad45b6 | !hbusreq2 & ad45c0;
assign c3d74b = hgrant2_p & c3d73c | !hgrant2_p & !c3d74a;
assign dc501d = hgrant4_p & adeca0 | !hgrant4_p & !adeca1;
assign c3cf1a = hready & c3cf19 | !hready & !v845542;
assign ad45b1 = hmaster2_p & v845542 | !hmaster2_p & !ad45b0;
assign c3ce64 = hbusreq1 & c3d379 | !hbusreq1 & v845542;
assign v9ea611 = hmaster0_p & v9ea3fc | !hmaster0_p & v9ea4b4;
assign c3d2e9 = locked_p & c3d2e8 | !locked_p & !v845542;
assign adec99 = hburst0 & adea97 | !hburst0 & adec98;
assign c3d373 = hgrant0_p & v845542 | !hgrant0_p & !c3d372;
assign c3d31f = hmaster2_p & adeaa5 | !hmaster2_p & c3d31e;
assign b57901 = hmaster0_p & b578fc | !hmaster0_p & b57900;
assign dc5040 = hbusreq4_p & dc503d | !hbusreq4_p & dc503f;
assign d35bef = hmaster0_p & d35bec | !hmaster0_p & d35bee;
assign b1c707 = decide_p & b1c82f | !decide_p & b1d013;
assign b574cb = hlock3 & b579e5 | !hlock3 & b574ca;
assign b0593f = hbusreq4_p & v9ea463 | !hbusreq4_p & v9f769c;
assign b1c5e8 = hgrant0_p & d355a8 | !hgrant0_p & v845542;
assign dc5076 = hmaster0_p & dc5073 | !hmaster0_p & dc5075;
assign v9ea4df = hmaster1_p & v9ea4de | !hmaster1_p & v9ea4bd;
assign v9f7d23 = hmaster2_p & v9f7d20 | !hmaster2_p & v9f7d22;
assign ad4f19 = hbusreq2 & ad4e65 | !hbusreq2 & !v845542;
assign v9f776a = hbusreq4_p & v9f7768 | !hbusreq4_p & !v9f7769;
assign b57443 = hgrant3_p & b57946 | !hgrant3_p & b57442;
assign b1c03c = hbusreq2 & b1c035 | !hbusreq2 & b1c03a;
assign ad4387 = hbusreq0_p & ad4f3e | !hbusreq0_p & v845542;
assign b573e2 = hbusreq1_p & b573e1 | !hbusreq1_p & b57942;
assign ad4257 = hbusreq2 & ad4ff5 | !hbusreq2 & v845542;
assign cc36bb = hlock3_p & v84556c | !hlock3_p & !cc36ba;
assign bd5881 = hgrant4_p & ade572 | !hgrant4_p & !bd574e;
assign ad46d3 = hmaster2_p & v845542 | !hmaster2_p & ad46d2;
assign c3cee4 = hready & c3cee2 | !hready & !c3cee3;
assign v9f77a6 = hbusreq1_p & v9f7797 | !hbusreq1_p & v9f77a5;
assign v9ea597 = hbusreq3 & v9ea593 | !hbusreq3 & v9ea596;
assign d35a43 = hlock0_p & d35a41 | !hlock0_p & !d35a42;
assign ad43ba = hmaster0_p & ad43b5 | !hmaster0_p & ad43b9;
assign v9f7671 = hlock3 & v9f7670 | !hlock3 & v9f766f;
assign c5c3be = hbusreq3_p & c5c3b7 | !hbusreq3_p & c5c9b5;
assign d35920 = hmaster1_p & d3590b | !hmaster1_p & d3591d;
assign b05a15 = hbusreq1_p & b05a0d | !hbusreq1_p & b05a14;
assign b1c71b = hmaster2_p & b1c70f | !hmaster2_p & b1c71a;
assign d35c01 = hmaster2_p & d35c00 | !hmaster2_p & !v84555a;
assign b5744d = hready_p & b5744b | !hready_p & b5744c;
assign df519b = hgrant1_p & v84556c | !hgrant1_p & !df519a;
assign ad414a = hgrant1_p & v845542 | !hgrant1_p & ad4e8e;
assign ad427d = hbusreq3 & ad427c | !hbusreq3 & v845542;
assign b1c76a = hbusreq0 & b1c769 | !hbusreq0 & !v845542;
assign ac148b = hbusreq1_p & ac145c | !hbusreq1_p & ac148a;
assign ad4fe8 = stateG10_4_p & ad4fe6 | !stateG10_4_p & ad4fe7;
assign aa4260 = jx2_p & aa425d | !jx2_p & !aa425f;
assign d356fb = hbusreq2 & d356b6 | !hbusreq2 & d356ad;
assign b579e4 = hgrant1_p & v845542 | !hgrant1_p & b579e3;
assign ade563 = hlock0_p & v84556c | !hlock0_p & !ade562;
assign c3d2de = hbusreq1 & v845564 | !hbusreq1 & v845542;
assign bd56d3 = hburst0 & dc5318 | !hburst0 & bd56d2;
assign ad4722 = hmaster1_p & ad4721 | !hmaster1_p & ad471b;
assign ad3cbf = hmaster1_p & ad3cbe | !hmaster1_p & ad43ba;
assign v9f787e = hlock2_p & v9f787a | !hlock2_p & v9f787d;
assign c3ce93 = hmaster0_p & c3ce13 | !hmaster0_p & c3ce92;
assign ad3cfd = hbusreq1_p & ad3cea | !hbusreq1_p & ad3cfc;
assign ad459b = hmaster2_p & adec93 | !hmaster2_p & v845542;
assign v9ea61b = hmaster1_p & v9ea61a | !hmaster1_p & v9ea3f0;
assign b05a04 = hmaster1_p & b05a03 | !hmaster1_p & b05943;
assign v9f765a = stateG10_4_p & v9f7658 | !stateG10_4_p & v9f7659;
assign d35524 = hbusreq1_p & d35514 | !hbusreq1_p & d35522;
assign b1c049 = hmaster1_p & b1c03d | !hmaster1_p & b1c048;
assign b058fa = hbusreq4 & b058f8 | !hbusreq4 & b058f9;
assign b058b4 = hlock2 & b058aa | !hlock2 & b058b3;
assign d3557a = hbusreq4_p & d354c0 | !hbusreq4_p & !d35aab;
assign ad4608 = hmaster2_p & adec93 | !hmaster2_p & ad4607;
assign c3cf01 = hmaster2_p & c3cf00 | !hmaster2_p & !v845542;
assign b1c07a = hgrant1_p & b1c078 | !hgrant1_p & b1c079;
assign ad4352 = hmaster0_p & ad4320 | !hmaster0_p & ad4293;
assign ad4301 = hmaster1_p & ad42fe | !hmaster1_p & ad4300;
assign c3ceb8 = hbusreq2_p & c3ce91 | !hbusreq2_p & c3ceb7;
assign c3d2ee = hmaster2_p & c3d2ed | !hmaster2_p & v845542;
assign v9e9fb4 = hready_p & v9ea436 | !hready_p & v9e9fb3;
assign ad4ed6 = hbusreq4_p & ad4ed3 | !hbusreq4_p & ad4ed5;
assign c3d672 = hmaster0_p & c3d66f | !hmaster0_p & c3d671;
assign ad439c = hmaster1_p & ad4391 | !hmaster1_p & ad439b;
assign c3d35e = hbusreq3 & c3d35d | !hbusreq3 & c3d306;
assign v9f77b3 = hbusreq3 & v9f77a5 | !hbusreq3 & v9f77b2;
assign v9f7dd1 = hgrant4_p & v9f7cd8 | !hgrant4_p & v9f7dd0;
assign ba7c76 = jx1_p & ba7c75 | !jx1_p & ba7c72;
assign v845549 = hbusreq0 & v845542 | !hbusreq0 & !v845542;
assign d357d1 = hbusreq1_p & d357d0 | !hbusreq1_p & v84554a;
assign ac146f = hgrant2_p & cc36d3 | !hgrant2_p & ac146d;
assign ad3d04 = hbusreq0 & ad3d03 | !hbusreq0 & v845542;
assign ad4fe5 = hbusreq0_p & v845542 | !hbusreq0_p & !ad4fe4;
assign d35652 = hlock0_p & d35651 | !hlock0_p & ade562;
assign ad4761 = hmaster1_p & ad4760 | !hmaster1_p & ad45a5;
assign b1c7c2 = hbusreq0 & b1c7c1 | !hbusreq0 & b1cfcc;
assign b05a9e = jx2_p & b0589f | !jx2_p & !b05a9d;
assign ade4cd = hbusreq4_p & ade4cc | !hbusreq4_p & !v845542;
assign d3549d = hmaster0_p & d3549b | !hmaster0_p & d3549c;
assign b1c615 = jx0_p & b1c86b | !jx0_p & b1c614;
assign b058bd = hready & b058bc | !hready & b058b8;
assign ad42aa = hlock1_p & ad42a9 | !hlock1_p & !v84554d;
assign b573f7 = hbusreq2_p & b573e0 | !hbusreq2_p & b573f6;
assign stateG3_2 = !v9e9fe9;
assign d35a21 = hmaster2_p & v84557a | !hmaster2_p & !adeca0;
assign bd57df = hgrant1_p & bd57de | !hgrant1_p & dc4fb0;
assign ad47f0 = hmaster1_p & ad47ef | !hmaster1_p & ad46ec;
assign v845564 = hmaster2_p & v845542 | !hmaster2_p & !v845542;
assign ad3d43 = hmaster0_p & ad3cc0 | !hmaster0_p & ad4488;
assign ad5045 = hmaster2_p & ad503d | !hmaster2_p & ad5044;
assign v8da5a6 = hgrant2_p & v845542 | !hgrant2_p & v8da5a4;
assign b573fb = hbusreq3 & b573e3 | !hbusreq3 & b57942;
assign b1c7b0 = hbusreq1 & b1c713 | !hbusreq1 & b1c718;
assign b1c768 = hbusreq0 & b1c767 | !hbusreq0 & !v845542;
assign b059a6 = hlock2_p & b059a2 | !hlock2_p & b059a5;
assign d357e1 = hgrant2_p & v84554a | !hgrant2_p & d357df;
assign v9ea5f6 = hmaster0_p & v9ea3fa | !hmaster0_p & v9ea4b7;
assign v8cc4a8 = hbusreq4 & v8cc4a6 | !hbusreq4 & v8cc4a7;
assign b05a66 = hgrant4_p & b058a3 | !hgrant4_p & b05a65;
assign bd5b90 = hbusreq2_p & bd5b8f | !hbusreq2_p & !v845542;
assign b57450 = jx1_p & b57405 | !jx1_p & b5744f;
assign dc53be = decide_p & dc53bd | !decide_p & v845542;
assign bd5ba2 = hbusreq2 & dc53a3 | !hbusreq2 & v845564;
assign v9f76bd = decide_p & v9f76b7 | !decide_p & v9f76bc;
assign cc36f3 = hgrant4_p & v845542 | !hgrant4_p & !cc36f2;
assign ade5be = hbusreq3 & ade548 | !hbusreq3 & !v845558;
assign ad4f6c = hmaster2_p & ad4f66 | !hmaster2_p & ad4f6b;
assign d3551c = hmaster1_p & d3542e | !hmaster1_p & d3551a;
assign b578f1 = hmaster2_p & v845542 | !hmaster2_p & b5b408;
assign bd5e9d = hlock4_p & bd5b88 | !hlock4_p & !d35a4f;
assign b5743b = hmaster1_p & b579b4 | !hmaster1_p & b5743a;
assign v9f7837 = hgrant1_p & v9f778c | !hgrant1_p & v9f7836;
assign v9ea483 = hlock1 & v9ea46d | !hlock1 & v9ea482;
assign v9f781a = hgrant0_p & v9f7785 | !hgrant0_p & v9f7743;
assign v9e9f85 = hlock3 & v9e9f84 | !hlock3 & v9e9f81;
assign c3d52d = hbusreq2 & c3d527 | !hbusreq2 & c3d52b;
assign b1c61c = hready_p & v845542 | !hready_p & b1c61b;
assign v8cc79c = hready & v8cc79b | !hready & v8ccb6b;
assign c3cef2 = hmaster2_p & c3cef1 | !hmaster2_p & v845542;
assign ad4315 = hgrant1_p & v845542 | !hgrant1_p & ad4314;
assign ad42b9 = hready & v9c81a4 | !hready & ad42b8;
assign v8cc130 = hgrant3_p & v8cc12b | !hgrant3_p & v8cc12f;
assign v9e9fb9 = hmaster0_p & v9e9fb8 | !hmaster0_p & v9e9ee9;
assign dc4f7d = hbusreq4_p & dc4f7c | !hbusreq4_p & !ade4d9;
assign b1c77a = hlock2_p & b1c776 | !hlock2_p & b1c779;
assign ac1470 = hlock2_p & ac146e | !hlock2_p & ac146f;
assign v9f785d = hbusreq4_p & v9f772a | !hbusreq4_p & v9f785c;
assign d359c0 = hburst0 & d359bb | !hburst0 & d359bf;
assign bd5b6a = hmastlock_p & bd5b69 | !hmastlock_p & v845542;
assign b05911 = hlock2 & b058d5 | !hlock2 & b05910;
assign v9f7881 = hbusreq0_p & v9f77be | !hbusreq0_p & v9f7880;
assign d35907 = hmastlock_p & d35906 | !hmastlock_p & !v845542;
assign b1c7ad = hbusreq0 & b1c7ac | !hbusreq0 & b1cfcc;
assign bb9bdd = hburst0_p & v845542 | !hburst0_p & bb9bdc;
assign bd5901 = decide_p & bd58f3 | !decide_p & !v845572;
assign v9f77af = hmaster2_p & v9f77ac | !hmaster2_p & v9f77ae;
assign v9f77e7 = hlock4_p & d35a0b | !hlock4_p & !v845542;
assign c3ce30 = hgrant3_p & c3ce28 | !hgrant3_p & c3ce2f;
assign ad4e6d = hgrant0_p & d3597f | !hgrant0_p & !ad4e6c;
assign v9f7888 = hbusreq0 & v9f7886 | !hbusreq0 & v9f7887;
assign b574cd = hlock2 & b579e5 | !hlock2 & b574cc;
assign v9f7d79 = hlock0_p & v9f7d78 | !hlock0_p & !v9f7c9f;
assign b1c7fe = hgrant3_p & b1c78a | !hgrant3_p & b1c7fd;
assign ad3cd9 = hgrant1_p & ad4411 | !hgrant1_p & ad3cd8;
assign ad503a = hgrant4_p & ad5016 | !hgrant4_p & cc36fc;
assign dc4f70 = hmaster2_p & ade4bf | !hmaster2_p & !ade4d9;
assign c3d5e3 = hbusreq0 & c3d5e0 | !hbusreq0 & c3d5e2;
assign b1c5f0 = hmaster1_p & b1cfb8 | !hmaster1_p & b1c5ef;
assign d35ab2 = hmaster2_p & d35ab1 | !hmaster2_p & d35aac;
assign bd5e1f = hbusreq2 & dc5317 | !hbusreq2 & bd5e1e;
assign b05a89 = hmaster1_p & b05a88 | !hmaster1_p & b058e1;
assign d354a8 = hlock4_p & v845542 | !hlock4_p & !d35a45;
assign bd57ff = hgrant4_p & bd572e | !hgrant4_p & bd57fe;
assign v8cc803 = hgrant1_p & v845542 | !hgrant1_p & v8cc802;
assign bd578b = hburst0 & d35617 | !hburst0 & bd578a;
assign ad43f9 = hbusreq0 & ad43f8 | !hbusreq0 & !v845542;
assign ad4413 = hready & b1c71d | !hready & !v845542;
assign b1c852 = hmaster0_p & b1cfb8 | !hmaster0_p & b1c851;
assign dc4fd0 = hmaster2_p & v84556c | !hmaster2_p & adec9a;
assign b1c037 = hbusreq4_p & ade4d9 | !hbusreq4_p & b1c036;
assign ad46da = hgrant0_p & ad4566 | !hgrant0_p & v845542;
assign v9f7d77 = hbusreq4_p & v9f7d75 | !hbusreq4_p & v9f7d76;
assign v9ea406 = hmaster1_p & v9ea3fd | !hmaster1_p & v9ea405;
assign b1c088 = hbusreq1_p & b1c7e1 | !hbusreq1_p & b1c087;
assign v9e9f63 = hbusreq2 & v9e9f61 | !hbusreq2 & v9e9f62;
assign bd5b7d = decide_p & bd5b7c | !decide_p & v845542;
assign b058a4 = stateG2_p & v845542 | !stateG2_p & !v857440;
assign dc504d = hmastlock_p & dc504c | !hmastlock_p & v845542;
assign v9f7cba = hlock4 & v9f7cb7 | !hlock4 & v9f7cb9;
assign d35a98 = hbusreq4_p & v845542 | !hbusreq4_p & v845548;
assign b05960 = hready & b0595f | !hready & b0595b;
assign c3d377 = hbusreq3 & c3d376 | !hbusreq3 & v845542;
assign v9e9f8f = hgrant4_p & v9e9f6a | !hgrant4_p & v9e9f74;
assign ad4359 = hmaster1_p & ad4358 | !hmaster1_p & ad42d9;
assign ad432c = hmaster1_p & ad432b | !hmaster1_p & ad42d9;
assign cc36c6 = hbusreq1_p & cc36c5 | !hbusreq1_p & !cc36b8;
assign ad4f08 = hbusreq4_p & ad4f07 | !hbusreq4_p & b1cfbe;
assign ad4f8c = hbusreq4_p & ad4f89 | !hbusreq4_p & ad4f8b;
assign d35415 = hbusreq2_p & d35411 | !hbusreq2_p & d35414;
assign b0597c = stateG10_4_p & v9f7d42 | !stateG10_4_p & b0597b;
assign d354af = locked_p & d354ae | !locked_p & v845542;
assign b059ac = hgrant2_p & b059a8 | !hgrant2_p & b059ab;
assign dc4fad = hmaster2_p & dc4fac | !hmaster2_p & dc4fa7;
assign d3542a = hmaster0_p & d35426 | !hmaster0_p & d35429;
assign ad42cb = hmaster0_p & ad42c8 | !hmaster0_p & ad42c3;
assign v8cc788 = hbusreq2 & v8cc786 | !hbusreq2 & v8cc787;
assign b1c5db = hmaster1_p & v845542 | !hmaster1_p & b1c5da;
assign bd583a = hbusreq1 & bd5839 | !hbusreq1 & !dc501a;
assign ad4277 = hlock1_p & ad4eca | !hlock1_p & ad4f62;
assign d359e3 = hgrant1_p & d359cc | !hgrant1_p & d359e2;
assign v9ea4af = hmaster0_p & v9ea4a9 | !hmaster0_p & v9ea4ae;
assign v9ea579 = hmaster0_p & v9ea576 | !hmaster0_p & v9ea578;
assign v9e9ea1 = hgrant1_p & v9ea3fc | !hgrant1_p & v9e9ea0;
assign ade59f = hlock4_p & ade59d | !hlock4_p & !ade59e;
assign d35997 = hlock0_p & d35995 | !hlock0_p & !d35996;
assign df518a = hbusreq2 & df5189 | !hbusreq2 & !v84554c;
assign v9ea613 = hmaster0_p & v9ea44a | !hmaster0_p & v9ea4cb;
assign v9f7705 = hgrant1_p & v9f7dbf | !hgrant1_p & v9f7704;
assign b0591d = hmaster2_p & b0591c | !hmaster2_p & b058a6;
assign v9e9f99 = hgrant1_p & v9e9ef0 | !hgrant1_p & v9e9f98;
assign b1c497 = hmaster2_p & v845542 | !hmaster2_p & b1c496;
assign b1c7bb = hgrant0_p & v84556c | !hgrant0_p & !bd574e;
assign v9f7d21 = hbusreq0_p & v9ea3ec | !hbusreq0_p & !v9f7cc6;
assign b1cfd2 = hbusreq3 & b1cfc9 | !hbusreq3 & b1cfd1;
assign ac1459 = hgrant4_p & v845542 | !hgrant4_p & ac1458;
assign b8f6e3 = hmaster0_p & b8f6e1 | !hmaster0_p & b8f6e2;
assign ad46fa = hbusreq2_p & ad46ef | !hbusreq2_p & !ad46f9;
assign b05957 = hlock4_p & b05955 | !hlock4_p & b05956;
assign v8ccb87 = hlock2_p & v8ccb82 | !hlock2_p & v8ccb84;
assign v9ea5e4 = hmaster1_p & v9ea5e3 | !hmaster1_p & v9ea583;
assign bd585b = hgrant4_p & bd5735 | !hgrant4_p & adec89;
assign d354cc = hbusreq4_p & d354cb | !hbusreq4_p & v845542;
assign df5150 = hbusreq1_p & df514f | !hbusreq1_p & v845542;
assign bd5849 = hgrant4_p & v84556c | !hgrant4_p & bd574e;
assign v9e9eba = hgrant1_p & v9ea4b7 | !hgrant1_p & v9e9eb9;
assign ade616 = hmaster0_p & ade615 | !hmaster0_p & ade541;
assign b579b8 = stateA1_p & b579b7 | !stateA1_p & b578f7;
assign b573e4 = hbusreq3 & b573e2 | !hbusreq3 & b573e3;
assign dc5028 = hgrant4_p & v845542 | !hgrant4_p & !adeca1;
assign b059d1 = hbusreq3 & b059cd | !hbusreq3 & b059d0;
assign ad46cd = hbusreq4 & ad46cc | !hbusreq4 & v845542;
assign b0ed8b = stateG2_p & v845542 | !stateG2_p & c74202;
assign v9f7cfc = hbusreq4 & v9f7cfa | !hbusreq4 & v9f7cfb;
assign v9f7e35 = hlock4 & v9f7e32 | !hlock4 & v9f7e34;
assign b05a77 = hlock2 & b05a74 | !hlock2 & b05a76;
assign d3562d = hbusreq2_p & d3562c | !hbusreq2_p & d35a97;
assign b579bd = hbusreq0 & b579bb | !hbusreq0 & b579bc;
assign d354ca = hbusreq1_p & d354c9 | !hbusreq1_p & d354c8;
assign v9ea3e1 = hmaster2_p & v845542 | !hmaster2_p & v9f21c5;
assign b05a6f = hlock1 & b05a69 | !hlock1 & b05a6e;
assign v8cc0df = hlock1 & v8cc494 | !hlock1 & v8cc0de;
assign c3d6cd = hgrant4_p & c3d689 | !hgrant4_p & c3d6cb;
assign c3d2ba = hbusreq1 & c3d2b2 | !hbusreq1 & c3d2b6;
assign v9e9eec = hlock0_p & v9e9eeb | !hlock0_p & v9ea4b6;
assign b1c08b = hmaster1_p & b1c076 | !hmaster1_p & b1c08a;
assign b1c799 = hgrant4_p & b1c731 | !hgrant4_p & !b1c797;
assign ad43bd = hmaster1_p & ad43bc | !hmaster1_p & ad43ba;
assign ad4775 = hbusreq4_p & ad4774 | !hbusreq4_p & !v845542;
assign v9e9ef7 = hready_p & v9ea3e3 | !hready_p & v9e9ef6;
assign bd58be = hgrant4_p & v84556c | !hgrant4_p & bd58bd;
assign df5187 = hgrant2_p & df5179 | !hgrant2_p & !df5186;
assign v9f7722 = hready_p & v9f7716 | !hready_p & !v9f7721;
assign v8cc822 = hlock3 & v8cc501 | !hlock3 & v8cc821;
assign ad42c9 = hmaster0_p & ad42c8 | !hmaster0_p & ad42a7;
assign dc53d8 = decide_p & dc53d7 | !decide_p & !v845542;
assign ad4e8c = hgrant4_p & v845542 | !hgrant4_p & b1cfcb;
assign v9f774d = hbusreq3 & v9f774b | !hbusreq3 & v9f774c;
assign c3d6f6 = hlock0_p & c3d6c7 | !hlock0_p & c3d6f5;
assign ad4153 = hbusreq4_p & ad4152 | !hbusreq4_p & ad4f38;
assign v9e9fa8 = hmaster1_p & v9e9fa7 | !hmaster1_p & v9e9ef1;
assign v9f7830 = hlock0 & v9f782f | !hlock0 & v9f782e;
assign v9f779e = hmaster2_p & v9f7785 | !hmaster2_p & !v9f779d;
assign dc500f = hgrant4_p & v845542 | !hgrant4_p & !ade563;
assign bd57b2 = hmaster1_p & bd5798 | !hmaster1_p & bd57b1;
assign v9f7d16 = hbusreq4 & v9f7d14 | !hbusreq4 & v9f7d15;
assign b57536 = jx1_p & b57509 | !jx1_p & b57535;
assign c3d67b = hmaster2_p & c3d678 | !hmaster2_p & c3d67a;
assign c3d4fb = hmaster2_p & v845542 | !hmaster2_p & c3d4fa;
assign d35a04 = hgrant4_p & d3598a | !hgrant4_p & d35a03;
assign b05948 = decide_p & b05935 | !decide_p & !b05947;
assign b058da = hready & b058d9 | !hready & b058d5;
assign ad47f2 = hlock2_p & ad47ed | !hlock2_p & !ad47f1;
assign b57aed = hready_p & b5799c | !hready_p & b57aec;
assign v9e9fcc = hgrant3_p & v9e9fbf | !hgrant3_p & v9e9fcb;
assign b57941 = locked_p & b578f9 | !locked_p & v845542;
assign v9f77f7 = hgrant2_p & v9f773b | !hgrant2_p & v9f77f5;
assign d35586 = hbusreq1_p & d354bb | !hbusreq1_p & !d35585;
assign v9f7d07 = hbusreq0 & v9f7d04 | !hbusreq0 & v9f7d06;
assign ad4eef = hgrant4_p & v845542 | !hgrant4_p & ad4ee3;
assign c3d526 = hready & c3d525 | !hready & v845542;
assign v8cc7f8 = hlock0_p & v8cc7bc | !hlock0_p & v8cc7f7;
assign v9f782a = hgrant0_p & v9f779d | !hgrant0_p & !v9f772f;
assign c3ce4f = hmaster1_p & c3ce45 | !hmaster1_p & c3ce4e;
assign v9f76a7 = hmaster1_p & v9f7691 | !hmaster1_p & v9f76a6;
assign ad4789 = hready_p & ad4763 | !hready_p & !ad4788;
assign v9f7de4 = hlock4_p & v9f7de2 | !hlock4_p & v9f7de3;
assign dc5045 = hbusreq4_p & dc5042 | !hbusreq4_p & dc5044;
assign ad5070 = hready_p & ad4ffb | !hready_p & ad506f;
assign d357f3 = hlock0_p & v845542 | !hlock0_p & !d357f2;
assign ba7c81 = jx2_p & ba7c77 | !jx2_p & ba7c80;
assign c3d72a = hbusreq2_p & c3d728 | !hbusreq2_p & c3d729;
assign v8cc0ee = hlock3 & v8ccbd8 | !hlock3 & v8cc0ec;
assign ad4484 = hbusreq0 & ad4483 | !hbusreq0 & v845542;
assign b05992 = hmaster2_p & b0598a | !hmaster2_p & !b05991;
assign bd58b6 = hbusreq1 & bd575e | !hbusreq1 & df513c;
assign ad4df1 = hbusreq3 & ad4df0 | !hbusreq3 & v845542;
assign b1c7d3 = stateG10_4_p & b1c7bc | !stateG10_4_p & b1c7d2;
assign ad4477 = hmaster0_p & ad43ab | !hmaster0_p & ad43a9;
assign v9e9ecc = hmaster0_p & v9e9e79 | !hmaster0_p & v9ea3fa;
assign d354a1 = hlock1_p & d3549f | !hlock1_p & !d354a0;
assign dc500a = hgrant4_p & v845542 | !hgrant4_p & !adec89;
assign ad437e = hmaster2_p & v845542 | !hmaster2_p & ad437d;
assign v9ea578 = hmaster2_p & v9ea4b9 | !hmaster2_p & v9ea577;
assign v9f77d2 = hbusreq3 & v9f77cf | !hbusreq3 & v9f77d1;
assign c3ce45 = hgrant1_p & v84554d | !hgrant1_p & c3ce44;
assign bd5762 = hmaster0_p & bd5760 | !hmaster0_p & bd5761;
assign ad4580 = hmaster1_p & ad4572 | !hmaster1_p & ad457f;
assign v9f7804 = hgrant1_p & v9f772c | !hgrant1_p & v9f77e1;
assign ad5068 = hgrant2_p & ad501f | !hgrant2_p & ad5067;
assign ad42c0 = hbusreq1 & ad4da1 | !hbusreq1 & v845542;
assign d35aa3 = hready_p & d35a94 | !hready_p & !d35aa2;
assign v8cc49f = stateG10_4_p & v845542 | !stateG10_4_p & v8cc49e;
assign v9e9ec2 = hbusreq3 & v9e9eb2 | !hbusreq3 & v9ea4cd;
assign d35768 = hready_p & d35767 | !hready_p & d35aa2;
assign ad4f62 = hbusreq1 & ad4f4c | !hbusreq1 & v845542;
assign v9f7cdd = hmaster2_p & v9f7cda | !hmaster2_p & v9f7cdc;
assign ade5cb = stateA1_p & ade5ca | !stateA1_p & !c74621;
assign b1cbf3 = hlock4_p & b1cfc6 | !hlock4_p & b1cffa;
assign ad4327 = hmaster1_p & ad4326 | !hmaster1_p & ad431c;
assign b05a49 = hmaster1_p & b05a48 | !hmaster1_p & b05943;
assign ad42bc = hbusreq1_p & ad42bb | !hbusreq1_p & v845542;
assign v9f76e7 = stateG10_4_p & v9f76e5 | !stateG10_4_p & v9f76e6;
assign ad474a = hmaster2_p & v845542 | !hmaster2_p & ad4749;
assign ad3cf9 = hmaster2_p & ad3ccc | !hmaster2_p & ad3cf8;
assign b1c7da = hgrant4_p & b1c734 | !hgrant4_p & b1c79d;
assign adec9e = hbusreq3 & adec8a | !hbusreq3 & adec93;
assign b1c733 = hbusreq0 & b1c732 | !hbusreq0 & v845542;
assign ad4135 = hgrant4_p & dc52fa | !hgrant4_p & v845542;
assign v9e9ea8 = hgrant1_p & v9ea4bc | !hgrant1_p & v9e9ea7;
assign b058c4 = hlock2 & b058b8 | !hlock2 & b058c3;
assign c3d3a4 = hbusreq1_p & c3d305 | !hbusreq1_p & c3d3a3;
assign c3cec2 = hbusreq0_p & v84556e | !hbusreq0_p & v845542;
assign ad4709 = hbusreq4 & ad4708 | !hbusreq4 & v845542;
assign v9f7e23 = hbusreq4 & v9f7e21 | !hbusreq4 & v9f7e22;
assign d35595 = hbusreq2_p & d3556f | !hbusreq2_p & !d35594;
assign dc4ffe = hbusreq1_p & dc4ffc | !hbusreq1_p & dc4ffd;
assign d35518 = hmaster2_p & v84555a | !hmaster2_p & d35517;
assign b058f1 = hbusreq1 & b058ef | !hbusreq1 & b058f0;
assign bd591a = hmaster1_p & bd5919 | !hmaster1_p & v84556c;
assign b1c564 = hbusreq4_p & b1d000 | !hbusreq4_p & !b1c85d;
assign d35a62 = hmaster2_p & d35a5b | !hmaster2_p & d35a61;
assign d35015 = hgrant1_p & d35805 | !hgrant1_p & d35014;
assign ad4eaf = hmaster2_p & v84557a | !hmaster2_p & !ad4eae;
assign c3cf25 = hmaster1_p & c3cf24 | !hmaster1_p & c3d36b;
assign c3d501 = hmaster2_p & adeaa5 | !hmaster2_p & c3d4f4;
assign b1c842 = hbusreq1_p & v845542 | !hbusreq1_p & b1c841;
assign c3d732 = hmaster0_p & c3d676 | !hmaster0_p & c3d66f;
assign ad3cc4 = hbusreq2_p & ad3cbd | !hbusreq2_p & ad3cc3;
assign ad4714 = hbusreq4 & ad4713 | !hbusreq4 & v845542;
assign b05975 = hbusreq2 & b05973 | !hbusreq2 & b05974;
assign b1c06c = hgrant4_p & v845542 | !hgrant4_p & b1c062;
assign c3ce89 = hready_p & c3ce87 | !hready_p & c3ce88;
assign v8cc7ff = hbusreq4 & v8cc7fd | !hbusreq4 & v8cc7fe;
assign ad47e8 = hbusreq2 & ad4576 | !hbusreq2 & v845542;
assign v9ea490 = hlock4 & v9ea43b | !hlock4 & v9ea48f;
assign b059ef = hgrant1_p & b058dc | !hgrant1_p & !b059ee;
assign bd577a = hmaster1_p & bd5774 | !hmaster1_p & bd5779;
assign b05924 = hlock0_p & b058a6 | !hlock0_p & !b058d3;
assign d358f4 = hbusreq3 & d358f3 | !hbusreq3 & v845542;
assign d35500 = hbusreq1_p & d35c0b | !hbusreq1_p & !d354ff;
assign ad5056 = hmaster2_p & ad5054 | !hmaster2_p & ad504e;
assign d35aac = hbusreq4_p & v845542 | !hbusreq4_p & !d35aab;
assign b574bb = hgrant1_p & b574ba | !hgrant1_p & b579b3;
assign d35509 = hbusreq4_p & d35508 | !hbusreq4_p & v845542;
assign ad435c = hbusreq2 & ad427c | !hbusreq2 & v845542;
assign d35a66 = hgrant4_p & v845542 | !hgrant4_p & d35a64;
assign dc502f = hgrant1_p & dc501c | !hgrant1_p & dc502e;
assign v845574 = hgrant3_p & v845542 | !hgrant3_p & !v845542;
assign ad4ebe = hbusreq0 & ad4eb8 | !hbusreq0 & ad4ebd;
assign ad3d4b = decide_p & ad3d40 | !decide_p & ad3d4a;
assign d355a7 = hburst0 & d355a6 | !hburst0 & d35a4d;
assign d356e2 = hbusreq1_p & d356e1 | !hbusreq1_p & v845542;
assign c3d741 = hgrant4_p & c3d669 | !hgrant4_p & !c3d740;
assign bd582b = hbusreq0 & bd5829 | !hbusreq0 & bd582a;
assign df5149 = hbusreq3 & df5146 | !hbusreq3 & df5148;
assign v8ccb67 = hburst0_p & bb9c5a | !hburst0_p & !v8ccb66;
assign v8cc7f0 = stateG10_4_p & v845542 | !stateG10_4_p & v8cc7ef;
assign v9ea425 = hmaster0_p & v9ea417 | !hmaster0_p & v9ea424;
assign c3d59a = hmaster1_p & c3d596 | !hmaster1_p & c3d599;
assign v8ccb6a = locked_p & v8ccb69 | !locked_p & v845542;
assign v9ea57f = hready_p & v9ea3e3 | !hready_p & v9ea57e;
assign b05a30 = hmaster1_p & b05a2f | !hmaster1_p & b05913;
assign c3d52a = hready & c3d529 | !hready & c3d47b;
assign d358ec = stateA1_p & c5c894 | !stateA1_p & v845542;
assign dc5055 = hgrant4_p & v84556c | !hgrant4_p & ade58d;
assign c3d74d = hmaster0_p & c3d701 | !hmaster0_p & c3d6e8;
assign ad43a6 = hbusreq0 & ad43a5 | !hbusreq0 & v845542;
assign b57ae9 = hmaster1_p & b579b4 | !hmaster1_p & b57ae8;
assign b05a42 = hbusreq1_p & b0591f | !hbusreq1_p & b05a40;
assign v8cc11f = hbusreq2_p & v8cc0eb | !hbusreq2_p & v8cc11e;
assign v9f7687 = hbusreq2_p & v9f7677 | !hbusreq2_p & v9f7686;
assign c3d6e3 = hbusreq4_p & c3d6e1 | !hbusreq4_p & c3d6e2;
assign b1c804 = hbusreq0 & b1c7b7 | !hbusreq0 & !d35a9c;
assign v9f7741 = busreq_p & v845542 | !busreq_p & v84557c;
assign v8cc7bc = hgrant0_p & v8cc796 | !hgrant0_p & v845542;
assign ad425f = hready_p & ad425c | !hready_p & ad425e;
assign c3d531 = hmaster0_p & c3d530 | !hmaster0_p & c3d2be;
assign b1c5b4 = hmaster0_p & v845542 | !hmaster0_p & b1c5b3;
assign d3599d = hmaster2_p & d3599c | !hmaster2_p & v845542;
assign v9f767d = hmaster1_p & v9f767c | !hmaster1_p & v9f7ce9;
assign d3541e = hlock4_p & v845542 | !hlock4_p & !dc5318;
assign b57a1e = hbusreq1_p & b578fb | !hbusreq1_p & b57a1c;
assign ad43b7 = hmaster2_p & ad43b6 | !hmaster2_p & v845542;
assign ad4de3 = hready & ad4de1 | !hready & !ad4de2;
assign v9f7d38 = hlock3_p & v9f7cf1 | !hlock3_p & v9f7d37;
assign d35983 = locked_p & v845542 | !locked_p & adeca0;
assign df5138 = hbusreq1 & df5137 | !hbusreq1 & v845542;
assign v9f7cae = hbusreq1 & v9f7cac | !hbusreq1 & v9f7cad;
assign b1cfb6 = hlock0_p & cc36fc | !hlock0_p & !v845542;
assign b1c580 = hbusreq0 & b1c4c9 | !hbusreq0 & b1c57f;
assign v9f7d1e = hlock2 & v9f7d1b | !hlock2 & v9f7d1d;
assign b1cf35 = hmaster1_p & v845542 | !hmaster1_p & b1cf34;
assign d35516 = hlock4_p & v845542 | !hlock4_p & !d35956;
assign ad46d4 = hbusreq0 & ad46d0 | !hbusreq0 & ad46d3;
assign c3d5f0 = hmaster2_p & c3d5e1 | !hmaster2_p & v845542;
assign b059dc = stateG10_4_p & b059da | !stateG10_4_p & !b059db;
assign b579c5 = hgrant1_p & b57942 | !hgrant1_p & b579b3;
assign dc53c7 = decide_p & dc53c4 | !decide_p & v845542;
assign b1c587 = hready_p & b1c56e | !hready_p & b1c586;
assign v9ea4bf = hmaster0_p & v9ea4b4 | !hmaster0_p & v9ea4b7;
assign dc5063 = hbusreq0 & dc5059 | !hbusreq0 & dc5062;
assign c3d37f = hgrant1_p & c3d2de | !hgrant1_p & c3d37e;
assign dc4f90 = hbusreq0 & dc4f7e | !hbusreq0 & dc4f8f;
assign ad4ff5 = hgrant1_p & v84556c | !hgrant1_p & ad4fc1;
assign d3590f = hbusreq3 & d3590e | !hbusreq3 & v845542;
assign c3d2cc = hbusreq3 & c3d2cb | !hbusreq3 & !v845542;
assign d35623 = hbusreq1 & d3560e | !hbusreq1 & d35618;
assign df51a1 = decide_p & df516c | !decide_p & d6ebca;
assign dc5032 = hbusreq4_p & c3d66d | !hbusreq4_p & !adeca0;
assign ad460e = hmaster0_p & ad460b | !hmaster0_p & ad460d;
assign c3d749 = hmaster0_p & c3d748 | !hmaster0_p & c3d6d1;
assign ad4fea = hmaster2_p & ad4fe3 | !hmaster2_p & ad4fe9;
assign v8cc4b9 = hbusreq2 & v8cc4b8 | !hbusreq2 & v8ccbd8;
assign v9f76c7 = hbusreq1_p & v9f7d3e | !hbusreq1_p & v9f76c6;
assign ad4ea4 = hmaster2_p & ad4e8a | !hmaster2_p & ad4ea3;
assign v9f7841 = hgrant4_p & v9f77ae | !hgrant4_p & !v9f780b;
assign df50d9 = hlock1_p & df50d8 | !hlock1_p & v845542;
assign df5178 = hmaster0_p & df5176 | !hmaster0_p & df5177;
assign v9e9ec9 = hbusreq2_p & v9e9ec6 | !hbusreq2_p & v9e9ec8;
assign v8cc7e3 = hbusreq4 & v8cc7e1 | !hbusreq4 & v8cc7e2;
assign b5744a = hready_p & b57446 | !hready_p & b57449;
assign v9f7daa = hbusreq1 & v9f7da8 | !hbusreq1 & v9f7da9;
assign ad4348 = hbusreq2_p & ad4342 | !hbusreq2_p & ad4347;
assign ad502b = hbusreq3 & ad502a | !hbusreq3 & ad5024;
assign b579d2 = hgrant4_p & v845542 | !hgrant4_p & b579d1;
assign ba7c6c = hgrant1_p & v845558 | !hgrant1_p & ba7c66;
assign v9ea3f9 = hlock3_p & v9ea3f4 | !hlock3_p & v9ea3f8;
assign ad4312 = hmaster1_p & ad4311 | !hmaster1_p & ad4297;
assign c5c891 = hmaster1_p & c5c890 | !hmaster1_p & v845542;
assign ad4740 = hgrant1_p & ad473e | !hgrant1_p & ad473f;
assign c3d326 = stateG10_4_p & v84556e | !stateG10_4_p & c3d2fd;
assign ade56d = locked_p & ade56c | !locked_p & adeca0;
assign v9f7dfe = hlock3 & v9f7da3 | !hlock3 & v9f7daa;
assign dc4f78 = hmastlock_p & adea86 | !hmastlock_p & !v845542;
assign c3ce82 = hgrant1_p & v84554d | !hgrant1_p & c3ce81;
assign c5c953 = decide_p & c5c92c | !decide_p & c5c952;
assign v9f7c9e = stateA1_p & v845542 | !stateA1_p & !v9f7c95;
assign ad4399 = hready & v845542 | !hready & ad4398;
assign bd5941 = jx0_p & bd5922 | !jx0_p & bd5940;
assign df54df = hmastlock_p & df54de | !hmastlock_p & v845542;
assign ad4f52 = hbusreq1_p & df5147 | !hbusreq1_p & !v845542;
assign dc4f83 = hmaster0_p & dc4f73 | !hmaster0_p & dc4f82;
assign hgrant2 = !bd5942;
assign d354e6 = hgrant1_p & d354e5 | !hgrant1_p & d354c4;
assign ade58f = locked_p & adec8f | !locked_p & !v845542;
assign b57504 = hready_p & b57a12 | !hready_p & b57503;
assign c3d70b = hbusreq1_p & c3d696 | !hbusreq1_p & c3d685;
assign dc4fd2 = hbusreq2 & dc4fcf | !hbusreq2 & dc4fd1;
assign ad46ae = hready & ad4697 | !hready & ad46ad;
assign v9f7715 = hbusreq2_p & v9f7710 | !hbusreq2_p & v9f7714;
assign c3ce66 = hgrant1_p & c3ce63 | !hgrant1_p & c3ce65;
assign v9f77ad = hbusreq0_p & v845542 | !hbusreq0_p & v9f779d;
assign d35a93 = hgrant3_p & d3597e | !hgrant3_p & d35a92;
assign df5171 = hbusreq1_p & df5170 | !hbusreq1_p & v845542;
assign c3d5b7 = hgrant0_p & v845542 | !hgrant0_p & !c3d5b1;
assign v9e9ee9 = hmaster2_p & v9e9ee7 | !hmaster2_p & v9ea3fb;
assign c3d589 = hgrant3_p & c3d535 | !hgrant3_p & c3d588;
assign b5741e = hmaster2_p & b57419 | !hmaster2_p & b5741d;
assign b1c70f = hlock0_p & bd572e | !hlock0_p & b1c70e;
assign ad4f98 = hmaster2_p & ad4f95 | !hmaster2_p & ad4f97;
assign d3563c = locked_p & d3563b | !locked_p & v845542;
assign c3d47e = hbusreq2 & c3d479 | !hbusreq2 & c3d47c;
assign v9f7dcc = stateG10_4_p & v9f7d42 | !stateG10_4_p & v9f7dcb;
assign ad4286 = hbusreq3 & ad4e65 | !hbusreq3 & !v845542;
assign c3d352 = hmaster0_p & c3d349 | !hmaster0_p & c3d351;
assign ad4ee5 = hgrant4_p & ad4ecd | !hgrant4_p & ad4ee3;
assign v9f7d0f = hlock2 & v9f7d05 | !hlock2 & v9f7d0e;
assign ba05cf = hready_p & v845550 | !hready_p & ba05ce;
assign b0595e = hlock4 & b0595b | !hlock4 & b0595d;
assign c3d713 = hmaster1_p & c3d712 | !hmaster1_p & c3d69b;
assign d3543e = hmaster0_p & d3542e | !hmaster0_p & d35429;
assign v9f77c8 = hmaster2_p & v9f77c7 | !hmaster2_p & !v845542;
assign ad3d2c = hmaster0_p & ad3d2b | !hmaster0_p & ad4411;
assign d356b6 = hbusreq1_p & d356b5 | !hbusreq1_p & v845542;
assign dc4f9c = hburst1 & dc4f9b | !hburst1 & v845566;
assign v9f7cc9 = hlock0 & v9f7cc8 | !hlock0 & v9f7cc4;
assign b1c6f8 = hbusreq1_p & b1c6b9 | !hbusreq1_p & b1c85f;
assign ad4800 = hgrant2_p & ad47fe | !hgrant2_p & ad47ff;
assign ad455d = hbusreq4_p & ad455c | !hbusreq4_p & v845542;
assign ad4dde = hburst0 & dc4f79 | !hburst0 & adea86;
assign b1c7e5 = hgrant2_p & b1c791 | !hgrant2_p & b1c7e4;
assign b05a91 = hmaster1_p & b05a90 | !hmaster1_p & b05a20;
assign cc36fb = hbusreq4_p & dc500e | !hbusreq4_p & cc36fa;
assign d35633 = hready_p & d355b0 | !hready_p & d35632;
assign d3552b = hmaster0_p & d35524 | !hmaster0_p & d3552a;
assign ad4567 = hlock4_p & ad4566 | !hlock4_p & v845542;
assign d357d4 = hlock1_p & d3577b | !hlock1_p & v84554a;
assign dc53ce = decide_p & dc53cb | !decide_p & v845542;
assign ade574 = hmaster2_p & v845558 | !hmaster2_p & ade573;
assign b1cc03 = hmaster1_p & b1cfb8 | !hmaster1_p & b1cc02;
assign d35771 = hbusreq0 & d35770 | !hbusreq0 & v845542;
assign d35ab9 = hbusreq2_p & d35aa9 | !hbusreq2_p & !d35ab8;
assign ade595 = hgrant0_p & adec9a | !hgrant0_p & v84556c;
assign ad42d1 = hbusreq1_p & ad42d0 | !hbusreq1_p & c3d2d9;
assign v8cc474 = hmaster2_p & v8cc473 | !hmaster2_p & v845542;
assign v9f76d5 = hmaster0_p & v9f7e0d | !hmaster0_p & v9f7d9f;
assign dc53b2 = decide_p & dc53a8 | !decide_p & v845542;
assign c3cf2d = hmaster0_p & c3d5ec | !hmaster0_p & c3d306;
assign v9f7ce3 = hlock1 & v9f7cdd | !hlock1 & v9f7ce2;
assign ad413b = hlock4_p & ad413a | !hlock4_p & !ad4e9a;
assign b05a93 = hmaster0_p & b0593d | !hmaster0_p & b05a0f;
assign ade5c4 = hbusreq3 & ade5ab | !hbusreq3 & !v845558;
assign c3d709 = hmaster2_p & c3d669 | !hmaster2_p & !c3d6e6;
assign dc53d1 = hbusreq3_p & dc53d0 | !hbusreq3_p & !dc5088;
assign c3d388 = hmaster0_p & v845555 | !hmaster0_p & v845551;
assign ad4f4f = hmaster0_p & ad4f47 | !hmaster0_p & ad4f4e;
assign dc4fa7 = hlock0_p & dc4f9d | !hlock0_p & !v845542;
assign v9f7d63 = hmaster2_p & v9f7d60 | !hmaster2_p & v9f7d62;
assign d35a56 = hmastlock_p & adea97 | !hmastlock_p & !d359ba;
assign v8cc604 = hbusreq3_p & v8cc5c9 | !hbusreq3_p & v8cc603;
assign c3d5eb = hbusreq4 & c3d5e8 | !hbusreq4 & !c3d5ea;
assign start = ac1495;
assign ad47f7 = hbusreq2_p & ad47f2 | !hbusreq2_p & !ad47f6;
assign v9f7c96 = stateG2_p & v845542 | !stateG2_p & v9f7c95;
assign bd593c = decide_p & bd593b | !decide_p & v845572;
assign ad43df = hlock1_p & ad43d9 | !hlock1_p & ad43de;
assign ad4fe2 = stateG10_4_p & v84556c | !stateG10_4_p & !ad4fe1;
assign v9f76fc = hbusreq1_p & v9f7db4 | !hbusreq1_p & v9f76f2;
assign c3d2d6 = hready & v845564 | !hready & !v845542;
assign ad4324 = hbusreq1_p & ad4323 | !hbusreq1_p & v845542;
assign ad4f58 = hgrant1_p & ad4f56 | !hgrant1_p & ad4f57;
assign ad446f = hlock2_p & ad446b | !hlock2_p & ad446e;
assign ad4587 = hbusreq3 & ad4586 | !hbusreq3 & !v845547;
assign v9ea5b1 = hbusreq2 & v9ea5b0 | !hbusreq2 & v9ea586;
assign c3d3ab = hready_p & c3d3aa | !hready_p & c3d393;
assign d3591b = hmaster2_p & adea8a | !hmaster2_p & !d3591a;
assign v8cc5bf = hbusreq3 & v8cc5bd | !hbusreq3 & v8cc5be;
assign b058d5 = hmaster2_p & b058d2 | !hmaster2_p & b058d4;
assign bd576e = hbusreq2 & bd576d | !hbusreq2 & v845542;
assign b57ae2 = hlock3 & b579c5 | !hlock3 & b579c4;
assign d356a6 = hbusreq1 & d356a5 | !hbusreq1 & v845542;
assign ad4e24 = hmaster1_p & ad4e21 | !hmaster1_p & ad4e23;
assign dc4fe0 = hmaster2_p & c3d66d | !hmaster2_p & v845542;
assign b05a82 = hmaster1_p & b05a78 | !hmaster1_p & b05a81;
assign ad43fa = hbusreq4 & ad43f5 | !hbusreq4 & !ad43f9;
assign bd56de = hbusreq2_p & bd56dd | !hbusreq2_p & v845542;
assign c3d5dc = hbusreq4_p & c3d5da | !hbusreq4_p & !c3d5db;
assign d3578e = hlock0_p & v845542 | !hlock0_p & !d35617;
assign adea92 = hgrant4_p & v84556c | !hgrant4_p & !v845542;
assign b1cfc1 = hlock0_p & b1cfc0 | !hlock0_p & !v845542;
assign v9f77ba = hready_p & v9f7740 | !hready_p & v9f77b9;
assign d35707 = hbusreq1 & d35a18 | !hbusreq1 & v845542;
assign ad475c = hmaster1_p & ad475b | !hmaster1_p & ad4591;
assign v9ea5a1 = hready & v9ea5a0 | !hready & v9ea59b;
assign c3d38e = hmaster0_p & c3d38c | !hmaster0_p & c3d38d;
assign bd5739 = stateA1_p & v8ccb68 | !stateA1_p & !bd5738;
assign b1cbfa = hmaster2_p & b1cfb7 | !hmaster2_p & b1cbf9;
assign dc4fb0 = hbusreq4 & dc4fab | !hbusreq4 & dc4faf;
assign v9ea476 = hbusreq0 & v9ea475 | !hbusreq0 & v9ea46d;
assign c3d739 = hgrant2_p & c3d738 | !hgrant2_p & !c3d735;
assign d3501d = hgrant1_p & d35018 | !hgrant1_p & d3501c;
assign v9ea590 = hbusreq4_p & v9ea458 | !hbusreq4_p & v9ea4c8;
assign ad43d0 = hlock0_p & d35616 | !hlock0_p & !ad43cf;
assign b05969 = hlock1_p & b058b1 | !hlock1_p & b058f1;
assign ad3cfb = hready & ad3cfa | !hready & !ad3cd7;
assign c3d712 = hmaster0_p & c3d697 | !hmaster0_p & c3d685;
assign c3d4fd = hbusreq0 & c3d4fb | !hbusreq0 & c3d4fc;
assign ad5034 = hready & ad5030 | !hready & !ad5033;
assign v8cc4ed = hbusreq4_p & v8d29fa | !hbusreq4_p & v8d29fb;
assign v9f76aa = hmaster1_p & v9f76a9 | !hmaster1_p & v9f7d64;
assign cc3706 = hgrant2_p & cc36d3 | !hgrant2_p & !cc3705;
assign b1c79f = hgrant4_p & c3d66d | !hgrant4_p & !b1c79d;
assign c3d753 = hgrant2_p & c3d751 | !hgrant2_p & c3d752;
assign v9f77e2 = hgrant1_p & v9f77d6 | !hgrant1_p & v9f77e1;
assign c3d6b5 = hmaster2_p & c3d669 | !hmaster2_p & !c3d6b4;
assign ad4700 = hbusreq4_p & ad46ff | !hbusreq4_p & v845542;
assign ad4148 = hmaster1_p & ad410c | !hmaster1_p & ad4147;
assign c3d717 = hgrant2_p & c3d713 | !hgrant2_p & c3d716;
assign d35796 = hmaster0_p & d35791 | !hmaster0_p & d35795;
assign ade61b = hbusreq2 & ade5ab | !hbusreq2 & !v845558;
assign c3ce1e = hbusreq2 & c3d37f | !hbusreq2 & c3d2de;
assign df54ed = hgrant2_p & df54eb | !hgrant2_p & df54db;
assign ad42df = hlock1_p & ad42de | !hlock1_p & ad4267;
assign v9f7cc2 = hbusreq2 & v9f7cc0 | !hbusreq2 & v9f7cc1;
assign v9ea461 = hbusreq2 & v9ea45f | !hbusreq2 & v9ea460;
assign ad5024 = hgrant1_p & v845547 | !hgrant1_p & ad5023;
assign b1c7bd = hgrant4_p & b1c720 | !hgrant4_p & !b1c7bc;
assign ad42b0 = hbusreq4_p & ad45ae | !hbusreq4_p & !v845542;
assign d354b3 = hgrant4_p & v845542 | !hgrant4_p & !d354b2;
assign ad4fc5 = hmaster0_p & ad4fc0 | !hmaster0_p & ad4fc4;
assign v8cc4db = hbusreq2_p & v8cc4b3 | !hbusreq2_p & v8cc4da;
assign dc5003 = hgrant4_p & adec89 | !hgrant4_p & ade563;
assign c3d6a5 = hgrant0_p & c3d66a | !hgrant0_p & !c3d669;
assign d35790 = hbusreq0 & d3578f | !hbusreq0 & v845542;
assign b1c03d = hmaster0_p & b1c03b | !hmaster0_p & b1c03c;
assign c3d513 = hgrant1_p & v845564 | !hgrant1_p & c3d512;
assign d35a5d = hlock0_p & d35a5c | !hlock0_p & !ade562;
assign df515a = hbusreq3 & df5157 | !hbusreq3 & df5159;
assign v9ea586 = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea585;
assign d35761 = hready_p & d35760 | !hready_p & d3575d;
assign d35688 = hgrant3_p & d35633 | !hgrant3_p & d35687;
assign ad42ef = hbusreq1 & ad4e91 | !hbusreq1 & v845542;
assign c3d33a = hmaster2_p & c3d339 | !hmaster2_p & v845542;
assign c3d72d = hmaster0_p & c3d685 | !hmaster0_p & c3d699;
assign b57946 = hready_p & b578f5 | !hready_p & b57945;
assign c3d2d1 = hmaster0_p & c3d2d0 | !hmaster0_p & c3d2be;
assign b57a21 = hbusreq2_p & b5790a | !hbusreq2_p & b57a20;
assign d35757 = hgrant2_p & d3574e | !hgrant2_p & !d35756;
assign c3d2b0 = hburst0 & c3d2ae | !hburst0 & c3d2af;
assign df5535 = hmaster0_p & df5534 | !hmaster0_p & df5532;
assign v9e9ea7 = hbusreq1_p & v9ea46d | !hbusreq1_p & v9ea4d9;
assign ad4faa = hlock3_p & ad4f32 | !hlock3_p & ad4fa9;
assign ad48b5 = hbusreq1 & ad48a6 | !hbusreq1 & ad48b1;
assign d35702 = hgrant1_p & v845542 | !hgrant1_p & d35701;
assign ad45a2 = hmaster2_p & v845542 | !hmaster2_p & ad45a1;
assign ad4375 = hbusreq2_p & ad4370 | !hbusreq2_p & ad4374;
assign b05916 = hmaster1_p & b05915 | !hmaster1_p & b05913;
assign ade548 = hbusreq4_p & c3d66d | !hbusreq4_p & v845542;
assign b57420 = hbusreq0 & b5741e | !hbusreq0 & b5741f;
assign ad506a = hmaster0_p & ad5013 | !hmaster0_p & ad5069;
assign v9e9f81 = hgrant1_p & v9e9f72 | !hgrant1_p & v9e9f80;
assign dc531e = hlock3_p & dc531d | !hlock3_p & v845542;
assign c3d5a7 = hbusreq2 & c3d5a0 | !hbusreq2 & v845542;
assign ad4db4 = hmaster2_p & ad4db2 | !hmaster2_p & ad4daf;
assign v9ea4d6 = hgrant4_p & v9ea4bb | !hgrant4_p & v9ea4d5;
assign c3d347 = hready & c3d346 | !hready & c3d300;
assign v8cc4b0 = hbusreq2 & v8cc4ae | !hbusreq2 & v8cc4af;
assign bd57f1 = hbusreq1 & bd574d | !hbusreq1 & v84556c;
assign ad4fd1 = hbusreq1_p & ad4fb0 | !hbusreq1_p & ad4fd0;
assign ad4db9 = hmaster0_p & ad4da4 | !hmaster0_p & ad4db8;
assign b573da = hlock3 & b579e5 | !hlock3 & b573d9;
assign c3cf1c = hbusreq3 & c3cf1b | !hbusreq3 & c3cee4;
assign ad42e8 = hmaster0_p & ad42e6 | !hmaster0_p & ad42e7;
assign c3d36a = hmaster0_p & c3d368 | !hmaster0_p & c3d369;
assign v9e9e7d = decide_p & v9e9e75 | !decide_p & v9e9e7c;
assign ad46b7 = hlock4_p & ad4ebf | !hlock4_p & v845542;
assign dc5019 = hmaster2_p & c3d66d | !hmaster2_p & !ade56d;
assign df517b = hbusreq1_p & df517a | !hbusreq1_p & v845542;
assign c3ce37 = hbusreq1_p & c3ce36 | !hbusreq1_p & !v845542;
assign dc5392 = hlock3_p & dc5391 | !hlock3_p & !v845542;
assign ad3d17 = hmaster1_p & ad3d16 | !hmaster1_p & ad4419;
assign d35752 = hgrant1_p & d35aa4 | !hgrant1_p & d35751;
assign c3d686 = hbusreq1_p & c3d683 | !hbusreq1_p & c3d685;
assign b57a20 = hmaster1_p & b57a1d | !hmaster1_p & b57a1f;
assign b1c7e3 = hmaster0_p & b1c7cb | !hmaster0_p & b1c7e2;
assign c3cefb = hmaster1_p & c3cef9 | !hmaster1_p & c3cefa;
assign c3d726 = decide_p & c3d720 | !decide_p & !c3d725;
assign d359fa = hlock4_p & d359f8 | !hlock4_p & d359f9;
assign b05a4c = hready_p & b05a37 | !hready_p & !b05a4b;
assign c3cebd = hgrant4_p & v845542 | !hgrant4_p & c3cebc;
assign v9f7d49 = hmaster0_p & v9f7d3b | !hmaster0_p & v9f7d3c;
assign b0592c = hmaster1_p & b0592b | !hmaster1_p & b05926;
assign b1c73b = hmaster0_p & b1c737 | !hmaster0_p & b1c73a;
assign d35646 = hbusreq1 & d355a3 | !hbusreq1 & d355a9;
assign ade5d5 = hlock0_p & ade5ce | !hlock0_p & ade4e7;
assign bd585d = hlock4_p & bd585b | !hlock4_p & bd585c;
assign v9f772c = hmaster2_p & v9f772b | !hmaster2_p & d359c4;
assign v845542 = 1;
assign v9f7cd8 = hlock0_p & v9f7cb4 | !hlock0_p & v9f7cd7;
assign b5798a = hmaster1_p & b5794b | !hmaster1_p & b57989;
assign b574fb = decide_p & b57940 | !decide_p & b574fa;
assign b1c612 = hgrant3_p & b1c5fe | !hgrant3_p & b1c611;
assign b1c78a = hready_p & b1c74c | !hready_p & !b1c789;
assign b1c81e = hbusreq0 & b1c81d | !hbusreq0 & !d35a9c;
assign c5c96e = hgrant0_p & c5c8e7 | !hgrant0_p & c5c896;
assign dc5081 = hbusreq2_p & dc5069 | !hbusreq2_p & dc5080;
assign v9f7ca0 = locked_p & v9f7c9d | !locked_p & !v9f7c9f;
assign v9ea627 = decide_p & v9ea61f | !decide_p & v9ea626;
assign c3d2df = hbusreq3 & c3d2dd | !hbusreq3 & c3d2de;
assign d357a7 = hmaster1_p & d35796 | !hmaster1_p & d357a6;
assign ad4300 = hmaster0_p & ad4f19 | !hmaster0_p & !ad42ff;
assign ad4589 = hmaster0_p & ad4587 | !hmaster0_p & ad4588;
assign v9f7de7 = hmaster2_p & v9f7ddc | !hmaster2_p & v9f7de6;
assign ad43fc = hmaster0_p & ad43e0 | !hmaster0_p & ad43fb;
assign c3d6af = stateG10_4_p & c3d6ac | !stateG10_4_p & !c3d6ae;
assign c3d6e6 = hbusreq4_p & c3d6e4 | !hbusreq4_p & c3d6e5;
assign v9f7ce9 = hmaster0_p & v9f7cd5 | !hmaster0_p & !v9f7ce8;
assign b05978 = hgrant4_p & b058a7 | !hgrant4_p & !b05954;
assign ad4752 = hmaster1_p & ad4751 | !hmaster1_p & ad460e;
assign v9e9f8b = hgrant4_p & v9e9f67 | !hgrant4_p & v9e9f74;
assign b1c736 = hbusreq0 & b1c735 | !hbusreq0 & !v845542;
assign v9f7d6e = hbusreq1_p & v9f7d6d | !hbusreq1_p & v9f7d0c;
assign v9e9fd1 = hmaster1_p & v9ea44a | !hmaster1_p & v9e9fd0;
assign v9ea40a = decide_p & v9ea3f9 | !decide_p & v9ea409;
assign v8cc0ec = hbusreq1 & v8cc0ce | !hbusreq1 & v8cc0cf;
assign dc5009 = hgrant4_p & v84556c | !hgrant4_p & adec89;
assign v8cc509 = hmaster1_p & v8cc475 | !hmaster1_p & v8cc508;
assign df51a8 = hbusreq3 & df5195 | !hbusreq3 & !v84554c;
assign b1c76c = hbusreq1_p & b1c766 | !hbusreq1_p & b1c76b;
assign d354c3 = hbusreq0 & d354c2 | !hbusreq0 & d354aa;
assign b1c04c = hready_p & b1c824 | !hready_p & !b1c04b;
assign d35735 = decide_p & d35734 | !decide_p & !v84556c;
assign ad4e6f = hlock0_p & ad4e6d | !hlock0_p & !ad4e6e;
assign bd5b95 = hbusreq3 & d35a50 | !hbusreq3 & bd5b94;
assign c3d2af = hburst1 & c3d2ae | !hburst1 & v845566;
assign v9f77fc = hbusreq3 & v9f77f9 | !hbusreq3 & v9f77fb;
assign stateG10_1 = !ad13e5;
assign d356f9 = hmaster0_p & d356f3 | !hmaster0_p & d356f8;
assign b058cb = hbusreq3 & b058c8 | !hbusreq3 & b058ca;
assign ad4560 = hready & ad4557 | !hready & ad455f;
assign ad4691 = hlock4_p & ad4e7c | !hlock4_p & b1cfcb;
assign b05a2f = hmaster0_p & b058e8 | !hmaster0_p & b058c7;
assign ad435a = decide_p & ad42ce | !decide_p & ad4359;
assign dc4f8c = hbusreq3 & dc4f8b | !hbusreq3 & v845542;
assign b5795a = hgrant2_p & v845542 | !hgrant2_p & b57958;
assign b574cf = hmaster0_p & b574bf | !hmaster0_p & b574ce;
assign ad4f3d = hmaster2_p & v845542 | !hmaster2_p & ad4f36;
assign d357fa = hmaster2_p & v845558 | !hmaster2_p & d35a9c;
assign v9f780e = hbusreq4_p & v9f780c | !hbusreq4_p & !v9f780d;
assign ad4f44 = hready & dc4fcb | !hready & v84556c;
assign dc507b = hbusreq1_p & dc5079 | !hbusreq1_p & dc507a;
assign ad4dac = hbusreq4_p & dc4f78 | !hbusreq4_p & !v845542;
assign d3575c = hbusreq3_p & d35725 | !hbusreq3_p & !d3575b;
assign bd58a3 = hgrant0_p & v84556c | !hgrant0_p & !bd58a2;
assign dc5052 = hgrant4_p & ade572 | !hgrant4_p & !adeca1;
assign df50cc = hlock1_p & df50cb | !hlock1_p & !v845542;
assign ade4b6 = hburst1_p & v8f2540 | !hburst1_p & !c74a04;
assign c5c8ee = hready_p & c5c893 | !hready_p & !c5c8ed;
assign ad4e53 = hmastlock_p & d359c8 | !hmastlock_p & v845542;
assign dc4ff9 = hbusreq4 & dc4fed | !hbusreq4 & dc4ff8;
assign v9f7dea = hlock4 & v9f7de7 | !hlock4 & v9f7de9;
assign c3d311 = hbusreq0 & v845542 | !hbusreq0 & v8da5a1;
assign c3ce72 = decide_p & c3ce40 | !decide_p & !c3ce71;
assign c3d30d = hgrant4_p & v845542 | !hgrant4_p & ade562;
assign ad475e = hmaster0_p & ad470d | !hmaster0_p & ad459e;
assign d35953 = hbusreq3 & d35952 | !hbusreq3 & v845542;
assign bd5b8e = hgrant2_p & bd5b8d | !hgrant2_p & !v845542;
assign ad45a0 = hbusreq1_p & ad459e | !hbusreq1_p & ad456f;
assign b05a05 = locked_p & b0591c | !locked_p & b05938;
assign c3d737 = hmaster0_p & c3d685 | !hmaster0_p & c3d682;
assign bd587e = hgrant4_p & bd587d | !hgrant4_p & adec89;
assign df51c5 = hgrant1_p & df5538 | !hgrant1_p & !df5183;
assign b1c4ae = hmaster0_p & v845542 | !hmaster0_p & b1c4a7;
assign ad3d37 = hmaster1_p & ad3d36 | !hmaster1_p & ad4469;
assign b1cf2c = hbusreq0 & b1cf2a | !hbusreq0 & b1cf2b;
assign ad40e9 = hlock2_p & ad4898 | !hlock2_p & !ad40e8;
assign ad4e90 = hbusreq4 & ad4e88 | !hbusreq4 & ad4e8f;
assign dc5014 = hbusreq4 & dc5008 | !hbusreq4 & dc5013;
assign bd5779 = hmaster0_p & bd5776 | !hmaster0_p & bd5778;
assign b1c84e = decide_p & b1c84d | !decide_p & v845542;
assign v8cc497 = hbusreq0_p & v8cc492 | !hbusreq0_p & v8cc496;
assign b05930 = hmaster1_p & b0591e | !hmaster1_p & b05926;
assign b579f1 = hmaster1_p & b579f0 | !hmaster1_p & v845542;
assign v8cc128 = hmaster0_p & v8cc127 | !hmaster0_p & v845542;
assign c5c89c = hbusreq4_p & c5c89b | !hbusreq4_p & !v845542;
assign v9f7665 = stateG10_4_p & v9f7663 | !stateG10_4_p & v9f7664;
assign b579b9 = hmastlock_p & b579b8 | !hmastlock_p & v845542;
assign v9e9f55 = stateG10_4_p & v9ea441 | !stateG10_4_p & v9e9f54;
assign c3d5d6 = stateG10_4_p & c3d5d4 | !stateG10_4_p & c3d5d5;
assign v9f7cca = hbusreq0 & v9f7cc4 | !hbusreq0 & v9f7cc9;
assign df51c8 = hgrant2_p & df51c2 | !hgrant2_p & !df51c7;
assign d35807 = hlock0_p & v845542 | !hlock0_p & !d35806;
assign v9ea605 = hbusreq1_p & v9ea43b | !hbusreq1_p & v9ea604;
assign dc4f6e = hbusreq1 & dc4f68 | !hbusreq1 & dc4f6a;
assign d35693 = hbusreq2 & d35aae | !hbusreq2 & d35ab4;
assign ad4426 = hmaster1_p & ad4422 | !hmaster1_p & ad4425;
assign b059ab = hmaster1_p & b059aa | !hmaster1_p & b059a0;
assign c3d5cf = hbusreq2 & c3d353 | !hbusreq2 & c3d32f;
assign bd5915 = hbusreq1 & d35a50 | !hbusreq1 & bd5b94;
assign ad501f = hmaster1_p & ad501a | !hmaster1_p & ad501e;
assign dc5035 = hbusreq1_p & dc5031 | !hbusreq1_p & dc5034;
assign v9e9f4f = hlock0_p & v9e9f4d | !hlock0_p & v9e9f4e;
assign df512d = decide_p & df511b | !decide_p & d6ebca;
assign c3d371 = hmastlock_p & c3d370 | !hmastlock_p & !v845542;
assign dc4fb4 = hbusreq3 & dc4fa3 | !hbusreq3 & v845542;
assign d359af = hlock1_p & d35991 | !hlock1_p & !d359ae;
assign v9e9e9f = hmaster2_p & v9e9e9e | !hmaster2_p & v9ea448;
assign v9f77f2 = hmaster2_p & v9f77ea | !hmaster2_p & !v9f77f1;
assign v8cc78e = decide_p & v8cc4f4 | !decide_p & v8cc782;
assign d359fe = hgrant4_p & d359c9 | !hgrant4_p & v845542;
assign ad4dea = hbusreq3 & ad4de9 | !hbusreq3 & !v845542;
assign v9e9ed9 = hbusreq3_p & v9e9ec1 | !hbusreq3_p & v9e9ed8;
assign v9e9eb5 = hbusreq2 & v9e9eb4 | !hbusreq2 & v9ea4cd;
assign v8cc7c1 = hlock0 & v8ccbf4 | !hlock0 & v8cc7c0;
assign ad42a6 = hbusreq3 & ad42a1 | !hbusreq3 & ad42a5;
assign ad43c8 = hbusreq0 & ad43c7 | !hbusreq0 & v845542;
assign v8cc620 = hbusreq3 & v8cc4ac | !hbusreq3 & v8cc61e;
assign c3d68e = hmaster1_p & c3d68d | !hmaster1_p & c3d68b;
assign c3ceaa = hready_p & c3ce9a | !hready_p & c3cea9;
assign ad4763 = decide_p & ad475d | !decide_p & !ad4762;
assign df5118 = hbusreq1_p & df5117 | !hbusreq1_p & v845542;
assign dc4fe2 = hbusreq1_p & dc4fdf | !hbusreq1_p & dc4fe1;
assign bd592e = hbusreq0_p & d35a58 | !hbusreq0_p & dc52fa;
assign b57a27 = hbusreq1_p & b5794a | !hbusreq1_p & b57a26;
assign v9f7799 = hbusreq3 & v9f7797 | !hbusreq3 & v9f7798;
assign d357bf = hlock1_p & d35778 | !hlock1_p & v84554a;
assign b058ee = hbusreq4 & b058ec | !hbusreq4 & b058ed;
assign ad13e4 = hready_p & ad13e2 | !hready_p & ad13e3;
assign c3cedd = hbusreq0_p & c3d59e | !hbusreq0_p & v845542;
assign b1c777 = hbusreq2 & b1c762 | !hbusreq2 & b1c764;
assign ad4ecf = hready & ad4ece | !hready & !v845542;
assign v9f7792 = hlock0 & v9f772d | !hlock0 & v9f7791;
assign d35a0e = hgrant4_p & v845542 | !hgrant4_p & d359f7;
assign b1d00e = hgrant1_p & v845542 | !hgrant1_p & v8da59f;
assign b05a5b = hgrant0_p & b058a3 | !hgrant0_p & b05a5a;
assign v9f7ce0 = hlock4 & v9f7cdd | !hlock4 & v9f7cdf;
assign ad4486 = hbusreq0 & ad4485 | !hbusreq0 & v845542;
assign bd5928 = hmaster0_p & v845542 | !hmaster0_p & bd5927;
assign ad46ed = hmaster1_p & ad46e9 | !hmaster1_p & ad46ec;
assign v9ea4cd = hbusreq1_p & v9ea3fa | !hbusreq1_p & v9ea4b4;
assign c3ce58 = hgrant1_p & v84554d | !hgrant1_p & c3ce57;
assign ad4372 = hmaster1_p & ad4371 | !hmaster1_p & ad4297;
assign d354eb = decide_p & d354ea | !decide_p & v84556c;
assign c3d386 = hready_p & c3d364 | !hready_p & c3d385;
assign v9f7d40 = hlock4_p & v9f7c9d | !hlock4_p & v9ea3ec;
assign d35a58 = locked_p & d35a57 | !locked_p & !v845542;
assign d35a36 = hbusreq2_p & d35a28 | !hbusreq2_p & !d35a35;
assign v9e9fc4 = hgrant2_p & v9e9fc1 | !hgrant2_p & v9e9fc3;
assign ad442c = hgrant4_p & b1c714 | !hgrant4_p & v845542;
assign c3d36c = hmaster1_p & c3d36a | !hmaster1_p & c3d36b;
assign d3570c = hmaster1_p & d35702 | !hmaster1_p & d3570b;
assign v9f7d2e = hbusreq2 & v9f7d2c | !hbusreq2 & !v9f7d2d;
assign ad46ec = hmaster0_p & ad46ea | !hmaster0_p & !ad46eb;
assign ad4d91 = hmastlock_p & ad4d90 | !hmastlock_p & v845542;
assign bd5850 = stateG10_4_p & bd5842 | !stateG10_4_p & !bd584f;
assign ad4f0d = hbusreq4_p & ad4f0c | !hbusreq4_p & adeaa4;
assign c3d2e7 = hburst1 & c3d2e6 | !hburst1 & v845542;
assign c5c8f3 = hgrant4_p & v845542 | !hgrant4_p & c5c8f2;
assign bd5818 = hmaster2_p & bd5817 | !hmaster2_p & dc500c;
assign b1c716 = hlock0_p & bd5744 | !hlock0_p & !b1c715;
assign ad4145 = hgrant1_p & ad40ff | !hgrant1_p & ad4144;
assign v9f7e3d = stateG10_4_p & v9f7dad | !stateG10_4_p & v9f7e3c;
assign dc531c = hmaster0_p & dc531b | !hmaster0_p & v845542;
assign v9f77cb = hlock4 & v9f77c8 | !hlock4 & v9f77ca;
assign b1c0b1 = hgrant3_p & b1c84f | !hgrant3_p & b1c0b0;
assign ad40f6 = hbusreq2 & ad501b | !hbusreq2 & v845542;
assign ad4dc6 = hready & ad4d96 | !hready & !ad4dc5;
assign ad4dd4 = hready & ad4dab | !hready & ad4dd3;
assign v9e9fc5 = hmaster0_p & v9e9eed | !hmaster0_p & v9e9fa6;
assign b579da = hmaster2_p & b579d8 | !hmaster2_p & b579d2;
assign ad45fa = hbusreq2 & ad45c6 | !hbusreq2 & ad45c9;
assign v8ccb76 = hlock1_p & v8d29fa | !hlock1_p & v8ccb75;
assign ad4731 = hbusreq4 & v845542 | !hbusreq4 & c3d327;
assign bd58fb = hmaster0_p & bd58fa | !hmaster0_p & bd5831;
assign df5196 = hbusreq2 & df5195 | !hbusreq2 & !v84554c;
assign df5131 = decide_p & df5130 | !decide_p & d6ebca;
assign dc5047 = hgrant4_p & ade581 | !hgrant4_p & ade59c;
assign ad46e7 = hbusreq2 & ad4586 | !hbusreq2 & !v845542;
assign v8cc7ef = hgrant4_p & v8cc7dd | !hgrant4_p & v845542;
assign v9f76ac = hmaster0_p & v9f7691 | !hmaster0_p & v9f76ab;
assign v9ea43a = hmaster2_p & v9ea439 | !hmaster2_p & v9ea3fb;
assign v8ccbd9 = hmaster0_p & v8ccbd8 | !hmaster0_p & v845542;
assign ad3d5e = jx1_p & ad3d5d | !jx1_p & ad48ca;
assign df50d0 = hmaster1_p & df54f4 | !hmaster1_p & df50cf;
assign d3561c = stateA1_p & d3561b | !stateA1_p & ade4b7;
assign dc5389 = hmaster2_p & v84556c | !hmaster2_p & adea9a;
assign ba7c64 = hbusreq4_p & v845542 | !hbusreq4_p & v845576;
assign b57a76 = hlock0 & b579ce | !hlock0 & b57a75;
assign df5533 = hbusreq1 & v84556c | !hbusreq1 & v845542;
assign bd58bb = hbusreq4_p & bd58ba | !hbusreq4_p & bd58aa;
assign v9f7650 = hlock2 & v9f764d | !hlock2 & v9f764f;
assign v8cc4ae = hbusreq3 & v8cc4ac | !hbusreq3 & v8cc4ad;
assign ac1478 = stateG10_4_p & ac1465 | !stateG10_4_p & !ac1477;
assign b8ef50 = hgrant3_p & b8f6e0 | !hgrant3_p & b8f74d;
assign v9f76f1 = hbusreq4_p & v9f7d86 | !hbusreq4_p & v9f76f0;
assign v9f7733 = hbusreq0_p & v845542 | !hbusreq0_p & !v9f772f;
assign d35717 = hlock1_p & d359ca | !hlock1_p & v845542;
assign bd58d4 = hgrant1_p & df5538 | !hgrant1_p & bd58d3;
assign ad480e = hbusreq2 & ad480d | !hbusreq2 & v845542;
assign d357ca = stateG10_4_p & d3576e | !stateG10_4_p & d357c8;
assign ad4f12 = hbusreq4 & ad4f06 | !hbusreq4 & ad4f11;
assign ad4fa8 = hgrant2_p & v845542 | !hgrant2_p & !ad4fa7;
assign ad3d1d = hgrant2_p & ad3d17 | !hgrant2_p & ad3d1c;
assign ad430d = hmaster0_p & ad42ee | !hmaster0_p & ad430c;
assign v9f764e = hlock3 & v9f764d | !hlock3 & v9f764a;
assign ad4582 = hmaster0_p & ad456c | !hmaster0_p & ad4581;
assign b57906 = hbusreq2_p & b57905 | !hbusreq2_p & b57904;
assign d359cf = hgrant4_p & d35983 | !hgrant4_p & d359ce;
assign b1cfce = hbusreq4_p & b1cfcc | !hbusreq4_p & !b1cfcd;
assign ade5a6 = hgrant2_p & ade546 | !hgrant2_p & ade5a5;
assign v9f7cfe = hlock1 & v9f7cf8 | !hlock1 & v9f7cfd;
assign b1c7f3 = hbusreq1 & b1c73e | !hbusreq1 & !v845542;
assign ad4811 = hbusreq3 & ad4810 | !hbusreq3 & v845542;
assign c3d6c1 = hgrant4_p & c3d66e | !hgrant4_p & !c3d6ac;
assign d35a18 = hbusreq4 & d35a0a | !hbusreq4 & d35a17;
assign dc4faa = hmaster2_p & dc4fa6 | !hmaster2_p & !dc4fa9;
assign adec98 = hburst1 & adea98 | !hburst1 & adec97;
assign c3ce7f = hbusreq1_p & c3ce43 | !hbusreq1_p & c3d3a3;
assign bd57ba = busreq_p & c5c88b | !busreq_p & ade4b8;
assign b05902 = hmaster0_p & b058f6 | !hmaster0_p & b05901;
assign ad4ef8 = hgrant4_p & v84556c | !hgrant4_p & ad4ef7;
assign b1cfc6 = hgrant4_p & v845542 | !hgrant4_p & !b1cfc5;
assign c5c999 = hgrant2_p & c5c97c | !hgrant2_p & c5c978;
assign adea93 = hlock4_p & adea92 | !hlock4_p & !v845542;
assign v9ea475 = hlock0 & v9ea46d | !hlock0 & v9ea474;
assign dc53c2 = hmaster0_p & dc53c1 | !hmaster0_p & v845542;
assign v9f7877 = hmaster1_p & v9f7876 | !hmaster1_p & v9f7736;
assign b05936 = stateA1_p & v845542 | !stateA1_p & !b058a0;
assign d359dd = stateG10_4_p & d359ce | !stateG10_4_p & d359dc;
assign v8cc0db = hbusreq0 & v8cc0da | !hbusreq0 & v8cc494;
assign v9e9f69 = hbusreq0_p & v9ea44c | !hbusreq0_p & v9ea4b3;
assign c3d75c = hmaster1_p & c3d75b | !hmaster1_p & c3d69b;
assign d35c03 = hmaster2_p & v84555a | !hmaster2_p & !d35c02;
assign b5794b = hgrant1_p & v845542 | !hgrant1_p & b5794a;
assign d35493 = hlock4_p & v845542 | !hlock4_p & dc52fa;
assign ad4825 = hmaster0_p & ad4823 | !hmaster0_p & ad4824;
assign c3ce14 = hbusreq2 & c3ce13 | !hbusreq2 & c3d368;
assign d359b9 = stateA1_p & v8ccb68 | !stateA1_p & !bb9bdd;
assign bd5834 = hbusreq1 & bd5768 | !hbusreq1 & !bd576c;
assign d35433 = hmaster2_p & v84555a | !hmaster2_p & d35432;
assign v9f7669 = hbusreq0 & v9f765c | !hbusreq0 & v9f7668;
assign c3d483 = decide_p & c3d482 | !decide_p & !c3d36c;
assign ad438d = hmaster2_p & ad4380 | !hmaster2_p & b1c714;
assign v9e9ef1 = hmaster0_p & v9e9eee | !hmaster0_p & v9e9ef0;
assign ad4288 = hbusreq3 & ad4287 | !hbusreq3 & v845542;
assign d35bf3 = hbusreq1_p & d35bed | !hbusreq1_p & d35bf2;
assign d356ab = hbusreq1_p & d356aa | !hbusreq1_p & v845542;
assign v9f7756 = hlock1 & v9f7751 | !hlock1 & v9f7755;
assign b1c867 = decide_p & b1c865 | !decide_p & b1c866;
assign bd5875 = hlock0_p & bd5871 | !hlock0_p & !bd5874;
assign bd58f0 = hmaster0_p & bd58ef | !hmaster0_p & bd5797;
assign ad5065 = hbusreq3 & ad5064 | !hbusreq3 & v845542;
assign d35025 = hbusreq3_p & d357e8 | !hbusreq3_p & d35024;
assign d3501a = hmaster2_p & d35019 | !hmaster2_p & d35aac;
assign v9f76ce = hmaster0_p & v9f7692 | !hmaster0_p & v9f7d5e;
assign ad4259 = hmaster1_p & ad4258 | !hmaster1_p & ad416b;
assign v8cc503 = hmaster1_p & v8cc500 | !hmaster1_p & v8cc502;
assign c3cee6 = hbusreq2 & c3cee0 | !hbusreq2 & c3cee4;
assign b57985 = hbusreq4_p & b5794f | !hbusreq4_p & b57984;
assign b1c860 = hbusreq1_p & b1c850 | !hbusreq1_p & b1c85f;
assign ad4e48 = hmaster2_p & d3597f | !hmaster2_p & ad4e47;
assign d354e4 = hlock1_p & d354e2 | !hlock1_p & !d354e3;
assign v9e9ed0 = hgrant2_p & v9e9ecd | !hgrant2_p & v9e9ecf;
assign d356bb = hbusreq1_p & d356ba | !hbusreq1_p & v845542;
assign df511b = hbusreq2_p & df511a | !hbusreq2_p & df552f;
assign v8cc47c = hlock0 & v8ccbd8 | !hlock0 & v8cc47b;
assign d35741 = hmaster1_p & d35740 | !hmaster1_p & d3570b;
assign c3ce25 = hgrant3_p & c3d5b0 | !hgrant3_p & c3ce24;
assign d35a1e = hbusreq2 & v84557a | !hbusreq2 & !v845542;
assign b1c740 = hbusreq3 & b1c73f | !hbusreq3 & !v845542;
assign c3cef4 = hgrant4_p & v845542 | !hgrant4_p & !c3ceee;
assign d354db = hmaster0_p & d354d9 | !hmaster0_p & !d354da;
assign df513d = hbusreq1 & df513c | !hbusreq1 & v845542;
assign c3d391 = hmaster1_p & c3d38e | !hmaster1_p & c3d390;
assign d35a11 = hmaster2_p & d35a0d | !hmaster2_p & d35a10;
assign v9ea5bb = hgrant3_p & v9ea57f | !hgrant3_p & v9ea5ba;
assign v8cc0e6 = hlock2 & v8cc4ad | !hlock2 & v8cc0e4;
assign d354f6 = hbusreq3 & d354f4 | !hbusreq3 & !d354f5;
assign d359a7 = hbusreq4_p & d359a5 | !hbusreq4_p & d359a6;
assign b1c4c5 = hbusreq4_p & b1c495 | !hbusreq4_p & !v845542;
assign v8cc623 = hmaster0_p & v8cc61c | !hmaster0_p & v8cc621;
assign c3d2ce = hmaster0_p & c3d2c8 | !hmaster0_p & c3d2cd;
assign b1c7ed = hgrant2_p & b1c7ec | !hgrant2_p & b1c7e4;
assign c3d699 = hmaster2_p & c3d669 | !hmaster2_p & !c3d675;
assign bd591c = hlock2_p & bd591b | !hlock2_p & !v845542;
assign v9f77c6 = stateG10_4_p & v9f77c4 | !stateG10_4_p & v9f77c5;
assign b57a8e = hready_p & b5799c | !hready_p & b57a8d;
assign v9f7d61 = hbusreq0_p & v9ea3fb | !hbusreq0_p & v9f7d5d;
assign d354f4 = hbusreq1_p & d354bd | !hbusreq1_p & d354f3;
assign v9f768a = hmaster1_p & v9f7689 | !hmaster1_p & v9f7d64;
assign c3d66d = hmastlock_p & c3d66b | !hmastlock_p & v84557a;
assign bd58cc = hbusreq0 & bd58c2 | !hbusreq0 & bd58cb;
assign ad5018 = hready & ad5017 | !hready & !v845564;
assign ad4fcf = hmaster2_p & v84556c | !hmaster2_p & !ad4fce;
assign c3d583 = hmaster1_p & c3d581 | !hmaster1_p & c3d582;
assign v9f7d7b = hgrant4_p & v9f7c9f | !hgrant4_p & !v9f7d79;
assign ad469b = hbusreq4_p & ad469a | !hbusreq4_p & v845542;
assign ad4e8a = hbusreq4_p & ad4e89 | !hbusreq4_p & b1cfb6;
assign ad4dbf = hmaster1_p & ad4dbe | !hmaster1_p & ad4db9;
assign c3d6c8 = hgrant0_p & c3d681 | !hgrant0_p & c3d66d;
assign bd583c = hgrant4_p & c3d674 | !hgrant4_p & !bd574e;
assign c73a9a = start_p & v845542 | !start_p & c76645;
assign ade5dc = hmaster1_p & ade5db | !hmaster1_p & ade5d9;
assign v9ea59b = hmaster2_p & v9ea4d2 | !hmaster2_p & v9ea59a;
assign v9ea618 = hready_p & v9ea436 | !hready_p & v9ea617;
assign d35a23 = hbusreq2 & d35a22 | !hbusreq2 & !v845542;
assign b8f6e1 = hgrant1_p & v845542 | !hgrant1_p & c3d2fd;
assign v9f784d = hlock2 & v9f784a | !hlock2 & v9f784c;
assign cc36c8 = stateG10_4_p & ade563 | !stateG10_4_p & dc500e;
assign v9e9ee6 = jx1_p & v9e9ed9 | !jx1_p & v9e9ee5;
assign cc36c1 = hmaster1_p & cc36bf | !hmaster1_p & cc36c0;
assign d6ebcc = hgrant3_p & d6ebc9 | !hgrant3_p & !d6ebcb;
assign v8cc035 = hgrant3_p & v8cc820 | !hgrant3_p & v8cc034;
assign c3d4f9 = hlock4_p & c3d319 | !hlock4_p & v845542;
assign ad4da8 = hlock4_p & v9f21c4 | !hlock4_p & v845542;
assign ad4711 = hgrant4_p & v845542 | !hgrant4_p & ad4fdc;
assign d359d8 = stateG10_4_p & v845542 | !stateG10_4_p & d359d6;
assign b059bd = hbusreq2 & b059bb | !hbusreq2 & b059bc;
assign bd58e9 = hmaster0_p & bd58e8 | !hmaster0_p & bd5773;
assign b1c761 = hmaster2_p & b1c755 | !hmaster2_p & !ade4df;
assign v9e9f6d = hlock4 & v9e9f68 | !hlock4 & v9e9f6c;
assign v9ea4c9 = hbusreq4_p & v9ea4c7 | !hbusreq4_p & v9ea4c8;
assign b1c722 = hbusreq0 & b1c721 | !hbusreq0 & v845542;
assign ade618 = hmaster0_p & ade5b4 | !hmaster0_p & ade569;
assign b57a1d = hbusreq1_p & b578fa | !hbusreq1_p & b57a1c;
assign adeaab = decide_p & adea8d | !decide_p & adeaa7;
assign b57a2b = hmaster1_p & b57a28 | !hmaster1_p & b57a2a;
assign ad47fb = hmaster1_p & ad47fa | !hmaster1_p & ad471b;
assign b1c4ca = hbusreq4_p & b1c4a3 | !hbusreq4_p & !v845542;
assign b1c77c = hmaster0_p & b1c75d | !hmaster0_p & b1c77b;
assign ade58c = hbusreq0_p & ade58a | !hbusreq0_p & !ade58b;
assign bd56cc = hready_p & bd5ea9 | !hready_p & !bd56cb;
assign v8cc7b4 = hlock3 & v8ccbe8 | !hlock3 & v8cc7b2;
assign ad474d = hgrant1_p & ad460d | !hgrant1_p & ad474c;
assign d357fd = hbusreq0 & d357fc | !hbusreq0 & d357fa;
assign dc4fa5 = hbusreq3 & dc4fa4 | !hbusreq3 & v845542;
assign b1d006 = hmaster1_p & b1cfb8 | !hmaster1_p & b1d005;
assign ad40fc = hready_p & ad4828 | !hready_p & ad40fb;
assign dc4f7f = hmaster2_p & dc4f7d | !hmaster2_p & !ade4e8;
assign ad4f6f = hgrant4_p & v845542 | !hgrant4_p & !ad4f36;
assign b57431 = hbusreq2 & b5742f | !hbusreq2 & b57430;
assign ad45a7 = hmaster0_p & ad459d | !hmaster0_p & ad456f;
assign ad4e84 = hmaster2_p & ad4e83 | !hmaster2_p & v845542;
assign c5c8e6 = hmastlock_p & c5c8e5 | !hmastlock_p & !v845542;
assign v9f7692 = hmaster2_p & v9f7d59 | !hmaster2_p & !v9f7e31;
assign b57502 = hmaster1_p & b57501 | !hmaster1_p & v845542;
assign d3573c = hready_p & d35735 | !hready_p & !d3573b;
assign v9e9f97 = hlock1 & v9e9f8e | !hlock1 & v9e9f96;
assign c3d34e = hbusreq4 & c3d34b | !hbusreq4 & !c3d34d;
assign c3d57e = hbusreq4 & c3d57a | !hbusreq4 & !c3d57d;
assign dc4fc0 = hmaster0_p & dc4fb8 | !hmaster0_p & dc4fbf;
assign ad4f20 = hbusreq2 & ad4f1f | !hbusreq2 & !v845542;
assign v9f7e04 = hlock1_p & v9f7ccf | !hlock1_p & v9f7d19;
assign b1c066 = hlock0_p & b1c7bb | !hlock0_p & !d3580b;
assign ad4293 = hbusreq1_p & ad4292 | !hbusreq1_p & v845542;
assign b1c5dd = hbusreq2_p & b1c5dc | !hbusreq2_p & b1c82f;
assign d356d2 = hbusreq1 & d3590e | !hbusreq1 & v845542;
assign c3d5c3 = hready & c3d5c2 | !hready & c3d313;
assign ad4e78 = stateG10_4_p & ad4e75 | !stateG10_4_p & !ad4e77;
assign b1c727 = hbusreq0 & b1c726 | !hbusreq0 & v845542;
assign c3ce52 = hbusreq1_p & c3ce51 | !hbusreq1_p & c3d305;
assign b57ac7 = hgrant1_p & b57ac6 | !hgrant1_p & b578f9;
assign ad46c7 = hlock4_p & ad4eec | !hlock4_p & ad4f36;
assign v9f7e1f = hmaster2_p & v9f7e1b | !hmaster2_p & !v9f7e1e;
assign v9f7d00 = hlock3 & v9f7cf8 | !hlock3 & v9f7cff;
assign ad3cc5 = decide_p & ad4476 | !decide_p & ad3cc4;
assign v9f76b5 = hmaster0_p & v9f7e01 | !hmaster0_p & v9f7d34;
assign v9f7e19 = hgrant4_p & v9f7ca5 | !hgrant4_p & v9f7d81;
assign b1c822 = hmaster1_p & b1c80c | !hmaster1_p & b1c821;
assign ad505a = stateG10_4_p & v845542 | !stateG10_4_p & ad5059;
assign v9f7682 = hlock2 & v9f767f | !hlock2 & v9f7681;
assign b1cf29 = hlock0_p & v845566 | !hlock0_p & !v845542;
assign v9f7db1 = hlock4_p & v9f7daf | !hlock4_p & v9f7db0;
assign v8cc0d7 = hgrant4_p & v8cc0c3 | !hgrant4_p & v845542;
assign b57957 = hmaster0_p & b5794e | !hmaster0_p & b57956;
assign ad4758 = hbusreq3 & ad46b4 | !hbusreq3 & !v845547;
assign d35a4a = hmaster2_p & d35a47 | !hmaster2_p & d35a49;
assign adea8b = hmaster2_p & adea8a | !hmaster2_p & !v845542;
assign ad504d = stateG10_4_p & ad504b | !stateG10_4_p & ad504c;
assign bd5759 = hbusreq3 & bd5758 | !hbusreq3 & v84556c;
assign bd5859 = hbusreq1 & c3d68a | !hbusreq1 & !v845542;
assign d356e5 = hmaster0_p & d356e2 | !hmaster0_p & d356e4;
assign ad4385 = hready & ad437f | !hready & ad4384;
assign b57445 = hmaster1_p & b57444 | !hmaster1_p & v845542;
assign b059f6 = hmaster1_p & b059bd | !hmaster1_p & b059f5;
assign b578f2 = hmaster0_p & b578f1 | !hmaster0_p & v845542;
assign ad4263 = jx0_p & ad48cb | !jx0_p & ad4262;
assign ad459d = hready & ad459a | !hready & ad459c;
assign v9f7e24 = hready & v9f7e23 | !hready & v9f7e1f;
assign ad40ec = hmaster0_p & ad40eb | !hmaster0_p & ad484c;
assign v9f7d1c = hlock3 & v9f7d1b | !hlock3 & v9f7d1a;
assign ad4f13 = hready & ad4ef2 | !hready & ad4f12;
assign c3cf31 = hgrant3_p & c3cf2c | !hgrant3_p & c3cf30;
assign d357f5 = hmaster2_p & d357f4 | !hmaster2_p & v84554a;
assign ad43ef = hlock4_p & ad43c6 | !hlock4_p & v845542;
assign b05a36 = hbusreq2_p & b05a33 | !hbusreq2_p & b05a35;
assign df54ff = decide_p & df54fd | !decide_p & d6ebca;
assign v9e9eab = hlock2 & v9e9ea8 | !hlock2 & v9e9eaa;
assign v9f776d = hmaster0_p & v9f7767 | !hmaster0_p & v9f776c;
assign b1c5fe = hready_p & b1c82d | !hready_p & b1c5fd;
assign ade660 = hready_p & ade65e | !hready_p & ade65f;
assign v9f7da5 = hbusreq0 & v9f7cf6 | !hbusreq0 & v9f7da4;
assign b57415 = hlock2 & b57983 | !hlock2 & b57414;
assign v9ea58e = hbusreq1 & v9ea58d | !hbusreq1 & v9ea586;
assign b05a47 = hmaster1_p & b05a46 | !hmaster1_p & b05943;
assign v9e9fca = decide_p & v9ea4b2 | !decide_p & v9e9fc9;
assign ade4f3 = hready_p & ade4b5 | !hready_p & ade4f2;
assign v9f7870 = hbusreq2 & v9f786e | !hbusreq2 & v9f786f;
assign ad4f31 = hgrant2_p & ad4f28 | !hgrant2_p & !ad4f30;
assign ad4467 = hready & ad445a | !hready & ad4466;
assign d354fb = hmaster0_p & d354f6 | !hmaster0_p & d354fa;
assign b57ad0 = hmaster0_p & b57acf | !hmaster0_p & b578fa;
assign v9ea449 = hmaster2_p & v9ea444 | !hmaster2_p & v9ea448;
assign c3ce62 = hbusreq1 & c3d2d9 | !hbusreq1 & v845542;
assign v9ea454 = hlock1 & v9ea3fa | !hlock1 & v9ea453;
assign v9f789a = hmaster1_p & v9f7892 | !hmaster1_p & v9f7899;
assign b05a0a = hgrant4_p & v9ea463 | !hgrant4_p & v9ea464;
assign v9f78a5 = hmaster0_p & v9f784e | !hmaster0_p & v9f7829;
assign df51b7 = hbusreq2_p & df51b4 | !hbusreq2_p & df51b6;
assign c3d6a0 = decide_p & c3d695 | !decide_p & c3d69f;
assign ad4f8a = hgrant4_p & v845542 | !hgrant4_p & !ad4f88;
assign v9f7dc0 = hbusreq1_p & v9f7d90 | !hbusreq1_p & v9f7db4;
assign ad4e68 = hburst0_p & c74202 | !hburst0_p & c74198;
assign b57903 = hmaster0_p & b578f9 | !hmaster0_p & b578fa;
assign ad3cda = hbusreq3 & ad3cd0 | !hbusreq3 & ad3cd9;
assign b57a83 = hgrant2_p & b579b0 | !hgrant2_p & b57a82;
assign b05a8b = hgrant2_p & b05a89 | !hgrant2_p & b05a8a;
assign c3d5bf = hgrant4_p & v845542 | !hgrant4_p & c3d5b7;
assign ad4405 = hmaster1_p & ad4404 | !hmaster1_p & ad43fc;
assign c5c8fe = hgrant4_p & v845542 | !hgrant4_p & !c5c8fd;
assign ade656 = hmaster1_p & v845542 | !hmaster1_p & ade655;
assign v9ea420 = hbusreq0_p & v9ea41e | !hbusreq0_p & v9ea41f;
assign v9f7861 = hlock4 & v9f785e | !hlock4 & v9f7860;
assign ad3d23 = hmaster1_p & ad3d22 | !hmaster1_p & ad43ba;
assign ad4460 = hlock0_p & adea99 | !hlock0_p & ad4387;
assign df51c1 = hmaster0_p & df51c0 | !hmaster0_p & df518f;
assign d3550e = hmaster0_p & d3542e | !hmaster0_p & d3550d;
assign b1c5e1 = hmaster0_p & b1cfb8 | !hmaster0_p & b1c5e0;
assign b05a40 = hmaster2_p & b05a3f | !hmaster2_p & !v9f7d42;
assign ad471a = hgrant1_p & ad45a4 | !hgrant1_p & ad4719;
assign ade587 = hburst1 & c3d66b | !hburst1 & v845542;
assign v9f7727 = hmaster0_p & d35aaa | !hmaster0_p & v9f7726;
assign d3559a = hbusreq0 & d35526 | !hbusreq0 & d35599;
assign ad4f39 = locked_p & ad4f38 | !locked_p & !v845542;
assign b1c5f1 = hgrant2_p & v845542 | !hgrant2_p & b1c5f0;
assign ad45ed = hbusreq4_p & ad45ec | !hbusreq4_p & v845542;
assign c3d4e1 = hbusreq4_p & c3d4e0 | !hbusreq4_p & !adeaa4;
assign b05923 = hbusreq4_p & b05922 | !hbusreq4_p & !v9f7d42;
assign jx0 = v9f78b1;
assign ad3cec = hgrant4_p & b1c714 | !hgrant4_p & ad3ceb;
assign ad4106 = hbusreq2 & ad4105 | !hbusreq2 & v845542;
assign b1c096 = decide_p & b1c095 | !decide_p & b1d013;
assign d35618 = hmaster2_p & dc5318 | !hmaster2_p & d35617;
assign v8cc801 = hlock1 & v8cc439 | !hlock1 & v8cc800;
assign d35a5b = hbusreq4_p & d35a5a | !hbusreq4_p & dc5010;
assign dc53a2 = hmaster1_p & dc53a1 | !hmaster1_p & v845542;
assign v9ea441 = hgrant0_p & v9ea3e6 | !hgrant0_p & v9f20a1;
assign ad4354 = hmaster0_p & ad4320 | !hmaster0_p & df5142;
assign b1cf3f = hmaster2_p & v845542 | !hmaster2_p & b1cf3e;
assign bd5826 = hbusreq1 & bd5749 | !hbusreq1 & dc4fcb;
assign ad41a6 = hbusreq2 & ad5064 | !hbusreq2 & v845542;
assign b1c090 = hready_p & b1c08e | !hready_p & !b1c08f;
assign ad41b3 = decide_p & ad481f | !decide_p & ad41b2;
assign c3ce8e = hmaster0_p & c3ce8c | !hmaster0_p & c3ce8d;
assign v9f7d5b = hmaster2_p & v9f7d59 | !hmaster2_p & !v9ea3fb;
assign v9e9fb2 = hbusreq2_p & v9e9fa1 | !hbusreq2_p & v9e9fb1;
assign v9f773f = hlock3_p & v9f773a | !hlock3_p & v9f773e;
assign dc52fb = hbusreq4_p & dc52fa | !hbusreq4_p & v84556c;
assign c3d304 = hbusreq0 & v845576 | !hbusreq0 & v845542;
assign ad3cbd = hgrant2_p & ad4478 | !hgrant2_p & ad3cbc;
assign bd5813 = hbusreq0 & bd5803 | !hbusreq0 & bd5812;
assign bd5754 = hbusreq2 & bd5752 | !hbusreq2 & v845542;
assign v9ea3ee = hlock0_p & v9f20a1 | !hlock0_p & v9ea3ed;
assign bd574d = hmaster2_p & bd572e | !hmaster2_p & adec89;
assign v9f7856 = hmaster0_p & v9f7779 | !hmaster0_p & v9f774f;
assign df507c = hmaster1_p & v845542 | !hmaster1_p & df507b;
assign ade621 = decide_p & ade620 | !decide_p & adeaa7;
assign v9f777e = hmaster1_p & v9f777d | !hmaster1_p & v9f776d;
assign d35590 = hbusreq1_p & d354d1 | !hbusreq1_p & d3558f;
assign d35a1b = hmaster0_p & d359e4 | !hmaster0_p & d35a1a;
assign v9f7868 = hbusreq3 & v9f7865 | !hbusreq3 & v9f7867;
assign v9f7708 = hlock2 & v9f7705 | !hlock2 & v9f7707;
assign v9e9f5f = hgrant1_p & v9e9ee9 | !hgrant1_p & v9e9f57;
assign v9f7779 = hbusreq2 & v9f7777 | !hbusreq2 & v9f7778;
assign b1c7af = hgrant1_p & b1c794 | !hgrant1_p & b1c7ae;
assign c3ce0a = decide_p & c3ce02 | !decide_p & c3ce09;
assign v9f781f = hlock0 & v9f77c8 | !hlock0 & v9f781e;
assign ad443b = hbusreq4 & ad443a | !hbusreq4 & ad4430;
assign ad4438 = hbusreq4_p & ad4437 | !hbusreq4_p & adeaa4;
assign d354b8 = hgrant1_p & d354a2 | !hgrant1_p & d354b7;
assign d35597 = hbusreq1_p & d3542f | !hbusreq1_p & d35522;
assign ac1454 = hready_p & ac1453 | !hready_p & !v845542;
assign v9ea3f4 = hbusreq2_p & v9ea3f1 | !hbusreq2_p & v9ea3f3;
assign b058e7 = locked_p & b058e6 | !locked_p & v9f7d42;
assign ad4f21 = hbusreq2 & ad4ecf | !hbusreq2 & v845542;
assign ad4578 = hbusreq3 & ad4577 | !hbusreq3 & v845542;
assign v9f77ed = hbusreq0_p & v845542 | !hbusreq0_p & !v9f77ec;
assign bd5828 = hbusreq1_p & bd5826 | !hbusreq1_p & bd5827;
assign ad4edc = hgrant4_p & ad4ecd | !hgrant4_p & ad4eda;
assign dc52f9 = hburst0 & dc52f8 | !hburst0 & adea98;
assign v9ea4b3 = locked_p & v9f20a1 | !locked_p & v9ea3ec;
assign v9f7db6 = hbusreq0 & v9f7dac | !hbusreq0 & v9f7db5;
assign ade584 = hbusreq1 & ade583 | !hbusreq1 & v9041a4;
assign b57ab4 = hbusreq2 & b57ab2 | !hbusreq2 & b57ab3;
assign dc5311 = hmaster1_p & dc5307 | !hmaster1_p & v84556c;
assign bd5832 = hmaster0_p & bd5825 | !hmaster0_p & bd5831;
assign ad4419 = hmaster0_p & ad4414 | !hmaster0_p & ad4418;
assign d35584 = hgrant1_p & d35578 | !hgrant1_p & d35583;
assign d354b1 = hgrant0_p & v845542 | !hgrant0_p & d354af;
assign c3d51f = hgrant2_p & c3d36c | !hgrant2_p & c3d51e;
assign c3ce19 = hmaster1_p & c3ce16 | !hmaster1_p & c3ce18;
assign b57a6d = hbusreq1 & b57a6c | !hbusreq1 & b57942;
assign ad4595 = hmaster1_p & ad4594 | !hmaster1_p & ad4591;
assign v9e9e6f = hready_p & v9ea436 | !hready_p & v9e9e6e;
assign v9ea4ad = hlock0_p & v9f20a1 | !hlock0_p & v9ea4ac;
assign b1c7a2 = hmaster2_p & b1c79b | !hmaster2_p & b1c7a1;
assign c3d338 = stateG10_4_p & c3d336 | !stateG10_4_p & c3d337;
assign b1cff6 = hgrant4_p & v845542 | !hgrant4_p & !b1cff5;
assign c3ce3b = hbusreq1 & c3d2b2 | !hbusreq1 & !v845542;
assign ad3cca = hgrant4_p & b1c714 | !hgrant4_p & c3cec2;
assign ade5df = hready_p & ade5c8 | !hready_p & ade5de;
assign ad45bc = hlock4_p & ad4d9a | !hlock4_p & !v845542;
assign b1c794 = hbusreq1_p & b1c792 | !hbusreq1_p & b1c793;
assign ade628 = hgrant3_p & ade5df | !hgrant3_p & ade627;
assign c3d594 = hbusreq2 & c3d592 | !hbusreq2 & v845555;
assign v9ea4e0 = hmaster1_p & v9ea4cb | !hmaster1_p & v9ea4db;
assign v9f76ed = hbusreq0_p & v9f7d82 | !hbusreq0_p & v9f76ec;
assign v9f7ca7 = hmaster2_p & v9f7ca5 | !hmaster2_p & !v9f7ca6;
assign v9f766b = hbusreq4 & v9f7669 | !hbusreq4 & v9f766a;
assign b1c7c4 = hgrant4_p & v845542 | !hgrant4_p & b1c7bc;
assign c3d2f6 = hmaster2_p & c3d2f5 | !hmaster2_p & v845576;
assign dc4fea = stateG10_4_p & ade557 | !stateG10_4_p & dc4fe9;
assign v9f7dc7 = hbusreq1_p & v9f7dc6 | !hbusreq1_p & !v9f7d2a;
assign v9ea42a = hgrant2_p & v9ea429 | !hgrant2_p & v9ea426;
assign v9f78a9 = hgrant2_p & v9f78a4 | !hgrant2_p & v9f78a8;
assign v9f7e0c = hlock2 & v9f7e09 | !hlock2 & v9f7e0b;
assign v9f77dd = hlock1 & v9f77d8 | !hlock1 & v9f77dc;
assign v8cc812 = hmaster0_p & v845542 | !hmaster0_p & v8cc810;
assign ad43f0 = hbusreq4_p & ad43ef | !hbusreq4_p & v845542;
assign ad45e5 = hmaster2_p & v845542 | !hmaster2_p & ad45e4;
assign d356ff = hbusreq1 & d35a4a | !hbusreq1 & v845542;
assign ad3d2d = hmaster1_p & ad3d2c | !hmaster1_p & ad4419;
assign ade59d = hgrant4_p & v84556c | !hgrant4_p & !ade59c;
assign dc53db = hready_p & v845542 | !hready_p & dc53da;
assign v9e9fae = hbusreq2 & v9e9fac | !hbusreq2 & v9e9fad;
assign c3ce02 = hbusreq2_p & c3cdfd | !hbusreq2_p & c3ce01;
assign bd5e9f = hmaster2_p & adec93 | !hmaster2_p & bd5e9e;
assign ad44a6 = hbusreq4_p & ad44a3 | !hbusreq4_p & ad44a5;
assign c3ce92 = hbusreq2 & c3d2d6 | !hbusreq2 & c3d2d9;
assign ade552 = hgrant0_p & c3d66d | !hgrant0_p & ade550;
assign b05a54 = hgrant2_p & b05a53 | !hgrant2_p & b05a50;
assign ad46f2 = hmaster1_p & ad46f1 | !hmaster1_p & ad46ec;
assign v9ea5d8 = hmaster1_p & v9ea5d7 | !hmaster1_p & v9ea579;
assign b57405 = hbusreq3_p & b573fa | !hbusreq3_p & b57404;
assign v8cc6b3 = decide_p & v8cc4f4 | !decide_p & v8cc626;
assign b058a2 = stateA1_p & v845542 | !stateA1_p & b058a1;
assign v9e9f78 = hmaster2_p & v9e9f52 | !hmaster2_p & v9e9f77;
assign bd5b9c = hlock3_p & bd5b90 | !hlock3_p & bd5b9b;
assign ad45f4 = hready & ad45e1 | !hready & ad45f3;
assign ad4292 = hbusreq1 & ad4fb3 | !hbusreq1 & v845542;
assign d3552d = hbusreq2_p & d3551d | !hbusreq2_p & d3552c;
assign dc531b = hbusreq3 & dc5317 | !hbusreq3 & dc531a;
assign c3ce07 = hmaster1_p & c3ce05 | !hmaster1_p & c3ce06;
assign b5799c = decide_p & b57982 | !decide_p & b5798b;
assign b1caf8 = hbusreq0 & b1caf5 | !hbusreq0 & b1caf7;
assign b058ad = hlock4 & b058aa | !hlock4 & b058ac;
assign b05a4e = hmaster1_p & b05a4d | !hmaster1_p & b058e1;
assign v9f783a = hlock3 & v9f7839 | !hlock3 & v9f7837;
assign b57950 = hlock4_p & b5794f | !hlock4_p & v845542;
assign v9ea4a6 = hmastlock_p & v9ea4a5 | !hmastlock_p & v845542;
assign v9f7848 = hgrant2_p & v9f7819 | !hgrant2_p & v9f7847;
assign v8cc7a2 = hbusreq2 & v8cc7a0 | !hbusreq2 & v8cc7a1;
assign bd5899 = hmaster1_p & bd5832 | !hmaster1_p & bd5898;
assign v9f7d28 = hready & v9f7d27 | !hready & !v9f7d23;
assign v9f7d87 = stateG10_4_p & v9f7d83 | !stateG10_4_p & v9f7d85;
assign bd5787 = hmaster2_p & bd5786 | !hmaster2_p & ade4c5;
assign b0590b = hbusreq4 & b05909 | !hbusreq4 & b0590a;
assign b0593c = hmaster0_p & b0593a | !hmaster0_p & b0593b;
assign ad41ae = hgrant3_p & ad40fc | !hgrant3_p & ad41ad;
assign d35be3 = hbusreq4_p & d35be2 | !hbusreq4_p & v845542;
assign c5c968 = locked_p & c5c967 | !locked_p & c5c896;
assign cc36f6 = hbusreq1_p & d35a49 | !hbusreq1_p & cc36f5;
assign d359b6 = hburst0 & d359b5 | !hburst0 & v845542;
assign d354a6 = hbusreq4_p & d354a5 | !hbusreq4_p & v845542;
assign d35420 = hmaster2_p & d3541f | !hmaster2_p & d3541b;
assign bd5796 = hmaster2_p & bd5786 | !hmaster2_p & !v845566;
assign ad4f0e = hgrant4_p & v845542 | !hgrant4_p & ad4f00;
assign ade63c = hbusreq2_p & adea8d | !hbusreq2_p & adeab1;
assign v9f7648 = hbusreq1 & v9f7646 | !hbusreq1 & v9f7647;
assign c3d5b8 = hgrant4_p & v845542 | !hgrant4_p & !c3d5b7;
assign ad484d = hmaster0_p & ad484b | !hmaster0_p & ad484c;
assign c3d309 = stateG10_4_p & ade562 | !stateG10_4_p & !c3d308;
assign ac1481 = hready_p & ac1480 | !hready_p & !v845542;
assign v9ea3fc = hmaster2_p & v9ea3e6 | !hmaster2_p & v9ea3fb;
assign v9e9fdb = decide_p & v9e9fda | !decide_p & v9ea409;
assign b1d018 = hready_p & b1d014 | !hready_p & b1d017;
assign v9f7e16 = stateG10_4_p & v9f7d78 | !stateG10_4_p & v9f7e15;
assign d354ad = hmastlock_p & ade54b | !hmastlock_p & !v845542;
assign v9f7659 = hgrant4_p & v9f7cd8 | !hgrant4_p & v9f7658;
assign b059f2 = hbusreq3 & b059ef | !hbusreq3 & b059f1;
assign df54e1 = hburst0 & df54dd | !hburst0 & df54e0;
assign ade4c7 = hmaster2_p & ade4c0 | !hmaster2_p & ade4c6;
assign b579c8 = hbusreq2 & b579c6 | !hbusreq2 & b579c7;
assign v8cc809 = hmaster0_p & v8cc7ee | !hmaster0_p & v8cc808;
assign ad4380 = hlock0_p & v84556c | !hlock0_p & v845542;
assign ad4fda = hgrant0_p & ad4fca | !hgrant0_p & v845542;
assign bd57cd = hbusreq2 & bd57c4 | !hbusreq2 & !v845542;
assign df54e6 = hbusreq1 & dc53a3 | !hbusreq1 & v845564;
assign d3558f = hbusreq0 & d3558c | !hbusreq0 & d3558e;
assign bd58c5 = hgrant0_p & df513b | !hgrant0_p & v84556c;
assign v9e9f9e = hbusreq2 & v9e9f9c | !hbusreq2 & v9e9f9d;
assign c3ced5 = hgrant2_p & v845551 | !hgrant2_p & c3ced4;
assign v8cc484 = hbusreq1 & v8cc483 | !hbusreq1 & v8ccbd8;
assign ade559 = hbusreq4_p & ade558 | !hbusreq4_p & !v845542;
assign v9ea414 = locked_p & v9ea413 | !locked_p & v845542;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hbusreq2_p = 0;
  hlock2_p = 0;
  hbusreq3_p = 0;
  hlock3_p = 0;
  hbusreq4_p = 0;
  hlock4_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmaster1_p = 0;
  hmaster2_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  hgrant2_p = 0;
  hgrant3_p = 0;
  hgrant4_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  stateG10_2_p = 0;
  stateG10_3_p = 0;
  stateG10_4_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hbusreq2_p = hbusreq2;
  hlock2_p = hlock2;
  hbusreq3_p = hbusreq3;
  hlock3_p = hlock3;
  hbusreq4_p = hbusreq4;
  hlock4_p = hlock4;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmaster1_p = hmaster1;
  hmaster2_p = hmaster2;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  hgrant2_p = hgrant2;
  hgrant3_p = hgrant3;
  hgrant4_p = hgrant4;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  stateG10_2_p = stateG10_2;
  stateG10_3_p = stateG10_3;
  stateG10_4_p = stateG10_4;
  jx0_p = jx0;
  jx1_p = jx1;
  jx2_p = jx2;
    end
endmodule

