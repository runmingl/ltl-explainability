module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hbusreq2, hlock2, hbusreq3, hlock3, hbusreq4, hlock4, hbusreq5, hlock5, hbusreq6, hlock6, hburst0, hburst1, hmaster0, hmaster1, hmaster2, hmastlock, start, decide, locked, hgrant0, hgrant1, hgrant2, hgrant3, hgrant4, hgrant5, hgrant6, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, stateG10_2, stateG10_3, stateG10_4, stateG10_5, stateG10_6, jx0, jx1, jx2, jx3);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v84561b;
  wire v845649;
  wire v22f9cb4;
  wire v23fb564;
  wire v230bf69;
  wire v84565f;
  wire v191a86f;
  wire v84563f;
  wire v22ec1cb;
  wire v23fc331;
  wire v2310c2b;
  wire bd757c;
  wire v2309295;
  wire v23fba6b;
  wire v23fcf46;
  wire v191a879;
  wire v10dbf64;
  wire v23f646e;
  wire v22eeb03;
  wire v2306d29;
  wire v23f476a;
  wire v23fb136;
  wire v191a876;
  wire v23126ae;
  wire v106af73;
  wire v23f4426;
  wire v23fbf37;
  wire v22f2f3e;
  wire v22f7176;
  wire v1aad6c8;
  wire v23fc378;
  wire v23f5cb3;
  wire v22f56d2;
  wire v230f63f;
  wire v23070c1;
  wire v22fdfde;
  wire v23f5d1a;
  wire v2311d0c;
  wire v22f666d;
  wire v23f55ea;
  wire v23f606c;
  wire v23fae84;
  wire v23fbfb9;
  wire v2302e32;
  wire v22eb1f5;
  wire v22fa870;
  wire v1aaddf4;
  wire v22fbb99;
  wire v231170f;
  wire v23046f7;
  wire v22fd25c;
  wire v22fae6e;
  wire v230a24c;
  wire v230889a;
  wire v22f00b6;
  wire v22f7d5d;
  wire v22f0e00;
  wire v2306fba;
  wire v22ef05d;
  wire v23fc904;
  wire v22f5e8c;
  wire v230320e;
  wire v23fc127;
  wire v22f8be5;
  wire v23125a8;
  wire v22ee47d;
  wire v230e40c;
  wire bc87ee;
  wire v22fccf1;
  wire v23f4201;
  wire v2392d61;
  wire v23fb8bf;
  wire v22eb5b3;
  wire v23fce86;
  wire v23fcc36;
  wire v23fbca3;
  wire v23fcf5b;
  wire b3d617;
  wire v23fbfaa;
  wire v22f18a3;
  wire v23f5474;
  wire v23fba4a;
  wire v23f724e;
  wire v23fcb29;
  wire v22f243b;
  wire v22f0e99;
  wire v230f133;
  wire v22ecb12;
  wire v22f4ef7;
  wire v23045dc;
  wire v22f5272;
  wire v230c4c3;
  wire v22eec47;
  wire v23f6ad0;
  wire v2304904;
  wire v22eec2a;
  wire v23fbe50;
  wire v23094c7;
  wire v23fcf62;
  wire v23fc541;
  wire v230e75b;
  wire v23fc3da;
  wire v23f95bd;
  wire v23fc29b;
  wire v22f7aff;
  wire v23fc757;
  wire v23fc3e8;
  wire v23f3d47;
  wire v230741d;
  wire v23fb8aa;
  wire v22f7dbc;
  wire v2305aa9;
  wire v22f46ff;
  wire v22f5808;
  wire v23fc7a7;
  wire v22f0a24;
  wire d49f2b;
  wire v2308b58;
  wire v23041ea;
  wire v230ca0f;
  wire v23fc963;
  wire v22ec354;
  wire v2309475;
  wire v23fb7c3;
  wire v23fc3aa;
  wire v22f7ec9;
  wire v23f39e6;
  wire v22f8a46;
  wire v2304082;
  wire v23117c1;
  wire v23fcc3d;
  wire v23fc372;
  wire b1e9fa;
  wire v22f0bb6;
  wire v230ccaf;
  wire v22f151d;
  wire v23f5429;
  wire v2392811;
  wire v22f5c1b;
  wire v23f38b7;
  wire v22fd364;
  wire v22eb02e;
  wire v23fb82a;
  wire v23fbe9d;
  wire v22f1744;
  wire v23fb143;
  wire v22fcdd3;
  wire v23f6c83;
  wire v23fc7c7;
  wire v2304a06;
  wire v23f74b7;
  wire v23fc4e2;
  wire v23fbf06;
  wire v230b77e;
  wire fc8c53;
  wire v22f639d;
  wire v23f42ec;
  wire v22f446b;
  wire v23fb533;
  wire v22fdf28;
  wire v23f52f2;
  wire v23fc0d4;
  wire v23113f5;
  wire v230a6c8;
  wire v2303d9e;
  wire v2392394;
  wire v22eb2ee;
  wire v2311031;
  wire v22ff29f;
  wire v23fc7d9;
  wire v2300995;
  wire v22fcabb;
  wire v23fc86a;
  wire v23067c9;
  wire v23f7c5a;
  wire v230418f;
  wire v2303554;
  wire v23fce1b;
  wire v230ad74;
  wire v23fc1ec;
  wire v23fbba0;
  wire v22f580c;
  wire v23fcae1;
  wire v230b93b;
  wire v23fc087;
  wire v2305141;
  wire v23fc7f2;
  wire v23fcd9b;
  wire v231228f;
  wire v230754e;
  wire v23123a3;
  wire v22f8639;
  wire v191ac63;
  wire v23fbe02;
  wire v2311b9e;
  wire v22f68f1;
  wire v23069b0;
  wire v23022d5;
  wire v1aae8d3;
  wire bd74e7;
  wire v23fcb75;
  wire v22f16bf;
  wire v22f334c;
  wire v1e8439a;
  wire v22f9396;
  wire v22f01b6;
  wire v23fc02a;
  wire v23fc26a;
  wire v23f6d65;
  wire v22eeab9;
  wire v22f2592;
  wire v22f45d7;
  wire v230dfa0;
  wire v2308d60;
  wire v23f5d39;
  wire v22ff21b;
  wire v23fc20d;
  wire v2394087;
  wire v22fa5f1;
  wire v1aad4c6;
  wire v23fc92f;
  wire v92eb35;
  wire v23f38f8;
  wire v23f3bde;
  wire v23013b5;
  wire v230200a;
  wire v2300362;
  wire v23f5066;
  wire v23fc01f;
  wire v23fce88;
  wire v23025e4;
  wire v23fb0f0;
  wire v23fcb6d;
  wire v23f259c;
  wire v22ed34b;
  wire v22f9d07;
  wire v230e932;
  wire v23130d6;
  wire v230d664;
  wire v23f3501;
  wire v22efe81;
  wire v22f91ef;
  wire v22f7fdd;
  wire v230170e;
  wire v22f8686;
  wire v22fa6f5;
  wire v2309d23;
  wire v23068f2;
  wire v2312ebb;
  wire v22eaf83;
  wire v23070ef;
  wire v23fcfb1;
  wire v22f8c01;
  wire v22f9cd9;
  wire v2302e7b;
  wire v23fc061;
  wire v22ff0de;
  wire bd8ac4;
  wire v23faade;
  wire v23f420c;
  wire v230f549;
  wire v22f0635;
  wire v22f32df;
  wire v23f7cec;
  wire v23132db;
  wire v23fb670;
  wire v22edc69;
  wire v231138f;
  wire c26df3;
  wire v8958ff;
  wire v23fb8b8;
  wire v23fbf7f;
  wire v23fcbaf;
  wire v23f6032;
  wire v23f8e1c;
  wire v230236f;
  wire e1c7f2;
  wire v2311ed2;
  wire v23f5dfd;
  wire v22ec2c0;
  wire v22fbb46;
  wire v23f7b9b;
  wire v23934ed;
  wire v230ccc4;
  wire v22fd907;
  wire v22f939d;
  wire v23f3d5b;
  wire v23fc324;
  wire v22efef6;
  wire v94e4a6;
  wire v22f021c;
  wire v23fc9c6;
  wire v22fb4e3;
  wire v22f7f74;
  wire v22fef4f;
  wire v22ec29a;
  wire v2307582;
  wire v22f7cab;
  wire v2307a0f;
  wire v22f1a02;
  wire v23127ef;
  wire v2312283;
  wire v22fe9b7;
  wire v22f3502;
  wire v13afa38;
  wire v22f0e5e;
  wire v22f08d0;
  wire v23f4855;
  wire v2303068;
  wire v22fcbcd;
  wire v23fcbb5;
  wire v106af4d;
  wire v23fbe4c;
  wire v22ec0d4;
  wire v22ff463;
  wire v23fba24;
  wire v23f8928;
  wire bd766b;
  wire v23fd033;
  wire v22f66bc;
  wire v23fb410;
  wire v2303d1d;
  wire v23fcccf;
  wire v23fc004;
  wire v230d4f1;
  wire v2312a23;
  wire v23fcd8e;
  wire v23f2553;
  wire v23fcd29;
  wire v23f94bc;
  wire v23f6865;
  wire v230a51c;
  wire v22f2b52;
  wire v23f0cbe;
  wire v22f8aea;
  wire v22f6dfa;
  wire v22fba0e;
  wire v22f5e59;
  wire v22efc2a;
  wire v2309377;
  wire v23fb849;
  wire v22fdbf7;
  wire v191b1f3;
  wire v22f42c9;
  wire v2300c5c;
  wire v23fc914;
  wire v2310c7c;
  wire v22ee34a;
  wire v230f050;
  wire v15072af;
  wire v938878;
  wire v22ee0db;
  wire v23f425f;
  wire v22f09ab;
  wire v230178e;
  wire v22fbb33;
  wire v230fd1d;
  wire v22f33c4;
  wire v22fcdf7;
  wire v1aae387;
  wire v22f8fb2;
  wire v230cfe2;
  wire v22f2958;
  wire v23f707f;
  wire v22ff64f;
  wire v23085df;
  wire v230ff13;
  wire v22f9c73;
  wire v23fb61f;
  wire v23fc9f1;
  wire v23fb4b6;
  wire v230f5e2;
  wire v230f222;
  wire v23fc7a4;
  wire v230e7e3;
  wire v22f08be;
  wire v230df19;
  wire v230a2b1;
  wire v23f069d;
  wire v2306ee6;
  wire v23fcb36;
  wire v23fc5a0;
  wire v22fc85f;
  wire v230521a;
  wire v23f0b4e;
  wire v23fcd84;
  wire v22fd2ec;
  wire v22faefb;
  wire v230219b;
  wire v23fa75a;
  wire v2312d11;
  wire v23048df;
  wire v23f1d8b;
  wire v23f0a0b;
  wire v23fc225;
  wire v23f5fcd;
  wire v191b04d;
  wire v23fb992;
  wire b9d0d2;
  wire v2303558;
  wire v23fbf10;
  wire v2308b4b;
  wire v2307852;
  wire v23fc821;
  wire v23fc802;
  wire v2305a69;
  wire a1fd46;
  wire v2312e03;
  wire v22f215c;
  wire v22ff6e8;
  wire v23fc7fb;
  wire v1aad586;
  wire v22ff404;
  wire v23fc782;
  wire v2312de4;
  wire v23fc94c;
  wire v2300338;
  wire v23003b8;
  wire v2308356;
  wire v2300bb2;
  wire v230d5be;
  wire v22f249f;
  wire v23060ed;
  wire v23f1109;
  wire v23fc2f1;
  wire v23035c1;
  wire v23fcd4f;
  wire b00a61;
  wire v23fba3f;
  wire v22f45ac;
  wire v2309bda;
  wire v23fb18e;
  wire v23f57c1;
  wire v2303061;
  wire v22f854f;
  wire v23f9d0b;
  wire v230a744;
  wire v22f9df1;
  wire v9bf2ce;
  wire v23fcbab;
  wire v23f75e9;
  wire v2304fae;
  wire v23fcb3c;
  wire v23f79b4;
  wire v22f067f;
  wire v22f6385;
  wire v22f220a;
  wire v22ec477;
  wire v23fc74f;
  wire v231343f;
  wire v23129e0;
  wire v23fcff6;
  wire v22ff9c3;
  wire v23fc2b7;
  wire v23fbd7e;
  wire v1aad421;
  wire v2300437;
  wire v22f18b4;
  wire v23fc2ba;
  wire v22efc42;
  wire v230db4e;
  wire v230160e;
  wire v23fcf74;
  wire v230aba5;
  wire v23fcd9f;
  wire v2301797;
  wire v23fbb73;
  wire v23f53e9;
  wire v23fc247;
  wire v22fb260;
  wire v23033d3;
  wire v22fee58;
  wire v191b18a;
  wire v22eeb42;
  wire v23f47ca;
  wire v22ed741;
  wire v23fcf89;
  wire v23f7a18;
  wire v86df86;
  wire v230788d;
  wire v22fda8c;
  wire v22f83d7;
  wire v239253c;
  wire v23fbe00;
  wire v22f6e29;
  wire v23f6d9c;
  wire v22f2a94;
  wire v22fd196;
  wire v23fcfb6;
  wire v23f9885;
  wire v23f4ff3;
  wire v230b7c8;
  wire v23fc550;
  wire v1aada8c;
  wire v23120a5;
  wire v22f1d46;
  wire v2308fc5;
  wire v22f94ba;
  wire v23041b6;
  wire v23fb8da;
  wire v22f39e3;
  wire v23000e2;
  wire v22fac2f;
  wire v22eee34;
  wire v22f4a4f;
  wire v2300fb4;
  wire v22f78b7;
  wire v953acf;
  wire v23fcd74;
  wire v2392868;
  wire v23fb526;
  wire v230e539;
  wire v23fca3e;
  wire v23067ba;
  wire v22fb8df;
  wire v2392229;
  wire v239342f;
  wire v23fcf38;
  wire v23fbd0e;
  wire v23fc847;
  wire v2303707;
  wire v23f8679;
  wire c0e31a;
  wire v22eb498;
  wire v22f6d45;
  wire v22efe01;
  wire v23fc854;
  wire v2304fc6;
  wire v22f83fb;
  wire v22f865d;
  wire v22ee75e;
  wire v23fc349;
  wire v22ff0ef;
  wire v23f83af;
  wire v2300b33;
  wire v861565;
  wire v23107cf;
  wire v230627c;
  wire v23fc430;
  wire v23fcf7a;
  wire v22eef92;
  wire v22ebe46;
  wire v230538c;
  wire v22eb9b4;
  wire v23fb4e5;
  wire v2312e39;
  wire ba1576;
  wire v230a0d1;
  wire v23f8efa;
  wire v23f7e3d;
  wire v23f9b49;
  wire bd74f4;
  wire v22f5125;
  wire v2311831;
  wire v23019f7;
  wire v2301463;
  wire v22ed5c5;
  wire v22fe2b6;
  wire v22ebe13;
  wire v22ee9bb;
  wire v230290f;
  wire v22fe4ea;
  wire v22f6228;
  wire v22ec934;
  wire v23007c9;
  wire v230ef73;
  wire v2312cf9;
  wire v22f8eb8;
  wire v23f8a89;
  wire v23fbfb6;
  wire v23f8fc1;
  wire v2310222;
  wire v191ab52;
  wire v22ee09a;
  wire v230913e;
  wire v23f18a1;
  wire v23fc473;
  wire v23f2bb6;
  wire v22fc6b9;
  wire v23fbf8e;
  wire v22fde04;
  wire v23f5dd2;
  wire v23fcebe;
  wire v23f4015;
  wire v23f9dba;
  wire v22f14d1;
  wire v2306bfb;
  wire v22fee9e;
  wire v23fbd71;
  wire v1aad4b7;
  wire v23fc42e;
  wire v23fc679;
  wire v23fceb5;
  wire v230183d;
  wire v22f81a7;
  wire v2311f44;
  wire v2302b93;
  wire v23068bb;
  wire v2310f12;
  wire b42c55;
  wire v22f10a7;
  wire v230a407;
  wire v23f55a4;
  wire v23f710c;
  wire v230b6fc;
  wire v22eb83a;
  wire v23f4fa9;
  wire v23fc618;
  wire v23fca40;
  wire v23f9193;
  wire v23fc2ff;
  wire v22eddfd;
  wire v873a56;
  wire v22f8917;
  wire v23fc7dd;
  wire v230ad5b;
  wire v23fad76;
  wire v23fb121;
  wire v23fb1d4;
  wire v22fa662;
  wire v22fe582;
  wire v23fb848;
  wire v22f4ef1;
  wire v23fadf4;
  wire v23f572e;
  wire v2305a05;
  wire v2307b9c;
  wire v23f9db0;
  wire v22f51ba;
  wire v22fd32a;
  wire v22ed725;
  wire v230e94e;
  wire v2393ecb;
  wire d49f32;
  wire v230717d;
  wire v935301;
  wire v1506fdd;
  wire v2308c4d;
  wire v191aa68;
  wire v22f2bab;
  wire v2303c9d;
  wire v23fc026;
  wire v23fc19b;
  wire v22f580d;
  wire v22fba38;
  wire v23fc151;
  wire v22ecc15;
  wire v2392d6d;
  wire v22fa5a5;
  wire v23f6cdb;
  wire v22fd559;
  wire v23fc347;
  wire v231253d;
  wire v22ec414;
  wire v239387a;
  wire v23f1688;
  wire v230eb13;
  wire v23fcb38;
  wire v23fc393;
  wire v23f6a8a;
  wire v2300032;
  wire a1fe27;
  wire v22fe62b;
  wire v2302a4d;
  wire v23117f5;
  wire v22fd6fb;
  wire v230833e;
  wire v23f9307;
  wire v23fb604;
  wire v23f8866;
  wire v230695e;
  wire v22ef983;
  wire v22fcd0f;
  wire v22f6a6e;
  wire v2308d09;
  wire v22eb840;
  wire v22f9d92;
  wire v23f3a16;
  wire v2309871;
  wire v23fb029;
  wire v22f7022;
  wire v22f7c2b;
  wire v2302c67;
  wire v22eaaa7;
  wire v22ef144;
  wire v22fd799;
  wire v22f57ea;
  wire v23fa3bb;
  wire v23fcc5e;
  wire v230dc43;
  wire v23fc8ba;
  wire v23f8d79;
  wire v22f56a5;
  wire v23f0eec;
  wire v23f1225;
  wire v22faa26;
  wire v23f8a49;
  wire v2311af8;
  wire v2312e4e;
  wire v2306088;
  wire v2304aae;
  wire v23fb701;
  wire v230a934;
  wire v23fcd24;
  wire v23008f3;
  wire v22f9b67;
  wire v22f68e5;
  wire v23fc152;
  wire v23f8d9f;
  wire v23fcd2a;
  wire v23122fa;
  wire v23f36a3;
  wire v230de82;
  wire v22ebedc;
  wire v23f4758;
  wire v23f5907;
  wire v23f58bb;
  wire v22f1895;
  wire v22fda61;
  wire v1e840b4;
  wire a9c602;
  wire v23efa84;
  wire v230fc64;
  wire v22fbbd0;
  wire v230f7ce;
  wire v230b8fe;
  wire v23f2837;
  wire v23f273b;
  wire v22fca64;
  wire v23fba12;
  wire v22ed6e1;
  wire v2305c54;
  wire v2312d03;
  wire v23fc7f4;
  wire v23fc776;
  wire v23f52f3;
  wire v23f6db4;
  wire v22f6759;
  wire v2307dfb;
  wire v23928ae;
  wire b59af9;
  wire v23fbc1b;
  wire v23fc4df;
  wire v23fc885;
  wire v22eba40;
  wire v2305933;
  wire v23f437e;
  wire v23fbe99;
  wire v22f65dd;
  wire v23fbf84;
  wire v230723b;
  wire v22fcea3;
  wire v23fc9d6;
  wire v23fc613;
  wire v23fcd97;
  wire v231324d;
  wire v22f0074;
  wire v22f9980;
  wire v22f5d84;
  wire v917514;
  wire v9eaa59;
  wire v22eef3f;
  wire v22fc2c1;
  wire v2309561;
  wire v23105ac;
  wire v23fc9be;
  wire v23f6f14;
  wire v23fc0ac;
  wire v22f1d1a;
  wire v22ec855;
  wire v23066bf;
  wire v23067c3;
  wire v97b313;
  wire v22eb397;
  wire v22fa440;
  wire v230bd96;
  wire v23fc484;
  wire v23f3915;
  wire v230d24a;
  wire v22f35e8;
  wire v23fc65d;
  wire v23fc7bb;
  wire v2312f4f;
  wire v230c3aa;
  wire v230f257;
  wire v230c83a;
  wire v2305eb1;
  wire v1e8408c;
  wire v22f257b;
  wire v22f8f5c;
  wire v23f443d;
  wire v22f4986;
  wire v23f2d31;
  wire v23fbcc8;
  wire v22f8f1e;
  wire v23fc282;
  wire v23041e2;
  wire v22fc5d2;
  wire v22f37e8;
  wire v230b3d5;
  wire v2309840;
  wire v22ef499;
  wire c20a75;
  wire v1e84b3d;
  wire v23f7bc9;
  wire v23f8529;
  wire v23094b2;
  wire v230bb08;
  wire v22fb062;
  wire v23fce06;
  wire v22ee3ca;
  wire v23fbc43;
  wire v23f3f24;
  wire v22eaaba;
  wire v22fde5c;
  wire v22eaf66;
  wire v22eafde;
  wire v2310969;
  wire v23fc267;
  wire v22f324a;
  wire v230ca62;
  wire v231045a;
  wire v23fcc1c;
  wire a9176f;
  wire v23fc162;
  wire v23faede;
  wire v23fcec8;
  wire v23f3c00;
  wire v22f0ea8;
  wire v22f771b;
  wire v22f9f2f;
  wire v23f2eff;
  wire v2310b15;
  wire aacd54;
  wire v230b3d2;
  wire v2302e0f;
  wire v23007de;
  wire v23fc0e7;
  wire v2393401;
  wire v22eef1f;
  wire v2312ebe;
  wire v22ff1cb;
  wire v2312b57;
  wire v23037f2;
  wire v2300474;
  wire v22ffc69;
  wire v91b2de;
  wire v22f8483;
  wire v2303f04;
  wire v22ef823;
  wire v23fca2d;
  wire v22f7d4e;
  wire v23fc851;
  wire v23034a4;
  wire v22f346d;
  wire v8a6d1a;
  wire v230c6f1;
  wire v23031f0;
  wire v23fc00a;
  wire v1aae9a1;
  wire v22eb664;
  wire v23f60d2;
  wire v22fea3f;
  wire v23f5f4d;
  wire bd772c;
  wire v23fcb62;
  wire v230262f;
  wire v23fb6ce;
  wire v23fc461;
  wire v919672;
  wire v2313230;
  wire v23fc89d;
  wire v22ef9ff;
  wire v2308e64;
  wire v23fc36b;
  wire v22ef962;
  wire v23fcab4;
  wire v23113f1;
  wire v22fbbd2;
  wire v230fe41;
  wire v23fb842;
  wire v230b516;
  wire v23f6d93;
  wire v230d2a8;
  wire v2310e40;
  wire v2302460;
  wire v2300dcb;
  wire v239158d;
  wire v1aae2e4;
  wire v23fb661;
  wire v230abb0;
  wire v1aad535;
  wire v2308a2f;
  wire v23fc740;
  wire v23fcaae;
  wire bd7b44;
  wire v23f5dfe;
  wire v22f758c;
  wire v23fb886;
  wire v23fc5ac;
  wire v23fc4d8;
  wire v230446b;
  wire v23f8294;
  wire v23099b2;
  wire v23fd018;
  wire v23f5df1;
  wire v23f84dc;
  wire v23f2af5;
  wire v23f5388;
  wire v22f70bf;
  wire v22fb631;
  wire v23f1221;
  wire v2307e41;
  wire v23fb8f7;
  wire v22fefde;
  wire v230749a;
  wire v1aae277;
  wire v2305b24;
  wire v23132e5;
  wire v23fc946;
  wire v22f1d1f;
  wire v2302e1b;
  wire v23f5893;
  wire v22ebbf2;
  wire v230ecb6;
  wire v23108bb;
  wire v2302a57;
  wire v2302b81;
  wire v22f0fcd;
  wire v23f9a3a;
  wire v22fc2d0;
  wire v230c94b;
  wire v22fa0b2;
  wire v22ec60b;
  wire v23f4f2c;
  wire v23fbb81;
  wire v23fa69e;
  wire v22fdc20;
  wire v22fb0cb;
  wire v22eb899;
  wire v2300d51;
  wire v22fbfe5;
  wire v23fb55a;
  wire v22ebe78;
  wire v230e2f9;
  wire v22f533e;
  wire f40dc0;
  wire v230b6a4;
  wire v23f7968;
  wire v22fd30c;
  wire v23fcf91;
  wire v23fcd3c;
  wire v2311dff;
  wire v230bd05;
  wire v22f954f;
  wire v2307701;
  wire v23f512e;
  wire v23fbc42;
  wire v22fc7c1;
  wire v23055b3;
  wire v22f6a6b;
  wire v22fb706;
  wire v23f4af5;
  wire v23071f6;
  wire bd7c3f;
  wire v23f9a56;
  wire v23f13f3;
  wire v2306d08;
  wire v2307ff5;
  wire v22ee750;
  wire v23fcccd;
  wire v22f9c42;
  wire v22f6cc8;
  wire v23fba79;
  wire v22f41ee;
  wire v23fc2a5;
  wire v23fcb9a;
  wire v230c2b1;
  wire v22fb773;
  wire v22feb8b;
  wire v22f2851;
  wire v22fafa5;
  wire v23037ac;
  wire v2308dbf;
  wire v23073e6;
  wire b159aa;
  wire v22ed49b;
  wire v2301709;
  wire v2304299;
  wire v230254a;
  wire v22ef3d4;
  wire v23108aa;
  wire v22fc9bf;
  wire f406c6;
  wire v22ffcb8;
  wire v23929d0;
  wire v230a644;
  wire v22ed9a9;
  wire v2311ec3;
  wire v22f5605;
  wire v23fc3a7;
  wire v23fc0ce;
  wire v23022f2;
  wire v23012e5;
  wire v23f520c;
  wire v2308592;
  wire v22f753d;
  wire v2313618;
  wire v12cda57;
  wire v23fc8ea;
  wire v23fb838;
  wire v22f61b1;
  wire v22ec20d;
  wire v22f04ac;
  wire v23f7aea;
  wire v23fcb3b;
  wire v22f4e9f;
  wire v231396f;
  wire v22ed4ea;
  wire v22f61d2;
  wire v23f56c0;
  wire v22fe260;
  wire v22eefc4;
  wire v23fa8d7;
  wire v23fba65;
  wire v23fbbb9;
  wire v22f13ad;
  wire v2303516;
  wire v2310e81;
  wire v23f6130;
  wire v22f6d58;
  wire v23fc362;
  wire v23fc750;
  wire v23fcbf3;
  wire v23fd051;
  wire v23fb720;
  wire v2311506;
  wire a5a279;
  wire a88394;
  wire v23f3ab0;
  wire v22ff9d9;
  wire v23f480d;
  wire v23f8036;
  wire v23fb9d0;
  wire b09263;
  wire v230e9d1;
  wire v23fbe7b;
  wire v2308b98;
  wire v22edb13;
  wire v22f79be;
  wire v230c727;
  wire v2391d99;
  wire v22fd150;
  wire v2312401;
  wire v23fb7b2;
  wire v22f2bc2;
  wire v22fa823;
  wire v22f0b45;
  wire v2391a62;
  wire v22eb6fc;
  wire v22ebedd;
  wire v22f2cb3;
  wire v2302693;
  wire adc67b;
  wire v23fc78e;
  wire v22f7879;
  wire v2304f67;
  wire v23f3bcb;
  wire v2313266;
  wire v2307646;
  wire v22f9049;
  wire v23f2a7c;
  wire v231007b;
  wire v23126b1;
  wire v2306e27;
  wire v23f2c8b;
  wire v23fb175;
  wire v23074aa;
  wire v23fc039;
  wire v22f4f06;
  wire v2301c2a;
  wire v12cd4be;
  wire v22fb49d;
  wire v23fbca1;
  wire v22f1b18;
  wire v23fbf02;
  wire v22f0a39;
  wire v23f8095;
  wire v2302608;
  wire v230c6c0;
  wire v22fd298;
  wire v23fb583;
  wire v22ed881;
  wire v2303acd;
  wire v23fc67b;
  wire v2304d08;
  wire v23fbbcb;
  wire v22fc32c;
  wire v23066e8;
  wire v22f9cee;
  wire v2391a45;
  wire v23fb7a3;
  wire v23fc4b7;
  wire v23f4edc;
  wire v23fce02;
  wire v230be28;
  wire v23f664b;
  wire v22f79a5;
  wire v22f3730;
  wire v23fcbfb;
  wire v23fbdd8;
  wire v2307170;
  wire v22ff30c;
  wire v23fb954;
  wire v22ec8dc;
  wire v106a7d3;
  wire v23fc90b;
  wire v22edb96;
  wire v22fec34;
  wire v22ff3c3;
  wire v22f04b5;
  wire v23f17ff;
  wire v22f04ff;
  wire v22ec960;
  wire fc8fcf;
  wire v23fcc89;
  wire v22fe84a;
  wire v22f7d00;
  wire v23f5deb;
  wire b6f226;
  wire v22f7f3f;
  wire v22f230d;
  wire v23fbe6c;
  wire v23fc45d;
  wire v239298e;
  wire a1fc4e;
  wire v22edaf2;
  wire v23fc1a7;
  wire v22fd136;
  wire v22f1aae;
  wire v23fc636;
  wire v22f1040;
  wire v23fce9c;
  wire v23fb188;
  wire v22f7524;
  wire v23fcb9c;
  wire v23fb5b9;
  wire v22f1969;
  wire v1507088;
  wire v23fbe51;
  wire e1dd6a;
  wire v23fc6f7;
  wire v1aad3ae;
  wire v23fced8;
  wire v23f1bbf;
  wire v23fc0ab;
  wire v23fad33;
  wire v2308f89;
  wire v230b68a;
  wire v23f56de;
  wire v23fbe6e;
  wire v23fb144;
  wire v230b5c7;
  wire v22f4284;
  wire v23f2c35;
  wire a1fcb8;
  wire v23f95ba;
  wire v22ecdc8;
  wire v22f6618;
  wire v22eb6e2;
  wire v23f5a6d;
  wire v22ff5c1;
  wire v230387b;
  wire v230f82f;
  wire v23f1c12;
  wire c20101;
  wire v23fcc42;
  wire v22ed711;
  wire v22eaf2a;
  wire v22f5c2b;
  wire v23f1a2b;
  wire v2301a7e;
  wire v2300048;
  wire v23fbdf6;
  wire v230af11;
  wire v23fc4d4;
  wire v23fb7c8;
  wire v22ef38d;
  wire v23fbced;
  wire v23044d2;
  wire v22fa0ec;
  wire v23fbdd2;
  wire v22f8c8d;
  wire v23f4117;
  wire v22fe76b;
  wire v23fa2b8;
  wire v22ebc26;
  wire v230bd1c;
  wire v23f44e8;
  wire v22fdc30;
  wire v23fbd56;
  wire v22f81ba;
  wire v2306e0e;
  wire v23fb094;
  wire v15074d0;
  wire v22f5db6;
  wire v23fbfc0;
  wire v22f789c;
  wire v22ecc3f;
  wire v23fccbe;
  wire v2302251;
  wire v23f1e5c;
  wire v23f6fa8;
  wire v23fb43a;
  wire v22f1d85;
  wire v230fbb3;
  wire v2307ab6;
  wire bfba4f;
  wire v230935d;
  wire v23f3e38;
  wire v22f6629;
  wire v9b93b3;
  wire v8b4671;
  wire v23f6c7c;
  wire v23f9fcf;
  wire v22ec39f;
  wire v23fb5f1;
  wire v22f86f3;
  wire af7272;
  wire v22fe426;
  wire v22efc9e;
  wire v23fc063;
  wire fc8fe6;
  wire v22fb4d8;
  wire v2391e8e;
  wire v22ee0c9;
  wire v230997a;
  wire v23fc5ce;
  wire v23f51a6;
  wire v23058b0;
  wire v22fbdb1;
  wire v23094ad;
  wire v23065ad;
  wire v230b4ad;
  wire v23f7039;
  wire v23fbc17;
  wire v23f11a3;
  wire v230f760;
  wire v22f00eb;
  wire v22f1f92;
  wire v2310fb9;
  wire v22eec68;
  wire v230fc8c;
  wire v2301ef1;
  wire v230b8fb;
  wire v22fb941;
  wire v22ee9d5;
  wire v23f83de;
  wire v23fbc0d;
  wire v230a688;
  wire v22fb40c;
  wire v22f6986;
  wire v11853ca;
  wire v230754a;
  wire v22f3eed;
  wire v23fa825;
  wire v22ed631;
  wire v23fbc89;
  wire v23f5e3d;
  wire v22ee681;
  wire bd0733;
  wire v23f4e90;
  wire v22fda63;
  wire v23fce89;
  wire v22f482d;
  wire v22f51b1;
  wire v23fb9bf;
  wire v230a87b;
  wire v22ff79d;
  wire v23115b1;
  wire v2304d0c;
  wire v23fca1b;
  wire v22f6d19;
  wire v23fb777;
  wire v2303fa7;
  wire v23f7632;
  wire v22f30dc;
  wire v22f4d28;
  wire v23fbd7d;
  wire v23f84f9;
  wire v23fcc83;
  wire v23096af;
  wire v1506a7a;
  wire v23f4f13;
  wire v2393769;
  wire v98d402;
  wire v22f2903;
  wire v230bf92;
  wire v22f1037;
  wire v230354e;
  wire v22f8943;
  wire v230aa0d;
  wire v23fbf8b;
  wire v22f61f6;
  wire v230bd36;
  wire v22f26f5;
  wire v22f25ae;
  wire v23f4f88;
  wire v2312050;
  wire v22ef757;
  wire v230c91d;
  wire v23fbf45;
  wire v22f659a;
  wire v23fcdd1;
  wire v23fc85b;
  wire v23fccaf;
  wire v23fb64a;
  wire v23f6079;
  wire v22ffc83;
  wire v22fa9de;
  wire v23fcf82;
  wire v22eeb7a;
  wire v23fbd46;
  wire v23133fe;
  wire v22ed291;
  wire v23f1824;
  wire v23f165d;
  wire v22fb0ac;
  wire bd74b6;
  wire v2301bda;
  wire v23056e9;
  wire v23fc374;
  wire v23fb80e;
  wire v23f5d36;
  wire v23fbbbd;
  wire v2312231;
  wire v13aff86;
  wire v22fa73a;
  wire v23f9d9a;
  wire v22faa39;
  wire v230f9b8;
  wire v23f864d;
  wire v23037b3;
  wire v23f3f36;
  wire v230186e;
  wire v23fb9f8;
  wire v23090fb;
  wire v23fb1e5;
  wire v22f4638;
  wire v22ec08f;
  wire a0b7a3;
  wire bd8ccb;
  wire v22ff08f;
  wire v23fb215;
  wire v22fe7f5;
  wire v23fc551;
  wire v22f9e3d;
  wire v23fb6a7;
  wire v2309456;
  wire v23f6927;
  wire e1df54;
  wire v23f3c84;
  wire v23fb07c;
  wire v23f6bba;
  wire v23fc689;
  wire v22fe147;
  wire v23fc08f;
  wire v22fe116;
  wire v230ea67;
  wire v23fd002;
  wire v23fa94e;
  wire v23fcd42;
  wire v23105b1;
  wire v230cfb5;
  wire v22ee4eb;
  wire v23fb92b;
  wire v150744b;
  wire v2308750;
  wire v22ed1d3;
  wire v22fca3a;
  wire v230313e;
  wire v2306119;
  wire v23009d5;
  wire v22fed90;
  wire v230b9fc;
  wire v23f77a4;
  wire v23fc7a6;
  wire v191afb7;
  wire v22f8f56;
  wire v23fc128;
  wire v2302d53;
  wire v22f48b7;
  wire v23f33b2;
  wire v23f724a;
  wire v22f62e3;
  wire v23fcfd1;
  wire v22f8f70;
  wire v22fee59;
  wire v23123b4;
  wire v23fc51c;
  wire v23fc35f;
  wire v22ffdc5;
  wire v23fbd48;
  wire v22f1a04;
  wire v23934f0;
  wire v22f0b8a;
  wire v230d00c;
  wire v23fc3f3;
  wire v22f2ffc;
  wire v23fc279;
  wire v23fbfb2;
  wire v230887b;
  wire v22ec686;
  wire v22f768b;
  wire v2311a4a;
  wire v23fc92c;
  wire v23f5bf3;
  wire v230e8a6;
  wire v23fc7e2;
  wire v2301a67;
  wire v23fcb0d;
  wire v230da69;
  wire v230f087;
  wire v230b82e;
  wire v22f3f9f;
  wire v23fbabc;
  wire v23067cd;
  wire v2304193;
  wire e1d3f0;
  wire v22f9392;
  wire v23f475e;
  wire v22ee2eb;
  wire v22fced7;
  wire v230abf3;
  wire v22ef659;
  wire v23fc207;
  wire v23fc336;
  wire v2393417;
  wire v22f1ae7;
  wire v22fa6ab;
  wire v23f4bc2;
  wire v22ee521;
  wire v22f0470;
  wire v15070d3;
  wire v23fb8fc;
  wire v22ed1e8;
  wire v23fc209;
  wire v23fc117;
  wire v23fc4a3;
  wire v23fb8d1;
  wire v230638a;
  wire v22fb87a;
  wire v22eb3fc;
  wire v1aae222;
  wire v22f7d67;
  wire v22f814e;
  wire v23fc745;
  wire v22fdca9;
  wire v23f7795;
  wire v23130a1;
  wire v22f94ea;
  wire v22fb272;
  wire v23fb5ec;
  wire v2310319;
  wire v23fc6af;
  wire v2307009;
  wire v23fb9ef;
  wire v22f1683;
  wire v23f7ff2;
  wire v22f07e0;
  wire v23fb8fd;
  wire v22f4bcf;
  wire v23f4bab;
  wire v22f4cf2;
  wire v23f8848;
  wire v22fd0fb;
  wire v23fbff5;
  wire v191b215;
  wire v845625;
  wire v17cf1d8;
  wire v23fbb0e;
  wire v2307d70;
  wire v23fb9d4;
  wire v230c771;
  wire v17cf286;
  wire v845629;
  wire v21eabbd;
  wire v23fbdf1;
  wire v23faaac;
  wire v23fc26e;
  wire v23fb5a2;
  wire v2302d9a;
  wire v230eaba;
  wire v22f166b;
  wire v2309543;
  wire v17a2d5a;
  wire v21ea5eb;
  wire v845635;
  wire v23f1ec4;
  wire v23f4ab4;
  wire v85fd50;
  wire b7d0f1;
  wire v22f30bb;
  wire v23f8e04;
  wire v22f50ae;
  wire v85e5cf;
  wire v23fced3;
  wire v231029e;
  wire v123d721;
  wire v845665;
  wire v230f4d3;
  wire v22f178d;
  wire v22f53f3;
  wire v22fa205;
  wire v23f4c9c;
  wire v2301d76;
  wire v22ef2c3;
  wire v22ede4d;
  wire v23fa882;
  wire v23fc684;
  wire v23fcbb0;
  wire v191ac87;
  wire v230a9ca;
  wire v230b5cc;
  wire v2309520;
  wire v2304568;
  wire v22f3628;
  wire v22f3091;
  wire v23f37bf;
  wire v2307b18;
  wire v23f8b6b;
  wire v22ef2c7;
  wire e1e7b0;
  wire v230c3f5;
  wire v23fd01e;
  wire v23fb11d;
  wire v2308225;
  wire v23039be;
  wire v22fca4e;
  wire v2306c16;
  wire v22f4e94;
  wire v22eb25c;
  wire v22f9a50;
  wire v23f6827;
  wire v2302e76;
  wire v2309d29;
  wire v230083b;
  wire v1507056;
  wire v23fbf6e;
  wire v2312ccb;
  wire v23f6658;
  wire v22f5421;
  wire v2300246;
  wire v231285b;
  wire v22fcabc;
  wire v2304987;
  wire v23fb323;
  wire a6c3d1;
  wire v23fcbbb;
  wire v22fd145;
  wire v22ed48c;
  wire v2391728;
  wire v23f40d6;
  wire v2393739;
  wire v230879e;
  wire v23109fb;
  wire v22f764d;
  wire v22f6066;
  wire v230dc56;
  wire v2308f80;
  wire v23fcbc8;
  wire v23fc120;
  wire v22eeea9;
  wire v230d836;
  wire v2305263;
  wire v23f1133;
  wire v2312dfa;
  wire v230f6d0;
  wire v2312a9e;
  wire v23fc32b;
  wire b09503;
  wire v23f9395;
  wire v23fbe24;
  wire v23fbfbb;
  wire v22f52c1;
  wire b00ad2;
  wire v2308627;
  wire v23f28de;
  wire v23fc76a;
  wire bd7c6a;
  wire v23fb704;
  wire v230a180;
  wire da38b9;
  wire v2304cc3;
  wire v23fc343;
  wire v22edd3f;
  wire v22f14bf;
  wire b9c976;
  wire v23f8caa;
  wire v2312196;
  wire v22f3519;
  wire v23fc941;
  wire v23f6c16;
  wire v23fc2cc;
  wire v23fc5a9;
  wire v22fa7b8;
  wire v2300aab;
  wire v2307061;
  wire v2311918;
  wire v191ae51;
  wire v2300cd4;
  wire v23fc7f9;
  wire v23f347b;
  wire v2306d2c;
  wire v22ffc31;
  wire v23fb4a9;
  wire v230812e;
  wire v22f98ca;
  wire v23fc1ac;
  wire v2302da4;
  wire v2303352;
  wire v22f0ecb;
  wire v22efb46;
  wire v23f51e3;
  wire v2393118;
  wire v23fb9a3;
  wire v22ef607;
  wire v2307f27;
  wire v22ec98c;
  wire v22f7f2a;
  wire v2304421;
  wire v22eb415;
  wire v22f8440;
  wire v2309a46;
  wire v2393900;
  wire v23086c5;
  wire v23126fc;
  wire v230b9b4;
  wire v22ef99b;
  wire v23134bf;
  wire v23f4f3b;
  wire v22fec16;
  wire v23f5558;
  wire v23f68d8;
  wire v23f77d5;
  wire v22f63cc;
  wire v22f82f1;
  wire v230716d;
  wire v230e817;
  wire v23fbe61;
  wire v22fc712;
  wire v23f5156;
  wire v23fcbd7;
  wire v23fc748;
  wire v230cea0;
  wire v22f3813;
  wire v23030e8;
  wire v23fcb44;
  wire v23fb883;
  wire bb324c;
  wire v1e84190;
  wire v23f619d;
  wire v22f42b0;
  wire v2302cce;
  wire v23f3b1d;
  wire v91c376;
  wire v22fd69b;
  wire v23919c0;
  wire v230d6fd;
  wire v23fcbb2;
  wire v23fcfbf;
  wire v2310075;
  wire v23fbe0b;
  wire v23f9033;
  wire v22f7588;
  wire v22effdc;
  wire v23fba4d;
  wire v23fbdc6;
  wire v230ca71;
  wire b00b0b;
  wire v845653;
  wire v22f217d;
  wire v22ecc0d;
  wire v22eec5f;
  wire v23f3051;
  wire v22fe60b;
  wire v22f5c70;
  wire v23fcb61;
  wire v230ec4b;
  wire v845641;
  wire v214cf31;
  wire v23fc8d7;
  wire v23f2216;
  wire v23fce65;
  wire v1b87673;
  wire v22f037a;
  wire v22f1f71;
  wire v2391d0b;
  wire v22f1b3b;
  wire v22f694d;
  wire v230226e;
  wire v22ec20e;
  wire v23039af;
  wire v2308506;
  wire v23fc23b;
  wire v23f1193;
  wire v22ed337;
  wire v22eb3aa;
  wire v23fcdb9;
  wire v23fc2d2;
  wire v230d23a;
  wire b84615;
  wire v22fa771;
  wire v23fb505;
  wire v23f8465;
  wire v23f5e22;
  wire v23fba1a;
  wire v22f0810;
  wire v23fb9ff;
  wire v23f9ca2;
  wire v22f0360;
  wire v2306bf9;
  wire v8abd93;
  wire v23fcd5f;
  wire v191b17f;
  wire ae3590;
  wire v23fbf87;
  wire v22f1ef6;
  wire v23f4761;
  wire v22f9078;
  wire v23f4e43;
  wire v2301e9c;
  wire v230f43d;
  wire v22fb6db;
  wire v230960c;
  wire bd7747;
  wire v23fcc50;
  wire v23058da;
  wire v22f4e2e;
  wire v22fba6d;
  wire v230aa17;
  wire v23021d9;
  wire v2304c95;
  wire v22fbab1;
  wire v22f35eb;
  wire v23fa4cb;
  wire v2304faf;
  wire v22ed07d;
  wire v23fc5d4;
  wire v2392803;
  wire v22f5696;
  wire v22ff4aa;
  wire v22f3dea;
  wire v23fc28d;
  wire v2309305;
  wire v23fbb58;
  wire v23efd8a;
  wire b9ca3d;
  wire v22f426a;
  wire v22f69eb;
  wire v23fb9fe;
  wire v231354e;
  wire v23fcba7;
  wire v2306d22;
  wire v2307c15;
  wire v23f7be0;
  wire v23fcc7c;
  wire v22ee4e7;
  wire v23061de;
  wire v22eec2d;
  wire v23fbd8c;
  wire v23f8e0b;
  wire v22f8105;
  wire v23fc3de;
  wire v23f32eb;
  wire v2302370;
  wire v230a775;
  wire v23f7344;
  wire v22ed53e;
  wire v22f6963;
  wire v23fc0b7;
  wire v22faf4e;
  wire v22ecb28;
  wire v2306656;
  wire v23f6afa;
  wire v2306a6f;
  wire v106a7bd;
  wire v2306c5e;
  wire v23f745f;
  wire v2306e8f;
  wire v23fcbe2;
  wire v23fc35e;
  wire v23fb4f0;
  wire v23fc772;
  wire v23f36f9;
  wire v22f9c37;
  wire v23fce3b;
  wire v23126be;
  wire v2305841;
  wire v23fa7ba;
  wire v22fe50f;
  wire v23fcce5;
  wire v23f8798;
  wire v96bd8b;
  wire v94701c;
  wire v23f35c2;
  wire v22fb151;
  wire v23ef987;
  wire v23fc617;
  wire v22f3a91;
  wire v23f741e;
  wire v2305aa1;
  wire v23f00cf;
  wire v22ee516;
  wire v1e8408b;
  wire v23fc0f5;
  wire v22ebccb;
  wire v12cd993;
  wire v22fdb4e;
  wire v23fc8be;
  wire v23fbe41;
  wire v23f38d5;
  wire v239154a;
  wire v23121aa;
  wire v2307edb;
  wire v2308be0;
  wire v23fb456;
  wire v23fb679;
  wire v22eed1b;
  wire v230a905;
  wire v2346b41;
  wire v22ff1ee;
  wire v23fcb53;
  wire bd9ec5;
  wire v22f6e47;
  wire v22eb6dd;
  wire v23fb4be;
  wire v23011c7;
  wire v23fb132;
  wire v23f7b85;
  wire v230cc50;
  wire v23fcaa7;
  wire v845647;
  wire v23fbfaf;
  wire v23fb481;
  wire v2307b4c;
  wire v23fcd71;
  wire v106ae74;
  wire fc8c68;
  wire v22fcad1;
  wire v23fac2d;
  wire v22ec5d6;
  wire v230440f;
  wire v2391cf8;
  wire v22f8499;
  wire v23fbf48;
  wire v23129fa;
  wire v22f118f;
  wire b11fc3;
  wire v23f9f71;
  wire v1b87890;
  wire v22f334e;
  wire v23fc2dd;
  wire v8d360e;
  wire v22fcdf6;
  wire v1aae56f;
  wire v23fc85c;
  wire v13afe8f;
  wire v106ae21;
  wire v230a759;
  wire v22f95c1;
  wire v84564d;
  wire v23f7af2;
  wire v23fc17d;
  wire v23fa931;
  wire v23f5bdc;
  wire v23fbeb4;
  wire v22f349a;
  wire v22faeec;
  wire v22f7f52;
  wire v22f9911;
  wire v23fb9c2;
  wire fc88ba;
  wire v23fc8a3;
  wire v23021e1;
  wire v2391ab6;
  wire v22fa5b4;
  wire v2302dd1;
  wire v230db9d;
  wire v23f6ac2;
  wire v230f5a3;
  wire v230a83f;
  wire v22f46b1;
  wire v23fb9d9;
  wire v230ad60;
  wire v2303a62;
  wire v230e1f2;
  wire v23fc476;
  wire v23fc8ad;
  wire v23fa524;
  wire v23fba7e;
  wire v1aae29a;
  wire v191ae42;
  wire v23f2873;
  wire v84563e;
  wire v2302ca3;
  wire v23fc2f3;
  wire v23f68bf;
  wire b9c92c;
  wire v230fdc7;
  wire v23f8364;
  wire v22f8ba5;
  wire v22fa36f;
  wire v2312faa;
  wire v23fcc05;
  wire v2305853;
  wire v231026b;
  wire v2392c72;
  wire v191aed3;
  wire a1fe40;
  wire v2393fc1;
  wire v2307150;
  wire v23fc7e7;
  wire v2302131;
  wire v23f74da;
  wire v23fbcc3;
  wire v22eeb4b;
  wire v23fa4ca;
  wire v23fc896;
  wire v22f60da;
  wire v2307b25;
  wire v22fc58a;
  wire v231228e;
  wire b06cee;
  wire v23fc22f;
  wire v2304070;
  wire v2312325;
  wire v2311944;
  wire c17811;
  wire v23faa93;
  wire v23fc7b5;
  wire v23fb732;
  wire v23f711a;
  wire v23f38b1;
  wire v22ebffc;
  wire v22f37c1;
  wire v22f60c6;
  wire v2300c3d;
  wire v2305252;
  wire v191abfa;
  wire v22f79c8;
  wire v2310c54;
  wire v22ec74f;
  wire v23fbcad;
  wire v23fc3a4;
  wire v23fc7d6;
  wire v23fc97a;
  wire v23fc822;
  wire v22ff727;
  wire v22f7d93;
  wire v22f4f0f;
  wire v23f645e;
  wire a1fd0b;
  wire v2309a10;
  wire v23065db;
  wire v2391f9b;
  wire v22fbb7f;
  wire v22fdb25;
  wire v2309094;
  wire v2303632;
  wire aaca7f;
  wire v23fbf1c;
  wire v22f2188;
  wire v22fa262;
  wire v23f7c8d;
  wire v230a66b;
  wire v22f6c3a;
  wire v2306514;
  wire v23f8a06;
  wire v230997b;
  wire v23f4d1c;
  wire v23fbdd4;
  wire v2309221;
  wire v23f20d7;
  wire v22efd1a;
  wire v23fc199;
  wire v22fa827;
  wire v230cb9d;
  wire v22f03aa;
  wire v22eaf7a;
  wire v23f89db;
  wire v22f852d;
  wire v22f78a9;
  wire v23054ba;
  wire v2307729;
  wire a68bda;
  wire v22fc96c;
  wire v23fcc8e;
  wire v2305128;
  wire v230d64e;
  wire v22fa345;
  wire v23efdd0;
  wire v230818b;
  wire v22f1133;
  wire v23f43af;
  wire v23fbec8;
  wire v22f8959;
  wire v22fb7bc;
  wire v22f264f;
  wire v23f529c;
  wire v2392534;
  wire v2392ed3;
  wire v23fc4b4;
  wire b50bc7;
  wire c24eac;
  wire v22eea9a;
  wire v22fa474;
  wire v23fcadf;
  wire v230abce;
  wire v22ebe7f;
  wire v22f9d69;
  wire v23fbe7e;
  wire v23f4cdc;
  wire v2309515;
  wire v22fa1af;
  wire v22ed898;
  wire v23fbb37;
  wire v23ef9c4;
  wire v22f9de9;
  wire v230baba;
  wire v23f23e8;
  wire v22ee269;
  wire v22fdb01;
  wire v22ec71a;
  wire v2303461;
  wire v230813c;
  wire v22ebc25;
  wire v230f538;
  wire v2391e8f;
  wire v230dcf6;
  wire v230f4e5;
  wire v23fbad3;
  wire v22f115b;
  wire v239208c;
  wire v90af77;
  wire v23f90c4;
  wire v230995b;
  wire v23fc1dc;
  wire v23f3a95;
  wire v22fd781;
  wire v22f39b0;
  wire v22fb5b1;
  wire v23fb649;
  wire v23fbed3;
  wire v22ece03;
  wire v23fb1e3;
  wire v2308c31;
  wire v9c12cb;
  wire bd9ab5;
  wire v22fb1f3;
  wire v230bbf8;
  wire v23fb92a;
  wire v230c12c;
  wire a8a256;
  wire v23f9a46;
  wire v230f863;
  wire v22ee03c;
  wire v23f32db;
  wire v22f5355;
  wire v23fcc90;
  wire v22fe362;
  wire v23f710d;
  wire v22f7fd1;
  wire v23fc96d;
  wire v23fc85e;
  wire v23f9110;
  wire v230a5e6;
  wire v23fc126;
  wire v23fcc24;
  wire e1dcf6;
  wire v23fbb74;
  wire v23f2a3d;
  wire v23fcb58;
  wire v230b7c1;
  wire v23fc125;
  wire v23fbae2;
  wire v23f1cd5;
  wire v231241e;
  wire v22f3b94;
  wire v23f4517;
  wire v22f8107;
  wire v22ef1a3;
  wire v23fafc1;
  wire v23f7372;
  wire v23fb4b1;
  wire v230e07e;
  wire v23fbddb;
  wire v23fb5db;
  wire v22f3f15;
  wire v23faaef;
  wire v230feae;
  wire v2307ab9;
  wire v22efa17;
  wire v23fc0c6;
  wire v22f28aa;
  wire v230eeb5;
  wire v2308c3d;
  wire v230e882;
  wire v23fc220;
  wire v23fbd76;
  wire v22f6e0c;
  wire v22f4d69;
  wire v23fc6ac;
  wire v22fb157;
  wire v23f65b4;
  wire v23009f0;
  wire v22fb09f;
  wire v22fcf55;
  wire v23f6f5c;
  wire v23f1b3d;
  wire v23f4872;
  wire v22ee8d8;
  wire v23fc92a;
  wire v23f8ade;
  wire v23fbd94;
  wire v22eea67;
  wire v23fcac8;
  wire v23f7d57;
  wire v23f3c3b;
  wire v22f7713;
  wire v230b464;
  wire v23f34d7;
  wire v2312524;
  wire v23fc4dd;
  wire v22f4bf5;
  wire v230aabf;
  wire v23fb793;
  wire v2302992;
  wire v23fcc2a;
  wire v23f73af;
  wire v23fb3f3;
  wire v23f05c0;
  wire v23fc6e0;
  wire v23fc989;
  wire v22f5ea8;
  wire v2301cf4;
  wire v23fc8f3;
  wire v22ee8ee;
  wire v22f4339;
  wire v22fef14;
  wire v22f7f12;
  wire v2312d2c;
  wire v230592c;
  wire v23038cc;
  wire v23f5f62;
  wire v23f15ba;
  wire v22f476c;
  wire v23fc116;
  wire v2309a51;
  wire v22f3294;
  wire v22fab99;
  wire v13afe3a;
  wire v23fc46b;
  wire v1e84038;
  wire v231008b;
  wire v22fca12;
  wire v23fccc6;
  wire v2308f7f;
  wire v23fbe89;
  wire v23fc5de;
  wire v23930d8;
  wire v86d5f2;
  wire v23fbab6;
  wire v22f9a6b;
  wire v23f7456;
  wire v23104db;
  wire v23fb4a4;
  wire v230177d;
  wire v2313264;
  wire v2306775;
  wire v23fcb5d;
  wire v22f0eec;
  wire v231066c;
  wire v22fed4e;
  wire v22f80ca;
  wire v191a90b;
  wire v22f0362;
  wire v23f8ecc;
  wire v23efe10;
  wire v22fa4dd;
  wire v2308d79;
  wire a1fd35;
  wire v2312f7e;
  wire v23fcd09;
  wire v23fb77e;
  wire v22faa1f;
  wire v230204f;
  wire v23f9904;
  wire v230b364;
  wire v23022b1;
  wire v12cdba9;
  wire v22fec20;
  wire v22f8db2;
  wire v23fba3a;
  wire v23131e8;
  wire v2302e73;
  wire v2306220;
  wire v22f1d96;
  wire v9ad58e;
  wire v23fb73d;
  wire v23f63b2;
  wire v23f8914;
  wire v23027e9;
  wire v230f578;
  wire v9bd8c6;
  wire v22f79de;
  wire v106a7d6;
  wire v22f91c9;
  wire v12ce195;
  wire v2392974;
  wire v22f8626;
  wire v23fcf5e;
  wire v23125ee;
  wire v22ff0da;
  wire v1506a4c;
  wire v23088ef;
  wire v22f9183;
  wire v23fc91c;
  wire v23fc7ca;
  wire v23fc514;
  wire v230cf2f;
  wire v23fad53;
  wire v230f2ef;
  wire v2309c9d;
  wire v230248b;
  wire v23fb9ad;
  wire v22febe7;
  wire v23101ee;
  wire v22f163a;
  wire v23fc02b;
  wire v230f165;
  wire v2300b80;
  wire v22ef109;
  wire v23fceb2;
  wire v22ffad4;
  wire v23fb7d7;
  wire v22f6315;
  wire v23fce25;
  wire v23fc1c4;
  wire v22f9414;
  wire v23f4a02;
  wire v23fc232;
  wire v23f2602;
  wire v23018ac;
  wire v23f8607;
  wire v22f1dc4;
  wire v22f8985;
  wire v22f38db;
  wire v22f444f;
  wire v2306e3c;
  wire v22fe44f;
  wire v22fa736;
  wire v191acbd;
  wire v2393f05;
  wire v23f28ed;
  wire v22f2b42;
  wire v22ecd3a;
  wire v23fbd08;
  wire v23f033c;
  wire v23f2fe0;
  wire v23f6bf3;
  wire v22f9369;
  wire v22f3959;
  wire v2391f3b;
  wire v23fb98d;
  wire v22f2d83;
  wire v230d630;
  wire v23fc8f9;
  wire v2308b7c;
  wire v22faee9;
  wire v231171d;
  wire v22f1cbc;
  wire v2307a62;
  wire v230de91;
  wire v23f1ccc;
  wire v22fe1d9;
  wire fc8c27;
  wire v23f616b;
  wire v230e821;
  wire v23f4bfc;
  wire v23f581f;
  wire v239160b;
  wire v23fbefa;
  wire v23f8f21;
  wire v2308ae2;
  wire v23fbbd2;
  wire v231339c;
  wire v23f8638;
  wire v2306885;
  wire v2310da0;
  wire v23fcf65;
  wire v23fba13;
  wire v2303393;
  wire v22fa055;
  wire v2309465;
  wire v230065b;
  wire v230a193;
  wire v23fa720;
  wire v22f3c9a;
  wire v2301a7d;
  wire v22f19a0;
  wire v23f73dd;
  wire v22fd311;
  wire v22fca75;
  wire v230cec5;
  wire v22ed2e5;
  wire v23f9bcf;
  wire v22fe9dc;
  wire v23f2698;
  wire v22fe19b;
  wire v2310bdf;
  wire e1de18;
  wire v23fac5a;
  wire v23f266b;
  wire v23f1eb7;
  wire v22fb147;
  wire v23fc449;
  wire v2309d0b;
  wire v22f25ed;
  wire v230913d;
  wire v22ebb85;
  wire v2311f99;
  wire v22f07ac;
  wire v23fcd91;
  wire v23f89f4;
  wire v23fc628;
  wire v23fc9eb;
  wire v23fc93b;
  wire v22fc90d;
  wire v22f87bf;
  wire v22f5019;
  wire bd94fd;
  wire v230649c;
  wire v22ec5f2;
  wire v230cd17;
  wire v23133be;
  wire v231016f;
  wire v22f6d27;
  wire v2301b38;
  wire v23f8a5e;
  wire v22f947f;
  wire v2306b99;
  wire v23f4928;
  wire v23fbedd;
  wire v23f818e;
  wire v2312bae;
  wire v22ef7a7;
  wire v23f4ad7;
  wire v23007d9;
  wire v845657;
  wire v2302c31;
  wire v13afc19;
  wire v22f975b;
  wire v22f7ad5;
  wire v230429d;
  wire v23f522c;
  wire v22ff12b;
  wire v23f90b2;
  wire v230bb92;
  wire v23fc549;
  wire v23f895d;
  wire v23fb1b9;
  wire v22ff882;
  wire v230dcf9;
  wire v23fc5f5;
  wire v2311629;
  wire v22f2c72;
  wire v23f6acc;
  wire v84562e;
  wire v23f06d7;
  wire v23fabb8;
  wire v2308a32;
  wire v230d2b0;
  wire v23fb5b7;
  wire v23f1391;
  wire v23075ce;
  wire v22fdaf3;
  wire v230c7f6;
  wire v22f7be4;
  wire v23f1354;
  wire v23fc139;
  wire v23f91bc;
  wire v23f2810;
  wire v2303fb2;
  wire v22fa9f7;
  wire v22ed494;
  wire v23fc1d3;
  wire v23fba28;
  wire v23f3dcc;
  wire v23fc1fc;
  wire v22f6277;
  wire v22f8cce;
  wire v23fb828;
  wire v23fc965;
  wire v23fa3b6;
  wire v23fb9fc;
  wire v84562d;
  wire v23f537e;
  wire v230fe27;
  wire v23040c8;
  wire v23f85b6;
  wire v230ecb1;
  wire abf9f6;
  wire v2309eb8;
  wire v22fd79d;
  wire v22ef76f;
  wire v2304856;
  wire v23fcb80;
  wire v23fbd92;
  wire v22ebe52;
  wire v230ed31;
  wire v23fca8a;
  wire v23f6da6;
  wire v23fba0d;
  wire v23f85a9;
  wire v2307e5a;
  wire v23067de;
  wire v106a888;
  wire v2303a58;
  wire v23fccc1;
  wire v23fcb24;
  wire v23fcec1;
  wire v23fc521;
  wire v2305a91;
  wire b61053;
  wire v23f9f9d;
  wire v23046be;
  wire v22f4af1;
  wire v23fc56c;
  wire v2310e5d;
  wire v23fc627;
  wire v22fb1d7;
  wire v23fc1a1;
  wire v22ebc8f;
  wire v22f95e4;
  wire v22f674b;
  wire v23fb671;
  wire v23018f1;
  wire v230aa94;
  wire v22f0bea;
  wire v2312fc4;
  wire v23f6b25;
  wire v230c963;
  wire v22fc020;
  wire v22eba71;
  wire v23fbaa2;
  wire v23fc22c;
  wire v23fcdb0;
  wire v23f4c50;
  wire v22f5828;
  wire v2308a7d;
  wire v23fb58e;
  wire v230c3ee;
  wire v23f6325;
  wire v1507a21;
  wire v22f4b6d;
  wire v23fbf73;
  wire v23fbf58;
  wire aca9e4;
  wire f4067f;
  wire v2391a57;
  wire v23f9fc1;
  wire v22ff4eb;
  wire v22fc9ad;
  wire v23f3d62;
  wire v23fbc82;
  wire v230c1dd;
  wire v23fbc6d;
  wire v23f7206;
  wire v22f19cb;
  wire v22f167b;
  wire v2309e42;
  wire v23f651a;
  wire v22ffa6e;
  wire v230e97b;
  wire v12cd570;
  wire v2305024;
  wire v22fe852;
  wire v2303154;
  wire f40ab9;
  wire v23fbb55;
  wire v23fbd69;
  wire v230b4c5;
  wire v22fe098;
  wire v22f1e46;
  wire v23f67fe;
  wire v23fb97c;
  wire v2302983;
  wire v22f2db6;
  wire v23fbe30;
  wire v23041ab;
  wire v2311761;
  wire v23fb9c7;
  wire e1df52;
  wire v2310c26;
  wire v23f2f5d;
  wire v23f439b;
  wire v230648c;
  wire v23f4dd0;
  wire v22f96f1;
  wire v23fc2c1;
  wire v23f2856;
  wire v2308c76;
  wire v23fbe91;
  wire v23fd008;
  wire v1aadcf6;
  wire v23f37b9;
  wire v22f6b4e;
  wire v2393909;
  wire v230a510;
  wire v230f857;
  wire v22fbe9e;
  wire v22ed8b0;
  wire v2300ce0;
  wire v22f779a;
  wire v22f1c40;
  wire v22eebf5;
  wire v2302812;
  wire v22f2286;
  wire v22efb8e;
  wire v2310d59;
  wire v230193c;
  wire v23fc3ca;
  wire v22eee15;
  wire v2311668;
  wire v23088a9;
  wire v23126b7;
  wire v2310538;
  wire v23fcfa1;
  wire v23fcd5c;
  wire v23fb622;
  wire v23fb062;
  wire v2300e92;
  wire v23fb8c7;
  wire v23fb565;
  wire v23f5d72;
  wire v12cd900;
  wire v22ebccd;
  wire v22f2e61;
  wire v23006ef;
  wire v23f95c3;
  wire v230a8b2;
  wire v22ed8a3;
  wire v22f3af7;
  wire v23f3856;
  wire v23f329a;
  wire v23fcefc;
  wire v23f60dc;
  wire v230e568;
  wire v23fc300;
  wire v23fc2f2;
  wire v230b7f4;
  wire v22f23a1;
  wire v230104a;
  wire v22eddd9;
  wire v22ecf6c;
  wire v23fb41a;
  wire v23fba81;
  wire v2307d30;
  wire v1aad8a4;
  wire v22f7b3e;
  wire v23fbe6d;
  wire v12cd66d;
  wire v22f95ec;
  wire v23091ce;
  wire v22f0dd3;
  wire v22eb629;
  wire v230a0e7;
  wire v22fe1e5;
  wire v2310e53;
  wire v23fc3b9;
  wire v22f0a19;
  wire v23f5927;
  wire v22f5088;
  wire v1aad67e;
  wire v22eaec3;
  wire v23fc25b;
  wire v22fd49d;
  wire v1aae1af;
  wire v22fdd6b;
  wire v2303841;
  wire v2313637;
  wire v22fbf19;
  wire v23fb88f;
  wire v23f9945;
  wire v23fc6f5;
  wire v23fbbec;
  wire fc8e3a;
  wire v23fc4f5;
  wire v22eec21;
  wire v22ecbb2;
  wire v22ec96a;
  wire v23fce7f;
  wire v22eb657;
  wire v23fbc28;
  wire v230b930;
  wire v845645;
  wire v22f5edf;
  wire v23f4540;
  wire v22f3196;
  wire v230664e;
  wire v23081e8;
  wire v22fa851;
  wire v231363a;
  wire v23fba5a;
  wire v1aad6a6;
  wire v23fb1c5;
  wire v2309cb5;
  wire v231009b;
  wire v12cd692;
  wire v23fc27c;
  wire v23ef915;
  wire v230e760;
  wire v230f92a;
  wire v2309733;
  wire v23fb593;
  wire v23fcb43;
  wire v22ef9aa;
  wire v23fcecb;
  wire v23f733f;
  wire v2304be0;
  wire v230042c;
  wire v2306540;
  wire v23fc1e1;
  wire v191ae90;
  wire v23fcd90;
  wire v2308e49;
  wire v23fc081;
  wire v191b0f9;
  wire v2392a17;
  wire v22f7e4a;
  wire v22ffe51;
  wire v23f3dd3;
  wire v23fb2e9;
  wire v23f31a9;
  wire v22f7c44;
  wire v191b0e4;
  wire v23fc017;
  wire v22fd8f6;
  wire v2303fd8;
  wire v23fb933;
  wire v22ed458;
  wire v22ef513;
  wire v23fa2d6;
  wire v22fb3ef;
  wire v2304899;
  wire v23fc3e1;
  wire v22f7375;
  wire v23f1fad;
  wire v23f1387;
  wire v23fc1fa;
  wire v230b267;
  wire v2307d7f;
  wire v23f3fb6;
  wire v230acb5;
  wire v2303c5b;
  wire v22f8aa0;
  wire v22f443a;
  wire v23047f9;
  wire v22f779f;
  wire v2302c4b;
  wire fc8ab7;
  wire v8c2b38;
  wire v230a3f5;
  wire v2307942;
  wire v2312cd5;
  wire v22ebd85;
  wire v1e84028;
  wire v230d1c3;
  wire v2312cad;
  wire v22ef848;
  wire v23fc2bc;
  wire v23fbba6;
  wire v2301b06;
  wire v23fc983;
  wire v23088b3;
  wire v23fcea3;
  wire v2307f3f;
  wire v2306eb5;
  wire v23fbb50;
  wire v2305797;
  wire v23fcf4b;
  wire v23fc0cd;
  wire v22ee41e;
  wire v23f9c7f;
  wire v230b713;
  wire v23f9666;
  wire v23f70c6;
  wire v23fccbf;
  wire v23fcb8d;
  wire v23f2e65;
  wire b533b5;
  wire v22ec5ac;
  wire v23fa08a;
  wire v23f9fb5;
  wire v2312cb7;
  wire v1aada6e;
  wire v23fb8f3;
  wire v23fb90b;
  wire v2311919;
  wire v22f43c9;
  wire v23fcdf8;
  wire v22f5033;
  wire v22ffde1;
  wire v1aad441;
  wire v23fbb27;
  wire v22f2939;
  wire v845655;
  wire v230b2a1;
  wire v22eda04;
  wire fc8c9b;
  wire v22fb386;
  wire v23fcb89;
  wire v23f7326;
  wire v23fb95d;
  wire v2307e48;
  wire v23fc722;
  wire v22f6e51;
  wire v845663;
  wire v22ed56a;
  wire v2307460;
  wire v2309891;
  wire v23fcb2b;
  wire v23fc296;
  wire v23f06c9;
  wire v23056b2;
  wire v23fc523;
  wire v23fc855;
  wire v23f3499;
  wire v230e3d1;
  wire v22ee274;
  wire v23fa599;
  wire v23fc9f2;
  wire v2311e03;
  wire v22f1697;
  wire v22f04c8;
  wire v8b5388;
  wire v230d4b4;
  wire v22f62dc;
  wire v22ff9d7;
  wire v23fb672;
  wire v23f0aec;
  wire v2310b8a;
  wire v22ec2cb;
  wire v23f854f;
  wire v230d82c;
  wire v22f69c6;
  wire v23ef4b1;
  wire v22ef3d1;
  wire a878fd;
  wire v2304edd;
  wire v22f43cf;
  wire v22f349c;
  wire v23036c1;
  wire v23fc856;
  wire v2303cc1;
  wire v2308cec;
  wire v22f725a;
  wire v23f6ba0;
  wire v2305114;
  wire v23fc907;
  wire v22f517e;
  wire v23f9ee2;
  wire v22feb20;
  wire v22f154e;
  wire v23fc943;
  wire v2301f50;
  wire v22f7b24;
  wire v22ff294;
  wire v23f88a1;
  wire v23fc5b7;
  wire v23f5109;
  wire v2307c06;
  wire bd770f;
  wire v23fbc19;
  wire v23f40fd;
  wire v22f380e;
  wire v22fc03b;
  wire v23124e2;
  wire v230471d;
  wire v23fc027;
  wire v23fc95c;
  wire ae1a21;
  wire bd953c;
  wire v2301400;
  wire v23f65b6;
  wire v2308748;
  wire v23fc5d9;
  wire v22fa3e9;
  wire v23f5d23;
  wire v22fb335;
  wire v22f2453;
  wire v2311899;
  wire v230cf0c;
  wire v22fd171;
  wire v2302cf5;
  wire v2304598;
  wire v22fc163;
  wire v22ed220;
  wire v22eb95e;
  wire v23fbd3a;
  wire v22f5898;
  wire v230adfa;
  wire v22fd030;
  wire bebe64;
  wire v22f3673;
  wire v1e83f7f;
  wire v2393e5c;
  wire v22f7ca0;
  wire v9526ac;
  wire v845667;
  wire v23f54be;
  wire v22ec87b;
  wire a1fba6;
  wire v22f00c6;
  wire v22fe2a8;
  wire v2302149;
  wire v22f5353;
  wire v23fbfe9;
  wire v230d58c;
  wire v231096b;
  wire v22fd796;
  wire v23fb861;
  wire v23134a0;
  wire v230efeb;
  wire v2305c24;
  wire v23fc002;
  wire a1fbb6;
  wire v238ae11;
  wire v23fb875;
  wire v23fc048;
  wire v22f207c;
  wire v23fc07e;
  wire v2311246;
  wire v230cc30;
  wire v230de17;
  wire v23f8fd7;
  wire v23f1eac;
  wire v230933a;
  wire a1fbc2;
  wire b00ac4;
  wire v22eb377;
  wire v23f8a97;
  wire v2300d5f;
  wire v22ee956;
  wire v230e857;
  wire v2391fc6;
  wire v23f972e;
  wire v1506fe9;
  wire v230fb96;
  wire v230ad18;
  wire v23fc1b9;
  wire v22f3ed0;
  wire v23f98ab;
  wire v22f368e;
  wire v22f8fe0;
  wire v22ff732;
  wire v230d8af;
  wire bf150c;
  wire v23fc975;
  wire v22ec150;
  wire v23fd00e;
  wire v1aad346;
  wire v23f0588;
  wire v23fba06;
  wire v23fca4b;
  wire v23fc69f;
  wire v23052dd;
  wire v23fba6a;
  wire v23f397b;
  wire v230abc9;
  wire v23fbf54;
  wire v230aa9b;
  wire v2304074;
  wire v22f8ee3;
  wire v230966c;
  wire v23f223a;
  wire v2393c3f;
  wire v231142b;
  wire v2301567;
  wire v230945e;
  wire v22f8420;
  wire v23fc329;
  wire v2310b4d;
  wire v22edcce;
  wire v230e1e0;
  wire v23fcd83;
  wire v22f1afb;
  wire v22f85f6;
  wire v2311810;
  wire v2311559;
  wire v23fcd28;
  wire v23fc6a1;
  wire v23fa967;
  wire v23fcae8;
  wire v23fb1c6;
  wire v22f9ac5;
  wire v23fb957;
  wire v22fa4a3;
  wire v2307ffd;
  wire v23fbd6c;
  wire v2304bcd;
  wire v2312e30;
  wire v23fbdf8;
  wire v912a31;
  wire v22fb427;
  wire a72160;
  wire v23f5ab1;
  wire v230aded;
  wire v23fbc3f;
  wire v2307e0c;
  wire v23fbfd5;
  wire v2306593;
  wire v230b38b;
  wire v22faa19;
  wire v22f6ae5;
  wire v23fc94d;
  wire v230be9e;
  wire v23fcf63;
  wire v22f41c4;
  wire v23fbebe;
  wire v230fe6b;
  wire v23013f8;
  wire v22f5429;
  wire v22fe0cb;
  wire v2306da6;
  wire v22fd841;
  wire v22eb563;
  wire v23fc2dc;
  wire v2308b9a;
  wire v23fc46c;
  wire v22f2b34;
  wire v23fbb85;
  wire v22f9f2a;
  wire v22fd445;
  wire v22fcb9d;
  wire v22f2d26;
  wire v22f75b0;
  wire v23f7f35;
  wire v2392867;
  wire v22f23e6;
  wire v2310047;
  wire v23f558b;
  wire v23fd02c;
  wire v23f5019;
  wire v1aadb95;
  wire v22f6058;
  wire v22fc835;
  wire v23fbcff;
  wire v22fa682;
  wire v2304283;
  wire v22eed66;
  wire v23fc3cb;
  wire v2391fae;
  wire v22f3754;
  wire v23001a4;
  wire v23101b1;
  wire v22fb4ab;
  wire v22f94a7;
  wire v22fd767;
  wire v90aa06;
  wire v22f3499;
  wire v22f3b3c;
  wire v23fbaaa;
  wire v23050c1;
  wire v23f447e;
  wire v2303e9a;
  wire v23fb57d;
  wire v22f288e;
  wire v13afeef;
  wire v230d61c;
  wire v22f7928;
  wire v22ecf87;
  wire v22ff58f;
  wire v23f243b;
  wire v22f01c1;
  wire v23fcfdb;
  wire v22ffdf8;
  wire v230a02b;
  wire v230dcef;
  wire v22f4855;
  wire v22f5eae;
  wire v231108b;
  wire v2310904;
  wire v23f8747;
  wire v22ee195;
  wire v23fca1e;
  wire v22f47fe;
  wire v22f8d11;
  wire v23fb993;
  wire f40a94;
  wire v2310434;
  wire v230b8ff;
  wire v22f0d2b;
  wire v23fb8a0;
  wire v23fc676;
  wire v23fbcf8;
  wire v22ffd22;
  wire v230aec0;
  wire v22ef469;
  wire v23fc054;
  wire v23fc388;
  wire v23fc8df;
  wire v23fbacb;
  wire v23fb53b;
  wire v23fb999;
  wire v230ebb1;
  wire v230b837;
  wire v22f95a4;
  wire v23fb5ba;
  wire v23fccb7;
  wire v23f69e4;
  wire v1507439;
  wire v23fc763;
  wire v22ecd54;
  wire v23fc0d8;
  wire v22f1874;
  wire v22fa20a;
  wire v22fb891;
  wire v22ee495;
  wire v230f105;
  wire v23fd060;
  wire v2391f3c;
  wire v23fbaa8;
  wire v2312f45;
  wire v23fc253;
  wire v230f453;
  wire v22f8387;
  wire v22f122e;
  wire v23106e3;
  wire v231140d;
  wire v15070fa;
  wire v23011a9;
  wire v87c96d;
  wire v23fb5ee;
  wire v230339f;
  wire v23f62d5;
  wire v23fb52d;
  wire v2301b70;
  wire v23fac09;
  wire v23f5fe3;
  wire v22fa6c0;
  wire v22fc1be;
  wire v23038a2;
  wire v23f8c7b;
  wire v22f2998;
  wire v23fcced;
  wire v23fbcd0;
  wire v22f6756;
  wire v2303a74;
  wire v22fc5d8;
  wire v2301b52;
  wire v22f43fb;
  wire v23f494b;
  wire v22ed495;
  wire v23fbddf;
  wire v23fcb6f;
  wire v23fc8d2;
  wire v23f01f8;
  wire v23f2504;
  wire v22eb49d;
  wire v23fbb42;
  wire v230b789;
  wire v23fc5ab;
  wire v23fc555;
  wire v230952f;
  wire v2312ad7;
  wire v23fc05d;
  wire v2307c9a;
  wire v230e4c7;
  wire v23028ef;
  wire baf3e5;
  wire v22f6dee;
  wire v22f1ab6;
  wire v23f7fe8;
  wire v23fb045;
  wire v22f7fed;
  wire v23125ab;
  wire v23fbeae;
  wire v230fe82;
  wire v2301937;
  wire v23fbb28;
  wire v22fc7e5;
  wire a89109;
  wire v1aae374;
  wire v23fc357;
  wire v86e576;
  wire v2300834;
  wire v22f6169;
  wire v23f781b;
  wire v230adbf;
  wire v2302348;
  wire v22f036f;
  wire v22fc66c;
  wire v2312919;
  wire v2307ee4;
  wire v22f5280;
  wire v23f0fd1;
  wire v23fcee2;
  wire v22f80b8;
  wire v23fcf5c;
  wire v230d5ab;
  wire v22f19a1;
  wire v2304e69;
  wire v22f20d3;
  wire v23fc4b2;
  wire v230972f;
  wire v23fb489;
  wire v23f8deb;
  wire v23f3472;
  wire v23fc8bb;
  wire v23fc22e;
  wire v22ee1b8;
  wire v23fc48e;
  wire v23064ce;
  wire v23fc79d;
  wire v22f4626;
  wire e1e1d4;
  wire v23fc798;
  wire v23f7066;
  wire v230c132;
  wire v22f149c;
  wire v22f24ca;
  wire v230c37d;
  wire v22feb5c;
  wire b0fad6;
  wire v22f7fcc;
  wire v22f1a8f;
  wire v23027b1;
  wire v22f248e;
  wire v22f0acc;
  wire v22f4af5;
  wire v22f8986;
  wire v23f5cfd;
  wire v22fc5ad;
  wire v23fa0aa;
  wire v23fc3d4;
  wire v231057b;
  wire v22ef648;
  wire v23fce64;
  wire v2309598;
  wire v2302c28;
  wire v22f2195;
  wire v22f7dd1;
  wire v22f469a;
  wire v22eb5dd;
  wire v239346f;
  wire v23fba42;
  wire v1507446;
  wire v23f88d9;
  wire v230a1c7;
  wire v22f2f16;
  wire v22fc3c7;
  wire v2310cbb;
  wire v22f803b;
  wire v230539c;
  wire v23050ee;
  wire v23fb64e;
  wire v22f317b;
  wire v90eab4;
  wire v23fc1d1;
  wire v2311790;
  wire v22fbc04;
  wire v22fca43;
  wire v23f147c;
  wire v23fce61;
  wire v2304e0f;
  wire v22ed7da;
  wire v2305992;
  wire v22f99e9;
  wire v230ff65;
  wire v23fc03d;
  wire v1507246;
  wire v23f87e4;
  wire v23fbf90;
  wire v23f1925;
  wire v22fe0b0;
  wire v230d4cc;
  wire v230a9f0;
  wire v23fbbcf;
  wire v23f9a06;
  wire v22fd7ea;
  wire v22f0295;
  wire v23fbd52;
  wire v22fb32a;
  wire v22eee99;
  wire v23fc71a;
  wire v2392254;
  wire v22f4727;
  wire v22faa40;
  wire v230074c;
  wire v230f27a;
  wire v23fbd11;
  wire v22ec8d1;
  wire v22ed212;
  wire v23f965c;
  wire v22ee60e;
  wire v23f0903;
  wire v230ba09;
  wire v23fb8d6;
  wire v23fc8d6;
  wire v230d921;
  wire be9b63;
  wire v23fcbc3;
  wire v230bd77;
  wire v23f8b5b;
  wire v22f5495;
  wire v230ba79;
  wire v23f7891;
  wire v2313504;
  wire v22f2a1b;
  wire v23fb89c;
  wire v22ee142;
  wire v23066bc;
  wire v22f5cd9;
  wire v22fbebb;
  wire v23084cc;
  wire v23fc39d;
  wire v23fc786;
  wire v2300e6b;
  wire v2306f00;
  wire v23f49b3;
  wire v23fcba5;
  wire v23fb0ce;
  wire v23f5e8a;
  wire v2300617;
  wire v22f482a;
  wire v22ff0d3;
  wire v22fd0b6;
  wire v2303fa1;
  wire v23fc815;
  wire v230c949;
  wire v23f34e1;
  wire v8f9141;
  wire v22f0f7c;
  wire v8dd9c7;
  wire aba695;
  wire v23f4cc5;
  wire v23009cc;
  wire v23fb83c;
  wire v23fba61;
  wire v22f04a6;
  wire v22ebc3c;
  wire v2312577;
  wire v2308a71;
  wire v231072a;
  wire v23f3c77;
  wire v1aad31a;
  wire v22fe869;
  wire v22ec88f;
  wire v2309939;
  wire v230e191;
  wire v23041c1;
  wire v23080ab;
  wire v230b4d9;
  wire v23f8e6b;
  wire v22f2e7b;
  wire v231147e;
  wire v22f6d6e;
  wire v23f3508;
  wire a1fdac;
  wire v22fae03;
  wire v230817b;
  wire v23f999c;
  wire v23fcb23;
  wire v23f80e9;
  wire v22f8594;
  wire v230a774;
  wire v23fc2e8;
  wire v22f7ec4;
  wire v23fc2c8;
  wire v23fb8be;
  wire v22f80b4;
  wire v2387c09;
  wire v23042b7;
  wire v22f2c8a;
  wire v22f59bd;
  wire v22ec1b1;
  wire v23f8d91;
  wire v2300e70;
  wire v2312009;
  wire v22fdb07;
  wire v230d82a;
  wire v22f6955;
  wire v23fcf6b;
  wire v23fbf83;
  wire v230e312;
  wire a1f79d;
  wire v230b282;
  wire v230abf9;
  wire v22ee3e8;
  wire v22fc837;
  wire v23a2d0a;
  wire v230cfe6;
  wire v230d2c2;
  wire v238c168;
  wire v22f17ca;
  wire v1506f9f;
  wire v22efee2;
  wire v231033b;
  wire v23f20d3;
  wire v22f0567;
  wire v23fa623;
  wire v2310d04;
  wire v23f99a0;
  wire v23f40ab;
  wire v23f58e5;
  wire v22f8f27;
  wire v2304990;
  wire v22effdf;
  wire v2301884;
  wire v230ef0b;
  wire v230829b;
  wire v23039c8;
  wire v22f85c2;
  wire bd7c9b;
  wire v2304b35;
  wire v23fbd53;
  wire bc96dd;
  wire v23f1b3c;
  wire v22fcce6;
  wire v22ff05e;
  wire v23fcc35;
  wire v22fea26;
  wire v23fc50a;
  wire v230beed;
  wire v23f1a1c;
  wire v22f40e3;
  wire v2307b06;
  wire v23fcaef;
  wire v15074eb;
  wire v23fcc72;
  wire v230dd28;
  wire v23fc00b;
  wire v2392cce;
  wire v23fbea0;
  wire b425f1;
  wire v22ec9fa;
  wire v23fc48f;
  wire v23fcc2e;
  wire v23f54f7;
  wire v2308e85;
  wire v23fc5ff;
  wire v23f93e7;
  wire bd7497;
  wire v22f5076;
  wire v23f9aa8;
  wire v23fc410;
  wire v23f89fd;
  wire v22f2214;
  wire v22f70b0;
  wire v22fd74b;
  wire v22f3dc7;
  wire v23107f5;
  wire v22f0cc4;
  wire v22f1d80;
  wire v22fb00c;
  wire v22f4b91;
  wire v22edc14;
  wire b00aa0;
  wire v2304abd;
  wire v22ff259;
  wire v2303051;
  wire v22ef100;
  wire v23fbe7d;
  wire v22ffa07;
  wire f40764;
  wire f40618;
  wire v23fb4cb;
  wire v23fb6ff;
  wire v22fe920;
  wire v22f8cb9;
  wire v23f052e;
  wire v23fc823;
  wire v23fc778;
  wire v23fbd89;
  wire v22eb404;
  wire v230da2f;
  wire v22efd02;
  wire v23fc11b;
  wire v12cd9f9;
  wire v23fb906;
  wire v22f40ef;
  wire v2312f1b;
  wire v23fca4e;
  wire v23065d3;
  wire v23fbace;
  wire v2393142;
  wire v22f4619;
  wire v23fba74;
  wire v22ff3e6;
  wire v23fc89b;
  wire v23f86a0;
  wire v2312b9e;
  wire v2308db0;
  wire v22f57d4;
  wire v22fa819;
  wire v230070e;
  wire v22fcd80;
  wire v23fbb53;
  wire v23f3e68;
  wire v23f0dc7;
  wire v23fc453;
  wire v23f8986;
  wire v22f24f8;
  wire v22fda59;
  wire v23f3346;
  wire v23f51da;
  wire v22f7ed8;
  wire v230fd1c;
  wire v2301105;
  wire v23fb818;
  wire v23fc9dd;
  wire v23fcd00;
  wire v23122cf;
  wire v22eb8ae;
  wire v23f598e;
  wire v2312cb9;
  wire v2311da7;
  wire a1fdd3;
  wire v230e896;
  wire v22eb015;
  wire v230ec04;
  wire v230b0f2;
  wire v23fc880;
  wire v9ed019;
  wire v2307eac;
  wire v2311d05;
  wire v230f18c;
  wire v1aad45d;
  wire v23fccb5;
  wire a8ec08;
  wire v23fc458;
  wire ad78c9;
  wire v22f8a0c;
  wire v908162;
  wire v230bf72;
  wire v2302dca;
  wire v22f5c1a;
  wire v2305a52;
  wire v191abed;
  wire v23f76fb;
  wire v23139c9;
  wire v22fe7ca;
  wire v23fbf31;
  wire v23fcaf6;
  wire v22f3832;
  wire v22f05b4;
  wire v22fe6f8;
  wire b0d6e5;
  wire v23fb555;
  wire v230ffae;
  wire v230d533;
  wire v23fb5cf;
  wire v9122cc;
  wire v22efadc;
  wire v22efd99;
  wire v2303efa;
  wire v23fccfd;
  wire v22f6534;
  wire v22f4ef0;
  wire v1aadad9;
  wire v2393495;
  wire v23f8d36;
  wire v23f41ec;
  wire v23f2f8d;
  wire v23fbc37;
  wire v23fcc52;
  wire v230f1d6;
  wire v22fb22e;
  wire v2300686;
  wire v2310852;
  wire v22fbd9a;
  wire v22ecc5a;
  wire v23fc15b;
  wire v2301dad;
  wire v2305a14;
  wire v22fb7e0;
  wire v23045ae;
  wire v22ee3a3;
  wire v230c2f3;
  wire v23fb922;
  wire v22fb417;
  wire v22eed25;
  wire v22f4db6;
  wire a9da2d;
  wire v22eb3bc;
  wire v23f50d9;
  wire v22ed363;
  wire v22f1aed;
  wire v977ddf;
  wire bd6575;
  wire v23f52c1;
  wire v22fae48;
  wire v23f80cc;
  wire v22eef66;
  wire v23f089b;
  wire v23fccd4;
  wire v22f4016;
  wire v23f8c22;
  wire v22f991d;
  wire v22f12e5;
  wire v23fced9;
  wire v22fe495;
  wire v23fb7fc;
  wire v22fba9a;
  wire v2304184;
  wire v23fc6ca;
  wire v22f8427;
  wire v23f4008;
  wire v23f39fb;
  wire v23fbbc3;
  wire v13afb6e;
  wire v2309783;
  wire v22fe370;
  wire v23fbedf;
  wire v23fcaf1;
  wire v230058a;
  wire v22f9801;
  wire v23f97c6;
  wire v2309459;
  wire v23fbb39;
  wire v23fa2eb;
  wire v23fb17e;
  wire v1aadf2f;
  wire v9799b6;
  wire v22ef3aa;
  wire v23fb4e6;
  wire v230b621;
  wire v23fbcae;
  wire v2303634;
  wire v23111c7;
  wire v22f015d;
  wire v22fbeb3;
  wire v231262f;
  wire v22fd827;
  wire v23015c7;
  wire v23109c8;
  wire v23fc1db;
  wire v22f8e08;
  wire v23fbfba;
  wire v22fc9cb;
  wire v2310f5b;
  wire v23fa1ad;
  wire v2312bd9;
  wire v23fb60e;
  wire v22f7273;
  wire v22f03b1;
  wire v230aa63;
  wire v23fab26;
  wire v22f98ad;
  wire v230ed8b;
  wire v22f389b;
  wire v22ef2b4;
  wire v22efa0f;
  wire v22fd2e8;
  wire v2303f7c;
  wire bd7a62;
  wire v22f118e;
  wire v22f07d5;
  wire v2309440;
  wire v9df685;
  wire v23fcf56;
  wire v22f5d0e;
  wire v23f426b;
  wire v23fb1b7;
  wire v22fc73a;
  wire v8ef087;
  wire v23f7d2e;
  wire v23fb61d;
  wire v23019b7;
  wire v23f4dc4;
  wire v23f8324;
  wire v23fb73e;
  wire v2303982;
  wire v23fb242;
  wire v230499e;
  wire v22efa95;
  wire v230ea78;
  wire v22ef78e;
  wire v22fc964;
  wire v9ed9e1;
  wire v22f1e6a;
  wire v23fc52e;
  wire v2311b96;
  wire v23fbf9a;
  wire v22ef292;
  wire v22ec1fc;
  wire v23f55c5;
  wire v23117d2;
  wire v23f592f;
  wire v23fbd50;
  wire v23fb6b9;
  wire v22f6db5;
  wire v22fbbcc;
  wire v2305339;
  wire v23f6013;
  wire v106aead;
  wire v23fb752;
  wire v22ec753;
  wire v23026f7;
  wire v230899e;
  wire v921155;
  wire v23f67dd;
  wire v23f8e1f;
  wire b00ad3;
  wire v22fbadb;
  wire v23fce22;
  wire v23f85d7;
  wire v22f7ad6;
  wire v23fc5cd;
  wire v23fca9c;
  wire v230ac33;
  wire v2391d17;
  wire v23fc4d1;
  wire d7df7e;
  wire v2309c45;
  wire v23010ae;
  wire v23f7c65;
  wire v2310c1a;
  wire v23f8e52;
  wire v23fcf49;
  wire v23f9dd1;
  wire v22ff9d4;
  wire v2301ad7;
  wire v2307a6d;
  wire v22ed7ba;
  wire v23fc04f;
  wire v23f5cd3;
  wire v2393abe;
  wire v2305e00;
  wire v2311e38;
  wire v22f9f68;
  wire v2304764;
  wire v23060eb;
  wire v23fc9b6;
  wire v23f34d5;
  wire v23fc33e;
  wire v230381a;
  wire v23fcaf8;
  wire v23fca35;
  wire v23fc15d;
  wire v22f7752;
  wire v23f3ccf;
  wire v23fc838;
  wire v230cb9a;
  wire v22ff3d1;
  wire v23064e4;
  wire v23f4c57;
  wire v23fbc78;
  wire v230ba85;
  wire v12cd54c;
  wire v22ed59e;
  wire v22fe573;
  wire v230bb63;
  wire v22ef46e;
  wire v23fcc08;
  wire v23fcc95;
  wire v22f336f;
  wire v22f30be;
  wire v22f8bd0;
  wire v23fca0f;
  wire v23fa71e;
  wire v22ebb51;
  wire v2311358;
  wire v23f626c;
  wire v23fc147;
  wire v23f593e;
  wire v22fae9f;
  wire v22fa8d7;
  wire v2301edd;
  wire v23fcb65;
  wire v23fc804;
  wire v23fc8b3;
  wire v23fbedc;
  wire v23fbd5d;
  wire v23f849c;
  wire v22ff043;
  wire v2300f25;
  wire v2305483;
  wire v22f484b;
  wire v230180d;
  wire v23f729b;
  wire v23f0206;
  wire v22f9a8b;
  wire v23f6710;
  wire v230ab7a;
  wire v23f9812;
  wire v2307403;
  wire v23f841d;
  wire v230ef1c;
  wire v23f0865;
  wire v23119a8;
  wire v22fd48a;
  wire v23efd4b;
  wire v9b1253;
  wire v23fc678;
  wire v2310d1e;
  wire v2305630;
  wire v22fd60f;
  wire v23fbd8e;
  wire v23fb1d7;
  wire v845651;
  wire v23fc9a4;
  wire v23000a8;
  wire v23fbc7b;
  wire v1e841b6;
  wire bbc337;
  wire v23fb0c2;
  wire v13afb18;
  wire v23fbca4;
  wire a8d315;
  wire v22f926d;
  wire v22ebce1;
  wire v23f820a;
  wire v23f98f8;
  wire v23fc0c9;
  wire v23fcd8d;
  wire v23fd037;
  wire v23f3bd2;
  wire v845637;
  wire v230a3c9;
  wire v845636;
  wire v23fcea8;
  wire v23fc98a;
  wire v22f4114;
  wire bd8af4;
  wire v22ee6ce;
  wire v230a555;
  wire v2302177;
  wire v22fc398;
  wire v230e9f8;
  wire v23f946b;
  wire v2304578;
  wire v23fa36c;
  wire v23fb935;
  wire v23fa1e7;
  wire v22f09a2;
  wire v23fbff3;
  wire v22f2718;
  wire v2311255;
  wire v23efbfd;
  wire v22ee918;
  wire v22f5ab0;
  wire v23f53a0;
  wire v23f26fc;
  wire v22ef39f;
  wire v22f1d6c;
  wire v1aae087;
  wire v22f1389;
  wire v2302048;
  wire v23f9c5f;
  wire v23fc001;
  wire v22f1f78;
  wire v23fbd38;
  wire v2307578;
  wire v230e860;
  wire v22ec8d7;
  wire v22ebbab;
  wire v23076e7;
  wire b15ae7;
  wire v23fc7c0;
  wire v84562f;
  wire v23fbad4;
  wire v23fc346;
  wire v2312dd2;
  wire v23f3d02;
  wire v23068a9;
  wire v22ec6e5;
  wire v22f5198;
  wire v22ef7a5;
  wire v2301135;
  wire v22ff1b9;
  wire v1aadb8e;
  wire v23f35ff;
  wire v230ab2e;
  wire v23f82b3;
  wire v22fcf04;
  wire v230e45a;
  wire v22f961e;
  wire v22f2ca2;
  wire v2308ef0;
  wire v22fd8a4;
  wire v22f9833;
  wire v23f7c32;
  wire v230f0d2;
  wire v2309a8c;
  wire v23f649a;
  wire v23113a4;
  wire v22fce73;
  wire v23fc176;
  wire v23059ee;
  wire v22fd9f5;
  wire v22f5218;
  wire v230af06;
  wire v23fd015;
  wire v87d737;
  wire v23f4d54;
  wire v23f3ca5;
  wire v23fc7db;
  wire v22ec2a4;
  wire v22ed942;
  wire v230fc36;
  wire da3103;
  wire v23090a6;
  wire v22f99e0;
  wire v230e322;
  wire v23fbd64;
  wire v23fbdb1;
  wire v23fcb9d;
  wire v23fc826;
  wire v2309e7a;
  wire v22ee281;
  wire v8f530a;
  wire v23fbdb9;
  wire v230b236;
  wire v2392e6c;
  wire v230158f;
  wire v23fcf96;
  wire v2309e9d;
  wire v13aff51;
  wire v23f0234;
  wire v22fb442;
  wire v2306728;
  wire v22ff982;
  wire v2304dc2;
  wire v23f34b8;
  wire v230f5a4;
  wire v23f5a68;
  wire v2305b34;
  wire v106af3a;
  wire v2308706;
  wire v23efce3;
  wire v23f1c9b;
  wire v23fbd8a;
  wire v23fc5b3;
  wire v22fdad1;
  wire v23fb948;
  wire v23f029a;
  wire v23f2298;
  wire v23fc01d;
  wire v2305aa7;
  wire v23f9737;
  wire v22fac35;
  wire v23fb52f;
  wire v23f2df5;
  wire v23fcd47;
  wire v2312a98;
  wire v22f0a76;
  wire v23fb578;
  wire v23f7680;
  wire v2308b14;
  wire v23078cb;
  wire v23f3d0e;
  wire v230fdf7;
  wire v2391c55;
  wire v22f6c01;
  wire v22fb74f;
  wire v23fbbef;
  wire v23fbbaa;
  wire v23fc49c;
  wire v22ee3c9;
  wire v23f7ad1;
  wire v23f39f2;
  wire v23fb51a;
  wire v23f965d;
  wire v22ed145;
  wire v22ff134;
  wire v22f755a;
  wire v23fc9cf;
  wire v23fbca2;
  wire v23fc24c;
  wire v2307add;
  wire v22f4ba1;
  wire v22f8c84;
  wire v230cc12;
  wire v869055;
  wire v2300d6c;
  wire v23fceb9;
  wire v2309945;
  wire v22f88aa;
  wire v1aad5ad;
  wire v23087d7;
  wire v22fafaa;
  wire v2307750;
  wire v2312775;
  wire v2303e4f;
  wire v22f4d77;
  wire v23fcea0;
  wire v84562b;
  wire a8b64b;
  wire v230a6a7;
  wire v23fbab2;
  wire v12cd4c6;
  wire v23fb5b4;
  wire v22fd696;
  wire v230e43d;
  wire v22ffdd1;
  wire v22eb338;
  wire v922c74;
  wire v2308b24;
  wire v22fa976;
  wire v22eaeab;
  wire v2302868;
  wire v23fb562;
  wire v17a34f9;
  wire v23fbe83;
  wire v23fc746;
  wire v230abf6;
  wire v23fbc65;
  wire v23fb9e5;
  wire v15072a7;
  wire v230f151;
  wire v23fca45;
  wire v23059c5;
  wire v23f7014;
  wire v23fcd56;
  wire v2301a75;
  wire v8a3511;
  wire v22ef062;
  wire v94e407;
  wire v23fbfe5;
  wire v23fc143;
  wire v22f5e91;
  wire v23f62a8;
  wire v23f0288;
  wire v23fcf94;
  wire v23fb2f5;
  wire v22f1585;
  wire v23fc6d3;
  wire v23065b6;
  wire v2308765;
  wire v2308331;
  wire v2305bb2;
  wire v230c8e9;
  wire v23030ad;
  wire v23fbdfd;
  wire v23f85b0;
  wire v230665f;
  wire v845627;
  wire v23070c0;
  wire v2310bf5;
  wire v22f2095;
  wire v22ff18a;
  wire v23f6326;
  wire v22f1faf;
  wire v23fb8e4;
  wire v23fcfa6;
  wire v22f7ef7;
  wire v23fbde1;
  wire v2309a1d;
  wire v23fcdda;
  wire v23f79d2;
  wire v23f44bd;
  wire v23fc630;
  wire v23f06a5;
  wire v23fb71a;
  wire v2367a45;
  wire v23fb22d;
  wire v23049d7;
  wire b50a75;
  wire v22f5fb4;
  wire v22ee124;
  wire v23fba25;
  wire v23f471a;
  wire v22f21bd;
  wire v22ff4af;
  wire v22fa3fa;
  wire v22fff2d;
  wire v23fb819;
  wire v23f111f;
  wire v22fc42e;
  wire v22ef810;
  wire v23f91a5;
  wire v22f16ef;
  wire v230038a;
  wire v23096f8;
  wire v23fb590;
  wire v2301509;
  wire v22ff1dd;
  wire v22ec2c4;
  wire v23fc29d;
  wire v23fcc6c;
  wire v22eb60c;
  wire v22ebd1b;
  wire v22eafaa;
  wire v22f07bb;
  wire v230fb9e;
  wire v23f96b0;
  wire a1fbcb;
  wire v23fa903;
  wire v23fc92e;
  wire v9cf5cf;
  wire v12cda11;
  wire v22ef079;
  wire v22ff80d;
  wire v23fb544;
  wire bfce54;
  wire v22fc90f;
  wire v22eaf73;
  wire v22f5941;
  wire v22f9160;
  wire v23f2bc0;
  wire v23f5046;
  wire v9442ad;
  wire v23fa215;
  wire v23f2d39;
  wire v230aedf;
  wire v23fc80c;
  wire v23f5cd7;
  wire v22ed35b;
  wire v22f3a1f;
  wire v845633;
  wire v191acb4;
  wire v23f07eb;
  wire v22fad67;
  wire v230ba49;
  wire v230184a;
  wire v22f4ecf;
  wire v2306cca;
  wire v22f7fc1;
  wire v22f6f2d;
  wire v23fbc46;
  wire v23fbd51;
  wire v23fbb35;
  wire v22fc8e5;
  wire v23fba70;
  wire v23f5be9;
  wire v22ee946;
  wire v22f49c4;
  wire v23f54ef;
  wire v23fc493;
  wire v22efb8c;
  wire v2301274;
  wire v845623;
  wire v22ffcbd;
  wire v845622;
  wire v22f878c;
  wire e1e72e;
  wire v23fbf36;
  wire fc8f90;
  wire v1aad354;
  wire v22f511c;
  wire v23f35a8;
  wire v22eedbb;
  wire v230f0c6;
  wire v150716b;
  wire v23017a9;
  wire v23faa11;
  wire v23fc917;
  wire v230efa0;
  wire v230089c;
  wire v2309c79;
  wire v23fcbf0;
  wire v23f5240;
  wire v23fb77d;
  wire v22eb651;
  wire v23051a9;
  wire e1e75d;
  wire v23f1c0b;
  wire v23fba66;
  wire v230c213;
  wire v23f4096;
  wire v22fe9e0;
  wire v2304ec7;
  wire v22f0fb9;
  wire v23f7698;
  wire v23021af;
  wire v23fce1e;
  wire v22f004e;
  wire v22f05f3;
  wire v23133fa;
  wire v22ec658;
  wire v22f2f87;
  wire v22f446e;
  wire v23fcedd;
  wire v2307788;
  wire v230f347;
  wire a476c2;
  wire v23fc9d2;
  wire v2312351;
  wire v23fc38f;
  wire d79b38;
  wire a1fbe9;
  wire v23f06ee;
  wire v23fc457;
  wire v2310ad7;
  wire v23fc669;
  wire v2307805;
  wire v23fbbc7;
  wire v23fc842;
  wire v23efe0a;
  wire v191ae6e;
  wire v22ef5c2;
  wire v23f5abd;
  wire v23f8689;
  wire v23fcc84;
  wire v22f09b1;
  wire v22f2965;
  wire v22eec14;
  wire v12cc317;
  wire v23095d8;
  wire v23fc12b;
  wire v22f3000;
  wire v22f85a0;
  wire v2310a9f;
  wire v23fc13a;
  wire v230bbb3;
  wire v22f9089;
  wire v23fc30d;
  wire v231398c;
  wire v23110b9;
  wire v22ff106;
  wire v230b089;
  wire v23063f8;
  wire v2303679;
  wire v22f39d3;
  wire v230efe0;
  wire v23f6532;
  wire v23f1f36;
  wire bee61a;
  wire v23004ba;
  wire v12cd540;
  wire c08bce;
  wire v2300070;
  wire v22ec763;
  wire v22eb6c8;
  wire v22fa23d;
  wire v230a15d;
  wire v2302943;
  wire v23fce29;
  wire v22ecf16;
  wire v22fcef4;
  wire v23f2dbb;
  wire v23fb8b7;
  wire v22fdbac;
  wire v23f23f4;
  wire v22f2009;
  wire v22f954a;
  wire v22fc92d;
  wire v22ed1b0;
  wire v23fb1bb;
  wire v23fb0a8;
  wire v230aa5d;
  wire v2312d9c;
  wire v230dcd9;
  wire v231243e;
  wire v23f9758;
  wire v2300c56;
  wire v2392f02;
  wire v23fc08e;
  wire v23fcf44;
  wire v22f7e19;
  wire bf7e60;
  wire v13afb04;
  wire v22f7b49;
  wire v23f46d8;
  wire v23fc68e;
  wire v22eb57a;
  wire v23916d5;
  wire v22ebb8e;
  wire v12cd552;
  wire v2307bcb;
  wire v2312ea4;
  wire v23121e0;
  wire v23fc4b0;
  wire v2310bf7;
  wire v22fccc4;
  wire ab2d7c;
  wire v22f8834;
  wire v23fc633;
  wire v22eda0b;
  wire v22ef026;
  wire v22ed01d;
  wire v23fcdf0;
  wire v22fa49d;
  wire v23fc0a3;
  wire v2303b0a;
  wire v22eb6e4;
  wire v23fc2da;
  wire v22f90d2;
  wire v230420d;
  wire v23f1495;
  wire v22f63e9;
  wire v230f069;
  wire v2307fee;
  wire v2308237;
  wire a3aa64;
  wire v23fc4e7;
  wire fc894d;
  wire v23f6fe7;
  wire v230af39;
  wire v22f1dec;
  wire v23f443c;
  wire v22fa631;
  wire v23f748c;
  wire v22ff789;
  wire v23f8dba;
  wire v22fb7e2;
  wire v23f2849;
  wire v2307de6;
  wire v23fcdfa;
  wire v230c81f;
  wire v106a7cd;
  wire v2308be7;
  wire v23fcbaa;
  wire v23fba1d;
  wire v22eec56;
  wire v22f08f1;
  wire v2309d59;
  wire v23fb4ae;
  wire v22f7ceb;
  wire v230c025;
  wire v23fc1c6;
  wire v2311cd1;
  wire v2304bc1;
  wire v230e869;
  wire v230aa99;
  wire v12cda15;
  wire v22f6b45;
  wire v2300d1d;
  wire v22eb32b;
  wire v23f3940;
  wire v23fb8a2;
  wire v2312d20;
  wire v23f5ce0;
  wire v230580d;
  wire v22f3aa1;
  wire v22f0538;
  wire v23925a8;
  wire v2309e57;
  wire v230f14b;
  wire v23fcd16;
  wire v23fbc5a;
  wire v23fcef5;
  wire v23059b0;
  wire v23fcdc1;
  wire v22f4ee6;
  wire v23fbe05;
  wire v22fc95b;
  wire v23fce8e;
  wire v23fcb2d;
  wire v230e28d;
  wire v23fca75;
  wire v230e40a;
  wire v23064ae;
  wire v22f4d68;
  wire v239302b;
  wire v22f7e37;
  wire v22ef424;
  wire v2307a5e;
  wire v2302bd3;
  wire v23f2abe;
  wire v2300d32;
  wire v23fc3fb;
  wire v22ecbbd;
  wire v2393321;
  wire v2312925;
  wire v22ef1eb;
  wire v22f2450;
  wire v23f120d;
  wire v23f4979;
  wire v22ece0d;
  wire v22f92f8;
  wire v230ae06;
  wire v22eeb19;
  wire v22ed8fe;
  wire v23f18da;
  wire v22ebed1;
  wire v23f3561;
  wire v23f81e6;
  wire v2310406;
  wire v191ac40;
  wire v23060ff;
  wire v230894d;
  wire v23f6ec1;
  wire v23fcbb6;
  wire v22ebe03;
  wire v22fa86d;
  wire v22fc903;
  wire v230db4d;
  wire v22fdabc;
  wire v23f1cd2;
  wire v22eec0e;
  wire v2308d5a;
  wire v23fbc3a;
  wire v22f9dab;
  wire v22f78c3;
  wire v23065fc;
  wire v22f23f6;
  wire v22f6090;
  wire v23f7796;
  wire v23108a7;
  wire v23fc957;
  wire v231022d;
  wire v23fc6a0;
  wire v2305296;
  wire v23f2d37;
  wire v2310eb0;
  wire v2393f08;
  wire v2300881;
  wire v22fb5a3;
  wire v23f883a;
  wire v230af38;
  wire v22fa5f9;
  wire v2305d89;
  wire v23fc587;
  wire v22f752e;
  wire v13afef6;
  wire v22ffdc3;
  wire v23f96d1;
  wire v22ee50f;
  wire v23fca5d;
  wire v22f4407;
  wire v85bd38;
  wire v230aef9;
  wire v23fcbde;
  wire v13aff5b;
  wire v23059d8;
  wire v2306785;
  wire v2394081;
  wire v22fd79e;
  wire d49f20;
  wire v191aea6;
  wire v2303535;
  wire v22fb4a1;
  wire v2310558;
  wire v23fc1bf;
  wire v22eb742;
  wire v23fbb5f;
  wire v230e618;
  wire v23fba07;
  wire v22f9b00;
  wire v23fbc75;
  wire v2305e86;
  wire v2308ee1;
  wire v23916d6;
  wire v23faacf;
  wire v23fb477;
  wire v23003a8;
  wire v23fc53e;
  wire v230e78c;
  wire v23ef8ef;
  wire v2306257;
  wire v9347cd;
  wire v895ae7;
  wire v22fd663;
  wire v22f3092;
  wire v23f6d92;
  wire v22f6265;
  wire bd74ba;
  wire v23f99cf;
  wire v2392c41;
  wire v2303f37;
  wire v23127fb;
  wire v2300a5a;
  wire v23f4ccb;
  wire v23f7a5f;
  wire v22edb0c;
  wire v22fc05f;
  wire b5e598;
  wire v23fba35;
  wire v22f17eb;
  wire v230f253;
  wire v23fb648;
  wire v23f3adc;
  wire v22eb72a;
  wire f40dab;
  wire v995fa2;
  wire v1e8471c;
  wire v23f832b;
  wire v22ef65b;
  wire v2310253;
  wire v2305cf5;
  wire v230e040;
  wire v230105d;
  wire v2301bcb;
  wire v23fa0a3;
  wire v23f240a;
  wire v22ebf17;
  wire v906d1d;
  wire v2312a8d;
  wire v23fb942;
  wire v2301f52;
  wire a1382d;
  wire v23fc974;
  wire v230fa92;
  wire v2306441;
  wire v22f0d8d;
  wire v230b78b;
  wire v23fbcef;
  wire v23f5d7f;
  wire v23fc303;
  wire v23f8979;
  wire v22f1992;
  wire v230bc0c;
  wire v230bb30;
  wire v22eaa94;
  wire v23fa9c5;
  wire v23035d7;
  wire v23f004a;
  wire v23fce4e;
  wire v22fb2c5;
  wire v230bdb9;
  wire v23fb9d6;
  wire v2304c86;
  wire v12cd534;
  wire v22edf79;
  wire v23fb7da;
  wire v191b212;
  wire v22fb081;
  wire v23fb958;
  wire v22f2ac8;
  wire v86374c;
  wire v23032db;
  wire v22f8b55;
  wire v22fd6f9;
  wire v230e872;
  wire v23fc064;
  wire v230b4af;
  wire v22ff8a6;
  wire v23fc828;
  wire v23f1f6f;
  wire v23f340b;
  wire v22fa654;
  wire v23f7d51;
  wire v2304415;
  wire v13affe0;
  wire v106ae69;
  wire v23f79a9;
  wire v22f8e10;
  wire v230df30;
  wire v23f8093;
  wire v23fac04;
  wire v2307dbf;
  wire v23fb80a;
  wire v23fb0cd;
  wire v23fca23;
  wire v22edf81;
  wire v2309263;
  wire v12cd9cd;
  wire v22f1e02;
  wire v2305792;
  wire v230abb1;
  wire v2305838;
  wire v23fb6a6;
  wire v230e1a3;
  wire v2307779;
  wire v22ff916;
  wire v23f5fa6;
  wire v230d134;
  wire v23fb1a1;
  wire v22faae8;
  wire v23f5c89;
  wire v22ffea8;
  wire v230840f;
  wire v239174c;
  wire v22f6ad2;
  wire v2392bc1;
  wire v2306c80;
  wire v23f15ec;
  wire v23fd045;
  wire v230a8ea;
  wire v231114e;
  wire v23fc4fd;
  wire v23fce98;
  wire v23fbcfc;
  wire v23f5d6f;
  wire v2303ee8;
  wire v230875c;
  wire v150736d;
  wire v23f0d46;
  wire v23fc03c;
  wire v23fce7b;
  wire v22f4a20;
  wire v2306de4;
  wire v230a891;
  wire v1aad4ef;
  wire v22f4089;
  wire v2304924;
  wire v23fcc58;
  wire v22f9e59;
  wire v23f53d0;
  wire e1e1ba;
  wire v23040a5;
  wire v230267d;
  wire v23f717f;
  wire v230a05f;
  wire v22f067b;
  wire v23115bd;
  wire v23133b3;
  wire v230d75a;
  wire f40d66;
  wire c16218;
  wire v22efc21;
  wire v23f9452;
  wire v23f35c7;
  wire v22fe2d5;
  wire v2312a52;
  wire v23fb1db;
  wire v23f3d0b;
  wire v2300142;
  wire v22f8d58;
  wire v22ee057;
  wire v230197f;
  wire v22f7371;
  wire v23fbe03;
  wire v23f957b;
  wire v23f5eba;
  wire v23f2704;
  wire v2393f1a;
  wire v23f200c;
  wire v23fbfee;
  wire v23936a3;
  wire v2307704;
  wire v230bead;
  wire v23102b0;
  wire v23f2b21;
  wire v23f2d1d;
  wire v23fbb98;
  wire v23f20d0;
  wire v23fc60a;
  wire v22f6cde;
  wire v231330b;
  wire v23fc846;
  wire v2310197;
  wire v23fb6b6;
  wire v22fa889;
  wire v22ee8bf;
  wire v23fc51e;
  wire v2303513;
  wire v2309889;
  wire v22eb01f;
  wire v22fd71a;
  wire v1e84195;
  wire a0de1c;
  wire v22f1117;
  wire v22fc27d;
  wire v23f942a;
  wire v230562d;
  wire v23f8100;
  wire v23fc459;
  wire v22fa646;
  wire v22f9ab6;
  wire v23faf72;
  wire v23f5983;
  wire v23fc030;
  wire v22ed925;
  wire v2302c6d;
  wire v191b10f;
  wire v23fcb8a;
  wire v2305aea;
  wire v12cde1b;
  wire v23fc1b3;
  wire v23008a6;
  wire v23fc9b7;
  wire be86f6;
  wire v22fa064;
  wire v23fcf8a;
  wire v22fe408;
  wire v230f072;
  wire v22f7098;
  wire v23fc3c2;
  wire v23f47a1;
  wire v23fbcd2;
  wire v22ff4bc;
  wire v22f5136;
  wire v23127ee;
  wire v230064b;
  wire v2303c5a;
  wire v23fb62d;
  wire v2304048;
  wire v23fc9b4;
  wire v22f2487;
  wire v2311f82;
  wire v23fa966;
  wire v903f7f;
  wire v23fc443;
  wire v23fc7e5;
  wire v22eefab;
  wire v22ebe99;
  wire v230a573;
  wire v23025ae;
  wire v23fcab6;
  wire v22f7859;
  wire v23f794b;
  wire v230e07d;
  wire v2310a7e;
  wire v230e311;
  wire v2309aa0;
  wire v23fbe81;
  wire bc5d21;
  wire v23f9c45;
  wire v23fc153;
  wire v230a42d;
  wire v22efa49;
  wire v9ec6b5;
  wire v1aadac4;
  wire v22ef750;
  wire v2311524;
  wire v22fe62a;
  wire v22f971b;
  wire v230e8a0;
  wire b72216;
  wire v23028be;
  wire v22f3cf2;
  wire v23fca50;
  wire v22f3d5a;
  wire v23fb97f;
  wire v23fc7ff;
  wire v2393f0d;
  wire v2308e98;
  wire v23fd06a;
  wire v23fcf98;
  wire v22fd6d8;
  wire v22f71ca;
  wire v2308bcd;
  wire v22fd124;
  wire v23fbda1;
  wire v23fb172;
  wire v23fcadd;
  wire v23fab8b;
  wire v23005e2;
  wire v22f3a6f;
  wire v22f7a0c;
  wire v23fcc22;
  wire v23fba03;
  wire v22f2319;
  wire v22f0218;
  wire v23fbf35;
  wire v22eef44;
  wire v23fca38;
  wire v23f0a6b;
  wire v23fcbc9;
  wire v960676;
  wire v23fbfca;
  wire v2393de1;
  wire v23f7950;
  wire v230201b;
  wire a03e3a;
  wire bd74c6;
  wire v230630c;
  wire v22f6397;
  wire v22f5fa1;
  wire v230b95f;
  wire v22f7efd;
  wire v22f7466;
  wire v23fbae8;
  wire v23fb1ab;
  wire v22f65b7;
  wire e1e250;
  wire v239228f;
  wire v23fb931;
  wire v230c104;
  wire v22fe0f9;
  wire v239254b;
  wire v23fc849;
  wire v22f65c0;
  wire v22ec1c3;
  wire v23fce4c;
  wire v23f5cfe;
  wire v22fd0fa;
  wire v23fcf9e;
  wire v22f10d6;
  wire v22f56c2;
  wire v230bdd9;
  wire v23fab9b;
  wire v22facd1;
  wire v23f6d80;
  wire v22f1e91;
  wire v230bbce;
  wire v12cd3aa;
  wire v23f4194;
  wire v22f063d;
  wire v23fcd03;
  wire v22ecaf6;
  wire v22f34bd;
  wire v22f516b;
  wire v230c428;
  wire v23f9f68;
  wire v22facbb;
  wire v230cb7a;
  wire v23f8970;
  wire v230bb21;
  wire v23fc203;
  wire bd7adc;
  wire v23f77b1;
  wire v23f0d8a;
  wire v23fc5c6;
  wire v2392fa6;
  wire v22f5120;
  wire v23fcc97;
  wire v22ef481;
  wire v23fb11b;
  wire v191b107;
  wire v23fb7b4;
  wire v230a65d;
  wire v23fb043;
  wire v23fc72c;
  wire v23f1a86;
  wire bdeff3;
  wire v23f507b;
  wire v2312164;
  wire v23fc79a;
  wire v22fbf21;
  wire a04d83;
  wire v22f7a1d;
  wire v2307206;
  wire v23f561c;
  wire v23fc937;
  wire v22f7277;
  wire v23f8a43;
  wire v23fbd2a;
  wire v23f74bf;
  wire v2392f25;
  wire v2302844;
  wire v23f4b9c;
  wire v23fc065;
  wire v22eddae;
  wire v22f36c5;
  wire v23f40d1;
  wire v22ec334;
  wire v23fcdb4;
  wire v23f44d0;
  wire v2312ac8;
  wire v23f77c5;
  wire v23f350b;
  wire v22ecdde;
  wire v23fca5c;
  wire v22ebf32;
  wire v23f15c1;
  wire abc0f5;
  wire v23f8124;
  wire v22fa5a6;
  wire e1e6ee;
  wire v22f5afa;
  wire v23fb145;
  wire v2307d93;
  wire v191b1ae;
  wire v23f35de;
  wire v22f1efd;
  wire v22f8acc;
  wire v22ed654;
  wire v23f7cbe;
  wire v22fa6ae;
  wire v22f9601;
  wire v2309c93;
  wire v2310589;
  wire v2305c7f;
  wire v23074d2;
  wire v23fbf16;
  wire v23f99ae;
  wire v23fc390;
  wire v2311027;
  wire v22f7ccb;
  wire v23f7b9e;
  wire v23f2041;
  wire c16602;
  wire v22fab2d;
  wire v230564d;
  wire v15075f0;
  wire v22f4eeb;
  wire v22f48a5;
  wire v2305071;
  wire v22ebfd7;
  wire v23fbd58;
  wire v2305d6e;
  wire v23fbae6;
  wire v2300ccc;
  wire v22efdae;
  wire v23fc1bc;
  wire v2307224;
  wire v23fc80d;
  wire v23f1643;
  wire v22ece6c;
  wire v23fc726;
  wire v23fc17b;
  wire v1aad571;
  wire v23f859a;
  wire v230b09e;
  wire v17a34ea;
  wire v23f9226;
  wire v23fba7c;
  wire v23fbb41;
  wire v230cb59;
  wire v23f111c;
  wire v23fb9a9;
  wire v23f50bd;
  wire v23f543d;
  wire v230b131;
  wire v22ed4b7;
  wire v2308d20;
  wire v23fc335;
  wire v230259f;
  wire v230c116;
  wire v23fb788;
  wire v23f7f0d;
  wire v230590b;
  wire v22f1899;
  wire v23fb592;
  wire v23fcba2;
  wire e1dbd6;
  wire v22f6e30;
  wire v8963c2;
  wire v23f5fc3;
  wire v23f5398;
  wire v22f5f28;
  wire v22f8894;
  wire v23f1032;
  wire v22faa4d;
  wire v23fb095;
  wire fc8f81;
  wire v231196d;
  wire v22f5f09;
  wire v23fc796;
  wire v23919bb;
  wire v1507529;
  wire da38ba;
  wire v22f36da;
  wire v23f58e1;
  wire v23056bf;
  wire v2392537;
  wire v22fe382;
  wire v23fb6c7;
  wire v23fb33a;
  wire v22f910f;
  wire v23131af;
  wire da310f;
  wire v22eedcd;
  wire v2302244;
  wire v239299c;
  wire v22f5f54;
  wire v23fcfd3;
  wire v23f8345;
  wire v23fb84a;
  wire v2301f9a;
  wire v23f84cc;
  wire v23f4f34;
  wire v2304443;
  wire v230d9cf;
  wire v230dd35;
  wire v2300d0f;
  wire v22fb379;
  wire v2303ba8;
  wire v23fb919;
  wire v8cded5;
  wire v23f5102;
  wire v23126de;
  wire v23030fc;
  wire v22efa93;
  wire v23f4cfb;
  wire v23fbf61;
  wire da310c;
  wire v22f575a;
  wire v22f42a5;
  wire v23f37c8;
  wire fc8fdb;
  wire v230e2bb;
  wire v230b4b4;
  wire v22fed4f;
  wire v23fb492;
  wire v23f56c3;
  wire v191a964;
  wire v23fced0;
  wire v23fcb87;
  wire v2301178;
  wire v22f4d20;
  wire v23934f3;
  wire v22f0050;
  wire v2312680;
  wire v23f56bc;
  wire v230a84b;
  wire v23fc2ae;
  wire v2309d7f;
  wire v23fbbc2;
  wire v2310682;
  wire v23f924a;
  wire v23139c3;
  wire v22eb952;
  wire v230629d;
  wire v23129c2;
  wire v22ef9ea;
  wire v23fc57c;
  wire v23fb947;
  wire v22f6fda;
  wire v23fbd5b;
  wire v22f76b3;
  wire v23fc4a2;
  wire v23119b0;
  wire a452a3;
  wire v23f215c;
  wire v23934b5;
  wire v23fb66d;
  wire v23f7714;
  wire v94f831;
  wire v22fa309;
  wire v2306838;
  wire v22f2590;
  wire v2391950;
  wire v868c84;
  wire v230118f;
  wire v22f3189;
  wire v22f8309;
  wire v23fb9c5;
  wire v22ecd97;
  wire v8f2065;
  wire v23fc513;
  wire v23f5ce2;
  wire v230b59f;
  wire v23f1a43;
  wire v23f087f;
  wire v23f8a0e;
  wire v2313059;
  wire v230a63b;
  wire v2391bb7;
  wire v230b8cd;
  wire v8bb259;
  wire v22ff890;
  wire v23fbe09;
  wire v230f537;
  wire v22f8093;
  wire v23fcb64;
  wire v23fbf12;
  wire v2308af4;
  wire v23f4ab8;
  wire v23139aa;
  wire v230ae19;
  wire v22ecec6;
  wire v22ff4c3;
  wire v230e6ea;
  wire v22f9452;
  wire v22edadc;
  wire v22ebc60;
  wire v2303e0d;
  wire v2312053;
  wire bd9dce;
  wire v22f536a;
  wire v22f3738;
  wire v22fc122;
  wire v23fc2ee;
  wire v22f8acf;
  wire v22fb5f7;
  wire b16326;
  wire v22f7dc7;
  wire v230156d;
  wire v23fc73e;
  wire v23fc686;
  wire v23fc19c;
  wire v23fc99f;
  wire v230ae1e;
  wire v230c233;
  wire v2346b6a;
  wire v230fc70;
  wire v22fadb0;
  wire v22f2639;
  wire v23fc7f5;
  wire v230bbe4;
  wire v23fcf79;
  wire v22efd62;
  wire v22fdd09;
  wire v22f4678;
  wire v22ee457;
  wire v1506ae6;
  wire v23f50bb;
  wire b10190;
  wire v230b19a;
  wire v23f3e42;
  wire v23f5461;
  wire v23f6d50;
  wire v22f2bb8;
  wire v1aae175;
  wire v2312187;
  wire v2310a9a;
  wire v23f6309;
  wire v23f7275;
  wire v23fba0c;
  wire v2305628;
  wire v23f5ed5;
  wire v22f18b1;
  wire v23fbd3e;
  wire v22ecced;
  wire v230ecac;
  wire v2393346;
  wire v230361d;
  wire v22f2d35;
  wire v230f790;
  wire v23fc013;
  wire v23f7b94;
  wire v23f96b7;
  wire v23f1f1e;
  wire v23fc947;
  wire v230037d;
  wire v22f4700;
  wire v230828c;
  wire fc8c57;
  wire v12cda32;
  wire v23fcf2d;
  wire v22efa67;
  wire v23f00ec;
  wire v23fbda4;
  wire v23f68c1;
  wire v23f2b6d;
  wire v22ec9ce;
  wire v2301e66;
  wire v23f79a7;
  wire v23f7637;
  wire v23fcc0c;
  wire v22f988a;
  wire v22f679a;
  wire v23fb9e7;
  wire v22ff66a;
  wire v230b0c6;
  wire v2302f2c;
  wire v23fa1e3;
  wire v23f9044;
  wire v22eb303;
  wire v23fbaac;
  wire v230a2c7;
  wire v23fcd49;
  wire v23fc783;
  wire v23132fc;
  wire v23020a2;
  wire v2305b2e;
  wire v2311c16;
  wire v230c499;
  wire v22ec0f7;
  wire a7fdb1;
  wire v23f8d5a;
  wire bcc479;
  wire v23f4168;
  wire v230ad0e;
  wire v2302dc1;
  wire v22f1cc5;
  wire v23fb166;
  wire v22faa4b;
  wire v23f36d3;
  wire v22ebfcf;
  wire v22f091e;
  wire v1aae362;
  wire v22fa4b4;
  wire v2300b96;
  wire v23fc40f;
  wire v23fb798;
  wire v23fa7ec;
  wire v23fcaf0;
  wire v22fa6a4;
  wire v23fbe12;
  wire v22faba3;
  wire v230f010;
  wire v22fad24;
  wire v22fc508;
  wire v22ed5c8;
  wire v22ed72b;
  wire v23fcaad;
  wire v15071c2;
  wire v23095fa;
  wire v15070e0;
  wire v22ff315;
  wire v2391e51;
  wire v23fbb0f;
  wire v22f2f44;
  wire v23f91e7;
  wire v23fb218;
  wire v230cd61;
  wire v22ffc55;
  wire v230bdd6;
  wire v22efd70;
  wire v2300e95;
  wire v230a4f1;
  wire v12cd538;
  wire v23040c7;
  wire v2393b5a;
  wire v23fa875;
  wire v231051e;
  wire v23010b3;
  wire v23fc753;
  wire v22fbdbc;
  wire v23fcce3;
  wire v23f6038;
  wire v23f368a;
  wire a136c1;
  wire v22f3262;
  wire v22fef6a;
  wire v230128e;
  wire v23fca5a;
  wire v2312aec;
  wire v23f0bd2;
  wire v23017ee;
  wire v22fa101;
  wire v23fc8ee;
  wire v23f34d4;
  wire v23fba09;
  wire v22fe0c1;
  wire v23112d5;
  wire v22f7564;
  wire v230aa0c;
  wire v2311967;
  wire v23fb821;
  wire v23fb99f;
  wire v22ff36f;
  wire v22fa8e6;
  wire a5d081;
  wire v2304583;
  wire v23fcec5;
  wire v191ad2f;
  wire bd74ad;
  wire v22fcf75;
  wire v23115e2;
  wire v23fbe63;
  wire v22f6176;
  wire v23fb673;
  wire v23fc3fe;
  wire v23f16f6;
  wire v2300edd;
  wire v23f2a1a;
  wire v22f4bdf;
  wire v23fc8f0;
  wire v2309099;
  wire d7db8a;
  wire v22f4cf3;
  wire v230cfc7;
  wire v22ee95f;
  wire v22f2eaf;
  wire v22f1ae9;
  wire ab5bb8;
  wire v23f8089;
  wire v2304009;
  wire v23f7024;
  wire v23fbc9a;
  wire v23fca55;
  wire v23f7158;
  wire v23fc529;
  wire v23fcaaa;
  wire v22f8088;
  wire v2311f53;
  wire v22f9a51;
  wire v23066df;
  wire v22fbb8a;
  wire v23118f7;
  wire v23f5fdb;
  wire v2309790;
  wire v23fc9e4;
  wire b9d038;
  wire v22f1d08;
  wire v23f60fb;
  wire v23fc6c2;
  wire v23fca7a;
  wire v22f2fe1;
  wire v22f968e;
  wire v12cd632;
  wire v23fb1aa;
  wire v230f9db;
  wire v23124c5;
  wire v230e02e;
  wire v22fc452;
  wire v230d5a9;
  wire v23133a7;
  wire v1507102;
  wire v23f41c2;
  wire v230c73d;
  wire v22ff6a8;
  wire v22f0de0;
  wire v230ae46;
  wire v2311645;
  wire v2312301;
  wire v23051cf;
  wire v23fbc40;
  wire v22ecc58;
  wire v23fb4d8;
  wire v23faee6;
  wire v23fcf40;
  wire v23fc416;
  wire v23fc6b0;
  wire v2304402;
  wire v23fc4d0;
  wire v23fc5d0;
  wire v230685f;
  wire v22f636a;
  wire v23fb9b2;
  wire e1e73c;
  wire v22fe0ef;
  wire v23f682a;
  wire v23fd025;
  wire v2301c02;
  wire v230eed2;
  wire v23f9507;
  wire a8e3ee;
  wire v22fc53d;
  wire v23f7429;
  wire v22ec0d1;
  wire v2301292;
  wire v2302245;
  wire v23fc2d7;
  wire v23f1279;
  wire v23fc6b6;
  wire v22f7c05;
  wire v23f5526;
  wire v12cc2ef;
  wire v230ae3f;
  wire v23f15a7;
  wire v22fecf3;
  wire v23f3e1b;
  wire v23f515d;
  wire v22f1383;
  wire v22fd83a;
  wire v22fafef;
  wire v13afed6;
  wire v22f023b;
  wire v23fca20;
  wire v23fa5d4;
  wire v22f4eab;
  wire v230eb5a;
  wire v23f1816;
  wire v2311fb5;
  wire v23fbca0;
  wire v230e9ef;
  wire v23fcf17;
  wire v22f061c;
  wire v23fbed7;
  wire fc8f74;
  wire v23f6dc8;
  wire v1aad847;
  wire v22fbdda;
  wire v2308364;
  wire v2301800;
  wire v23119e3;
  wire v23fccf5;
  wire v22f95c3;
  wire v95ca80;
  wire v22efeb6;
  wire v2301992;
  wire v2302c02;
  wire v22f0cf9;
  wire v23fbd28;
  wire v23fd019;
  wire v22ef5f1;
  wire v239157f;
  wire v23fcec4;
  wire v23fb657;
  wire v23fbe38;
  wire v23fc83e;
  wire v23fc006;
  wire v230e7d2;
  wire v22ff89d;
  wire v2303e60;
  wire v23fc658;
  wire v22f2c8b;
  wire v230308e;
  wire v23fc1d2;
  wire v230b125;
  wire v230f70d;
  wire v23f939f;
  wire v23fae9e;
  wire v22efc04;
  wire v22f0546;
  wire v2301c51;
  wire v23f7789;
  wire v23f301a;
  wire v22f4d97;
  wire v22fd387;
  wire v23f9127;
  wire v230547a;
  wire v23f5ace;
  wire v22f383c;
  wire v230694d;
  wire v23f7f51;
  wire v22ee8dd;
  wire v230e703;
  wire v22ed01c;
  wire v22ecd9e;
  wire v2392d0d;
  wire v1506aab;
  wire v22f9793;
  wire v23fb9b9;
  wire v23fce8d;
  wire v2311a1d;
  wire v22eda36;
  wire a1fcc3;
  wire v23fc35a;
  wire v22f83e8;
  wire v23f5a88;
  wire v230536c;
  wire v23f3cb8;
  wire v23f4ed3;
  wire v23fc0e0;
  wire v23fbe27;
  wire v22f4fb8;
  wire v22fc6ca;
  wire v22f2e75;
  wire v22f0f15;
  wire v2304910;
  wire v2302d97;
  wire v23fc5be;
  wire v22edf29;
  wire v230ef38;
  wire v22fd6c8;
  wire v2312d71;
  wire v23037d3;
  wire v22fc2eb;
  wire v23fb576;
  wire v22f96e9;
  wire v230c805;
  wire v230a890;
  wire v22fa857;
  wire v22f53e2;
  wire v230f3e5;
  wire v22f2de3;
  wire v23f692f;
  wire v22fd522;
  wire v22f83fd;
  wire v23fb5d7;
  wire v22eddf2;
  wire v15071f0;
  wire v22fc745;
  wire v23faa16;
  wire v23f8772;
  wire v23f6e45;
  wire v23fc04c;
  wire ae78a6;
  wire v2310104;
  wire v22fc5fd;
  wire v1507317;
  wire v23fc02e;
  wire v2346b79;
  wire v23f917f;
  wire v22ee920;
  wire v23f282d;
  wire v2300936;
  wire v23f6cef;
  wire v22f7e59;
  wire v230ced0;
  wire v230fbc5;
  wire v2300c80;
  wire v22f316b;
  wire v22f6671;
  wire v23fcd70;
  wire v2307b17;
  wire v22fdcc5;
  wire v23fc8a9;
  wire v22f01b2;
  wire v23f7a8e;
  wire e1e35b;
  wire v22f2835;
  wire v22ff6f9;
  wire v2312057;
  wire v230bdd0;
  wire v23001c7;
  wire v23fcb83;
  wire v2306f3c;
  wire v22fa56f;
  wire v23fa4bd;
  wire v22fe2dc;
  wire v22f8ad5;
  wire v23faaa0;
  wire v22f7659;
  wire v23111d5;
  wire v22ef21f;
  wire v2303bc3;
  wire v22ff0be;
  wire v23fc84a;
  wire v230206c;
  wire v230e44a;
  wire v230c95c;
  wire v23fcccb;
  wire v23fc270;
  wire v22f5242;
  wire v230859e;
  wire v22ec63d;
  wire v12cd903;
  wire v22f21f6;
  wire b00a78;
  wire v22f5235;
  wire v23fc9ee;
  wire v23fa66e;
  wire v22f696f;
  wire v12cc310;
  wire v230928c;
  wire v22f0c59;
  wire v22f1963;
  wire v23fc31a;
  wire v23fc511;
  wire v22f971f;
  wire v2303822;
  wire v23fb91d;
  wire v22eff53;
  wire b0fc7a;
  wire v23f613e;
  wire v23fc105;
  wire v2304060;
  wire v22ebb5c;
  wire v9c1abc;
  wire v22f3aac;
  wire a1fdb9;
  wire v22efafa;
  wire v22fdc63;
  wire v23f1cf2;
  wire v23fc446;
  wire v22f1971;
  wire v22ef354;
  wire v22f1d4f;
  wire v23128f3;
  wire v23091d2;
  wire v22ff483;
  wire v23fbb00;
  wire v1aaddcb;
  wire v22f568c;
  wire v23fbaf0;
  wire v22f76c2;
  wire v23fcc3c;
  wire v22ef4f0;
  wire v23f0cce;
  wire v22f91a6;
  wire v2301a6d;
  wire v23f4937;
  wire v230174f;
  wire v231131d;
  wire v22f0d4e;
  wire v22f78b4;
  wire v23fcf10;
  wire v22ff8ea;
  wire v22f17bb;
  wire v22fe59a;
  wire v22fc2bd;
  wire v230ca57;
  wire v23fc18a;
  wire v230a671;
  wire v22f5cf0;
  wire v22fec56;
  wire v230a6ed;
  wire v2306d47;
  wire v23fb1ca;
  wire v23faca5;
  wire v2302225;
  wire v230be4a;
  wire v23084ce;
  wire b16aac;
  wire v23f38c4;
  wire b1e86b;
  wire v23fbfcd;
  wire v22f8f2b;
  wire v1aadc9e;
  wire v23fbcc2;
  wire c16bc3;
  wire v23fce79;
  wire b9c969;
  wire v230e13a;
  wire v230f9f1;
  wire v23fb231;
  wire v23fba62;
  wire v2302f72;
  wire v2302e80;
  wire v23fbb6a;
  wire v230a050;
  wire v23fca52;
  wire v22ec1f4;
  wire v22f98e7;
  wire v23fc19e;
  wire v230ce74;
  wire v22f6b57;
  wire v22edfb7;
  wire v23f200b;
  wire v23fba49;
  wire v23f2b14;
  wire v2301d23;
  wire v230d4d9;
  wire v23fc4a8;
  wire v23f4926;
  wire v23f5f78;
  wire v23f74bc;
  wire v23fc738;
  wire v23f29f5;
  wire v23097f5;
  wire v1aae9b5;
  wire v23f1db4;
  wire v2300b76;
  wire v2300a04;
  wire v22f4bae;
  wire v23fbe6a;
  wire v230a4ef;
  wire v22f4810;
  wire v23fc27a;
  wire v23fbc64;
  wire v12cd5e1;
  wire v12cd9e0;
  wire a090d5;
  wire v23f1cdf;
  wire v22ec5e3;
  wire v2310537;
  wire v1aacf10;
  wire f405e4;
  wire v23f60ba;
  wire v23fb139;
  wire v23fb70e;
  wire v10dbf63;
  wire v22f7728;
  wire v23fce08;
  wire v230430f;
  wire v23016dc;
  wire v2302de2;
  wire v1e840fa;
  wire v23fb62c;
  wire v23fab11;
  wire v23fce46;
  wire v2304b9d;
  wire v2302b3f;
  wire v22f61ac;
  wire v230468d;
  wire v23f62a3;
  wire v23fc940;
  wire v2303f9a;
  wire bd5342;
  wire v231155f;
  wire v2392e9d;
  wire v23f9c30;
  wire fc8f72;
  wire v23fc190;
  wire v22eaaef;
  wire v23ef8bb;
  wire v22efce2;
  wire v23f3c28;
  wire v22ecb5c;
  wire v2308848;
  wire v2301f3a;
  wire v22f7e80;
  wire v23fcafe;
  wire v22f4bec;
  wire v2311c5d;
  wire v23f880f;
  wire v23135fa;
  wire v230a44f;
  wire v23f7aba;
  wire v2301392;
  wire v22f2d10;
  wire v23fbe94;
  wire v23fc9c2;
  wire v23fbb3c;
  wire c25c58;
  wire v2392fd0;
  wire v23fbe44;
  wire v2310e89;
  wire v22ee2b4;
  wire v23f5868;
  wire v22eba12;
  wire v22f1393;
  wire v22fe940;
  wire v2300523;
  wire v23fbcac;
  wire v23fbd62;
  wire v23940ce;
  wire v23fbcc0;
  wire v23fcd3a;
  wire v230d4c3;
  wire v23094a3;
  wire v23fbe22;
  wire add85b;
  wire v2310e05;
  wire v230b00c;
  wire v22f18df;
  wire v230d8c2;
  wire v22f5bca;
  wire v22f331e;
  wire v23fc9de;
  wire v22f9124;
  wire v22f6894;
  wire v22f6bae;
  wire v23fb9cb;
  wire v23f9a4d;
  wire v23fcffd;
  wire v23131eb;
  wire v23f1f3f;
  wire v22ee913;
  wire v22ebd80;
  wire v17a34ff;
  wire v22f6917;
  wire v2304744;
  wire v22ef255;
  wire v22f288d;
  wire v23934cb;
  wire v230e71f;
  wire v997ca9;
  wire v8a0e71;
  wire v22f74f7;
  wire e1dcf1;
  wire v2307758;
  wire v23f4b99;
  wire v2393c48;
  wire v22ed2f0;
  wire v23fb5fa;
  wire v22fff04;
  wire v23f5a8b;
  wire v22fb74c;
  wire v22f1491;
  wire v23fc6a7;
  wire a1fd78;
  wire v22ff0d2;
  wire v22f5d15;
  wire v230dd9e;
  wire v22f9c2f;
  wire v23109c3;
  wire v23135cc;
  wire v22ecde7;
  wire v22eb292;
  wire bd7c53;
  wire v23fb159;
  wire v1aad5c9;
  wire v22ef217;
  wire v22f5204;
  wire v230f099;
  wire v2311eb3;
  wire v23fce6f;
  wire v231353a;
  wire v22ed42c;
  wire v22f19c3;
  wire v17a2d5b;
  wire v84563a;
  wire v845632;
  wire v845626;
  wire v84562a;
  wire v23f40ba;
  wire v23fc85a;
  wire bd7bf6;
  wire v2304db3;
  wire v845661;
  wire v106a782;
  wire v22f6ba1;
  wire v230cff9;
  wire v191accc;
  wire v22f3a11;
  wire v22f051d;
  wire v23f1f21;
  wire v23fcaa6;
  wire v22ebca0;
  wire v23fc93e;
  wire v23f3115;
  wire v22fb3c1;
  wire v22f9248;
  wire v2393aca;
  wire v23fb624;
  wire v991952;
  wire v23fcf35;
  wire v22f160c;
  wire v239174b;
  wire v22eedf9;
  wire v23fc1de;
  wire v2302d85;
  wire v22f442c;
  wire v23f94e5;
  wire v2302bb2;
  wire v2392842;
  wire v22f5b27;
  wire v1aad98e;
  wire v23fcfbc;
  wire v23127ff;
  wire v23fca66;
  wire v2301c57;
  wire v22ebb82;
  wire v191b1d9;
  wire v2311da1;
  wire v230702c;
  wire v22f7241;
  wire v23fba9a;
  wire v23f0872;
  wire v9ad48f;
  wire v23fb877;
  wire v23fc08c;
  wire v2300c4a;
  wire v22ebf47;
  wire v230bf6d;
  wire v919ce6;
  wire v23fc9c1;
  wire v22fab80;
  wire v2306d9e;
  wire v23043b8;
  wire v22f0380;
  wire v22ede16;
  wire v23fc1ce;
  wire b9ff2b;
  wire d962e3;
  wire v2306e28;
  wire v23fafaf;
  wire v23f5043;
  wire v2301933;
  wire v23f44b1;
  wire v23f6765;
  wire v22f84ff;
  wire v1aad4b2;
  wire v22fe74e;
  wire v22eb3ad;
  wire v23fc3f5;
  wire v23f53bd;
  wire v23fc254;
  wire v2301f92;
  wire v23f79a0;
  wire v22f5e36;
  wire b9eb75;
  wire v23fc799;
  wire v23933e8;
  wire v22f4301;
  wire v23fc96b;
  wire v23f69a3;
  wire baa1eb;
  wire v22fab90;
  wire v22fa711;
  wire v23fba3e;
  wire v23f83f3;
  wire v22f9f26;
  wire v22f6949;
  wire v22ed067;
  wire v22fdd56;
  wire v22fdbbb;
  wire v106ae3a;
  wire v22f9b3f;
  wire v23f31d3;
  wire v23fb3d1;
  wire v2301d45;
  wire v23051c4;
  wire v23fb1fc;
  wire e1e1cb;
  wire b5e222;
  wire v230c52a;
  wire v23fc161;
  wire v22fab50;
  wire v23fb81f;
  wire v230d3a4;
  wire v22eb0b1;
  wire v23fbf1e;
  wire v2311c98;
  wire v22fe775;
  wire v23f0e65;
  wire v23f04f2;
  wire v230b9f3;
  wire v22f5944;
  wire v23fbbf8;
  wire v22f0b0d;
  wire v23fcb0b;
  wire v22ef945;
  wire v2307e2c;
  wire v23fce91;
  wire v23fb24f;
  wire v22f14ed;
  wire v22ffb12;
  wire v22f3c3d;
  wire v23fc382;
  wire v22ecaef;
  wire v23007a1;
  wire v23f8a99;
  wire v22fe346;
  wire v22edcf4;
  wire v230bdad;
  wire v23f8787;
  wire v2310f77;
  wire v22ef998;
  wire a6db07;
  wire v23fbf68;
  wire v23f8ba7;
  wire v230f0de;
  wire v230a241;
  wire v22f07cd;
  wire v98c729;
  wire v22edbd4;
  wire v22feff6;
  wire v22f397b;
  wire v22ee499;
  wire v23fbe9a;
  wire v230297f;
  wire v23fc78b;
  wire v23f9f07;
  wire v22f69aa;
  wire v22eb1a8;
  wire v23fc77d;
  wire v2308b2e;
  wire a20348;
  wire v2301cee;
  wire v22f8551;
  wire v23fb964;
  wire v23fc2f6;
  wire v230aa7a;
  wire v22eb711;
  wire v23fc029;
  wire v23064bf;
  wire v230327d;
  wire v22f46ab;
  wire v23f5f07;
  wire v22f03b8;
  wire v23fb10d;
  wire v22ffaff;
  wire v23f730c;
  wire v2303c12;
  wire v23f4d72;
  wire v2310d6a;
  wire v23fccb0;
  wire v22f6d61;
  wire v2301484;
  wire v845620;
  wire v22ee59c;
  wire v23f2eb5;
  wire v22f1412;
  wire v239171e;
  wire v23f6e64;
  wire v23f7094;
  wire v23fccca;
  wire v230115b;
  wire v22fe150;
  wire v23f9a37;
  wire v22fc7c2;
  wire v88c9bf;
  wire v1506add;
  wire v23fc9e5;
  wire v22f7914;
  wire v22f3699;
  wire v22f6fa9;
  wire v23fc88f;
  wire v23fbd21;
  wire v23fcdcb;
  wire v22fe188;
  wire v22fe907;
  wire v23f2a15;
  wire v2309c55;
  wire a37ffd;
  wire v22fd008;
  wire v230fcad;
  wire v22f9fe0;
  wire v23126f2;
  wire v2311a34;
  wire v22f14ff;
  wire v1aad5a0;
  wire v23f8536;
  wire v22fc741;
  wire v23fbd79;
  wire v22fe181;
  wire v23fbfd8;
  wire v22fe542;
  wire v23915e9;
  wire v23000a6;
  wire v23fc993;
  wire v2308e0b;
  wire v22fd61b;
  wire v230764f;
  wire v23fc8bc;
  wire v23fcbe3;
  wire v23fb9b7;
  wire v23f6b11;
  wire v2301e10;
  wire v22ef1f3;
  wire bd1c32;
  wire v22f668b;
  wire v23071f4;
  wire v22ed127;
  wire v22faa24;
  wire v23fbdb7;
  wire v22fbb54;
  wire v231025b;
  wire v22ebc9f;
  wire v23fcbdc;
  wire v12cda8f;
  wire v2310fde;
  wire v22fbda1;
  wire v22f06fc;
  wire v23fc1e3;
  wire v23faf60;
  wire v2309ba2;
  wire v23fd022;
  wire v22f4bf4;
  wire v23fc539;
  wire v23effa5;
  wire v2304691;
  wire v23fc925;
  wire v22fb6f9;
  wire v22fb9eb;
  wire v2391670;
  wire v230432b;
  wire v2305498;
  wire v2305847;
  wire v22efbe2;
  wire bdac8b;
  wire v22f3e40;
  wire v2309b3a;
  wire v22fb403;
  wire v22f923c;
  wire v23f24d1;
  wire v22fdfd9;
  wire v230c4e8;
  wire v23f14e1;
  wire v22fe7b0;
  wire v23f3ff9;
  wire v22ec350;
  wire v23fc5dc;
  wire v22f1713;
  wire v23044f6;
  wire v23130da;
  wire v22ec92b;
  wire v22fc231;
  wire v231210f;
  wire v230bc37;
  wire v23fb5d0;
  wire v22f950e;
  wire v2300b4f;
  wire v230c910;
  wire v22f8afa;
  wire v23fb483;
  wire b3772b;
  wire v23fca10;
  wire v22f7ee5;
  wire v23fc0b9;
  wire v23fc932;
  wire v12cd4da;
  wire v2310037;
  wire v23fc3d8;
  wire v23fbb84;
  wire v23fab82;
  wire v23025aa;
  wire v22fb727;
  wire v22fea89;
  wire v230397f;
  wire v22ed6ac;
  wire v230192f;
  wire v23fc21a;
  wire v22ff308;
  wire v22ebee0;
  wire a92d05;
  wire v23fbcc7;
  wire v230eb8d;
  wire v22ef9df;
  wire v91ba6f;
  wire v23fc9c4;
  wire v230d8fa;
  wire v22ffe8d;
  wire v2312ae4;
  wire v2310895;
  wire v239315b;
  wire v22eaf16;
  wire v22fa7f5;
  wire v23fb913;
  wire v23fab20;
  wire v22ff33b;
  wire v23fc384;
  wire v2301d40;
  wire v23fbc06;
  wire v2304339;
  wire v23919d4;
  wire v23031b6;
  wire v23f2e42;
  wire v1507045;
  wire v22f407c;
  wire v22f2281;
  wire v2312290;
  wire bd74a3;
  wire v23fc16f;
  wire v22f3bc9;
  wire v22fc3c4;
  wire v23f133b;
  wire v2304fe7;
  wire v22f1f3f;
  wire v22ed756;
  wire v23fc953;
  wire v22f1dc9;
  wire v23fba19;
  wire a1fd70;
  wire v2303ce3;
  wire v22f0c75;
  wire v23fcb16;
  wire v22fd411;
  wire v22fef4c;
  wire v22fcc70;
  wire v2311a24;
  wire v230890f;
  wire v230de5a;
  wire v23fbdcc;
  wire v230efb1;
  wire v22ed8c2;
  wire v22ee0c4;
  wire v23fc112;
  wire v2302aac;
  wire v1506fbf;
  wire v23f30cf;
  wire v23fb084;
  wire v23fc905;
  wire v22fda6e;
  wire v96c563;
  wire v23fc887;
  wire v2310eb6;
  wire v23fba93;
  wire v230a3e6;
  wire v230c781;
  wire v23fc593;
  wire v23fbf85;
  wire a1fdf8;
  wire v2310747;
  wire v22f4828;
  wire v2309499;
  wire v23fb5b3;
  wire v23fba99;
  wire v23f9714;
  wire v23f49cd;
  wire v23f8180;
  wire v23036d1;
  wire v22ef867;
  wire v2392897;
  wire v23f4e36;
  wire v22fc3b1;
  wire v22edaa4;
  wire v2305a94;
  wire v230ac22;
  wire v23fcc21;
  wire v22f9527;
  wire v106ae43;
  wire v23f8466;
  wire v23fcf21;
  wire v230f911;
  wire v23fba32;
  wire v23fc827;
  wire v22ee657;
  wire v23fcdd8;
  wire v2311d6b;
  wire v2304a2d;
  wire v22f1498;
  wire v22ee524;
  wire v23fb681;
  wire v230deb1;
  wire v230477b;
  wire v23fbd9c;
  wire v1507157;
  wire v23fc948;
  wire v23fbf0a;
  wire v230a91b;
  wire v23fc67c;
  wire v230d667;
  wire v23fd038;
  wire v2392898;
  wire v22fe08f;
  wire v22fc0ec;
  wire v230814d;
  wire v22f3466;
  wire v23fc067;
  wire v23fcf4c;
  wire v231246b;
  wire v22f5b18;
  wire v23007f9;
  wire v22f4fb2;
  wire v2393031;
  wire v23fcc09;
  wire v23fc47e;
  wire v2300290;
  wire v191ad69;
  wire b9d049;
  wire v2305606;
  wire v22f6611;
  wire v23fc3fd;
  wire v23fcdf6;
  wire v191a905;
  wire v2311b32;
  wire v23f5fb9;
  wire v23f8062;
  wire v22eab03;
  wire v23fd016;
  wire v22ed928;
  wire v2312990;
  wire v22ed533;
  wire v23f9f89;
  wire v230e2d4;
  wire v898be2;
  wire a296f8;
  wire v2306b06;
  wire v23fce60;
  wire v23089cd;
  wire v23f8895;
  wire v22f9ca3;
  wire v23fbf08;
  wire v22ecff8;
  wire v23fc646;
  wire v23fce6b;
  wire v23f21c1;
  wire v23fc5e8;
  wire v23f3a5b;
  wire v23fc23a;
  wire v23fc1c0;
  wire bd7669;
  wire v22f831d;
  wire v22ede66;
  wire v23fb8fb;
  wire abfa28;
  wire v22f5820;
  wire v23fbddc;
  wire v23f61ba;
  wire v23008e6;
  wire v23f7f9d;
  wire v9e23c0;
  wire v9d1fa2;
  wire v2309248;
  wire v2311f22;
  wire v23fbb7b;
  wire v22f457a;
  wire v23080be;
  wire v23fca48;
  wire v23f0699;
  wire v230153c;
  wire v22f6f16;
  wire v23f2ec0;
  wire v23079bc;
  wire v23fbdc0;
  wire v2309b63;
  wire v22fab02;
  wire f40628;
  wire v22ef377;
  wire v23fcc44;
  wire v1b87776;
  wire v22f1f55;
  wire v23f3768;
  wire v23fc76e;
  wire v22fcf35;
  wire v23fa031;
  wire v23fbe85;
  wire v22f509a;
  wire v230524c;
  wire v22ffc85;
  wire v8d07e3;
  wire v23fc7ab;
  wire v22fdd65;
  wire v22f4266;
  wire v23fb90a;
  wire v23fbe95;
  wire v23f193e;
  wire v22f313c;
  wire v2302ca7;
  wire v23fc721;
  wire v22ef734;
  wire v22fd169;
  wire v23fcc25;
  wire v22f6bba;
  wire v230790b;
  wire v22fb011;
  wire bd74cf;
  wire v23f24d5;
  wire v2304965;
  wire v2300c23;
  wire v239162d;
  wire v23f1908;
  wire v23104a1;
  wire v22fe605;
  wire v2311771;
  wire v2301934;
  wire v22f5a56;
  wire v2312186;
  wire v22f47c6;
  wire v23fca36;
  wire b0df38;
  wire v22ee703;
  wire v23fc275;
  wire v23f91d0;
  wire v2312885;
  wire v23fcfed;
  wire v22fb42c;
  wire v22ec240;
  wire v23fb9c1;
  wire v23fc009;
  wire v1aae124;
  wire e1e34d;
  wire v22ef35b;
  wire v23fb13c;
  wire v22eaf27;
  wire v22ebc38;
  wire v2310a50;
  wire v23046a7;
  wire v22eb4b3;
  wire v23fba11;
  wire v23fbcaa;
  wire v2302b5b;
  wire v230cb83;
  wire v2308980;
  wire v22f2aff;
  wire v23fccf0;
  wire v15071f7;
  wire v23f6ec6;
  wire v23fc647;
  wire v23fbfa5;
  wire v2306cad;
  wire v23f78c4;
  wire v2300420;
  wire v23f7822;
  wire v22f800e;
  wire v2311cea;
  wire v22eb8fb;
  wire v22f0945;
  wire v230c469;
  wire v23fc249;
  wire v23fcaa1;
  wire v2305b74;
  wire v22f2d05;
  wire v230105a;
  wire v22f1691;
  wire v230164e;
  wire v2391b49;
  wire v23f4ca0;
  wire v23121b5;
  wire f40d9e;
  wire v230d5aa;
  wire v23fa463;
  wire v23f2a5b;
  wire v22ed5be;
  wire v1aad31c;
  wire v23f0776;
  wire v230af0f;
  wire v22f9554;
  wire v85c335;
  wire v22f064a;
  wire v23f3724;
  wire v2309c52;
  wire v22ef350;
  wire v2310b0b;
  wire v23fa8c7;
  wire v22ed975;
  wire v106a831;
  wire v983a4e;
  wire v23fb1e0;
  wire v22fd6c0;
  wire v22f8e09;
  wire v22fcf52;
  wire v23f76dc;
  wire v22f908b;
  wire v23fc891;
  wire v22edbc3;
  wire v23fc07d;
  wire v22ff123;
  wire v23f4e3d;
  wire v23fcff1;
  wire v23fc8eb;
  wire v23f51a4;
  wire v23fb98a;
  wire v22f2cf1;
  wire v23fbd0d;
  wire v22fb744;
  wire a2e978;
  wire v22f3b2e;
  wire v22ec2e9;
  wire v22fd693;
  wire v22f85f2;
  wire v230d1ff;
  wire v22f5378;
  wire b7427f;
  wire v23f6045;
  wire v2310812;
  wire v8e4c22;
  wire v230a035;
  wire v230a56a;
  wire v2312ef7;
  wire v23051eb;
  wire v23095df;
  wire v23fbc3d;
  wire v23f8410;
  wire v23fca7d;
  wire v23fba08;
  wire v23919ec;
  wire v230439f;
  wire v93dace;
  wire v230c0b8;
  wire v22ef6ce;
  wire v230299b;
  wire v22f1e67;
  wire e1e358;
  wire v2310db9;
  wire v23fb94a;
  wire v23057a4;
  wire v23f3ce8;
  wire v22f5d45;
  wire v23fbe8f;
  wire v22ef0a0;
  wire v22ee9be;
  wire v23fbeaa;
  wire v2310657;
  wire v22ebf1f;
  wire v22fd0cd;
  wire v230f9e8;
  wire v23f08a4;
  wire v2312cc9;
  wire v23f4fcd;
  wire v23fbd90;
  wire v22f2ffd;
  wire v22f8e53;
  wire v23fc8e6;
  wire v23f53c1;
  wire v23fb998;
  wire v22ece21;
  wire v230caee;
  wire v1e841ad;
  wire v23fbd91;
  wire v230fbe2;
  wire v1506af9;
  wire v22ed6c5;
  wire v22f0785;
  wire v23fcd73;
  wire bd74c0;
  wire v23919a5;
  wire v22f2db0;
  wire v22fc99c;
  wire v13affaa;
  wire v230a2bd;
  wire v23fb104;
  wire v1aae98c;
  wire v23089c5;
  wire v23f67e2;
  wire v15072de;
  wire v23fa2ec;
  wire b3cfb7;
  wire v2301aa7;
  wire v22f0073;
  wire v230de81;
  wire v23fa1f4;
  wire v15074fb;
  wire v22fce8b;
  wire v22ef270;
  wire v23fcab8;
  wire v22f7efa;
  wire v22f343b;
  wire v230446f;
  wire v23018a8;
  wire v22f814a;
  wire v2301655;
  wire v22ff4e2;
  wire v22fc0a4;
  wire v23fcf07;
  wire v22ffea0;
  wire v2305031;
  wire v22ee7a7;
  wire v23fca06;
  wire v22f4527;
  wire v22fa68b;
  wire v2308a75;
  wire v231181c;
  wire v23fc110;
  wire v230882d;
  wire v22fc569;
  wire v22f15fe;
  wire v23f3c12;
  wire v23025ab;
  wire v23f60ef;
  wire v23efe71;
  wire v22ef8a9;
  wire v23f7564;
  wire v22fc4d8;
  wire v9585ce;
  wire v2302071;
  wire v23fcdc9;
  wire v23036ca;
  wire v23f366d;
  wire v23f5218;
  wire v23fcf70;
  wire v22ec3c3;
  wire v22ee0d5;
  wire v2392fa3;
  wire v230af81;
  wire v2309d55;
  wire v22ff914;
  wire v22fb89a;
  wire v23fbd16;
  wire v230be24;
  wire v2393ac5;
  wire v22fb8d6;
  wire v23fbe66;
  wire v2311ef7;
  wire v23f039f;
  wire b9c9ef;
  wire v22ef816;
  wire v22fc13d;
  wire e1e70f;
  wire v23fa9b8;
  wire v22f90af;
  wire v230560c;
  wire v2302c45;
  wire v22ff244;
  wire v22ebdbc;
  wire v2304922;
  wire v23f6470;
  wire v23fb083;
  wire v230f2dc;
  wire v22fda32;
  wire v23f789c;
  wire v23f23fb;
  wire v2311756;
  wire v23fcfb4;
  wire v22f0698;
  wire v230cb53;
  wire v22f4a16;
  wire v2392f6b;
  wire v2393508;
  wire v22f05b9;
  wire v22fd7d4;
  wire v87cfb8;
  wire v23fc530;
  wire v2306405;
  wire v22f2bf1;
  wire ad6e26;
  wire v23fb865;
  wire v22fdd8a;
  wire v2301a99;
  wire v924a36;
  wire v2307aeb;
  wire bd7476;
  wire v22f13e3;
  wire v23f4c8c;
  wire v23fce3a;
  wire v23f4fa4;
  wire v2302907;
  wire v23f5c9b;
  wire v23fc4f7;
  wire v230f5ee;
  wire v22ec782;
  wire v23fb9c6;
  wire v2310641;
  wire v230e551;
  wire v230828b;
  wire v23067c1;
  wire v22fa700;
  wire v2311214;
  wire v22ecbc3;
  wire v231089e;
  wire v23f608b;
  wire a1fe5a;
  wire v230fd1b;
  wire v23fb98b;
  wire v23f24c0;
  wire v2303481;
  wire v23135cf;
  wire v1aae22e;
  wire v22ee0d6;
  wire v2312f81;
  wire v22ec7e8;
  wire v230c398;
  wire v23fc790;
  wire v23fc180;
  wire v1aad988;
  wire v23f89fc;
  wire v23fc98b;
  wire v23fb9c4;
  wire v22f3d4b;
  wire v22f92a2;
  wire v22fdf3c;
  wire v22ff1d8;
  wire v22f2a2f;
  wire v23fcb7c;
  wire v22ef0de;
  wire v230554d;
  wire v230ec4a;
  wire v1e84170;
  wire v22f125c;
  wire v23fc0bf;
  wire v239345a;
  wire v23fb994;
  wire v22f5840;
  wire v22faac8;
  wire v2306070;
  wire v23109e9;
  wire v22fca61;
  wire v23fccfe;
  wire f40d2a;
  wire v23fc6fe;
  wire v22fd533;
  wire v23050c3;
  wire v2391a4f;
  wire v23f76a5;
  wire v23faa5c;
  wire v2301a04;
  wire v230df28;
  wire v230dec9;
  wire v2312be4;
  wire v23fad13;
  wire v22f1866;
  wire v22f799b;
  wire v23060e3;
  wire v23f925b;
  wire v22ed12b;
  wire v22f6f0c;
  wire v191afde;
  wire v22f0ceb;
  wire v22f82ea;
  wire v23117c5;
  wire v23fbdf3;
  wire v23f84b5;
  wire v230a941;
  wire v22eeb7d;
  wire v22f1244;
  wire b00aa6;
  wire v2303a7f;
  wire v23fc2a7;
  wire v23fcbba;
  wire v22f8f0b;
  wire v23f4462;
  wire v230979f;
  wire v23fb8a7;
  wire v22f70f4;
  wire v23007f2;
  wire v23fb3cf;
  wire v23fbb1c;
  wire v230415a;
  wire e1dcf4;
  wire v23fbe0a;
  wire v22ffa10;
  wire v23fb809;
  wire v22fc1df;
  wire v23f552d;
  wire v22ebddc;
  wire v22edd99;
  wire v22f04eb;
  wire v12cda44;
  wire v23fc200;
  wire v2307a75;
  wire v230d7b7;
  wire v22f3de9;
  wire v23fbb70;
  wire v2391545;
  wire v22fbd4b;
  wire v23fc632;
  wire v230a753;
  wire v23fafc5;
  wire bd762f;
  wire v22f64de;
  wire v230e3a0;
  wire v23f3f59;
  wire v239281b;
  wire v23fc6a3;
  wire v23fc341;
  wire v23f99f6;
  wire v23fcd63;
  wire v23fb949;
  wire v2312bfb;
  wire v22fec92;
  wire v23f446c;
  wire v22f8f5f;
  wire v23fcec3;
  wire v22fa945;
  wire v230a2bb;
  wire v22f411f;
  wire v22f9eb0;
  wire v23f963f;
  wire v2309b33;
  wire v22f4062;
  wire v23f85b5;
  wire v230cd1c;
  wire aa51ef;
  wire v2307ec5;
  wire v2312be1;
  wire v1e84057;
  wire v23066fe;
  wire v230936c;
  wire v22fdf59;
  wire v22ef4de;
  wire v22f6053;
  wire v22fa39e;
  wire v22f1962;
  wire v2308bfc;
  wire v2308ba7;
  wire v22f2e20;
  wire v23f2f40;
  wire v230e534;
  wire v23fc8d1;
  wire v23fb8ee;
  wire bf8fe1;
  wire v22ebbea;
  wire v22fa245;
  wire v22eab01;
  wire v23fc9db;
  wire v23f6f99;
  wire v230b0d6;
  wire v23086ef;
  wire v22f4d37;
  wire v230a735;
  wire v23fc7ad;
  wire v2300dab;
  wire v22f7e7a;
  wire v230681b;
  wire v230c5eb;
  wire v23f3e81;
  wire v2301997;
  wire v230fc03;
  wire v23fb498;
  wire v23f9c72;
  wire v23fcd76;
  wire v22f3e94;
  wire v2302779;
  wire v230c4a4;
  wire v22f5e60;
  wire v22ef27f;
  wire v230333f;
  wire v23fc0fc;
  wire v17a34e6;
  wire v22f2f04;
  wire v23023b3;
  wire v22f91f3;
  wire v106a7a0;
  wire v22fd29a;
  wire v22ef0b3;
  wire v23f2862;
  wire v22f79fb;
  wire v22fafd7;
  wire v230ace0;
  wire v23fc383;
  wire v22f12cd;
  wire v22ff399;
  wire v2311d9d;
  wire v2308b6b;
  wire v230d9d9;
  wire v22f3e93;
  wire v2308880;
  wire v23fcd9e;
  wire v23fb44f;
  wire v22fcc32;
  wire v1e845ac;
  wire v23fb5ad;
  wire v22fe009;
  wire v230f5d0;
  wire v230088c;
  wire v23019e7;
  wire v12cd523;
  wire v23fb054;
  wire v22faef8;
  wire v150755e;
  wire v230f1a7;
  wire v23f08e5;
  wire v2307725;
  wire v13afe7d;
  wire v22f5137;
  wire v23fb6c6;
  wire af6dff;
  wire v23051f6;
  wire v22ee44f;
  wire v23f2cbe;
  wire v23fbb8d;
  wire v23fbbb0;
  wire v2306b74;
  wire v23f9ce3;
  wire v22ee4fe;
  wire v23fb1a6;
  wire v2393c3a;
  wire v21b0f6a;
  wire v23f43cf;
  wire v22ffba8;
  wire v230a25a;
  wire v22fc80c;
  wire v23f97a7;
  wire v22f29e5;
  wire v191ad8e;
  wire bd7a67;
  wire v230ed08;
  wire v230cb0f;
  wire v23fbef6;
  wire v2307553;
  wire v23fb95f;
  wire v23f2353;
  wire v23fc083;
  wire v22ed598;
  wire v22eecbb;
  wire v23fc6f1;
  wire v2311a27;
  wire v2309897;
  wire v23121ff;
  wire v23fc32d;
  wire v23f36e9;
  wire v230e874;
  wire v87d84c;
  wire v22ec616;
  wire v22ee6cb;
  wire v230ca7c;
  wire v2303147;
  wire v23fc5a8;
  wire v230942e;
  wire v23f6890;
  wire v22f58f9;
  wire v23fc5b0;
  wire v22fb68b;
  wire v2392a0d;
  wire v2307205;
  wire v22f291f;
  wire v2304c77;
  wire v23031eb;
  wire v22f035c;
  wire v239379c;
  wire v23fcf92;
  wire v23f4eb4;
  wire v2310283;
  wire v23916fa;
  wire v23fc14d;
  wire v23fbd00;
  wire a1fe3e;
  wire v2305a79;
  wire v22fab30;
  wire v23122cd;
  wire v22fe415;
  wire v23f600f;
  wire v22f0dc3;
  wire v230d235;
  wire v23fac6d;
  wire v8c875e;
  wire v22f97fe;
  wire v230bf27;
  wire v23fc284;
  wire v230e7d6;
  wire v231248c;
  wire v23f9bd1;
  wire v2303bfd;
  wire v23fc0a4;
  wire v230fa21;
  wire v23fca96;
  wire a1fe03;
  wire v23fca0c;
  wire v23f596f;
  wire v23fcf9d;
  wire v230e100;
  wire v23117af;
  wire v22ee145;
  wire v23fc250;
  wire v230e71c;
  wire v2308fe7;
  wire v2310d44;
  wire v22fe165;
  wire v22fc997;
  wire v23fc0da;
  wire v22f7d41;
  wire v23f4fa1;
  wire v23f8383;
  wire v23fbb8a;
  wire da30f9;
  wire v231206c;
  wire v22f90bf;
  wire v150748b;
  wire v2391b6f;
  wire v23f1281;
  wire v23f0c9a;
  wire v22f1e96;
  wire v22f30fe;
  wire v23f83ef;
  wire v23f680b;
  wire v230c69b;
  wire v23fcaff;
  wire v230ed3d;
  wire v22f2429;
  wire v23f76f4;
  wire v23050a2;
  wire v22fead6;
  wire v23f909e;
  wire v22f8593;
  wire v230360b;
  wire v2307836;
  wire v23fc14e;
  wire v22f6518;
  wire v23f3d39;
  wire v23fc22d;
  wire v2307743;
  wire v22f69b7;
  wire v2391ada;
  wire v23fb096;
  wire v13b0055;
  wire v23fbeb3;
  wire v23fc6d6;
  wire v23f79f6;
  wire v22fdc37;
  wire v23fc301;
  wire v23039ea;
  wire v22fb428;
  wire v23f5057;
  wire v2303226;
  wire v22f728a;
  wire v230bb69;
  wire v22f5521;
  wire v23fca4a;
  wire v22fb592;
  wire f40a8f;
  wire v22fd9eb;
  wire v1aae19c;
  wire v23f022d;
  wire v22fa48a;
  wire v230a9a0;
  wire v23f6380;
  wire v22f5243;
  wire v2307ab1;
  wire v23fbf1a;
  wire v23fc5c7;
  wire v23fc0c2;
  wire v22ec522;
  wire v9e8d9f;
  wire v23fce57;
  wire v23125fd;
  wire v230aaa7;
  wire v22f4593;
  wire v1507009;
  wire v1aae2be;
  wire v22ed7a5;
  wire v22f709c;
  wire v23fafca;
  wire v23f855f;
  wire v22f5734;
  wire v23fb5d1;
  wire v23fb669;
  wire v22fce06;
  wire v22f0ac0;
  wire v2393f52;
  wire v23fbd03;
  wire v23f3b00;
  wire v23fcd81;
  wire v230b52c;
  wire v23faece;
  wire v22f0332;
  wire v22f3c6b;
  wire v230ce98;
  wire v23f54de;
  wire v191abd1;
  wire v22f1d05;
  wire v22eb12e;
  wire v2393f3f;
  wire v22fca63;
  wire v22fef21;
  wire v23fc63a;
  wire v191b1a1;
  wire v22f12c8;
  wire v23f7ae7;
  wire v22fac26;
  wire v23fc1df;
  wire v8d83bb;
  wire v23fbcba;
  wire v2302e98;
  wire v2391f85;
  wire v23f7370;
  wire v22fb769;
  wire v23fc43d;
  wire v22fcd49;
  wire v23fcdb1;
  wire v23efe7d;
  wire v22ffffa;
  wire v2311729;
  wire v23fc04a;
  wire v231256a;
  wire v23070de;
  wire v2301da2;
  wire v22fe036;
  wire v22f54a0;
  wire v230f75b;
  wire v23f20a8;
  wire v23f8328;
  wire v22fdb97;
  wire v22f9ef0;
  wire v23934e0;
  wire v88bc32;
  wire v23f19b4;
  wire v23fcdce;
  wire v2310fcd;
  wire v22ef0b4;
  wire v23f1160;
  wire v191b160;
  wire v230d680;
  wire v106ae25;
  wire v2312020;
  wire v106af55;
  wire v23098c0;
  wire v23f6e9c;
  wire v230a574;
  wire v22f9d19;
  wire v22ebaa4;
  wire v230e5da;
  wire v22f70bd;
  wire v2392d8a;
  wire v22fe315;
  wire v22fc690;
  wire v230960d;
  wire v23fcd6d;
  wire v23fc3f6;
  wire v23f7073;
  wire v2306854;
  wire v23fb47d;
  wire v8b7fb1;
  wire v22f9d85;
  wire v23fb966;
  wire v22ef043;
  wire v23fcd1e;
  wire v23f384c;
  wire v2303ebe;
  wire v23f2426;
  wire v23f99bb;
  wire v23f58ed;
  wire v22fe792;
  wire v23049f8;
  wire v22f8e0c;
  wire v23fc91d;
  wire v2303886;
  wire v22f52f0;
  wire v23fb9be;
  wire v2300711;
  wire v22fce66;
  wire v230b739;
  wire v106ae8b;
  wire v22f39f4;
  wire v23fc263;
  wire v23fa2c3;
  wire v231156b;
  wire v230bdd4;
  wire v23fc781;
  wire v22eff0e;
  wire v22fdb21;
  wire af3c3f;
  wire v22eced4;
  wire v230ec21;
  wire v22f63e8;
  wire v22eeaaf;
  wire v230d70b;
  wire b8656c;
  wire v23f7605;
  wire v23fca58;
  wire v2308e63;
  wire v23f2422;
  wire v22fe5b1;
  wire v23fcfcd;
  wire v23fa63b;
  wire v2393420;
  wire v23fc1c7;
  wire v230e032;
  wire v2342fc3;
  wire v23fbb7f;
  wire v2311072;
  wire v2307c2a;
  wire v23fcbdb;
  wire v22f5037;
  wire v22f993e;
  wire v22f9927;
  wire v23f111b;
  wire v22ee1d1;
  wire v230f375;
  wire v2303831;
  wire b63b0c;
  wire v22f0860;
  wire v22fc7b7;
  wire v22f2eba;
  wire v2309569;
  wire v23fc761;
  wire v23fbe6f;
  wire v2304b4d;
  wire v23f3978;
  wire v23120a3;
  wire v22ee91d;
  wire v22f517c;
  wire v23f4f9f;
  wire v1aae385;
  wire v23fca1d;
  wire v2304b2a;
  wire v230cf1d;
  wire v23fb115;
  wire v2306aef;
  wire v22ffe30;
  wire v22f525a;
  wire v23fa8aa;
  wire v22f931d;
  wire v22fbbb8;
  wire v22f9880;
  wire v23f9a81;
  wire v22ffc44;
  wire v23fb900;
  wire v2311374;
  wire v23fc98e;
  wire v23fce7e;
  wire v230fb43;
  wire v23027f9;
  wire v22ed8c4;
  wire v23fc5dd;
  wire v23fc8b2;
  wire v23f82e4;
  wire v2309d97;
  wire v23fcaab;
  wire v230d2a3;
  wire v23f20e8;
  wire v22ed645;
  wire v23fcf15;
  wire v23fc920;
  wire v23f95e1;
  wire v22ecee2;
  wire v23fc066;
  wire v23f296d;
  wire v23fcd52;
  wire v22feb0d;
  wire v23f7b33;
  wire v230cdfb;
  wire v230da35;
  wire v23fbd5c;
  wire v23fb4c7;
  wire v23fb479;
  wire v22f13cb;
  wire v230f947;
  wire v22f1fec;
  wire v22f3789;
  wire v22fbeea;
  wire v2301271;
  wire v23fbd99;
  wire bd9c50;
  wire v22fe145;
  wire v23f8013;
  wire v22fe820;
  wire v230e54d;
  wire v22fdfdd;
  wire v23fbd04;
  wire v230e1bd;
  wire v230e794;
  wire v230c58d;
  wire v23f5dab;
  wire v23fba4f;
  wire v23fbade;
  wire v22edeb5;
  wire v22fc430;
  wire v23fcd05;
  wire v23f8241;
  wire v22f9321;
  wire b8c90d;
  wire v23f6e68;
  wire v23087e9;
  wire v239308e;
  wire v22fd747;
  wire v2392adb;
  wire v23000cf;
  wire v23fc4c0;
  wire v22edcf1;
  wire v22f7484;
  wire v22fbc73;
  wire v2303811;
  wire v23f740f;
  wire v22faa86;
  wire v23fc330;
  wire v230be37;
  wire v2307a9e;
  wire v23fbb1b;
  wire v2306b1d;
  wire v23f1ff1;
  wire v22fab6a;
  wire v22ee9c4;
  wire v23f4963;
  wire v23fd021;
  wire v22f4168;
  wire v12cd3bc;
  wire b8a8d7;
  wire v22ffaef;
  wire v23fa823;
  wire v2306473;
  wire v2306f4e;
  wire v2306967;
  wire v23fd01f;
  wire v230b6d9;
  wire v23f6404;
  wire v2391e3e;
  wire v22f86d2;
  wire v23fc8a2;
  wire v22fa3f5;
  wire v23fcf14;
  wire v23fb66a;
  wire v22f8d2b;
  wire v22eddb2;
  wire v23f7ffc;
  wire v23f16fd;
  wire v2308ecc;
  wire v2307abc;
  wire v890cdd;
  wire v23fcdcf;
  wire v23fc370;
  wire v23fcbe1;
  wire v23fc30e;
  wire v22fec81;
  wire v23fbfb5;
  wire b9d0ca;
  wire v22f02bd;
  wire v22f37e5;
  wire v2312edb;
  wire v23fad54;
  wire v22edccd;
  wire v2387c0f;
  wire v230b30c;
  wire v23fab81;
  wire v2392ec8;
  wire a1bfd6;
  wire v22f06fb;
  wire v23f7f8d;
  wire v23055c3;
  wire v22fd3b1;
  wire v23f809b;
  wire v230b313;
  wire v23f5269;
  wire v150708b;
  wire v2302094;
  wire v23103e6;
  wire v2309410;
  wire v22f6d0b;
  wire v22f1841;
  wire v23fbc71;
  wire v2393501;
  wire v22f15b7;
  wire v23f69cd;
  wire v22f3e2e;
  wire v23fc840;
  wire v22f2d93;
  wire v22eea15;
  wire v23f3ab8;
  wire v2306d36;
  wire v22f2d88;
  wire v23098ce;
  wire v22fd02d;
  wire v23102b2;
  wire v23fb76c;
  wire v12cc321;
  wire v2307419;
  wire v23fc59e;
  wire v23fbe11;
  wire v230363f;
  wire v11853d9;
  wire v84564f;
  wire v22f6c1b;
  wire v22fbe6a;
  wire v231242a;
  wire v23fc577;
  wire v23fc205;
  wire v22faf60;
  wire v22ed0d9;
  wire v22f20c0;
  wire v22ee0c0;
  wire v2308a60;
  wire v230e991;
  wire v22ec2d6;
  wire v2302c42;
  wire v2309aca;
  wire v23fbf1d;
  wire v23fb54f;
  wire v22fd621;
  wire v2300562;
  wire v23fc970;
  wire v231185e;
  wire v1aae6ba;
  wire v1aae9dc;
  wire v22f65e3;
  wire v22f1d7b;
  wire v23f193c;
  wire v845643;
  wire v10dbf78;
  wire v845631;
  wire e1e78b;
  wire v22ed287;
  wire v22fd679;
  wire v1128cd1;
  wire v2308b8e;
  wire v22f4e3c;
  wire v22f4cca;
  wire v23fca94;
  wire e1df2d;
  wire v22eedac;
  wire v22fff51;
  wire v22efd39;
  wire v8fac11;
  wire v22f7722;
  wire v23fc942;
  wire v23f0b27;
  wire v23f2d6c;
  wire v22f88ee;
  wire v23fcd7a;
  wire v230b199;
  wire v2303972;
  wire v23fb0e3;
  wire v22f7378;
  wire v2302e9e;
  wire v22f2d7c;
  wire v23f525c;
  wire v2307ff9;
  wire v22ed7d3;
  wire v22ec6d9;
  wire v23fc454;
  wire v23f307c;
  wire v23fb5d6;
  wire afb25b;
  wire v22f092c;
  wire v22f21d0;
  wire v22f991b;
  wire v2313372;
  wire v230834c;
  wire v22fca2f;
  wire v23fcee9;
  wire v230c4bb;
  wire v231326a;
  wire v22f23e7;
  wire v2304962;
  wire v22fede6;
  wire bd8367;
  wire v22f09fe;
  wire v22eddc0;
  wire v22fea77;
  wire v22f5d89;
  wire v22f5e18;
  wire v23fc74c;
  wire v23fce11;
  wire v2391b46;
  wire v23fc432;
  wire v23f580c;
  wire v23f7ef3;
  wire v23fbe0e;
  wire v231003e;
  wire v2310a5e;
  wire v22feecb;
  wire v230de93;
  wire v2300815;
  wire v23fc4ca;
  wire v23fcd69;
  wire v22fa36d;
  wire v230b18b;
  wire v23f9c66;
  wire v22f86fc;
  wire v230371b;
  wire v22fdc60;
  wire bd3bb2;
  wire v23f61f7;
  wire da38c1;
  wire v230129b;
  wire v2301e9a;
  wire v23f4338;
  wire v23fbafd;
  wire v22f25c6;
  wire v23fc07c;
  wire a1fe5e;
  wire v23fc0a5;
  wire e1deb1;
  wire v230f613;
  wire v23058ba;
  wire v23fce3d;
  wire v230ac9e;
  wire v230a22e;
  wire v22f0126;
  wire v230052f;
  wire v22f065f;
  wire v22fdda4;
  wire v23034c9;
  wire v23014b0;
  wire v23fb0c7;
  wire v2306291;
  wire v22f4ab3;
  wire v191b147;
  wire v22faa0e;
  wire v2313549;
  wire v2306875;
  wire v23f468c;
  wire v91ff8a;
  wire v230020c;
  wire v23f3545;
  wire v23102f3;
  wire v230720b;
  wire v23fcc82;
  wire v23017b3;
  wire v23f3d7d;
  wire v23fc8a1;
  wire v22fd6ad;
  wire v23fb9ec;
  wire f40d81;
  wire v2302ea0;
  wire v22f06ac;
  wire v23f4572;
  wire v22ff5ea;
  wire v23fc5d3;
  wire v23f05e3;
  wire v9ee8a4;
  wire v23fc8a8;
  wire v22fe3f6;
  wire v230e1f3;
  wire v22fd283;
  wire v22f8d0c;
  wire v22f2564;
  wire v22f2817;
  wire v23022c5;
  wire v22f0870;
  wire v22f9d95;
  wire v23fbb5b;
  wire v2303507;
  wire v23fc7fe;
  wire v22f5f72;
  wire v23046fe;
  wire v23fc5f4;
  wire v22f7e09;
  wire v23fa893;
  wire v23fca17;
  wire v230d65b;
  wire v23fc4e0;
  wire v22f49e4;
  wire v23f7499;
  wire v2308f3d;
  wire v23f2513;
  wire v1aad8c1;
  wire v230e4da;
  wire v230fe8e;
  wire v22fd029;
  wire v2302022;
  wire v22f274e;
  wire v22f90a5;
  wire v23fce52;
  wire v23028fa;
  wire v23fbf2a;
  wire v22eb771;
  wire v23fbb89;
  wire v23fc58e;
  wire v1aae09e;
  wire v2303c10;
  wire v230b111;
  wire v230db01;
  wire v23f8a36;
  wire v22f2430;
  wire v23fc0d0;
  wire v23fb586;
  wire v23115f8;
  wire v22f7d5c;
  wire v2300bc5;
  wire v23051ab;
  wire v23f14c7;
  wire da3129;
  wire v22f5d49;
  wire v2305af1;
  wire v23060d4;
  wire v22f5611;
  wire v23fb49a;
  wire v2309e12;
  wire v22f1b31;
  wire v22ec5f6;
  wire v230e8d3;
  wire v22f0393;
  wire v22f6844;
  wire v23f87f4;
  wire v22eb184;
  wire v23fb786;
  wire v22f31b2;
  wire v22f925b;
  wire v2304f32;
  wire v22f19cc;
  wire v22f893a;
  wire v230aa96;
  wire v230e651;
  wire v23f4e8c;
  wire v230e167;
  wire v23fcf77;
  wire v230bc39;
  wire v22f3998;
  wire v22f882c;
  wire v23f420e;
  wire v97b973;
  wire v230ea6d;
  wire v23110a4;
  wire fc8f82;
  wire v230aef0;
  wire v23f47b3;
  wire v22ff94b;
  wire v23087bc;
  wire v22efae1;
  wire v23fb710;
  wire v22eeb07;
  wire v23f0178;
  wire v23fca37;
  wire v23f75db;
  wire v22f05ac;
  wire v22ec4d6;
  wire v22f0dc0;
  wire v22f9d79;
  wire v22f7885;
  wire v23930d2;
  wire v22f4d61;
  wire v22f621f;
  wire v150745f;
  wire e1bfb3;
  wire v23fbdc2;
  wire v230b5ad;
  wire v23fb527;
  wire v23facc2;
  wire v2310c6d;
  wire v23fbf32;
  wire v230cbf6;
  wire v23fbe18;
  wire v22fbe28;
  wire v2301319;
  wire v150718d;
  wire c1f7e4;
  wire v23fb980;
  wire v23fb796;
  wire v23fc0de;
  wire v23fbf53;
  wire v2306b9f;
  wire v22f2e9f;
  wire v97808c;
  wire v23f5d5f;
  wire v230bd8f;
  wire v22f2623;
  wire v23f89d9;
  wire v2311196;
  wire v22fa65d;
  wire v22f03ec;
  wire v23fb3c7;
  wire v22f9f88;
  wire v22eeece;
  wire v23f1afd;
  wire v2308bbe;
  wire v23f6836;
  wire abf6b6;
  wire v22fa76f;
  wire v230e916;
  wire v230eca1;
  wire v2312b99;
  wire v23fbe14;
  wire v23fc273;
  wire v23fcfa5;
  wire v2302d56;
  wire v2309add;
  wire v230c70b;
  wire c043dc;
  wire v13afeb1;
  wire v22f448b;
  wire v23f63ab;
  wire v23fccd8;
  wire bd7f79;
  wire v23fbbeb;
  wire v2307c0c;
  wire v22f8e4d;
  wire v231242d;
  wire v22f990d;
  wire v22f0768;
  wire v23fc4e8;
  wire v2310051;
  wire v2313077;
  wire aeff78;
  wire v2303db8;
  wire v23fb9b6;
  wire v1e8413d;
  wire v22f5b4b;
  wire v230dc73;
  wire v23f7d1a;
  wire bd75f3;
  wire bda6cc;
  wire v230025c;
  wire v2309d7a;
  wire v23f11ae;
  wire v230e2bd;
  wire v23fbfb7;
  wire v23facb5;
  wire v22ee394;
  wire v22fe5f9;
  wire v2303cda;
  wire v23fc30a;
  wire v23fc442;
  wire v23fcb67;
  wire v23f209f;
  wire v9d7c04;
  wire v22f11cc;
  wire v23fbe1c;
  wire v2304cd0;
  wire v22f3879;
  wire v23fbf3f;
  wire v22fd0f1;
  wire v23fc121;
  wire v2309ca8;
  wire v22f1b30;
  wire v23f8692;
  wire v2310934;
  wire v22fd532;
  wire v23fbbbf;
  wire v230b292;
  wire v23fb899;
  wire v23fbf5f;
  wire v2303fb9;
  wire v230a92e;
  wire v22f61bb;
  wire v22f1acb;
  wire v22f2ff1;
  wire v22f15e8;
  wire v2306f5b;
  wire v2309dca;
  wire v22fdc16;
  wire v23115a7;
  wire v23fc7b9;
  wire v22f848f;
  wire v23fc6ce;
  wire v23fcf51;
  wire v22fcaa6;
  wire v2306bc5;
  wire v230cff8;
  wire v2301b0c;
  wire v23103f4;
  wire v2392d45;
  wire v23fcfaa;
  wire v22fdb5c;
  wire v23fc810;
  wire v22eb8ad;
  wire v2301a90;
  wire v230e19d;
  wire v23fc2df;
  wire v23f5dca;
  wire v23fbc6b;
  wire v2306690;
  wire v22f03a7;
  wire v23029bb;
  wire v22f75d4;
  wire v22f77e4;
  wire v23f8357;
  wire v22f68fe;
  wire v2300c5a;
  wire v23fc9cb;
  wire v22ec92f;
  wire v2309280;
  wire v2307a27;
  wire v2301aab;
  wire v22f36ba;
  wire v23fc5ec;
  wire v230766b;
  wire v23f73a4;
  wire v22fba61;
  wire v22eb2f1;
  wire v22f8062;
  wire v22fb2f7;
  wire v22ff0a6;
  wire v191ad4f;
  wire v23082bc;
  wire v22f8c2f;
  wire v231271d;
  wire v23127b3;
  wire v23fc55f;
  wire v23f36a5;
  wire v230d379;
  wire v23fc945;
  wire v23efc12;
  wire v23f3a55;
  wire v230d16b;
  wire v13aff30;
  wire v2303e06;
  wire v230eb18;
  wire v23fbaf3;
  wire v2392ece;
  wire v8819d8;
  wire v230a951;
  wire v230ef5b;
  wire v23fbf2c;
  wire v2301e20;
  wire v22f6183;
  wire v230d509;
  wire v22fcf3e;
  wire v23fa91a;
  wire v230c0e9;
  wire v23007a2;
  wire v22fe097;
  wire v22f9cd7;
  wire v23fb619;
  wire v22eff6d;
  wire v191aada;
  wire v23fc921;
  wire v22f9023;
  wire v23fc6a8;
  wire v23fbf17;
  wire v22f2d2a;
  wire v23f149d;
  wire v2307a49;
  wire v23fb97a;
  wire v22fbb07;
  wire v22fd19c;
  wire v23fb820;
  wire v22f4e0b;
  wire v22efa3b;
  wire v22f8209;
  wire e1ddd0;
  wire v23fd049;
  wire v191b096;
  wire v191b0a2;
  wire v23f36f1;
  wire v22ee92e;
  wire v22fe963;
  wire v230bd6c;
  wire v23f58d2;
  wire v23fc900;
  wire v23fcc28;
  wire v22f4594;
  wire v22f03ce;
  wire v2391a89;
  wire v22f0105;
  wire v23f6f4d;
  wire v231055e;
  wire v2306b05;
  wire v22f7b8b;
  wire v23fb0d9;
  wire v22f1166;
  wire v2307a21;
  wire v23f5ae4;
  wire v2309eab;
  wire v23f9a5b;
  wire v2306c0c;
  wire e1e7a3;
  wire v2305400;
  wire v22f1324;
  wire v23fc864;
  wire v230d7e4;
  wire v230282c;
  wire v230b0f6;
  wire v230c034;
  wire v22f4809;
  wire v230464b;
  wire v230e514;
  wire v23f9370;
  wire v23f4b35;
  wire v22f0af2;
  wire v2308a4b;
  wire v230159e;
  wire v230ae4f;
  wire v23f9e9f;
  wire v23fcd8a;
  wire v23fcfa8;
  wire v23fc0f8;
  wire v9a4fb4;
  wire v1506a9c;
  wire v23fc572;
  wire v22f57e8;
  wire v231106e;
  wire v23fc77b;
  wire v2310f61;
  wire v22f3586;
  wire v230d0ed;
  wire v22eb15f;
  wire v23fb925;
  wire v23f4ce2;
  wire v2304919;
  wire v22f2957;
  wire v23f6858;
  wire v23fc6b1;
  wire v2313131;
  wire v2308c50;
  wire v23fc8a4;
  wire v22f866f;
  wire v1507464;
  wire v22eb097;
  wire v23fc3b3;
  wire v2304d64;
  wire v230067a;
  wire v23f4e63;
  wire bc65c8;
  wire v23f3ac9;
  wire v1e84072;
  wire v2309fb1;
  wire v230e165;
  wire v22fa999;
  wire v230f2d6;
  wire a84b89;
  wire v2302075;
  wire v22f92b8;
  wire v23fb928;
  wire v23077e6;
  wire v22f64e0;
  wire v23fb12a;
  wire v230d6c1;
  wire v22fc11b;
  wire v2311e62;
  wire v230679a;
  wire v23041c3;
  wire v22eb682;
  wire v2304bd1;
  wire v23fc923;
  wire v230e598;
  wire v22edc4f;
  wire v22ee184;
  wire v23f6a00;
  wire v22f8556;
  wire v22f069f;
  wire v23fc6e5;
  wire v23fc460;
  wire v23fb8ec;
  wire v23006f8;
  wire v22fb653;
  wire v1aad527;
  wire v23f7688;
  wire v23fb137;
  wire v23fccec;
  wire v230571c;
  wire v22f766b;
  wire v2309130;
  wire v23fcafd;
  wire v2312da9;
  wire v23f40da;
  wire v230e185;
  wire v2304574;
  wire v22edf62;
  wire v23fc06c;
  wire v22fc374;
  wire v23038dd;
  wire v23fc2fe;
  wire v22f35fd;
  wire v22fa69c;
  wire v22ee36e;
  wire v23fb196;
  wire v23fc8d3;
  wire v23fbdc1;
  wire v23fbf8d;
  wire v22fe627;
  wire v2310a35;
  wire v23f4cf7;
  wire v23fbee9;
  wire v23055fd;
  wire v1aadb61;
  wire v2303350;
  wire v2307ff1;
  wire v23fb8e7;
  wire v2306997;
  wire v2304a45;
  wire v23fba45;
  wire v23f66ec;
  wire v23f37ba;
  wire v230383e;
  wire v23fcfdf;
  wire addc42;
  wire v23fbf0d;
  wire v23f704d;
  wire v2305719;
  wire v22f743b;
  wire v230f904;
  wire v2312a3d;
  wire v2307483;
  wire v23fa21b;
  wire v23fbf07;
  wire v22fbf38;
  wire v23f7fcb;
  wire v2305b5a;
  wire v23f6ace;
  wire v22ecaeb;
  wire v23fcaa5;
  wire v23135ec;
  wire v230fd50;
  wire v23fcb3f;
  wire v22ec978;
  wire v2309bab;
  wire v23f66db;
  wire v22f88bb;
  wire v22fb8c0;
  wire v22f19dd;
  wire v22ef772;
  wire v2392ea0;
  wire bd8382;
  wire v23f5872;
  wire v23f2ecd;
  wire v22eec02;
  wire v22fff6e;
  wire v23fbe7a;
  wire v2391f87;
  wire v230c55d;
  wire v22ee338;
  wire v22f34d8;
  wire v230d25c;
  wire v22fe552;
  wire v22fb5da;
  wire v22f0fe4;
  wire v23fc1ef;
  wire v22ebc57;
  wire v230fe65;
  wire v22edf86;
  wire v23faa39;
  wire v23100d2;
  wire v230c24b;
  wire v2393f41;
  wire v22f561a;
  wire v23046d0;
  wire v22fb4de;
  wire bd761f;
  wire v230b08d;
  wire v22f135c;
  wire v22f0b42;
  wire v22fb802;
  wire v23fcf60;
  wire v23f6adf;
  wire v231220c;
  wire v22fc365;
  wire v22f4d17;
  wire e1dea8;
  wire v191a8f7;
  wire v230996e;
  wire v22f2852;
  wire v23f51cc;
  wire v230eb8e;
  wire v23fbf9d;
  wire v2309c70;
  wire da38bd;
  wire v2303046;
  wire v22f358f;
  wire b13467;
  wire v23f9a04;
  wire v22fb890;
  wire v23faaa7;
  wire v22f1d92;
  wire v2311106;
  wire v2312ad2;
  wire v22f3b00;
  wire v23fc1ab;
  wire v23fa837;
  wire v22eb359;
  wire v2304913;
  wire v22ec21e;
  wire v22f89c7;
  wire v22f0a7b;
  wire v23fb8de;
  wire v23f5c03;
  wire v230d7e2;
  wire v23f98d2;
  wire v23fd067;
  wire v23fb6e3;
  wire v22fb17b;
  wire v2312696;
  wire v23fbfc3;
  wire v230b504;
  wire v2310a40;
  wire v23fc661;
  wire v23f2c05;
  wire v23fc439;
  wire v22fcfed;
  wire v1506ffd;
  wire v963922;
  wire v22f1ece;
  wire v22ff6a2;
  wire v23fb84b;
  wire v23070d5;
  wire v22feb6e;
  wire v2309464;
  wire v22ee9ac;
  wire v22f0e2f;
  wire v230b740;
  wire v23fb0b6;
  wire v23fbcfd;
  wire v22ef3e8;
  wire v23fb71f;
  wire v22fafe4;
  wire b62970;
  wire v22f9567;
  wire v2310475;
  wire v23fa345;
  wire v23f68ab;
  wire v230ccff;
  wire v23f982d;
  wire v230cffc;
  wire v2304ec9;
  wire v23f2bfa;
  wire v2313394;
  wire v22fe8a4;
  wire v22f155f;
  wire v22f19ce;
  wire v22f3c27;
  wire v2393635;
  wire v22f8864;
  wire v22f3fec;
  wire v2309b7e;
  wire v230bd81;
  wire v230466d;
  wire v8be441;
  wire v191aec6;
  wire v23fc114;
  wire v22faef4;
  wire v22fb759;
  wire v23fb910;
  wire v2310a05;
  wire v230cae4;
  wire v23fbf97;
  wire v2302c91;
  wire v23fbdf5;
  wire v23f84f8;
  wire v22f43d7;
  wire v23f07c2;
  wire v23fb598;
  wire ab4e4e;
  wire v22ec745;
  wire v23f3ebd;
  wire v230ea4c;
  wire v9a6a67;
  wire v23fb561;
  wire v22f383b;
  wire v23fced1;
  wire v22f2bf8;
  wire a39dae;
  wire v23fc8d8;
  wire v22f8bcf;
  wire v2312025;
  wire v23f2bb9;
  wire v23fc624;
  wire af5f08;
  wire v22fe0a8;
  wire v22f28df;
  wire ab39f4;
  wire v23fbc6e;
  wire v22fdb73;
  wire v22ffb91;
  wire v22f9a85;
  wire v22f2ed0;
  wire v23fc277;
  wire v230113d;
  wire v23fb58b;
  wire v22fe22b;
  wire v12cc2ff;
  wire v22f3272;
  wire v23f1608;
  wire v22f68c3;
  wire v23fcd6e;
  wire v23fc747;
  wire v23fd055;
  wire v23fcd96;
  wire v23fc7ce;
  wire v23efb4d;
  wire v23fbbc9;
  wire v23fa397;
  wire v22f54cb;
  wire v23f0ba3;
  wire v2393742;
  wire v23f6b2f;
  wire v2305741;
  wire v2393efc;
  wire v23f1609;
  wire v22fc4a3;
  wire v1aad4fc;
  wire v23f3a07;
  wire v22f6cec;
  wire v22ec326;
  wire v23f817b;
  wire v23fb5e9;
  wire v22fc6e6;
  wire v2301bdf;
  wire v230306f;
  wire v23130de;
  wire v23fcafc;
  wire v22ed55a;
  wire v2313189;
  wire v22fbe9c;
  wire v2300962;
  wire v22f8ac3;
  wire v23fb914;
  wire v230154b;
  wire v23084c9;
  wire v2309e8e;
  wire v22fd2a3;
  wire v23fca3b;
  wire v23f8299;
  wire v23fb8d7;
  wire v191ac91;
  wire v230330a;
  wire v23f6a11;
  wire v23f5acd;
  wire v23060b1;
  wire v230fdd7;
  wire v1aad815;
  wire b031da;
  wire v22f658e;
  wire v23fb202;
  wire v2309bcf;
  wire v22ed30e;
  wire v22eb2fd;
  wire v23086ec;
  wire v22ec9a7;
  wire v23fbf9f;
  wire v23fcf43;
  wire v2310e4a;
  wire v22f5215;
  wire v23fb495;
  wire v22f847c;
  wire v230a77a;
  wire v230b780;
  wire v22fc6d7;
  wire v23fc7e9;
  wire v23037b2;
  wire v22ffacb;
  wire v23f1325;
  wire v2303102;
  wire v2310c61;
  wire v23041ed;
  wire v22eb69b;
  wire v22f7063;
  wire v230969a;
  wire v22f5e09;
  wire v845671;
  wire v23fc512;
  wire v23fbfe0;
  wire v23fb6bb;
  wire v230c6c7;
  wire v22f25ac;
  wire v106a84c;
  wire e1bacb;
  wire v23f99ec;
  wire v23fcc31;
  wire v23fcd2d;
  wire v23f5513;
  wire v2311290;
  wire v2301fc9;
  wire v23f82bb;
  wire v23916b5;
  wire v23f54e8;
  wire v23133b7;
  wire v23fbf14;
  wire v191b037;
  wire b355fd;
  wire v23fa3e0;
  wire v230fe54;
  wire v23f3d09;
  wire v23055f4;
  wire v22ff1f8;
  wire v23fb4cd;
  wire v22f1b23;
  wire v22eb75e;
  wire v230c15a;
  wire v2312e04;
  wire v2304d7a;
  wire v22f4642;
  wire v23f6b18;
  wire v230ce2b;
  wire v22ed1c4;
  wire v23fc75a;
  wire v22ffcb0;
  wire v22ff184;
  wire v22fc481;
  wire v23fbc95;
  wire v23f7933;
  wire v22f9bb3;
  wire v8920c5;
  wire v230bb9f;
  wire v22eb970;
  wire v23fbbc5;
  wire bd7ae5;
  wire v23111a4;
  wire v23f1a1f;
  wire v23fc966;
  wire v23fcfab;
  wire v23fbae0;
  wire v23f1b7a;
  wire v22f4ae7;
  wire v22edd9f;
  wire v23fc720;
  wire v22eba1d;
  wire v2304dc4;
  wire v23fb0ee;
  wire v2307c3d;
  wire v2306790;
  wire v230b77c;
  wire v22ef55f;
  wire v22f4507;
  wire v23fccc5;
  wire v23f0db6;
  wire v106a7d8;
  wire v22ebf90;
  wire v2308dcf;
  wire v23fbd41;
  wire v2309fdb;
  wire ae7427;
  wire v191ae4a;
  wire v23f302c;
  wire v23f8534;
  wire v22f0052;
  wire v23103f8;
  wire v23fc1c2;
  wire f4066e;
  wire v2302efc;
  wire v23f9b8f;
  wire v23fccd3;
  wire v22ec6f1;
  wire v22ffcae;
  wire v230892a;
  wire v22ff205;
  wire v1aad34c;
  wire v22ef507;
  wire v22fa4ea;
  wire v22f32b9;
  wire v23f5b67;
  wire v231329e;
  wire v9aa6cf;
  wire v2300791;
  wire v22ff70d;
  wire v2392122;
  wire v2309b67;
  wire v1aae9e1;
  wire v23049cc;
  wire v2300359;
  wire v22f97f5;
  wire bb5cd7;
  wire v2304da3;
  wire v230d14d;
  wire v12cd673;
  wire v23fb2ba;
  wire v23fc234;
  wire v23f3b8f;
  wire v191ab29;
  wire v23f72fe;
  wire v2312be0;
  wire v230c3d2;
  wire v22f4e48;
  wire v23fcfb2;
  wire v22fdf30;
  wire v1b87672;
  wire v230c117;
  wire v23f18f2;
  wire v22f320d;
  wire v12cd5f2;
  wire v23fb635;
  wire v23fcb90;
  wire v22f037f;
  wire v23fb482;
  wire v22f8c70;
  wire v22fe71e;
  wire v23089a5;
  wire v23f2bc5;
  wire v23f88e6;
  wire v22eda3a;
  wire v23fc6ab;
  wire v23fc546;
  wire v23f93b5;
  wire v2305f49;
  wire v22f2ece;
  wire v22eafd6;
  wire v22f367c;
  wire v22ec552;
  wire v22f39b4;
  wire v23fa14e;
  wire v2309192;
  wire v230d8b2;
  wire v1aad8ea;
  wire v23f7fb6;
  wire v22f14ee;
  wire v230a58f;
  wire v230d66e;
  wire v2312162;
  wire v22f5d62;
  wire v2391d8a;
  wire v23ef95f;
  wire v230156f;
  wire v22f372e;
  wire v23f1e80;
  wire v23fbcb1;
  wire v23fb550;
  wire v22ec330;
  wire v2392258;
  wire v2300479;
  wire v22fdbbe;
  wire v23124aa;
  wire v23fceca;
  wire v22fbc05;
  wire v22f0dd6;
  wire v22f67ef;
  wire v2311dcb;
  wire v22fd713;
  wire v2305799;
  wire v22f049f;
  wire v23fc0bc;
  wire v1506ad8;
  wire v22f549a;
  wire v22f481f;
  wire v23fcf71;
  wire v230d814;
  wire v23075a5;
  wire v22f3b33;
  wire v23fc2bf;
  wire v23fbdef;
  wire v22f898b;
  wire v2303e13;
  wire v23fb94d;
  wire v1aad63a;
  wire v23fb7e0;
  wire v23fc094;
  wire v230cd87;
  wire v22f17ed;
  wire v22f0102;
  wire v230b781;
  wire v22edf4f;
  wire v23fbcc4;
  wire v22ee10b;
  wire v22f91a8;
  wire v2306494;
  wire v23f6ac5;
  wire v230c5ea;
  wire v23f847c;
  wire v230af72;
  wire v22f2d51;
  wire v23f38ff;
  wire v23fcb47;
  wire v23fc198;
  wire v12cc6e0;
  wire fc8fd5;
  wire f4061f;
  wire v23f3dd7;
  wire v230ddf3;
  wire v23f344d;
  wire v23fb869;
  wire v230e9a6;
  wire v22f2f19;
  wire v22fba66;
  wire v23fc4f9;
  wire v2302e87;
  wire v23f66a4;
  wire v2301fe9;
  wire v2306e35;
  wire v23fc9a1;
  wire v22f20b4;
  wire v23049ad;
  wire v23f7921;
  wire v230b011;
  wire v23fbf46;
  wire v23f89f6;
  wire v23fc972;
  wire v230fcf6;
  wire v22f9b46;
  wire v23fc834;
  wire v22ebe86;
  wire v23fc2ab;
  wire v23fb04e;
  wire v23fc0e4;
  wire v2302c68;
  wire v23fb85c;
  wire v23089ec;
  wire v22f1427;
  wire v2392cdd;
  wire v23fc1fb;
  wire v94dcdf;
  wire v23efdd4;
  wire v2304937;
  wire a1fee6;
  wire v23f680a;
  wire v23f3e7f;
  wire v23fb2e5;
  wire v22f4d04;
  wire v22fa5c9;
  wire v2309963;
  wire v2308c0b;
  wire v22f2e64;
  wire v22f33d3;
  wire v23f8884;
  wire v22f7634;
  wire v23052c9;
  wire v230e579;
  wire v22f609b;
  wire v23f0734;
  wire v23389c8;
  wire v2303d95;
  wire v22fec30;
  wire v23f54f3;
  wire v23f46b3;
  wire v23fc437;
  wire v2301e43;
  wire b9d0a0;
  wire v23fbe26;
  wire v22f8cd9;
  wire v2306a5d;
  wire v23fcd0e;
  wire v22f0755;
  wire v22ee889;
  wire v2310da2;
  wire v22ee26d;
  wire v22fa05c;
  wire v22f5e57;
  wire v2309550;
  wire v22f03a0;
  wire v1aada96;
  wire v23fcfd9;
  wire v23074dd;
  wire v23fc49b;
  wire v23fb2d6;
  wire v23108db;
  wire v22f6d82;
  wire v89e88b;
  wire v23fc11a;
  wire v23001a6;
  wire v22ed0f0;
  wire ac10e3;
  wire v2309b3c;
  wire v22f53b4;
  wire v22f6ac9;
  wire v22fa652;
  wire v23083d6;
  wire v23fc102;
  wire v2307d4e;
  wire v23fcb99;
  wire v22f7e21;
  wire v23fb63f;
  wire v23fbbee;
  wire a3ace7;
  wire v22ec4ce;
  wire v2305148;
  wire v23fc6bd;
  wire v2391665;
  wire v22f5164;
  wire v22f4b2c;
  wire v23f9cc4;
  wire v230a534;
  wire v230ecba;
  wire v2305aee;
  wire v23fb736;
  wire v22f89d5;
  wire v191abf8;
  wire v230cf9a;
  wire v22f6c36;
  wire v23f4d0d;
  wire v23135a4;
  wire v22eb3fd;
  wire v2303d87;
  wire v23fbe56;
  wire v22fab7b;
  wire v23fc6a6;
  wire v23fb89b;
  wire v2393d28;
  wire v230efee;
  wire v23fafe3;
  wire v2308609;
  wire v23fba71;
  wire v95ca19;
  wire v22fccf0;
  wire v2303a2d;
  wire v23fb4e8;
  wire v23022c3;
  wire v23f2e5d;
  wire v22f6e56;
  wire v22ecce6;
  wire v22fc0ee;
  wire v23f8ca8;
  wire v23fc2b4;
  wire v230d513;
  wire v23f1faa;
  wire v22fe908;
  wire v239158e;
  wire v23f4d86;
  wire v230e628;
  wire v23fc4ce;
  wire v23125e2;
  wire v2312ea0;
  wire v22ee345;
  wire v2306126;
  wire v23fc53d;
  wire v22eb8e1;
  wire v23fce7a;
  wire v22feb39;
  wire v191aa98;
  wire v22f3834;
  wire v15075a6;
  wire v23fb99d;
  wire v230df81;
  wire v2392fc4;
  wire v22eaed2;
  wire v23fc104;
  wire v22f3c10;
  wire v22f4cb3;
  wire v23f5a4e;
  wire v1aadeea;
  wire v23f82dd;
  wire v23063de;
  wire v22f235b;
  wire v23f273d;
  wire v2302e47;
  wire v23fc63e;
  wire v9d8aae;
  wire v23f55ae;
  wire v8c25df;
  wire v23f7d9f;
  wire v22f2e41;
  wire v22f9add;
  wire v22ebd88;
  wire v23fca78;
  wire v23f65eb;
  wire v22fe19a;
  wire v230e689;
  wire v23fcfe4;
  wire v23fce9a;
  wire v22eb6ab;
  wire v23f90bc;
  wire v23fca63;
  wire v22eba97;
  wire v23f3c20;
  wire v230493b;
  wire v23fcdc4;
  wire v23fbc7d;
  wire v22f8f91;
  wire v23f6969;
  wire v22f7078;
  wire v23fcfa4;
  wire v23f1316;
  wire v23069f2;
  wire v2308a4c;
  wire v8912cf;
  wire v2303da9;
  wire v22fa628;
  wire v23f1432;
  wire v22f9db5;
  wire v23f9ae7;
  wire v230ac1b;
  wire v2312268;
  wire v23f4900;
  wire v22f7832;
  wire v22edf7b;
  wire v23f486d;
  wire v22eb06f;
  wire v23130ac;
  wire v22f2883;
  wire v23035f1;
  wire v22f4989;
  wire v23084c2;
  wire v22fdc17;
  wire v23fbff6;
  wire v22fd314;
  wire v22f5753;
  wire v22fa768;
  wire v23f2a25;
  wire v23f790a;
  wire v230eaa1;
  wire v106af1c;
  wire v230fe99;
  wire v22f98d3;
  wire v23fcc2f;
  wire v23fca89;
  wire v22fa1a2;
  wire v22f0492;
  wire v23f6646;
  wire v2301adf;
  wire v22ef44c;
  wire v12cd2e3;
  wire v23fb201;
  wire v1e840fd;
  wire v23915cb;
  wire v23f9a8e;
  wire v2313134;
  wire v23fcba6;
  wire v2303cfd;
  wire v23f8c1f;
  wire v23fca31;
  wire v23131fd;
  wire v230daec;
  wire v23f0958;
  wire v230648e;
  wire v22f53a0;
  wire v23fb21c;
  wire v23fcdca;
  wire v2302ffc;
  wire v84565b;
  wire f4076d;
  wire v23f2fb7;
  wire v23fb724;
  wire v85fc1a;
  wire v22fa655;
  wire v22fa202;
  wire v23f6a42;
  wire v862ce7;
  wire v23fcb28;
  wire v22ee413;
  wire v8632f2;
  wire v23000a7;
  wire v23f4a0f;
  wire v23f906a;
  wire v239298c;
  wire v23f7ffb;
  wire v150742d;
  wire v106ae19;
  wire v2309c8a;
  wire v23f5af5;
  wire v23f6411;
  wire v23044cf;
  wire v23f41b9;
  wire v2312189;
  wire v863ce5;
  wire v22ef862;
  wire v106ae1c;
  wire v22f8271;
  wire b5f51c;
  wire v230f2af;
  wire v22ed7a4;
  wire v22eb5a9;
  wire v23094c6;
  wire v23004f9;
  wire v22f5fa8;
  wire v23056b1;
  wire v2309057;
  wire v1b87732;
  wire v23fa95c;
  wire v22fbdcf;
  wire v23f6653;
  wire v1506fa4;
  wire v22ff6c5;
  wire v230377f;
  wire v22f3a35;
  wire v23fc4c3;
  wire v2301e4f;
  wire v2300f82;
  wire v2309317;
  wire v23f1206;
  wire v23fbda8;
  wire v23108cb;
  wire v23f1cc0;
  wire v2303ce0;
  wire v845621;
  wire v23fc755;
  wire v230463a;
  wire v23fbb0c;
  wire v23f651e;
  wire v22f695c;
  wire baa026;
  wire v2313463;
  wire v230fec6;
  wire v22f5de1;
  wire v23f3c98;
  wire v2305cac;
  wire v230f8f4;
  wire v2310c98;
  wire v23fc97f;
  wire v2305b35;
  wire v230c2f4;
  wire v22f31b9;
  wire v22f6f8f;
  wire v23f908f;
  wire b95000;
  wire v23fc3ac;
  wire v2308d63;
  wire v23f632e;
  wire v22fd15a;
  wire v230d32a;
  wire v23f6ef7;
  wire v23f0bbc;
  wire v230dd4d;
  wire v23f7a6d;
  wire v2382e8c;
  wire v22ff114;
  wire v230a0ad;
  wire v23fc640;
  wire v22f251d;
  wire v230fe87;
  wire v22feb04;
  wire v23fc575;
  wire v22fc2ca;
  wire v23fc944;
  wire v23fbd19;
  wire v23117cd;
  wire v23f216d;
  wire v23fb8f4;
  wire v2305c43;
  wire bd7535;
  wire v23fce39;
  wire v22f52a4;
  wire v23fb8c9;
  wire v23fc6be;
  wire v2303b1a;
  wire v23fb63e;
  wire v23f98a9;
  wire v12cd586;
  wire v230095f;
  wire v22ec37c;
  wire v22f2b59;
  wire a54167;
  wire v22eaee1;
  wire v22ec882;
  wire v23f317c;
  wire v23fc58b;
  wire v23007a4;
  wire v22f7830;
  wire v23fc4a1;
  wire v2309b0f;
  wire v23fc7df;
  wire v2310116;
  wire v23fba29;
  wire v106ae4a;
  wire v2308a30;
  wire b9888a;
  wire v230d346;
  wire v22f5515;
  wire v23fceb0;
  wire v230a9d5;
  wire v22f64b2;
  wire b3865a;
  wire bd7c1c;
  wire v2303e1a;
  wire v22f1f6f;
  wire v22ee581;
  wire v23f76c2;
  wire v23f51b1;
  wire v15071a5;
  wire v22f012b;
  wire v23f5276;
  wire v23f595d;
  wire v22fe497;
  wire v22ffe44;
  wire v22f2f26;
  wire v23f43d6;
  wire v22f1a14;
  wire a1ff0e;
  wire v2304118;
  wire v23f688e;
  wire v22f05a0;
  wire v13afad9;
  wire v23fbb20;
  wire v22ff92f;
  wire v23fa2e7;
  wire v22fb8d3;
  wire v230cf1a;
  wire v2304e9c;
  wire v22ef458;
  wire v22f6de3;
  wire v23fcc9a;
  wire v22fbde2;
  wire v23f3eda;
  wire v23f567b;
  wire v23f9150;
  wire v2393392;
  wire v23fb62b;
  wire v2303598;
  wire v2311df1;
  wire v2312be7;
  wire v23fbc12;
  wire be4ff1;
  wire v22ffb52;
  wire v23effbc;
  wire v22f3b18;
  wire v23f6575;
  wire v230573f;
  wire v23fba3d;
  wire v23077c2;
  wire v23fccf8;
  wire v22fb850;
  wire v23fc2ce;
  wire v2304b1d;
  wire v2311826;
  wire v2311be2;
  wire v23f1561;
  wire v22ebc28;
  wire v230dd17;
  wire v22fc8e1;
  wire v23125fb;
  wire v23091e0;
  wire v12cd5dd;
  wire v22f6ba0;
  wire v230f0a1;
  wire v22f532c;
  wire v22f9092;
  wire v1e84124;
  wire v23fc463;
  wire v22fbe99;
  wire v22fa2dd;
  wire v23fcc81;
  wire v1aada71;
  wire v23f3c2a;
  wire v23f75ce;
  wire v22f742b;
  wire v2312f44;
  wire v23f3bc9;
  wire v2312236;
  wire v22ef31d;
  wire v23fd01b;
  wire v22eec8b;
  wire v23fc0f3;
  wire v22f9acf;
  wire v2305f58;
  wire v2302d1f;
  wire v12cd9c9;
  wire v22f4a7a;
  wire v12ce9b8;
  wire v2309c2c;
  wire v979b7c;
  wire v23fc019;
  wire v22fa0d4;
  wire v2306e6f;
  wire v23fc610;
  wire v22fe551;
  wire v23fc5b4;
  wire v23f87be;
  wire v23104cf;
  wire v1aad420;
  wire v23f39d9;
  wire v23fcc1e;
  wire v13afe72;
  wire v2309f1a;
  wire v230965a;
  wire v23fcea2;
  wire v2309a44;
  wire v23fbbf6;
  wire v22f1000;
  wire v23925af;
  wire v23fcd34;
  wire v2306cae;
  wire v23fce3f;
  wire v22ed000;
  wire v230f47e;
  wire v23fcc11;
  wire v23fbb77;
  wire v23f424b;
  wire v22ef5cd;
  wire v22ee0ea;
  wire v22ee4b6;
  wire v23f354c;
  wire v22ed346;
  wire v23fc6d9;
  wire v2306d37;
  wire v22f316f;
  wire v23fba9b;
  wire v22f2730;
  wire v23fc6b3;
  wire v23fbf92;
  wire v23fc7c4;
  wire v23115ff;
  wire v22ecab8;
  wire b84511;
  wire v22fd152;
  wire v22f0d28;
  wire a15268;
  wire v23f4be7;
  wire v9932c2;
  wire v23fb540;
  wire v23fcec2;
  wire v23fc706;
  wire v22fa16b;
  wire v23fbf9c;
  wire v22f8235;
  wire v22f3ad4;
  wire v22eb67a;
  wire v2310271;
  wire v23fcfae;
  wire v22f3b15;
  wire bd94ed;
  wire v230f480;
  wire v22f5fb8;
  wire v23f47d5;
  wire v2392fbd;
  wire v230ee35;
  wire v2307c5d;
  wire v23fb487;
  wire v23005ea;
  wire v23f904c;
  wire v22f9f67;
  wire v22f2005;
  wire v23fb965;
  wire v23fcf99;
  wire v23085b7;
  wire v23fbe7c;
  wire v23f8f24;
  wire v23fcf45;
  wire v99005c;
  wire v2308277;
  wire v22f6f7e;
  wire v1e83f8d;
  wire v23fcd66;
  wire v23f2578;
  wire v23107f0;
  wire v22fe4bb;
  wire v2301a3f;
  wire v23f403e;
  wire v23f593d;
  wire v22eccfc;
  wire v23038ea;
  wire v22ed8e2;
  wire v230beb6;
  wire v23f084d;
  wire v22f8cd8;
  wire v2304cc4;
  wire v106a81a;
  wire v230697e;
  wire v22f031f;
  wire v23f4fe1;
  wire v23fc81b;
  wire v23f810b;
  wire v230b11a;
  wire v231321e;
  wire v23faa52;
  wire v22f1553;
  wire v22fa7f7;
  wire v23fbf66;
  wire v23f1e9c;
  wire v23f9fdc;
  wire v22edc8d;
  wire v2310c11;
  wire v2309b80;
  wire v230c97c;
  wire v23fa6eb;
  wire v22f8f49;
  wire v23fb4a5;
  wire v22f6c46;
  wire v23f9bcc;
  wire v23efa39;
  wire v2312060;
  wire v23f3d38;
  wire v22f166c;
  wire v2304b4e;
  wire a5666b;
  wire v22fed40;
  wire v23fc485;
  wire v23f6c8f;
  wire v22ee24a;
  wire v230ad95;
  wire v23f723b;
  wire v23f6042;
  wire v23f3f46;
  wire v23105b6;
  wire b9c955;
  wire v22f8549;
  wire v23139e3;
  wire v22f92fa;
  wire v1e8404d;
  wire v23f9fc6;
  wire v23fbbf9;
  wire v23fb975;
  wire v22f60ce;
  wire v23f6949;
  wire v230e80e;
  wire v23fb9d3;
  wire v22f244d;
  wire v22f4950;
  wire v22ecea2;
  wire v22f43ec;
  wire v2313328;
  wire v23f8263;
  wire v2391b34;
  wire v2312628;
  wire v23f5500;
  wire v23fc73b;
  wire v2302553;
  wire v22f9532;
  wire v23106c2;
  wire v22fda35;
  wire v23fbfb1;
  wire v2303cae;
  wire v23fc32e;
  wire v2308ef6;
  wire v22f658c;
  wire v23f5201;
  wire v230b91d;
  wire v23fd03b;
  wire v23f46ba;
  wire v23f4c32;
  wire v23089b2;
  wire v22f902d;
  wire v2303b9a;
  wire v230d1a6;
  wire v23fc503;
  wire v23fc578;
  wire v22f0de9;
  wire v22f7b29;
  wire v12cdab5;
  wire v22f18b5;
  wire v22ecbc1;
  wire v22f38ab;
  wire v22fef36;
  wire v22feb95;
  wire e1e73a;
  wire v22f3ca0;
  wire v2306f7b;
  wire v22feafc;
  wire v23fc0a0;
  wire v23fa577;
  wire v23f677f;
  wire v23f1c0f;
  wire e1e65a;
  wire v23fae22;
  wire v22f67fb;
  wire v2312839;
  wire v230bb2a;
  wire v2313339;
  wire v230f573;
  wire v230b62c;
  wire v22f22ec;
  wire v22f0b62;
  wire v2307d0e;
  wire v191aeb3;
  wire v2306779;
  wire v23fccd5;
  wire v2305522;
  wire v22ebd62;
  wire f40c9d;
  wire v23fd057;
  wire v23f5596;
  wire v23fbce0;
  wire v230df5c;
  wire v23fb86a;
  wire v23f5f18;
  wire v2307309;
  wire v22f9c34;
  wire v23f50dd;
  wire v2307479;
  wire v230ed07;
  wire v2307fd0;
  wire v23fcda1;
  wire v238b0d7;
  wire v23f3e19;
  wire v2391c8a;
  wire v22f7100;
  wire v22ed035;
  wire v22eeef8;
  wire v2312c62;
  wire b535c6;
  wire v22f9faa;
  wire v22fd048;
  wire b00a55;
  wire bd77c5;
  wire v22ee7e0;
  wire v23f73d7;
  wire v22f6a1b;
  wire v22fcbbb;
  wire v23078ff;
  wire v22fcc89;
  wire v230ba0a;
  wire v2312343;
  wire v22f5a6c;
  wire v23051fd;
  wire v2304781;
  wire v22f7d9a;
  wire v230017e;
  wire v23fcb60;
  wire v230b6e3;
  wire v23031c5;
  wire v23fc7cb;
  wire v22f73a9;
  wire v23fbb63;
  wire v2309cda;
  wire v23f64d3;
  wire v22faa42;
  wire v22f8c8b;
  wire v191a965;
  wire v23f960d;
  wire v22ed48a;
  wire v1e83fd9;
  wire v2308815;
  wire v22fee46;
  wire v230f08b;
  wire v1506eb2;
  wire v230538a;
  wire v22fe261;
  wire v230eb9b;
  wire v23fc365;
  wire v23fcab7;
  wire v22fbf74;
  wire v23077ec;
  wire v22fdd29;
  wire v22ee73b;
  wire v23f931e;
  wire v23fbe2d;
  wire v23f835c;
  wire v23f5c95;
  wire v22fed78;
  wire v2300cc2;
  wire v2310482;
  wire v22fc767;
  wire v2311e9f;
  wire v22eb47c;
  wire v22f6953;
  wire v22ee7ee;
  wire v22fa4c3;
  wire v23fcd13;
  wire v22fc212;
  wire v230056c;
  wire v22efce1;
  wire v23fb14d;
  wire v22f2123;
  wire v22fab33;
  wire v23fba96;
  wire v23fc616;
  wire v22eea0f;
  wire v22f438c;
  wire v230128b;
  wire v22f811e;
  wire v23f3c86;
  wire v23fbb15;
  wire v23fbeec;
  wire v23fc020;
  wire v22f3f06;
  wire v23f8395;
  wire v191a973;
  wire v23f4938;
  wire v230bdf9;
  wire v2391dfa;
  wire v23fbcfb;
  wire v22f5471;
  wire v15072cc;
  wire v22f2271;
  wire v23133bb;
  wire v22edba6;
  wire v23f65bb;
  wire v2302167;
  wire v2311a3e;
  wire v2302353;
  wire v2303a53;
  wire v230e0c0;
  wire v23f4694;
  wire v22fd106;
  wire v22eb5cc;
  wire v12cd931;
  wire v23fbfea;
  wire v2304883;
  wire v22f6fb8;
  wire v23f8825;
  wire v230313a;
  wire v22fe204;
  wire v230fb4c;
  wire v22f3d79;
  wire v22f6a0e;
  wire v230b12a;
  wire v22eedd0;
  wire v23916c0;
  wire v22f7bb9;
  wire v22ee68f;
  wire a75533;
  wire v23f42a6;
  wire v23fcc94;
  wire v22ec078;
  wire v23fa8bb;
  wire v23f1ca8;
  wire v22fd06d;
  wire v231200e;
  wire adb81d;
  wire v22ff120;
  wire v23fbc97;
  wire v2302b2c;
  wire v22fb10b;
  wire v22ec61a;
  wire v2302386;
  wire v2305d15;
  wire v22f9dd0;
  wire v23fc84e;
  wire v22fb27b;
  wire v230da3e;
  wire v23fc17f;
  wire v23fbb48;
  wire v23f8988;
  wire v22f5c4c;
  wire v22ee93b;
  wire v22f4bca;
  wire v23fc133;
  wire v23f5622;
  wire v22f071b;
  wire v23fcb10;
  wire v23fcd0c;
  wire v106ae87;
  wire v230ad0f;
  wire v23fb314;
  wire v23f0162;
  wire v230e8d0;
  wire v23fc3a1;
  wire v23f1861;
  wire v23fd034;
  wire v23fc03f;
  wire v2310ab6;
  wire v23fc327;
  wire v86a21a;
  wire v23fcdde;
  wire v23fc092;
  wire v23fb0ab;
  wire v22fe985;
  wire v2306822;
  wire v23fc4eb;
  wire v23fc8ac;
  wire v22eef3b;
  wire v2311e58;
  wire v23f6dfb;
  wire v23fc8ce;
  wire v22febdb;
  wire v106a8b9;
  wire v22f8e29;
  wire v230a1fa;
  wire v23047dd;
  wire v23fc75d;
  wire v2305abd;
  wire v22f853d;
  wire v231254f;
  wire v23f56b1;
  wire v23fc4a7;
  wire v23fc42c;
  wire v23031bc;
  wire v22f664f;
  wire v22f7988;
  wire v22f6d51;
  wire v23f87ea;
  wire v23f4b28;
  wire v23fcfb8;
  wire v22ff38e;
  wire v22fc091;
  wire b9c8ff;
  wire v23fbffe;
  wire v22f65d5;
  wire v22f9c5f;
  wire v22fb554;
  wire v22f5583;
  wire v23fc671;
  wire v2305196;
  wire v22fb77d;
  wire v23082ec;
  wire v22fc5f0;
  wire v23021b9;
  wire v23fbaae;
  wire v22ebe16;
  wire a1fde3;
  wire v23108b7;
  wire v230dc17;
  wire v2310b27;
  wire v22ecbf0;
  wire v22fda49;
  wire v23fc89a;
  wire v2306b2e;
  wire v230e473;
  wire v23f69ba;
  wire v23fbbf2;
  wire v230c0e6;
  wire v23fb9ca;
  wire v22f87a1;
  wire v22fc19c;
  wire v23f75aa;
  wire v22f03cf;
  wire v2305e79;
  wire v22fdaa5;
  wire v23fc596;
  wire v22eb3e5;
  wire v8fafbf;
  wire v22f748c;
  wire v23fc567;
  wire v22ef509;
  wire v22f98e3;
  wire v2300d93;
  wire v23fc265;
  wire v23fc3f2;
  wire v23f3297;
  wire v230cdc1;
  wire v933ab1;
  wire v230da4a;
  wire v22f4587;
  wire a1f77b;
  wire v22efcd6;
  wire v23f5a2e;
  wire v239383d;
  wire v22fee78;
  wire v2301044;
  wire v23fc839;
  wire v23fc614;
  wire v230fc56;
  wire v23fbeeb;
  wire v22eb22e;
  wire v23f2c89;
  wire v22fe37c;
  wire v2308110;
  wire v23fcb14;
  wire v22fdf25;
  wire v23fb98e;
  wire v2308d80;
  wire v23fc8a6;
  wire v22f7929;
  wire v23fcbeb;
  wire v22fc564;
  wire v23fc016;
  wire v22f0a22;
  wire a1fd0e;
  wire v23fb7ea;
  wire v23fcddd;
  wire v23fb91a;
  wire v22fb0b7;
  wire v23fbf6c;
  wire v22f8ad3;
  wire v23f1e38;
  wire v22f99e3;
  wire v23002bf;
  wire v22fce2e;
  wire v23f9fc8;
  wire v23fcf88;
  wire v230bff5;
  wire v2312d33;
  wire v230ed77;
  wire v22f860b;
  wire v23fca9e;
  wire v2307f2b;
  wire v23fc89e;
  wire v23fc64c;
  wire v22f03c8;
  wire v22f9a75;
  wire v23fbb5a;
  wire v22fccbd;
  wire v23fcab3;
  wire bd7530;
  wire v230144a;
  wire v2309b39;
  wire v2311606;
  wire v22ffff6;
  wire v23025d8;
  wire v2302783;
  wire v22f73fb;
  wire v22fa58f;
  wire v2310ec5;
  wire v22edff5;
  wire v22f0d5a;
  wire v23f01d5;
  wire v2311470;
  wire v1aae1de;
  wire v1aad517;
  wire v22f1892;
  wire v2393705;
  wire v22f01b7;
  wire a7e154;
  wire v23122b0;
  wire v2312397;
  wire v23f1a83;
  wire v2306b33;
  wire v22ec303;
  wire v22fb71d;
  wire v22f679f;
  wire v2300059;
  wire v22f74de;
  wire v22ff90b;
  wire v2307eb9;
  wire v22ffb9d;
  wire v22efeed;
  wire v230feb2;
  wire v23fbe4d;
  wire v230b20b;
  wire v22f409f;
  wire v230b9ad;
  wire v230080a;
  wire v230d910;
  wire v230e71d;
  wire v23fb66f;
  wire v2311b7c;
  wire v22f8c0b;
  wire v22f61b6;
  wire v23fbac0;
  wire v23fce2c;
  wire v23f2cbb;
  wire v23f7961;
  wire v23fc51f;
  wire v23fb1f1;
  wire v22fbea4;
  wire b094ff;
  wire v2306bb2;
  wire ba569c;
  wire v22f2c2c;
  wire v23037d2;
  wire v23fce72;
  wire v2305d2f;
  wire v22f3c11;
  wire v23fb976;
  wire v9ae938;
  wire v23f9773;
  wire bab0c9;
  wire v22f9b95;
  wire v23f660f;
  wire v23f5948;
  wire v231101b;
  wire v23106ba;
  wire v2305050;
  wire v22fb155;
  wire v22f6187;
  wire v22f0678;
  wire v23f65c8;
  wire v23f08af;
  wire v191ae7e;
  wire v22fc4af;
  wire v23039fa;
  wire v230a3b3;
  wire v2309532;
  wire v2306538;
  wire v23112ad;
  wire v2310389;
  wire v22ffea6;
  wire v22f3feb;
  wire v23fb6d7;
  wire v22ff538;
  wire v22eeff5;
  wire v23f5382;
  wire v230c439;
  wire v23fbd34;
  wire v22f5992;
  wire v230e3c5;
  wire v22ff92c;
  wire v23115f4;
  wire v230c2c5;
  wire v230e0b7;
  wire v23fb8ae;
  wire v22fe6b3;
  wire v22ed614;
  wire v23f14bc;
  wire v230545b;
  wire v22f0d4b;
  wire v22eaff1;
  wire v2303329;
  wire v22f0b79;
  wire v22ee6e8;
  wire v23f35ea;
  wire v22f4a1f;
  wire v23fcab0;
  wire v23fbb4e;
  wire v23060a6;
  wire v230a580;
  wire v22f4d65;
  wire v1b8769e;
  wire v23fc870;
  wire v231262c;
  wire v22f068b;
  wire v230ea57;
  wire v230fb0a;
  wire v22f44cc;
  wire v230322f;
  wire v23051fc;
  wire v22fc723;
  wire v2311be9;
  wire v22f9445;
  wire v231151a;
  wire v22f6ac3;
  wire v22fe657;
  wire v23fca70;
  wire v22f5b75;
  wire v23fc664;
  wire v2311094;
  wire v23fc519;
  wire v22ec894;
  wire v22f33e0;
  wire v22ff7d0;
  wire v23f6721;
  wire v2312441;
  wire v230f755;
  wire v22fe343;
  wire v23fbce6;
  wire v22f909b;
  wire v22ec9b2;
  wire v2303f50;
  wire v22f1fdb;
  wire v23fc169;
  wire v22fc98d;
  wire v23fb93c;
  wire v22ec7cf;
  wire v23fba92;
  wire v23fc261;
  wire v23fbe7f;
  wire v23fbeb2;
  wire v2391568;
  wire v23f2199;
  wire v22eb674;
  wire v23fca4d;
  wire v2301e40;
  wire v23f6aab;
  wire v22ebd72;
  wire v22f7347;
  wire v17a3514;
  wire v22ed2f5;
  wire v22f6aa3;
  wire v230b4f9;
  wire v22fcc62;
  wire v2391d2f;
  wire v2305345;
  wire v23fc136;
  wire v22f176d;
  wire v23fb6b5;
  wire v23fcfc4;
  wire v23f5e84;
  wire v23f7393;
  wire v15071ed;
  wire v2391cf3;
  wire v23f9e87;
  wire v22f58e8;
  wire v23071be;
  wire v1506a9e;
  wire v9bc7cb;
  wire v230848d;
  wire v23fc3ee;
  wire v22f62ae;
  wire be29ff;
  wire v23f9870;
  wire v2300382;
  wire v22eb52b;
  wire v22f595f;
  wire v2310476;
  wire v2311268;
  wire v239367b;
  wire v230a58e;
  wire v22fdc74;
  wire v22f2e82;
  wire v22f53c0;
  wire v23f439a;
  wire v23fc525;
  wire e1e353;
  wire v23fbee2;
  wire v22fe052;
  wire v23fce78;
  wire v230842d;
  wire v22f7c42;
  wire v23078f5;
  wire v22fb051;
  wire v22fc61a;
  wire v2312dc1;
  wire v22f891a;
  wire v23035b0;
  wire bda6a0;
  wire v191b187;
  wire v22fb95e;
  wire v22f8629;
  wire v23fcd0a;
  wire v23f75e5;
  wire v230e831;
  wire v230edb2;
  wire v23fb6cf;
  wire v2301585;
  wire v22f859d;
  wire v15075e0;
  wire v23fc566;
  wire v23fc246;
  wire v23f67bd;
  wire v23fb4a8;
  wire v23f9d5f;
  wire v22fd973;
  wire v23f4bbd;
  wire v23fc545;
  wire v23001d6;
  wire v2300004;
  wire v23f80c9;
  wire v22f065b;
  wire v23fbf3b;
  wire v22fbb0f;
  wire v23f12d0;
  wire v23f83d7;
  wire c098a9;
  wire v23f41af;
  wire v23fc642;
  wire v22f58c2;
  wire v23f9fa4;
  wire v23003f5;
  wire v2312846;
  wire v23fca6c;
  wire v2305f8e;
  wire v2304332;
  wire v22f8f64;
  wire v2311b1e;
  wire v23fc607;
  wire v23f59dc;
  wire v23f4b8f;
  wire v2308d9e;
  wire v23fbb64;
  wire v2309320;
  wire v23f70cf;
  wire v2303fec;
  wire v22fe4f6;
  wire v23fb652;
  wire v22efcc1;
  wire v23f2184;
  wire v23086b9;
  wire v23099de;
  wire v23fb47c;
  wire v22f0fd7;
  wire v230aa1f;
  wire v22f4b50;
  wire v2312608;
  wire v2392ff9;
  wire v23075dd;
  wire v2308955;
  wire v230d674;
  wire v99b664;
  wire v23f4160;
  wire v2300985;
  wire v23fc106;
  wire v23fbb99;
  wire v23f1891;
  wire v23fbfcb;
  wire v23fc9bf;
  wire v23fbc61;
  wire v2311011;
  wire v23fb384;
  wire v23013d7;
  wire v1aae37a;
  wire v23f196c;
  wire v2303650;
  wire v2308ae7;
  wire v22f2db9;
  wire v23018c4;
  wire v23fcdd7;
  wire v15072a9;
  wire v23fc387;
  wire v22ed309;
  wire v23075ba;
  wire v2301450;
  wire v22f419a;
  wire v2309dc4;
  wire v23fcdb2;
  wire v23fcdbe;
  wire fc8f95;
  wire v22ffcbf;
  wire v2311c0b;
  wire v1e840d4;
  wire v230dd15;
  wire v23fbf5c;
  wire v23fb299;
  wire v2305819;
  wire v2306597;
  wire v23f2d28;
  wire v22f595b;
  wire v22f91f1;
  wire v23027c2;
  wire v2305568;
  wire v22f28d6;
  wire v2301e50;
  wire v22f04d8;
  wire v22f483c;
  wire v23f6a95;
  wire v2308164;
  wire v230259a;
  wire v23fbe60;
  wire v22f0953;
  wire v22fadf8;
  wire v23fbf6d;
  wire v22f118a;
  wire v2313370;
  wire v23fba34;
  wire v23fc696;
  wire v99a622;
  wire v23fcb2a;
  wire v23fcc68;
  wire v23130f6;
  wire v22ef040;
  wire v22f62a9;
  wire v23f534c;
  wire v23fcfd2;
  wire v22f216d;
  wire v22fb2b4;
  wire v22f8e9a;
  wire v23010d9;
  wire v230be8f;
  wire v23fb20f;
  wire v12cd63d;
  wire v23f427e;
  wire fc8f5a;
  wire v22f6fba;
  wire v23fcabd;
  wire v23fc5bc;
  wire v22fb30f;
  wire v22ffa4c;
  wire v22ec702;
  wire v23f7086;
  wire v23fc9b9;
  wire v230dde9;
  wire v22f7ab4;
  wire v22ef9d0;
  wire v23fbb30;
  wire v230c404;
  wire v23f869a;
  wire v23063b0;
  wire v23fcff5;
  wire v23fb599;
  wire v1aae2c1;
  wire v23f9887;
  wire v22fa8c6;
  wire v23fc9d8;
  wire v2302a58;
  wire v22fd720;
  wire v22ef92c;
  wire v23fb811;
  wire v22f76ae;
  wire v23029ed;
  wire v230ef09;
  wire v230d25d;
  wire v2311568;
  wire v23f4a2c;
  wire v23fb89e;
  wire v23fa69c;
  wire v23faa19;
  wire v22fb3f4;
  wire v23f7997;
  wire v23fb1c0;
  wire v23f2df7;
  wire v191a8e5;
  wire v23f05ee;
  wire v9ce77e;
  wire v23fc23c;
  wire v23fd04d;
  wire v22ffaf3;
  wire v230f1d9;
  wire v22ec66d;
  wire v2302f85;
  wire v2306292;
  wire bdf576;
  wire bafb17;
  wire v230a579;
  wire v22ff2bf;
  wire v23f232a;
  wire v22fde54;
  wire v22efe1b;
  wire v22f9374;
  wire v23fbf0f;
  wire v23fb591;
  wire v90b913;
  wire v22eafb2;
  wire v23fbb0b;
  wire v22f3be4;
  wire v23fbcb2;
  wire v23f450b;
  wire v22ee2bb;
  wire v22ee1e6;
  wire v23024b6;
  wire v23f2eec;
  wire v22f2703;
  wire v23fbc20;
  wire v230ff42;
  wire v22f0ddd;
  wire v230db14;
  wire v230ff7d;
  wire v23015be;
  wire v23ef93c;
  wire v22fd8e1;
  wire v22eea63;
  wire v230e606;
  wire v23fc2fd;
  wire v2300597;
  wire v23f0ded;
  wire v22fddc8;
  wire v230e72d;
  wire v23fa9dd;
  wire v2368b8a;
  wire v22f3999;
  wire v2300387;
  wire v22f8c43;
  wire v230426b;
  wire v230f75a;
  wire v22f2624;
  wire v23107b6;
  wire v23fca0a;
  wire v23f55c0;
  wire v2313a33;
  wire v23fb1c8;
  wire bdac8d;
  wire v23088a4;
  wire v22f1905;
  wire v23fb1d1;
  wire v23fc3dd;
  wire v23fc63b;
  wire v22ff745;
  wire v2313041;
  wire v22ef575;
  wire v22f5e97;
  wire v239353f;
  wire fc907f;
  wire v23074c0;
  wire v23fc561;
  wire v23f10a4;
  wire v2313965;
  wire v22fa594;
  wire v23fbfd9;
  wire v23fc2fc;
  wire v22eb66f;
  wire v2310af0;
  wire v2305979;
  wire v23f39e5;
  wire v13afb01;
  wire v2310a41;
  wire v15071d8;
  wire v191afad;
  wire v1aae490;
  wire v2303e03;
  wire v23fd035;
  wire v230e779;
  wire v23f0c76;
  wire v23fc5eb;
  wire v230bb2d;
  wire v22f174d;
  wire v230dfff;
  wire v22f3579;
  wire v23fb4a3;
  wire bd7f18;
  wire v22fb23d;
  wire v23fcb6c;
  wire v23fc873;
  wire v23fcf9c;
  wire v2308dd1;
  wire v22fdce0;
  wire v23fb69d;
  wire v13b0013;
  wire v2300c97;
  wire v22ec6e7;
  wire v2393f17;
  wire v22f6056;
  wire v23fb98c;
  wire v22f6410;
  wire v2308058;
  wire v2391f4b;
  wire v23f62fe;
  wire v2392077;
  wire v23f6d19;
  wire v23fb25c;
  wire v23fb682;
  wire v22fcc0d;
  wire v98d297;
  wire v22f946f;
  wire v23fc37d;
  wire v23fc6ed;
  wire v22fd762;
  wire v23111da;
  wire v22f995e;
  wire v22eaea8;
  wire v23fc098;
  wire v2306703;
  wire v23f513d;
  wire v230f4d0;
  wire v230bba4;
  wire v22f3027;
  wire v23fc1fe;
  wire v23113e8;
  wire v22fe367;
  wire v2305258;
  wire v23efed1;
  wire v23f96f7;
  wire v23fce8b;
  wire v23fc788;
  wire v2308aef;
  wire v22ebfa3;
  wire v22f8694;
  wire v22ee06a;
  wire e1e659;
  wire v22f6721;
  wire c24c97;
  wire v22f0869;
  wire v22ff6ba;
  wire v1aadb45;
  wire v22f515e;
  wire v22ed809;
  wire v2305d6f;
  wire v23f9546;
  wire v22fb8f1;
  wire v230f846;
  wire b8cd18;
  wire v22fe95c;
  wire v23fbd26;
  wire v2308a42;
  wire v2393364;
  wire v2310251;
  wire v23f7ea0;
  wire v23fce66;
  wire v230e851;
  wire e1beab;
  wire v231050f;
  wire v22fed24;
  wire v2391b88;
  wire bc2a58;
  wire v2305748;
  wire v23fc355;
  wire v230345c;
  wire v22ec09c;
  wire v230e2d8;
  wire v23f9680;
  wire v230dcba;
  wire v22eed68;
  wire v23010f6;
  wire v23f8f1d;
  wire a7b623;
  wire v97f5b6;
  wire v23efcfb;
  wire v2308a1b;
  wire v22f128d;
  wire v23087e8;
  wire v22ee62f;
  wire v22f8477;
  wire v231324f;
  wire v23f28a1;
  wire v22f5fe4;
  wire v1aae12f;
  wire v23047e5;
  wire v23f5b7b;
  wire v2309a71;
  wire v8ce364;
  wire v23fb82c;
  wire v23f8e93;
  wire v23fbee6;
  wire v2391c72;
  wire v22fd2e2;
  wire a6a2f9;
  wire v23facdf;
  wire v2305e51;
  wire v22f0acd;
  wire v23f14e6;
  wire a1fc74;
  wire v23f3c1b;
  wire v2303a76;
  wire v22fb29c;
  wire v23fce5f;
  wire v2301ac0;
  wire v230f691;
  wire v230b3ec;
  wire v2307e4c;
  wire v23f07f9;
  wire v2312679;
  wire v22ec6c7;
  wire v22f0445;
  wire v22f6403;
  wire v23fa1cd;
  wire v23fb6a0;
  wire v22ef3f8;
  wire v23fbe36;
  wire v22fd3c7;
  wire v22faa7a;
  wire v22ff7ef;
  wire v22f20a2;
  wire v22f867e;
  wire v23fbf13;
  wire v22fede1;
  wire v2303b17;
  wire v22eedcf;
  wire v22f1ae5;
  wire v230d804;
  wire v22f2c87;
  wire v23fbc0c;
  wire v22f9d17;
  wire v23f537c;
  wire v230aeb3;
  wire v22eb74d;
  wire v230e979;
  wire v23f6723;
  wire v22f2ee3;
  wire v106af28;
  wire v2392eb5;
  wire v23f9545;
  wire v22f59e9;
  wire v23111c0;
  wire v943604;
  wire v22f6870;
  wire v23fca08;
  wire v230753a;
  wire v230e8a7;
  wire v23f53e4;
  wire v23f328e;
  wire v1aad641;
  wire v23089fa;
  wire v23fd032;
  wire v231005a;
  wire v191b038;
  wire v23082c9;
  wire v23fcb09;
  wire v23094cb;
  wire v22faa21;
  wire v23f21cf;
  wire v2311748;
  wire v22f37de;
  wire v230330d;
  wire v23072f3;
  wire v2304e28;
  wire v23fcea5;
  wire v23105aa;
  wire v230f03c;
  wire v2391b52;
  wire v231188f;
  wire v2307fb2;
  wire v2309066;
  wire v23fbc48;
  wire v23fce31;
  wire v2304d59;
  wire v230b573;
  wire v22ec41b;
  wire v22f661c;
  wire v22fd41b;
  wire v231141f;
  wire v23fc888;
  wire v22fd079;
  wire v23f886a;
  wire v23f7ba2;
  wire v22efcbf;
  wire v23fc5ca;
  wire v230f82b;
  wire v23fcad4;
  wire v22ed493;
  wire v23fba0b;
  wire v23fc047;
  wire v230eafe;
  wire v22fed5c;
  wire v22eb0b3;
  wire v22f3f2d;
  wire v23f3f40;
  wire v22f5568;
  wire v23f62ee;
  wire v1aad703;
  wire v23fc8e5;
  wire v230bbaf;
  wire v1aae296;
  wire v2301a76;
  wire v22fbd0e;
  wire v22fb214;
  wire v23fc811;
  wire v22f49ac;
  wire v22f9b6f;
  wire v23642d5;
  wire v22eb4a6;
  wire v23fb4cf;
  wire v22ff0ce;
  wire b208fd;
  wire v23f5ae3;
  wire v2392023;
  wire v22fb3c8;
  wire v23fc976;
  wire v22fa70c;
  wire v22f18ad;
  wire v2306932;
  wire v230b68b;
  wire v13aff3b;
  wire adf3a3;
  wire v22f5b73;
  wire v23f4722;
  wire v23fb2f8;
  wire v22ed83b;
  wire v230e4ef;
  wire v22f1de1;
  wire v2391d40;
  wire v22f8d38;
  wire v23091ef;
  wire v23fc14b;
  wire v1507134;
  wire v23f9424;
  wire aa6574;
  wire v23109e5;
  wire v2305bf7;
  wire v23111b2;
  wire v231347a;
  wire b572e8;
  wire v2304ed3;
  wire v22f2481;
  wire v23f763f;
  wire v23efdcb;
  wire v106a846;
  wire v23fb081;
  wire v22fc3d9;
  wire v22fc945;
  wire v230aa2f;
  wire v23fc91a;
  wire v22f591c;
  wire v1507631;
  wire v23fb5f6;
  wire v23fc46d;
  wire v230def2;
  wire v23f64dd;
  wire v22eccee;
  wire v22ec335;
  wire v23fc01e;
  wire v22f78ee;
  wire v23fbfce;
  wire v1aad518;
  wire v22fcbac;
  wire v23fbde0;
  wire v2312917;
  wire v8d030a;
  wire b7b244;
  wire v23fc9d1;
  wire v1e840f2;
  wire v23fcfcf;
  wire v22fecb6;
  wire v23f8e34;
  wire v23f70e3;
  wire v23fbf80;
  wire v22f2a24;
  wire v23015f8;
  wire v230ece0;
  wire v23fbe80;
  wire v15074df;
  wire v22f4e7f;
  wire v230e23c;
  wire v23043ec;
  wire v23fbc86;
  wire v1aad39a;
  wire v23f65ae;
  wire a1b75e;
  wire v23f5d34;
  wire v23fc4fc;
  wire v23f361e;
  wire v22fff0a;
  wire v23fbfd3;
  wire v12cd8ed;
  wire v22f1e81;
  wire v23efc03;
  wire v23f12fa;
  wire v22f6f2b;
  wire v22f654e;
  wire v2300a72;
  wire v230ac29;
  wire v23fc3fa;
  wire v22f654a;
  wire v23f1228;
  wire v23fb28e;
  wire v23fb574;
  wire v22eece2;
  wire v2308b19;
  wire v230f046;
  wire v2312ec4;
  wire v22f2e92;
  wire v22ebad7;
  wire v23fbe39;
  wire v22fd1a7;
  wire v1b876be;
  wire v2307081;
  wire v2307c44;
  wire v230c4ae;
  wire v23fc44d;
  wire v23fb946;
  wire v22fc531;
  wire v23fb708;
  wire v23fc1ea;
  wire v22f45a5;
  wire v2303c39;
  wire v2310900;
  wire v22eb05f;
  wire v23fc982;
  wire v22f5e45;
  wire v23f76d0;
  wire v22f73a3;
  wire v23fbffa;
  wire v23fb93f;
  wire v23f98d4;
  wire v22f903f;
  wire v23fb102;
  wire v22eede3;
  wire v23efb3a;
  wire v230585c;
  wire v230d5af;
  wire v22fbaf1;
  wire v22eb14c;
  wire v22f5768;
  wire v23fb50c;
  wire v23f8b2b;
  wire v22fb638;
  wire v23fb0c9;
  wire v15070ca;
  wire v239223a;
  wire v23fcb35;
  wire v23f83ff;
  wire v23fbadd;
  wire v22f19f7;
  wire v230e37a;
  wire v23122cb;
  wire v22ecb08;
  wire v23fb53c;
  wire v23f6396;
  wire v2307c17;
  wire v23126e2;
  wire v23fb545;
  wire v22fce1f;
  wire v22f4442;
  wire v23fcb57;
  wire v22febf8;
  wire v230a571;
  wire v23f1328;
  wire v1aad4d7;
  wire v23fccb2;
  wire v23fb073;
  wire v23fb1b5;
  wire v2303bf6;
  wire v22ebe70;
  wire v23f9a36;
  wire v23f763a;
  wire v23f712d;
  wire v22fcfee;
  wire v23063db;
  wire v12cc315;
  wire v22f006c;
  wire bd76c5;
  wire bd785e;
  wire v230b3a5;
  wire b7ab40;
  wire v22fe1c8;
  wire v22fd271;
  wire v22ffb6b;
  wire v23fc5b6;
  wire v22f4bea;
  wire v2393485;
  wire v23f846c;
  wire v23f8186;
  wire v22f65c9;
  wire v23f12d3;
  wire v22ede51;
  wire v22f6af6;
  wire v86c49f;
  wire v22f2a85;
  wire v23085c5;
  wire b79a15;
  wire v23fce16;
  wire v231258e;
  wire v23fc4d3;
  wire v230bf51;
  wire v2304bcb;
  wire v22f0b75;
  wire v22feca2;
  wire v23f66cf;
  wire v23fc7d4;
  wire v22fa4f7;
  wire v22ed92a;
  wire v22fa63e;
  wire v2308e08;
  wire v22fb112;
  wire v2312282;
  wire v2305b67;
  wire v230677d;
  wire v23fc0eb;
  wire v2306798;
  wire d49f4d;
  wire v23fb522;
  wire v8eb4b5;
  wire v23fc403;
  wire v23f4b56;
  wire b9d013;
  wire v23fc88c;
  wire v23fb4ba;
  wire v22f37ba;
  wire b9d00f;
  wire v22f1b4e;
  wire v230a9eb;
  wire v23fb879;
  wire v239196f;
  wire v22ee4ab;
  wire v230cc18;
  wire v12cd3f4;
  wire v22fc9cf;
  wire v23f14ce;
  wire v23fc5db;
  wire v230650d;
  wire v23f86f0;
  wire v23f7659;
  wire v2310b47;
  wire v23fd010;
  wire v23f78a4;
  wire v23fb2f7;
  wire v23fbea6;
  wire v2309a78;
  wire v22ffbb3;
  wire v2304f4c;
  wire v22efcee;
  wire v23fa511;
  wire v23fc0c7;
  wire v23fcfe9;
  wire v22ff457;
  wire v23f807d;
  wire v23fbf3e;
  wire v22fd5dd;
  wire v230f848;
  wire v2304b49;
  wire v23faada;
  wire v22fc37d;
  wire v22efcad;
  wire v23f3922;
  wire v23041a6;
  wire v231304d;
  wire v23fb9c9;
  wire v2391e26;
  wire v23f623e;
  wire v230f161;
  wire v230aec3;
  wire v22efa0a;
  wire v9bcd2e;
  wire v23fc8e4;
  wire v8fb6b6;
  wire v23fc3b8;
  wire v95fb82;
  wire v22faba5;
  wire v23008a1;
  wire v23fcc9f;
  wire v23f5c2f;
  wire v22f2cd3;
  wire v22f1259;
  wire v23fcca7;
  wire v23fb4b4;
  wire v23fc1f8;
  wire v22ed8b5;
  wire v230a092;
  wire v23f3f38;
  wire v23fcbe8;
  wire v106a7a1;
  wire v23f741d;
  wire v23f805c;
  wire v22f324c;
  wire v1aad671;
  wire v230607d;
  wire v22f57e9;
  wire v231363c;
  wire v22f07d3;
  wire v23fd00d;
  wire v23fb920;
  wire v23fc1c1;
  wire v22ef4ce;
  wire v2305926;
  wire v23fb0dd;
  wire v2309943;
  wire v2312c13;
  wire v22fb589;
  wire v2310256;
  wire v2312d0e;
  wire b9c985;
  wire v22fc88a;
  wire v230ce52;
  wire v22f6ee2;
  wire v23fc68c;
  wire v22ede7f;
  wire v22ed7d1;
  wire v23fb0ba;
  wire v23fc882;
  wire v2308e3c;
  wire v23f8176;
  wire v23f6b0f;
  wire v23fba17;
  wire v23f15af;
  wire v23026c8;
  wire v23f9081;
  wire v22f85c0;
  wire v22fbfe3;
  wire v23fcb56;
  wire v22f1ee0;
  wire v231125d;
  wire v22eb933;
  wire v22ed933;
  wire v22f0098;
  wire v23fc564;
  wire v23fc4fb;
  wire v23f3a8b;
  wire v23045ac;
  wire v230411f;
  wire v22ec5e6;
  wire v22f7f91;
  wire v23f8017;
  wire v191ab30;
  wire v23fbbe7;
  wire v230c521;
  wire v22f2805;
  wire v22f2677;
  wire v23fbf6b;
  wire v230bf1e;
  wire v23fb936;
  wire v22f41c0;
  wire v23fbba8;
  wire v230c342;
  wire v230e336;
  wire v22ed467;
  wire v22f5e63;
  wire v2308b08;
  wire v23fbde8;
  wire v230ff63;
  wire v230faa5;
  wire v230b50c;
  wire v23004f1;
  wire v23fc5a4;
  wire v22fe4be;
  wire v22f66b0;
  wire v23fcaf7;
  wire v23fc23e;
  wire v22ef9db;
  wire v230a2c6;
  wire v2310303;
  wire v231350d;
  wire f40761;
  wire v23081f5;
  wire v22fc517;
  wire v23f64e5;
  wire v22f302f;
  wire v23fc1c8;
  wire v2303ce2;
  wire v2305f5e;
  wire v22fd50f;
  wire v23fbb4b;
  wire v23efb5a;
  wire v23fcd0d;
  wire v22fe56f;
  wire v1aad8a8;
  wire v23f16dc;
  wire v23f61e5;
  wire v8d1fa5;
  wire v23006a1;
  wire v23fba52;
  wire v2311d16;
  wire v23fccb8;
  wire v23fce4d;
  wire v230ff8a;
  wire v231269d;
  wire v23f0f9a;
  wire v1aadf44;
  wire bd837d;
  wire v23fb60a;
  wire v2303cd6;
  wire v2302f63;
  wire v23fc411;
  wire v230ceb6;
  wire v2392067;
  wire v22fe816;
  wire v22f0e4e;
  wire v22ff400;
  wire v23f55fb;
  wire v23130dd;
  wire v2309f3f;
  wire v22eda7c;
  wire v23fcdc0;
  wire v1e840d3;
  wire v22ef56f;
  wire v23fcc70;
  wire v23fcebf;
  wire v23fc20e;
  wire v23fb8cc;
  wire v8f3940;
  wire v22f053b;
  wire v2308ddf;
  wire v23fbec3;
  wire v2303d2e;
  wire v23fc0f0;
  wire v2300af8;
  wire v23f6d39;
  wire v22f1c57;
  wire v230d6ca;
  wire v22f4f42;
  wire v22eff51;
  wire v94778a;
  wire v23002d1;
  wire v22f44d0;
  wire f405eb;
  wire v23fc7e3;
  wire v230e04a;
  wire v23f3166;
  wire v2305c74;
  wire v22fb406;
  wire v23fc053;
  wire v23fcb94;
  wire v23fb189;
  wire v230a413;
  wire v23fc219;
  wire v230e58e;
  wire v22ed7a8;
  wire v2306660;
  wire v23fc46e;
  wire v22f299d;
  wire e1e5c9;
  wire v2305ce8;
  wire v23fc8d9;
  wire v23006c2;
  wire v23fcb0e;
  wire v22fcb7b;
  wire v230ce72;
  wire v2308d06;
  wire v23fcf04;
  wire v23fd013;
  wire v23fb5c0;
  wire afffd9;
  wire v23f1c14;
  wire v22f0d07;
  wire v106af57;
  wire v23fbc4a;
  wire v22f1279;
  wire v23fbe8b;
  wire v23fb155;
  wire v22ff83d;
  wire v23fce75;
  wire v23f292d;
  wire v23fcab1;
  wire v23fc6f3;
  wire v22fdaa0;
  wire v23fb98f;
  wire v22eb9e7;
  wire v23fbada;
  wire v23f770f;
  wire v23fb9cf;
  wire v23fc194;
  wire v2392ef6;
  wire v22f583d;
  wire v12cd3a7;
  wire v23129e8;
  wire v23083ee;
  wire v23f957f;
  wire v22f3483;
  wire v22f8ccb;
  wire v2393327;
  wire a1fcc9;
  wire v12cd68e;
  wire v22fcf7a;
  wire v23fc59a;
  wire v22eb3e3;
  wire v23008c7;
  wire v23fbf49;
  wire v22f1682;
  wire v23f2b0b;
  wire v22ec7a2;
  wire v22f6d06;
  wire v22f277f;
  wire v2304a64;
  wire a1fe52;
  wire v23f89fe;
  wire v2304deb;
  wire v23fade4;
  wire v22fedf7;
  wire v23fb94b;
  wire v23fc7d1;
  wire v23fbe77;
  wire v23fc09c;
  wire v22f638b;
  wire v23fc34a;
  wire v22f07fc;
  wire v2302d68;
  wire v23065d6;
  wire v1aadd09;
  wire v23fc5c5;
  wire v23fbab3;
  wire v22f691e;
  wire v2306595;
  wire ae2bc6;
  wire v23fcad0;
  wire a07f9b;
  wire v22fdafe;
  wire v23faacb;
  wire v22f5b58;
  wire v23f1a8d;
  wire v2309270;
  wire v2309ffa;
  wire v23fcb69;
  wire v22f0552;
  wire v230d6b2;
  wire v230e449;
  wire f406a3;
  wire v22f94c1;
  wire bdab35;
  wire a4c73f;
  wire v2309856;
  wire v23f18fc;
  wire v230c155;
  wire v22f7070;
  wire v22fba10;
  wire v23fc884;
  wire v22f42d3;
  wire v23fcf6a;
  wire v22f2ce7;
  wire v22f7083;
  wire v230a8eb;
  wire v22f65b0;
  wire v22f3206;
  wire v230f330;
  wire v23f15fe;
  wire v23fcf8f;
  wire v23fc612;
  wire v22f46a6;
  wire v23fcd22;
  wire v2392d4f;
  wire v23f0bf1;
  wire v2308b33;
  wire v2302d69;
  wire v22fa5a0;
  wire v2302514;
  wire v2307ed4;
  wire v23fb5e8;
  wire v23f72ff;
  wire v23fcffa;
  wire v22f2653;
  wire v22f5a29;
  wire v22fa155;
  wire v23fcae5;
  wire v23f0b47;
  wire v23f6650;
  wire v22ffa1b;
  wire v22eea08;
  wire v2307b93;
  wire v23f9283;
  wire v230fd86;
  wire v22f5ca6;
  wire v2306298;
  wire v230d976;
  wire v23f2f42;
  wire v1aae9e2;
  wire bd951f;
  wire v2300d2f;
  wire v23facc9;
  wire v230792c;
  wire v23fcb9f;
  wire v23062fe;
  wire v1506ea6;
  wire v22f1dab;
  wire v150705a;
  wire v22ee561;
  wire v23fa9df;
  wire v22ebb7b;
  wire v22f802b;
  wire v231256b;
  wire v230e8ea;
  wire v230f5b9;
  wire v23fcb40;
  wire v23f51ac;
  wire v191b085;
  wire v23057f1;
  wire v22ee9d2;
  wire v22fb31a;
  wire v2311491;
  wire v2305f67;
  wire v23fb9aa;
  wire v23f1a76;
  wire b9ca52;
  wire v845639;
  wire b8f86b;
  wire v2304373;
  wire v85d975;
  wire v23fbe1f;
  wire v23fc548;
  wire b910da;
  wire v2305fe0;
  wire v22ef26f;
  wire v22f52a0;
  wire v23086d9;
  wire v23fca34;
  wire v22f9d57;
  wire v9d0518;
  wire v23f0b74;
  wire v22fac3f;
  wire v22ee09d;
  wire v23fbac3;
  wire v2393527;
  wire v231124e;
  wire v23fc338;
  wire v23f614a;
  wire v22fa88a;
  wire v230d2c7;
  wire v23f5fb5;
  wire v23fbadb;
  wire v2301f63;
  wire v23fc21d;
  wire v23fc29c;
  wire v23f316e;
  wire v22f322a;
  wire v230278e;
  wire v191ae81;
  wire v23fc3bf;
  wire v2305c1f;
  wire v230c79d;
  wire v23110f1;
  wire v23fc621;
  wire v23001e2;
  wire v22fb841;
  wire v230207d;
  wire v1aad4fb;
  wire v23f1f3e;
  wire v22fa068;
  wire v23fc21b;
  wire v23fc2ca;
  wire v23fb9a0;
  wire v23fcddb;
  wire v2308d51;
  wire v23f86dc;
  wire v23faae7;
  wire v22f16ad;
  wire v22f29e6;
  wire v23f3d91;
  wire v23fcb78;
  wire v23fc733;
  wire v23fc178;
  wire v22fd379;
  wire v23fb107;
  wire v2303539;
  wire v23fbd2e;
  wire v22f619f;
  wire v22f70d2;
  wire v23fa600;
  wire v23f5ac2;
  wire v862ae0;
  wire v22f6a93;
  wire v2309aaa;
  wire v23fcea9;
  wire v22f6607;
  wire v23fc637;
  wire v23039c0;
  wire v22f5317;
  wire v230ce9d;
  wire v22fa616;
  wire v22fff3a;
  wire v1aad3bf;
  wire v22faf11;
  wire v2305ea5;
  wire v23055b0;
  wire v23fc351;
  wire v22f366a;
  wire v23fbc07;
  wire v23fc843;
  wire v2303388;
  wire v22f8da5;
  wire v22f4998;
  wire v23fa3c0;
  wire v23f710b;
  wire v22fb1d6;
  wire v23fc2ea;
  wire v2303245;
  wire v23fc680;
  wire v230aa2c;
  wire v23fbd14;
  wire v22f0b50;
  wire v23fb9f0;
  wire v22f4f1e;
  wire v230404f;
  wire v2391b32;
  wire v23ef89d;
  wire v23f797b;
  wire e1e707;
  wire v23f6fed;
  wire v22f421a;
  wire v23119a4;
  wire v23f699c;
  wire v23068bf;
  wire v23fcead;
  wire v2346bd3;
  wire v22ed85a;
  wire v22fd8a6;
  wire v23f4d58;
  wire v23f15ac;
  wire v2300071;
  wire v2300829;
  wire v23fc192;
  wire v23fc008;
  wire v23119e0;
  wire v23f7992;
  wire v22f39a1;
  wire v22ee0e1;
  wire v230a3ec;
  wire v22fa2de;
  wire v230358b;
  wire v230de4d;
  wire v12cd995;
  wire v23fca93;
  wire v22ee959;
  wire v23f984b;
  wire v22fbf54;
  wire v23fcc10;
  wire v1e84184;
  wire v2308f46;
  wire v23f9e4f;
  wire v23fbe8e;
  wire v2312ea7;
  wire v22fd6ba;
  wire v23fc491;
  wire v15071da;
  wire v230c899;
  wire v22ff090;
  wire v230b04e;
  wire v191ae28;
  wire v22ff0d7;
  wire v22ed5a5;
  wire v22edc85;
  wire v2310a58;
  wire v2313476;
  wire v22ec060;
  wire v22ee4d5;
  wire v23f48a1;
  wire v230f795;
  wire v23fb0bb;
  wire v22fc5a9;
  wire v23fb0f3;
  wire v9ae0d1;
  wire v2391e5e;
  wire v1aad5ee;
  wire v22fb88d;
  wire v230c440;
  wire v23fc48a;
  wire v22fe62e;
  wire e1dd71;
  wire v2312999;
  wire v23fa3b8;
  wire v23045f5;
  wire v23fb5a7;
  wire v23fbc9c;
  wire v23fc478;
  wire v23f3970;
  wire a0f5d5;
  wire v22f0c90;
  wire v22f654f;
  wire v2304432;
  wire v22fdd92;
  wire v22ec77a;
  wire v230c0dd;
  wire v22fabad;
  wire v23f496d;
  wire v23fc380;
  wire v230eae5;
  wire v2306d5c;
  wire v2301d2f;
  wire v23f8486;
  wire v23fbda6;
  wire v22f7919;
  wire v8e28ac;
  wire v23fc23d;
  wire v23056bc;
  wire v23f9319;
  wire v23fbe5d;
  wire v2304f11;
  wire v22fb7ef;
  wire v23083ed;
  wire v23f8134;
  wire v22fc63c;
  wire v23fbdb0;
  wire v23fc48b;
  wire v23fb8e0;
  wire v23fc7b4;
  wire v22fe74a;
  wire v22fc34e;
  wire v22f9657;
  wire v239213c;
  wire v23fcc99;
  wire v22f0d89;
  wire v2306667;
  wire v22f5eee;
  wire v22febb1;
  wire v22f8d74;
  wire v230c65f;
  wire v230d20f;
  wire v23fbc1a;
  wire v23fbcbf;
  wire v191ac53;
  wire v22f4ebc;
  wire v22f0331;
  wire a1fd9c;
  wire v23f460c;
  wire v22feb47;
  wire v2310d2f;
  wire e1de6f;
  wire v22f79fd;
  wire v23f2be7;
  wire v23fba94;
  wire v2306b35;
  wire v230d7b4;
  wire v22eed0b;
  wire v23fb554;
  wire v22fa77b;
  wire v2302f60;
  wire v23040af;
  wire v230f6a7;
  wire v22f337b;
  wire v23fc69b;
  wire v22f5767;
  wire v22f9552;
  wire v23fa950;
  wire v230d849;
  wire v2305811;
  wire v1507071;
  wire v23f97bb;
  wire v22ed805;
  wire v23fbfd4;
  wire v2307b39;
  wire v23fb6a4;
  wire v230bf9f;
  wire v230391b;
  wire v2302db0;
  wire v22f28c4;
  wire v23fc15f;
  wire v230e295;
  wire v23003cc;
  wire v23071cd;
  wire v191b1e4;
  wire v22eb41e;
  wire v23f7aa3;
  wire v2300de3;
  wire da3886;
  wire v23facab;
  wire v22f8a7e;
  wire v22fa0e4;
  wire v23f2daf;
  wire v2309b5d;
  wire v23f6659;
  wire v2310ff6;
  wire v22f0719;
  wire v23f7d43;
  wire v230c749;
  wire v22f83f2;
  wire v230c9f0;
  wire v23f79ba;
  wire v23fc33a;
  wire v23fcb63;
  wire v22ff414;
  wire v22ee772;
  wire v22edb43;
  wire v949c12;
  wire v22eec11;
  wire v2302a2c;
  wire v22f8cb7;
  wire v22f9dfb;
  wire v23fc8f6;
  wire v22f9340;
  wire v23f8fd0;
  wire v23fce49;
  wire v22f45e9;
  wire v23f3b81;
  wire v22f0284;
  wire v230994d;
  wire v23fca59;
  wire v23fc4f4;
  wire v23fc631;
  wire v22f28f7;
  wire v22f4a68;
  wire v23fd011;
  wire v23053fb;
  wire v2300503;
  wire v23fc522;
  wire v23026db;
  wire v23f894b;
  wire v2313118;
  wire v23fa2f1;
  wire v2306944;
  wire v23f1879;
  wire v2301e1a;
  wire v2309726;
  wire v22fb757;
  wire v23fc32a;
  wire v22f5576;
  wire v22f91b6;
  wire v23fc369;
  wire v23f7e8f;
  wire v22fbc0e;
  wire v23092cd;
  wire v22f10c8;
  wire v23f5446;
  wire v231065b;
  wire v23f58a6;
  wire v22fe285;
  wire v22f2254;
  wire v23fb862;
  wire v230a942;
  wire v23fceb8;
  wire v23f7cea;
  wire v230851f;
  wire v230e962;
  wire v23088db;
  wire v23fc7dc;
  wire v22fdd61;
  wire v23fcb02;
  wire bad6eb;
  wire v22fa080;
  wire v22eb58b;
  wire v23fbcbe;
  wire v22f5dc1;
  wire v22fcf46;
  wire v892c49;
  wire v2308a8f;
  wire v23fa3fc;
  wire v23fc293;
  wire v23fbb83;
  wire v23fb8f1;
  wire v23fc99e;
  wire v2303fe4;
  wire b08eee;
  wire v22f03c1;
  wire v23fcf11;
  wire v22f1125;
  wire v22f8cee;
  wire v22edbd5;
  wire v23f8d53;
  wire v22f8ec8;
  wire v23fbc53;
  wire v22f58a9;
  wire bf9ce3;
  wire v2303b2a;
  wire v22f8001;
  wire v22f1e8e;
  wire v2393bce;
  wire v22f9b42;
  wire v22fc8c8;
  wire v23fc91f;
  wire v22fe421;
  wire v23fcc91;
  wire v23fc27d;
  wire v230ad15;
  wire v22fd7dd;
  wire v12cd8c9;
  wire v22eb334;
  wire v23fcb5b;
  wire v23fce77;
  wire v23fb581;
  wire v22fdaa1;
  wire v22f8214;
  wire v191aa95;
  wire v230dae4;
  wire v22f8b12;
  wire v230fe14;
  wire v8bc4e1;
  wire v23f7ef4;
  wire v23f65f3;
  wire v23fb924;
  wire v22ec644;
  wire v22f5a27;
  wire v23122bc;
  wire v22ed65e;
  wire v2311c4d;
  wire v23fca1c;
  wire v23f756e;
  wire v23007b3;
  wire v23f6b67;
  wire v22fea98;
  wire v23fb810;
  wire v230ae4e;
  wire v23fbab4;
  wire v23fc25a;
  wire v23fc412;
  wire a1fc9e;
  wire v230e9be;
  wire v2304c8b;
  wire v2313429;
  wire v2304d26;
  wire v23fb97e;
  wire v23fca56;
  wire v23fbf44;
  wire v23102d5;
  wire v22f1d8b;
  wire v22f94ec;
  wire v230e115;
  wire v22f5f7e;
  wire v22f0132;
  wire v23fc340;
  wire v2307f77;
  wire v22f5664;
  wire v23fc744;
  wire v2310c62;
  wire v23fbd9b;
  wire v13afc17;
  wire v23f4154;
  wire v23f7eaa;
  wire v230a355;
  wire v22fee3b;
  wire v22fccd1;
  wire v230bafe;
  wire v22ff1b0;
  wire v23f5ead;
  wire v23fa2b5;
  wire v22f9bc8;
  wire v22fffa6;
  wire v23fcb96;
  wire v23f77e8;
  wire v23f445f;
  wire v230d291;
  wire bd9c35;
  wire v22f46d3;
  wire v22ed491;
  wire v2310e10;
  wire v23fcd7f;
  wire v23fc7c6;
  wire v22f475e;
  wire v23fc723;
  wire v23024e8;
  wire v1aad9cb;
  wire v23f19ee;
  wire v22f6aa1;
  wire v23f682c;
  wire v22ebd0b;
  wire v23f910c;
  wire v23f93ee;
  wire v22f2efc;
  wire v2312580;
  wire v23fc72d;
  wire v22fa27c;
  wire v230d109;
  wire v99d709;
  wire v22ffb2b;
  wire v23f9f77;
  wire v2301216;
  wire v2309ce6;
  wire v23fb21a;
  wire v23f6478;
  wire dab2cc;
  wire v23f6114;
  wire v2308aa9;
  wire v23f8561;
  wire v2312a18;
  wire v23f7123;
  wire v2312888;
  wire v94508c;
  wire v22eb38b;
  wire v23fc497;
  wire v22f28eb;
  wire v22f451b;
  wire v23fb808;
  wire v23fc0c3;
  wire v2311476;
  wire v23f9c7b;
  wire v23fc342;
  wire v22f8d80;
  wire v22eefd1;
  wire v1507161;
  wire v85d110;
  wire v23f8edc;
  wire v23fbb9b;
  wire v2304474;
  wire v1506a4d;
  wire v23fbef7;
  wire v23f1ca1;
  wire v23f0169;
  wire v23f14ef;
  wire v230d32d;
  wire v22edd64;
  wire v230d529;
  wire v2304536;
  wire v22f9280;
  wire v230fa04;
  wire v9b33d9;
  wire v23fcfbe;
  wire v22fc70a;
  wire v230c0da;
  wire v2303fa0;
  wire v23fc890;
  wire v23f1812;
  wire v23f4007;
  wire v23fcef8;
  wire v23fca14;
  wire v23fc50e;
  wire a0e5e2;
  wire v23f45d2;
  wire v22fec8c;
  wire v12cd4c5;
  wire a25b7d;
  wire v2305a2a;
  wire v23fc4c2;
  wire v23fc87a;
  wire v23f5dcc;
  wire v23fc5fb;
  wire v22f7997;
  wire v87eb7a;
  wire v8902b0;
  wire v230b27c;
  wire v23fcba1;
  wire v23fb926;
  wire v23fca9d;
  wire v2303b86;
  wire v23fb08d;
  wire v23139b9;
  wire v963cc3;
  wire v22f8bd7;
  wire v1507118;
  wire v23f89b6;
  wire v22fdc2b;
  wire fc88bb;
  wire v23f89f0;
  wire v2307816;
  wire v22f6b3e;
  wire v2301f8c;
  wire v22f8613;
  wire v23fcc39;
  wire v2301968;
  wire v22f20cf;
  wire v22ff09a;
  wire v22ffffd;
  wire v23fb537;
  wire v22eaeaf;
  wire v2312ba0;
  wire v230ae14;
  wire v2304e51;
  wire v22f9f01;
  wire v2303ebc;
  wire v22eda43;
  wire v23f2e61;
  wire v23062f0;
  wire v1aae2a8;
  wire v230fce3;
  wire v23f082a;
  wire v23fbd13;
  wire v22f5b7c;
  wire v23f9789;
  wire v23f4526;
  wire v22f9f47;
  wire v230ba92;
  wire v23f8f18;
  wire v2300c85;
  wire v22f884c;
  wire v2312dc5;
  wire v22f09c4;
  wire v22f7303;
  wire v23043b1;
  wire v23929fd;
  wire v230efa2;
  wire v2305d50;
  wire v22edb60;
  wire v22f1754;
  wire v22f90c3;
  wire v23fcdc5;
  wire v23132cd;
  wire v2312c3f;
  wire v2304b8d;
  wire v22ece29;
  wire v22f0974;
  wire v23fbaed;
  wire v23fbbbe;
  wire v230d532;
  wire a05106;
  wire v230e800;
  wire v2304ccc;
  wire v23fcae0;
  wire v23105eb;
  wire v23fcfd0;
  wire v84571e;
  wire v2303d65;
  wire v23fcc5f;
  wire v22fb44a;
  wire v2393091;
  wire v22fab7c;
  wire v22edf31;
  wire v23f3de0;
  wire v23f3e77;
  wire v23fc5e5;
  wire v22eea6a;
  wire v23f43db;
  wire v22f8312;
  wire v22eca5d;
  wire v23fb074;
  wire v2306837;
  wire v23f883c;
  wire v23fbb9d;
  wire v22f71ee;
  wire v23fc56a;
  wire v23fbf94;
  wire v22f606c;
  wire v1aae2a5;
  wire v22f4abc;
  wire v23f15e7;
  wire v23fc5bf;
  wire v9ce189;
  wire v23fce9d;
  wire v2309b75;
  wire f4064b;
  wire v23116cd;
  wire v22ec6a7;
  wire v230e437;
  wire v2308363;
  wire v23fcc49;
  wire v23fc40a;
  wire v22eb23c;
  wire b1d009;
  wire v23f62f2;
  wire v23126b8;
  wire v22f5216;
  wire v22f297d;
  wire v23fb0bf;
  wire v23fbc9e;
  wire v230fca8;
  wire v966100;
  wire v22ee7cf;
  wire v23fbb11;
  wire v22f47b0;
  wire v23f7e43;
  wire e1e5c7;
  wire v2304fdd;
  wire bfde5b;
  wire v2311928;
  wire v22fb2dc;
  wire v2312f82;
  wire v1aae6b5;
  wire v23fc7a1;
  wire c242c8;
  wire v22ecca9;
  wire v23f182c;
  wire v2300d67;
  wire v23f2d33;
  wire v23f5ef2;
  wire v23f4861;
  wire v230fb76;
  wire v23fb745;
  wire v23fb9a7;
  wire v22fe58b;
  wire v22ed121;
  wire v23fb625;
  wire v231128c;
  wire v23f54ac;
  wire v230474b;
  wire v9052d9;
  wire v23f7cba;
  wire v230ea7f;
  wire v22f824f;
  wire v23fb973;
  wire v23fbbf3;
  wire v23fb4a6;
  wire v230f776;
  wire v22f1ca0;
  wire ac37a1;
  wire v23fb912;
  wire v22fcf71;
  wire v2311089;
  wire v23fbd80;
  wire v23060c7;
  wire v2310f46;
  wire v22ecba3;
  wire v230e6ba;
  wire v23fba97;
  wire v2303d00;
  wire v23f7218;
  wire v23fc19d;
  wire v23f3eed;
  wire v23f2a86;
  wire v23fc9aa;
  wire v22f214f;
  wire v23f3206;
  wire v22f8857;
  wire fc8c3f;
  wire v23fb099;
  wire v22eb99d;
  wire v2304189;
  wire v2305ee5;
  wire v2303c07;
  wire v22ee024;
  wire v12cd9b6;
  wire v230ab24;
  wire v23fc7b2;
  wire v22f53a6;
  wire v23f0ce0;
  wire v22ef8af;
  wire v23fb567;
  wire v23f450d;
  wire v23fc55d;
  wire v23fc818;
  wire v23fb4fd;
  wire v23f7efd;
  wire v23fb9ac;
  wire v230561d;
  wire v22fe46b;
  wire v22f1681;
  wire v23f4bcd;
  wire v23fc1c9;
  wire v23f404a;
  wire v23fc042;
  wire v2303dd7;
  wire v230fae0;
  wire a678c9;
  wire v22f0faf;
  wire v230f485;
  wire v231160e;
  wire a6b8e0;
  wire v230ec1c;
  wire v23fc6a2;
  wire v2308d83;
  wire v230eafa;
  wire v22f7861;
  wire v23139ef;
  wire v22ec0d9;
  wire v23fc709;
  wire v23fbdfc;
  wire v23fc0c1;
  wire v22fc9cd;
  wire v23934d5;
  wire v22f586f;
  wire v1aad323;
  wire v22fe924;
  wire v23fb743;
  wire v22f7b83;
  wire v22ee884;
  wire v2312c3c;
  wire v22f0bb4;
  wire v23fba0f;
  wire v22f25e6;
  wire v2393b93;
  wire v22fa002;
  wire v15070f7;
  wire v23fc243;
  wire v23fc583;
  wire v22ec53b;
  wire v23fc3f7;
  wire v22fe73f;
  wire v8ebd5d;
  wire v22edbe0;
  wire v23fc356;
  wire v23fc9ef;
  wire v85f4fd;
  wire v22fea74;
  wire v22f56ce;
  wire v22fe01a;
  wire v230cdf2;
  wire v230ae9d;
  wire v2301e8c;
  wire v22fc477;
  wire v23129d7;
  wire v23015a7;
  wire v95adb3;
  wire v230094d;
  wire v23fbba4;
  wire v22f2aa4;
  wire v23fca61;
  wire v22f1943;
  wire v22f6683;
  wire v2305d69;
  wire v23f4067;
  wire v23081eb;
  wire v230a117;
  wire v2302973;
  wire v230d2d1;
  wire v23f4254;
  wire v22f70a0;
  wire v23fc526;
  wire v22fe948;
  wire v231164b;
  wire v23fcd38;
  wire v22f542d;
  wire v23018f2;
  wire v230709c;
  wire v23f022a;
  wire v22eaafd;
  wire v22fa195;
  wire v230158e;
  wire v23fb4bd;
  wire v22f8e5d;
  wire v23fb968;
  wire v22f39a8;
  wire v23fcc8c;
  wire v23f80c1;
  wire v22f4e64;
  wire a83396;
  wire v22f9b0c;
  wire v22f969f;
  wire v231345a;
  wire v12cd6a1;
  wire v22f4faf;
  wire v230cfba;
  wire v230e4ae;
  wire v22feae3;
  wire v22f3e14;
  wire v22f0139;
  wire v2392d52;
  wire v23f21e5;
  wire v23f617e;
  wire v23fb109;
  wire v23f59e0;
  wire v22f099c;
  wire v23928cd;
  wire f40aac;
  wire v23fc228;
  wire v22f1b11;
  wire v23fbf26;
  wire v23fc56f;
  wire v23fbb8b;
  wire v23fbd42;
  wire v23fb8fa;
  wire v239383b;
  wire v22fe6c8;
  wire v22f5a08;
  wire v23f3b1e;
  wire v191b041;
  wire v22fbf28;
  wire v2311c26;
  wire v23fbb7e;
  wire v22f2c30;
  wire v23fc732;
  wire v2303c9e;
  wire v23043af;
  wire v23fc70c;
  wire v2303dcb;
  wire v23f024e;
  wire v23f57a2;
  wire v23fb873;
  wire v22eed4c;
  wire v23f87b7;
  wire v230abfb;
  wire v230e547;
  wire v22f8aeb;
  wire v230f2f5;
  wire v230faaf;
  wire v22ef725;
  wire v230ebff;
  wire v230d793;
  wire v230c124;
  wire v22eef57;
  wire v2300271;
  wire v2306fb7;
  wire v23f408c;
  wire v22f732c;
  wire v99ce01;
  wire v230dce6;
  wire v23f1e1b;
  wire v230c93a;
  wire v23fb2ea;
  wire v1e83f7c;
  wire v23fcb76;
  wire v2310b6a;
  wire v2309c14;
  wire v23fb9dc;
  wire v23f35c4;
  wire v23fb1b4;
  wire v22f7e16;
  wire v2302c08;
  wire v23fb473;
  wire v23fb4d1;
  wire v22edee1;
  wire v2304049;
  wire v2392833;
  wire v23fc8ef;
  wire v23f730d;
  wire v2304ee5;
  wire v22f26fc;
  wire v2305d92;
  wire v23fcb31;
  wire v22f603b;
  wire v23fc11e;
  wire v22f3643;
  wire v22ecfe0;
  wire v230283f;
  wire v2303b4f;
  wire v12cc72f;
  wire v2312392;
  wire v2309126;
  wire v22f9690;
  wire v23f89df;
  wire v22fca28;
  wire v23fcd6b;
  wire v2304669;
  wire v2313405;
  wire a04dcc;
  wire v23f5bf7;
  wire v22f41ab;
  wire v22f082c;
  wire v23fc050;
  wire v230522a;
  wire v22f4f40;
  wire v23fc853;
  wire v23fc90f;
  wire v2302136;
  wire bd9916;
  wire v22f4ace;
  wire v23fcf9b;
  wire v230b913;
  wire v23fcbd3;
  wire v22f4008;
  wire v23fbaef;
  wire v23f1227;
  wire v23fc5d5;
  wire v2391c58;
  wire v22f0326;
  wire v23045e7;
  wire v22f61cc;
  wire v22fb3df;
  wire v230c5ad;
  wire v23fb217;
  wire v230ee28;
  wire v23fb84f;
  wire v23f8cd3;
  wire v22fe96a;
  wire v23fbadc;
  wire v23fb8a8;
  wire v2311aad;
  wire v22fe144;
  wire v23f6a76;
  wire v23fc82c;
  wire v230a2ae;
  wire v22f3982;
  wire a4e378;
  wire v22f95c8;
  wire v2302b44;
  wire v22fb6bf;
  wire v22f9ae9;
  wire v23fbacc;
  wire v22efda2;
  wire v23fc96e;
  wire v22eb6ba;
  wire v22ed751;
  wire v23f619e;
  wire v23f761c;
  wire v22fcd7c;
  wire v22fa156;
  wire v1aad31f;
  wire b9c9d4;
  wire v23fbc77;
  wire v22f8af0;
  wire v22f7800;
  wire v2310516;
  wire f405d5;
  wire v230ef7c;
  wire v22f9894;
  wire v22f7159;
  wire v22ecc25;
  wire v22fcceb;
  wire v2302933;
  wire v23fc1a3;
  wire v2305a1c;
  wire v22eb3c2;
  wire v22f5d1e;
  wire v23fcefd;
  wire v22ed267;
  wire v23f8d76;
  wire v23f8913;
  wire v230d0a3;
  wire v230646f;
  wire v230faec;
  wire v22f5a2a;
  wire v23f01d2;
  wire v23f0030;
  wire v2308d66;
  wire v2308be5;
  wire v23f6bf0;
  wire v23f8274;
  wire v2311fc9;
  wire v22fecf2;
  wire v22f518e;
  wire v23f9682;
  wire v23f374e;
  wire v2303edc;
  wire v23059e1;
  wire v23fc469;
  wire v23f7b32;
  wire v23096e7;
  wire bda69e;
  wire v230dacd;
  wire v22eeecc;
  wire c0084f;
  wire v22f7319;
  wire v23f8c92;
  wire v230c0b4;
  wire v238ab71;
  wire v22fc56c;
  wire v23f6f06;
  wire v23fbad9;
  wire v2302f12;
  wire v12ce4ac;
  wire v22f88c3;
  wire v23fa005;
  wire v895d68;
  wire v22fe2ae;
  wire v23fbe76;
  wire v23facd7;
  wire v9bcad3;
  wire v23f441d;
  wire v22f5d73;
  wire v23fcb17;
  wire v22f5437;
  wire v230c872;
  wire v23064ad;
  wire v2301bdb;
  wire v2303e23;
  wire v23fb138;
  wire v22f52d4;
  wire v230cbc4;
  wire v22f753f;
  wire v230e9ea;
  wire v230932e;
  wire v23fca19;
  wire v22efdb1;
  wire v23fcf25;
  wire v23fbb10;
  wire v191b155;
  wire v23fcdac;
  wire v23f7898;
  wire v8a7512;
  wire v22ee323;
  wire v239233a;
  wire v22fa4df;
  wire v239288d;
  wire v23f2fd2;
  wire v22f8b41;
  wire v22eef9f;
  wire v23fcff0;
  wire v230d5f4;
  wire v22ef0fe;
  wire v17a34f8;
  wire v23f0eeb;
  wire v22f8603;
  wire v231032d;
  wire v22ef769;
  wire v23114d2;
  wire v2391b6c;
  wire v23fb8e5;
  wire v230a730;
  wire v230345b;
  wire v23fc089;
  wire v23fbf0b;
  wire v13afc0b;
  wire v23fce54;
  wire v23fb85a;
  wire v23fcffb;
  wire v23fb18d;
  wire v1aadf33;
  wire v2305cc1;
  wire v22ede0b;
  wire v23fc898;
  wire v12cd6a2;
  wire v23057ba;
  wire v2300aa8;
  wire v22fd666;
  wire v23fc994;
  wire v2307a72;
  wire v23f6843;
  wire v230ad1e;
  wire v23082fe;
  wire v2310aee;
  wire v23f4451;
  wire v23f8d1a;
  wire v23fce7d;
  wire v23034f8;
  wire v23925e9;
  wire v22efc7f;
  wire v23fb615;
  wire v231232b;
  wire v23fc44a;
  wire v23fc140;
  wire a1fda8;
  wire v22f6124;
  wire v23fca95;
  wire v2301312;
  wire v22f3692;
  wire v22f39af;
  wire v22f1bec;
  wire v22edaad;
  wire v2310430;
  wire v22ee339;
  wire v23f4a16;
  wire v22f792a;
  wire v23126c9;
  wire v23fc9d3;
  wire v23fcedb;
  wire v23fc034;
  wire v230ed7d;
  wire v23fc1a2;
  wire v22f8da4;
  wire a4c16b;
  wire v23f30b2;
  wire v23fbc6a;
  wire v22f2884;
  wire v23fce0d;
  wire v22ff066;
  wire v23f35d5;
  wire v22f2a4f;
  wire v22f3bb0;
  wire aa26cc;
  wire v2312a93;
  wire v23044e1;
  wire v1aae206;
  wire v22fc8fb;
  wire v23fc366;
  wire v23fc498;
  wire v230f1c8;
  wire v23fc2b8;
  wire v23f5055;
  wire a1ba8b;
  wire v23fc230;
  wire v23916ef;
  wire v22fb790;
  wire v22f8d2f;
  wire v22ee957;
  wire v230f654;
  wire v22f50bf;
  wire v2309310;
  wire v2391bc1;
  wire v2306996;
  wire v2392a3a;
  wire v22fe831;
  wire v23fc5f8;
  wire v230c20b;
  wire v230704c;
  wire v23fd017;
  wire v23fbaa7;
  wire v230f4a8;
  wire v23f0135;
  wire v22fdf5b;
  wire v2310d74;
  wire v230df15;
  wire v22fda30;
  wire v2312fc7;
  wire v230011a;
  wire v22f5109;
  wire v22f7c09;
  wire v22ef45e;
  wire bdc4e2;
  wire v8f8537;
  wire v2307375;
  wire v23f4a00;
  wire v22efd4a;
  wire v230bae0;
  wire v230c03a;
  wire v2393775;
  wire v23f5787;
  wire v23fb8e3;
  wire v22ff13f;
  wire v22ec89f;
  wire v22f227e;
  wire v23920d8;
  wire v230b756;
  wire v22f53df;
  wire v22ed148;
  wire v23006e9;
  wire v22f6358;
  wire v23fcbe9;
  wire v23fcedf;
  wire v23f592d;
  wire v2391e0c;
  wire v230a226;
  wire v239313a;
  wire v22f690f;
  wire v8a34ca;
  wire v150730e;
  wire v23fc78a;
  wire v2306844;
  wire v230d6b6;
  wire b23404;
  wire v23fc88b;
  wire v23f47e1;
  wire v23fcf22;
  wire v23fcdcd;
  wire v22ec0de;
  wire v230199e;
  wire v22f8da3;
  wire v230f933;
  wire v22ff613;
  wire v23fba98;
  wire v2312e57;
  wire v23fcb0f;
  wire v22f3324;
  wire v22f94b6;
  wire v22fe32b;
  wire v23f2713;
  wire v22f53d4;
  wire v23f22d2;
  wire v23f2768;
  wire v2301cc6;
  wire v23fb200;
  wire v23f38a5;
  wire v22fa3df;
  wire v22f6219;
  wire v230df7b;
  wire v22f8b43;
  wire v1aad9a6;
  wire v23f1e72;
  wire v2393723;
  wire v22ecb9d;
  wire v230c649;
  wire v23044e2;
  wire v23111ee;
  wire v23f850a;
  wire v22f66cf;
  wire v23f7db2;
  wire v22fa371;
  wire v22f15ef;
  wire v22f6b7d;
  wire v23f2c65;
  wire v23fc02d;
  wire v22f0f36;
  wire v23fc61d;
  wire v23f78df;
  wire v230cc95;
  wire v23fc638;
  wire v23fcca2;
  wire v22eccde;
  wire v1b8771f;
  wire v22fb36e;
  wire v22f58cd;
  wire v2307cdf;
  wire v2311504;
  wire v23080f9;
  wire v23f60e8;
  wire v23fc32f;
  wire v22fb4a6;
  wire v22fa9ce;
  wire v22efe2f;
  wire v22f0c6d;
  wire v22fe675;
  wire v1e845a7;
  wire v230713e;
  wire v23fcbd8;
  wire v22ec1a8;
  wire v230c1e1;
  wire v22ec2e6;
  wire v230e0d6;
  wire v22fb068;
  wire v23fcfba;
  wire v231024c;
  wire v22efa8c;
  wire v239407e;
  wire v990272;
  wire v22f639a;
  wire v23f532f;
  wire v2392222;
  wire v22f9b30;
  wire v22ec012;
  wire v23fcb8f;
  wire v22eaf81;
  wire v2305bf5;
  wire v1506ff4;
  wire v22ff5bd;
  wire v23f4c5b;
  wire v23fbff9;
  wire v23f232d;
  wire v23109e3;
  wire v23fb078;
  wire v22fee33;
  wire v22ef094;
  wire v23fb843;
  wire v2312e50;
  wire v22f0646;
  wire v15071a6;
  wire v23f4a48;
  wire v2305866;
  wire v23fbb9c;
  wire v23fcfce;
  wire v23f62c2;
  wire v22f856d;
  wire v22f8e2f;
  wire v23fc320;
  wire v23fc98c;
  wire v230ccd6;
  wire v22fdbdb;
  wire v2301818;
  wire v23f66fd;
  wire v23075bd;
  wire v23130ea;
  wire v23fbb44;
  wire v13afad7;
  wire v23fc92d;
  wire v23f3d14;
  wire v239214a;
  wire v23fc197;
  wire v23127b2;
  wire b9c9cc;
  wire v23f836b;
  wire v22f0ad8;
  wire v23fcabe;
  wire v230a5f5;
  wire v22fd7ee;
  wire v22f4321;
  wire v23fc99c;
  wire v23f9c04;
  wire v22faf41;
  wire v22f53b1;
  wire v230a36f;
  wire v230124d;
  wire v22ecb49;
  wire v22ec992;
  wire v23fb5d8;
  wire v230fac9;
  wire v22f4b44;
  wire v230716c;
  wire v2310a55;
  wire v23f4a07;
  wire v23fca46;
  wire v239174f;
  wire v23125a2;
  wire v23fcc45;
  wire v22fa987;
  wire v22ee665;
  wire v22ed674;
  wire v2301a42;
  wire v22fde18;
  wire v22ed12a;
  wire v1506ec2;
  wire v22f88f9;
  wire v23104c1;
  wire v23f3ac8;
  wire v22f7289;
  wire v2393bcf;
  wire v230c480;
  wire v22f1153;
  wire v23fccbc;
  wire v23fcd0b;
  wire v191ad59;
  wire v23fa0bf;
  wire v22f3f32;
  wire v23fbc96;
  wire v22f082f;
  wire v23fcbed;
  wire v2302b3e;
  wire v23fc318;
  wire v2392d97;
  wire v23f66e6;
  wire v2309ff9;
  wire v23fc3ff;
  wire v2304ad5;
  wire v23fb709;
  wire v22f8fa4;
  wire v23052a8;
  wire v2306f84;
  wire v2312c77;
  wire v2311675;
  wire v23faa23;
  wire v22f3d00;
  wire v23f4808;
  wire v12cda0a;
  wire v23113d2;
  wire v22fb465;
  wire v2305c78;
  wire v231140b;
  wire v23f482d;
  wire v22f09c5;
  wire v22ed4c6;
  wire v2308235;
  wire v23fbfe2;
  wire v22f10cc;
  wire v22fc7e6;
  wire v230e32f;
  wire v22f7c6f;
  wire v230ec2b;
  wire v23f63dc;
  wire v22fd8c5;
  wire v22ede9f;
  wire v23fbd33;
  wire v230979d;
  wire v2313595;
  wire v22f7d33;
  wire v23fbff0;
  wire v2393064;
  wire v22f6719;
  wire v22f0aea;
  wire v22fd372;
  wire v23095b3;
  wire v2309cb0;
  wire v23fcbca;
  wire v23fcf7c;
  wire v23fc820;
  wire v22f0dc9;
  wire v2300487;
  wire v23fbc83;
  wire b0fe84;
  wire v23fc1ee;
  wire v23087f2;
  wire v2300cbb;
  wire v23fb1e1;
  wire v23fbfa7;
  wire v22f3dab;
  wire v22f76c6;
  wire v2300c06;
  wire v2311d04;
  wire v23fb667;
  wire v23f03d2;
  wire v23fbf0e;
  wire v2306625;
  wire v23fd026;
  wire v230278d;
  wire v23fc8cf;
  wire v23fcb03;
  wire v1e84183;
  wire v23fbf55;
  wire v22fb28f;
  wire v22f609f;
  wire v23fc235;
  wire v23fc570;
  wire v23fcfd6;
  wire v23f4634;
  wire b9d061;
  wire v22f7110;
  wire v22ef9f7;
  wire v23fc808;
  wire v2392f11;
  wire ba4552;
  wire v23fc43e;
  wire v230b5b8;
  wire v23fcd7c;
  wire v23fca90;
  wire v23f6729;
  wire v2303270;
  wire v22f7758;
  wire v22ede8c;
  wire v23045fa;
  wire v23f6739;
  wire v22eb665;
  wire v2309d09;
  wire v23fc2a0;
  wire a1ff39;
  wire v23027bf;
  wire v22fcb45;
  wire v22fce0a;
  wire v230eb9e;
  wire v2300621;
  wire v23fcdd9;
  wire v23fcb1a;
  wire v23f2dd4;
  wire v22fb373;
  wire v2310ab0;
  wire b52881;
  wire v23f839a;
  wire v230a742;
  wire v230e262;
  wire v230a71c;
  wire v23fc3c3;
  wire v23f23f1;
  wire v23fc9c8;
  wire v22ebbf1;
  wire v22f5d87;
  wire v22f4bb5;
  wire v2392836;
  wire v22ed10d;
  wire v2312948;
  wire v22f4a40;
  wire v22f84f8;
  wire v22eb6ee;
  wire v23fca15;
  wire v23fcfb7;
  wire v2308786;
  wire v2310731;
  wire v23fcca1;
  wire v22ec64d;
  wire v23f4f43;
  wire v22eb8b6;
  wire v230cc4c;
  wire fc9434;
  wire v230f256;
  wire v22f3f68;
  wire v22eb2a2;
  wire v23fbc94;
  wire v23fc3f1;
  wire v23f7853;
  wire v23022d0;
  wire v23fc060;
  wire v2391982;
  wire v22ed03d;
  wire b6c104;
  wire v22ee5fb;
  wire v230c849;
  wire b9d041;
  wire v2313279;
  wire v230cfa5;
  wire v239300d;
  wire v23fbea4;
  wire v23fb1a0;
  wire v23f7f02;
  wire v2301f5c;
  wire v230e966;
  wire v23fba9f;
  wire v230272d;
  wire v23fc040;
  wire v2302179;
  wire v2303415;
  wire v23f25c8;
  wire v22f8d8e;
  wire v23f4491;
  wire v23fc315;
  wire v22ed6bc;
  wire v2303996;
  wire a51d7a;
  wire v230b161;
  wire v22ed984;
  wire v23084cf;
  wire v22ec801;
  wire v2392f21;
  wire v230edde;
  wire v23f6155;
  wire v22f83cf;
  wire v230ae09;
  wire v23f7f77;
  wire v23f0625;
  wire v23f7148;
  wire v2303978;
  wire v22fe992;
  wire v23f81cf;
  wire v22fa766;
  wire v12cddb2;
  wire v22f8b9c;
  wire v23fb501;
  wire v22f78de;
  wire v2391f2b;
  wire v22fea3e;
  wire v23f95ef;
  wire v23f84b2;
  wire v2300cb6;
  wire v22f11fe;
  wire v23fc256;
  wire v23fb8cb;
  wire v23f3955;
  wire v22efdfe;
  wire v23fc25e;
  wire v23f1ad7;
  wire v23f6283;
  wire v230448f;
  wire v22eefe2;
  wire v22fbe82;
  wire v230fa1a;
  wire v2346b8a;
  wire v22f05a9;
  wire v22f9f44;
  wire v230f554;
  wire v23fcd33;
  wire v230a562;
  wire v22f2114;
  wire v230389f;
  wire v1507437;
  wire v23fc5e9;
  wire v23fba73;
  wire v230eac0;
  wire v2307020;
  wire v2306d33;
  wire v230379f;
  wire v191a909;
  wire v2301bb5;
  wire v23074c9;
  wire v23f8976;
  wire v22fcea7;
  wire v23fc9f3;
  wire v1aae262;
  wire v23fce81;
  wire v23f1515;
  wire v22f2a76;
  wire v23f24c5;
  wire v22f4e1f;
  wire v23fc605;
  wire v22fb450;
  wire v230d709;
  wire v2312526;
  wire v23f32a6;
  wire v230916d;
  wire v22f55fa;
  wire v23fc316;
  wire v23fc2db;
  wire v23fcecc;
  wire v22fcc78;
  wire v1aad46b;
  wire v23f8ddb;
  wire e1e258;
  wire v23fbeb5;
  wire v230afed;
  wire v23f2380;
  wire v2306f2e;
  wire v23fba39;
  wire v2302a77;
  wire v23f99bc;
  wire v22f0de4;
  wire v23120b1;
  wire v23fbe06;
  wire v2306fae;
  wire v23fc70f;
  wire v22ecab2;
  wire v22edd4c;
  wire v23fcdbd;
  wire b20f9d;
  wire v230e6ad;
  wire v23fb476;
  wire v21b35f9;
  wire v2300755;
  wire v23fc4a4;
  wire v22ed878;
  wire v230ec10;
  wire v23fc71d;
  wire v23fbfd0;
  wire v2305338;
  wire v230910b;
  wire v230806a;
  wire v23fce71;
  wire v191ab5f;
  wire v22f197e;
  wire v22f0add;
  wire v2310a63;
  wire a1fcbb;
  wire v230b981;
  wire v23fcd6a;
  wire v23fb4a0;
  wire v22fe34f;
  wire v22f803d;
  wire v2302d3c;
  wire v23fbbf0;
  wire v230502a;
  wire v2304494;
  wire v22fc4d3;
  wire b9c8dc;
  wire v23fced7;
  wire v2301505;
  wire v230f2d1;
  wire v23fc7d5;
  wire v23f391e;
  wire v23fc739;
  wire v9f4f45;
  wire v23fb978;
  wire v22f0d22;
  wire v230f9c8;
  wire b60876;
  wire v23fc41e;
  wire v230aca2;
  wire v23fba85;
  wire v2305dde;
  wire v23fc7c8;
  wire v2392b3d;
  wire v230a7c3;
  wire v23fcaec;
  wire v23fc6f0;
  wire v1e84b3e;
  wire v23938ff;
  wire bd9e8b;
  wire v2312142;
  wire v22f05a7;
  wire v23fc585;
  wire v230ae24;
  wire v23f8a9d;
  wire v22f99ee;
  wire v230153d;
  wire v992f98;
  wire v23f2d8c;
  wire v23014fb;
  wire v2306414;
  wire v22f8543;
  wire v23efac1;
  wire v1aae294;
  wire v23128a1;
  wire v230e509;
  wire v22fd3f9;
  wire v23fc9f8;
  wire v23fc931;
  wire v23fb96b;
  wire v23fb4af;
  wire v12cd4f6;
  wire v23fa392;
  wire v230774f;
  wire v23f7b0a;
  wire v23fbba5;
  wire v231251d;
  wire v23fcc64;
  wire v23f8da8;
  wire v22f1762;
  wire v8a894a;
  wire v2304ea9;
  wire v23fa8d8;
  wire v23fc01a;
  wire v23fa492;
  wire v2302365;
  wire v22f6741;
  wire v23fbcce;
  wire v23f4364;
  wire v23fb4a1;
  wire v23f6f49;
  wire v230e8b8;
  wire v23f2508;
  wire b9d02f;
  wire v12cd69f;
  wire v22f11f6;
  wire v22edfa7;
  wire v2305b58;
  wire v2311656;
  wire v22f0b56;
  wire v23fce15;
  wire v23fc260;
  wire v23920aa;
  wire v23013a2;
  wire v22edec8;
  wire v22f6a3a;
  wire v13aff46;
  wire v2312b5a;
  wire v22fda85;
  wire e1cfe5;
  wire v23fcb68;
  wire v23f5ba9;
  wire v22f839c;
  wire v23f3e44;
  wire v23f1e3f;
  wire v230197e;
  wire v23fc9a5;
  wire v2311eaa;
  wire v22f721f;
  wire v230dffa;
  wire v2308a0c;
  wire v22f3101;
  wire v23fc7e6;
  wire v23fbfc9;
  wire v22f8aba;
  wire v22f60dd;
  wire v230f9d5;
  wire v23f8a41;
  wire v23fc4a5;
  wire v23fbf67;
  wire v230f1ae;
  wire v22f5110;
  wire v22fe59c;
  wire v23fa9d0;
  wire v23fb636;
  wire v22ed236;
  wire v1aad609;
  wire v230f693;
  wire v22f6e67;
  wire v230287e;
  wire v23fc023;
  wire v230adb7;
  wire v23135ca;
  wire v22fb511;
  wire v2312067;
  wire v230c876;
  wire v932767;
  wire v23f8bef;
  wire v2303674;
  wire v22ef0c8;
  wire v23fccd6;
  wire v23fa175;
  wire v22f6f5c;
  wire v22f9f33;
  wire v2307320;
  wire v23fb81d;
  wire v22fca36;
  wire v23fc038;
  wire v22f0f76;
  wire v22faa66;
  wire v23fc867;
  wire v23053bd;
  wire v23024ed;
  wire v2306bed;
  wire v23f1726;
  wire v230aa0b;
  wire v2308669;
  wire v23fc364;
  wire v230334d;
  wire v23fcfe8;
  wire v22f5d5e;
  wire v22eaafa;
  wire v22fa415;
  wire v23107f9;
  wire v22f231d;
  wire v2306d26;
  wire v230a67e;
  wire v23f2f45;
  wire v23f1207;
  wire v230f370;
  wire v230b1ac;
  wire v22f35f5;
  wire v23fcc67;
  wire v22fc893;
  wire v23fcfad;
  wire v23fc75c;
  wire v230c041;
  wire v23055d4;
  wire v22ed5e6;
  wire v23fbdfe;
  wire v22eafea;
  wire v23fb90c;
  wire v23070cf;
  wire v23fcd4b;
  wire v23f7ce8;
  wire v22ff9c5;
  wire v22fe1ad;
  wire v23f2b69;
  wire v23043b7;
  wire v23090fd;
  wire v2393116;
  wire v191ae6a;
  wire v23fc7ee;
  wire v23fc086;
  wire v23f7dbe;
  wire v2305bbb;
  wire v22f42bd;
  wire v22ee660;
  wire v23fbf24;
  wire v22f34c1;
  wire b6f86d;
  wire f40cd3;
  wire v22fb7a5;
  wire v22f98fd;
  wire v23f8c0b;
  wire v22ff969;
  wire v23fb3a3;
  wire v230d99c;
  wire v22fffe4;
  wire v23041ee;
  wire v239350a;
  wire v22f9bed;
  wire v23fc7b7;
  wire c173c8;
  wire v230f70f;
  wire v22fe81e;
  wire v23016d9;
  wire v22f84a0;
  wire v23070dd;
  wire v23f6e78;
  wire v23f88a9;
  wire v23fce9e;
  wire v2309282;
  wire v22f640a;
  wire v23f54a0;
  wire v2304452;
  wire v23fc9fb;
  wire v23fbf74;
  wire v22eb265;
  wire v2308abb;
  wire v22f6463;
  wire v23fba18;
  wire v23fca7e;
  wire v23fb938;
  wire v23015c2;
  wire a7482d;
  wire v2301652;
  wire v2310ffa;
  wire v23fba04;
  wire v1aae99f;
  wire v23fc785;
  wire v23040a8;
  wire v23f673b;
  wire v230b1ab;
  wire v23fcd45;
  wire v95aaca;
  wire v23052b7;
  wire v22f1f9f;
  wire v23fbccc;
  wire v23f5470;
  wire v23f2324;
  wire v2308e2e;
  wire v23fcf83;
  wire v23fbb95;
  wire v23f4cb5;
  wire v23fbe96;
  wire v2308b2f;
  wire v22f0128;
  wire v22f985c;
  wire v230ef5e;
  wire v23fcb0a;
  wire v2300b6b;
  wire v899296;
  wire v230ca2b;
  wire v23fb63c;
  wire v23f5ad6;
  wire v23f659c;
  wire v1b87690;
  wire v230fab4;
  wire v22f5d52;
  wire v22eea17;
  wire v22fafe5;
  wire v22f3b02;
  wire v2303199;
  wire v23fc468;
  wire a33e98;
  wire v230708b;
  wire v22f2822;
  wire v22feee5;
  wire v22ecdfe;
  wire v2306fdd;
  wire v230a7a5;
  wire v230b2a4;
  wire v230e95c;
  wire v2307aad;
  wire v2307e4f;
  wire v22f35fa;
  wire v9180fe;
  wire v23fcf54;
  wire v191b186;
  wire v23fcd5d;
  wire aa8bd6;
  wire v23fc850;
  wire v2305c2e;
  wire v230835d;
  wire v22ecff3;
  wire v22efdf3;
  wire v2311dc5;
  wire v2301306;
  wire v22f5efe;
  wire v2304a1e;
  wire v22fe740;
  wire v22fba3f;
  wire v22f2363;
  wire v230b23c;
  wire v2302831;
  wire v230cbdd;
  wire v23f353e;
  wire v22fa502;
  wire v22f7152;
  wire v23fc844;
  wire v230fe71;
  wire v22fd86e;
  wire v23fd050;
  wire v22f881b;
  wire v22f1ee5;
  wire c086a6;
  wire v22edcfc;
  wire v23124cc;
  wire v22f5834;
  wire v2311e39;
  wire v23fc99a;
  wire v23028f6;
  wire v22f8012;
  wire v230e0d5;
  wire v23fc969;
  wire v2307632;
  wire v230a919;
  wire v230a70a;
  wire v23fb12f;
  wire v2311302;
  wire v22eaee7;
  wire v231261b;
  wire v2312a90;
  wire v23fcb7e;
  wire v230e7e4;
  wire v230f713;
  wire v230ff52;
  wire d97946;
  wire v22f3068;
  wire v12cd9b5;
  wire v22f2f33;
  wire v2309023;
  wire v2304b5d;
  wire v230c0b2;
  wire v23fb4d3;
  wire v23fbe1b;
  wire v230eeb6;
  wire v9e3170;
  wire v23fb7d1;
  wire v23fb856;
  wire v22fa027;
  wire v23078cd;
  wire v230ca2e;
  wire v22f791d;
  wire v22f18f3;
  wire v22fb6df;
  wire v22eb856;
  wire v23f96d0;
  wire v23f33c7;
  wire v23f669d;
  wire v22f69ed;
  wire v22fc588;
  wire v22f7c32;
  wire v23f5767;
  wire v22fbd02;
  wire v22fd00f;
  wire v22fef20;
  wire v23fb236;
  wire v23002e0;
  wire v22fe300;
  wire v23f50ec;
  wire v22fabd2;
  wire v2310238;
  wire v22ef2be;
  wire v2313351;
  wire v230f7ff;
  wire v22eea5b;
  wire v22fd9a5;
  wire v23f2843;
  wire v23f1d35;
  wire v23045fb;
  wire v2300f96;
  wire v23064ff;
  wire v22fe428;
  wire v22eb599;
  wire v23f3f73;
  wire e1e722;
  wire v230886c;
  wire v2300bb5;
  wire v23fc67f;
  wire v22f4627;
  wire a7dd55;
  wire v22f50f0;
  wire v22f8f3d;
  wire v23fbc55;
  wire v22f15fd;
  wire v23fcaeb;
  wire v2301eb1;
  wire v2310108;
  wire v2313144;
  wire v23077dc;
  wire v22f165f;
  wire v22f8ce6;
  wire v22f3385;
  wire v191b1ba;
  wire v22fef65;
  wire v2312e80;
  wire v22ed999;
  wire v22f8c6b;
  wire v23023aa;
  wire v22f16d8;
  wire v23f416b;
  wire v23fbc1d;
  wire v23fc3c9;
  wire v23f22a1;
  wire v23fb122;
  wire v23fb8c1;
  wire v22f5f1c;
  wire v23f6250;
  wire v23fab18;
  wire v2310782;
  wire v1506f02;
  wire v23f4e25;
  wire v23102bf;
  wire v230dbc9;
  wire v22efa5e;
  wire v23fc7f0;
  wire v230de92;
  wire v23022b3;
  wire v22fc23d;
  wire v191ae7d;
  wire v23f9465;
  wire v23fc52d;
  wire v23fa77d;
  wire v23f31d6;
  wire v2303075;
  wire a1b802;
  wire v230ed27;
  wire v22efb25;
  wire v12ce0d0;
  wire v23928d0;
  wire v22ed48e;
  wire v230c84d;
  wire v9a3d0c;
  wire v22f0c5f;
  wire v22fa299;
  wire v23faa0a;
  wire v22ebebe;
  wire v23fba16;
  wire v23fc26c;
  wire v23fb0a1;
  wire v1aad65a;
  wire v22ffdc9;
  wire v230eed5;
  wire v23f437d;
  wire v2301190;
  wire v23fb52e;
  wire v230984f;
  wire v23089f7;
  wire v22fb009;
  wire v22efceb;
  wire v23f5fd9;
  wire v231182b;
  wire v230251b;
  wire v23fcdb6;
  wire v23fbad7;
  wire v23fcc43;
  wire v23fcfda;
  wire v22f97c3;
  wire v23083c1;
  wire v23130b0;
  wire v23093e2;
  wire v23fbc9f;
  wire v22ebe20;
  wire v22fa6b2;
  wire v106ae5a;
  wire v22ef242;
  wire v22eebd6;
  wire v22f3b8c;
  wire v23fc39f;
  wire v22f8824;
  wire v1506a62;
  wire v23fba0a;
  wire v23fc60e;
  wire v22febe1;
  wire v23fb5e3;
  wire v23fcac2;
  wire v22fa9be;
  wire v1aad481;
  wire v23128ab;
  wire v23fbd1a;
  wire v23f50e0;
  wire v22f1e0b;
  wire v23fc7ef;
  wire v2300df6;
  wire v23f6588;
  wire v23fc6ef;
  wire v23fbec5;
  wire v9c8a7f;
  wire v2305a26;
  wire v2307fcd;
  wire v22f825a;
  wire v230d1de;
  wire v22f1376;
  wire v1aad38a;
  wire v22f8ed1;
  wire v23fcd6c;
  wire v23060bb;
  wire v23fb813;
  wire v22edb40;
  wire v230b08b;
  wire v2303ae3;
  wire v2300b7b;
  wire v23f3958;
  wire v22fa5fd;
  wire v23027cd;
  wire v22fc1e9;
  wire v23fbcca;
  wire v23fc18b;
  wire v22fec1c;
  wire v2308b02;
  wire v22efbd5;
  wire v22fd2ac;
  wire v22ffcec;
  wire v22ef116;
  wire v230b1a3;
  wire v2307eee;
  wire v23fceec;
  wire v23126c6;
  wire v2300c47;
  wire v191ace8;
  wire v22f5039;
  wire v23046b5;
  wire v22f01c5;
  wire v22f4d74;
  wire v22f7144;
  wire v2308455;
  wire v22fd655;
  wire v1aadf17;
  wire v23f58f9;
  wire v2310bd4;
  wire v22fc963;
  wire v2392aaa;
  wire v23f2d60;
  wire v22fdf70;
  wire v230296a;
  wire v230075e;
  wire v23f6f88;
  wire v23fbf93;
  wire v23fc7ba;
  wire v230a435;
  wire v23fb436;
  wire v230e635;
  wire v22ede6c;
  wire v23fc5ad;
  wire v23f3af2;
  wire v230cdc7;
  wire v2309ae3;
  wire v23094a1;
  wire v230e880;
  wire v22fabaf;
  wire v23fc2d8;
  wire v22fbc4e;
  wire v230884d;
  wire v231086d;
  wire v23f7700;
  wire v23faa78;
  wire v22ef62d;
  wire v230a434;
  wire v23fc683;
  wire v230cb1f;
  wire v22f3e8d;
  wire v23fbbb2;
  wire v23fcdaa;
  wire v22f0c5d;
  wire v230f974;
  wire v22edf54;
  wire v22f1a26;
  wire v230b1db;
  wire v22ef403;
  wire v2301e25;
  wire v230aa54;
  wire v22f0593;
  wire v230880f;
  wire v22eb6ca;
  wire v23fceb3;
  wire v23fb8c0;
  wire v2312d48;
  wire v230fff1;
  wire v22f4f14;
  wire v2302937;
  wire v23fb1a4;
  wire v23129bb;
  wire v23f8490;
  wire v230d854;
  wire v2309751;
  wire v23fbd1b;
  wire v22eefaf;
  wire v2301be6;
  wire v23fc622;
  wire v23fbb80;
  wire v22fb07c;
  wire v23fcda9;
  wire v22ed1b5;
  wire v12cda51;
  wire v22eeb06;
  wire v22ee36d;
  wire v2301d4e;
  wire v2306a0e;
  wire v23f363f;
  wire v2302fbc;
  wire v23f936e;
  wire v22fdba7;
  wire v23fc068;
  wire v23f7e51;
  wire v2302cfa;
  wire v22f3d67;
  wire v23f493a;
  wire v2300827;
  wire v22ff5af;
  wire v23fb0c0;
  wire v23fc8a5;
  wire v22f9403;
  wire v23fb504;
  wire v22ed1a8;
  wire v2305a37;
  wire a48bb0;
  wire v23013a6;
  wire v23fc3eb;
  wire v22f48ce;
  wire v2301f5d;
  wire v85b90c;
  wire v22eb7cc;
  wire v23fc34b;
  wire v23fbdbe;
  wire v23fba78;
  wire v230d96b;
  wire v23fbb4a;
  wire v2303314;
  wire v23fca6f;
  wire v230ab72;
  wire v2308ced;
  wire v230caac;
  wire v23fc816;
  wire v23f5af8;
  wire v2300de1;
  wire v22f9e08;
  wire v230f403;
  wire v22ff78b;
  wire v2308fb4;
  wire v23fba1c;
  wire v2301511;
  wire v23fd05d;
  wire v23fccdb;
  wire v2306d07;
  wire v2305a12;
  wire v90c400;
  wire v2309599;
  wire v22efc3c;
  wire v22ec921;
  wire v2302e43;
  wire v23f8db0;
  wire v23fbfa0;
  wire v22f54a4;
  wire v22f30df;
  wire v22feec8;
  wire v9e764b;
  wire v2309c28;
  wire v23fb5a4;
  wire v22f0db9;
  wire v23f6635;
  wire v22ebfd3;
  wire v23f4961;
  wire v1aae5da;
  wire c17224;
  wire v23fbaf6;
  wire v23f7db8;
  wire v22ebb79;
  wire v23f73ba;
  wire v230ea9f;
  wire v22f0c1b;
  wire v22f3618;
  wire v23f9593;
  wire v2303b6a;
  wire v23079d8;
  wire v22f72ff;
  wire v23f97de;
  wire v23fc71b;
  wire v23f7561;
  wire v23f6cc2;
  wire ad06d5;
  wire v2312f85;
  wire v23f5eb6;
  wire v22ffd0e;
  wire v22ff45e;
  wire v23f940c;
  wire v23f3f65;
  wire v22ff192;
  wire v22f670f;
  wire v22f0210;
  wire v22f448e;
  wire v23f79e9;
  wire v22ebe5c;
  wire v22f8026;
  wire v23f6bc1;
  wire v22fba41;
  wire v230a9a3;
  wire v23fcf05;
  wire v23fca2a;
  wire v23fc681;
  wire v22f0824;
  wire v22fbdd6;
  wire v23f5b31;
  wire v23fc2e0;
  wire v23fc84b;
  wire v23fa8c8;
  wire v23fcf52;
  wire v22fd5fc;
  wire v230d30a;
  wire v23100c8;
  wire v15071c7;
  wire v23fb6ed;
  wire v22ed335;
  wire v23fb937;
  wire v23fc17c;
  wire v23927e4;
  wire v230049a;
  wire v230dbcc;
  wire v22fc68e;
  wire v22ff3c6;
  wire v2302ba4;
  wire v230eab7;
  wire v23f4cc1;
  wire ad89b5;
  wire v230fe9b;
  wire v23fb6bd;
  wire v22f2849;
  wire v22fc67e;
  wire v22fab21;
  wire v2391655;
  wire v23efec0;
  wire v23fc0a7;
  wire v2300cf1;
  wire v23fbce4;
  wire v23fc0b3;
  wire v22fc0a2;
  wire v22f8839;
  wire v23131a6;
  wire v22ed7b6;
  wire v2307572;
  wire v23fc1be;
  wire v22ed4e1;
  wire v22f1fca;
  wire v230801c;
  wire v23faa94;
  wire v22f0545;
  wire v22f5388;
  wire v23fbab9;
  wire v2306b0a;
  wire v230e086;
  wire v23055d9;
  wire v230c32e;
  wire v230bd1b;
  wire fc90a8;
  wire v2313111;
  wire v23050fb;
  wire v2302abd;
  wire v22fd67c;
  wire v22ffc90;
  wire v22fb43e;
  wire v22fc689;
  wire v23fc6b2;
  wire v22fc493;
  wire v23f6789;
  wire v2309df7;
  wire v23fbe21;
  wire v22f7c9a;
  wire v23fc926;
  wire v230bc8b;
  wire v230230d;
  wire v23058ae;
  wire v23fa997;
  wire v22f8b01;
  wire v23f37c6;
  wire v23fbac1;
  wire v2312acc;
  wire v22f264a;
  wire v23f3fca;
  wire v23fc39c;
  wire v23fcd0f;
  wire v23f7b86;
  wire v23fcb5e;
  wire v12cd93a;
  wire v22f8fc0;
  wire b30f07;
  wire v23080ec;
  wire v9bbf5d;
  wire v23fd069;
  wire v23fbc7e;
  wire v22fb877;
  wire v2301d10;
  wire v22fd3f7;
  wire v23052cc;
  wire v23f987b;
  wire v106a7a3;
  wire v2305055;
  wire v22fba03;
  wire v15072b7;
  wire v22ed907;
  wire v23928f2;
  wire v22f52c3;
  wire v22fcd06;
  wire v23fc841;
  wire v23fbbc0;
  wire v230e7d4;
  wire v22fd8fc;
  wire v230658d;
  wire v23fc58a;
  wire v23fc323;
  wire v2392d6f;
  wire v230b961;
  wire v23f5b39;
  wire v23f3310;
  wire v22f299f;
  wire v22f45ff;
  wire v22ff469;
  wire v23099c5;
  wire v23fceb6;
  wire v23fb14b;
  wire v23fc268;
  wire v23f9bf9;
  wire v230e8a8;
  wire v23fc9dc;
  wire v23fb790;
  wire v22f25fa;
  wire v230f073;
  wire v230cbde;
  wire v230b23b;
  wire v230a3af;
  wire v1e84174;
  wire v23fa1f9;
  wire v230e89f;
  wire v22fe4a1;
  wire v23fbe74;
  wire v23fcb5c;
  wire v23fbd93;
  wire b2aff2;
  wire v22fc10a;
  wire v22fb88e;
  wire v23111c2;
  wire v2312cdf;
  wire v23fbab0;
  wire v22f3be2;
  wire v23064ca;
  wire v106aeed;
  wire v2312007;
  wire v230824c;
  wire v22f0542;
  wire v22eca17;
  wire v22f8ad4;
  wire v22fd0e6;
  wire v12cd3e7;
  wire v230ed6b;
  wire v23f6849;
  wire v23ef95a;
  wire v22febde;
  wire v22f25c5;
  wire v23f22f9;
  wire v2303943;
  wire v23fc997;
  wire v22f1403;
  wire v22f08b7;
  wire v23fb47e;
  wire v2392809;
  wire v230de50;
  wire v23101b0;
  wire v22fbef0;
  wire v23fc58d;
  wire e1d75b;
  wire v22ed1f3;
  wire v2309ab5;
  wire v22f6246;
  wire v22fa105;
  wire v23fc16b;
  wire v22f4667;
  wire v22f28e6;
  wire v22ffab6;
  wire v22eb701;
  wire v23fc8f8;
  wire v23fce10;
  wire v879c1f;
  wire v23098d3;
  wire v2367a5a;
  wire v2307480;
  wire v230d282;
  wire v22f0e84;
  wire v2305782;
  wire v22ff179;
  wire v231185d;
  wire v22fd825;
  wire v22f8463;
  wire v23fb23b;
  wire v22fdcc7;
  wire v23fc34f;
  wire v23015de;
  wire v230c653;
  wire v2301c48;
  wire v23fcd35;
  wire v23fbdf9;
  wire v23fbe15;
  wire v23fc787;
  wire v23f240c;
  wire v23fbb9e;
  wire v23045c3;
  wire v13afbf0;
  wire v22fc908;
  wire v23036a1;
  wire v23f0db7;
  wire v22f2e0c;
  wire v22ed4b0;
  wire v2391dd6;
  wire v230c2ff;
  wire v2309be5;
  wire v230c66e;
  wire v23fd040;
  wire v23fc619;
  wire v23fc81c;
  wire v23fa155;
  wire v23fcd4a;
  wire v23fb5a1;
  wire v22f69cc;
  wire v230c6eb;
  wire v23f4268;
  wire b15a69;
  wire v23f0329;
  wire v22f324f;
  wire v9f009f;
  wire v9ab66e;
  wire v23012c6;
  wire v22f108e;
  wire v22f7b47;
  wire v22f25da;
  wire v23929ca;
  wire v23fcbd0;
  wire v22fb842;
  wire v23fba6c;
  wire v98151e;
  wire v22fdc80;
  wire v230c437;
  wire v23fc334;
  wire v23f7a92;
  wire v22f39a5;
  wire v23f8d64;
  wire v22eb16b;
  wire v23f1e1a;
  wire v191aa89;
  wire v22f129b;
  wire v23fcd30;
  wire v2392d9f;
  wire v22eaee8;
  wire v23f72e4;
  wire v23f1974;
  wire v22ebc86;
  wire v22fa821;
  wire v23fc556;
  wire v2391aa0;
  wire v22f181c;
  wire v22ee247;
  wire bd7786;
  wire v23f3dc2;
  wire v23fcb1f;
  wire v23fc19a;
  wire v2309c07;
  wire v22fbc47;
  wire v23fbe2a;
  wire v2307dae;
  wire v23fcb71;
  wire f40c98;
  wire v2308f5d;
  wire v2305660;
  wire v23f9dd8;
  wire v22f7ce8;
  wire v23fc4ef;
  wire v23fc517;
  wire v106af01;
  wire v230d02b;
  wire v23fb699;
  wire v23fbf28;
  wire v2302fbf;
  wire v2391fb2;
  wire v23f3073;
  wire v22f9b75;
  wire v23fb70f;
  wire v22f3e5b;
  wire v23fbcf0;
  wire v23fc588;
  wire v23fbcde;
  wire v230d3c2;
  wire v22ff2c4;
  wire v23101dc;
  wire v2309573;
  wire v23fb845;
  wire v2310ada;
  wire v2309dce;
  wire v230786e;
  wire v23fbf00;
  wire v23f0489;
  wire v23f7ed6;
  wire v23f47ae;
  wire v230d45f;
  wire v230de87;
  wire v23fb0d0;
  wire v22f7d04;
  wire v22ebbde;
  wire v23135f8;
  wire v22ec502;
  wire v22f341f;
  wire v22fd032;
  wire v2301b99;
  wire v23f3ed0;
  wire v23f6d75;
  wire v22f1154;
  wire v230e50f;
  wire v230b49b;
  wire v22ff257;
  wire v2302c88;
  wire v22fd549;
  wire v230941d;
  wire v23fcb55;
  wire v23f7b1d;
  wire v2392d14;
  wire v23fcba3;
  wire v2300ab9;
  wire v23fc879;
  wire v23f6d6c;
  wire v2310754;
  wire c0aa95;
  wire v22f12fb;
  wire v23f1a14;
  wire v23fbf59;
  wire v230c579;
  wire v23fc164;
  wire v23f5a02;
  wire v23094f0;
  wire v23f1a4c;
  wire v230b086;
  wire v22f25a1;
  wire v22ff650;
  wire v23fc438;
  wire v22fd72d;
  wire v23061d7;
  wire v2313255;
  wire v23f47e3;
  wire v22fbde3;
  wire v22f4864;
  wire v22fafa3;
  wire v191abc5;
  wire v23113b5;
  wire v22f9056;
  wire v23f6fe8;
  wire v23107fc;
  wire v23fbea2;
  wire v23021ec;
  wire v23fca67;
  wire v22fb49a;
  wire v23fcc4e;
  wire v22fbd15;
  wire v2308f85;
  wire v23fc0fd;
  wire v230841a;
  wire v22f8278;
  wire a1ff27;
  wire v230d04a;
  wire v23efa52;
  wire v23011cb;
  wire v230f8b2;
  wire v22f3396;
  wire v23f280c;
  wire v22efc50;
  wire v23fc096;
  wire v23fc5a3;
  wire v23026ed;
  wire v230cfed;
  wire v230d8f3;
  wire v22f0fe5;
  wire v23130c9;
  wire v23001d0;
  wire v23fc005;
  wire v23f29e9;
  wire v23f3715;
  wire v13afebe;
  wire v22eecf9;
  wire v22f5974;
  wire v22ec562;
  wire v150715d;
  wire v230971e;
  wire b194d1;
  wire v230810c;
  wire v23f3321;
  wire v2309294;
  wire v22f3411;
  wire v23f5aa7;
  wire v23fccb3;
  wire v230b0f9;
  wire v23fcdb8;
  wire v23933b0;
  wire v2300687;
  wire v191ab12;
  wire v2392f80;
  wire v23018b7;
  wire v23fbb3e;
  wire v2307946;
  wire v2303125;
  wire v191ab91;
  wire v22fe51f;
  wire v2312912;
  wire v23f8f25;
  wire v22ed6ee;
  wire v22f1a1b;
  wire v23f8c71;
  wire v23f92d5;
  wire v23929a6;
  wire v23fbdac;
  wire v22f8aec;
  wire v230ed85;
  wire v23fbd5f;
  wire v23fc949;
  wire v230fa13;
  wire v23fcc7a;
  wire b7029b;
  wire v2391eaa;
  wire v23919f9;
  wire v230216e;
  wire v23fc956;
  wire v22f49ff;
  wire v22f78ef;
  wire v23fb59e;
  wire v22f4d46;
  wire v22f383e;
  wire v231007d;
  wire v22f7ef4;
  wire v22f6b4c;
  wire v22f6529;
  wire v230cd34;
  wire v22f737d;
  wire v22f263c;
  wire v22efe6e;
  wire f40cfd;
  wire v94116b;
  wire v22f877e;
  wire v23fc24a;
  wire v2301482;
  wire v2304c4c;
  wire v230b375;
  wire v2311ed4;
  wire v230f331;
  wire v22fc5e2;
  wire v97ba8e;
  wire v22f3ac3;
  wire v231049c;
  wire v22f6edc;
  wire v22ee43f;
  wire v23f9ba6;
  wire b9c90c;
  wire v23f1bd6;
  wire v230e94c;
  wire v22faf49;
  wire v22fe939;
  wire v22f161f;
  wire v2304253;
  wire v22eb993;
  wire v2303220;
  wire v23063fa;
  wire v23fb825;
  wire v230031f;
  wire v23f96aa;
  wire v22fa48c;
  wire v22fb1bc;
  wire v23fc53b;
  wire v22f4c34;
  wire v23f732a;
  wire v23f2278;
  wire v22f6bd4;
  wire v22f587e;
  wire v23105cd;
  wire v22eb332;
  wire v230de18;
  wire v23fbdec;
  wire v22ece0e;
  wire v23f71c9;
  wire v22f97e9;
  wire v230e1fc;
  wire v22f36ff;
  wire v23fb4e1;
  wire v2300934;
  wire v23fbedb;
  wire v23fc687;
  wire v22fe723;
  wire v230a4b6;
  wire v2308967;
  wire v23fcc5a;
  wire v22fef02;
  wire v23fc1bb;
  wire v23fcd14;
  wire v22f8838;
  wire v22f4bc7;
  wire v2303ae8;
  wire v23fc3cd;
  wire v23fbe4b;
  wire v23fbb25;
  wire v2311d38;
  wire v23fb553;
  wire v2311a61;
  wire v23019e9;
  wire v22efd33;
  wire v23fbb94;
  wire v22f009f;
  wire v23f5a39;
  wire v22f20df;
  wire v2392066;
  wire v230385f;
  wire v23fc754;
  wire v22f2ed7;
  wire v22fbeb1;
  wire v23fbe4f;
  wire v22f36a0;
  wire v23fce0b;
  wire v2301b00;
  wire v22f0069;
  wire v22f4858;
  wire v12cd51b;
  wire v230d90f;
  wire v22fe22a;
  wire v22f2158;
  wire v23fc9b2;
  wire v2302d12;
  wire v23fbf9b;
  wire v22f1172;
  wire v2308aec;
  wire v2305a09;
  wire v2312eaa;
  wire v23fc281;
  wire v22f4bcc;
  wire v23fc04e;
  wire v23fc142;
  wire v23068cd;
  wire v23fa460;
  wire v23fcc8f;
  wire v230edc0;
  wire v23fb1c3;
  wire v22f7793;
  wire a507a6;
  wire v22efbaa;
  wire v22ec531;
  wire v23f5686;
  wire v230eef7;
  wire v23fc4f8;
  wire v22f5405;
  wire v2303bee;
  wire v230bed2;
  wire v23fcbcd;
  wire v23f535c;
  wire v230d91f;
  wire v22f0677;
  wire v2312259;
  wire v23f8a70;
  wire v22ff29c;
  wire v2307b42;
  wire v230d56c;
  wire v2308818;
  wire v22f2e69;
  wire v2312cf2;
  wire v22f4163;
  wire v2310ec8;
  wire v23f52b9;
  wire v23fc60b;
  wire v22fc399;
  wire v23fb66e;
  wire v2301c10;
  wire v23916d8;
  wire v23fba9c;
  wire v23fa6f1;
  wire v23f9414;
  wire v2309c99;
  wire v23fc361;
  wire v2309cdc;
  wire v2311d52;
  wire v22f2abb;
  wire v23fc252;
  wire v23f7ab7;
  wire v230fc1f;
  wire v2302875;
  wire v22ffc07;
  wire v23f5f5f;
  wire v230a709;
  wire v23f67fa;
  wire v22fcab7;
  wire v23fc1f0;
  wire v23fcfbb;
  wire v22ede34;
  wire v22feb98;
  wire v23f3997;
  wire v23fc95a;
  wire v23fc1aa;
  wire v22fe392;
  wire v23fb787;
  wire v23f594f;
  wire v22f8291;
  wire v2303253;
  wire v230f6e9;
  wire v2312248;
  wire v22f979e;
  wire v23076ca;
  wire v23f6077;
  wire v22edb22;
  wire v23fb67c;
  wire v22f092f;
  wire v22eb659;
  wire v23035ba;
  wire v22f62ea;
  wire v230b7fc;
  wire v23fca4f;
  wire v23fbeb0;
  wire v23099fc;
  wire v23054d5;
  wire v2307707;
  wire v230f34c;
  wire v2303115;
  wire v23f173d;
  wire v238aeb0;
  wire v22f4aa2;
  wire v22efb77;
  wire v22f82cd;
  wire v2301a5f;
  wire v8ea3a5;
  wire v23fbeaf;
  wire v23f1686;
  wire v22f9188;
  wire v22fca1d;
  wire v2346b90;
  wire v23fc31c;
  wire v2308ac3;
  wire v23f4edf;
  wire b00ac7;
  wire v23fca43;
  wire v230466c;
  wire v22f0104;
  wire v23fb1d6;
  wire v22fb9ad;
  wire v2301c2e;
  wire v23f9e84;
  wire v23fcdef;
  wire v23fc3c7;
  wire v22eb51e;
  wire v230930b;
  wire v23034e5;
  wire v23f6591;
  wire v23fcf5d;
  wire v2305fbf;
  wire v231359f;
  wire v22ebb15;
  wire ae0418;
  wire v2300ba2;
  wire v2309efb;
  wire v2392697;
  wire v230b4d4;
  wire v22f03a2;
  wire v2308fe5;
  wire v231171e;
  wire v239268e;
  wire v231160c;
  wire v22fa99c;
  wire v2392f52;
  wire v23116b7;
  wire v230444c;
  wire v22fa1ab;
  wire v23f0dd4;
  wire v22ff67c;
  wire v22f25e0;
  wire v2310317;
  wire v2303efe;
  wire v22ef61b;
  wire v23f1803;
  wire v231094e;
  wire v1aae9f4;
  wire a2cc4e;
  wire v22f8c55;
  wire v23fbff1;
  wire v23fa4bb;
  wire v23f2bbf;
  wire v22fbd88;
  wire v23fcf1f;
  wire v23fcc1f;
  wire v23023c9;
  wire c258f4;
  wire v23fc660;
  wire v23fbfe4;
  wire v23057e6;
  wire v2313247;
  wire v22febaf;
  wire v2306e5a;
  wire v23fc54f;
  wire v2302a8c;
  wire v230b611;
  wire v23fbacf;
  wire v23fb1c1;
  wire b67ed5;
  wire v22ef751;
  wire v23fcd1b;
  wire v22fa707;
  wire v22f0051;
  wire v2311d12;
  wire v22ec299;
  wire v22f7808;
  wire v22eb895;
  wire v23fca07;
  wire v22eee6a;
  wire v22ec191;
  wire v23017f0;
  wire v23fcdd5;
  wire v22ef683;
  wire v230ee7d;
  wire v23fbdea;
  wire v23f71d5;
  wire v23fd064;
  wire v22f7b13;
  wire v22f2a60;
  wire v23fc6c0;
  wire v23fb4d7;
  wire v22fb0c7;
  wire v22fc8d0;
  wire v22f9ddc;
  wire v23f6215;
  wire v23017c7;
  wire v23f5f94;
  wire v8da3ef;
  wire v2306873;
  wire v231363b;
  wire v22fd9be;
  wire v23114a6;
  wire v2312bd0;
  wire v23f9a93;
  wire v2306fa2;
  wire v23fc01c;
  wire v1e84012;
  wire v23fb9ea;
  wire v23f4e99;
  wire v23f134a;
  wire v2309729;
  wire v230be96;
  wire v2311b20;
  wire v2393b99;
  wire v23065e7;
  wire v23fd00f;
  wire v23fcaea;
  wire v23f9ef5;
  wire v191b1b9;
  wire v230df44;
  wire v22fc22b;
  wire v22f24a3;
  wire v23042ca;
  wire v23fb0eb;
  wire v2312e02;
  wire v23fb584;
  wire v23006de;
  wire v2307742;
  wire v2300ac2;
  wire f40c96;
  wire v22f3b08;
  wire v2303376;
  wire v22f931f;
  wire v2303b76;
  wire v230af3a;
  wire v230b02b;
  wire v23fcca4;
  wire v23f0652;
  wire v23fa3a4;
  wire v22f6e70;
  wire v8f4f78;
  wire v2305833;
  wire v22f5815;
  wire v22feb6b;
  wire v23f9864;
  wire v22eeb27;
  wire v22f3840;
  wire v230f94d;
  wire v23022ab;
  wire v8bbb53;
  wire v230591e;
  wire v23005a9;
  wire v230bece;
  wire v22ff63a;
  wire v23fbc74;
  wire v2391735;
  wire v1aae0dc;
  wire v23fbce3;
  wire v23fc0a6;
  wire v23fbfcf;
  wire v22f0323;
  wire v22fd699;
  wire v22eec6e;
  wire v230e85f;
  wire v230beb8;
  wire v2392ff0;
  wire v23fd014;
  wire v22f915d;
  wire v230a44c;
  wire f40a9e;
  wire v23fbed5;
  wire v22f2ffe;
  wire v23fc21c;
  wire v2313367;
  wire v2307d08;
  wire be7d90;
  wire v23101f4;
  wire v2305684;
  wire v230b750;
  wire v23fb952;
  wire v230ce60;
  wire v230f9c2;
  wire v23f6769;
  wire v22ed8bc;
  wire v22fdbd2;
  wire v23fbcd4;
  wire v23f1e4f;
  wire v23f4e1c;
  wire v230988d;
  wire v23fbd75;
  wire v23fbc7f;
  wire v2393f95;
  wire v22ffd9a;
  wire v23f1703;
  wire v23fc30b;
  wire v22fd2f5;
  wire v2306e1a;
  wire v2305ebc;
  wire v22f1796;
  wire v23f6089;
  wire v230e41f;
  wire v23fa23d;
  wire v22f6ed4;
  wire v23fb727;
  wire v23f50f8;
  wire v2302c0e;
  wire v23fb960;
  wire v2311891;
  wire v22f6372;
  wire v23f5caf;
  wire v23f988f;
  wire v23f7031;
  wire v23fc26f;
  wire v23fc765;
  wire v12cc2f8;
  wire v23915d8;
  wire v22f4e77;
  wire v23087b6;
  wire v23f6c84;
  wire v23fc881;
  wire v2393c38;
  wire v23030ae;
  wire v1b87752;
  wire v230c589;
  wire v22f8b0a;
  wire v22f6ac8;
  wire v22ee8f3;
  wire v22f3b24;
  wire v23084fa;
  wire v2301de9;
  wire v23fbe82;
  wire v22f4f19;
  wire c60af7;
  wire v23f8e25;
  wire v22ec339;
  wire v23074cd;
  wire v2393dd2;
  wire v2305194;
  wire b5b985;
  wire v2304477;
  wire v23fc528;
  wire v22f1ef1;
  wire v22ff129;
  wire v23fcb5a;
  wire v23faab2;
  wire v230fe15;
  wire v22fa11e;
  wire v23f65cd;
  wire v23f6954;
  wire v23049af;
  wire v230437d;
  wire v22f9ebc;
  wire v230f883;
  wire v230db5e;
  wire v22ef0ab;
  wire v230062b;
  wire v23f9d8e;
  wire v22fc351;
  wire v23f3ff7;
  wire v22f3cc0;
  wire v22ebfcb;
  wire v23fc5fe;
  wire v23fbe0d;
  wire v23003fc;
  wire v23f7de2;
  wire b79082;
  wire v22f8f8c;
  wire v23fc223;
  wire v230da9b;
  wire v23f78a3;
  wire v22f7a20;
  wire v23fbce1;
  wire v22f3550;
  wire v23fca2f;
  wire v23fc999;
  wire v23fbea7;
  wire v230cb63;
  wire v23fccc2;
  wire v23fccd7;
  wire v2301565;
  wire v23f7503;
  wire v2310385;
  wire v23f87e1;
  wire v22fbd4f;
  wire v22eee95;
  wire v2307c63;
  wire v23fc598;
  wire v23fbcd8;
  wire v2310d79;
  wire v22f2e48;
  wire v22f89b9;
  wire v23f0dd1;
  wire v22fd55f;
  wire v22f04bf;
  wire v22f9734;
  wire v22ec2ba;
  wire v23028fc;
  wire da30fb;
  wire f405c6;
  wire v22f9497;
  wire v23fc5ba;
  wire v2301b2d;
  wire v22f7004;
  wire v230f860;
  wire v22f22b2;
  wire v22fb5bd;
  wire v22f7da7;
  wire v22efd4d;
  wire v22f7195;
  wire v23f7254;
  wire v230ec39;
  wire v22ed684;
  wire v23fbd2f;
  wire v2312637;
  wire v22f2879;
  wire v2312336;
  wire v23fb6c2;
  wire v230173a;
  wire v230522c;
  wire v22f2b78;
  wire v23fc404;
  wire v86c778;
  wire v12cc30c;
  wire v23fc6db;
  wire v230b879;
  wire v22f3839;
  wire v23fcf81;
  wire v23f67d3;
  wire v191a912;
  wire v2308a91;
  wire v23fc908;
  wire v23f333e;
  wire v2309c1f;
  wire v230dde6;
  wire v2304928;
  wire v23073e4;
  wire v23fcd88;
  wire v23fbffc;
  wire v23fab2c;
  wire v23fc5c4;
  wire v2302520;
  wire v23fb691;
  wire v23fb5c4;
  wire v2308813;
  wire v22f958d;
  wire v23093a7;
  wire v2303f89;
  wire v2392095;
  wire v2313564;
  wire f4066f;
  wire v23fc57e;
  wire c16191;
  wire v23f6926;
  wire v22fb00d;
  wire v22fd794;
  wire v23fc8c3;
  wire v23fc36e;
  wire a0d50a;
  wire v22f5836;
  wire v230cef0;
  wire v23fc741;
  wire e1e726;
  wire v22fd002;
  wire v9f5c3c;
  wire v22f13d8;
  wire v22f3d18;
  wire v230a3e2;
  wire v22efc28;
  wire v23fbb8f;
  wire v23fc505;
  wire v23f8368;
  wire v2311c65;
  wire v2301972;
  wire v23fc5ea;
  wire v22f26d2;
  wire v23fbe79;
  wire v8c495d;
  wire v23fc7e8;
  wire v23fa590;
  wire v23fc6cc;
  wire v23fcb1b;
  wire v23f5c60;
  wire v23fb569;
  wire v22fa8e8;
  wire v23f23bf;
  wire v22ffed0;
  wire v230ada5;
  wire v230d2d8;
  wire v22f8f34;
  wire v23fc673;
  wire v22eb748;
  wire v22f7ad4;
  wire v23f0978;
  wire v23fb95a;
  wire v23fcc9e;
  wire v230f31f;
  wire a28a9e;
  wire v1aaddfe;
  wire v22ef3fe;
  wire v23fbf5d;
  wire v230c322;
  wire v23fc297;
  wire v23fbe69;
  wire v23f420d;
  wire v23fb92f;
  wire v22feac9;
  wire v23100e9;
  wire v230d5ca;
  wire v23fc8b8;
  wire v230cc70;
  wire v23fcb01;
  wire v23fc095;
  wire v23f8a29;
  wire v22faf3a;
  wire v2393332;
  wire v23fcd39;
  wire v22f1cb7;
  wire v23fb99b;
  wire v22fcf5b;
  wire v23fc742;
  wire v22eefcf;
  wire v23f36c8;
  wire v22ef2aa;
  wire v2310826;
  wire v23fc4b1;
  wire v23f4f1e;
  wire v23f4fbf;
  wire v23fbef9;
  wire v23f66a8;
  wire v23f4da0;
  wire v23fc988;
  wire v2311bc4;
  wire v23f179d;
  wire v22ed400;
  wire v23fbf63;
  wire v23f19e4;
  wire v23031c2;
  wire v23f4827;
  wire v23ef951;
  wire v230b304;
  wire v22ef663;
  wire v230891d;
  wire v230f96f;
  wire v23f9492;
  wire v23fba43;
  wire v22f8d6a;
  wire v23fbcbb;
  wire v230d3f5;
  wire v23fc66d;
  wire v230e01b;
  wire v23f412d;
  wire v23fcf4d;
  wire v23fc44e;
  wire v230e1e4;
  wire v23f64db;
  wire v23f7423;
  wire v2305b70;
  wire v230875f;
  wire v22f959d;
  wire v23130d9;
  wire v22eea52;
  wire v22f16d5;
  wire v23fc215;
  wire v22ffb10;
  wire v23fc2b1;
  wire v23fb923;
  wire v22fd6a4;
  wire v230104e;
  wire v230b0f5;
  wire v22fe326;
  wire v23fc68a;
  wire v2304b05;
  wire v23fbf27;
  wire v1507557;
  wire v22fb5f1;
  wire v22fa05b;
  wire v22f8e1b;
  wire v23fbe1d;
  wire da38c9;
  wire v22f7cbf;
  wire v230c616;
  wire v22f7a60;
  wire v23065ee;
  wire v23fce12;
  wire v2307949;
  wire v22f2759;
  wire v13afbf5;
  wire v23fbc8c;
  wire v230e6ee;
  wire v2309cfe;
  wire v23fb0ea;
  wire v23f7114;
  wire v22f92f9;
  wire v22fc3ed;
  wire v231086f;
  wire v23fb56e;
  wire v22eed5b;
  wire v22ef542;
  wire v23083e6;
  wire v23f17e2;
  wire v23fc6c4;
  wire v23efcf8;
  wire v23f5ede;
  wire v230557c;
  wire v22fefa1;
  wire v22eb134;
  wire v22f8e56;
  wire v239310f;
  wire v22f9e5b;
  wire v22fe0ee;
  wire v2312f3c;
  wire v23faf8a;
  wire v23f4cd4;
  wire v22fbc63;
  wire v23f6c41;
  wire v23f8ca4;
  wire v23fc8d4;
  wire v2311743;
  wire v22f3add;
  wire v22ec1ef;
  wire v22f8ebe;
  wire v23fc3af;
  wire v230e352;
  wire v22f0e6b;
  wire v22faa7c;
  wire v2300774;
  wire v23fce05;
  wire v23fb31d;
  wire v23f2650;
  wire v2307b64;
  wire v22f8013;
  wire v2306bd7;
  wire v23f6623;
  wire v22ec1ae;
  wire v22fa934;
  wire v230727f;
  wire afc788;
  wire v23fcabb;
  wire v230fb99;
  wire v2303d8f;
  wire v23fb4d4;
  wire v22f76f0;
  wire v22fbfaf;
  wire v230bdbb;
  wire v2311ed7;
  wire v2304672;
  wire a3cb61;
  wire v230cd57;
  wire v22f1339;
  wire v22f8240;
  wire v22f92ec;
  wire v23fc8a0;
  wire v23f5140;
  wire v231192e;
  wire v13afaae;
  wire v22f9b5b;
  wire v23f9b8d;
  wire v191abee;
  wire bd7b37;
  wire v22fa16d;
  wire v23fcfcc;
  wire v23f0386;
  wire v23062f8;
  wire v22f9f27;
  wire v23fc716;
  wire bfb87c;
  wire v22ed5fd;
  wire v23fbe3a;
  wire v23f1263;
  wire v23f4ae1;
  wire v22f6735;
  wire v22f9838;
  wire v2305de3;
  wire v22f8dea;
  wire v23fc7d7;
  wire v230e897;
  wire v23fcf69;
  wire v23f5207;
  wire v2305507;
  wire v23112a4;
  wire v23fbafc;
  wire v230c4ea;
  wire acdb9d;
  wire v22ff50f;
  wire v22ebeb2;
  wire v22fd1ba;
  wire v1aad69f;
  wire v22f1b63;
  wire v22fcd0c;
  wire v22f96f2;
  wire v2391a43;
  wire v23041a1;
  wire v230065d;
  wire v23fca72;
  wire v23f9631;
  wire v22fcc05;
  wire v22ecc3b;
  wire v2301073;
  wire v22f9ab1;
  wire v23fbf41;
  wire v23fbd70;
  wire v22ec890;
  wire v23fb90f;
  wire v22eca65;
  wire v22fad0f;
  wire v23fc3e7;
  wire v23fc9e8;
  wire v2301abc;
  wire v23fca32;
  wire v2306609;
  wire v23040f3;
  wire v23035a3;
  wire v230a989;
  wire v23f08d9;
  wire v230fdb8;
  wire v22fc979;
  wire v2309033;
  wire v23f4267;
  wire v2309b3e;
  wire v12cd920;
  wire v23fc44c;
  wire f40d2d;
  wire v23fc2c6;
  wire v23fcf87;
  wire v230fae1;
  wire v230c995;
  wire v23fcf0e;
  wire v2303a32;
  wire v2311b78;
  wire v191afef;
  wire v2307517;
  wire v230bbda;
  wire v22edd3d;
  wire v23f6a5b;
  wire v22f836e;
  wire v22fa61c;
  wire v22f1a0e;
  wire v2310291;
  wire v23fb8bd;
  wire v23052a2;
  wire v23fc6dd;
  wire v22ef530;
  wire v2300f19;
  wire v2304258;
  wire v2391935;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hbusreq2_p;
  input hbusreq2;
  reg hlock2_p;
  input hlock2;
  reg hbusreq3_p;
  input hbusreq3;
  reg hlock3_p;
  input hlock3;
  reg hbusreq4_p;
  input hbusreq4;
  reg hlock4_p;
  input hlock4;
  reg hbusreq5_p;
  input hbusreq5;
  reg hlock5_p;
  input hlock5;
  reg hbusreq6_p;
  input hbusreq6;
  reg hlock6_p;
  input hlock6;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmaster1_p;
  output hmaster1;
  reg hmaster2_p;
  output hmaster2;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg hgrant2_p;
  output hgrant2;
  reg hgrant3_p;
  output hgrant3;
  reg hgrant4_p;
  output hgrant4;
  reg hgrant5_p;
  output hgrant5;
  reg hgrant6_p;
  output hgrant6;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg stateG10_2_p;
  output stateG10_2;
  reg stateG10_3_p;
  output stateG10_3;
  reg stateG10_4_p;
  output stateG10_4;
  reg stateG10_5_p;
  output stateG10_5;
  reg stateG10_6_p;
  output stateG10_6;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;
  reg jx2_p;
  output jx2;
  reg jx3_p;
  output jx3;

assign v22fc399 = hmaster0_p & v22f2e69 | !hmaster0_p & v23fc60b;
assign v2305aa7 = hbusreq3_p & v23efbfd | !hbusreq3_p & v23fc01d;
assign v22ecbc1 = hbusreq3_p & v12cdab5 | !hbusreq3_p & v22f18b5;
assign v23fc9be = hmaster2_p & v22f9980 | !hmaster2_p & !v2392d6d;
assign v22ebfd3 = hmaster0_p & v22feec8 | !hmaster0_p & v23f6635;
assign v84571e = hbusreq3 & v23fcfd0 | !hbusreq3 & v84561b;
assign v23fc9de = hgrant1_p & v23fb6ff | !hgrant1_p & v22f331e;
assign v22eea6a = hbusreq4_p & v23fc5e5 | !hbusreq4_p & v23f3e77;
assign v23fbe12 = hbusreq5 & fc8ab7 | !hbusreq5 & !v84561b;
assign v921155 = hmaster1_p & v84561b | !hmaster1_p & v230899e;
assign v23fbb8d = hbusreq1_p & v22ee44f | !hbusreq1_p & !v23f2cbe;
assign v23fca38 = hgrant3_p & v23fca50 | !hgrant3_p & v22eef44;
assign v2308d09 = hlock1_p & v191aa68 | !hlock1_p & v191a86f;
assign v2308d63 = hmaster2_p & v106a782 | !hmaster2_p & !v23f908f;
assign v23f28de = hmaster0_p & v23fbfbb | !hmaster0_p & v2308627;
assign f40cfd = hmaster0_p & v22f49ff | !hmaster0_p & v22efe6e;
assign v1aadf17 = hmaster2_p & v22fd655 | !hmaster2_p & v84561b;
assign v23058ba = hbusreq2_p & da38c1 | !hbusreq2_p & v84561b;
assign v22f7fcc = hbusreq4 & v22f24ca | !hbusreq4 & b0fad6;
assign v23fbe24 = hbusreq3_p & b09503 | !hbusreq3_p & v23f9395;
assign v2307a72 = hbusreq4_p & v23fc994 | !hbusreq4_p & v84561b;
assign v23f7ffb = hmastlock_p & v239298c | !hmastlock_p & v84561b;
assign v22fd9f5 = hbusreq3_p & v23059ee | !hbusreq3_p & v84561b;
assign v22f483c = hmaster2_p & v15072a9 | !hmaster2_p & v22f04d8;
assign v23fc73e = hbusreq0_p & v23fc513 | !hbusreq0_p & v845629;
assign v23fc1de = hgrant2_p & v84562a | !hgrant2_p & v22eedf9;
assign v191a8f7 = hmaster0_p & v22f4d17 | !hmaster0_p & e1dea8;
assign v23088a9 = hbusreq4_p & v230193c | !hbusreq4_p & v2311668;
assign v230f578 = hmaster2_p & v2312f7e | !hmaster2_p & v23027e9;
assign v230f2af = hmaster2_p & v22f8271 | !hmaster2_p & b5f51c;
assign v22f9880 = hbusreq1_p & v22f5037 | !hbusreq1_p & v22fbbb8;
assign v2393f05 = hgrant3_p & v191acbd | !hgrant3_p & v22fe44f;
assign v23f1d35 = hbusreq0 & v23f8da8 | !hbusreq0 & v84561b;
assign v23fc215 = hbusreq1_p & v22f16d5 | !hbusreq1_p & v84561b;
assign v22fc8d0 = hbusreq3 & v23fb4d7 | !hbusreq3 & v22fb0c7;
assign v23fca61 = hlock0_p & v23fbba4 | !hlock0_p & v22f2aa4;
assign v22ed287 = hgrant6_p & v845631 | !hgrant6_p & e1e78b;
assign v230d2c7 = hgrant5_p & v22fa88a | !hgrant5_p & v23fc338;
assign v2304b4d = hbusreq2 & v23022b1 | !hbusreq2 & !v84561b;
assign v23fb2d6 = hbusreq3 & v23fc49b | !hbusreq3 & v84564d;
assign v23fce0b = hbusreq3_p & v22f36a0 | !hbusreq3_p & v84561b;
assign v22f5b18 = hmaster2_p & v22ee0c4 | !hmaster2_p & !v84561b;
assign v22f825a = hbusreq0 & v2301505 | !hbusreq0 & v84561b;
assign v23f1cd2 = hbusreq5_p & v22fdabc | !hbusreq5_p & v84561b;
assign v22f60da = hmaster2_p & v23fa4ca | !hmaster2_p & v23fc896;
assign v22f39a1 = stateA1_p & v84561b | !stateA1_p & v23f7992;
assign v22f91c9 = hmastlock_p & v106a7d6 | !hmastlock_p & v84561b;
assign v23fb937 = hmaster2_p & v23f4b28 | !hmaster2_p & v84561b;
assign v845632 = hbusreq4 & v84561b | !hbusreq4 & !v84561b;
assign v23f12d0 = hbusreq6_p & v230edb2 | !hbusreq6_p & v22fbb0f;
assign v2306b99 = hbusreq6_p & v22f947f | !hbusreq6_p & v23133be;
assign v22eea5b = hbusreq3 & v2313351 | !hbusreq3 & v230f7ff;
assign v23f19ee = hmaster2_p & v22f337b | !hmaster2_p & v2310e10;
assign b08eee = hbusreq4 & v2303fe4 | !hbusreq4 & v84561b;
assign v23fc098 = hbusreq3_p & v230426b | !hbusreq3_p & v22eaea8;
assign v12cd586 = hbusreq4_p & v23f98a9 | !hbusreq4_p & v23fb63e;
assign v23fccfe = hlock2_p & v22fca61 | !hlock2_p & v23f6b25;
assign v22f5d0e = hgrant1_p & v12cd9f9 | !hgrant1_p & !v23fa1ad;
assign v23fbf02 = hmaster0_p & v2313266 | !hmaster0_p & v22f1b18;
assign v23087b6 = hbusreq1_p & v23915d8 | !hbusreq1_p & v22f4e77;
assign v230d1c3 = hbusreq3 & v1e84028 | !hbusreq3 & v845645;
assign v23fbcbb = hbusreq1_p & v22f8d6a | !hbusreq1_p & v84561b;
assign v22fc3d9 = hmaster0_p & v231347a | !hmaster0_p & !v23fb081;
assign v23fc787 = hmaster0_p & v23fc34f | !hmaster0_p & v23fbe15;
assign v23fb7e0 = hgrant5_p & v1aad63a | !hgrant5_p & v22fe097;
assign v23045ac = hgrant0_p & v2309b0f | !hgrant0_p & v23f3a8b;
assign v23fc5a8 = hbusreq0 & v22fc4d8 | !hbusreq0 & !v22eedf9;
assign v23f36c8 = hmaster2_p & v23fc742 | !hmaster2_p & v2310754;
assign v22f7885 = hbusreq5 & v230882d | !hbusreq5 & !v84561b;
assign v22f753d = hlock0_p & v22fd30c | !hlock0_p & v2308592;
assign v23fc393 = busreq_p & v230eb13 | !busreq_p & !v23fcb38;
assign v230426b = hmaster2_p & v230ff7d | !hmaster2_p & v22f8c43;
assign v2301fc9 = hbusreq5_p & v2311290 | !hbusreq5_p & !v84561b;
assign v22f9e59 = hbusreq3_p & v23fcc58 | !hbusreq3_p & v84561b;
assign v22f2998 = hgrant1_p & v22f3ed0 | !hgrant1_p & v23f8c7b;
assign v22fd49d = hbusreq6_p & v230e97b | !hbusreq6_p & v230a0e7;
assign v22f7ad5 = hbusreq3 & v22f975b | !hbusreq3 & v84561b;
assign v2310754 = hgrant1_p & v84561b | !hgrant1_p & v23f6d6c;
assign v22fce0a = hgrant3_p & v2309d09 | !hgrant3_p & v22fcb45;
assign v22f9ddc = hmaster2_p & v23fc6c0 | !hmaster2_p & v23fb1c1;
assign v23f81cf = hgrant0_p & v84561b | !hgrant0_p & v22fe992;
assign v23fcd35 = hbusreq4_p & v2301c48 | !hbusreq4_p & v84561b;
assign v2308a1b = hmaster0_p & v22eed68 | !hmaster0_p & v23efcfb;
assign v230ce98 = hmaster2_p & v22fab30 | !hmaster2_p & v22f3c6b;
assign v23fb323 = hmaster0_p & v2304987 | !hmaster0_p & v22f9a50;
assign v23fc6fe = hbusreq2_p & f40d2a | !hbusreq2_p & v84561b;
assign v2304deb = hgrant1_p & v22ffbb3 | !hgrant1_p & v23f89fe;
assign v106ae74 = hgrant5_p & v23fcd71 | !hgrant5_p & v23fcb53;
assign v22f9b42 = hbusreq2 & v2393bce | !hbusreq2 & v84561b;
assign v22f47b0 = hbusreq2 & v23fbb11 | !hbusreq2 & v84561b;
assign v23fc300 = jx0_p & v22f779a | !jx0_p & v230e568;
assign v22ed491 = hbusreq6 & v22f46d3 | !hbusreq6 & v84561b;
assign a1bfd6 = hgrant0_p & v84561b | !hgrant0_p & !v845653;
assign v23fbc46 = hbusreq6_p & v22f6f2d | !hbusreq6_p & !v84561b;
assign v23fbab3 = stateG2_p & v84561b | !stateG2_p & !v230f0a1;
assign v15071a5 = hgrant0_p & v22f1f6f | !hgrant0_p & v23f51b1;
assign v2391b6f = hgrant1_p & v23fca0c | !hgrant1_p & v150748b;
assign v23f8b6b = hgrant0_p & v84561b | !hgrant0_p & v2307b18;
assign v23125a2 = hmaster0_p & v239174f | !hmaster0_p & v23f3d14;
assign abc0f5 = hbusreq4 & v23f15c1 | !hbusreq4 & v845627;
assign v22fe71e = hbusreq1_p & v1aae56f | !hbusreq1_p & v13affaa;
assign v230a22e = hbusreq5_p & da38c1 | !hbusreq5_p & v230ac9e;
assign v230aef9 = hbusreq5 & v22f2718 | !hbusreq5 & v84561b;
assign v22f66bc = hlock0_p & v106af73 | !hlock0_p & v191a879;
assign v23fc355 = hlock1_p & bc2a58 | !hlock1_p & v2305748;
assign v23135cf = jx2_p & v2303481 | !jx2_p & v84561b;
assign v2308592 = hbusreq0_p & v22fd30c | !hbusreq0_p & v22f6a6b;
assign v22f5110 = hbusreq5_p & v230f1ae | !hbusreq5_p & !v84561b;
assign v23fbffe = hbusreq0 & v13affaa | !hbusreq0 & v84561b;
assign b50a75 = hbusreq1_p & v845627 | !hbusreq1_p & !v84561b;
assign v23071f6 = hgrant5_p & v23055b3 | !hgrant5_p & v23f4af5;
assign v23050fb = hbusreq6_p & fc90a8 | !hbusreq6_p & v2313111;
assign v2307742 = hbusreq1_p & v23fb584 | !hbusreq1_p & v23006de;
assign v23008f3 = hbusreq3_p & v230a934 | !hbusreq3_p & v23fcd24;
assign v23075bd = hmaster1_p & v23fb843 | !hmaster1_p & v23f66fd;
assign v23fca2d = hbusreq0_p & v22ecc15 | !hbusreq0_p & v2392d6d;
assign v230c83a = hmaster2_p & v22f9980 | !hmaster2_p & !v22f35e8;
assign v23fb8cb = hbusreq3_p & v22fea3e | !hbusreq3_p & v23fc256;
assign v22f25ac = hgrant4_p & v84561b | !hgrant4_p & v230c6c7;
assign v23f029a = hmaster1_p & v23f649a | !hmaster1_p & v23fb948;
assign v23f8490 = hbusreq5_p & v23129bb | !hbusreq5_p & !v84561b;
assign v2301400 = stateG10_5_p & v84561b | !stateG10_5_p & v2307e48;
assign v23f7cea = hbusreq4 & v23fba94 | !hbusreq4 & v23fba11;
assign v22ebe86 = hlock6_p & v23f3dd7 | !hlock6_p & v23fc834;
assign v23efd8a = hbusreq6_p & v23fbb58 | !hbusreq6_p & v2309305;
assign v2300de1 = hmaster2_p & v84561b | !hmaster2_p & v23fbb80;
assign v23fc67c = hbusreq3 & v23f8466 | !hbusreq3 & v230a91b;
assign v22fef20 = hbusreq1_p & v22fd00f | !hbusreq1_p & v84561b;
assign v2393705 = jx1_p & v22f1892 | !jx1_p & v23047dd;
assign v23084cc = hmaster0_p & v23fc357 | !hmaster0_p & v22fbebb;
assign v239379c = hbusreq0 & v23036ca | !hbusreq0 & v22eedf9;
assign v22f2abb = hbusreq3_p & v2309c99 | !hbusreq3_p & v2311d52;
assign v23f8299 = jx1_p & v22fbe9c | !jx1_p & v23fca3b;
assign v230679a = hlock0_p & v23f3a55 | !hlock0_p & v2311e62;
assign v230a8ea = hbusreq0 & v1aadb8e | !hbusreq0 & v84561b;
assign v22f69c6 = hgrant1_p & v84561b | !hgrant1_p & v230d82c;
assign v2300e92 = hmaster1_p & v23126b7 | !hmaster1_p & v23fb062;
assign v230b0f2 = hbusreq4_p & v22f8cb9 | !hbusreq4_p & v230ec04;
assign v23fbac0 = hmaster2_p & v22f61b6 | !hmaster2_p & v22ff90b;
assign v2393401 = hmaster0_p & v22fda61 | !hmaster0_p & v23efa84;
assign v22ede51 = hmaster0_p & v23f12d3 | !hmaster0_p & v22fe1c8;
assign v230ed6b = hbusreq3 & v12cd3e7 | !hbusreq3 & v84561b;
assign v22fb769 = hmaster2_p & v23f7370 | !hmaster2_p & v22f1244;
assign bd953c = hbusreq6_p & ae1a21 | !hbusreq6_p & a878fd;
assign v22f421a = hmaster0_p & v23fb9f0 | !hmaster0_p & v23f6fed;
assign v23f8d5a = hmaster0_p & v23132fc | !hmaster0_p & a7fdb1;
assign v230f4d3 = stateG3_0_p & v845665 | !stateG3_0_p & !v845665;
assign v23f62c2 = hlock4_p & v2305866 | !hlock4_p & v23fcfce;
assign v22f28eb = hbusreq6 & v23fc497 | !hbusreq6 & v84561b;
assign v23f7950 = hmaster0_p & v23fca38 | !hmaster0_p & v2393de1;
assign v2311761 = hmaster0_p & v23fbe30 | !hmaster0_p & v23041ab;
assign v23070dd = hmaster0_p & v23090fd | !hmaster0_p & v22f84a0;
assign v22f732c = hbusreq3_p & v23f408c | !hbusreq3_p & v84561b;
assign v23fca1d = hbusreq6 & v23f4f9f | !hbusreq6 & !v1aae385;
assign v23f5a2e = hbusreq5_p & v23fbbf2 | !hbusreq5_p & v22efcd6;
assign v230b77c = hlock6_p & v2306790 | !hlock6_p & !v84561b;
assign v2310731 = hmaster2_p & v22feae3 | !hmaster2_p & v2308786;
assign v23f5dca = hmaster2_p & v97b973 | !hmaster2_p & v22efae1;
assign v23f4f88 = hmaster0_p & v22f25ae | !hmaster0_p & !v22feb8b;
assign v2306775 = hburst1 & v230177d | !hburst1 & v2313264;
assign v230ed08 = hbusreq3 & v23fc180 | !hbusreq3 & !v1aad988;
assign v22f92f9 = hmastlock_p & v23f7114 | !hmastlock_p & v84561b;
assign v2303b86 = hmaster0_p & v23fb926 | !hmaster0_p & v23fca9d;
assign v23fc6e5 = hbusreq3 & v2307c0c | !hbusreq3 & v845636;
assign v23fb92f = hmaster0_p & v22f82cd | !hmaster0_p & v23f420d;
assign v23fccbc = hbusreq3 & v230c480 | !hbusreq3 & v22f1153;
assign v2310108 = hbusreq1_p & v2301eb1 | !hbusreq1_p & v84561b;
assign v22eaafd = hlock0_p & v23fbb35 | !hlock0_p & !v845622;
assign a75533 = hgrant3_p & a1fbc2 | !hgrant3_p & v22ee68f;
assign v2313965 = hbusreq1_p & v23fc561 | !hbusreq1_p & v23f10a4;
assign v2307a62 = hbusreq1 & v23131e8 | !hbusreq1 & v2306220;
assign v23fc7f9 = hmaster2_p & v84561b | !hmaster2_p & v2311918;
assign v22febaf = hmaster2_p & v2313247 | !hmaster2_p & v22f8b01;
assign v23fc1aa = hmaster0_p & v22ede34 | !hmaster0_p & v23fc95a;
assign b6f86d = hready & v84561b | !hready & !v23f2508;
assign v23fcf46 = locked_p & v84561b | !locked_p & !v23fba6b;
assign v22fe097 = hgrant0_p & v230d509 | !hgrant0_p & v23007a2;
assign v23fc005 = hbusreq6_p & v23001d0 | !hbusreq6_p & v84561b;
assign v23f5b31 = hmaster0_p & v230a9a3 | !hmaster0_p & v22fbdd6;
assign v23fb708 = hlock0_p & v22f654e | !hlock0_p & v84561b;
assign v22edf81 = hgrant1_p & v230b4af | !hgrant1_p & v23fca23;
assign v22ed684 = hgrant3_p & f405c6 | !hgrant3_p & v230ec39;
assign v13afe7d = stateG10_5_p & v23f08e5 | !stateG10_5_p & v2307725;
assign v2307d08 = hgrant3_p & v23fc0a6 | !hgrant3_p & v2313367;
assign v23fb4e6 = hgrant1_p & v12cd9f9 | !hgrant1_p & !v22f991d;
assign v22ef0b3 = hmastlock_p & v22fd29a | !hmastlock_p & !v84561b;
assign v23f4e99 = hbusreq5_p & v23fb9ea | !hbusreq5_p & v84561b;
assign v22f37ba = stateG2_p & v84561b | !stateG2_p & !v863ce5;
assign v230e185 = hbusreq3_p & v22f069f | !hbusreq3_p & !v23f40da;
assign v231008b = hmaster0_p & v84561b | !hmaster0_p & !v1e84038;
assign stateG3_0 = !da3129;
assign v2309d09 = hlock3_p & v22eb665 | !hlock3_p & !v84561b;
assign v230c0da = hbusreq3_p & v22fc70a | !hbusreq3_p & v845620;
assign v23fcabd = jx1_p & v22ef040 | !jx1_p & v22f6fba;
assign v22f1ae5 = hlock0_p & v22eedcf | !hlock0_p & !v84561b;
assign v22f2ed0 = hmaster2_p & v22ec745 | !hmaster2_p & !v22f9a85;
assign v230b59f = hgrant0_p & v84561b | !hgrant0_p & v23f5ce2;
assign abfa28 = busreq_p & v845661 | !busreq_p & v84565f;
assign v22f5ab0 = hbusreq3_p & v22ee918 | !hbusreq3_p & v84561b;
assign v2307a5e = hgrant1_p & v230e28d | !hgrant1_p & v22ef424;
assign v2392a3a = hbusreq3 & v22ee957 | !hbusreq3 & v2306996;
assign v23f1faa = hmaster0_p & v84561b | !hmaster0_p & !v230d513;
assign v23fc850 = hmaster2_p & v84561b | !hmaster2_p & aa8bd6;
assign v22ec61a = hgrant0_p & v22fbf74 | !hgrant0_p & !v23fcda1;
assign v23fca90 = hgrant5_p & v23fcd7c | !hgrant5_p & v230fae0;
assign v230105d = hbusreq3_p & v230e040 | !hbusreq3_p & v84561b;
assign v23fbed3 = hgrant0_p & v23f3a95 | !hgrant0_p & v23fb649;
assign v23f4f3b = hmaster1_p & v22ef607 | !hmaster1_p & v23134bf;
assign v2393508 = hbusreq1_p & v230446f | !hbusreq1_p & !v2301655;
assign v2305128 = hbusreq1 & v191a86f | !hbusreq1 & !v84561b;
assign v230971e = hgrant1_p & v23fbb80 | !hgrant1_p & v150715d;
assign v2311470 = hmaster0_p & v22f73fb | !hmaster0_p & !v23f01d5;
assign v23f745f = hgrant1_p & v84561b | !hgrant1_p & v2306c5e;
assign v23f60e8 = hmaster0_p & v2311504 | !hmaster0_p & v23080f9;
assign v230e100 = hlock5_p & v23f596f | !hlock5_p & v23fcf9d;
assign v8cded5 = hlock3_p & v23fb919 | !hlock3_p & v2303ba8;
assign v22f053b = hmaster0_p & v8f3940 | !hmaster0_p & v23130dd;
assign v2306728 = hmaster2_p & v1aae087 | !hmaster2_p & v23fcf96;
assign v22feb5c = hgrant3_p & v2312919 | !hgrant3_p & v230c37d;
assign v23f4dd0 = hbusreq3 & v230648c | !hbusreq3 & v84561b;
assign v23fc684 = hmaster0_p & v84561b | !hmaster0_p & v23fa882;
assign v2394081 = hlock2_p & v2311255 | !hlock2_p & v22f2718;
assign v22f45a5 = hbusreq5 & v23fb708 | !hbusreq5 & v23fc1ea;
assign v12cd5e1 = hmaster1_p & v22f6b57 | !hmaster1_p & v23fbc64;
assign v23f84f9 = hbusreq4_p & v22f30dc | !hbusreq4_p & v23fbd7d;
assign a7482d = hmaster2_p & v845620 | !hmaster2_p & v22f98fd;
assign v23fa2f1 = hmaster2_p & v2313118 | !hmaster2_p & v84561b;
assign v230d291 = hmaster2_p & v23f77e8 | !hmaster2_p & v23f445f;
assign v23fbddc = hmaster2_p & v22f5820 | !hmaster2_p & !v84561b;
assign v1e83f7c = hbusreq5 & v23fbdb0 | !hbusreq5 & v84561b;
assign v8e28ac = locked_p & v84561b | !locked_p & v22f7919;
assign v191ad59 = hbusreq1 & v845620 | !hbusreq1 & v22ee9be;
assign stateG2 = !v1b87890;
assign v22f16d8 = hlock6_p & v22f8ce6 | !hlock6_p & v23023aa;
assign v23fb89e = hgrant5_p & v84561b | !hgrant5_p & !v23f4a2c;
assign v230b6a4 = hgrant5_p & v22ebe78 | !hgrant5_p & f40dc0;
assign v2308b98 = stateG10_5_p & v22fb706 | !stateG10_5_p & v23126ae;
assign v22f41c4 = hmaster0_p & v22f368e | !hmaster0_p & v23fcf63;
assign v22f9f2a = hmaster0_p & v22f368e | !hmaster0_p & v22eb563;
assign v191abc5 = hgrant1_p & v84561b | !hgrant1_p & v22fafa3;
assign v23fbe74 = hgrant3_p & v84561b | !hgrant3_p & v22fe4a1;
assign v23fa4cb = hmaster2_p & v23fc2d2 | !hmaster2_p & v1b87673;
assign v22fc11b = hlock0_p & v23fc6ac | !hlock0_p & v230d6c1;
assign v2302d69 = hmaster2_p & v23f0bf1 | !hmaster2_p & v23fbaaa;
assign v22ffdc9 = hmaster0_p & v23fb0a1 | !hmaster0_p & !v1aad65a;
assign v22fccf0 = hmaster1_p & v95ca19 | !hmaster1_p & v84561b;
assign v23fc2ff = hbusreq4_p & v23f18a1 | !hbusreq4_p & v23f9193;
assign hgrant3 = !fc8c9b;
assign v23fccd5 = hlock0_p & v2303b9a | !hlock0_p & v2306779;
assign v230a941 = hgrant0_p & v84561b | !hgrant0_p & !v23f84b5;
assign v23f58a6 = hbusreq4_p & v231065b | !hbusreq4_p & v84561b;
assign v23f8988 = hgrant3_p & v23fba96 | !hgrant3_p & v23fbb48;
assign v22edba6 = stateG10_5_p & v23133bb | !stateG10_5_p & a1fbc2;
assign v2305a94 = hmaster2_p & v22edaa4 | !hmaster2_p & !v84561b;
assign v23fbf53 = hbusreq1_p & v22eeb07 | !hbusreq1_p & v23fc0de;
assign v23f659c = hbusreq5 & v23f1207 | !hbusreq5 & v230b1ac;
assign v191ae7e = hgrant3_p & v22f8e29 | !hgrant3_p & v23f08af;
assign v22f8e53 = hmaster0_p & v22f2ffd | !hmaster0_p & !v96c563;
assign v2312c3f = hbusreq3_p & v23132cd | !hbusreq3_p & v84561b;
assign v22ee561 = hbusreq5_p & v22ff732 | !hbusreq5_p & v150705a;
assign v22f583d = hmaster0_p & v23fcab1 | !hmaster0_p & v2392ef6;
assign e1e1ba = hgrant3_p & v84561b | !hgrant3_p & v23f53d0;
assign v22ebc60 = hgrant3_p & v2308af4 | !hgrant3_p & v22edadc;
assign v22f2429 = hbusreq3 & v23f789c | !hbusreq3 & v23fa2ec;
assign v22f5836 = hbusreq5_p & v22f4163 | !hbusreq5_p & a0d50a;
assign v23f7dbe = hbusreq3_p & v23fc01a | !hbusreq3_p & v23fc086;
assign v22fc430 = hbusreq5 & v22f931d | !hbusreq5 & v23fb900;
assign v22ffdd1 = hmaster2_p & v22fd696 | !hmaster2_p & !v84561b;
assign v2300d32 = hgrant5_p & v2302bd3 | !hgrant5_p & v23f2abe;
assign v23fd032 = hmaster0_p & v22f8e29 | !hmaster0_p & v23089fa;
assign v23f3fca = hbusreq5_p & v22f264a | !hbusreq5_p & v84561b;
assign a3ace7 = hbusreq5_p & v84564d | !hbusreq5_p & v23fbbee;
assign v2312919 = hbusreq3_p & v23f558b | !hbusreq3_p & v22fc66c;
assign v23f63dc = hbusreq3 & v22fa9ce | !hbusreq3 & v84561b;
assign v23fbae6 = hmaster2_p & v230665f | !hmaster2_p & v23f79d2;
assign v23fc026 = hbusreq3_p & v22f2bab | !hbusreq3_p & v2303c9d;
assign v22f2a85 = hmaster1_p & v22fe1c8 | !hmaster1_p & v22ede51;
assign v23f1816 = hmaster2_p & v1aae362 | !hmaster2_p & !v13afe3a;
assign v22eea9a = hmaster2_p & v22fc96c | !hmaster2_p & c24eac;
assign v2309ce6 = hbusreq6 & v2301216 | !hbusreq6 & v84561b;
assign v23004f1 = hlock1_p & v22f1b4e | !hlock1_p & !v23056b1;
assign b09263 = hbusreq3_p & v23f3ab0 | !hbusreq3_p & v23fb9d0;
assign v2301274 = hmaster0_p & v22fc8e5 | !hmaster0_p & v22efb8c;
assign v22faba3 = hlock5_p & v84561b | !hlock5_p & !v23fbe12;
assign v22ffc07 = hbusreq1 & v22f36ff | !hbusreq1 & !v84561b;
assign v23f2508 = stateG2_p & v84561b | !stateG2_p & v230e8b8;
assign v23098c0 = hgrant5_p & v84561b | !hgrant5_p & v106af55;
assign v23f9a93 = hbusreq2 & v23105cd | !hbusreq2 & v2312bd0;
assign a476c2 = hgrant2_p & v22f2f87 | !hgrant2_p & v84564d;
assign v23fc646 = hbusreq5_p & v84561b | !hbusreq5_p & v22ecff8;
assign v23fb0eb = hbusreq6_p & v23fcaea | !hbusreq6_p & v23042ca;
assign v22f0c59 = hbusreq1_p & v230928c | !hbusreq1_p & v84561b;
assign v23fc4fc = hmaster2_p & v23f5d34 | !hmaster2_p & !v23043ec;
assign v23fb0e3 = hgrant0_p & v84561b | !hgrant0_p & v2303972;
assign v230299b = hmaster2_p & v230c0b8 | !hmaster2_p & v84561b;
assign v23fbfb6 = hbusreq4_p & v22f6228 | !hbusreq4_p & v23f8a89;
assign v238aeb0 = hbusreq6_p & v23054d5 | !hbusreq6_p & v23f173d;
assign v22f7070 = hmaster2_p & v23f1a8d | !hmaster2_p & v22ff732;
assign v2391d0b = hmaster0_p & v84561b | !hmaster0_p & !v22f1f71;
assign v23022ab = hmaster0_p & v22f3b08 | !hmaster0_p & v230f94d;
assign v23f1803 = hmaster2_p & v2312259 | !hmaster2_p & !v22f4163;
assign v230de5a = stateA1_p & v23fc8d7 | !stateA1_p & !v845649;
assign v2302b5b = hmaster0_p & v23fbcaa | !hmaster0_p & !v96c563;
assign v22f8278 = locked_p & v230841a | !locked_p & v84561b;
assign v94dcdf = hbusreq0 & v23117af | !hbusreq0 & v84564d;
assign v22f1d4f = hbusreq4_p & v22ee8dd | !hbusreq4_p & v22ecd9e;
assign v2310a50 = jx2_p & v2311771 | !jx2_p & v22ebc38;
assign v23fb554 = hbusreq6 & v2306b35 | !hbusreq6 & v22eed0b;
assign v2303efe = hmaster2_p & v23fcbcd | !hmaster2_p & v22f4163;
assign v23fc593 = hbusreq3 & v230a3e6 | !hbusreq3 & v230c781;
assign v23fc01d = hmaster2_p & v2311255 | !hmaster2_p & v22f1389;
assign v23078cd = hlock2_p & v23128a1 | !hlock2_p & v22fa027;
assign v23fcd5f = hmaster2_p & v84561b | !hmaster2_p & v8abd93;
assign v22ffc44 = hbusreq2_p & v22f9927 | !hbusreq2_p & !v84561b;
assign v22f603b = hbusreq3_p & v23fcb31 | !hbusreq3_p & v84561b;
assign v2307e41 = jx0_p & v23f8294 | !jx0_p & v23f1221;
assign v23fba1a = hgrant3_p & v22ed337 | !hgrant3_p & v23f5e22;
assign v23fbad4 = hbusreq6 & v23fc7c0 | !hbusreq6 & v84562f;
assign v22ee7ee = jx3_p & v84561b | !jx3_p & v22f6953;
assign v191b107 = hgrant4_p & v22f08f1 | !hgrant4_p & v23fb11b;
assign v230e191 = hgrant0_p & v22ee956 | !hgrant0_p & v2309939;
assign v23f77c5 = hmaster0_p & v22eddae | !hmaster0_p & v2312ac8;
assign v23051cf = hmaster2_p & v84561b | !hmaster2_p & v845627;
assign v22f04ff = jx1_p & v23fc90b | !jx1_p & v23f17ff;
assign v230749a = hmaster2_p & v2310e40 | !hmaster2_p & v23fc127;
assign v23fc05d = hmaster0_p & v2301b52 | !hmaster0_p & v2312ad7;
assign v22f34bd = hbusreq1_p & v22f7859 | !hbusreq1_p & v17a34f9;
assign v22eeb27 = hmaster2_p & v23080ec | !hmaster2_p & v22f5815;
assign v230cec5 = hbusreq1 & v23fc514 | !hbusreq1 & !v22f91c9;
assign v2312ea0 = hmaster2_p & v22f8ac3 | !hmaster2_p & v84561b;
assign b00a61 = hgrant3_p & v23035c1 | !hgrant3_p & v23fcd4f;
assign v1507118 = hmaster1_p & a0e5e2 | !hmaster1_p & v22f8bd7;
assign v230e0b7 = hbusreq6_p & v230c439 | !hbusreq6_p & v230c2c5;
assign v23fbf37 = hmaster2_p & v22eeb03 | !hmaster2_p & v23f4426;
assign v22ffcbf = hbusreq3_p & v23fc387 | !hbusreq3_p & fc8f95;
assign v2308fb4 = hmaster1_p & v23fc816 | !hmaster1_p & v22ff78b;
assign v22ec98c = hbusreq5_p & v22ede4d | !hbusreq5_p & v2307f27;
assign busreq = v1506af9;
assign v23103f8 = hbusreq6_p & v22f0052 | !hbusreq6_p & !v84561b;
assign v23f880f = hbusreq1_p & v2302b3f | !hbusreq1_p & v2311c5d;
assign v22f52f0 = jx1_p & v23f58ed | !jx1_p & v2303886;
assign v2305792 = hbusreq1 & v84561b | !hbusreq1 & !v22f1e02;
assign v230c963 = hmaster2_p & v23f6b25 | !hmaster2_p & v84564d;
assign v23fceb8 = hbusreq6 & v230a942 | !hbusreq6 & v84561b;
assign v23f7b9b = jx1_p & c26df3 | !jx1_p & v22fbb46;
assign v23fc664 = hbusreq3 & v22f9445 | !hbusreq3 & v22f5b75;
assign v22ef3aa = hmaster0_p & v23fbbc3 | !hmaster0_p & v9799b6;
assign v230d2d1 = hgrant2_p & v2305d69 | !hgrant2_p & v2302973;
assign v12cd8c9 = hlock2_p & v230358b | !hlock2_p & v22fd7dd;
assign v22fe188 = jx1_p & v230327d | !jx1_p & v23fcdcb;
assign v22f3b3c = hgrant5_p & v22f3499 | !hgrant5_p & v22fd767;
assign v23fa2b5 = hbusreq1_p & v23f5ead | !hbusreq1_p & v84561b;
assign v23fcbaa = hbusreq6_p & v106a7cd | !hbusreq6_p & v2308be7;
assign v239154a = hmaster0_p & v23f38d5 | !hmaster0_p & v22f1f71;
assign v22f9bb3 = hbusreq6 & v23fbcad | !hbusreq6 & v23f7933;
assign v23fbeaf = hmaster0_p & v22f82cd | !hmaster0_p & v8ea3a5;
assign v23f82dd = hmaster1_p & v1aadeea | !hmaster1_p & v84561b;
assign v22f4b2c = hmaster0_p & v23fb63f | !hmaster0_p & v22f5164;
assign v2300f19 = hgrant6_p & v23f4edf | !hgrant6_p & v22ef530;
assign v1aae99f = hmaster0_p & v23090fd | !hmaster0_p & v23fba04;
assign v106a7cd = hbusreq4_p & v230c81f | !hbusreq4_p & v84562b;
assign v22f8f27 = hbusreq1 & v23fb9c2 | !hbusreq1 & v84561b;
assign v22f4ef1 = hgrant5_p & v22fe582 | !hgrant5_p & v23fb848;
assign v23f0489 = hbusreq4_p & v2309dce | !hbusreq4_p & v23fbf00;
assign v22f3483 = stateG10_5_p & v22f532c | !stateG10_5_p & !v22ed7a8;
assign v2309c70 = hlock0_p & v22f49c4 | !hlock0_p & v22f2590;
assign v22f88ee = hmaster2_p & v84561b | !hmaster2_p & e1df2d;
assign v23f62d5 = hmaster2_p & v23fbaaa | !hmaster2_p & v22f122e;
assign v2306593 = hbusreq3_p & v2307e0c | !hbusreq3_p & v23fbfd5;
assign v9ce189 = hmaster2_p & v22f337b | !hmaster2_p & v22f8cb7;
assign v22fd6f9 = hbusreq6_p & v23f240a | !hbusreq6_p & v22f8b55;
assign v22ebb51 = hbusreq6 & v23fca0f | !hbusreq6 & !v23fa71e;
assign v2307f2b = hmaster2_p & v22f860b | !hmaster2_p & v23fca9e;
assign v22f2817 = hgrant0_p & e1df2d | !hgrant0_p & v84561b;
assign v230e4ef = hbusreq0 & v23131e8 | !hbusreq0 & !v84561b;
assign v23fb8d6 = hmaster2_p & v230ba09 | !hmaster2_p & v22f6756;
assign v23fcc4e = jx1_p & v22fb49a | !jx1_p & v84561b;
assign v23f5ad6 = hgrant3_p & v23fb63c | !hgrant3_p & v2308b2f;
assign v230997a = hbusreq6_p & v23fbdd2 | !hbusreq6_p & v22fe76b;
assign v2300827 = hbusreq5_p & v23f5043 | !hbusreq5_p & v84564d;
assign v23fc68a = hgrant3_p & v23fc95a | !hgrant3_p & v22fe326;
assign v2312186 = hgrant1_p & v845626 | !hgrant1_p & v22f5a56;
assign v23fbc82 = hlock3_p & v23f3d62 | !hlock3_p & !v84561b;
assign v23f9bcc = jx1_p & v85e5cf | !jx1_p & !v22f6c46;
assign v2312637 = hgrant2_p & v22ee59c | !hgrant2_p & !v23fbd2f;
assign v22f725a = hgrant3_p & v84561b | !hgrant3_p & v2308cec;
assign v22f302f = hlock0_p & v23f51b1 | !hlock0_p & v23f64e5;
assign v23fb89b = hmaster2_p & v23fce22 | !hmaster2_p & v84561b;
assign v22fd41b = hmaster2_p & v230f9db | !hmaster2_p & !v22f661c;
assign v231321e = hbusreq6_p & v22ed8e2 | !hbusreq6_p & v230b11a;
assign v2309192 = hbusreq4_p & v2305f49 | !hbusreq4_p & v23fa14e;
assign v23f6dfb = jx2_p & v23f4a0f | !jx2_p & v2311e58;
assign v22f1553 = stateG10_5_p & v22f532c | !stateG10_5_p & !a1fbb6;
assign c258f4 = hgrant0_p & v22f3643 | !hgrant0_p & v23023c9;
assign v230f713 = hbusreq6 & v23fcb7e | !hbusreq6 & v230e7e4;
assign v23f3e81 = hlock3_p & v23fc7ad | !hlock3_p & v230c5eb;
assign v23fb4a1 = hbusreq3_p & v23f4364 | !hbusreq3_p & v84561b;
assign v23fb6b5 = hgrant3_p & v84561b | !hgrant3_p & v22f176d;
assign v23fab2c = hbusreq5 & v23fcbcd | !hbusreq5 & v23fbffc;
assign v23fb77d = hmaster2_p & v84561b | !hmaster2_p & v23f5240;
assign v23fc343 = hbusreq5_p & b09503 | !hbusreq5_p & v2304cc3;
assign v2301f3a = hbusreq0_p & v84564d | !hbusreq0_p & v2308848;
assign v23fcb9f = hgrant3_p & v22f368e | !hgrant3_p & v230792c;
assign v22f39a8 = hbusreq5_p & bbc337 | !hbusreq5_p & v23fb968;
assign v23046b5 = hlock1_p & v191ace8 | !hlock1_p & v22f5039;
assign v22f9a50 = hgrant3_p & v84561b | !hgrant3_p & v22eb25c;
assign v22f35f5 = hmaster2_p & v845620 | !hmaster2_p & v230b1ac;
assign acdb9d = hbusreq3 & v23fbafc | !hbusreq3 & v230c4ea;
assign v23f2184 = hbusreq4 & v22f8ad3 | !hbusreq4 & v22f5583;
assign v23efed1 = hgrant0_p & v22ffb9d | !hgrant0_p & !v2305258;
assign v22fdb07 = jx3_p & v22f0f7c | !jx3_p & v2312009;
assign v230ed31 = hmaster1_p & v230c7f6 | !hmaster1_p & v22ebe52;
assign v23fcb53 = hgrant0_p & v23fbe41 | !hgrant0_p & v22ff1ee;
assign v23fc21b = hbusreq5_p & v84561b | !hbusreq5_p & v22fa068;
assign v22f9801 = hmaster2_p & v23fb7fc | !hmaster2_p & v230058a;
assign v22ff6f9 = hbusreq1 & v22f4cf3 | !hbusreq1 & !v84561b;
assign v230b4f9 = hbusreq4_p & v22ebd72 | !hbusreq4_p & v22f6aa3;
assign v22ffd9a = hbusreq3 & v2393f95 | !hbusreq3 & v84561b;
assign v23fbb35 = hbusreq0 & v84564d | !hbusreq0 & v84561b;
assign v97b313 = hbusreq4_p & v23f6f14 | !hbusreq4_p & v23067c3;
assign v22f1125 = hlock4_p & v23fbb83 | !hlock4_p & v23fcf11;
assign v23f2b0b = hlock0_p & v22f1b4e | !hlock0_p & v22f1682;
assign v23fcfbc = hbusreq1_p & v23fcaa6 | !hbusreq1_p & v1aad98e;
assign v2302693 = hgrant1_p & f406c6 | !hgrant1_p & !v22f2cb3;
assign v231269d = jx2_p & v23fc403 | !jx2_p & v230ff8a;
assign v23fcd30 = hbusreq1_p & b15a69 | !hbusreq1_p & v22f108e;
assign v231304d = hbusreq6_p & v23041a6 | !hbusreq6_p & !v23f3922;
assign v2304dc2 = hbusreq6 & v22ff982 | !hbusreq6 & v84562f;
assign v22f7b49 = hmaster0_p & v23fb1bb | !hmaster0_p & v13afb04;
assign v22f0635 = hbusreq4_p & v23f420c | !hbusreq4_p & !v230f549;
assign v23fca19 = hmastlock_p & v230932e | !hmastlock_p & !v84561b;
assign v2300004 = hmaster2_p & v22f53c0 | !hmaster2_p & v23001d6;
assign v22f0a24 = hmaster2_p & v106af73 | !hmaster2_p & v230320e;
assign a25b7d = hbusreq6 & v12cd4c5 | !hbusreq6 & v84561b;
assign v23f9789 = hlock5_p & v22f0945 | !hlock5_p & !v845636;
assign v22f37e8 = hmaster0_p & v23fc282 | !hmaster0_p & v22fc5d2;
assign v23fb720 = stateG10_5_p & v22f41ee | !stateG10_5_p & v22f56d2;
assign bd9c50 = hbusreq2_p & v23fbd99 | !hbusreq2_p & v84561b;
assign v23fcb36 = hbusreq3_p & bd766b | !hbusreq3_p & v2306ee6;
assign v12cc315 = hgrant4_p & v84561b | !hgrant4_p & v23fcb57;
assign v23fc52d = hmaster2_p & v845620 | !hmaster2_p & v230dbc9;
assign v2307632 = hmaster2_p & v23fc969 | !hmaster2_p & v23124cc;
assign a51d7a = hbusreq0_p & v2303996 | !hbusreq0_p & v84561b;
assign v23fc679 = jx1_p & v23fcebe | !jx1_p & v23fc42e;
assign v23099fc = hmaster2_p & v23fbeb0 | !hmaster2_p & v23035ba;
assign v22feb47 = hready & v22f7919 | !hready & !v84561b;
assign f40dab = hbusreq5_p & v23f4ccb | !hbusreq5_p & v22eb72a;
assign v191aa95 = hbusreq2_p & v22f8214 | !hbusreq2_p & v84561b;
assign v22fe0ee = hbusreq0_p & v22f9e5b | !hbusreq0_p & !v22fc3ed;
assign v23f439b = hgrant3_p & v84564d | !hgrant3_p & !v23f2f5d;
assign f40dc0 = hbusreq5_p & v22f533e | !hbusreq5_p & v22fbfe5;
assign v2302875 = hmaster0_p & v22f2abb | !hmaster0_p & v230fc1f;
assign v23fc243 = hlock5_p & v84561b | !hlock5_p & v15070f7;
assign v23f70e3 = hlock3_p & v22fecb6 | !hlock3_p & v23f8e34;
assign v2306de4 = hbusreq3_p & v22f39d3 | !hbusreq3_p & v84561b;
assign v23f4827 = hmaster2_p & v23031c2 | !hmaster2_p & v2310754;
assign v23fc0a7 = hmaster1_p & v23fb6bd | !hmaster1_p & v23efec0;
assign v23f53e4 = hbusreq5_p & v22f1ae5 | !hbusreq5_p & v22f9d17;
assign v230f4e5 = hbusreq3 & v230dcf6 | !hbusreq3 & !v84561b;
assign v23fbca1 = hbusreq3_p & v12cd4be | !hbusreq3_p & v22fb49d;
assign v230db14 = hgrant5_p & v230ff42 | !hgrant5_p & !v22f0ddd;
assign v2392868 = hbusreq3_p & v22f4a4f | !hbusreq3_p & v23fcd74;
assign v230e551 = hbusreq0_p & v84562a | !hbusreq0_p & v22eedf9;
assign v23f1c0f = hmaster2_p & v106ae19 | !hmaster2_p & !v22feafc;
assign v22f3998 = hbusreq6 & v230aa96 | !hbusreq6 & !v230bc39;
assign v22f15fe = hbusreq2 & v22fc569 | !hbusreq2 & !v84561b;
assign v2303edc = hbusreq3 & v23f374e | !hbusreq3 & v84561b;
assign v23fcba7 = hlock0_p & v1b87673 | !hlock0_p & !v84561b;
assign v22fb009 = hmaster2_p & v23128a1 | !hmaster2_p & v230984f;
assign v23fc8a2 = hlock6_p & v230b6d9 | !hlock6_p & v22f86d2;
assign v23f3297 = hmaster2_p & v23fc3f2 | !hmaster2_p & v845622;
assign v22f8b55 = hbusreq4_p & v2304c86 | !hbusreq4_p & v23032db;
assign e1c7f2 = hmaster0_p & v230741d | !hmaster0_p & !v23130d6;
assign v22f7564 = hmaster2_p & v23fcaf0 | !hmaster2_p & v23112d5;
assign v230b573 = hlock0_p & v2309066 | !hlock0_p & !v230e40a;
assign v22ef9d0 = hgrant3_p & v84561b | !hgrant3_p & v22f7ab4;
assign v2312ae4 = hmaster2_p & v22ff308 | !hmaster2_p & v22ffe8d;
assign v23f6404 = hmaster2_p & v84561b | !hmaster2_p & !v23fd021;
assign v23fb922 = hmaster2_p & v230c2f3 | !hmaster2_p & v2310d04;
assign v23fcd28 = hmaster2_p & v2311810 | !hmaster2_p & v22eb377;
assign v23fc8f3 = hbusreq4_p & v2301cf4 | !hbusreq4_p & !v84561b;
assign v2301bda = hmaster1_p & bd74b6 | !hmaster1_p & !v106a7d3;
assign v230faaf = hbusreq2_p & v22f8aeb | !hbusreq2_p & !v230f2f5;
assign v23f9a8e = hlock6_p & v23fcc2f | !hlock6_p & v23915cb;
assign v23fc3f7 = hlock0_p & v22ec53b | !hlock0_p & v845620;
assign v23052cc = hgrant0_p & v2301e25 | !hgrant0_p & v22fd3f7;
assign v230a91b = hmaster2_p & v106ae43 | !hmaster2_p & v84561b;
assign v23f6f14 = hmaster0_p & v22eef3f | !hmaster0_p & !v23fc9be;
assign v23f4201 = hbusreq1_p & v191a86f | !hbusreq1_p & !v23f55ea;
assign v2309871 = hlock0_p & v191aa68 | !hlock0_p & v23fce86;
assign v22edec8 = hmaster0_p & v23fa8d8 | !hmaster0_p & v23013a2;
assign v23fbe50 = hbusreq3_p & v2304904 | !hbusreq3_p & v22eec2a;
assign v22edf62 = hbusreq1_p & v2309fb1 | !hbusreq1_p & v2304574;
assign v23fc404 = hmaster2_p & v22f2b78 | !hmaster2_p & v22f7b47;
assign f40c96 = hmaster2_p & v84561b | !hmaster2_p & v2300ac2;
assign v23fcdca = jx2_p & v191aa98 | !jx2_p & v23fb21c;
assign v23f3561 = hmaster0_p & v22ef1eb | !hmaster0_p & v22ebed1;
assign v23068bb = hbusreq4_p & v23fb670 | !hbusreq4_p & !v2302b93;
assign v22f44d0 = hmaster0_p & v230d6ca | !hmaster0_p & v23002d1;
assign v22f8e29 = hbusreq3_p & v84561b | !hbusreq3_p & v12cc2ef;
assign v2302348 = hbusreq4_p & v2300834 | !hbusreq4_p & v230adbf;
assign v2306b35 = hlock3_p & v23fba94 | !hlock3_p & !v84561b;
assign v23fc1ea = hlock0_p & v2300a72 | !hlock0_p & v84561b;
assign v191ac40 = hbusreq3_p & v2302177 | !hbusreq3_p & v2304bc1;
assign v231066c = hmastlock_p & v22f0eec | !hmastlock_p & v84561b;
assign v230c79d = hmaster2_p & v84561b | !hmaster2_p & v2305c1f;
assign v23f5201 = jx0_p & v2303cae | !jx0_p & !v22f658c;
assign v23126b1 = hmaster2_p & v22f954f | !hmaster2_p & v231007b;
assign v23f55ae = hmaster2_p & v9d8aae | !hmaster2_p & !v2312f7e;
assign v2306838 = hmaster2_p & v22fc8e5 | !hmaster2_p & v23f5be9;
assign v23f494b = hbusreq5_p & v22ff732 | !hbusreq5_p & v22f43fb;
assign v2308a32 = hbusreq3 & v23f2873 | !hbusreq3 & !v84561b;
assign v23fc5d3 = hgrant3_p & v84561b | !hgrant3_p & v22ff5ea;
assign v22fe76b = hmaster0_p & v22fa0ec | !hmaster0_p & !v23fb661;
assign v22fb4de = hgrant1_p & v84561b | !hgrant1_p & !v23046d0;
assign b9d049 = hbusreq1_p & v22ee0c4 | !hbusreq1_p & v191ad69;
assign v22ec191 = hgrant3_p & v22fbd88 | !hgrant3_p & v22eee6a;
assign v23fc40a = hbusreq4 & v23fcc49 | !hbusreq4 & v84561b;
assign v23f2dd4 = hmaster2_p & v84561b | !hmaster2_p & v23fcb1a;
assign v23fcaab = hbusreq3_p & v2306aef | !hbusreq3_p & v2309d97;
assign v22f13cb = hbusreq0 & v23fa63b | !hbusreq0 & !v23f3978;
assign v23fb935 = hbusreq4_p & v845637 | !hbusreq4_p & v23fa36c;
assign v23019b7 = hgrant3_p & v22f118e | !hgrant3_p & !v23fb61d;
assign v2311b9e = hmaster0_p & v22f2f3e | !hmaster0_p & v23fbe02;
assign v22fdce0 = hbusreq1 & v22f4587 | !hbusreq1 & !v23fc614;
assign v23fc03d = hbusreq4_p & v22f41c4 | !hbusreq4_p & v230ff65;
assign v230a1fa = hbusreq4_p & v84561b | !hbusreq4_p & v22f8e29;
assign v2307dae = hmaster0_p & v23f72e4 | !hmaster0_p & v23fbe2a;
assign v23f7c32 = hbusreq6 & v22f9833 | !hbusreq6 & v22f2ca2;
assign v22fa652 = hgrant1_p & v12cd9f9 | !hgrant1_p & v22f6ac9;
assign v22f64de = hgrant5_p & v84561b | !hgrant5_p & v230979f;
assign v12cda8f = hmaster0_p & v23fcbdc | !hmaster0_p & v230f0de;
assign v23f8772 = hbusreq1 & v23fc35a | !hbusreq1 & v23f3cb8;
assign v23fc369 = hbusreq4 & v22f91b6 | !hbusreq4 & v84561b;
assign v23fb04e = hbusreq3 & v23089a5 | !hbusreq3 & v84564d;
assign v22f1fca = hbusreq3 & v22ed4e1 | !hbusreq3 & v84561b;
assign v23f5af8 = hbusreq4 & v23fb0c0 | !hbusreq4 & v84561b;
assign v22f2ffd = hgrant3_p & v22ee657 | !hgrant3_p & v23fbd90;
assign v23fc2fc = hbusreq0 & e1ddd0 | !hbusreq0 & v84561b;
assign v230560c = hmaster0_p & v22fb89a | !hmaster0_p & !v22f90af;
assign v23fa71e = hmaster2_p & v23f4c57 | !hmaster2_p & !v22f8bd0;
assign v22f4ae7 = hlock6_p & v23f1b7a | !hlock6_p & !v84561b;
assign v23f4d72 = hgrant5_p & v2303c12 | !hgrant5_p & v23fb10d;
assign v23035d7 = hgrant1_p & v2312a8d | !hgrant1_p & v23fa9c5;
assign v22f297d = hmaster0_p & v2308363 | !hmaster0_p & v22f5216;
assign v2301c2e = hmaster2_p & v2300934 | !hmaster2_p & !v23fcd14;
assign v23132cd = hbusreq3 & v23fcdc5 | !hbusreq3 & v84561b;
assign v230c91d = hmaster1_p & v22ef757 | !hmaster1_p & !v231396f;
assign d49f2b = hbusreq3_p & v23fc7a7 | !hbusreq3_p & v22f0a24;
assign v23f420d = hmaster2_p & v23fbeb0 | !hmaster2_p & v84561b;
assign v23fc01e = hlock0_p & v23fc976 | !hlock0_p & v22ec335;
assign v23fc4ce = hbusreq6_p & v230e628 | !hbusreq6_p & v84561b;
assign v23019e7 = hbusreq2 & v230088c | !hbusreq2 & v84562b;
assign v22f5235 = hmaster2_p & b50a75 | !hmaster2_p & b00a78;
assign v22ebf1f = hbusreq0_p & v2310657 | !hbusreq0_p & v84561b;
assign v22f5388 = hbusreq3 & v22f0545 | !hbusreq3 & !v84561b;
assign v23102d5 = hbusreq1_p & v23fbf44 | !hbusreq1_p & v84561b;
assign v230abb1 = hbusreq1 & v84561b | !hbusreq1 & !v23068a9;
assign v23fc970 = hmaster0_p & v2300562 | !hmaster0_p & v231242a;
assign v230d2d8 = hmaster2_p & v84561b | !hmaster2_p & v22f3643;
assign v22ec060 = hmaster2_p & v845620 | !hmaster2_p & v2313476;
assign v23fc8bb = hbusreq1 & v23f8deb | !hbusreq1 & v23f3472;
assign v22fdcc5 = hmaster0_p & v230fbc5 | !hmaster0_p & v2307b17;
assign v22fd00f = hbusreq1 & v23fbfd0 | !hbusreq1 & v84561b;
assign v230f18c = hgrant3_p & v84561b | !hgrant3_p & !v23f3346;
assign v23fb6e3 = hbusreq5_p & v23fd067 | !hbusreq5_p & !v84561b;
assign v230f848 = hlock0_p & v106ae19 | !hlock0_p & v22fd5dd;
assign v23fc9d8 = hbusreq6 & v22fa8c6 | !hbusreq6 & v22f7347;
assign v22ec522 = hgrant5_p & v23fbf1a | !hgrant5_p & v23fc0c2;
assign v23fbb42 = hgrant3_p & v230d8af | !hgrant3_p & v22eb49d;
assign v23125ee = hgrant3_p & v23fcf5e | !hgrant3_p & v230f578;
assign v22f57d4 = hbusreq3_p & v23fba74 | !hbusreq3_p & v23fb906;
assign v23fb5a2 = hgrant5_p & v23fc26e | !hgrant5_p & v23fbdf1;
assign v23f6927 = hmaster2_p & v22f954f | !hmaster2_p & v2309456;
assign v2306fb7 = hmaster2_p & v23f024e | !hmaster2_p & v2300271;
assign v23fca0c = hbusreq1_p & v23fca96 | !hbusreq1_p & a1fe03;
assign v22f70bd = hmaster0_p & b00aa6 | !hmaster0_p & v230e5da;
assign v22ff6a8 = hbusreq3_p & v23fc6c2 | !hbusreq3_p & v23f41c2;
assign v23fb73d = hbusreq3_p & v22fec20 | !hbusreq3_p & v9ad58e;
assign v906d1d = hlock1_p & v23fbfe5 | !hlock1_p & v22ebf17;
assign v23f8536 = hbusreq1_p & v1aad5a0 | !hbusreq1_p & v22f7241;
assign v22edd3f = hbusreq1_p & b09503 | !hbusreq1_p & v23fc343;
assign v23f67d3 = hbusreq6 & v22ed684 | !hbusreq6 & v23fcf81;
assign v23051ab = hgrant6_p & v23fca17 | !hgrant6_p & v2300bc5;
assign v2309221 = hbusreq0 & v8d360e | !hbusreq0 & !v84561b;
assign v23f57a2 = hbusreq1_p & v23f7eaa | !hbusreq1_p & !v84561b;
assign v22eb01f = hmaster0_p & v2303513 | !hmaster0_p & v2309889;
assign v23f24c0 = jx1_p & v84561b | !jx1_p & v23fb98b;
assign v23fc89d = hmaster0_p & v919672 | !hmaster0_p & v230b8fe;
assign v22f8da4 = hbusreq3 & v22f8cb7 | !hbusreq3 & v84561b;
assign v2392f6b = hbusreq5_p & v230446f | !hbusreq5_p & !v2301655;
assign v230bbda = hgrant3_p & v8ea3a5 | !hgrant3_p & v2307517;
assign v2310ad7 = hlock2_p & v22f60c6 | !hlock2_p & !v84561b;
assign v23107f9 = hbusreq3 & v22eaafa | !hbusreq3 & v22fa415;
assign v2306d5c = stateA1_p & v22ec1cb | !stateA1_p & v84561b;
assign v12cd4da = hmaster0_p & v23fc932 | !hmaster0_p & v230f0de;
assign v23fb624 = hgrant1_p & v845626 | !hgrant1_p & v2393aca;
assign v22f8e08 = hbusreq3 & v23fc48f | !hbusreq3 & v23fcc2e;
assign v230e962 = hmaster0_p & v23fceb8 | !hmaster0_p & v230851f;
assign v2309377 = hlock2_p & v23f5cb3 | !hlock2_p & v23fbfb9;
assign v22ec150 = hmaster0_p & v22f368e | !hmaster0_p & v23fc975;
assign v231324f = hgrant3_p & v22ee62f | !hgrant3_p & v22f8477;
assign v23f412d = hmaster2_p & v2310754 | !hmaster2_p & v230d3f5;
assign v230fe71 = hmaster1_p & v23f5470 | !hmaster1_p & v23fc844;
assign v230dc56 = hlock0_p & v22ede4d | !hlock0_p & v84561b;
assign v106ae5a = hbusreq6 & v22fa6b2 | !hbusreq6 & !v84561b;
assign v23fc263 = hbusreq4 & v22f39f4 | !hbusreq4 & v22ef5f1;
assign v2302b81 = hbusreq4_p & v22f8c01 | !hbusreq4_p & v8958ff;
assign v22eeab9 = hmaster0_p & v2392d61 | !hmaster0_p & v23f6d65;
assign v23089c5 = hmaster2_p & bd74c0 | !hmaster2_p & v1aae98c;
assign v23fbebe = hmaster2_p & v1506fe9 | !hmaster2_p & v22ff732;
assign v23f90b2 = hbusreq3_p & v22ff12b | !hbusreq3_p & v84561b;
assign v23fb9b2 = hbusreq0 & v13afe3a | !hbusreq0 & !v22fbb8a;
assign v2313549 = hbusreq1_p & v22faa0e | !hbusreq1_p & v84561b;
assign v22f7277 = hlock4_p & v22f7a1d | !hlock4_p & v23fc937;
assign v23fba3f = hmaster0_p & v23fc802 | !hmaster0_p & b00a61;
assign v22ff2c4 = hbusreq6 & v230d3c2 | !hbusreq6 & v84561b;
assign v23fb4b4 = hmaster2_p & v22f1b4e | !hmaster2_p & v22ffbb3;
assign v23f4bfc = hmaster2_p & fc8c27 | !hmaster2_p & v230e821;
assign v230308e = hbusreq5 & v13afe3a | !hbusreq5 & !v22f9a51;
assign v22f2835 = jx0_p & v13afed6 | !jx0_p & e1e35b;
assign v23107cf = hbusreq3_p & v23fb18e | !hbusreq3_p & !v861565;
assign v22f0102 = hgrant3_p & v23fceca | !hgrant3_p & v22f17ed;
assign v22fbd88 = hbusreq3_p & v23fa4bb | !hbusreq3_p & v23f2bbf;
assign v23007f9 = hmaster2_p & v22ee0c4 | !hmaster2_p & v84561b;
assign v23fcb8f = jx1_p & v22ec012 | !jx1_p & v84561b;
assign v17a34ff = locked_p & v84561b | !locked_p & !v845647;
assign v22f803d = hmaster2_p & v23fc71d | !hmaster2_p & v23f9789;
assign v238ab71 = hgrant3_p & v84561b | !hgrant3_p & v230c0b4;
assign v191ae81 = hbusreq5_p & v84561b | !hbusreq5_p & v230278e;
assign v23fcc91 = hmaster2_p & v22fc8c8 | !hmaster2_p & v22fe421;
assign v22f7ec9 = hmaster2_p & v191a86f | !hmaster2_p & v22eb5b3;
assign v23fcb2b = hmaster2_p & v2309891 | !hmaster2_p & v84561b;
assign v22f46ff = hbusreq3_p & v22f7dbc | !hbusreq3_p & v2305aa9;
assign v23fcd3a = hgrant5_p & v23fbcc0 | !hgrant5_p & fc8f72;
assign v23f6765 = hgrant2_p & v84562a | !hgrant2_p & v23f44b1;
assign v23f23f4 = hmaster1_p & v23fce29 | !hmaster1_p & v22fdbac;
assign v2303fa7 = hbusreq6_p & v23fca1b | !hbusreq6_p & v23fb777;
assign v23f1ca1 = hbusreq0_p & v23fbef7 | !hbusreq0_p & v84561b;
assign v22fa0b2 = hmaster1_p & v23f9a3a | !hmaster1_p & v230c94b;
assign v23fb47d = hgrant6_p & v23135cf | !hgrant6_p & v2306854;
assign a452a3 = jx1_p & v23fc57c | !jx1_p & v23119b0;
assign v22fb428 = hbusreq3 & v23fcfb4 | !hbusreq3 & v23fa2ec;
assign v2310283 = hbusreq5 & v23f366d | !hbusreq5 & v2392fa3;
assign v23018ac = hgrant3_p & v23f2602 | !hgrant3_p & v23f4a02;
assign v2312da9 = hgrant3_p & v23fb137 | !hgrant3_p & v23fcafd;
assign v23f0625 = hbusreq1_p & v230ae09 | !hbusreq1_p & v23f7f77;
assign v23fcf9d = hbusreq5 & v22f0073 | !hbusreq5 & !v22f4527;
assign v23fb886 = hbusreq4_p & v23f5dfe | !hbusreq4_p & v22f758c;
assign v23fce1e = hlock3_p & v23021af | !hlock3_p & !v84561b;
assign v2304070 = hmaster0_p & v2307b25 | !hmaster0_p & v23fc22f;
assign v22f8aa0 = hbusreq4_p & v22f7375 | !hbusreq4_p & v2303c5b;
assign v2313230 = hmaster0_p & v919672 | !hmaster0_p & v23efa84;
assign v22ff882 = hbusreq3_p & v23fb1b9 | !hbusreq3_p & v84561b;
assign v22f742b = hgrant1_p & v23f3c2a | !hgrant1_p & v23f75ce;
assign v22ecde7 = hgrant3_p & v17a34ff | !hgrant3_p & v23135cc;
assign da3886 = hmaster2_p & v22ed85a | !hmaster2_p & v2300de3;
assign v23f73ba = hmaster2_p & v2310d04 | !hmaster2_p & v22ebb79;
assign v23f5df1 = hbusreq6_p & v22fd364 | !hbusreq6_p & v22f758c;
assign v22fdabc = hlock5_p & v84561b | !hlock5_p & v230db4d;
assign v22fdb25 = hmaster1_p & v23f38b1 | !hmaster1_p & v22fbb7f;
assign v230ed27 = hlock1_p & a1b802 | !hlock1_p & !v84561b;
assign v23fbc86 = hmaster2_p & v23fbe80 | !hmaster2_p & !v23043ec;
assign v22fab6a = hbusreq1 & v2304009 | !hbusreq1 & v23fb966;
assign v23fc5ff = hbusreq1_p & v2308e85 | !hbusreq1_p & v84561b;
assign v23f1207 = hready & v84561b | !hready & v23f2f45;
assign v2392aaa = hbusreq4 & v23f1812 | !hbusreq4 & v22fc963;
assign v22eb83a = jx0_p & v22fbb46 | !jx0_p & v230b6fc;
assign v22f3dab = hmaster2_p & v2312c77 | !hmaster2_p & v23fbfa7;
assign v22f4faf = stateG10_5_p & v23f3eed | !stateG10_5_p & v22f0945;
assign v23fcea9 = hbusreq5_p & v84561b | !hbusreq5_p & !v2309aaa;
assign v23036ca = hbusreq2_p & v2301655 | !hbusreq2_p & !v84561b;
assign v22f6683 = hbusreq2 & v22feb47 | !hbusreq2 & v845620;
assign v912a31 = stateA1_p & v23f54be | !stateA1_p & v84561b;
assign v2309840 = hmaster0_p & v23fc282 | !hmaster0_p & v230b3d5;
assign v23fc34b = jx1_p & v2306a0e | !jx1_p & v22eb7cc;
assign v2392b3d = hmaster2_p & v23f9789 | !hmaster2_p & b60876;
assign v22f9554 = hmaster1_p & v230af0f | !hmaster1_p & !v23f49cd;
assign v2305c43 = hbusreq4_p & v23fb8f4 | !hbusreq4_p & !v23f216d;
assign v23f88e6 = hbusreq6 & v23f2bc5 | !hbusreq6 & v84561b;
assign v23fc75c = hbusreq4 & v230a67e | !hbusreq4 & v23fcfad;
assign v2302ca3 = hburst1 & v84561b | !hburst1 & v84563e;
assign v22f6f2d = hlock6_p & v84561b | !hlock6_p & v23fc8f3;
assign v23fbdd2 = hmaster0_p & v22fa0ec | !hmaster0_p & v22ecb12;
assign v2305719 = hbusreq3_p & v23f704d | !hbusreq3_p & v2313131;
assign v23fb62c = hbusreq3_p & v84564d | !hbusreq3_p & !v1e840fa;
assign v23fc676 = hmaster2_p & v2310434 | !hmaster2_p & v23fb8a0;
assign v23fc329 = hmaster0_p & v2300d5f | !hmaster0_p & v22f8420;
assign v2302efc = hmaster0_p & f4066e | !hmaster0_p & v2308dcf;
assign v22f0c1b = hbusreq1 & v22f1a26 | !hbusreq1 & v84561b;
assign v2312ea7 = hready & v22fa2de | !hready & !v22fe9e0;
assign v22ffb52 = hgrant2_p & v2310116 | !hgrant2_p & be4ff1;
assign v2312325 = hbusreq4_p & v2304070 | !hbusreq4_p & v84561b;
assign v22eb57a = hbusreq3_p & v22f7e19 | !hbusreq3_p & !v84561b;
assign v23f7d1a = hbusreq3_p & v2307c0c | !hbusreq3_p & v230dc73;
assign v23018a8 = hmaster2_p & v22f343b | !hmaster2_p & v230446f;
assign v23fba24 = hgrant5_p & v22ff463 | !hgrant5_p & v23fbe4c;
assign v230fbc5 = hbusreq3_p & ae78a6 | !hbusreq3_p & v230ced0;
assign v23f2a7c = hgrant5_p & v22f9049 | !hgrant5_p & !v2313618;
assign v23f60ba = hmaster0_p & v84561b | !hmaster0_p & !f405e4;
assign v22ecd97 = hbusreq1_p & v23fb9c5 | !hbusreq1_p & v2309c93;
assign v23fbb4a = hbusreq4 & v23f363f | !hbusreq4 & v84561b;
assign v1e8471c = hgrant1_p & v2303f37 | !hgrant1_p & v995fa2;
assign v23fc0ce = hlock0_p & v22fd30c | !hlock0_p & v23fc3a7;
assign v23fba5a = hbusreq3 & v22febe7 | !hbusreq3 & v84561b;
assign v230d91f = hmaster0_p & v2303bee | !hmaster0_p & v23f535c;
assign v230177d = hburst0_p & v23fc116 | !hburst0_p & !v23fb4a4;
assign v23f3d5b = hmaster2_p & v2311d0c | !hmaster2_p & v23fbfb9;
assign v22f0db9 = hmaster0_p & v22feec8 | !hmaster0_p & v23fb5a4;
assign v230d533 = hgrant1_p & v230ffae | !hgrant1_p & !v84561b;
assign v230b516 = hready_p & v2308c4d | !hready_p & !v23fb842;
assign v8920c5 = hmaster0_p & v84564d | !hmaster0_p & v22f9bb3;
assign v22fe56f = hmaster0_p & v23fc23e | !hmaster0_p & v23fcd0d;
assign v22fddc8 = hgrant0_p & v23fbcb2 | !hgrant0_p & !v23f0ded;
assign v22f59bd = hmaster0_p & v22f2c8a | !hmaster0_p & v23fc815;
assign v230ba79 = hgrant3_p & v23fc975 | !hgrant3_p & v22f5495;
assign v22f3c11 = hmaster2_p & v22ff90b | !hmaster2_p & v2305d2f;
assign a0b7a3 = hmaster2_p & v23fb1e5 | !hmaster2_p & !v22ec08f;
assign v22f9657 = hmaster2_p & v23fcc10 | !hmaster2_p & v22fc34e;
assign v22fd2f5 = stateG10_5_p & v22fa707 | !stateG10_5_p & v22f3643;
assign v23fb1a4 = hready & v22f4f14 | !hready & v2302937;
assign v230fff1 = hmastlock_p & v2312d48 | !hmastlock_p & !v84561b;
assign v23fb873 = hbusreq5 & v22fc34e | !hbusreq5 & v84561b;
assign v230f5d0 = hlock0_p & v23fb5ad | !hlock0_p & v22fe009;
assign v2310812 = hbusreq1 & v23f3724 | !hbusreq1 & v84561b;
assign v22f13e3 = hbusreq1_p & v2392f6b | !hbusreq1_p & bd7476;
assign v23046a7 = hgrant6_p & v84563a | !hgrant6_p & v2310a50;
assign v23fb084 = hbusreq3 & v2302aac | !hbusreq3 & v23f30cf;
assign v22ed220 = hmaster1_p & bd953c | !hmaster1_p & v22fc163;
assign v22eaaef = hbusreq1_p & v2312351 | !hbusreq1_p & v23fc190;
assign v22f09b1 = hlock6_p & v84561b | !hlock6_p & v23fcc84;
assign v22ec339 = hgrant3_p & v84561b | !hgrant3_p & v23f8e25;
assign e1e75d = hlock6_p & v84561b | !hlock6_p & v23051a9;
assign v23efdd4 = hbusreq0 & v22f7f74 | !hbusreq0 & v84561b;
assign v23034c9 = hlock3_p & v22f065f | !hlock3_p & v22fdda4;
assign v23fbc6e = hmaster0_p & v23fced1 | !hmaster0_p & ab39f4;
assign v22ff38e = hbusreq0 & v1aae56f | !hbusreq0 & v84561b;
assign v22f53a6 = hready & v22fbf54 | !hready & v230c899;
assign v22f8f91 = hmastlock_p & v23fbc7d | !hmastlock_p & v84561b;
assign v23f47b3 = hmaster2_p & v97b973 | !hmaster2_p & !v230aef0;
assign v22f2487 = hbusreq4_p & v23fbcd2 | !hbusreq4_p & v23fc9b4;
assign v23f0865 = hbusreq1_p & v230ef1c | !hbusreq1_p & !v84561b;
assign v23122cf = hmaster2_p & v23fb906 | !hmaster2_p & v23fcd00;
assign v23fbaf6 = jx0_p & v23fc34b | !jx0_p & c17224;
assign v1aad3ae = hbusreq5_p & v2313618 | !hbusreq5_p & v23fc6f7;
assign v191b212 = hgrant3_p & v22f2ca2 | !hgrant3_p & v23fb7da;
assign v2304494 = hready & v84561b | !hready & v13afe3a;
assign v22f9280 = hmaster2_p & v2304536 | !hmaster2_p & v84561b;
assign v23fca55 = hbusreq3_p & v23fbc9a | !hbusreq3_p & v84561b;
assign v22edf79 = hbusreq3_p & v22f3092 | !hbusreq3_p & v23fc957;
assign v23f4bc2 = hbusreq3_p & v22f61f6 | !hbusreq3_p & v22fa6ab;
assign v22f766b = hgrant1_p & v230571c | !hgrant1_p & !v23fc3b3;
assign v230f0de = hgrant3_p & v84562e | !hgrant3_p & v23fba9a;
assign v22f8ad5 = hbusreq3 & v2306f3c | !hbusreq3 & v22fe2dc;
assign v22eb0b1 = hbusreq3_p & v23fb81f | !hbusreq3_p & v230d3a4;
assign v230d680 = hbusreq0_p & v23934e0 | !hbusreq0_p & v23f4462;
assign v230ba09 = hgrant1_p & v22f3ed0 | !hgrant1_p & v23f0903;
assign v2311a1d = hbusreq2_p & v23fce8d | !hbusreq2_p & v84561b;
assign v23fbe44 = hgrant1_p & v23fb6ff | !hgrant1_p & v2392fd0;
assign v23fbec8 = hbusreq2 & v191a86f | !hbusreq2 & !v84561b;
assign v230c84d = hlock4_p & v23f9465 | !hlock4_p & v22ed48e;
assign v2393c3a = hgrant0_p & v22ee4fe | !hgrant0_p & !v23fb1a6;
assign v23fc556 = hbusreq2_p & v22fa821 | !hbusreq2_p & !v84561b;
assign v230e9f8 = hlock6_p & v22fc398 | !hlock6_p & v845637;
assign v2313504 = hbusreq4_p & v23f8b5b | !hbusreq4_p & v23f7891;
assign v23f2422 = hbusreq2 & v2308e63 | !hbusreq2 & !v84561b;
assign v22f6228 = hmaster0_p & v22ebe46 | !hmaster0_p & v22fe4ea;
assign v22efa8c = hbusreq4 & v2312888 | !hbusreq4 & v22f475e;
assign v22f13d8 = hgrant3_p & v2310ec8 | !hgrant3_p & v9f5c3c;
assign v22ed335 = hmaster0_p & v15071c7 | !hmaster0_p & v23fb6ed;
assign v22f0c90 = hbusreq1_p & v2313476 | !hbusreq1_p & v845620;
assign v23fc320 = hbusreq4 & v22f8e2f | !hbusreq4 & v23fbcbf;
assign v23fccf8 = hgrant5_p & v23fba3d | !hgrant5_p & v23077c2;
assign v23fb24f = hbusreq5_p & v845636 | !hbusreq5_p & v23fce91;
assign v22f6917 = hmaster2_p & v845647 | !hmaster2_p & !v17a34ff;
assign v22f5218 = hbusreq3_p & v84564d | !hbusreq3_p & v84561b;
assign v90aa06 = stateG10_5_p & v22fd767 | !stateG10_5_p & v22eb377;
assign v23facdf = hgrant5_p & v2391c72 | !hgrant5_p & !a6a2f9;
assign bd75f3 = hbusreq6 & v23f7d1a | !hbusreq6 & v150718d;
assign v2310d44 = hlock2_p & v22f7f74 | !hlock2_p & v84561b;
assign v230397f = hbusreq5 & v22fea89 | !hbusreq5 & !v84561b;
assign v12cd3a7 = hmaster2_p & b9d013 | !hmaster2_p & !v23fb9cf;
assign v23f8410 = hmaster1_p & v23fbc3d | !hmaster1_p & !v23f49cd;
assign v23f5cfe = hmaster2_p & v1aadac4 | !hmaster2_p & v23fce4c;
assign v22fe5b1 = hbusreq2_p & v23f2422 | !hbusreq2_p & !v84561b;
assign v22fd79e = hbusreq2 & v2394081 | !hbusreq2 & v84561b;
assign v23111a4 = hbusreq4_p & v23fbbc5 | !hbusreq4_p & bd7ae5;
assign v2304d64 = hgrant1_p & v22eb097 | !hgrant1_p & !v23fc3b3;
assign bf7e60 = hlock3_p & v22f7e19 | !hlock3_p & !v84561b;
assign v22eed25 = hmaster0_p & v22fb7e0 | !hmaster0_p & v22fb417;
assign v22f5d1e = stateG10_5_p & v2305a1c | !stateG10_5_p & v22eb3c2;
assign v23fc7dc = hmaster0_p & v845632 | !hmaster0_p & v23088db;
assign v23fb0a8 = hbusreq4 & v23f3d02 | !hbusreq4 & v84562f;
assign v230bb92 = hbusreq6 & v230429d | !hbusreq6 & v23f90b2;
assign v23f7ef3 = hgrant1_p & v23f580c | !hgrant1_p & v84561b;
assign v23fbcae = hmaster2_p & v23fb4e6 | !hmaster2_p & v230b621;
assign v230e97b = hgrant3_p & v22ffa6e | !hgrant3_p & !v84561b;
assign v23fce16 = hgrant4_p & v845635 | !hgrant4_p & b79a15;
assign v8c25df = hmaster2_p & v9d8aae | !hmaster2_p & v230e032;
assign v2306405 = hmaster2_p & v230446f | !hmaster2_p & v23fc530;
assign v22f2592 = hlock4_p & v23fc26a | !hlock4_p & !v22eeab9;
assign v22ef823 = hlock3_p & v22f8483 | !hlock3_p & v2303f04;
assign v22fc588 = hmaster1_p & v12cd9b5 | !hmaster1_p & v22f69ed;
assign v23fca72 = hgrant1_p & v23035ba | !hgrant1_p & v230065d;
assign a7fdb1 = hgrant3_p & v2311c16 | !hgrant3_p & v22ec0f7;
assign v22edf54 = locked_p & v230f974 | !locked_p & !v84561b;
assign v1aad609 = hbusreq3 & v22ed236 | !hbusreq3 & v84561b;
assign v230230d = hbusreq5 & v230bc8b | !hbusreq5 & v84561b;
assign v22fbaf1 = hmaster1_p & v22f1e81 | !hmaster1_p & !v230d5af;
assign v230aec0 = hlock0_p & v22eed66 | !hlock0_p & v22ffd22;
assign v22ecd3a = hbusreq4_p & v22f2b42 | !hbusreq4_p & !v84561b;
assign v230e95c = hbusreq4 & v23f5ad6 | !hbusreq4 & v230b2a4;
assign v23fb533 = hmaster0_p & v230741d | !hmaster0_p & v22f0a24;
assign v22ed494 = hbusreq3_p & v22fa9f7 | !hbusreq3_p & v84561b;
assign v23fb9a3 = hgrant3_p & v84561b | !hgrant3_p & v2393118;
assign v23fc14d = hbusreq5_p & v23fbbb0 | !hbusreq5_p & v23916fa;
assign v23f7275 = stateG10_5_p & v23f6309 | !stateG10_5_p & v22f878c;
assign v22f3e40 = hbusreq5 & v22f3a11 | !hbusreq5 & !v84561b;
assign v22ef3fe = hmaster1_p & v22eb748 | !hmaster1_p & v1aaddfe;
assign v22fe9dc = hbusreq3_p & v23f73dd | !hbusreq3_p & v23f9bcf;
assign v23f8a41 = hbusreq3_p & v230f9d5 | !hbusreq3_p & v84561b;
assign v23f8848 = jx2_p & v23fd002 | !jx2_p & v22f4cf2;
assign v2306609 = hbusreq5 & v23fbeb0 | !hbusreq5 & v23fca32;
assign v23fcc2f = hbusreq4_p & v23f2a25 | !hbusreq4_p & v22f98d3;
assign v23fbd58 = hmaster2_p & v22ef062 | !hmaster2_p & !v22ebfd7;
assign v22f167b = hgrant3_p & v22f19cb | !hgrant3_p & !v84561b;
assign v22faeec = stateG2_p & v84561b | !stateG2_p & v22f349a;
assign v23fcd76 = hbusreq0 & bd74c0 | !hbusreq0 & v23fa2ec;
assign v22ebaa4 = hbusreq3_p & v22ef0b4 | !hbusreq3_p & v22f9d19;
assign v22fd145 = hlock5_p & v22ede4d | !hlock5_p & v84561b;
assign v23f216d = hmaster0_p & v106ae19 | !hmaster0_p & v2309057;
assign v230f92a = hbusreq3 & v230e760 | !hbusreq3 & !v84561b;
assign v23fbb0c = hmaster0_p & v23fc755 | !hmaster0_p & v230463a;
assign v2308abb = hlock4_p & v23070dd | !hlock4_p & !v22eb265;
assign v22fd533 = hmaster2_p & v23fc6fe | !hmaster2_p & v23fa2ec;
assign v23929ca = hbusreq3_p & v22f324f | !hbusreq3_p & v22f25da;
assign v22fb3df = hbusreq5 & v22f337b | !hbusreq5 & v845620;
assign v2304a06 = hbusreq3_p & v23fc7c7 | !hbusreq3_p & v22eec47;
assign v23f5c89 = hlock3_p & v23fb1a1 | !hlock3_p & v22faae8;
assign v2304b2a = hmaster0_p & v23fc761 | !hmaster0_p & !v23fca1d;
assign v230b236 = hlock3_p & v23fbdb9 | !hlock3_p & !v84561b;
assign v23fb946 = hmaster0_p & v2312ec4 | !hmaster0_p & !v23fc44d;
assign f4061f = hbusreq6 & fc8fd5 | !hbusreq6 & v84561b;
assign v22ec782 = hbusreq1_p & v23fc530 | !hbusreq1_p & v230f5ee;
assign v22eaf73 = hmaster2_p & v22fc90f | !hmaster2_p & !v84561b;
assign v230af06 = hlock3_p & v22fd9f5 | !hlock3_p & v22f5218;
assign v23073e4 = hbusreq6_p & v23f333e | !hbusreq6_p & v2304928;
assign v23099b2 = jx1_p & v23fc4d8 | !jx1_p & v23f8294;
assign v23f292d = hbusreq3_p & v22ff83d | !hbusreq3_p & v23fce75;
assign v22f85c0 = hgrant3_p & v230ce52 | !hgrant3_p & v23f9081;
assign v230649c = hmaster1_p & v84561b | !hmaster1_p & bd94fd;
assign v22ed30e = jx1_p & v23fb202 | !jx1_p & v2309bcf;
assign v23f80c1 = hgrant1_p & v23fc9dd | !hgrant1_p & v23fcc8c;
assign v23fc1bc = hmaster2_p & v845627 | !hmaster2_p & !v23fcfa6;
assign v23fb960 = hbusreq5 & v23105cd | !hbusreq5 & v2312bd0;
assign v22f4810 = hmaster0_p & v22f4bae | !hmaster0_p & v230a4ef;
assign v22f7588 = hmaster0_p & v230d6fd | !hmaster0_p & v23f9033;
assign v23fbf80 = hbusreq0 & v84561b | !hbusreq0 & !v845629;
assign v23132fc = hgrant3_p & v22f2bb8 | !hgrant3_p & v23fc783;
assign v23f5f62 = jx2_p & v230aabf | !jx2_p & v23038cc;
assign v23f259c = hlock4_p & v23fc01f | !hlock4_p & !v23fcb6d;
assign v22f0677 = hbusreq2 & v22f36ff | !hbusreq2 & !v84561b;
assign v230cb1f = start_p & v84561b | !start_p & !v230a434;
assign v23f6f88 = hbusreq1_p & v2300c47 | !hbusreq1_p & v230075e;
assign v22fb051 = hbusreq5_p & v84561b | !hbusreq5_p & !v23078f5;
assign v22ee9bb = hbusreq3_p & v230200a | !hbusreq3_p & v23fce88;
assign v23fbdea = stateG10_5_p & v230ee7d | !stateG10_5_p & v845620;
assign v22feb95 = hgrant0_p & b5f51c | !hgrant0_p & v22fef36;
assign v22f9de9 = hgrant0_p & v23f4cdc | !hgrant0_p & v23ef9c4;
assign v23130c9 = hbusreq6 & v22f0fe5 | !hbusreq6 & v84561b;
assign v23fb8ae = stateG10_5_p & v2306b33 | !stateG10_5_p & !v84561b;
assign v22fdc2b = jx3_p & v84561b | !jx3_p & v23f89b6;
assign v230a5e6 = hbusreq1 & v231026b | !hbusreq1 & v84564d;
assign v23fbc61 = hmaster0_p & v2300985 | !hmaster0_p & !v23fc9bf;
assign v2302973 = hready & v230a117 | !hready & !v84561b;
assign v22f4ebc = hbusreq3_p & v191ac53 | !hbusreq3_p & v84561b;
assign v22ecea2 = jx3_p & v84561b | !jx3_p & v22f4950;
assign v2312060 = hbusreq3_p & v23efa39 | !hbusreq3_p & v106a782;
assign v23f54f3 = hmaster2_p & v22f7634 | !hmaster2_p & v22fec30;
assign v22ed898 = hbusreq2_p & v2309515 | !hbusreq2_p & !v22fa1af;
assign hgrant1 = !v1e841b6;
assign v23fbb98 = hgrant3_p & v23102b0 | !hgrant3_p & v23f2d1d;
assign v23fc30e = hbusreq5_p & v23f16fd | !hbusreq5_p & v23fcbe1;
assign v23fc1c4 = hlock4_p & v23fc7ca | !hlock4_p & v23fce25;
assign v22febe7 = hmaster2_p & v23fc514 | !hmaster2_p & v23fb9ad;
assign v22f6edc = hgrant3_p & v23fb6ed | !hgrant3_p & v231049c;
assign v22fb23d = hmaster2_p & v230fc56 | !hmaster2_p & v22fc564;
assign v23f024e = hgrant1_p & v23fbb7e | !hgrant1_p & v2303dcb;
assign v23fcdb2 = hbusreq1_p & v2306538 | !hbusreq1_p & bab0c9;
assign v22f2a94 = hgrant1_p & v23f79b4 | !hgrant1_p & v23f6d9c;
assign v23f6c41 = hgrant5_p & v22f8b0a | !hgrant5_p & v22fbc63;
assign v22f1b11 = hbusreq2 & v23f7efd | !hbusreq2 & v23fc228;
assign v22f79de = hburst1 & v22f3294 | !hburst1 & v9bd8c6;
assign v230f5a3 = locked_p & v23f6ac2 | !locked_p & !v84561b;
assign v23fc96b = hbusreq3 & v22f4301 | !hbusreq3 & v23fba9a;
assign v22f6277 = hbusreq3_p & v23fc1fc | !hbusreq3_p & v84561b;
assign v22fb42c = hmaster1_p & v12cda8f | !hmaster1_p & v23fbd21;
assign v2304b9d = hgrant0_p & v23133fa | !hgrant0_p & v84564d;
assign v23fb64a = hbusreq6_p & v23fc85b | !hbusreq6_p & v23fccaf;
assign d962e3 = hbusreq3 & b9ff2b | !hbusreq3 & v23fba9a;
assign v230a774 = hbusreq5_p & v9526ac | !hbusreq5_p & v22f8594;
assign v22f1892 = hmaster1_p & v23fb91a | !hmaster1_p & v1aad517;
assign v22f19a1 = hlock0 & v230d5ab | !hlock0 & v23fcf5c;
assign v2300dab = hmaster2_p & v22f343b | !hmaster2_p & v22ffea0;
assign v23f9887 = hbusreq6 & v2391d2f | !hbusreq6 & v23fcfd2;
assign c043dc = hmaster2_p & v84561b | !hmaster2_p & v230c70b;
assign v22f8e1b = hgrant3_p & v22fe392 | !hgrant3_p & v22fa05b;
assign v23f39e5 = hbusreq5 & v22f03cf | !hbusreq5 & !v845622;
assign v23094b2 = hbusreq3_p & v23fc19b | !hbusreq3_p & v23f7bc9;
assign v2306540 = hlock3_p & v23f733f | !hlock3_p & v230042c;
assign v2301f5d = hmaster0_p & v22f9403 | !hmaster0_p & v22f48ce;
assign v23fcf91 = hgrant0_p & v2306d29 | !hgrant0_p & v22fd30c;
assign v23fb436 = hbusreq3_p & v22f4d74 | !hbusreq3_p & v230a435;
assign v2300474 = hbusreq0_p & v191a876 | !hbusreq0_p & v191a879;
assign v23fcaf0 = hbusreq5_p & v23fa7ec | !hbusreq5_p & v84561b;
assign v23fb565 = hbusreq2_p & v84564d | !hbusreq2_p & v84561b;
assign v230812e = hready_p & v230f6d0 | !hready_p & v23fb4a9;
assign v23fc63e = hmastlock_p & v2302e47 | !hmastlock_p & v84561b;
assign v22ec53b = hbusreq0 & v230358b | !hbusreq0 & v22f8d74;
assign v22f3d4b = hmaster2_p & v1aae98c | !hmaster2_p & v84561b;
assign v230f133 = hbusreq3_p & v22f243b | !hbusreq3_p & v22f0e99;
assign v2306cae = hbusreq5_p & v230fec6 | !hbusreq5_p & v23fcd34;
assign v23130ea = hbusreq4 & v23fbb9b | !hbusreq4 & v84561b;
assign v23fcdde = hmaster2_p & v22ff120 | !hmaster2_p & v23fc03f;
assign v22fb272 = hgrant1_p & f406c6 | !hgrant1_p & !v22f94ea;
assign v23fb682 = hlock0_p & v23f55c0 | !hlock0_p & v23fb25c;
assign v22ff538 = hbusreq3 & v23112ad | !hbusreq3 & v22f61b6;
assign v22fe181 = hgrant3_p & v84562e | !hgrant3_p & v23fbd79;
assign v23fc931 = hmaster2_p & v23fc9f8 | !hmaster2_p & v22f8543;
assign v23fb5d0 = stateG10_5_p & v23f3115 | !stateG10_5_p & v845636;
assign v230d667 = hbusreq4 & v23fc67c | !hbusreq4 & v22ee657;
assign v23fbb7b = hbusreq4_p & v22fe08f | !hbusreq4_p & v22f3466;
assign v23f67dd = stateA1_p & v22f79de | !stateA1_p & v22f3294;
assign v23fcbd0 = hgrant3_p & v230c66e | !hgrant3_p & v23929ca;
assign v15072a7 = hbusreq6_p & v22eaeab | !hbusreq6_p & v23fb9e5;
assign v23fcc82 = hbusreq4_p & v230720b | !hbusreq4_p & v23102f3;
assign v22fbe9c = hmaster1_p & v84561b | !hmaster1_p & !v2313189;
assign v22eb5dd = hgrant5_p & v22f469a | !hgrant5_p & v22f2195;
assign v2392ff0 = hbusreq3_p & v230beb8 | !hbusreq3_p & v23fba11;
assign v23f763a = jx0_p & v23f9a36 | !jx0_p & v23fcb57;
assign v22f4aa2 = hbusreq5_p & v23f4b28 | !hbusreq5_p & v23035ba;
assign v23fc1f8 = hmaster0_p & v23fbea6 | !hmaster0_p & v23fb4b4;
assign v23fc3fd = hbusreq3 & v2305606 | !hbusreq3 & v22f6611;
assign v23fcd8e = hbusreq2_p & v23126ae | !hbusreq2_p & v191a876;
assign v23fbf93 = hbusreq1 & v22ee9be | !hbusreq1 & v2310a55;
assign v23fbb9b = hbusreq3_p & v23f8edc | !hbusreq3_p & v22eefd1;
assign v23fc234 = hbusreq4 & v23fb2ba | !hbusreq4 & v84564d;
assign v230b18b = hmaster1_p & v22f5d89 | !hmaster1_p & v22fa36d;
assign v22f8838 = hmaster2_p & v23f87f4 | !hmaster2_p & v23fcd14;
assign v23113f1 = jx1_p & v23fcab4 | !jx1_p & aacd54;
assign v23fb55a = stateG10_5_p & v22fbfe5 | !stateG10_5_p & v23f646e;
assign b9c92c = stateA1_p & v2302ca3 | !stateA1_p & v23f68bf;
assign v23fccb8 = jx1_p & v85e5cf | !jx1_p & v2311d16;
assign v230371b = start_p & v84561b | !start_p & v845663;
assign v230499e = hbusreq6_p & v230ec04 | !hbusreq6_p & v23fb242;
assign bd766b = hmaster2_p & v23f4855 | !hmaster2_p & v23f8928;
assign v22fa1ab = hmaster1_p & v230444c | !hmaster1_p & v84561b;
assign v22fff3a = hgrant4_p & v22fac3f | !hgrant4_p & v22fa616;
assign v23fc9e8 = hbusreq6_p & v23fbf41 | !hbusreq6_p & v23fc3e7;
assign v2301e25 = hbusreq2_p & v23f5043 | !hbusreq2_p & v84564d;
assign v22fbd4b = hgrant2_p & v2391545 | !hgrant2_p & !v84561b;
assign v2310826 = hbusreq1 & v22fd699 | !hbusreq1 & v84561b;
assign v23fcd14 = hbusreq5_p & v23fc1bb | !hbusreq5_p & v84561b;
assign v230972f = stateG10_5_p & v23fc4b2 | !stateG10_5_p & a1fba6;
assign v22f3b18 = hlock0_p & b9888a | !hlock0_p & v23effbc;
assign v23fba19 = hmaster0_p & v22ed756 | !hmaster0_p & v22f1dc9;
assign v23094c6 = stateG3_2_p & v84561b | !stateG3_2_p & v845663;
assign v22f8e10 = hgrant2_p & v13affe0 | !hgrant2_p & v23f79a9;
assign v2392ff9 = hmaster0_p & v23f2184 | !hmaster0_p & v2312608;
assign v23f7f51 = hlock4_p & v84561b | !hlock4_p & v230694d;
assign v23fbf0a = hmaster0_p & v23fc948 | !hmaster0_p & !v96c563;
assign v23fbc77 = hbusreq3_p & b9c9d4 | !hbusreq3_p & v84561b;
assign v22f9a85 = hbusreq1_p & v9a6a67 | !hbusreq1_p & !v22ffb91;
assign v1aada96 = hgrant3_p & v22f8cd9 | !hgrant3_p & v22f03a0;
assign v23fb6c6 = hgrant5_p & v22f5137 | !hgrant5_p & v23f08e5;
assign v23f40ba = hgrant0_p & v845622 | !hgrant0_p & v84562a;
assign bd7c6a = hmaster0_p & v23fbfbb | !hmaster0_p & v23fc76a;
assign v23fcf15 = hbusreq6_p & v230cf1d | !hbusreq6_p & v22ed645;
assign v23fc723 = hbusreq6 & v23fcd7f | !hbusreq6 & v22f475e;
assign v22ff244 = hbusreq6_p & v23fc110 | !hbusreq6_p & v2302c45;
assign v23fcf70 = hbusreq1_p & v2301655 | !hbusreq1_p & v23f5218;
assign v2391dfa = hgrant5_p & v230bdf9 | !hgrant5_p & v191a973;
assign ad6e26 = hmaster0_p & v22fd7d4 | !hmaster0_p & v22f2bf1;
assign v22f0393 = hmaster2_p & v23060d4 | !hmaster2_p & v230e8d3;
assign v2311cd1 = hbusreq3 & v2309d59 | !hbusreq3 & v23fc1c6;
assign v22f1962 = hgrant3_p & v84561b | !hgrant3_p & v22f9eb0;
assign v23f1703 = hbusreq3_p & v22ffd9a | !hbusreq3_p & v84561b;
assign v22fd0e6 = hgrant1_p & v84564d | !hgrant1_p & v22f8ad4;
assign v2311e39 = hbusreq3 & v22f881b | !hbusreq3 & v22f5834;
assign v23f7014 = hbusreq1 & v2311255 | !hbusreq1 & v84561b;
assign v23011a9 = hmaster2_p & v23101b1 | !hmaster2_p & v15070fa;
assign v22eed0b = hlock3_p & v230d7b4 | !hlock3_p & !v84561b;
assign v22eb02e = hmaster2_p & v23f646e | !hmaster2_p & v2306d29;
assign v230178e = hmaster0_p & v22f8aea | !hmaster0_p & v22f09ab;
assign v23fca4d = hbusreq6_p & v23fc169 | !hbusreq6_p & v22eb674;
assign v23f05e3 = hmaster0_p & v23fb9ec | !hmaster0_p & v23fc5d3;
assign v22f9bed = hgrant3_p & v239350a | !hgrant3_p & v22fffe4;
assign v2312d71 = hmaster0_p & v22fc6ca | !hmaster0_p & v22fd6c8;
assign v23f9773 = hbusreq5_p & v22fb71d | !hbusreq5_p & v22efeed;
assign v22f9b75 = hmaster2_p & v23fc71b | !hmaster2_p & !v23f940c;
assign v22fca2f = hlock0_p & v2303972 | !hlock0_p & v230834c;
assign v22f10d6 = hbusreq3_p & v23fceb9 | !hbusreq3_p & v22fd696;
assign v1aae387 = hmaster0_p & v22f8aea | !hmaster0_p & v22fcdf7;
assign v22fd696 = hbusreq1_p & v84562b | !hbusreq1_p & v23fb5b4;
assign v22f6986 = jx3_p & v22fbdb1 | !jx3_p & v22fb40c;
assign v22f8235 = hgrant1_p & v2305b35 | !hgrant1_p & !v23fbf9c;
assign v2302177 = hmaster2_p & v84561b | !hmaster2_p & v13afb18;
assign v2310b27 = hbusreq6 & v23021b9 | !hbusreq6 & !v230dc17;
assign v230baba = hbusreq5 & v13afe8f | !hbusreq5 & v84561b;
assign v23fcfdf = hbusreq5_p & v230383e | !hbusreq5_p & !v84561b;
assign v23fbb5b = hgrant3_p & v84561b | !hgrant3_p & v22f9d95;
assign v23fbe03 = hmaster1_p & v22fd6f9 | !hmaster1_p & v22f7371;
assign v22f7fed = hgrant3_p & v230b38b | !hgrant3_p & v23011a9;
assign v23fc3ff = hbusreq1_p & v2309ff9 | !hbusreq1_p & v84561b;
assign v23fb1f1 = hbusreq5 & v23fc51f | !hbusreq5 & v22fb71d;
assign v23029ed = hmaster2_p & v22f76ae | !hmaster2_p & v22f7ab4;
assign v22ed363 = hbusreq4_p & v22eed25 | !hbusreq4_p & v23f50d9;
assign v23fb094 = hmaster0_p & v22f81ba | !hmaster0_p & !v230abb0;
assign v23fc7f4 = hbusreq4_p & v22fca64 | !hbusreq4_p & v2312d03;
assign v23fbc55 = hbusreq2 & v23fc4a5 | !hbusreq2 & v23f391e;
assign v23fcf10 = hmaster1_p & v22f568c | !hmaster1_p & v22f78b4;
assign v22f8af0 = hlock3_p & a4e378 | !hlock3_p & v23fbc77;
assign v23f4fcd = hmaster2_p & v23f08a4 | !hmaster2_p & v84561b;
assign v2302ca7 = hbusreq3 & v22f8afa | !hbusreq3 & v22fab50;
assign v2308f7f = hmaster1_p & v84561b | !hmaster1_p & v23fccc6;
assign v230ccaf = hlock6_p & v23041ea | !hlock6_p & !v22f0bb6;
assign v22fbeb1 = hbusreq1_p & v84564d | !hbusreq1_p & v22f3643;
assign v22fc98d = hbusreq3_p & v23f35ea | !hbusreq3_p & v23f660f;
assign v22fb406 = jx1_p & v85e5cf | !jx1_p & v2305c74;
assign v2307b06 = hbusreq1_p & v22f40e3 | !hbusreq1_p & v84561b;
assign v23f5043 = hready & v84564d | !hready & v84561b;
assign v22ebe03 = hgrant1_p & v23fcbb6 | !hgrant1_p & v230580d;
assign v230c849 = hgrant3_p & v84561b | !hgrant3_p & v22ee5fb;
assign v23fb98e = hbusreq1_p & v22f03cf | !hbusreq1_p & v22fdf25;
assign v2302e1b = hmaster2_p & v2310e40 | !hmaster2_p & v230320e;
assign v23fc4f7 = hlock0_p & v230446f | !hlock0_p & v23f5c9b;
assign v845635 = hbusreq5_p & v84561b | !hbusreq5_p & !v84561b;
assign v23fbb63 = hmaster1_p & bd77c5 | !hmaster1_p & !v22f73a9;
assign v2346b79 = hmaster2_p & v84562b | !hmaster2_p & v22fc5fd;
assign v2310a58 = hmaster0_p & v23fc008 | !hmaster0_p & v22edc85;
assign v1aad45d = hmaster2_p & v23f052e | !hmaster2_p & v22fe920;
assign v23fbd99 = hbusreq2 & v22ef513 | !hbusreq2 & v84561b;
assign v23fb1db = hbusreq3_p & v23fcc58 | !hbusreq3_p & v23fc957;
assign v23fc491 = hmastlock_p & v22ee959 | !hmastlock_p & v84561b;
assign v22ec2ba = hmaster1_p & v23fbcd8 | !hmaster1_p & v22f9734;
assign v23f43db = hbusreq6_p & v230e800 | !hbusreq6_p & v22eea6a;
assign v23fc4e7 = hbusreq4 & a3aa64 | !hbusreq4 & v22f2ca2;
assign v2308818 = hbusreq1_p & v23fa2ec | !hbusreq1_p & v23fc4f8;
assign v2312ccb = hbusreq5_p & v23f8b6b | !hbusreq5_p & v23fbf6e;
assign v23fc796 = hgrant1_p & v845625 | !hgrant1_p & v22f5f09;
assign v23fcb96 = hmaster0_p & v22f5664 | !hmaster0_p & v22fffa6;
assign v22f65e3 = hgrant4_p & v84561b | !hgrant4_p & !v1aae9dc;
assign v22ef350 = hmaster2_p & v2309c52 | !hmaster2_p & !v84561b;
assign v230988d = hgrant3_p & v84561b | !hgrant3_p & v23f4e1c;
assign v22edbd4 = hmaster0_p & v98c729 | !hmaster0_p & v230f0de;
assign v22f6735 = hbusreq0_p & v23f4ae1 | !hbusreq0_p & v23fcdd5;
assign v230379f = hgrant3_p & v2307020 | !hgrant3_p & v2306d33;
assign v22f01b7 = jx3_p & v23047dd | !jx3_p & v2393705;
assign v2312bfb = hbusreq3_p & v23fb949 | !hbusreq3_p & v23f3f59;
assign v230c589 = stateG10_5_p & v23fa3a4 | !stateG10_5_p & v22fef02;
assign v23074cd = hbusreq4 & v23fbe82 | !hbusreq4 & v22ec339;
assign v23fc887 = hmaster0_p & v23fb084 | !hmaster0_p & !v96c563;
assign v23faee6 = hlock5_p & v23fb4d8 | !hlock5_p & !v84561b;
assign v231026b = hbusreq5_p & v1aae56f | !hbusreq5_p & v106ae21;
assign v23fce71 = hready & v23fb95d | !hready & !v2302c4b;
assign v22ed85a = hready & v84561b | !hready & v84564d;
assign v23fce2c = hgrant3_p & v84561b | !hgrant3_p & v23fbac0;
assign v23fbff3 = hmastlock_p & v84561b | !hmastlock_p & !v84565f;
assign v22f5039 = hbusreq1 & v22ee9be | !hbusreq1 & v23f3d14;
assign v22fec92 = hlock3_p & v23fc6a3 | !hlock3_p & v2312bfb;
assign v23fcdb4 = hbusreq1_p & v22ec334 | !hbusreq1_p & v84561b;
assign v2312a90 = hbusreq6 & v22f8012 | !hbusreq6 & v231261b;
assign v22fac3f = hmaster1_p & v84561b | !hmaster1_p & v23f0b74;
assign v22fd1ba = hbusreq4 & v23f1263 | !hbusreq4 & v22ebeb2;
assign v22fc4d3 = hlock2_p & v23fbfd0 | !hlock2_p & v2304494;
assign v2392adb = hbusreq0_p & v230f947 | !hbusreq0_p & !v22fd747;
assign v23021d9 = hmaster0_p & v230960c | !hmaster0_p & v230aa17;
assign v22ee6ce = hbusreq4_p & v845637 | !hbusreq4_p & bd8af4;
assign v22f4d68 = hgrant0_p & v845623 | !hgrant0_p & v23064ae;
assign v23fb4cd = hmaster2_p & v230d7b7 | !hmaster2_p & v84564d;
assign v23f9864 = hgrant3_p & v22f8838 | !hgrant3_p & v22feb6b;
assign v22f8f56 = hmaster2_p & v23065ad | !hmaster2_p & v23f11a3;
assign v23f1e4f = hbusreq3 & v23fbcd4 | !hbusreq3 & v84561b;
assign v23fb20f = hgrant3_p & v22f8e29 | !hgrant3_p & v230be8f;
assign v23fc50e = hmaster0_p & v2303fa0 | !hmaster0_p & v22fb88d;
assign v23fc2e8 = stateG10_5_p & v23f80e9 | !stateG10_5_p & v22fd767;
assign v1e84190 = hgrant3_p & v84561b | !hgrant3_p & bb324c;
assign v2311290 = hlock5_p & v23f820a | !hlock5_p & v23fb4ae;
assign v230764f = hbusreq4_p & v23fbfd8 | !hbusreq4_p & v22fd61b;
assign v22ee3a3 = hbusreq1 & v23f6b25 | !hbusreq1 & v84561b;
assign v22f62dc = hgrant5_p & v84561b | !hgrant5_p & v230d4b4;
assign v22f56d2 = hbusreq2_p & v2306d29 | !hbusreq2_p & v23126ae;
assign v22f8d80 = hbusreq0 & v22ed85a | !hbusreq0 & v84561b;
assign v2312839 = stateG10_5_p & v22f532c | !stateG10_5_p & !v22f8271;
assign v22fff2d = hmaster0_p & v22ee124 | !hmaster0_p & v22fa3fa;
assign b9c955 = hlock1_p & v845661 | !hlock1_p & !v84561b;
assign b535c6 = hmaster0_p & v2307fd0 | !hmaster0_p & !v2312c62;
assign v22fb8f1 = hbusreq1 & v22f860b | !hbusreq1 & !v845622;
assign v23fc873 = hbusreq3_p & v2306292 | !hbusreq3_p & v23fcb6c;
assign v23fb820 = hbusreq1_p & v22fbb07 | !hbusreq1_p & v22fd19c;
assign v2309320 = hmaster2_p & v239383d | !hmaster2_p & !v23fb98e;
assign v22f0d4e = hlock6_p & v84561b | !hlock6_p & v231131d;
assign v12cd3f4 = hbusreq2_p & v106ae19 | !hbusreq2_p & b9d013;
assign v22f2e92 = hmaster2_p & v2306932 | !hmaster2_p & !v22f1ae5;
assign v23043af = stateG10_5_p & v23fc732 | !stateG10_5_p & !v2303c9e;
assign v2311da1 = hbusreq4_p & v239174b | !hbusreq4_p & v191b1d9;
assign v22f69b7 = hlock0_p & v230f1a7 | !hlock0_p & v2307743;
assign v23fbedc = hbusreq1_p & v23fc8b3 | !hbusreq1_p & v84561b;
assign v2312de4 = hbusreq0_p & v23fbfb9 | !hbusreq0_p & !v23046f7;
assign v23f8f18 = hlock4_p & v23fbd13 | !hlock4_p & v230ba92;
assign v22eec68 = hbusreq6_p & v22f00eb | !hbusreq6_p & v2310fb9;
assign v22f2849 = hmaster2_p & v22ef403 | !hmaster2_p & v23fcda9;
assign v23f65f3 = hbusreq3_p & v23fba11 | !hbusreq3_p & v845620;
assign v22ffe8d = hgrant1_p & v845626 | !hgrant1_p & v230d8fa;
assign v23fb590 = hbusreq1 & v23f3ca5 | !hbusreq1 & v84561b;
assign v2303dcb = hgrant5_p & v23fc70c | !hgrant5_p & v23fc732;
assign v23f0dd1 = hgrant3_p & v22f7793 | !hgrant3_p & v22f89b9;
assign v23f1281 = hbusreq1 & v22f0073 | !hbusreq1 & !v23fc9db;
assign v23fc7e7 = hmaster2_p & v84561b | !hmaster2_p & v2307150;
assign v22fd06d = stateG10_5_p & v23f1ca8 | !stateG10_5_p & v230eb9b;
assign v22f69ed = hbusreq4_p & v23f669d | !hbusreq4_p & v23f33c7;
assign v22f591c = hmaster0_p & v231347a | !hmaster0_p & !v23fc91a;
assign v23f366d = hlock0_p & v2301655 | !hlock0_p & v23036ca;
assign v23919a5 = hbusreq2 & v1aae56f | !hbusreq2 & v84561b;
assign v1aad6a6 = hbusreq3_p & v23fba5a | !hbusreq3_p & v84561b;
assign v23f832b = hmaster2_p & v84561b | !hmaster2_p & v1e8471c;
assign v22fecf2 = hbusreq5_p & v22f5a2a | !hbusreq5_p & v2311fc9;
assign v2309a46 = hgrant3_p & v84561b | !hgrant3_p & v22f8440;
assign v22ef3d1 = hgrant3_p & v84561b | !hgrant3_p & v23ef4b1;
assign v22efa93 = hgrant1_p & v84561b | !hgrant1_p & v23030fc;
assign v23fc22e = hgrant1_p & v2307ee4 | !hgrant1_p & v23fc8bb;
assign v23fac5a = hlock0_p & e1de18 | !hlock0_p & !v84561b;
assign v22f18a3 = hmaster0_p & v2392d61 | !hmaster0_p & !v23fbfaa;
assign v23fb137 = hbusreq3_p & v23fb925 | !hbusreq3_p & v23f7688;
assign v23fcd6c = hmaster2_p & v23fc7ef | !hmaster2_p & v1aad38a;
assign v23f5596 = hgrant1_p & v22f3a35 | !hgrant1_p & v23fd057;
assign v22edc4f = hgrant1_p & v22fa999 | !hgrant1_p & !v230e598;
assign v23fbf07 = hlock3_p & v2307483 | !hlock3_p & v23fa21b;
assign v23fc22c = hmaster0_p & v22f674b | !hmaster0_p & v23fbaa2;
assign v22f446b = hmaster0_p & v23fc3e8 | !hmaster0_p & v22f7dbc;
assign v23fba9c = jx0_p & v22f1172 | !jx0_p & v23916d8;
assign v22f83fb = hmaster2_p & v23129e0 | !hmaster2_p & v23f8679;
assign v23fbd94 = stateG10_5_p & v23fc92a | !stateG10_5_p & v23f8ade;
assign v12ce9b8 = hbusreq5_p & v23fc0f3 | !hbusreq5_p & v22f4a7a;
assign v22f069f = hbusreq3 & v23fc273 | !hbusreq3 & v23f87f4;
assign v22fe495 = hbusreq1_p & v23fced9 | !hbusreq1_p & v84561b;
assign v23f4fbf = hmaster2_p & v23fc742 | !hmaster2_p & v23f4f1e;
assign v23f99cf = hbusreq1 & v23fc346 | !hbusreq1 & v84561b;
assign v22fc837 = hgrant6_p & v84561b | !hgrant6_p & v22ee3e8;
assign v2301c51 = hgrant3_p & v22f0546 | !hgrant3_p & v22f2c8b;
assign v23f36a3 = hbusreq4_p & v22f9b67 | !hbusreq4_p & v23122fa;
assign v23fc3c7 = hmaster1_p & v22f0104 | !hmaster1_p & v23fcdef;
assign v23fbfd8 = hmaster0_p & v22f14ff | !hmaster0_p & v22fe181;
assign v22fa851 = hbusreq3 & v230f578 | !hbusreq3 & v84561b;
assign v23fc282 = hlock3_p & v23fbcc8 | !hlock3_p & v22f8f1e;
assign v23f5d36 = hbusreq5_p & v22fdc30 | !hbusreq5_p & v23fb80e;
assign v22eb32b = hlock5_p & v84561b | !hlock5_p & v2300d1d;
assign v22f5d62 = hmaster1_p & v23fb482 | !hmaster1_p & v2312162;
assign v22f3e93 = hgrant5_p & v230d9d9 | !hgrant5_p & v22ff399;
assign v2301c57 = hbusreq3_p & v991952 | !hbusreq3_p & v23fca66;
assign v230521a = hbusreq4_p & v1aae387 | !hbusreq4_p & v22fc85f;
assign v23f68c1 = hbusreq1 & v23f5be9 | !hbusreq1 & v2391950;
assign e1bfb3 = hmaster2_p & v150745f | !hmaster2_p & v845636;
assign v23fbba6 = hbusreq4_p & v22ebd85 | !hbusreq4_p & v23fc2bc;
assign v23fc896 = hbusreq1_p & v191a86f | !hbusreq1_p & !v13afe8f;
assign v22f83e8 = hmaster2_p & v2311a1d | !hmaster2_p & v23fc35a;
assign v22f3a1f = hmaster1_p & v23f111f | !hmaster1_p & v22ed35b;
assign v22f7ab4 = hgrant1_p & v84561b | !hgrant1_p & v230dde9;
assign v23f004a = hmaster2_p & v23035d7 | !hmaster2_p & v1e8471c;
assign v230c749 = hbusreq3 & v23f7d43 | !hbusreq3 & v84561b;
assign v22f28c4 = hlock3_p & v23fbfd4 | !hlock3_p & v2302db0;
assign v2302b3f = hgrant5_p & v22f05f3 | !hgrant5_p & v2304b9d;
assign v2304583 = hmaster2_p & v22fa8e6 | !hmaster2_p & a5d081;
assign v23fc2df = hbusreq3_p & v23fc810 | !hbusreq3_p & v230e19d;
assign v22ffcae = hlock6_p & bd7ae5 | !hlock6_p & !v84561b;
assign v977ddf = jx1_p & v22f1aed | !jx1_p & v84561b;
assign v22f47fe = hbusreq5_p & v9526ac | !hbusreq5_p & v23fca1e;
assign v23f2843 = hlock3_p & v22fd9a5 | !hlock3_p & v22eea5b;
assign v22fb7e0 = hbusreq4 & v23fc48f | !hbusreq4 & v23fcc2e;
assign a1fbb6 = hmastlock_p & v23f54be | !hmastlock_p & v84561b;
assign v22f8b0a = hbusreq5_p & v22fef02 | !hbusreq5_p & v230c589;
assign v23934b5 = hbusreq6 & v23127ee | !hbusreq6 & v2303c5a;
assign v23fce7a = hmaster1_p & v22eb8e1 | !hmaster1_p & v84561b;
assign v23fc388 = hbusreq5_p & v22ff732 | !hbusreq5_p & v23fc054;
assign v2307c63 = hmaster0_p & v23f78a3 | !hmaster0_p & v22eee95;
assign v1e84174 = hgrant1_p & v84564d | !hgrant1_p & v230a3af;
assign v22f17bb = hlock0_p & v84561b | !hlock0_p & !v22ff8ea;
assign v23fc112 = hbusreq5 & v22ee0c4 | !hbusreq5 & !v84561b;
assign v230083b = hbusreq0_p & v2307b18 | !hbusreq0_p & v2309d29;
assign v23fcf05 = hbusreq0 & v22f1a26 | !hbusreq0 & v84561b;
assign v22fe551 = hlock3_p & v23fc610 | !hlock3_p & v106ae19;
assign v23fb948 = hbusreq6_p & v23f5a68 | !hbusreq6_p & v22fdad1;
assign v22ffad4 = hbusreq3_p & v22ef109 | !hbusreq3_p & v23fceb2;
assign v2392122 = hmaster0_p & v1aad34c | !hmaster0_p & v22ff70d;
assign v23fc2c1 = hgrant3_p & v84564d | !hgrant3_p & !v22f96f1;
assign v23f64db = hmaster2_p & v23f4f1e | !hmaster2_p & v230d3f5;
assign v23fcf52 = hmaster0_p & v230a9a3 | !hmaster0_p & !v23fa8c8;
assign v22edaa4 = hready & v22fc3b1 | !hready & !v84561b;
assign v23fcec4 = hlock4_p & v84561b | !hlock4_p & !v239157f;
assign v230feb2 = stateG10_5_p & v22efeed | !stateG10_5_p & !v845623;
assign v23f6309 = hgrant0_p & v22f878c | !hgrant0_p & v2310a9a;
assign v2301e40 = hmaster1_p & v230e0b7 | !hmaster1_p & v23fca4d;
assign fc8fdb = hlock3_p & v23f37c8 | !hlock3_p & v22f42a5;
assign v23f15a7 = hbusreq3_p & v84561b | !hbusreq3_p & !v230ae3f;
assign v23f8deb = hgrant5_p & v23fb489 | !hgrant5_p & v23fc4b2;
assign v2302e98 = hmaster0_p & b00aa6 | !hmaster0_p & v23fbcba;
assign v23fa8c7 = hbusreq3_p & v2310b0b | !hbusreq3_p & v22ee657;
assign v23070cf = hmaster2_p & v23fb90c | !hmaster2_p & v230b1ac;
assign v23fb635 = hmaster0_p & bd7ae5 | !hmaster0_p & v12cd5f2;
assign v23fc3b8 = hlock4_p & v9bcd2e | !hlock4_p & !v8fb6b6;
assign v230c428 = hgrant0_p & v22f516b | !hgrant0_p & v23fab8b;
assign v23fba0b = hbusreq1 & v23f301a | !hbusreq1 & v22ed493;
assign v23f5c95 = hlock0_p & v84561b | !hlock0_p & v23f835c;
assign v22f84ff = hgrant0_p & v845622 | !hgrant0_p & v23f6765;
assign v191afef = hgrant3_p & v8ea3a5 | !hgrant3_p & v2311b78;
assign v230f755 = hgrant5_p & v84561b | !hgrant5_p & !v2312441;
assign v23fc9d6 = hmaster0_p & v23f58bb | !hmaster0_p & v230f7ce;
assign v2302c08 = hbusreq2 & v22f7e16 | !hbusreq2 & v84561b;
assign v22f19cc = hlock5_p & v2304f32 | !hlock5_p & bbc337;
assign v2311656 = hbusreq3_p & v2305b58 | !hbusreq3_p & v84561b;
assign v22ece03 = hbusreq5 & v191ae42 | !hbusreq5 & !v84561b;
assign v23f3f38 = hlock4_p & v23fc1f8 | !hlock4_p & !v230a092;
assign v2307ab1 = stateG10_5_p & v23f6380 | !stateG10_5_p & !v22f5243;
assign v23015a7 = hbusreq1 & v22feb47 | !hbusreq1 & v84561b;
assign v2391f2b = hgrant1_p & v23f0625 | !hgrant1_p & v22f78de;
assign v23f3051 = hgrant5_p & v22eec5f | !hgrant5_p & !v22f217d;
assign v23fbd8c = hready_p & v22f35eb | !hready_p & !v22eec2d;
assign v22f78a9 = hbusreq5 & v8d360e | !hbusreq5 & !v84561b;
assign v23fbfee = hbusreq3_p & v23f2704 | !hbusreq3_p & v23f200c;
assign v230184a = hlock4_p & v23f965d | !hlock4_p & !v84561b;
assign v23fb501 = hbusreq5_p & v23f7148 | !hbusreq5_p & v22f8b9c;
assign v23132e5 = hmaster1_p & v22fefde | !hmaster1_p & v2305b24;
assign v21b35f9 = hmastlock_p & v23fb476 | !hmastlock_p & v84561b;
assign v22f6176 = hbusreq4_p & v23fb99f | !hbusreq4_p & v23fbe63;
assign v2304abd = hbusreq6 & b00aa0 | !hbusreq6 & v845625;
assign v2306414 = hlock5_p & v22f99ee | !hlock5_p & v23014fb;
assign v23018f2 = hmaster2_p & v22f542d | !hmaster2_p & v84561b;
assign v230d709 = hgrant1_p & v23fce81 | !hgrant1_p & v22fb450;
assign v23fc4c2 = hbusreq6 & v2305a2a | !hbusreq6 & v84561b;
assign v22f5808 = hmaster0_p & v23fb8aa | !hmaster0_p & v22f46ff;
assign v2300d51 = hgrant2_p & v23f646e | !hgrant2_p & !v22ec29a;
assign v22eaeaf = hbusreq4 & v845620 | !hbusreq4 & v84561b;
assign v22ef61b = hmaster0_p & v22f2e69 | !hmaster0_p & v2303efe;
assign v23f1974 = hbusreq0_p & v2305a12 | !hbusreq0_p & !v22ec921;
assign v230037d = hbusreq0_p & v230a63b | !hbusreq0_p & v84561b;
assign v2391e51 = hbusreq5 & v22ff315 | !hbusreq5 & v84561b;
assign v22f6de3 = hgrant5_p & v22ef458 | !hgrant5_p & v230cf1a;
assign v22f0567 = hbusreq3_p & v1506f9f | !hbusreq3_p & v23f20d3;
assign v23fc64c = hmaster2_p & v2306b2e | !hmaster2_p & v84561b;
assign v239308e = hbusreq3_p & v23fb479 | !hbusreq3_p & v23087e9;
assign v22f65b0 = hmaster2_p & a07f9b | !hmaster2_p & v23f1a8d;
assign v23077e6 = hbusreq5_p & v23fb928 | !hbusreq5_p & !v84561b;
assign v23045dc = hbusreq3_p & v22ecb12 | !hbusreq3_p & v22f4ef7;
assign v12cc321 = decide_p & v2392ec8 | !decide_p & v23fb76c;
assign v23fc7bb = hmaster0_p & v23f3915 | !hmaster0_p & v23fc65d;
assign v23022c3 = hmaster2_p & b00ad3 | !hmaster2_p & v84561b;
assign v22f1969 = hbusreq6_p & v23fb5b9 | !hbusreq6_p & v23f664b;
assign v22fc2d0 = hmaster0_p & v230741d | !hmaster0_p & v2302e1b;
assign v1507529 = hgrant1_p & v845625 | !hgrant1_p & v23919bb;
assign v23f2041 = hbusreq6_p & v22f7ccb | !hbusreq6_p & v23f7b9e;
assign v230753a = hbusreq3_p & v22f6870 | !hbusreq3_p & v23fca08;
assign v2300059 = hbusreq5_p & v22f679f | !hbusreq5_p & v22fb71d;
assign stateG10_5 = !d49f4d;
assign v22f0d22 = hbusreq5 & v23fb978 | !hbusreq5 & v84561b;
assign v22ee195 = hgrant0_p & v2310904 | !hgrant0_p & v23f8747;
assign v22ff123 = hbusreq2 & v23fc07d | !hbusreq2 & !v845620;
assign v22f7b3e = hbusreq3_p & v1aad8a4 | !hbusreq3_p & !v84561b;
assign v22f6aa3 = hgrant3_p & v22f8e29 | !hgrant3_p & v22ed2f5;
assign v23fc844 = hbusreq4_p & v22f7152 | !hbusreq4_p & v84561b;
assign v23fc7d4 = jx0_p & v23f66cf | !jx0_p & v22f2a85;
assign v22fab21 = hmaster2_p & v23f8490 | !hmaster2_p & !v23fcda9;
assign v2303cae = jx1_p & v85e5cf | !jx1_p & !v23fbfb1;
assign v2312336 = hgrant0_p & v23fc4f8 | !hgrant0_p & v22f2879;
assign v23fb85a = hlock3_p & v23fce54 | !hlock3_p & !v84561b;
assign v231164b = hbusreq5_p & v230094d | !hbusreq5_p & v22fe948;
assign v23fbb9d = hbusreq3 & v23f883c | !hbusreq3 & v84561b;
assign v23019f7 = hbusreq3_p & v23fc20d | !hbusreq3_p & !v23fc92f;
assign v23fb1bb = hbusreq4 & v23fc7c0 | !hbusreq4 & v84562f;
assign v23fba12 = hmaster2_p & v191a876 | !hmaster2_p & !v23f3a16;
assign fc8f74 = hlock2_p & v22f9a51 | !hlock2_p & v84561b;
assign v23fc3a7 = hbusreq0_p & v22fd30c | !hbusreq0_p & v23f512e;
assign v23f6e64 = hgrant0_p & v845622 | !hgrant0_p & v239171e;
assign v22ed614 = hgrant5_p & v22fe6b3 | !hgrant5_p & !v2306b33;
assign v22f99e0 = hmaster2_p & v22f1389 | !hmaster2_p & v23f3ca5;
assign v2311944 = hbusreq6_p & v22eeb4b | !hbusreq6_p & v2312325;
assign v23fbf55 = hmaster2_p & v84561b | !hmaster2_p & v2312ea7;
assign v23fcff0 = hbusreq2 & v2313118 | !hbusreq2 & v23fc228;
assign v2307707 = hbusreq0 & v22f36ff | !hbusreq0 & !v84561b;
assign v23f58e5 = hbusreq1_p & v23f40ab | !hbusreq1_p & v84561b;
assign v23fbd42 = hbusreq5 & v23fbb8b | !hbusreq5 & v84561b;
assign v22f482d = hmaster0_p & v23fbdf6 | !hmaster0_p & !v23fc20d;
assign v22f4bae = hbusreq3_p & v23fc4a8 | !hbusreq3_p & v2300a04;
assign v23041b6 = hbusreq5_p & v23fbe4c | !hbusreq5_p & v22f94ba;
assign v919672 = hmaster2_p & v23fb6ce | !hmaster2_p & v23fc461;
assign v22fd3b1 = stateG10_5_p & a1bfd6 | !stateG10_5_p & v84561b;
assign v2302e0f = hmaster0_p & v22f56a5 | !hmaster0_p & !v23fcd24;
assign v22fd8c5 = hbusreq3 & v22fe675 | !hbusreq3 & v84561b;
assign v22f92f8 = hgrant5_p & v23f4979 | !hgrant5_p & v22ece0d;
assign v2393f3f = hbusreq6_p & v23fca4a | !hbusreq6_p & v22eb12e;
assign v23f4722 = hlock0_p & v13aff3b | !hlock0_p & v22f5b73;
assign v230f613 = hlock6_p & a1fe5e | !hlock6_p & e1deb1;
assign v2309248 = hmaster0_p & v9d1fa2 | !hmaster0_p & !v96c563;
assign v23fb31d = hbusreq4 & v22faa7c | !hbusreq4 & v23fce05;
assign v23fc908 = hbusreq6 & v2308a91 | !hbusreq6 & v230c437;
assign v22f051d = hbusreq5 & v22f3a11 | !hbusreq5 & v23f40ba;
assign v22ede0b = hbusreq4 & v2305cc1 | !hbusreq4 & v84561b;
assign v22fd713 = hbusreq5 & v23fba6b | !hbusreq5 & !v84561b;
assign v9347cd = hgrant5_p & v22f05f3 | !hgrant5_p & v2306257;
assign v22f9552 = hbusreq6 & v22f5767 | !hbusreq6 & v22eed0b;
assign v2302bd3 = hbusreq5_p & v23f5ce0 | !hbusreq5_p & !v84561b;
assign v22efcad = hmaster0_p & v23fbf3e | !hmaster0_p & v22fc37d;
assign v2309fdb = hlock1_p & v23fbd41 | !hlock1_p & !v2304ec7;
assign v22f1fec = hbusreq0 & v22f5037 | !hbusreq0 & v22f9927;
assign v1aad65a = hbusreq6 & v23fb978 | !hbusreq6 & v84561b;
assign v2309c28 = hlock0_p & v2301511 | !hlock0_p & v9e764b;
assign v2303393 = hlock0_p & v23fba13 | !hlock0_p & v2306885;
assign v23fcb3c = hmaster2_p & v2304fae | !hmaster2_p & v23f8928;
assign v22f4af5 = hbusreq6_p & v22f248e | !hbusreq6_p & v22f0acc;
assign v22ef0ab = hmaster2_p & v22eec6e | !hmaster2_p & v22fd0e6;
assign v231324d = hbusreq4_p & v23fc613 | !hbusreq4_p & v23fcd97;
assign v23f4ed3 = hmaster2_p & v2311a1d | !hmaster2_p & v23f3cb8;
assign v22efdae = hbusreq3_p & v2305d6e | !hbusreq3_p & v2300ccc;
assign v23fc983 = hmaster2_p & v84561b | !hmaster2_p & !v230913d;
assign v22f1ae7 = hgrant1_p & v23065ad | !hgrant1_p & v2393417;
assign v1506ae6 = hgrant5_p & v23fcf79 | !hgrant5_p & v22ee457;
assign v191aea6 = hbusreq2_p & v22fd79e | !hbusreq2_p & d49f20;
assign v23037b3 = hmaster0_p & v23f9d9a | !hmaster0_p & !v23f864d;
assign v22f609f = hbusreq3_p & v22fb28f | !hbusreq3_p & v22fe831;
assign v230c124 = hbusreq5_p & v23fb873 | !hbusreq5_p & v230d793;
assign v230db01 = hgrant0_p & v23fc5f4 | !hgrant0_p & v84561b;
assign v230f8b2 = hready & v22f8278 | !hready & v23011cb;
assign v22f7d04 = hmaster0_p & v230a9a3 | !hmaster0_p & v23fb0d0;
assign v230e1a3 = hbusreq1_p & v2305838 | !hbusreq1_p & v23fb6a6;
assign v1aae2e4 = hmaster1_p & v239158d | !hmaster1_p & bc87ee;
assign v23fcf1f = hbusreq5 & v84561b | !hbusreq5 & v845620;
assign v22fa5a0 = hbusreq3_p & v2308b33 | !hbusreq3_p & v2302d69;
assign v22fa6a4 = hmaster2_p & v23fc40f | !hmaster2_p & v23fcaf0;
assign v23fc250 = hbusreq2 & v22ee145 | !hbusreq2 & v84561b;
assign v22eb334 = hbusreq2 & v12cd8c9 | !hbusreq2 & v84561b;
assign v23fbe1c = hmaster2_p & v230e8d3 | !hmaster2_p & v22f893a;
assign v23f1279 = hbusreq3_p & v23fbc40 | !hbusreq3_p & v23fc2d7;
assign v22fa16b = hbusreq5_p & v84561b | !hbusreq5_p & v23fc706;
assign v230788d = hbusreq3_p & v23f7a18 | !hbusreq3_p & v86df86;
assign v23fcb69 = locked_p & v230e58e | !locked_p & a1fbb6;
assign v2302d53 = hbusreq6_p & v191afb7 | !hbusreq6_p & v23fc128;
assign v23f723b = hmaster0_p & v23f3d38 | !hmaster0_p & v230ad95;
assign v22fbbb8 = hbusreq5_p & v22f5037 | !hbusreq5_p & v22f931d;
assign v2302071 = hbusreq5_p & v22f343b | !hbusreq5_p & v9585ce;
assign v23fc513 = hbusreq0 & v22f446e | !hbusreq0 & v84561b;
assign v230d134 = hbusreq3 & v23f5fa6 | !hbusreq3 & v84561b;
assign v22ed7a4 = hmaster0_p & v2312189 | !hmaster0_p & v230f2af;
assign v22f8bd7 = hbusreq6_p & v963cc3 | !hbusreq6_p & v23139b9;
assign v23fb968 = stateG10_5_p & v23fb4bd | !stateG10_5_p & !v22f8e5d;
assign v23083ee = hmaster0_p & v23fcab1 | !hmaster0_p & !v23129e8;
assign v23f6836 = hlock0_p & v1aae56f | !hlock0_p & v2308bbe;
assign v22f6169 = hgrant3_p & v22f368e | !hgrant3_p & v2303a74;
assign v22ef3f8 = jx3_p & v230f1d9 | !jx3_p & v23fb6a0;
assign v23fc484 = hbusreq1_p & v2308d09 | !hbusreq1_p & !v22f9980;
assign v2303d95 = hbusreq1_p & v23fcf71 | !hbusreq1_p & v23fb7e0;
assign v2307553 = hmaster2_p & af6dff | !hmaster2_p & v230e3a0;
assign v23fc91c = hbusreq6 & v23125ee | !hbusreq6 & !v22f9183;
assign v23094cb = hbusreq0 & v13afe3a | !hbusreq0 & !b00ad3;
assign v22f946f = stateG10_5_p & v22fcc0d | !stateG10_5_p & v98d297;
assign v2312f7e = hmastlock_p & a1fd35 | !hmastlock_p & v84565f;
assign v230dc73 = hmaster2_p & v23fbf32 | !hmaster2_p & !v22f5b4b;
assign v22f0de9 = hgrant5_p & v23fc578 | !hgrant5_p & v230d1a6;
assign v22f469a = hbusreq5_p & v22ff732 | !hbusreq5_p & v22f7dd1;
assign v23fc228 = hlock2_p & v23f1879 | !hlock2_p & v845620;
assign v23fcf77 = hbusreq5_p & v230e167 | !hbusreq5_p & !v84561b;
assign v23fc44a = hbusreq4_p & v231232b | !hbusreq4_p & v84561b;
assign v22fe0b0 = hmaster2_p & a1fba6 | !hmaster2_p & v230945e;
assign v23fcdf0 = hbusreq4 & v23fc4b0 | !hbusreq4 & v22ed01d;
assign v22f118e = hbusreq3_p & v2303f7c | !hbusreq3_p & !bd7a62;
assign v2311e9f = hbusreq4_p & v2300cc2 | !hbusreq4_p & v22fc767;
assign v23122cb = hbusreq3_p & v230e37a | !hbusreq3_p & v15070ca;
assign v230a0e7 = hbusreq4_p & v2310538 | !hbusreq4_p & v23fcd5c;
assign v2306291 = hbusreq6_p & v230f613 | !hbusreq6_p & v23fb0c7;
assign v230262f = stateG10_5_p & v22f7f74 | !stateG10_5_p & v22ffc69;
assign v23fbe4b = hbusreq4_p & v22f4bc7 | !hbusreq4_p & v23fc3cd;
assign v23fcc5a = hbusreq0_p & v84564d | !hbusreq0_p & v22f3643;
assign e1dd71 = hbusreq1_p & v2300071 | !hbusreq1_p & v23f15ac;
assign v23007f2 = hbusreq2 & v2310ad7 | !hbusreq2 & !v22f70f4;
assign v230dd9e = hgrant5_p & v22f5d15 | !hgrant5_p & !v997ca9;
assign v87c96d = hbusreq3_p & v23106e3 | !hbusreq3_p & v23011a9;
assign v1aae6ba = jx1_p & v231185e | !jx1_p & v230e991;
assign v23015be = hbusreq1 & v22fc091 | !hbusreq1 & v22f5583;
assign v23f5a88 = hlock2_p & v84561b | !hlock2_p & !fc8ab7;
assign v230e94c = hbusreq4_p & v22ee43f | !hbusreq4_p & v23f1bd6;
assign v22f5b27 = hbusreq5_p & v22f051d | !hbusreq5_p & v22f442c;
assign v23f50bb = hbusreq1_p & v23fbe09 | !hbusreq1_p & v1506ae6;
assign v23013d7 = hmaster1_p & v22efcc1 | !hmaster1_p & v23fb384;
assign v22ecc15 = hbusreq2_p & v23fc151 | !hbusreq2_p & !v191a876;
assign v23f86dc = hmaster2_p & v2308d51 | !hmaster2_p & v84561b;
assign v23f87f4 = hbusreq5_p & bbc337 | !hbusreq5_p & v84561b;
assign v23fc855 = jx1_p & v23056b2 | !jx1_p & v23fc523;
assign v231228f = hmaster1_p & v23fc7f2 | !hmaster1_p & v23fcd9b;
assign v2309543 = hgrant6_p & v845629 | !hgrant6_p & v22f166b;
assign v23f6fe8 = hmaster0_p & v22fbde3 | !hmaster0_p & v22f9056;
assign baa026 = hbusreq3_p & v22f695c | !hbusreq3_p & v106a782;
assign v23133fa = hlock0_p & v84564d | !hlock0_p & !v84561b;
assign v23fc0fd = stateG2_p & v84561b | !stateG2_p & v2308f85;
assign v230bbe4 = stateG10_5_p & v23fc7f5 | !stateG10_5_p & v22f878c;
assign v22f70bf = hmaster1_p & v23f5388 | !hmaster1_p & v23fbba0;
assign v230128e = hbusreq4_p & v12cd538 | !hbusreq4_p & v22fef6a;
assign v23fc8c3 = hlock0_p & v23fd040 | !hlock0_p & v22fd794;
assign v23fbaae = hbusreq0 & v22ebbea | !hbusreq0 & !v84561b;
assign afc788 = hbusreq0 & v84561b | !hbusreq0 & v845620;
assign v22fe2ae = hmaster2_p & v84561b | !hmaster2_p & v845620;
assign v22f9fe0 = hbusreq1_p & v230fcad | !hbusreq1_p & v22f7241;
assign v23f5a8b = hgrant5_p & v22fff04 | !hgrant5_p & v22ed2f0;
assign c17811 = hmaster1_p & v2305853 | !hmaster1_p & v2311944;
assign v23129d7 = hmaster1_p & v22fc9cd | !hmaster1_p & v22fc477;
assign v22ffe51 = hbusreq1 & v2312f7e | !hbusreq1 & !v231009b;
assign v22f4f1e = hgrant0_p & v2305fe0 | !hgrant0_p & !v84561b;
assign v230c3ee = hmaster0_p & v23fcdb0 | !hmaster0_p & !v23fb58e;
assign v22f7997 = hmaster0_p & a25b7d | !hmaster0_p & v23fc5fb;
assign v22eaee1 = hmaster2_p & v23f5af5 | !hmaster2_p & v22f8271;
assign v22f0073 = hbusreq2_p & v2301aa7 | !hbusreq2_p & v84561b;
assign v22f96f2 = hgrant0_p & v84561b | !hgrant0_p & v22fcd0c;
assign v230b50c = hgrant1_p & v230e336 | !hgrant1_p & v230faa5;
assign v23f1515 = hbusreq5 & v23f0169 | !hbusreq5 & v2304536;
assign v23fb495 = hlock6_p & v23086ec | !hlock6_p & v22f5215;
assign v23f08d9 = hbusreq5 & v2303125 | !hbusreq5 & v230fa13;
assign v231343f = hgrant5_p & v23fc74f | !hgrant5_p & v23fcccf;
assign v22fbdd6 = hmaster2_p & v23fca2a | !hmaster2_p & v22f0824;
assign v22f1afb = hbusreq6_p & v2391fc6 | !hbusreq6_p & v23f397b;
assign v23f3970 = hmaster0_p & v23fa3b8 | !hmaster0_p & v23fc478;
assign v22f251d = hbusreq4_p & v23fc640 | !hbusreq4_p & !v230a0ad;
assign v23fc235 = hlock3_p & v22f609f | !hlock3_p & v22fe831;
assign v22f7d9a = hmaster2_p & v84561b | !hmaster2_p & v2304781;
assign v2300142 = hlock3_p & v23fb1db | !hlock3_p & v23f3d0b;
assign v23fb0bf = hlock4_p & v22f297d | !hlock4_p & v22eaeaf;
assign v23fb0dd = hbusreq5_p & v23fc4a1 | !hbusreq5_p & v2305926;
assign v22f679f = hbusreq5 & v2306b33 | !hbusreq5 & v22fb71d;
assign v23fcdc4 = stateA1_p & v23fc8d7 | !stateA1_p & !v230493b;
assign v230e5da = hgrant3_p & v84561b | !hgrant3_p & v22ebaa4;
assign v231089e = hbusreq6 & v2310641 | !hbusreq6 & v22ecbc3;
assign v22f0c5d = stateG2_p & v84561b | !stateG2_p & v23fcdaa;
assign v22fca61 = locked_p & v23109e9 | !locked_p & !v84561b;
assign v23fbcbe = hlock4_p & v22eb58b | !hlock4_p & !v23fc7dc;
assign a1ff27 = stateA1_p & v22f178d | !stateA1_p & !v84561b;
assign v23fc23b = hmaster2_p & v84561b | !hmaster2_p & !v22f037a;
assign v23fbd26 = hlock5_p & b8cd18 | !hlock5_p & v22fe95c;
assign v22f4321 = hmaster0_p & v23130ea | !hmaster0_p & v22fd7ee;
assign v23fb0b6 = hbusreq3_p & v230b740 | !hbusreq3_p & v23fb84b;
assign v23fc8d6 = hgrant3_p & v22f368e | !hgrant3_p & v23fb8d6;
assign v2302131 = hmaster2_p & v84561b | !hmaster2_p & v84564d;
assign v230f860 = stateG10_5_p & v22f7004 | !stateG10_5_p & v23fc4f8;
assign v22f5495 = hmaster2_p & v23fbaaa | !hmaster2_p & be9b63;
assign v22fb335 = hgrant3_p & v84561b | !hgrant3_p & v23f5d23;
assign v23fbce3 = hbusreq3 & v84561b | !hbusreq3 & v23fba11;
assign v191b18a = hbusreq1_p & v23126ae | !hbusreq1_p & v191a876;
assign v22fdf25 = hbusreq5_p & v22f03cf | !hbusreq5_p & v23fcb14;
assign v23f756e = hbusreq6 & v23fca1c | !hbusreq6 & v84561b;
assign v2300774 = hmaster2_p & v22f1796 | !hmaster2_p & v23f8ca4;
assign v230e58e = hmastlock_p & v23fc219 | !hmastlock_p & v84561b;
assign v22f8427 = hgrant1_p & v84564d | !hgrant1_p & !v23fc6ca;
assign v22fb1d7 = hbusreq4 & v23fc627 | !hbusreq4 & v84562d;
assign v23fbbaa = hlock4_p & v23fbbef | !hlock4_p & !v84561b;
assign v22f658e = hmaster0_p & b031da | !hmaster0_p & !v84561b;
assign v22ec855 = hbusreq3_p & v23fc19b | !hbusreq3_p & v23fc0ac;
assign v23f8cd3 = hgrant5_p & v23fb217 | !hgrant5_p & v23fb84f;
assign v23fb1aa = hbusreq5_p & v84561b | !hbusreq5_p & v23064ae;
assign v94f831 = hbusreq6_p & v23f1f36 | !hbusreq6_p & v23f7714;
assign v23fbc4a = stateG10_5_p & v106af57 | !stateG10_5_p & v23f5af5;
assign v22fa9f7 = hbusreq3 & v2303fb2 | !hbusreq3 & v84561b;
assign v23f3e7f = hbusreq2_p & a1fee6 | !hbusreq2_p & !v23f680a;
assign v23115f8 = hmaster0_p & v230b111 | !hmaster0_p & v23fb586;
assign v23fc1fc = hbusreq3 & v23f3dcc | !hbusreq3 & v84561b;
assign a9c602 = hmaster2_p & v191aa68 | !hmaster2_p & v23f3a16;
assign v22f859d = hmaster2_p & v2301585 | !hmaster2_p & v22f53c0;
assign v23fba93 = hbusreq1_p & v1506fbf | !hbusreq1_p & v2310eb6;
assign v23fce8d = hbusreq2 & v23fb9b9 | !hbusreq2 & v84561b;
assign v230174f = hlock4_p & v22f91a6 | !hlock4_p & v23f4937;
assign v23f3b1e = hgrant1_p & v22f0139 | !hgrant1_p & v22f5a08;
assign v22fd50f = hgrant5_p & v2305f5e | !hgrant5_p & v23fc1c8;
assign v22f2d05 = stateG2_p & v84561b | !stateG2_p & !v230efb1;
assign v230f9db = hbusreq1_p & v84561b | !hbusreq1_p & v23fb1aa;
assign v23920aa = hlock3_p & v2311656 | !hlock3_p & v23fc260;
assign v22fee46 = locked_p & v106ae1c | !locked_p & a1fbb6;
assign v22ec5d6 = hmaster0_p & v23fac2d | !hmaster0_p & !v23fcbe2;
assign v23fc42c = hbusreq4_p & v84561b | !hbusreq4_p & v23fc75d;
assign v23f4fe1 = hbusreq3_p & v23fcd66 | !hbusreq3_p & v230697e;
assign v23fcb58 = hbusreq0 & v23f2a3d | !hbusreq0 & v84564d;
assign v230a510 = hgrant3_p & v23f651a | !hgrant3_p & !v23fd008;
assign v230c94b = hbusreq4_p & v23f7cec | !hbusreq4_p & v22fc2d0;
assign v23fc256 = hmaster2_p & v22f83cf | !hmaster2_p & v22f11fe;
assign v22ebbab = hlock3_p & v84561b | !hlock3_p & !v22ec8d7;
assign v23096e7 = hmaster0_p & v22f7800 | !hmaster0_p & v23f7b32;
assign v22eeb07 = hlock5_p & v23fb710 | !hlock5_p & !v845636;
assign v1aad8a8 = hbusreq3_p & v23fa511 | !hbusreq3_p & v22fc37d;
assign v22fe775 = hbusreq3_p & v2311c98 | !hbusreq3_p & v23fba9a;
assign v22f8cb9 = hgrant3_p & v84561b | !hgrant3_p & !v22fe920;
assign v23f9885 = hgrant3_p & v230a744 | !hgrant3_p & v23fcfb6;
assign v1507161 = hbusreq0_p & v22f8d80 | !hbusreq0_p & v84561b;
assign v23fc5ec = hbusreq2 & v22ed6c5 | !hbusreq2 & v84564d;
assign v22f3e5b = hbusreq4_p & v23f3073 | !hbusreq4_p & v23fb70f;
assign v23f9414 = hbusreq1_p & v23fa6f1 | !hbusreq1_p & v845620;
assign v23f3de0 = hbusreq4 & v22edf31 | !hbusreq4 & v84561b;
assign v23fab18 = hbusreq1_p & v23f6250 | !hbusreq1_p & v84561b;
assign v23f6ac5 = hbusreq1 & v2302e32 | !hbusreq1 & !v84561b;
assign v2303245 = hbusreq5_p & v2305fe0 | !hbusreq5_p & !v23fc2ea;
assign v230d8fa = hgrant5_p & v23fc9c4 | !hgrant5_p & v230eb8d;
assign v2302075 = hgrant0_p & a84b89 | !hgrant0_p & v23fc55f;
assign v22f5605 = hlock0_p & v23f5cb3 | !hlock0_p & v2311ec3;
assign v23f67fa = hmaster0_p & v22f2abb | !hmaster0_p & !v230a709;
assign v22fb88e = stateG10_5_p & v23052cc | !stateG10_5_p & v2301e25;
assign v2307c5d = hgrant1_p & v23f908f | !hgrant1_p & v230ee35;
assign v230bd6c = hlock0_p & v22ee92e | !hlock0_p & v22fe963;
assign v230aa63 = hbusreq3 & v22fb00c | !hbusreq3 & !v845625;
assign v23f77e8 = hlock1_p & v22feb47 | !hlock1_p & !v84561b;
assign v2305522 = hgrant0_p & v22f8271 | !hgrant0_p & v23fccd5;
assign v23fbb28 = hgrant3_p & v22f6ae5 | !hgrant3_p & v23fb52d;
assign v230c949 = hmaster0_p & v22f6169 | !hmaster0_p & v23fc815;
assign v2308786 = hgrant1_p & v12cd6a1 | !hgrant1_p & v23fcfb7;
assign v23f41b9 = hmaster2_p & v23f5af5 | !hmaster2_p & !v106ae19;
assign v23fbd7d = hmaster0_p & v22f789c | !hmaster0_p & v22f4d28;
assign v23f72fe = hbusreq4 & v191ab29 | !hbusreq4 & v2302131;
assign e1e353 = hmaster2_p & v22f53c0 | !hmaster2_p & v23f660f;
assign v1aad9a6 = hbusreq5 & v23f6b67 | !hbusreq5 & v84561b;
assign v23f1a1c = hbusreq1_p & v230beed | !hbusreq1_p & !v84561b;
assign v22f5828 = hbusreq3 & v23f4c50 | !hbusreq3 & !v84561b;
assign v22ebc8f = hbusreq4_p & v23fc56c | !hbusreq4_p & v23fc1a1;
assign v22fc96c = hgrant1_p & v230997b | !hgrant1_p & a68bda;
assign v230160e = hmaster2_p & v23f8928 | !hmaster2_p & v230db4e;
assign v22ec921 = hbusreq2_p & v22efc3c | !hbusreq2_p & !v84561b;
assign v22f666d = hmaster2_p & v2311d0c | !hmaster2_p & v191a86f;
assign v23126f2 = hgrant1_p & v845626 | !hgrant1_p & v22f9fe0;
assign v2301292 = hlock4_p & v230eed2 | !hlock4_p & v22ec0d1;
assign v23fcd00 = hgrant1_p & v23fc9dd | !hgrant1_p & !v84561b;
assign v22f5204 = hmaster2_p & v2307758 | !hmaster2_p & v22ef217;
assign v23fc2ee = hbusreq0 & v845629 | !hbusreq0 & !v84561b;
assign v23f74bf = hbusreq3_p & v2307206 | !hbusreq3_p & v23fbd2a;
assign v230a1c7 = hmaster2_p & v23fbaaa | !hmaster2_p & v239346f;
assign v2393c48 = hgrant3_p & v845647 | !hgrant3_p & v23f4b99;
assign v23fcc6c = hmaster0_p & v23096f8 | !hmaster0_p & v23fc29d;
assign v2308609 = hmaster0_p & v84561b | !hmaster0_p & !v23fafe3;
assign v22eafd6 = hbusreq6 & v22f2ece | !hbusreq6 & v84561b;
assign v9a3d0c = hbusreq4_p & v230c84d | !hbusreq4_p & v22ed48e;
assign v895d68 = hmaster2_p & v22feb47 | !hmaster2_p & v22f337b;
assign v230fe9b = hmaster0_p & v22ef62d | !hmaster0_p & ad89b5;
assign v23fbafd = hlock2_p & da38c1 | !hlock2_p & v84561b;
assign v23f2bc5 = hbusreq4 & v23089a5 | !hbusreq4 & v84564d;
assign v191aada = hgrant5_p & v23efc12 | !hgrant5_p & !v22eff6d;
assign v23f6cc2 = hmaster0_p & v230ea9f | !hmaster0_p & !v23f7561;
assign v22f792a = hlock1_p & v23f4a16 | !hlock1_p & v845620;
assign v231363c = hbusreq3_p & v230607d | !hbusreq3_p & !v22f57e9;
assign v22ffcec = hmaster0_p & v22fec1c | !hmaster0_p & v22fd2ac;
assign v22f709c = hgrant3_p & f40a8f | !hgrant3_p & v22ed7a5;
assign v23f4b8f = hmaster0_p & v22f58c2 | !hmaster0_p & v23f59dc;
assign v22ec303 = hlock0_p & v23fbb35 | !hlock0_p & !v84561b;
assign v22fab90 = hmaster0_p & v23fafaf | !hmaster0_p & baa1eb;
assign v23fbf0d = hgrant1_p & v84561b | !hgrant1_p & !addc42;
assign v23fb0c7 = hbusreq4_p & e1deb1 | !hbusreq4_p & v23014b0;
assign e1e1d4 = hmaster2_p & v23fc22e | !hmaster2_p & v23fbaaa;
assign v22f95c1 = hbusreq3_p & v23fc85c | !hbusreq3_p & v230a759;
assign v22f1e6a = hbusreq6_p & v9ed9e1 | !hbusreq6_p & v23fb242;
assign v22fb850 = hbusreq1_p & v230a9d5 | !hbusreq1_p & v23fccf8;
assign v22fc3c4 = hbusreq5_p & v845636 | !hbusreq5_p & v22f3bc9;
assign v230b4af = hbusreq1_p & v23fc064 | !hbusreq1_p & v230e872;
assign v22f6cde = hbusreq3_p & v23fc001 | !hbusreq3_p & v23fc60a;
assign v23fbf5d = hmaster2_p & v23f4b28 | !hmaster2_p & v23035ba;
assign v23fcb0d = hmaster0_p & v23fc92c | !hmaster0_p & v2301a67;
assign v230d2b0 = hbusreq3_p & v2308a32 | !hbusreq3_p & !v84561b;
assign v22fa5a5 = hbusreq5_p & v22ecc15 | !hbusreq5_p & v2392d6d;
assign v23fb586 = hgrant3_p & v84561b | !hgrant3_p & v23fc0d0;
assign v22fc1e9 = hbusreq3 & v23fc6ef | !hbusreq3 & v23027cd;
assign v2308f46 = hlock5_p & v230de4d | !hlock5_p & v1e84184;
assign b1d009 = hlock4_p & v22eb23c | !hlock4_p & v22eaeaf;
assign v88c9bf = hgrant1_p & v845626 | !hgrant1_p & v22fc7c2;
assign v23f6827 = hmaster0_p & v23fd01e | !hmaster0_p & v22f9a50;
assign v22f1762 = hmaster2_p & v23f8da8 | !hmaster2_p & v84561b;
assign v23f3a5b = hbusreq3 & v23f21c1 | !hbusreq3 & v23fc5e8;
assign v22ebedd = hgrant1_p & v22f7aff | !hgrant1_p & !v22eb6fc;
assign v230ec2b = hmaster0_p & v22fb465 | !hmaster0_p & v22f7c6f;
assign v23fce78 = hmaster0_p & v23fc525 | !hmaster0_p & v22fe052;
assign v22ec2c0 = hbusreq4_p & v23f5dfd | !hbusreq4_p & !v22edc69;
assign v2307a9e = hbusreq6_p & v230e794 | !hbusreq6_p & v230be37;
assign v22f69aa = hmaster2_p & v23f9f07 | !hmaster2_p & v22fe346;
assign v23fbc9f = hbusreq6 & v23093e2 | !hbusreq6 & v84561b;
assign v2307081 = hmaster0_p & v2312ec4 | !hmaster0_p & v1b876be;
assign v23f1ff1 = jx0_p & v22f52f0 | !jx0_p & v2306b1d;
assign v230eed5 = hlock6_p & v23fc26c | !hlock6_p & !v22ffdc9;
assign v2311106 = hgrant5_p & v22f1d92 | !hgrant5_p & !v84561b;
assign v22ed6ac = stateG10_5_p & v230397f | !stateG10_5_p & v845636;
assign v2304ed3 = hbusreq0 & v23fb9ad | !hbusreq0 & v84561b;
assign v23f9d0b = hbusreq3_p & v22f854f | !hbusreq3_p & v23f57c1;
assign v2306b74 = hbusreq0 & v1aae98c | !hbusreq0 & v23fa2ec;
assign v23f8a29 = hmaster2_p & v23f9414 | !hmaster2_p & v23f7ab7;
assign v22ed01c = hbusreq3_p & v23051cf | !hbusreq3_p & v23fc2d7;
assign v23fbada = hbusreq5_p & v230a9eb | !hbusreq5_p & v22eb9e7;
assign v2392023 = hbusreq6_p & v23f5ae3 | !hbusreq6_p & v1aae296;
assign v2301a5f = hmaster0_p & v22f82cd | !hmaster0_p & v23fb937;
assign v2303a7f = hgrant2_p & v23fbbc7 | !hgrant2_p & !v84561b;
assign v2301a76 = hbusreq6_p & v2304e28 | !hbusreq6_p & v1aae296;
assign v22f6d27 = jx1_p & v230649c | !jx1_p & v231016f;
assign v22fd19c = hbusreq1 & v22eeb07 | !hbusreq1 & !v845636;
assign v2304edd = stateG10_5_p & v84561b | !stateG10_5_p & v2309891;
assign v22fc365 = jx1_p & v23f6adf | !jx1_p & v231220c;
assign v23fc541 = hmaster2_p & v23046f7 | !hmaster2_p & !v2302e32;
assign v230ccc4 = hmaster2_p & v22eeb03 | !hmaster2_p & !v23f5cb3;
assign v23f3ed0 = hmaster1_p & v22ebbde | !hmaster1_p & v2301b99;
assign v22ef31d = hlock3_p & v2312236 | !hlock3_p & !v106ae19;
assign v2301b52 = hgrant3_p & v22f368e | !hgrant3_p & v22fc5d8;
assign v23f391e = hready & v23f7326 | !hready & v22f197e;
assign v22f6f7e = hgrant6_p & v23f7a6d | !hgrant6_p & v2308277;
assign v2305de3 = hgrant0_p & v230fb99 | !hgrant0_p & v22f9838;
assign v1aadf33 = hbusreq3_p & v23fcffb | !hbusreq3_p & v23fb18d;
assign v23fc6a2 = hgrant3_p & v230ab24 | !hgrant3_p & v230ec1c;
assign v1aae9f4 = hbusreq4_p & v22ef61b | !hbusreq4_p & v231094e;
assign v22f5b58 = hbusreq3_p & v22fdafe | !hbusreq3_p & v23faacb;
assign v23fb9ff = hbusreq2_p & v22f0810 | !hbusreq2_p & !v84561b;
assign v230a2b1 = hbusreq1_p & v22f08d0 | !hbusreq1_p & v230df19;
assign v23fc198 = hgrant1_p & v230c5ea | !hgrant1_p & v23fcb47;
assign v22f2b52 = hmaster2_p & v23f4855 | !hmaster2_p & v230a51c;
assign v23fba65 = hgrant1_p & v23fcf46 | !hgrant1_p & v23fa8d7;
assign v23025e4 = hmaster2_p & v191a879 | !hmaster2_p & !v22eb1f5;
assign v863ce5 = stateG3_2_p & v84561b | !stateG3_2_p & v22f476c;
assign v2392c41 = hlock1_p & v23fc6d3 | !hlock1_p & v23f99cf;
assign v15074d0 = hbusreq6_p & v2306e0e | !hbusreq6_p & v23fb094;
assign v22f1e81 = hbusreq6_p & v1507631 | !hbusreq6_p & v12cd8ed;
assign v230020c = hmaster0_p & v2306875 | !hmaster0_p & v91ff8a;
assign v23f493a = hbusreq6_p & v22fdba7 | !hbusreq6_p & v22f3d67;
assign v2303535 = hgrant2_p & v191aea6 | !hgrant2_p & v84561b;
assign v23f7aba = hbusreq3_p & v230468d | !hbusreq3_p & v230a44f;
assign a1fba6 = hmastlock_p & v22ec87b | !hmastlock_p & v84561b;
assign v22fb74c = hgrant1_p & v17a34ff | !hgrant1_p & v23f5a8b;
assign v23f34d7 = hbusreq4_p & v230b464 | !hbusreq4_p & v84561b;
assign v230f43d = hgrant1_p & v2301e9c | !hgrant1_p & !v84561b;
assign v23124e2 = hgrant5_p & v84561b | !hgrant5_p & v22fc03b;
assign v23079bc = hmaster2_p & v23f2ec0 | !hmaster2_p & v84561b;
assign v9c12cb = hgrant5_p & v2308c31 | !hgrant5_p & v23fbed3;
assign v191b187 = hlock0_p & bda6a0 | !hlock0_p & !v84561b;
assign v23f317c = hbusreq3_p & v22eaee1 | !hbusreq3_p & !v22ec882;
assign v23f9dd8 = hmaster1_p & v23f7a92 | !hmaster1_p & v2305660;
assign v230ee7d = hbusreq5 & v845620 | !hbusreq5 & v22ef683;
assign v22fc8c8 = hbusreq2_p & v22f9b42 | !hbusreq2_p & v84561b;
assign a0d50a = stateG10_5_p & v23fc36e | !stateG10_5_p & v22f4163;
assign v231033b = hbusreq1_p & v22efee2 | !hbusreq1_p & v84561b;
assign v23fcb29 = hmaster1_p & v22f00b6 | !hmaster1_p & v23f724e;
assign v23f2278 = stateG2_p & v84561b | !stateG2_p & v23f732a;
assign v23f513d = hbusreq3 & v2309320 | !hbusreq3 & v230fc56;
assign v23ef915 = hbusreq3_p & v23fc27c | !hbusreq3_p & !v84561b;
assign v22f8a46 = hbusreq3_p & v22f7ec9 | !hbusreq3_p & v23f39e6;
assign v23f1387 = hbusreq3 & v23f1fad | !hbusreq3 & !v84561b;
assign v23f8d1a = hmaster0_p & v22fa4df | !hmaster0_p & v23f4451;
assign v23001a6 = hbusreq6 & v23fc11a | !hbusreq6 & v84561b;
assign v2393392 = hlock3_p & v23f9150 | !hlock3_p & v106ae19;
assign v230b02b = hbusreq0 & v23023c9 | !hbusreq0 & v23fcd1b;
assign v22f8594 = stateG10_5_p & v23f80e9 | !stateG10_5_p & v23fb1c6;
assign v23f6032 = hlock4_p & v23fcbaf | !hlock4_p & !v230f549;
assign v2311df1 = hmaster0_p & v22f1a14 | !hmaster0_p & !v2303598;
assign v2302dca = hmaster0_p & v230bf72 | !hmaster0_p & v9ed019;
assign v22f2214 = hbusreq4_p & v22f5076 | !hbusreq4_p & v23f89fd;
assign v2393064 = hbusreq3 & v23fc72d | !hbusreq3 & v84561b;
assign v23f9395 = hmaster2_p & b09503 | !hmaster2_p & v84561b;
assign v2312301 = hbusreq6_p & v12cd632 | !hbusreq6_p & v2311645;
assign v2305aee = jx3_p & v230ecba | !jx3_p & v84561b;
assign v22f4bec = hbusreq5_p & v2304b9d | !hbusreq5_p & v23fcafe;
assign v22ed5e6 = stateG2_p & v84561b | !stateG2_p & v23055d4;
assign v23f7456 = hmaster1_p & v84561b | !hmaster1_p & v22f9a6b;
assign v2309efb = hbusreq3_p & v2300ba2 | !hbusreq3_p & v84561b;
assign v23fa7ec = hlock5_p & v84561b | !hlock5_p & v23fb798;
assign v2300df6 = hmaster2_p & v23fcac2 | !hmaster2_p & v23fc7ef;
assign v22f8aba = hbusreq1_p & v23fbfc9 | !hbusreq1_p & v845620;
assign v23fc152 = hbusreq3_p & v22f2bab | !hbusreq3_p & v22f68e5;
assign v22f7371 = hbusreq6_p & v230267d | !hbusreq6_p & v230197f;
assign v23fc70f = jx3_p & v23fbea4 | !jx3_p & v2306fae;
assign v22f2f26 = hmaster2_p & v22f64b2 | !hmaster2_p & !v106ae19;
assign v23fc133 = hbusreq5_p & v84561b | !hbusreq5_p & v22f4bca;
assign v23f1e72 = hbusreq0 & v23fcb5b | !hbusreq0 & v191aa95;
assign v22f9b3f = hbusreq6_p & v22fab90 | !hbusreq6_p & v106ae3a;
assign v23fcab3 = hmaster0_p & v23fc89e | !hmaster0_p & !v22fccbd;
assign v22ebed1 = hgrant3_p & v23f120d | !hgrant3_p & v23f18da;
assign v23f4b9c = hbusreq4_p & v22f7277 | !hbusreq4_p & v2302844;
assign v23fccbe = hlock0_p & v2306d29 | !hlock0_p & v22ecc3f;
assign v23f54e8 = hmaster0_p & v23f99ec | !hmaster0_p & v23916b5;
assign v230049a = hmaster1_p & v22fd5fc | !hmaster1_p & v23927e4;
assign v94116b = hbusreq6_p & v22f737d | !hbusreq6_p & f40cfd;
assign v2301a04 = hmaster2_p & v23f60ef | !hmaster2_p & v84562a;
assign v230d0ed = hbusreq4_p & v22f1324 | !hbusreq4_p & v22f3586;
assign v2312ad2 = hgrant1_p & v84561b | !hgrant1_p & !v2311106;
assign v230f330 = hbusreq3_p & v22f65b0 | !hbusreq3_p & v22f3206;
assign v23fb526 = hgrant3_p & v1aada8c | !hgrant3_p & v2392868;
assign v2303996 = hbusreq0 & v23f54ac | !hbusreq0 & v84561b;
assign v22fc4a3 = hmaster2_p & v23fc658 | !hmaster2_p & !v84561b;
assign v23f841d = hbusreq1 & v13afe3a | !hbusreq1 & !fc8e3a;
assign fc88bb = jx0_p & v23fc342 | !jx0_p & v22fdc2b;
assign v23fc08c = hmaster1_p & v230702c | !hmaster1_p & v23fb877;
assign bdab35 = jx0_p & v22f94c1 | !jx0_p & !v23f623e;
assign v2312be4 = hbusreq4_p & v2391a4f | !hbusreq4_p & v230dec9;
assign v22f1683 = hmaster0_p & v2310319 | !hmaster0_p & v23fb9ef;
assign v23f64d3 = jx3_p & v84561b | !jx3_p & v2309cda;
assign v23f273d = hmastlock_p & v22f235b | !hmastlock_p & !v84565f;
assign v23fce15 = hbusreq3 & v22f0b56 | !hbusreq3 & v84561b;
assign v2313131 = hgrant1_p & v84561b | !hgrant1_p & !v23fc6b1;
assign v22f7a20 = hgrant3_p & v22eb51e | !hgrant3_p & v230f9c2;
assign v22fc0a4 = hbusreq3_p & v23018a8 | !hbusreq3_p & v22ff4e2;
assign v2308706 = hbusreq6 & v106af3a | !hbusreq6 & v22f2ca2;
assign v22f8694 = hbusreq1_p & v191afad | !hbusreq1_p & v22ebfa3;
assign v22fbc4e = jx2_p & v23f5767 | !jx2_p & v23fc2d8;
assign v23123b4 = hbusreq1_p & v22f79be | !hbusreq1_p & v22f6d58;
assign v2391fb2 = hmaster2_p & v22f3618 | !hmaster2_p & v23f940c;
assign v230e1e4 = hmaster0_p & v23fba43 | !hmaster0_p & v23fc44e;
assign v23f99f6 = hgrant1_p & v84561b | !hgrant1_p & v23fc341;
assign v22f1412 = hgrant2_p & v84562a | !hgrant2_p & !v23f2eb5;
assign v22fb8c0 = hbusreq4_p & v23f66db | !hbusreq4_p & v22f88bb;
assign b63b0c = hmaster2_p & v22fe5b1 | !hmaster2_p & !v2303831;
assign v22ef750 = hmaster2_p & v23f9c45 | !hmaster2_p & v1aadac4;
assign v22f7ca0 = stateG2_p & v84561b | !stateG2_p & v2393e5c;
assign v22f97c3 = hbusreq6 & v230b23c | !hbusreq6 & v84561b;
assign v22f0ecb = hgrant0_p & v84561b | !hgrant0_p & v2303352;
assign v23fcd0b = hmaster2_p & v23f77e8 | !hmaster2_p & v22f337b;
assign v23fc02a = hmaster2_p & v23f5cb3 | !hmaster2_p & !v23fc127;
assign v22fa889 = hmaster2_p & v895ae7 | !hmaster2_p & v23fc38f;
assign v22fa345 = hbusreq5 & v1aae56f | !hbusreq5 & v84564d;
assign v230dd17 = hbusreq6_p & v23f567b | !hbusreq6_p & v22ebc28;
assign v2310747 = hbusreq4_p & v23fc887 | !hbusreq4_p & a1fdf8;
assign v22f7466 = hgrant1_p & v23f794b | !hgrant1_p & v22f7efd;
assign v2312526 = hbusreq1 & v23f0169 | !hbusreq1 & v2304536;
assign v23fcdd8 = hbusreq3_p & v230ac22 | !hbusreq3_p & v22ee657;
assign v22fb011 = hbusreq4_p & v230790b | !hbusreq4_p & v230f0de;
assign v23fb8fc = hgrant0_p & v23f11a3 | !hgrant0_p & !v15070d3;
assign v23fba06 = hbusreq3_p & v230e857 | !hbusreq3_p & v23f0588;
assign v23fb029 = hbusreq5_p & v23f3a16 | !hbusreq5_p & v2309871;
assign v230cb59 = hlock1_p & v23fbb41 | !hlock1_p & v2312351;
assign v22ed1a8 = hbusreq3 & v23fb504 | !hbusreq3 & v84561b;
assign v22f1866 = hmaster2_p & v22fb8d6 | !hmaster2_p & !v22ec782;
assign v22ed291 = hbusreq4_p & v23fbd46 | !hbusreq4_p & v23133fe;
assign v23fc8e5 = hbusreq6_p & v22eb0b3 | !hbusreq6_p & v1aad703;
assign v231181c = hmaster0_p & v23fcf07 | !hmaster0_p & v2308a75;
assign v23fbb89 = hgrant5_p & v22eb771 | !hgrant5_p & v84561b;
assign v22fd0b6 = hmaster0_p & v22ff0d3 | !hmaster0_p & v22f1ab6;
assign v23fbe41 = locked_p & v22ebccb | !locked_p & v23fc8be;
assign v23fcfa5 = hbusreq6 & v23fc273 | !hbusreq6 & v23f87f4;
assign v23fceca = hlock3_p & v22ec330 | !hlock3_p & v23124aa;
assign fc90a8 = hmaster0_p & v23fccdb | !hmaster0_p & v230bd1b;
assign v22ffaf3 = hbusreq6_p & v23f2df7 | !hbusreq6_p & v23fd04d;
assign v22faef8 = hbusreq2 & v23fb054 | !hbusreq2 & v84561b;
assign fc8f82 = hbusreq5 & v191a876 | !hbusreq5 & !v84561b;
assign v22f1992 = hgrant2_p & v23f5d7f | !hgrant2_p & v23f8979;
assign v23fcd83 = jx1_p & v22edcce | !jx1_p & v230e1e0;
assign v23fbe3a = hbusreq3_p & v22f8240 | !hbusreq3_p & v22ed5fd;
assign v23fa4bd = hbusreq1_p & v22fa56f | !hbusreq1_p & v84561b;
assign v230f4d0 = hbusreq3_p & v23f0c76 | !hbusreq3_p & !v23f513d;
assign v23fbcac = hgrant3_p & v22ffa6e | !hgrant3_p & v2300523;
assign v935301 = hgrant4_p & v22eb83a | !hgrant4_p & v230717d;
assign v23f29f5 = hlock4_p & v23f5f78 | !hlock4_p & v23fc738;
assign v23f14bc = hgrant1_p & v84561b | !hgrant1_p & v22ed614;
assign v23f5269 = hgrant1_p & v84561b | !hgrant1_p & v230b313;
assign v23f0903 = hbusreq1_p & v23f8c7b | !hbusreq1_p & f40a94;
assign v22f00c6 = hmaster2_p & v9526ac | !hmaster2_p & a1fba6;
assign v22ebd85 = hmaster0_p & v2312cd5 | !hmaster0_p & v84561b;
assign v23fbe26 = hbusreq3 & v22f7ec9 | !hbusreq3 & !v84561b;
assign v22f7859 = hlock1_p & v23fceb9 | !hlock1_p & v84562b;
assign v845657 = hgrant4_p & v84561b | !hgrant4_p & !v84561b;
assign v22f8894 = hmaster0_p & v230b131 | !hmaster0_p & v22f5f28;
assign v2393c3f = hmaster1_p & v23f223a | !hmaster1_p & v23fd00e;
assign v23fc31c = jx3_p & v23076ca | !jx3_p & v2346b90;
assign v23fc5be = hmaster2_p & v2302d97 | !hmaster2_p & v84561b;
assign v23fafc1 = stateG10_5_p & v22f8107 | !stateG10_5_p & !v22ef1a3;
assign v23130d6 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v230320e;
assign v191a912 = hmaster2_p & v23fb5a1 | !hmaster2_p & v84561b;
assign v23fc1a3 = hgrant0_p & v22ecc25 | !hgrant0_p & v2302933;
assign v150705a = stateG10_5_p & v22f1dab | !stateG10_5_p & v22ff732;
assign v23fcb6d = hmaster0_p & v23f6ad0 | !hmaster0_p & !v23fb0f0;
assign v22eb69b = jx3_p & v230a77a | !jx3_p & v23041ed;
assign v23fc04c = hbusreq1_p & v23f6e45 | !hbusreq1_p & v84562b;
assign v23925e9 = hgrant3_p & v23034f8 | !hgrant3_p & v23fcd6b;
assign v2309a78 = hbusreq0_p & v23f6411 | !hbusreq0_p & !b9d013;
assign v23f6e78 = hmaster2_p & v84561b | !hmaster2_p & !v23fc7d5;
assign v2302f85 = hmaster2_p & v22f5583 | !hmaster2_p & !v23108b7;
assign v23fc5ca = jx0_p & v23fcb09 | !jx0_p & v22efcbf;
assign v22f4d77 = hbusreq6 & v23087d7 | !hbusreq6 & v2303e4f;
assign v230b3d5 = hmaster2_p & v191a86f | !hmaster2_p & v23041e2;
assign fc8f72 = hbusreq5_p & v23fc9d2 | !hbusreq5_p & v23f9c30;
assign v2311891 = hbusreq5 & c258f4 | !hbusreq5 & v22fa707;
assign v1aae2a5 = hbusreq4 & v949c12 | !hbusreq4 & v84562f;
assign v23fcfe4 = hbusreq3_p & v230e689 | !hbusreq3_p & v22ebd88;
assign c0e31a = hmaster2_p & v23f8928 | !hmaster2_p & v23f8679;
assign v22ed49b = hgrant0_p & v230219b | !hgrant0_p & b159aa;
assign v23fc8d9 = jx0_p & v2305ce8 | !jx0_p & !v23f623e;
assign v23fb3cf = hbusreq2_p & v23007f2 | !hbusreq2_p & !v84561b;
assign v230ebb1 = hmaster2_p & v23101b1 | !hmaster2_p & v23fb999;
assign v230eae5 = hmaster1_p & v22fe62e | !hmaster1_p & v23fc380;
assign v23fc761 = hlock3_p & v230f375 | !hlock3_p & v2309569;
assign v23f5e8a = hmaster2_p & v23fb0ce | !hmaster2_p & v23101b1;
assign v23131a6 = hbusreq3 & v22f8839 | !hbusreq3 & v84561b;
assign v1aae56f = locked_p & v84561b | !locked_p & v191a86f;
assign adf3a3 = hbusreq0 & v23022b1 | !hbusreq0 & !v84561b;
assign v23fc0c6 = hmaster2_p & v23fb5db | !hmaster2_p & v22efa17;
assign v23fa720 = hbusreq5 & v23fc514 | !hbusreq5 & !v23022b1;
assign v22f2bf8 = hbusreq5 & v2310da0 | !hbusreq5 & v84561b;
assign v230beb8 = hbusreq3 & v230e85f | !hbusreq3 & v23fba11;
assign v23faaac = stateG10_5_p & v23fbdf1 | !stateG10_5_p & v845629;
assign v2312f85 = hbusreq1 & v2300827 | !hbusreq1 & v84561b;
assign v22ef6ce = hmaster2_p & v230c0b8 | !hmaster2_p & !v84561b;
assign v230ad95 = hmaster2_p & v106a782 | !hmaster2_p & v2304b4e;
assign v23fbd5f = hbusreq0 & v2308848 | !hbusreq0 & v84561b;
assign v2312608 = hbusreq4 & v23086b9 | !hbusreq4 & v22f4b50;
assign v23fbc48 = hlock0_p & v2309066 | !hlock0_p & !v84561b;
assign v23f9aa8 = hmaster2_p & v231033b | !hmaster2_p & v23fc5ff;
assign v231170f = hlock6_p & v23f5d1a | !hlock6_p & !v22fbb99;
assign v23064ff = hlock1_p & v23045fb | !hlock1_p & !v2300f96;
assign v22f0dd6 = hbusreq1 & v23fba6b | !hbusreq1 & !v84561b;
assign v23fc40f = hbusreq5_p & v2300b96 | !hbusreq5_p & v84561b;
assign v230fae0 = hgrant0_p & v22f824f | !hgrant0_p & v2303dd7;
assign v22f067b = stateG10_5_p & v22f4d68 | !stateG10_5_p & !v84561b;
assign v23fd064 = hbusreq5 & c258f4 | !hbusreq5 & v22ef683;
assign v22fdcc7 = hgrant3_p & v231185d | !hgrant3_p & v23fb23b;
assign v23fc8ef = stateG10_5_p & v2304049 | !stateG10_5_p & v2392833;
assign v22f52a0 = hmaster0_p & v84561b | !hmaster0_p & !v22ef26f;
assign v23026c8 = hgrant1_p & v23fc68c | !hgrant1_p & v23f15af;
assign v22ec21e = hmaster1_p & v23fbf8d | !hmaster1_p & v2304913;
assign v2301392 = hgrant3_p & v22ffa6e | !hgrant3_p & v23f7aba;
assign v22eedcd = hgrant3_p & v23fb6c7 | !hgrant3_p & da310f;
assign v22fa857 = hmaster2_p & v230a890 | !hmaster2_p & v22fd696;
assign v22f009f = hmaster0_p & v2311a61 | !hmaster0_p & v23fbb94;
assign v23f9bf9 = hmaster0_p & v23fc323 | !hmaster0_p & v23fc268;
assign v23fb743 = hbusreq1 & v23f9e4f | !hbusreq1 & v22ff0d7;
assign v23fb1d4 = hgrant0_p & v23127ef | !hgrant0_p & v23fb121;
assign v23fb8fd = jx1_p & v22f07e0 | !jx1_p & v2304193;
assign v23fb8b7 = hbusreq4_p & v22fcef4 | !hbusreq4_p & v23fa36c;
assign v22f3502 = hgrant2_p & v2312283 | !hgrant2_p & !v22fe9b7;
assign v22f0104 = hbusreq6_p & v23fca43 | !hbusreq6_p & v230466c;
assign v23fb622 = hbusreq4_p & v230e97b | !hbusreq4_p & v23fcd5c;
assign v230e1fc = hmastlock_p & v22f97e9 | !hmastlock_p & v84561b;
assign v230b62c = hgrant1_p & v23f6653 | !hgrant1_p & v230f573;
assign v23f4a16 = hbusreq1 & v2313118 | !hbusreq1 & v23f1879;
assign v239298c = stateG2_p & v84561b | !stateG2_p & !v23f906a;
assign v23fca7a = hbusreq3_p & v23fc6c2 | !hbusreq3_p & !v84561b;
assign v23fbd79 = hmaster2_p & v23126f2 | !hmaster2_p & v22fc741;
assign v22f274e = hgrant1_p & v84561b | !hgrant1_p & v2302022;
assign v2300c85 = hbusreq4 & v845620 | !hbusreq4 & v23fb0bb;
assign v230440f = hbusreq6_p & v22ec5d6 | !hbusreq6_p & v23f7b85;
assign v23fcf22 = hmaster0_p & v23f592d | !hmaster0_p & v23f47e1;
assign v22f39b4 = hbusreq6 & v22ec552 | !hbusreq6 & !v84561b;
assign v23fcedb = hmaster2_p & v22ee339 | !hmaster2_p & v23fc9d3;
assign v9799b6 = hgrant3_p & v23fb17e | !hgrant3_p & !v1aadf2f;
assign v22ff184 = hbusreq6_p & v22ffcb0 | !hbusreq6_p & !v84561b;
assign v23fb669 = hbusreq0 & v23fbd16 | !hbusreq0 & v23f039f;
assign v22fd72d = hbusreq1 & v22f1403 | !hbusreq1 & v84561b;
assign v23f3d62 = hbusreq3_p & v22fc9ad | !hbusreq3_p & !v84561b;
assign v23fc3d8 = hmaster1_p & v230bc37 | !hmaster1_p & v2310037;
assign v22fa631 = hmaster2_p & v23fceb9 | !hmaster2_p & v84561b;
assign v23fbdc2 = hbusreq6 & v22f4d61 | !hbusreq6 & e1bfb3;
assign v22fa440 = stateG10_5_p & v22f7f74 | !stateG10_5_p & v22f9980;
assign v22fa682 = hgrant5_p & v23fbcff | !hgrant5_p & v22f6058;
assign b42c55 = hmaster1_p & v2311f44 | !hmaster1_p & v2310f12;
assign v2308d80 = hmaster2_p & v2308110 | !hmaster2_p & !v23fb98e;
assign v23130d9 = hmaster0_p & v23fba43 | !hmaster0_p & v22f959d;
assign v23f5207 = hmaster2_p & v23fcf69 | !hmaster2_p & v23f8f25;
assign v22ed2e5 = hbusreq1_p & v230cec5 | !hbusreq1_p & !v84561b;
assign v23fc8a9 = hbusreq4_p & v22ee920 | !hbusreq4_p & v22fdcc5;
assign v23f5ac2 = hgrant3_p & v84561b | !hgrant3_p & v23fa600;
assign v230cffc = hmaster0_p & v23fbcfd | !hmaster0_p & !v23f982d;
assign v2392d0d = hbusreq4_p & v23f7f51 | !hbusreq4_p & v22ecd9e;
assign v23f9c30 = hgrant0_p & v23133fa | !hgrant0_p & v2392e9d;
assign v1aadeea = hbusreq6_p & v23f5a4e | !hbusreq6_p & v84561b;
assign v23074c0 = hlock3_p & fc907f | !hlock3_p & v239353f;
assign v2307460 = stateG2_p & v84561b | !stateG2_p & v22ed56a;
assign v2310ec5 = hbusreq3_p & v23fbb5a | !hbusreq3_p & v22fa58f;
assign v230cfb5 = hmaster0_p & v22f6629 | !hmaster0_p & !v23105b1;
assign v23065fc = hbusreq3_p & v2304bc1 | !hbusreq3_p & !v23f946b;
assign v23fc2b7 = hgrant3_p & v230a744 | !hgrant3_p & v22ff9c3;
assign bd757c = stateG2_p & v23fc331 | !stateG2_p & v2310c2b;
assign v23fbb8b = hgrant0_p & v23fb109 | !hgrant0_p & v23fc56f;
assign v22efd1a = hbusreq2 & v22fcdf6 | !hbusreq2 & v84564d;
assign v22fcf75 = hmaster2_p & v22f4114 | !hmaster2_p & bd74ad;
assign v23fbf31 = hbusreq3_p & v23fba74 | !hbusreq3_p & v22fe7ca;
assign v22fdd61 = hlock4_p & v230e962 | !hlock4_p & !v23fc7dc;
assign v23fb1e1 = hbusreq1_p & v2300cbb | !hbusreq1_p & v84561b;
assign v23fcdbe = hgrant1_p & v12cc2ef | !hgrant1_p & v23fcdb2;
assign v23fcf6b = jx2_p & v23fb64e | !jx2_p & v22f6955;
assign v23f07c2 = hbusreq6_p & v22f155f | !hbusreq6_p & v22f43d7;
assign v2304be0 = hbusreq3 & v22fe44f | !hbusreq3 & !v84561b;
assign v23f1bd6 = hmaster0_p & v22f3ac3 | !hmaster0_p & b9c90c;
assign v230d4b4 = hgrant0_p & v84561b | !hgrant0_p & v8b5388;
assign v2311eaa = hmaster0_p & v23fa8d8 | !hmaster0_p & v23fc9a5;
assign v230be4a = hmaster2_p & v22fc2bd | !hmaster2_p & v2302225;
assign v23f5513 = hmaster2_p & v23fcd2d | !hmaster2_p & v84564d;
assign v2309b33 = hbusreq3_p & v22f9eb0 | !hbusreq3_p & v23f963f;
assign v23fcd5d = hbusreq0 & v23f1207 | !hbusreq0 & v230b1ac;
assign v2311919 = hbusreq6_p & v23fb90b | !hbusreq6_p & v23fc2bc;
assign v23fcc28 = hbusreq2 & v230882d | !hbusreq2 & v23f8364;
assign v22fbbd2 = jx3_p & v23037f2 | !jx3_p & v23113f1;
assign v2307483 = hbusreq3_p & v2312a3d | !hbusreq3_p & v2313131;
assign v2302a2c = hbusreq0_p & v845620 | !hbusreq0_p & v22f79fd;
assign v22fcd49 = hmaster0_p & v23fc43d | !hmaster0_p & b00aa6;
assign v22ed6c5 = locked_p & v84561b | !locked_p & v23fba6b;
assign v2300829 = hmaster2_p & v23f15ac | !hmaster2_p & v2300071;
assign v22edb0c = hbusreq0 & v23fc346 | !hbusreq0 & v84561b;
assign a4c16b = hbusreq3_p & v23fc1a2 | !hbusreq3_p & v22f8da4;
assign v22ff1ee = hgrant2_p & v23fbe41 | !hgrant2_p & v23fc2d2;
assign v22f6b57 = hbusreq6_p & v23fbcc2 | !hbusreq6_p & v230ce74;
assign v22f448e = hbusreq4_p & v22ff192 | !hbusreq4_p & v22f0210;
assign v23f894b = hmastlock_p & v23026db | !hmastlock_p & v84561b;
assign v22f3b94 = hbusreq2_p & v23fbae2 | !hbusreq2_p & v84564d;
assign v22f0dc3 = hbusreq3 & v23fcb7c | !hbusreq3 & v230554d;
assign v23f8b5b = hmaster0_p & v23fc8d6 | !hmaster0_p & v230bd77;
assign v23010d9 = hmaster2_p & v22f8e9a | !hmaster2_p & v23f660f;
assign v22ef9ea = hbusreq6_p & v23fb492 | !hbusreq6_p & v23129c2;
assign v963cc3 = hlock6_p & v87eb7a | !hlock6_p & v23139b9;
assign v2302cf5 = hgrant3_p & v84561b | !hgrant3_p & v22fd171;
assign v2312fc4 = hmastlock_p & v22f0bea | !hmastlock_p & v84561b;
assign v2307de6 = hmaster2_p & v1aad5ad | !hmaster2_p & v23fceb9;
assign v17a34e6 = hbusreq2 & v23fc0fc | !hbusreq2 & v84562b;
assign aeff78 = hmaster2_p & v84561b | !hmaster2_p & !v2301319;
assign v23fab81 = jx2_p & v23f1ff1 | !jx2_p & v230b30c;
assign v230f08b = hmaster2_p & v22fee46 | !hmaster2_p & a1fbc2;
assign v23fbf08 = hbusreq0_p & v84561b | !hbusreq0_p & v2310fde;
assign v22f40ef = hmaster2_p & v23fb906 | !hmaster2_p & v22eb404;
assign v22f122e = hgrant1_p & v22ee956 | !hgrant1_p & v22f8387;
assign v23fc636 = stateG10_5_p & v22f41ee | !stateG10_5_p & v22f1aae;
assign v23fbdef = hbusreq1_p & v22f3b33 | !hbusreq1_p & !v23fc2bf;
assign v23fbe7d = hmaster1_p & v23fbea0 | !hmaster1_p & v22ef100;
assign v22f518e = hgrant5_p & v22fecf2 | !hgrant5_p & v23f6bf0;
assign v231140d = hgrant5_p & v230d61c | !hgrant5_p & v22f288e;
assign v23f2eec = hgrant0_p & v23fbcb2 | !hgrant0_p & !v23024b6;
assign v22fc231 = hlock6_p & v23fc5dc | !hlock6_p & v22ec92b;
assign v22ff92c = hgrant3_p & v22f8e29 | !hgrant3_p & v230e3c5;
assign a1fe40 = hbusreq6 & v191aed3 | !hbusreq6 & v84564d;
assign e1e35b = jx1_p & v22f9793 | !jx1_p & v23f7a8e;
assign v23f904c = hmaster0_p & v22f3b15 | !hmaster0_p & v23005ea;
assign v22ff3e6 = hbusreq3_p & v23fba74 | !hbusreq3_p & v23f052e;
assign v23f374e = hmaster2_p & v23f024e | !hmaster2_p & v23f9682;
assign v2392842 = hbusreq5_p & v845636 | !hbusreq5_p & v2302bb2;
assign v22f1d46 = stateG10_5_p & v23f1d8b | !stateG10_5_p & v23046f7;
assign v23fcd81 = hbusreq5_p & v230360b | !hbusreq5_p & v23f3b00;
assign v23fca06 = hlock2_p & v22ee7a7 | !hlock2_p & v84561b;
assign v23fc07c = hmaster2_p & da38c1 | !hmaster2_p & v22f25c6;
assign v230ea78 = hbusreq6_p & ad78c9 | !hbusreq6_p & v22efa95;
assign v23f55c0 = hbusreq0 & v23007a2 | !hbusreq0 & v84561b;
assign v23f864d = hgrant3_p & v22f6d19 | !hgrant3_p & v230f9b8;
assign v23f3321 = hbusreq6 & v230810c | !hbusreq6 & v84561b;
assign v23fc945 = hlock5_p & bbc337 | !hlock5_p & !v230d379;
assign v23fba0c = hbusreq5_p & v8f2065 | !hbusreq5_p & v23f7275;
assign v2392e9d = hlock0_p & a476c2 | !hlock0_p & v231155f;
assign v23fc9c6 = hbusreq2_p & v23f646e | !hbusreq2_p & !v10dbf64;
assign v230edde = hbusreq5_p & v23fc315 | !hbusreq5_p & v2392f21;
assign v2309f3f = hmaster0_p & v2302f63 | !hmaster0_p & v23130dd;
assign v22f6949 = hmaster2_p & v22f9f26 | !hmaster2_p & v23fba9a;
assign v23fcfbe = hlock0_p & v845620 | !hlock0_p & !v84561b;
assign v97ba8e = hmaster2_p & v230b375 | !hmaster2_p & v22fc5e2;
assign v2305ce8 = jx1_p & v85e5cf | !jx1_p & e1e5c9;
assign v22fb062 = hmaster0_p & v230bb08 | !hmaster0_p & !c20a75;
assign v2306d33 = hmaster2_p & v22f11fe | !hmaster2_p & v230a562;
assign v22f35fd = hmaster0_p & v2312da9 | !hmaster0_p & v23fc2fe;
assign v22ebc86 = hlock0_p & v2305a12 | !hlock0_p & v23f1974;
assign v23fc04a = hgrant1_p & v84561b | !hgrant1_p & v2311729;
assign v22fcce6 = hbusreq1 & v13afe8f | !hbusreq1 & !v84561b;
assign v23f794b = hbusreq1_p & v22f7859 | !hbusreq1_p & v84562b;
assign v23f7632 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v23fccbe;
assign v23fc21d = hlock2_p & v2305fe0 | !hlock2_p & v84564d;
assign v23fcec5 = hbusreq3_p & v22fa101 | !hbusreq3_p & v2304583;
assign v22edb40 = hmaster2_p & v22ee9be | !hmaster2_p & v1aad38a;
assign v23f730c = stateG10_5_p & v22ffaff | !stateG10_5_p & v845636;
assign v23fb670 = hlock4_p & v23f7cec | !hlock4_p & !v23132db;
assign v23fc85a = hbusreq5 & v23f40ba | !hbusreq5 & !v84561b;
assign v23f712d = hgrant4_p & v84561b | !hgrant4_p & v23f763a;
assign v23fbbec = hmaster2_p & v84561b | !hmaster2_p & !v23fc46b;
assign v23095d8 = stateG10_5_p & v23fc9d2 | !stateG10_5_p & !v84561b;
assign v23f9fc6 = hmaster0_p & v23139e3 | !hmaster0_p & v1e8404d;
assign v22ef27f = busreq_p & v22f5e60 | !busreq_p & v22f03aa;
assign v22f5033 = jx1_p & v23fcdf8 | !jx1_p & v22ec5ac;
assign v23fcd33 = hgrant5_p & v230f554 | !hgrant5_p & v2346b8a;
assign v23fc016 = hmaster2_p & v22fc564 | !hmaster2_p & v230fc56;
assign v23f35ea = hbusreq3 & v230545b | !hbusreq3 & v22ee6e8;
assign v2302d85 = hlock0_p & v84562a | !hlock0_p & v23fc1de;
assign v23f01f8 = hgrant1_p & v22ff732 | !hgrant1_p & v23fc8d2;
assign v23fca58 = hmastlock_p & v23f7605 | !hmastlock_p & v84561b;
assign v23fcb9d = hbusreq6 & v23fbdb1 | !hbusreq6 & v23fd015;
assign v23fc5b6 = hmaster2_p & v22ffb6b | !hmaster2_p & b7ab40;
assign v23f6591 = hmaster0_p & v2311a61 | !hmaster0_p & v23034e5;
assign v2304bc1 = hlock5_p & v84561b | !hlock5_p & !v845636;
assign v23f7066 = hlock3 & v23fc798 | !hlock3 & e1e1d4;
assign v23fb6a7 = hgrant5_p & v22f9e3d | !hgrant5_p & !v22fe7f5;
assign v23f7039 = hbusreq3_p & c20101 | !hbusreq3_p & v230b4ad;
assign v22fa5b4 = hburst0 & v23fc8a3 | !hburst0 & !v2391ab6;
assign v23f0030 = hlock0_p & v23f01d2 | !hlock0_p & !v84561b;
assign v23130de = hbusreq4 & v23fb5e9 | !hbusreq4 & v230306f;
assign v23fc5dc = hmaster0_p & v23f14e1 | !hmaster0_p & v22ec350;
assign v191abd1 = hgrant3_p & v23f855f | !hgrant3_p & v23f54de;
assign v2300c97 = hlock0_p & v23f450b | !hlock0_p & v13b0013;
assign v22f8549 = hbusreq1_p & b9c955 | !hbusreq1_p & v106a782;
assign v1aad3bf = hgrant6_p & v22f9d57 | !hgrant6_p & v22fff3a;
assign v23fcd63 = hmaster2_p & v22f1244 | !hmaster2_p & v23f99f6;
assign v23fc68c = hbusreq1_p & v22f6ee2 | !hbusreq1_p & !v12cd3f4;
assign v22f09a2 = hmaster1_p & v230a555 | !hmaster1_p & v23fa1e7;
assign v23f8986 = hlock1_p & v23fc453 | !hlock1_p & !v84561b;
assign v230abf9 = hgrant3_p & v84561b | !hgrant3_p & v230b282;
assign v22f3959 = hmastlock_p & v22f9369 | !hmastlock_p & v84561b;
assign v23fbf7f = hbusreq4_p & v23fb8b8 | !hbusreq4_p & !v23fc061;
assign v23fbe89 = hmaster2_p & v13afe3a | !hmaster2_p & !v84561b;
assign v22eb6e2 = jx1_p & v23f17ff | !jx1_p & v22f6618;
assign v22ee338 = hbusreq5 & v84564d | !hbusreq5 & v23fa2ec;
assign v23f1316 = stateA1_p & v22f0362 | !stateA1_p & v230493b;
assign v2391a4f = hmaster0_p & v23fb994 | !hmaster0_p & v23050c3;
assign v23f3f65 = hmaster2_p & v22ebb79 | !hmaster2_p & v23f940c;
assign v23f781b = hgrant3_p & v23fc975 | !hgrant3_p & v23fc555;
assign v22f5e8c = hbusreq0_p & v2306d29 | !hbusreq0_p & v106af73;
assign v23fc023 = hlock0_p & v230287e | !hlock0_p & v845620;
assign v22f4442 = hmaster1_p & v239223a | !hmaster1_p & v22fce1f;
assign v23f5ace = hbusreq3_p & v22f4d97 | !hbusreq3_p & v230547a;
assign v22f67fb = hbusreq6_p & v23f677f | !hbusreq6_p & v23fae22;
assign v23fbacc = hbusreq5_p & v22fb6bf | !hbusreq5_p & v22f9ae9;
assign v23fce61 = hmaster1_p & v22fd841 | !hmaster1_p & v23f147c;
assign v22ebf47 = hmastlock_p & v2300c4a | !hmastlock_p & !v84561b;
assign v23f50bd = hmaster2_p & v23f859a | !hmaster2_p & v23fb9a9;
assign v23f4007 = hbusreq6 & v23fc890 | !hbusreq6 & v23f1812;
assign v22f61b1 = hmaster2_p & v22f954f | !hmaster2_p & v23fb838;
assign v23f4a07 = hbusreq1_p & v23f3d14 | !hbusreq1_p & v22ee9be;
assign v22fe145 = hmaster2_p & bd9c50 | !hmaster2_p & v22fbeea;
assign v23126ae = locked_p & v84561b | !locked_p & v191a876;
assign v23133b7 = hlock6_p & v23f54e8 | !hlock6_p & !v84561b;
assign v230abce = hbusreq1_p & v22fa474 | !hbusreq1_p & !v23fcadf;
assign v23fbf85 = hbusreq3_p & v23fb084 | !hbusreq3_p & v23fc593;
assign v23013a2 = hbusreq6 & v23f6f49 | !hbusreq6 & v23920aa;
assign v23fc468 = hbusreq5 & v23f1207 | !hbusreq5 & b6f86d;
assign v23f5fb5 = hgrant1_p & v84561b | !hgrant1_p & v230d2c7;
assign v22fd841 = hbusreq6_p & v22fe0cb | !hbusreq6_p & v2306da6;
assign v23fc785 = hbusreq4 & v22fda85 | !hbusreq4 & !v84561b;
assign v22ebe46 = hgrant3_p & v23fc430 | !hgrant3_p & v22eef92;
assign v22faa4b = hgrant4_p & v15075f0 | !hgrant4_p & v23fb166;
assign v22fd3f9 = hlock5_p & v230e509 | !hlock5_p & v2310a63;
assign v2303841 = jx1_p & v22fdd6b | !jx1_p & v2310e53;
assign v23f8d9f = hbusreq3_p & v23fc19b | !hbusreq3_p & v22f68e5;
assign v2312d03 = hmaster0_p & v1e840b4 | !hmaster0_p & !v2305c54;
assign v23fc8d4 = hmaster2_p & v1e84174 | !hmaster2_p & v23f8ca4;
assign v22ecb5c = hgrant3_p & v23fab11 | !hgrant3_p & v23f3c28;
assign v2304402 = hbusreq1_p & v23fc6b0 | !hbusreq1_p & !v84561b;
assign v23fbc74 = hmaster0_p & v22f3b08 | !hmaster0_p & v22ff63a;
assign v2308813 = hgrant5_p & v2302520 | !hgrant5_p & v23fb5c4;
assign v230cc4c = hlock5_p & v22eb8b6 | !hlock5_p & !v84561b;
assign v23fbe56 = hlock6_p & v2303d87 | !hlock6_p & v84561b;
assign v22f0785 = hlock2_p & v22ed6c5 | !hlock2_p & v84564d;
assign v23fbe05 = hmaster0_p & v23925a8 | !hmaster0_p & v22f4ee6;
assign v22f3982 = hbusreq3 & v230a2ae | !hbusreq3 & v84561b;
assign v23916ef = hlock4_p & v23044e1 | !hlock4_p & v23fc230;
assign v22fa155 = hgrant5_p & v22f5a29 | !hgrant5_p & v23fcffa;
assign v2311eb3 = hmaster0_p & v22ecde7 | !hmaster0_p & v230f099;
assign v230cc12 = hmaster1_p & v22ee3c9 | !hmaster1_p & v22f8c84;
assign v22eb95e = hmaster1_p & ae1a21 | !hmaster1_p & v2304598;
assign v23fc0a5 = hmaster2_p & v84561b | !hmaster2_p & v22f25c6;
assign v2306b33 = hgrant0_p & v23133fa | !hgrant0_p & !v84561b;
assign e1bacb = decide_p & v22f5e09 | !decide_p & v106a84c;
assign v23071f4 = hmaster1_p & v23fc8bc | !hmaster1_p & v22f668b;
assign v22f4fb8 = hbusreq3_p & v23fc0e0 | !hbusreq3_p & v23fbe27;
assign v23031b6 = hbusreq1_p & v23fc21a | !hbusreq1_p & v23919d4;
assign v22f9ae9 = stateG10_5_p & v12cc72f | !stateG10_5_p & !v84561b;
assign v23066fe = hmaster0_p & b00aa6 | !hmaster0_p & v1e84057;
assign v23fc81b = hlock3_p & v22f031f | !hlock3_p & v23f4fe1;
assign v23f200c = hbusreq3 & v2393f1a | !hbusreq3 & v84561b;
assign v23fc089 = hmaster2_p & v84564d | !hmaster2_p & v23fcc10;
assign v23033d3 = hbusreq3_p & v230200a | !hbusreq3_p & v23025e4;
assign v22efdf3 = hbusreq3_p & v23fc850 | !hbusreq3_p & v22ecff3;
assign v23fc6ab = hmaster2_p & v22fca61 | !hmaster2_p & v84564d;
assign v22fd9a5 = hbusreq3_p & v22ef2be | !hbusreq3_p & v22eea5b;
assign v22f0cc4 = hbusreq1 & v231228e | !hbusreq1 & v84561b;
assign v23066e8 = hbusreq3_p & v22fc32c | !hbusreq3_p & v23fc750;
assign v23fc6b1 = hgrant5_p & v23f6858 | !hgrant5_p & !v84561b;
assign v23fb84b = hbusreq3 & v963922 | !hbusreq3 & v22ff6a2;
assign v230be37 = hbusreq4_p & v22fe820 | !hbusreq4_p & v23fc330;
assign v230e44a = hmaster0_p & v23111d5 | !hmaster0_p & v230206c;
assign v23f2ec0 = hbusreq0_p & v22f6f16 | !hbusreq0_p & v84561b;
assign v23f79b4 = hbusreq1_p & v23f646e | !hbusreq1_p & !v10dbf64;
assign v22fa262 = hmaster2_p & v8d360e | !hmaster2_p & !v1aae29a;
assign v22fc767 = hmaster0_p & v23fbe2d | !hmaster0_p & v2310482;
assign v23fbb44 = hmaster2_p & v85d110 | !hmaster2_p & v22eefd1;
assign v230c4a4 = stateG2_p & v84561b | !stateG2_p & !v22f349a;
assign v22fa3e9 = hgrant1_p & v2307e48 | !hgrant1_p & v84561b;
assign v22fb09f = hbusreq0 & v23f65b4 | !hbusreq0 & !v23009f0;
assign v2306e5a = hmaster2_p & v2313247 | !hmaster2_p & v23080ec;
assign v22f8062 = hbusreq5 & v22eb2f1 | !hbusreq5 & v84561b;
assign e1e5c7 = hmaster2_p & v23f7e43 | !hmaster2_p & v84561b;
assign v23f3166 = hbusreq4_p & f405eb | !hbusreq4_p & v230e04a;
assign v2313266 = hgrant3_p & v23fb8aa | !hgrant3_p & v23f3bcb;
assign v23faab2 = hgrant3_p & v84561b | !hgrant3_p & v23fcb5a;
assign v22f42b0 = stateG10_5_p & v84561b | !stateG10_5_p & v23f68d8;
assign v22f7cab = hgrant0_p & v22f021c | !hgrant0_p & v2307582;
assign v85d975 = hmaster1_p & v2304373 | !hmaster1_p & v845639;
assign v22f8551 = hgrant3_p & v84562e | !hgrant3_p & v2301cee;
assign v230766b = hbusreq2 & v23fba6b | !hbusreq2 & !v84561b;
assign v230cd61 = hlock5_p & v84561b | !hlock5_p & !v23fb218;
assign v22fe426 = hbusreq1_p & v23fc904 | !hbusreq1_p & v230320e;
assign v23134bf = hmaster0_p & v2309a46 | !hmaster0_p & v22ef99b;
assign v22f1339 = hmaster2_p & a3cb61 | !hmaster2_p & v23919f9;
assign v2304b5d = hbusreq5_p & v2309023 | !hbusreq5_p & v845620;
assign v22eefd1 = hlock0_p & v22f8d80 | !hlock0_p & v84561b;
assign v23f24d5 = hbusreq4 & v23f3ff9 | !hbusreq4 & v230f0de;
assign v23fbd2a = hmaster2_p & v2367a45 | !hmaster2_p & v23f471a;
assign v23fae9e = hbusreq1_p & v23f939f | !hbusreq1_p & !v84561b;
assign v22ef734 = hgrant3_p & v84562e | !hgrant3_p & v23fc721;
assign v23fcae8 = hbusreq0_p & v9526ac | !hbusreq0_p & v23f972e;
assign v8bb259 = stateG10_5_p & v230b8cd | !stateG10_5_p & v2309c93;
assign v23130da = hbusreq6 & v230c4e8 | !hbusreq6 & v23044f6;
assign v22ffed0 = jx1_p & v23f23bf | !jx1_p & v84561b;
assign v22ee36e = hbusreq6_p & v1aad527 | !hbusreq6_p & v22fa69c;
assign v23fc3c2 = hgrant3_p & v23fc457 | !hgrant3_p & v22f7098;
assign v23fc8a0 = hbusreq0_p & v22f92ec | !hbusreq0_p & v84561b;
assign v22f4cf3 = busreq_p & v22f4bdf | !busreq_p & d7db8a;
assign v23054ba = stateG10_5_p & v22f852d | !stateG10_5_p & v22f78a9;
assign v23fbc20 = stateG10_5_p & v23f2eec | !stateG10_5_p & !v22f2703;
assign v2310434 = hgrant1_p & v22f3ed0 | !hgrant1_p & f40a94;
assign v2313279 = hmaster0_p & v23fc060 | !hmaster0_p & b9d041;
assign v87d84c = hbusreq3_p & v230b0d6 | !hbusreq3_p & v230e874;
assign v22fe326 = hmaster2_p & v23fcb55 | !hmaster2_p & v230b0f5;
assign v23126c6 = hlock5_p & v2307eee | !hlock5_p & v23fceec;
assign v22fb5f7 = hlock0_p & v845622 | !hlock0_p & v22f8acf;
assign v2305bbb = hgrant3_p & v23f7dbe | !hgrant3_p & v23fc01a;
assign v23f4117 = hbusreq4_p & v23fbdd2 | !hbusreq4_p & v22f8c8d;
assign v23f9a56 = hmaster2_p & v23f7968 | !hmaster2_p & bd7c3f;
assign v23fcaf7 = hmaster2_p & v230b50c | !hmaster2_p & v22f66b0;
assign v22f5164 = hbusreq6 & v2391665 | !hbusreq6 & v84561b;
assign v230345b = hmaster0_p & v22fa4df | !hmaster0_p & v230a730;
assign v23f7326 = stateG2_p & v84561b | !stateG2_p & v23fcb89;
assign v230a6c8 = hlock6_p & v22fdf28 | !hlock6_p & !v23113f5;
assign v23fc721 = hbusreq3_p & v2302ca7 | !hbusreq3_p & v230d3a4;
assign v23f73dd = hmaster2_p & v22f3c9a | !hmaster2_p & v22f19a0;
assign v22f36ff = hready & v2304ec7 | !hready & v230e1fc;
assign v2310f46 = hgrant5_p & v230ea7f | !hgrant5_p & v23060c7;
assign v22f753f = hbusreq2_p & v84561b | !hbusreq2_p & v845620;
assign v22ecc25 = hlock0_p & v22ec53b | !hlock0_p & v22f7159;
assign v22f2e75 = hmaster2_p & v23fc35a | !hmaster2_p & v84561b;
assign v23f35d5 = hgrant5_p & v84561b | !hgrant5_p & v22ff066;
assign v23fcfcf = hbusreq3 & v2312917 | !hbusreq3 & v1e840f2;
assign v23fb92a = hmaster0_p & v22ebc25 | !hmaster0_p & v230bbf8;
assign v23fbf9f = hbusreq5_p & v22ff89d | !hbusreq5_p & v22ec9a7;
assign v22f1bec = stateG10_5_p & v84561b | !stateG10_5_p & v845620;
assign v23fbc06 = hbusreq5_p & v845636 | !hbusreq5_p & v2301d40;
assign v12cd6a1 = hbusreq1_p & v22f1d8b | !hbusreq1_p & b7427f;
assign v23fb299 = hbusreq4_p & v2301450 | !hbusreq4_p & v23fbf5c;
assign v22ee9be = hbusreq0 & v845620 | !hbusreq0 & v84561b;
assign v23100d2 = jx0_p & v23f6ace | !jx0_p & v23faa39;
assign v22f54a0 = hbusreq6_p & v22fe036 | !hbusreq6_p & v22f6053;
assign f405eb = hlock4_p & v94778a | !hlock4_p & v22f44d0;
assign v23fb49a = hbusreq5_p & v22f5611 | !hbusreq5_p & v84561b;
assign v2300de3 = hlock0_p & v22ed85a | !hlock0_p & v23f7aa3;
assign v23fb202 = hmaster1_p & v84561b | !hmaster1_p & !v22f658e;
assign v2304691 = hbusreq1_p & v22fbb54 | !hbusreq1_p & v23effa5;
assign v23fc14b = hbusreq3_p & v22ed83b | !hbusreq3_p & v23091ef;
assign v23fc442 = hbusreq4 & v22ff94b | !hbusreq4 & !v845636;
assign v23fc293 = hbusreq6 & v23fa3fc | !hbusreq6 & v84561b;
assign v22f34d8 = hlock5_p & v22ee338 | !hlock5_p & !v84561b;
assign v22f43fb = stateG10_5_p & v23fc8df | !stateG10_5_p & v22ff732;
assign v23f18a1 = hmaster0_p & v191ab52 | !hmaster0_p & v230913e;
assign v23f7cec = hmaster0_p & v23fc3e8 | !hmaster0_p & !v230e932;
assign v23f69a3 = hbusreq3_p & v23fc96b | !hbusreq3_p & v23fba9a;
assign v23098d3 = hgrant3_p & v84561b | !hgrant3_p & v879c1f;
assign v230d0a3 = hbusreq3 & v23f8913 | !hbusreq3 & v84561b;
assign v22fe0f9 = hlock0_p & v230c104 | !hlock0_p & v84562b;
assign v23f5fa6 = hmaster2_p & v22edf81 | !hmaster2_p & v22ff916;
assign v23f353e = hbusreq4 & v230cbdd | !hbusreq4 & v84561b;
assign v2312a23 = hlock0_p & v23126ae | !hlock0_p & v191a876;
assign v23f60dc = hmaster1_p & v23fcefc | !hmaster1_p & v230e97b;
assign v23f6013 = hgrant6_p & f40618 | !hgrant6_p & v2305339;
assign v23f182c = hmaster2_p & v84561b | !hmaster2_p & v22ff0d7;
assign v23f91a5 = hbusreq1_p & v22ef810 | !hbusreq1_p & v84561b;
assign da3129 = decide_p & v23f3d7d | !decide_p & v23f14c7;
assign v23fc054 = stateG10_5_p & v22ef469 | !stateG10_5_p & v22ff732;
assign v230a555 = hbusreq6_p & v230a3c9 | !hbusreq6_p & v22ee6ce;
assign v23fbd89 = hbusreq1_p & v23fc778 | !hbusreq1_p & !v84561b;
assign v231396f = hbusreq4_p & v22f04ac | !hbusreq4_p & v22f4e9f;
assign v230fce3 = hmaster2_p & v1aae2a8 | !hmaster2_p & v84561b;
assign v23fd049 = hgrant0_p & v23133fa | !hgrant0_p & e1ddd0;
assign v23fc180 = hmaster2_p & v230446f | !hmaster2_p & v84561b;
assign v230330d = hbusreq4 & v22f37de | !hbusreq4 & v22f383c;
assign v23f23fb = hbusreq6 & v23f789c | !hbusreq6 & v23fa2ec;
assign da310f = hbusreq3_p & v23f5398 | !hbusreq3_p & v23131af;
assign v23fc993 = hbusreq3_p & v2311a34 | !hbusreq3_p & v23000a6;
assign v23f81e6 = hbusreq4_p & v23fbe05 | !hbusreq4_p & v23f3561;
assign hgrant5 = !e1bacb;
assign v22f8b12 = hbusreq6 & v23fce77 | !hbusreq6 & v230dae4;
assign v22fa080 = hbusreq6 & bad6eb | !hbusreq6 & v23fba11;
assign v23f29e9 = hbusreq6 & v23045c3 | !hbusreq6 & v84561b;
assign a39dae = hbusreq5_p & v22f2bf8 | !hbusreq5_p & v84561b;
assign v23f1032 = hmaster2_p & v23fb71a | !hmaster2_p & v23fba25;
assign v230f0d2 = hmaster0_p & v2308ef0 | !hmaster0_p & v23f7c32;
assign v23f5156 = hgrant5_p & v84561b | !hgrant5_p & v22fc712;
assign v23fc66d = hmaster2_p & v23fcb55 | !hmaster2_p & v230d3f5;
assign v2301a3f = hbusreq2_p & v22fe4bb | !hbusreq2_p & a1fbb6;
assign v9cf5cf = hmaster0_p & v23f96b0 | !hmaster0_p & v23fc92e;
assign v23fcc52 = hmaster0_p & v23f41ec | !hmaster0_p & v23fbc37;
assign v8dd9c7 = hmaster2_p & v2311810 | !hmaster2_p & v9526ac;
assign v23fc963 = hbusreq1_p & v191a86f | !hbusreq1_p & !v191a876;
assign v2305aa9 = hmaster2_p & v2306d29 | !hmaster2_p & v230320e;
assign v23f65b6 = hbusreq5_p & v2307e48 | !hbusreq5_p & v2301400;
assign v23fb4d7 = hmaster2_p & v23fc6c0 | !hmaster2_p & v22f8b01;
assign v23f1a8d = locked_p & b9d00f | !locked_p & a1fbb6;
assign v23f8e1c = hbusreq4_p & v23f6032 | !hbusreq4_p & !v230f549;
assign v23f7cba = hlock5_p & v84561b | !hlock5_p & v9052d9;
assign v23fca32 = hbusreq0_p & v2301abc | !hbusreq0_p & v84561b;
assign v23f6089 = hmaster2_p & v22f1796 | !hmaster2_p & v230ce60;
assign v23f942a = hgrant3_p & v22fc27d | !hgrant3_p & v23f004a;
assign v23015de = hgrant3_p & v2300cf1 | !hgrant3_p & v22f3be2;
assign v22f62ea = hmaster2_p & v23fb67c | !hmaster2_p & v23035ba;
assign v230c2f3 = hbusreq1_p & v22ee3a3 | !hbusreq1_p & v84561b;
assign v230833e = hbusreq3_p & v23fc19b | !hbusreq3_p & v23117f5;
assign v23fbe21 = hmaster2_p & v23f87f4 | !hmaster2_p & !v23f8490;
assign v22f4594 = hbusreq2_p & v23fc900 | !hbusreq2_p & !v23fcc28;
assign v22fd7d4 = hbusreq6 & v22f05b9 | !hbusreq6 & !v84562a;
assign v22f9f26 = hgrant1_p & v845626 | !hgrant1_p & v23f83f3;
assign v2312912 = hgrant5_p & v22fe51f | !hgrant5_p & v2303125;
assign v23118f7 = hmaster2_p & v22fbb8a | !hmaster2_p & !v2304009;
assign v23f1eb7 = hgrant3_p & v23f266b | !hgrant3_p & v2310bdf;
assign v23fca93 = hburst0_p & v230371b | !hburst0_p & v12cd995;
assign v231096b = hmaster0_p & v22fe2a8 | !hmaster0_p & v230d58c;
assign v22ed9a9 = hgrant3_p & v2306fba | !hgrant3_p & v230a644;
assign v22f516b = hlock0_p & v230c104 | !hlock0_p & v2302868;
assign v2300af8 = hbusreq5_p & v2303d2e | !hbusreq5_p & !v23fc0f0;
assign v22f0069 = hbusreq3 & v2301b00 | !hbusreq3 & v84561b;
assign v23fbc89 = hmaster1_p & v22ed631 | !hmaster1_p & !v2305b24;
assign v23fbdd4 = hbusreq0 & v22fcdf6 | !hbusreq0 & v84564d;
assign v23fbb80 = hlock0_p & v23f5043 | !hlock0_p & v23fc622;
assign v8f9141 = hbusreq6_p & v23fc39d | !hbusreq6_p & v23f34e1;
assign bd7530 = hbusreq4_p & v22f9a75 | !hbusreq4_p & v23fcab3;
assign v23fba07 = hbusreq3 & v230e618 | !hbusreq3 & v84561b;
assign v23f3c3b = hmaster2_p & v84561b | !hmaster2_p & v23f7d57;
assign v23041ea = hbusreq4_p & v22f5808 | !hbusreq4_p & v2308b58;
assign v230d56c = hbusreq5_p & v23fa2ec | !hbusreq5_p & v23fc4f8;
assign v22eba71 = hbusreq3_p & v22fc020 | !hbusreq3_p & v84561b;
assign v23f165d = hmaster0_p & v23fcdd1 | !hmaster0_p & !v230be28;
assign v23f033c = hbusreq5 & v2312f7e | !hbusreq5 & !v23022b1;
assign v2302db0 = hbusreq3_p & v230391b | !hbusreq3_p & v84561b;
assign v89e88b = hmaster2_p & v23fc094 | !hmaster2_p & v2309550;
assign v1aad441 = jx0_p & v23fa08a | !jx0_p & v22ffde1;
assign v2300ce0 = hmaster1_p & e1df52 | !hmaster1_p & v22ed8b0;
assign v23fcefd = hbusreq5_p & v230ef7c | !hbusreq5_p & v22f5d1e;
assign v9e8d9f = hbusreq1_p & v150748b | !hbusreq1_p & v22ec522;
assign v23f5e3d = hmaster0_p & v23fbdf6 | !hmaster0_p & !v2394087;
assign v22fdbd2 = hgrant3_p & v84561b | !hgrant3_p & v22ed8bc;
assign v22f7bb9 = hgrant1_p & a1fbc2 | !hgrant1_p & v23916c0;
assign v12cd692 = hmaster2_p & v231009b | !hmaster2_p & !v23027e9;
assign v1b87673 = hmastlock_p & v23fce65 | !hmastlock_p & !v84561b;
assign e1df54 = hgrant3_p & v2302251 | !hgrant3_p & v23f6927;
assign v22ee516 = hmastlock_p & v23f00cf | !hmastlock_p & !v84561b;
assign v22f0b75 = hmaster0_p & v2304bcb | !hmaster0_p & v22fe1c8;
assign v22ed337 = hlock3_p & v23f1193 | !hlock3_p & v84561b;
assign v191ac91 = hbusreq1 & v23fc658 | !hbusreq1 & v23fa397;
assign v22f2a76 = hbusreq5 & v23f3d14 | !hbusreq5 & v22ee9be;
assign v23fc925 = hgrant1_p & v845626 | !hgrant1_p & v2304691;
assign v23fcad0 = busreq_p & v22f691e | !busreq_p & ae2bc6;
assign v23fd055 = hbusreq5 & v13afe3a | !hbusreq5 & !v23fce22;
assign v2346b8a = hgrant0_p & v84561b | !hgrant0_p & v230fa1a;
assign v23f9a4d = hbusreq4_p & v23fbd62 | !hbusreq4_p & v23fb9cb;
assign v2312cb9 = hmaster0_p & v23f598e | !hmaster0_p & v22fcd80;
assign v22f654a = stateG10_5_p & v230ac29 | !stateG10_5_p & v23fc3fa;
assign afb25b = hmaster2_p & v84561b | !hmaster2_p & v23fb5d6;
assign v22f015d = hgrant1_p & v12cd9f9 | !hgrant1_p & !v23fcaf1;
assign f40aac = hbusreq2_p & v22f099c | !hbusreq2_p & v23928cd;
assign v23fc4a7 = hbusreq6_p & v84561b | !hbusreq6_p & v23f56b1;
assign v22fb3ef = hbusreq3 & v23fa2d6 | !hbusreq3 & v84561b;
assign v23121e0 = hbusreq4 & v230af06 | !hbusreq4 & v23fd015;
assign v22f45ff = hbusreq5 & v22f299f | !hbusreq5 & v84561b;
assign v23fb862 = hbusreq3_p & v22fe285 | !hbusreq3_p & v22f2254;
assign v22fb27b = hmaster2_p & v84561b | !hmaster2_p & v23fc84e;
assign v1aad420 = hbusreq4_p & v2306e6f | !hbusreq4_p & v23104cf;
assign v231242d = hmaster0_p & v13afeb1 | !hmaster0_p & !v22f8e4d;
assign v22f5f28 = hgrant3_p & v23f5fc3 | !hgrant3_p & v23f5398;
assign v22ec0d9 = hlock3_p & v23139ef | !hlock3_p & v22f7861;
assign v191ab91 = stateG10_5_p & v2303125 | !stateG10_5_p & v23f4b28;
assign v22f2d93 = hmaster1_p & v23055c3 | !hmaster1_p & v23fc840;
assign v22ecc3b = hmaster2_p & v23919f9 | !hmaster2_p & v23fca72;
assign v23f1608 = hmaster0_p & v23fc277 | !hmaster0_p & v22f3272;
assign v2312b9e = hgrant3_p & v84561b | !hgrant3_p & !v23f86a0;
assign v23fb10d = hgrant0_p & v845622 | !hgrant0_p & v22f03b8;
assign v23fb5f6 = hmaster2_p & v230e4ef | !hmaster2_p & !v23f763f;
assign v230e8a7 = hmaster0_p & v84561b | !hmaster0_p & v230753a;
assign v23f84cc = hbusreq1 & v23fca23 | !hbusreq1 & v84561b;
assign v191acbd = hbusreq3_p & v22fe44f | !hbusreq3_p & v22fa736;
assign v22fa299 = jx1_p & v22f0c5f | !jx1_p & v84561b;
assign f40a9e = hgrant5_p & v230a44c | !hgrant5_p & v22ef683;
assign v2309c45 = hbusreq3_p & d7df7e | !hbusreq3_p & v23fc4d1;
assign v23fcdc5 = hmaster2_p & v22ed85a | !hmaster2_p & v22fc34e;
assign v23fb66a = hbusreq0 & v22ff315 | !hbusreq0 & v23fb966;
assign v23fb81d = hbusreq3_p & v2307320 | !hbusreq3_p & v84561b;
assign v23fcca2 = jx0_p & v2302f12 | !jx0_p & v23fc638;
assign v22ef35b = jx1_p & e1e34d | !jx1_p & v22f0c75;
assign v2303e06 = hlock5_p & v13aff30 | !hlock5_p & v230d379;
assign v22edf29 = hbusreq6 & v22f2e75 | !hbusreq6 & v23fc5be;
assign v23059ee = hbusreq3 & v23fc176 | !hbusreq3 & v84561b;
assign v23fca66 = hmaster2_p & v23127ff | !hmaster2_p & v23fb624;
assign v23f51a6 = jx1_p & v22ee0c9 | !jx1_p & v23fc5ce;
assign v239174c = hlock1_p & v23fb590 | !hlock1_p & v230840f;
assign v22fd5dd = hbusreq0_p & v106ae19 | !hbusreq0_p & b9d013;
assign v22fd30c = hgrant2_p & v2306d29 | !hgrant2_p & !v191a86f;
assign v1507557 = hbusreq4 & v23fc68a | !hbusreq4 & v23fbf27;
assign v23f78a3 = hbusreq6 & v22ebfcb | !hbusreq6 & v230da9b;
assign v1aae294 = hmastlock_p & v23fcb89 | !hmastlock_p & v84561b;
assign v230377f = hbusreq0_p & v23f6411 | !hbusreq0_p & !v106ae19;
assign v23f52b9 = hmaster0_p & v22f2e69 | !hmaster0_p & v2310ec8;
assign v23fc9c1 = hgrant2_p & v84562a | !hgrant2_p & !v919ce6;
assign v23fb808 = hbusreq4_p & v22eb38b | !hbusreq4_p & v22f451b;
assign v23fc953 = hmaster2_p & v22ffe8d | !hmaster2_p & v23fba9a;
assign v230158f = hbusreq0_p & v84561b | !hbusreq0_p & v1aae087;
assign v22f4828 = hbusreq6_p & v23fc887 | !hbusreq6_p & v2310747;
assign v22f3411 = hmaster2_p & v22fd0e6 | !hmaster2_p & v230971e;
assign v23fbae8 = hbusreq1 & v1aad5ad | !hbusreq1 & v22eefab;
assign v22fe7f5 = hgrant0_p & v22f5605 | !hgrant0_p & !v23fb215;
assign v2307fb2 = hmaster1_p & v23fbf13 | !hmaster1_p & v231188f;
assign v23fc864 = hmaster2_p & v23facc2 | !hmaster2_p & !v23fb796;
assign v23f5eba = hmaster2_p & v84561b | !hmaster2_p & !v22f1e02;
assign v23fbdf5 = hbusreq6 & v230cae4 | !hbusreq6 & v2302c91;
assign v22ee345 = hbusreq6 & v22ebb85 | !hbusreq6 & !v2312ea0;
assign v23f8d91 = hbusreq4_p & v22f59bd | !hbusreq4_p & v22ec1b1;
assign v22f6a6b = hgrant2_p & v23126ae | !hgrant2_p & v191a876;
assign v230cb53 = hmaster0_p & v23fb083 | !hmaster0_p & v22f0698;
assign v23fb9a9 = hgrant1_p & v84561b | !hgrant1_p & v23f111c;
assign v23fbe30 = hgrant3_p & v22f2db6 | !hgrant3_p & !v2303154;
assign v899296 = hbusreq1_p & v2300b6b | !hbusreq1_p & v845620;
assign v230e8a6 = hgrant1_p & v22fe426 | !hgrant1_p & v23f5bf3;
assign v23f97a7 = hmaster2_p & v2308880 | !hmaster2_p & v22fc80c;
assign v2303115 = hmaster2_p & v230f34c | !hmaster2_p & !v23035ba;
assign v22f9911 = locked_p & v22f7f52 | !locked_p & v191a86f;
assign v230a9f0 = hgrant0_p & v230aded | !hgrant0_p & v1aadb95;
assign v23f5109 = hmaster1_p & v84561b | !hmaster1_p & v22f6e51;
assign v22f9d69 = hbusreq0 & v106ae21 | !hbusreq0 & v84564d;
assign v22f4858 = hbusreq3_p & v22f0069 | !hbusreq3_p & v84561b;
assign v22f4593 = hbusreq1_p & v23fb6c6 | !hbusreq1_p & a1fe3e;
assign v22fec16 = hgrant4_p & v23fc1ac | !hgrant4_p & v23f4f3b;
assign v23f2b21 = hmaster2_p & v23fbb5f | !hmaster2_p & v23035d7;
assign v230e6ee = hready & v23fbc8c | !hready & !v84561b;
assign v2305f8e = hmaster2_p & v2306b2e | !hmaster2_p & v22f03cf;
assign v23f1c9b = hlock3_p & v23efce3 | !hlock3_p & !v84561b;
assign v22ff64f = stateA1_p & v84561b | !stateA1_p & v230cfe2;
assign v22eede3 = hbusreq4 & v23f98d4 | !hbusreq4 & v23fb102;
assign v23f7123 = hlock1_p & v22f8cb7 | !hlock1_p & !v84561b;
assign v22f181c = hbusreq0_p & v2391aa0 | !hbusreq0_p & v23fd040;
assign v23fc19d = hgrant0_p & v22f824f | !hgrant0_p & v23f7218;
assign v23fc194 = hmaster2_p & v22f7b29 | !hmaster2_p & v23fb9cf;
assign v2303e4f = hmaster2_p & v2312775 | !hmaster2_p & v84561b;
assign v23f8a70 = hmaster2_p & v2312259 | !hmaster2_p & !v84561b;
assign v2391d40 = hbusreq0 & v2306220 | !hbusreq0 & !v84561b;
assign v23f6a11 = hlock5_p & v22ff89d | !hlock5_p & !v230330a;
assign v22f8ce6 = hmaster0_p & v22f50f0 | !hmaster0_p & v22f165f;
assign v23fbeb5 = hmaster2_p & v2391f2b | !hmaster2_p & v84561b;
assign v23fbf26 = hbusreq2_p & v22f1b11 | !hbusreq2_p & v845620;
assign v23fcf81 = hbusreq4 & v22ed684 | !hbusreq4 & v22f3839;
assign v23123a3 = jx3_p & v2305141 | !jx3_p & v230754e;
assign v23007c9 = hgrant3_p & v23f9b49 | !hgrant3_p & v22ec934;
assign v23f87e1 = hgrant3_p & v22f3643 | !hgrant3_p & v23f6089;
assign v23f8689 = hgrant3_p & v23fc457 | !hgrant3_p & v23f5abd;
assign v22fdbac = hbusreq6_p & v23f2dbb | !hbusreq6_p & v23fb8b7;
assign v22eb899 = hbusreq3_p & v230ccc4 | !hbusreq3_p & v22fb0cb;
assign v23fb98a = hgrant1_p & v84561b | !hgrant1_p & v23f51a4;
assign v23f8dba = hbusreq4_p & v22ff789 | !hbusreq4_p & v84562b;
assign v22ee269 = hbusreq5_p & v22ebe7f | !hbusreq5_p & v23f23e8;
assign v230e779 = hmaster0_p & v22ef575 | !hmaster0_p & v23fd035;
assign v23fccd8 = hmaster2_p & v230ea6d | !hmaster2_p & v23f63ab;
assign v230fe14 = hmaster0_p & v230ad15 | !hmaster0_p & v22f8b12;
assign v23108db = hbusreq3 & v23117c1 | !hbusreq3 & v84561b;
assign v22fd9eb = hbusreq1 & bd7476 | !hbusreq1 & !v230af81;
assign v22f1403 = hgrant5_p & v2303943 | !hgrant5_p & v23fc997;
assign v230ae09 = hbusreq1 & v85d110 | !hbusreq1 & v84561b;
assign v22f8f64 = hmaster0_p & v23fca6c | !hmaster0_p & v2304332;
assign v23fd026 = hmaster0_p & v22f0dc9 | !hmaster0_p & v2306625;
assign v22fd720 = stateG10_5_p & v23fc9b9 | !stateG10_5_p & !v84561b;
assign v2305c7f = hbusreq4_p & v2310589 | !hbusreq4_p & v2309c93;
assign v230f9e8 = hgrant5_p & v84561b | !hgrant5_p & v22fd0cd;
assign v22ee8bf = hgrant3_p & v23fce1e | !hgrant3_p & v22fa889;
assign v2309eb8 = hmaster2_p & v13afe8f | !hmaster2_p & !v231228e;
assign v23f75ce = hbusreq1_p & v23f595d | !hbusreq1_p & !v106ae19;
assign v23f6470 = hmaster2_p & v22ebdbc | !hmaster2_p & v2304922;
assign v23f3e1b = hlock3_p & v23f15a7 | !hlock3_p & !v22fecf3;
assign v2306b06 = hbusreq4_p & v22ed928 | !hbusreq4_p & a296f8;
assign v22f03b1 = hbusreq3 & v23f93e7 | !hbusreq3 & v2310d04;
assign v2392f21 = stateG10_5_p & v23084cf | !stateG10_5_p & v22ec801;
assign v22ef424 = hbusreq1_p & v23f3940 | !hbusreq1_p & v22f7e37;
assign v22f85f6 = hmaster1_p & v22f1afb | !hmaster1_p & v23fd00e;
assign v22ec745 = hbusreq5_p & ab4e4e | !hbusreq5_p & !v84561b;
assign v23fc030 = hbusreq3 & v23fbdb9 | !hbusreq3 & v84561b;
assign v230463a = hmaster2_p & v23fc755 | !hmaster2_p & !v84561b;
assign v22ec4ce = hgrant5_p & a3ace7 | !hgrant5_p & v2302075;
assign v2304744 = hmaster1_p & v22f6917 | !hmaster1_p & !v17a34ff;
assign v22efd99 = hmaster1_p & v22fe6f8 | !hmaster1_p & v22efadc;
assign v23928f2 = hmaster0_p & v23fbc7e | !hmaster0_p & v22ed907;
assign v230be28 = hgrant3_p & v2300362 | !hgrant3_p & v22fd150;
assign v230e04a = hmaster0_p & v230d6ca | !hmaster0_p & v23fc7e3;
assign v230e8b8 = stateA1_p & v23fc116 | !stateA1_p & v22f3294;
assign v23f9dba = hbusreq4_p & v23f4015 | !hbusreq4_p & v23f8a89;
assign v23f3f59 = hmaster2_p & v22f1244 | !hmaster2_p & v230e3a0;
assign v22eb184 = hbusreq6 & v22f6844 | !hbusreq6 & v23f87f4;
assign v22f61d2 = hmaster2_p & v23f646e | !hmaster2_p & v2310e40;
assign v22f63cc = hmaster0_p & v84561b | !hmaster0_p & v23f77d5;
assign v22f98e3 = hlock0_p & v22ef509 | !hlock0_p & v845622;
assign v239367b = hbusreq5_p & v84561b | !hbusreq5_p & !v2311268;
assign v8d83bb = hmaster2_p & v22f1244 | !hmaster2_p & v23fc1df;
assign v84562a = hbusreq2 & v84561b | !hbusreq2 & !v84561b;
assign v23f4fa4 = hbusreq3_p & v22f05b9 | !hbusreq3_p & v23fce3a;
assign v23faa19 = hmaster2_p & v22f7ab4 | !hmaster2_p & v23fa69c;
assign v2311d9d = hbusreq5 & v22f343b | !hbusreq5 & !v84562a;
assign f406c6 = hbusreq1_p & v23f5cb3 | !hbusreq1_p & !v2310e40;
assign v8d030a = hlock0_p & v2391d40 | !hlock0_p & v84561b;
assign v2391a57 = locked_p & f4067f | !locked_p & v84561b;
assign v22f19c3 = hready_p & v84564d | !hready_p & v22ed42c;
assign v22ffdc3 = hbusreq6_p & v22f9dab | !hbusreq6_p & v13afef6;
assign v8abd93 = hgrant1_p & v84561b | !hgrant1_p & v2306bf9;
assign v22ed309 = hgrant3_p & v84561b | !hgrant3_p & v23fc387;
assign v23f83ff = hbusreq5_p & v84561b | !hbusreq5_p & !v23fcb35;
assign v230b3ec = hbusreq3_p & v22f128d | !hbusreq3_p & !v230f691;
assign v23f73a4 = hbusreq2_p & v23fc5ec | !hbusreq2_p & v230766b;
assign v23f8e25 = hbusreq3_p & c60af7 | !hbusreq3_p & v84561b;
assign v22f174d = hlock3_p & v230bb2d | !hlock3_p & !v23fc5eb;
assign v2393f95 = hmaster2_p & v22eec6e | !hmaster2_p & v230ce60;
assign v23fc454 = hgrant0_p & v84561b | !hgrant0_p & v22ec6d9;
assign v23fb958 = hbusreq3_p & v230e040 | !hbusreq3_p & v23fc957;
assign v23f5ba9 = hlock3_p & v2312b5a | !hlock3_p & !v23fcb68;
assign v22fc70a = hmaster2_p & v845620 | !hmaster2_p & v23fcfbe;
assign v22f8864 = hmaster0_p & v23fbcfd | !hmaster0_p & v2393635;
assign v23fcb23 = hlock0_p & v84561b | !hlock0_p & v23f999c;
assign v23f5102 = hbusreq1 & v150736d | !hbusreq1 & v84561b;
assign v2392ed3 = stateG10_5_p & v23f529c | !stateG10_5_p & v2392534;
assign v23fc96d = hbusreq3 & v191aed3 | !hbusreq3 & v84564d;
assign v239214a = hmaster2_p & v22ee9be | !hmaster2_p & v23f3d14;
assign v22eee95 = hbusreq6 & v2310385 | !hbusreq6 & v22fbd4f;
assign v22f6607 = hgrant5_p & v23fcea9 | !hgrant5_p & !v22f6a93;
assign v23fa9df = hgrant5_p & v22ee561 | !hgrant5_p & v22f1dab;
assign v2304c77 = hgrant1_p & v2303147 | !hgrant1_p & v22f291f;
assign v23efc12 = hbusreq5_p & v23fc945 | !hbusreq5_p & !v84561b;
assign v23125ab = hmaster0_p & v23fb045 | !hmaster0_p & v22f7fed;
assign v2393364 = hlock0_p & v2308a42 | !hlock0_p & v2300597;
assign v230cbc4 = hlock3_p & v22f52d4 | !hlock3_p & v22fe2ae;
assign v2309cda = jx1_p & v23f651e | !jx1_p & v23fbb63;
assign v23f9fc8 = hmaster0_p & v23f1e38 | !hmaster0_p & v22fce2e;
assign v230d921 = hbusreq1_p & v22ed495 | !hbusreq1_p & v23fc8d2;
assign v23fc80c = hmaster0_p & v23f5046 | !hmaster0_p & v230aedf;
assign v23f7db8 = hbusreq1 & v23f5043 | !hbusreq1 & v84561b;
assign v22ef26f = hmaster2_p & v2305fe0 | !hmaster2_p & !v84561b;
assign v191b085 = hbusreq4_p & v230e8ea | !hbusreq4_p & v23f51ac;
assign v23f6c83 = hmaster0_p & v22fcdd3 | !hmaster0_p & v2304904;
assign v23fc526 = hbusreq5 & v22feb47 | !hbusreq5 & v84561b;
assign v2312067 = hbusreq0 & v23fc4a5 | !hbusreq0 & v22f0add;
assign v23fb5ad = hbusreq0 & v22f2db0 | !hbusreq0 & v23fa2ec;
assign v23fbc65 = hmaster0_p & v230e43d | !hmaster0_p & v230abf6;
assign v230697e = hmaster2_p & v106a81a | !hmaster2_p & a1fbb6;
assign v23fbea6 = hmaster2_p & v23f78a4 | !hmaster2_p & v23fb2f7;
assign v230d25d = hbusreq6 & v2391d2f | !hbusreq6 & v230ef09;
assign v191a905 = hmaster0_p & v23fcdf6 | !hmaster0_p & !v96c563;
assign v23f6729 = hgrant1_p & v12cd6a1 | !hgrant1_p & v23fca90;
assign v230d24a = hbusreq0_p & v191a86f | !hbusreq0_p & !v22f9980;
assign v23fc748 = hmaster2_p & v23fcbd7 | !hmaster2_p & v84561b;
assign v23f680a = hbusreq2 & v22f7f74 | !hbusreq2 & v84561b;
assign v2391b46 = hgrant1_p & v84561b | !hgrant1_p & v23fce11;
assign v23fc357 = hgrant3_p & v22f368e | !hgrant3_p & v23fbcd0;
assign v2303c5a = hgrant3_p & v84562d | !hgrant3_p & v230064b;
assign v23fbb6a = hlock0_p & v84561b | !hlock0_p & v2302e80;
assign v22f1d85 = hbusreq4_p & v23f1e5c | !hbusreq4_p & v23fb43a;
assign v23042ca = hmaster0_p & v231363b | !hmaster0_p & v22f24a3;
assign v23fc275 = hmaster2_p & v22ee703 | !hmaster2_p & v23fba9a;
assign v22f9a8b = hmaster0_p & v23fc804 | !hmaster0_p & !v23f0206;
assign v23fc788 = hbusreq5_p & v22fa594 | !hbusreq5_p & !v23fce8b;
assign v22fee58 = hlock3_p & v23033d3 | !hlock3_p & v23fb0f0;
assign v23055f4 = hlock3_p & v23f90b2 | !hlock3_p & v23f53a0;
assign bd7f18 = hmaster2_p & a1f77b | !hmaster2_p & !v2308110;
assign v22f9321 = hbusreq1_p & v22feb0d | !hbusreq1_p & v23f8241;
assign v22f1f55 = hbusreq6_p & v2309b63 | !hbusreq6_p & v1b87776;
assign v230477b = jx1_p & v23f8180 | !jx1_p & v230deb1;
assign v23fcba5 = hgrant5_p & v23f49b3 | !hgrant5_p & v22f6058;
assign v22fe4f6 = hmaster0_p & v2308d9e | !hmaster0_p & !v2303fec;
assign v22f74de = hgrant5_p & v84561b | !hgrant5_p & !v2300059;
assign v22f639d = hbusreq4_p & v230b77e | !hbusreq4_p & fc8c53;
assign v23fc20e = hbusreq3_p & b9d00f | !hbusreq3_p & v23fcebf;
assign v22f7e4a = hbusreq5_p & v2392a17 | !hbusreq5_p & !v22faee9;
assign v23fbca3 = hbusreq5_p & v22eb5b3 | !hbusreq5_p & v23fcc36;
assign v2303fb2 = hmaster2_p & v1aae56f | !hmaster2_p & v2307150;
assign v2308a30 = locked_p & v106ae4a | !locked_p & !v2309c8a;
assign v231350d = hbusreq1_p & v2310303 | !hbusreq1_p & !v230f848;
assign v23fbd56 = hmaster2_p & v23fc393 | !hmaster2_p & !v22fdc30;
assign v22ece29 = hbusreq4 & v2304b8d | !hbusreq4 & v84561b;
assign v2301800 = hgrant3_p & v2308364 | !hgrant3_p & v23f7024;
assign v22f2883 = hbusreq1_p & v23130ac | !hbusreq1_p & !v2307a62;
assign v22eef44 = hbusreq3_p & v22ef750 | !hbusreq3_p & v23fbf35;
assign v22f2271 = hgrant2_p & v22fee46 | !hgrant2_p & a1fbb6;
assign b59af9 = hmaster0_p & v23928ae | !hmaster0_p & v23f0eec;
assign v23fc811 = stateG10_5_p & v23f301a | !stateG10_5_p & v22faa21;
assign v230e534 = hmaster1_p & v22fa39e | !hmaster1_p & v23f2f40;
assign v23fb9b9 = hlock2_p & v84561b | !hlock2_p & !v1aae362;
assign v22f9d57 = hmaster1_p & v23fca34 | !hmaster1_p & v84561b;
assign v2308750 = hmaster2_p & v2310e40 | !hmaster2_p & v22fe426;
assign v22f0492 = hmaster2_p & v22ef513 | !hmaster2_p & v2310bdf;
assign v230a9a3 = hbusreq3_p & v22fba41 | !hbusreq3_p & v23f4b28;
assign v22f58f9 = hbusreq5 & v9585ce | !hbusreq5 & !v2392fa3;
assign v23039ea = hmaster0_p & v230ed3d | !hmaster0_p & v23fc301;
assign v22fd6ba = hbusreq5 & v2312ea7 | !hbusreq5 & v84561b;
assign v23fce4d = jx0_p & v23fccb8 | !jx0_p & !v23f623e;
assign v23fc498 = hbusreq3 & v2303fe4 | !hbusreq3 & v84561b;
assign v23f6a00 = hgrant3_p & v1e84072 | !hgrant3_p & v22ee184;
assign v22fd973 = hbusreq5_p & v22fb95e | !hbusreq5_p & v23f67bd;
assign v23fb2ba = hbusreq3_p & v230d14d | !hbusreq3_p & v12cd673;
assign v2309130 = hmaster2_p & v2313131 | !hmaster2_p & v22f766b;
assign v903f7f = hmaster2_p & v23fceb9 | !hmaster2_p & v1aad5ad;
assign v230f34c = hbusreq0_p & v2307707 | !hbusreq0_p & !v84561b;
assign v1aad4c6 = hmaster2_p & v191a86f | !hmaster2_p & v2302e32;
assign v22f8603 = hbusreq0 & v230d5f4 | !hbusreq0 & v23f0eeb;
assign v22fd621 = hmaster2_p & v23fb54f | !hmaster2_p & v22fbe6a;
assign v23080be = hmaster1_p & v22f457a | !hmaster1_p & !v23f49cd;
assign v23f86a0 = hbusreq3_p & v22fe920 | !hbusreq3_p & v23f052e;
assign v23129e0 = hgrant1_p & v22ec477 | !hgrant1_p & v231343f;
assign v22fd283 = hgrant1_p & e1df2d | !hgrant1_p & v84561b;
assign v22fdb73 = hbusreq4_p & af5f08 | !hbusreq4_p & v23fbc6e;
assign v22ff0d3 = hgrant3_p & v23f558b | !hgrant3_p & v22f482a;
assign v23126de = hlock1_p & v23f5102 | !hlock1_p & v23063f8;
assign v22f2a60 = hgrant5_p & v23f71d5 | !hgrant5_p & v22f7b13;
assign bd7ae5 = hbusreq6 & v84564d | !hbusreq6 & v84561b;
assign a37ffd = hbusreq1_p & v2309c55 | !hbusreq1_p & v22f7241;
assign v23fcb40 = hgrant3_p & v23fc975 | !hgrant3_p & v230f5b9;
assign v22eed66 = hgrant2_p & a1fbc2 | !hgrant2_p & a1fbb6;
assign v23f8928 = hgrant1_p & v2303068 | !hgrant1_p & v23fba24;
assign v2301933 = hbusreq2 & v84561b | !hbusreq2 & v23f5043;
assign v23fcb2d = hlock3_p & v22fc95b | !hlock3_p & v23fce8e;
assign v22fe852 = hbusreq3 & v2305024 | !hbusreq3 & v84561b;
assign v13afaae = hbusreq5_p & v23035ba | !hbusreq5_p & v231192e;
assign v1506eb2 = hmaster0_p & v2308815 | !hmaster0_p & v230f08b;
assign v23103e6 = hmaster0_p & v2302094 | !hmaster0_p & v23055c3;
assign v22fb4ab = hmaster2_p & v2304283 | !hmaster2_p & v23101b1;
assign e1e258 = hbusreq3_p & v1aad46b | !hbusreq3_p & v23f8ddb;
assign v22f3e14 = hbusreq1 & v23f2be7 | !hbusreq1 & v84561b;
assign v2301e4f = hmaster0_p & v22ff6c5 | !hmaster0_p & v23fc4c3;
assign v23fca31 = hmaster0_p & v84561b | !hmaster0_p & !v23f8c1f;
assign v23065b6 = hlock1_p & v23fc6d3 | !hlock1_p & v84564d;
assign v22f4cf2 = hgrant4_p & v22fee59 | !hgrant4_p & v23f4bab;
assign v230ad0f = hgrant3_p & v23fbe2d | !hgrant3_p & v106ae87;
assign v22f6bae = hgrant3_p & v22ffa6e | !hgrant3_p & v22f6894;
assign v23fb60a = hmaster2_p & b9d00f | !hmaster2_p & a1fbb6;
assign v23f5872 = hbusreq2 & bd8382 | !hbusreq2 & v84561b;
assign v22f215c = hlock0_p & v23f5cb3 | !hlock0_p & v2312e03;
assign v22f3ac3 = hgrant3_p & v15071c7 | !hgrant3_p & v97ba8e;
assign v22ed809 = hbusreq3 & v2307f2b | !hbusreq3 & !v845622;
assign v230e9ea = hgrant2_p & v22f753f | !hgrant2_p & v845620;
assign v2306703 = hgrant3_p & v2308dd1 | !hgrant3_p & v23fc098;
assign v22f5db6 = hbusreq5_p & v2306d29 | !hbusreq5_p & v22fdc30;
assign v230389f = hgrant3_p & v23f6283 | !hgrant3_p & v22f2114;
assign v23fb9c1 = hmaster0_p & v22f7ee5 | !hmaster0_p & v22ec350;
assign v230e07e = hbusreq5_p & v23f529c | !hbusreq5_p & v23fb4b1;
assign v22fafe4 = hbusreq2_p & v23fb71f | !hbusreq2_p & !v23f8914;
assign v106a7d3 = hbusreq4_p & v2307170 | !hbusreq4_p & v22ec8dc;
assign v22f25da = hmaster2_p & v23fb5a1 | !hmaster2_p & v22f7b47;
assign v23f8100 = hmaster0_p & v23f20d0 | !hmaster0_p & v230562d;
assign v23fbc5a = hlock5_p & v84561b | !hlock5_p & v23fcd16;
assign a9da2d = hmaster2_p & v23f1a1c | !hmaster2_p & !v22f1d80;
assign v22f2d83 = stateA1_p & v2302ca3 | !stateA1_p & v23fb98d;
assign v2312e03 = hbusreq0_p & v23fbfb9 | !hbusreq0_p & !v22fd25c;
assign v22f8cd8 = hlock0_p & v106ae4a | !hlock0_p & v23f084d;
assign v22eea15 = jx1_p & v22f2d93 | !jx1_p & v2309410;
assign a1ba8b = hbusreq4 & v23f5055 | !hbusreq4 & v84561b;
assign v22ffffa = jx1_p & v23fcdb1 | !jx1_p & v23efe7d;
assign v22fd60f = jx0_p & v2307403 | !jx0_p & !v2305630;
assign a33e98 = hlock5_p & v23fc468 | !hlock5_p & v1b87690;
assign v23f3dd7 = hmaster0_p & v230b781 | !hmaster0_p & f4061f;
assign v22f5137 = hbusreq5_p & v1e845ac | !hbusreq5_p & v13afe7d;
assign v230a66b = hbusreq3 & v22fa262 | !hbusreq3 & !v23f7c8d;
assign f40c98 = hgrant3_p & v23f6635 | !hgrant3_p & v23fcb71;
assign v22f071b = hgrant1_p & v22ee73b | !hgrant1_p & !v23f5622;
assign v2312164 = hlock4_p & v23fc72c | !hlock4_p & v23f507b;
assign v2312007 = hgrant3_p & v84561b | !hgrant3_p & v106aeed;
assign v22fb155 = hgrant5_p & v23fbe4d | !hgrant5_p & !v2305050;
assign v2306d2c = hlock4_p & v2300cd4 | !hlock4_p & v23f347b;
assign v230af3a = hbusreq0 & v23fc926 | !hbusreq0 & v2308848;
assign v23fcf8f = hgrant2_p & a07f9b | !hgrant2_p & v23f15fe;
assign v23112d5 = hbusreq5_p & v22fe0c1 | !hbusreq5_p & v84561b;
assign v23fc3ac = hmaster0_p & v22f31b9 | !hmaster0_p & b95000;
assign v150716b = hbusreq6_p & v1aad354 | !hbusreq6_p & v230f0c6;
assign v22f80b4 = hbusreq1_p & v9526ac | !hbusreq1_p & v23fb1c6;
assign v23f946b = hmaster2_p & v84561b | !hmaster2_p & !v22f4114;
assign v2304919 = hbusreq3_p & v23fb925 | !hbusreq3_p & v23f4ce2;
assign v22efb77 = hbusreq1_p & v23f4b28 | !hbusreq1_p & v23035ba;
assign v2310db9 = hmaster0_p & e1e358 | !hmaster0_p & !v96c563;
assign v22f6ac9 = hgrant5_p & v22f53b4 | !hgrant5_p & v23f36a5;
assign v23f0978 = hbusreq6 & ae0418 | !hbusreq6 & v84561b;
assign v22f349a = stateA1_p & v84561b | !stateA1_p & !v23fbeb4;
assign v23fa599 = hbusreq4_p & v22f6e51 | !hbusreq4_p & v23fc296;
assign bd770f = jx3_p & v23fc5b7 | !jx3_p & v2307c06;
assign v23fc0d4 = hmaster0_p & v23fb7c3 | !hmaster0_p & !v23fcc3d;
assign v2306996 = hmaster2_p & v84561b | !hmaster2_p & v2391bc1;
assign v23fbaed = hbusreq4 & v2310d2f | !hbusreq4 & v84561b;
assign v22f5280 = locked_p & v9526ac | !locked_p & a1fba6;
assign v23fc59a = hbusreq1_p & v22f0de9 | !hbusreq1_p & !b9d013;
assign v230a3e6 = hmaster2_p & v23fba93 | !hmaster2_p & !v84561b;
assign v23fc26f = hgrant5_p & v23f5caf | !hgrant5_p & v23f7031;
assign v23fc53d = hlock6_p & v2306126 | !hlock6_p & v84561b;
assign v191ae42 = hbusreq2_p & v191a86f | !hbusreq2_p & !v13afe8f;
assign v239345a = hbusreq6_p & v23fb9c4 | !hbusreq6_p & v23fc0bf;
assign v22ec1fc = hmaster0_p & v230f18c | !hmaster0_p & v23fcaf6;
assign v22f383e = stateG10_5_p & v22f4d46 | !stateG10_5_p & v22f0824;
assign v22f21d0 = hmaster0_p & v23f525c | !hmaster0_p & v22f092c;
assign v99ce01 = hlock3_p & v2311c26 | !hlock3_p & v22f732c;
assign v12cd673 = hmaster2_p & v22ed6c5 | !hmaster2_p & v13affaa;
assign v23f1160 = hgrant3_p & v84561b | !hgrant3_p & v22ef0b4;
assign v22fc90f = hbusreq1_p & v230fb9e | !hbusreq1_p & !v84561b;
assign v22ec7e8 = hbusreq4 & v22ee0d6 | !hbusreq4 & v2312f81;
assign v230e7d2 = hbusreq6_p & v23fbe38 | !hbusreq6_p & v23fc006;
assign v2391950 = hlock0_p & v84561b | !hlock0_p & !v22f2590;
assign v23fc8be = busreq_p & v22ee516 | !busreq_p & !v22fdb4e;
assign v230547a = hmaster2_p & v84561b | !hmaster2_p & !v23f9127;
assign v230283f = hbusreq2_p & v22ecfe0 | !hbusreq2_p & !v84562a;
assign v23fbf13 = hbusreq6_p & v84561b | !hbusreq6_p & v22f867e;
assign v86c778 = hbusreq3 & v22efd4d | !hbusreq3 & v23fc404;
assign v230e3d1 = jx0_p & v23056b2 | !jx0_p & v23f3499;
assign v22fb00d = hlock0_p & c16191 | !hlock0_p & v23f6926;
assign v22f1d08 = hmaster0_p & v22f1ae9 | !hmaster0_p & b9d038;
assign v23fc5d5 = hready & v2302136 | !hready & !v84561b;
assign v23f6bf0 = hgrant0_p & v23f0030 | !hgrant0_p & v2308be5;
assign v23fcea5 = hbusreq4_p & v23072f3 | !hbusreq4_p & v2304e28;
assign v230b4c5 = hgrant3_p & v23fc139 | !hgrant3_p & !v23fbd69;
assign v22fc03b = hgrant0_p & v84561b | !hgrant0_p & v22f380e;
assign v22f06ac = hgrant5_p & v84561b | !hgrant5_p & v2302ea0;
assign v22ecf6c = hbusreq3 & v230b7f4 | !hbusreq3 & v22eddd9;
assign v2309cb0 = hlock1_p & v22fd372 | !hlock1_p & v23095b3;
assign v22faba5 = hmaster2_p & b9d013 | !hmaster2_p & !v230a9eb;
assign v23fc7fb = hlock0_p & v106af4d | !hlock0_p & v22ff6e8;
assign v23f3ac8 = jx1_p & v23104c1 | !jx1_p & v84561b;
assign v23035b0 = hgrant3_p & v84561b | !hgrant3_p & v22f891a;
assign v22ff4af = hbusreq3_p & v23f44bd | !hbusreq3_p & v22f21bd;
assign v2392067 = hmaster2_p & b9d00f | !hmaster2_p & v230ceb6;
assign v23fc064 = hlock1_p & v22fc42e | !hlock1_p & v230e872;
assign v23fc327 = hgrant3_p & v22fed78 | !hgrant3_p & v2310ab6;
assign v22f8d2f = hmaster1_p & v23fc140 | !hmaster1_p & v22fb790;
assign v22f15b7 = hgrant1_p & v84561b | !hgrant1_p & v2393501;
assign v2391982 = hbusreq5_p & v84561b | !hbusreq5_p & v22fa002;
assign v2312577 = hgrant5_p & v22ebc3c | !hgrant5_p & v23fba61;
assign v23f5c03 = hgrant4_p & v84561b | !hgrant4_p & v23fb8de;
assign v23f1db4 = hbusreq1_p & v23fba49 | !hbusreq1_p & v1aae9b5;
assign v231025b = hgrant1_p & v845626 | !hgrant1_p & v22fbb54;
assign v22ef079 = hbusreq6 & v12cda11 | !hbusreq6 & v845627;
assign v23fcb7e = hmaster2_p & v23fd050 | !hmaster2_p & v84561b;
assign v230ea7f = hbusreq5_p & v23f7cba | !hbusreq5_p & v84561b;
assign v2309943 = hgrant5_p & v23fb0dd | !hgrant5_p & v22ef4ce;
assign v231131d = hbusreq4_p & v230174f | !hbusreq4_p & v23f4937;
assign v23fc60a = hbusreq3 & v2312dd2 | !hbusreq3 & v84561b;
assign v23fb819 = hbusreq4_p & v23f06a5 | !hbusreq4_p & v22fff2d;
assign v23fb5db = hgrant1_p & v23fcc24 | !hgrant1_p & v23fbddb;
assign v191a86f = hmastlock_p & v230bf69 | !hmastlock_p & v84565f;
assign v23f82e4 = hbusreq3_p & v23fb115 | !hbusreq3_p & v23fc8b2;
assign v22ee7e0 = hbusreq5_p & v2313463 | !hbusreq5_p & !v23fb540;
assign v22f758c = hmaster0_p & v23fb82a | !hmaster0_p & v230abb0;
assign v22f7fd1 = hbusreq6_p & v230c12c | !hbusreq6_p & v23f710d;
assign v2300032 = hbusreq0_p & v22fef4f | !hbusreq0_p & v23f6a8a;
assign v23fc4d4 = hmaster0_p & v23fbdf6 | !hmaster0_p & !v1aad535;
assign v2311771 = hgrant4_p & v845632 | !hgrant4_p & v22fe605;
assign v22f9d07 = hbusreq6_p & v23013b5 | !hbusreq6_p & v22ed34b;
assign v22f5dc1 = hbusreq6_p & v23fcb02 | !hbusreq6_p & v23fbcbe;
assign v23fc867 = hbusreq3 & v22faa66 | !hbusreq3 & v84561b;
assign v23038ea = hmaster0_p & v23107f0 | !hmaster0_p & v22eccfc;
assign v23fbdc0 = hbusreq3 & v230153c | !hbusreq3 & v23079bc;
assign v2307375 = hbusreq1_p & v8f8537 | !hbusreq1_p & b7427f;
assign a92d05 = hbusreq0_p & v22ebee0 | !hbusreq0_p & v84562a;
assign v22f580c = hmaster0_p & v22ec354 | !hmaster0_p & !v23117c1;
assign v23fbee6 = stateG10_5_p & v23fb82c | !stateG10_5_p & v23f8e93;
assign v22eb134 = hmaster0_p & v23fc223 | !hmaster0_p & v84561b;
assign v23106ba = hgrant3_p & v22f8e29 | !hgrant3_p & v231101b;
assign v22f021c = hlock0_p & v23f646e | !hlock0_p & !v10dbf64;
assign v1b87752 = hgrant3_p & v84561b | !hgrant3_p & v23030ae;
assign v23055b0 = hmaster1_p & v84561b | !hmaster1_p & v22f52a0;
assign v23916b5 = hbusreq6 & v23f5513 | !hbusreq6 & !v23f82bb;
assign v23f3a55 = hgrant2_p & v22f8959 | !hgrant2_p & v1aae56f;
assign v23f0386 = stateG10_5_p & v23fcfcc | !stateG10_5_p & v23035ba;
assign v230ae24 = hbusreq0 & v23fbfd0 | !hbusreq0 & v23fce71;
assign v23fcb76 = hbusreq0 & v23fbdb0 | !hbusreq0 & v84561b;
assign v23fcb03 = jx1_p & v23fc8cf | !jx1_p & v84561b;
assign v230a2c6 = hlock3_p & v22ef9db | !hlock3_p & !v2304b49;
assign v230d2c2 = hbusreq1_p & v230cfe6 | !hbusreq1_p & v84561b;
assign v2300815 = hgrant1_p & v84561b | !hgrant1_p & v230de93;
assign v230913d = hbusreq2_p & v13afe3a | !hbusreq2_p & v845647;
assign v23023b3 = stateA1_p & v84561b | !stateA1_p & v23fb98d;
assign v23fc459 = hlock4_p & v23f8100 | !hlock4_p & v22eb01f;
assign v230bb9f = hbusreq6 & v23fbcad | !hbusreq6 & !v230c15a;
assign v23f733f = hbusreq3_p & v23fcecb | !hbusreq3_p & !v84561b;
assign v23fcc89 = hbusreq6_p & v22f8c01 | !hbusreq6_p & v23fcbaf;
assign v23f5f78 = hmaster0_p & v23fc4a8 | !hmaster0_p & v23f4926;
assign v22f5515 = stateG10_5_p & v230d346 | !stateG10_5_p & !v2309c8a;
assign v191b10f = hgrant3_p & v2302c6d | !hgrant3_p & v23f5fa6;
assign v23066bc = hmaster0_p & v23fb89c | !hmaster0_p & v230fe82;
assign v23056bc = hmaster2_p & v23fc23d | !hmaster2_p & v84561b;
assign v23fa3fc = hbusreq4 & v2308a8f | !hbusreq4 & v84561b;
assign v23fc7ce = hbusreq5_p & v23fcd96 | !hbusreq5_p & !v84561b;
assign v23fbba4 = hbusreq0 & v23fc23d | !hbusreq0 & v84561b;
assign v22f4b50 = hmaster2_p & v230aa1f | !hmaster2_p & v84561b;
assign a68bda = hgrant5_p & v2307729 | !hgrant5_p & v22f852d;
assign v22ee8f3 = hgrant1_p & v22fef02 | !hgrant1_p & v22f6ac8;
assign v23045f5 = hmaster2_p & v2300071 | !hmaster2_p & v23f15ac;
assign v22fdc17 = hbusreq5_p & v2310da0 | !hbusreq5_p & v23084c2;
assign a1b75e = hbusreq5_p & v2391d40 | !hbusreq5_p & v23f65ae;
assign v22fce8b = hmaster2_p & v15074fb | !hmaster2_p & v84561b;
assign v23fc739 = hready & v23f7326 | !hready & !v84561b;
assign v22fbbd0 = hmaster0_p & v1e840b4 | !hmaster0_p & v230fc64;
assign v23fbf45 = hmaster2_p & v23fbf8b | !hmaster2_p & !v23fc362;
assign v231330b = hlock3_p & v22f6cde | !hlock3_p & v23fc60a;
assign v22f2c8b = hmaster2_p & v23fc658 | !hmaster2_p & v23f9dd1;
assign v23fbd8e = jx2_p & v23fc15d | !jx2_p & !v22fd60f;
assign v23fcc39 = hbusreq4 & v230f795 | !hbusreq4 & v84561b;
assign v23fbfd3 = hmaster0_p & v23f70e3 | !hmaster0_p & v22fff0a;
assign v2306690 = hbusreq3 & v23f5dca | !hbusreq3 & !v23fbc6b;
assign v23f4451 = hbusreq4 & v2310aee | !hbusreq4 & v23fb8e5;
assign v1e8413d = hbusreq5_p & v23f63ab | !hbusreq5_p & v84561b;
assign v22f690f = hlock3_p & v239313a | !hlock3_p & v230a226;
assign v23f2abe = hbusreq5_p & v23f5ce0 | !hbusreq5_p & v22f4d68;
assign v1aad481 = hbusreq0_p & v22fa9be | !hbusreq0_p & v84561b;
assign v23f28a1 = hmaster0_p & v22eed68 | !hmaster0_p & v231324f;
assign v22f6fa9 = hbusreq4_p & v2301484 | !hbusreq4_p & v22f3699;
assign v2310a9a = hlock0_p & v845622 | !hlock0_p & v2312187;
assign v2306a6f = hgrant2_p & v23f6afa | !hgrant2_p & !v84561b;
assign v23f6e9c = hbusreq1_p & v23fcdce | !hbusreq1_p & v23098c0;
assign v22ee1b8 = hmaster2_p & v23fc22e | !hmaster2_p & v23101b1;
assign v23f5fd9 = hbusreq6 & v22efceb | !hbusreq6 & v84561b;
assign v23fcdcf = hbusreq0 & v890cdd | !hbusreq0 & v23fb966;
assign v2307206 = hmaster2_p & v2310bf5 | !hmaster2_p & v22f1faf;
assign v22f95c3 = hbusreq3_p & v23119e3 | !hbusreq3_p & v23fccf5;
assign v2305853 = hbusreq6_p & v230ad60 | !hbusreq6_p & v23fcc05;
assign v23093a7 = hbusreq1_p & v23fcbcd | !hbusreq1_p & !v2312259;
assign v23fc3c9 = hbusreq5 & v23fbfd0 | !hbusreq5 & v22f0add;
assign v22f9124 = hmaster2_p & v23ef8bb | !hmaster2_p & v23fc9de;
assign v22f3f68 = hgrant1_p & v84561b | !hgrant1_p & v230f256;
assign v22f4089 = hmaster0_p & v22ffea8 | !hmaster0_p & v1aad4ef;
assign v22f9396 = hbusreq4_p & v1e8439a | !hbusreq4_p & !v22f334c;
assign v23fc55f = hgrant2_p & v2303f9a | !hgrant2_p & v84564d;
assign v230115b = hbusreq5_p & v845636 | !hbusreq5_p & v23fccca;
assign v22ec7a2 = hbusreq0_p & v2303b9a | !hbusreq0_p & !b9d013;
assign v230995b = hbusreq0 & v23fb9c2 | !hbusreq0 & v84564d;
assign v22f1ee0 = hlock3_p & v23fcb56 | !hlock3_p & v23fcc9f;
assign v2368b8a = hbusreq5_p & v22eea63 | !hbusreq5_p & !v23fa9dd;
assign v22f7273 = hgrant3_p & v22fc9cb | !hgrant3_p & !v23fb60e;
assign a1fc9e = hbusreq4_p & v230ae4e | !hbusreq4_p & v23fc412;
assign v22fc163 = hbusreq6_p & v2304598 | !hbusreq6_p & v2301f50;
assign v230d630 = hmastlock_p & v22f2d83 | !hmastlock_p & v84561b;
assign v22f3f15 = hbusreq1 & v22f9911 | !hbusreq1 & v230f5a3;
assign v22fb4e3 = hmastlock_p & v22f7176 | !hmastlock_p & v84565f;
assign v230e1e0 = hmaster1_p & v2391fc6 | !hmaster1_p & v23fd00e;
assign v23f4da0 = hgrant1_p & v84561b | !hgrant1_p & v23f66a8;
assign v2302abd = hmaster2_p & v2305a12 | !hmaster2_p & v2309c28;
assign v23f2af5 = hmaster1_p & v23f5df1 | !hmaster1_p & v23f84dc;
assign v23fc46c = hbusreq4_p & v22f41c4 | !hbusreq4_p & v2308b9a;
assign v2303a74 = hmaster2_p & v2310434 | !hmaster2_p & v22f6756;
assign v230c116 = hbusreq1 & v995fa2 | !hbusreq1 & v84561b;
assign v23111ee = hbusreq5_p & v1aad9a6 | !hbusreq5_p & v23044e2;
assign v1aad31f = hmaster2_p & v22eb6ba | !hmaster2_p & v22fa156;
assign v22f2db9 = hbusreq1_p & v2308ae7 | !hbusreq1_p & v22f8c0b;
assign v22fe62a = hbusreq3_p & v22fa631 | !hbusreq3_p & v84562b;
assign v22f476c = stateG3_0_p & v84561b | !stateG3_0_p & v845665;
assign v230a65d = hmaster2_p & v22ef062 | !hmaster2_p & v2308765;
assign v23000a7 = jx1_p & v862ce7 | !jx1_p & v8632f2;
assign v22f41ee = hgrant0_p & v22f56d2 | !hgrant0_p & !v23fba79;
assign v230ca2b = hmaster2_p & v230ef5e | !hmaster2_p & v899296;
assign v23f4c50 = hmaster2_p & v1aae29a | !hmaster2_p & !v231228e;
assign v23fb11b = jx0_p & v23f957b | !jx0_p & v22ef481;
assign v230835d = hlock0_p & v2305c2e | !hlock0_p & v845620;
assign v23003cc = hlock0_p & v22ed85a | !hlock0_p & v230e295;
assign v2301a90 = hmaster2_p & v845636 | !hmaster2_p & v150745f;
assign v23f600f = hgrant3_p & v22ee6cb | !hgrant3_p & v22fe415;
assign v22ef769 = hgrant5_p & v84561b | !hgrant5_p & v231032d;
assign v23fc110 = hlock6_p & v23fcab8 | !hlock6_p & v231181c;
assign v22f6f16 = hbusreq0 & v22ee0c4 | !hbusreq0 & v84561b;
assign v22f1cc5 = jx3_p & v22fa309 | !jx3_p & v2302dc1;
assign v22ed000 = hgrant1_p & v230fec6 | !hgrant1_p & v23fce3f;
assign v22fdf28 = hbusreq4_p & v22f446b | !hbusreq4_p & v23fb533;
assign v23f6635 = hmaster2_p & v23fa2ec | !hmaster2_p & v2309c28;
assign v2391e0c = hbusreq3 & v23fcc49 | !hbusreq3 & v84561b;
assign v2304e28 = hmaster0_p & v84561b | !hmaster0_p & v23fca08;
assign v230834c = hbusreq0_p & v2303972 | !hbusreq0_p & v2313372;
assign v2301a99 = hmaster0_p & v22fd7d4 | !hmaster0_p & !v22fdd8a;
assign v23fc013 = hmaster0_p & v23f5461 | !hmaster0_p & v230f790;
assign v2300ac2 = hgrant1_p & v2312e02 | !hgrant1_p & v2307742;
assign v23f350b = hbusreq4 & v230fb9e | !hbusreq4 & v845627;
assign v22fbf74 = hbusreq2_p & v84561b | !hbusreq2_p & v230eb9b;
assign v2305841 = hmaster2_p & v22f9c37 | !hmaster2_p & !v23126be;
assign v86c49f = hmaster1_p & v22fe1c8 | !hmaster1_p & v22f6af6;
assign v12cd523 = hbusreq2_p & v23019e7 | !hbusreq2_p & !v84561b;
assign v2309733 = hbusreq3_p & v230f92a | !hbusreq3_p & !v84561b;
assign v1aada8c = hbusreq3_p & v23fc3e8 | !hbusreq3_p & !v23fb7c3;
assign v1507631 = hlock6_p & v22fc3d9 | !hlock6_p & v22f591c;
assign v22f9ab6 = hgrant3_p & v22f2ca2 | !hgrant3_p & v22fa646;
assign v230b68b = hmaster2_p & v22fa70c | !hmaster2_p & !v2306932;
assign v2311790 = hmaster1_p & v22fd841 | !hmaster1_p & v23fc1d1;
assign v22fb4d8 = hmaster0_p & af7272 | !hmaster0_p & fc8fe6;
assign v22eb332 = hbusreq5 & v23105cd | !hbusreq5 & v84561b;
assign v23fa69e = jx1_p & v22fa0b2 | !jx1_p & v23fbb81;
assign v239158e = hmaster0_p & v84561b | !hmaster0_p & !v22fe908;
assign v22ed5c8 = hmaster2_p & v23fc40f | !hmaster2_p & v2304bc1;
assign v2393909 = hgrant3_p & v23f651a | !hgrant3_p & !v23f2f5d;
assign v23f06ee = hbusreq3_p & v2302131 | !hbusreq3_p & !v84561b;
assign v22ef92c = hbusreq5_p & v84561b | !hbusreq5_p & !v22fd720;
assign c20a75 = hmaster2_p & v22f4986 | !hmaster2_p & !v23041e2;
assign v2308765 = hbusreq1_p & v23065b6 | !hbusreq1_p & v84561b;
assign v23fc6dd = hgrant4_p & v23fc095 | !hgrant4_p & v23052a2;
assign v23f8465 = hgrant1_p & v84561b | !hgrant1_p & v23fb505;
assign v22f586f = hbusreq1_p & v23f9789 | !hbusreq1_p & v22f0945;
assign v23fad54 = hmaster1_p & v2312edb | !hmaster1_p & v84561b;
assign v23135ca = hbusreq3 & v230adb7 | !hbusreq3 & v84561b;
assign v22eda7c = hbusreq2_p & b9d00f | !hbusreq2_p & a1fba6;
assign v230fbe2 = hready_p & v23046a7 | !hready_p & !v23fbd91;
assign v22fa8d7 = hbusreq6_p & v2311358 | !hbusreq6_p & v22fae9f;
assign v2306885 = hbusreq0_p & v231339c | !hbusreq0_p & !v23f8638;
assign v23f20d7 = hlock0_p & v23fbdd4 | !hlock0_p & v2309221;
assign v22f3189 = hbusreq3_p & v230118f | !hbusreq3_p & v2309c93;
assign v23fbe94 = hbusreq4_p & v23fc940 | !hbusreq4_p & v22f2d10;
assign v23fc128 = hmaster0_p & v23f7039 | !hmaster0_p & !v22f8f56;
assign v23f79ba = hbusreq6 & v230c9f0 | !hbusreq6 & v84561b;
assign v230bb2d = hbusreq3_p & v23f0c76 | !hbusreq3_p & !v23fc5eb;
assign v230979d = hmaster2_p & v23f4808 | !hmaster2_p & v22fc7e6;
assign v23fcc8e = hbusreq1 & v1aae56f | !hbusreq1 & v84564d;
assign v23fcbde = hlock5_p & v85bd38 | !hlock5_p & v230aef9;
assign v230f2f5 = hbusreq2 & v84561b | !hbusreq2 & !v230abfb;
assign v2300bb5 = hbusreq3 & v2313351 | !hbusreq3 & v230886c;
assign v22ebe16 = hbusreq0 & v230f5a3 | !hbusreq0 & v84561b;
assign v230716d = hmaster1_p & v84561b | !hmaster1_p & v22f63cc;
assign v22ed0d9 = hgrant1_p & v84561b | !hgrant1_p & v22faf60;
assign v22f7a1d = hmaster0_p & v23fb7b4 | !hmaster0_p & a04d83;
assign v23fc827 = hmaster0_p & v23fba32 | !hmaster0_p & !v96c563;
assign v23f0aec = hgrant3_p & v22f04c8 | !hgrant3_p & v23fb672;
assign v23fbd70 = hmaster2_p & v23f9b8d | !hmaster2_p & v23fca72;
assign v23015f8 = hlock0_p & v230e4ef | !hlock0_p & v22f2a24;
assign v22f35eb = hgrant6_p & v230226e | !hgrant6_p & v22fbab1;
assign v22f5d5e = jx1_p & v23fcc64 | !jx1_p & v23fcfe8;
assign v22ff21b = hmaster2_p & v2306d29 | !hmaster2_p & v22f56d2;
assign b7d0f1 = jx1_p & v85fd50 | !jx1_p & v84561b;
assign v22f7b47 = hgrant1_p & v23fa2ec | !hgrant1_p & v22f108e;
assign v22f1ef6 = hbusreq5_p & v23fbf87 | !hbusreq5_p & !v84561b;
assign v230b04e = hbusreq5 & v22ff090 | !hbusreq5 & v84561b;
assign v22ef026 = hbusreq3_p & v22eda0b | !hbusreq3_p & v84561b;
assign v23fc7ca = hmaster0_p & v23fb73d | !hmaster0_p & !v23fc91c;
assign v22eeb7d = hgrant5_p & v84561b | !hgrant5_p & v230a941;
assign v230685f = hbusreq3_p & v23fc5d0 | !hbusreq3_p & v23051cf;
assign v23fc162 = hmaster2_p & v2302a4d | !hmaster2_p & !v191a876;
assign v23f3997 = hbusreq1_p & v22feb98 | !hbusreq1_p & v84561b;
assign v230415a = hgrant0_p & v84561b | !hgrant0_p & !v23fbb1c;
assign v23065ee = hmaster1_p & v22eea52 | !hmaster1_p & v22f7a60;
assign v230259a = hbusreq1_p & v22ed614 | !hbusreq1_p & bab0c9;
assign v9ae938 = hmaster0_p & v23fce2c | !hmaster0_p & v23fb976;
assign v23fb9be = hlock2_p & b00ad3 | !hlock2_p & v84561b;
assign v230942e = hlock0_p & v23fcd76 | !hlock0_p & v23fc5a8;
assign v22ee41e = jx0_p & v23047f9 | !jx0_p & v23fc0cd;
assign v22f7ef4 = hgrant5_p & v231007d | !hgrant5_p & v22f4d46;
assign v22ee142 = hmaster0_p & v23fb89c | !hmaster0_p & v22f1ab6;
assign v22eb629 = hbusreq6_p & v23fc3ca | !hbusreq6_p & v22f0dd3;
assign v22f20d3 = hbusreq5 & v2304e69 | !hbusreq5 & v22f6058;
assign v22ff89d = hbusreq5 & v13afe3a | !hbusreq5 & !fc8ab7;
assign v23fb53b = hgrant5_p & v23fc388 | !hgrant5_p & v23fbacb;
assign v23f9a81 = hmaster2_p & v22fe5b1 | !hmaster2_p & v22f9880;
assign v23fb07c = hmaster2_p & v2312231 | !hmaster2_p & v2309456;
assign v22f664f = hmaster1_p & v23fc4a7 | !hmaster1_p & v23031bc;
assign v230665f = hlock1_p & v22f2718 | !hlock1_p & !v84561b;
assign v231108b = hbusreq6_p & v230a02b | !hbusreq6_p & v22f5eae;
assign v2302386 = stateG10_5_p & v22ec61a | !stateG10_5_p & v22fbf74;
assign v2305b2e = hbusreq3_p & v2309c93 | !hbusreq3_p & v22f511c;
assign v22f2430 = hgrant1_p & v84561b | !hgrant1_p & v23f8a36;
assign v2308356 = hgrant0_p & v23fc94c | !hgrant0_p & !v23003b8;
assign v2306844 = hbusreq3 & v23126b8 | !hbusreq3 & v84561b;
assign v23f4c5b = hbusreq6 & v22ff5bd | !hbusreq6 & v84561b;
assign v2309c8a = busreq_p & v106ae19 | !busreq_p & !v23f7ffb;
assign v2308f85 = stateA1_p & v23fc683 | !stateA1_p & v23fbbb2;
assign v22f2e20 = hmaster0_p & v2308ba7 | !hmaster0_p & b00aa6;
assign v22fd699 = hgrant5_p & v22f0323 | !hgrant5_p & c258f4;
assign v23fc884 = hmaster2_p & v23fcb69 | !hmaster2_p & v22ff732;
assign v23fb138 = hbusreq3 & v2301bdb | !hbusreq3 & v2303e23;
assign v22fa5c9 = hbusreq5 & v230882d | !hbusreq5 & v23f8364;
assign v22ee920 = hlock4_p & v23fc02e | !hlock4_p & v23f917f;
assign v22f2c2c = hlock5_p & v23fb1f1 | !hlock5_p & ba569c;
assign v2306070 = stateG2_p & v84561b | !stateG2_p & !v22faac8;
assign v845655 = hgrant3_p & v84561b | !hgrant3_p & !v84561b;
assign v23fc2f2 = hgrant4_p & v23fbf73 | !hgrant4_p & !v23fc300;
assign v22eb3ad = hbusreq5_p & v845636 | !hbusreq5_p & v22fe74e;
assign v22f587e = locked_p & v22f6bd4 | !locked_p & !v84561b;
assign v12cd5f2 = hbusreq6 & v2302131 | !hbusreq6 & v84561b;
assign v949c12 = hlock3_p & v22edb43 | !hlock3_p & !v84561b;
assign v23fcc45 = hlock4_p & v230716c | !hlock4_p & v23125a2;
assign v230a730 = hbusreq4 & v22eef9f | !hbusreq4 & v23fb8e5;
assign v2305b35 = hbusreq5_p & v84561b | !hbusreq5_p & !v106a782;
assign v23f3ff9 = hgrant3_p & v84562e | !hgrant3_p & v22fe7b0;
assign v22f1efd = hbusreq6_p & v22fa5a6 | !hbusreq6_p & v23f35de;
assign v2392bc1 = hbusreq5 & v23f3ca5 | !hbusreq5 & v84561b;
assign v23fd010 = hbusreq6_p & v23fc5db | !hbusreq6_p & !v2310b47;
assign v22f288d = hmaster0_p & v17a34ff | !hmaster0_p & !v22f6917;
assign v230b82e = hmaster0_p & v23fc92c | !hmaster0_p & v230f087;
assign v2310e4a = hbusreq6 & v22fc4a3 | !hbusreq6 & v23fcf43;
assign v22ec2a4 = hbusreq3 & v23fc7db | !hbusreq3 & v84561b;
assign v845637 = hlock5_p & v84561b | !hlock5_p & !v84561b;
assign v23fc3fb = hbusreq1_p & v230580d | !hbusreq1_p & v2300d32;
assign v191aa68 = hmastlock_p & v1aad6c8 | !hmastlock_p & v84565f;
assign v23017f0 = hgrant2_p & v845620 | !hgrant2_p & v84561b;
assign v23fb98c = hbusreq5_p & v23fbb0b | !hbusreq5_p & !v22f6056;
assign v2311d38 = hmaster2_p & v22f3643 | !hmaster2_p & v84561b;
assign v22f20cf = hlock4_p & v2301f8c | !hlock4_p & v2301968;
assign v22f334c = hmaster0_p & v23fae84 | !hmaster0_p & !v22f16bf;
assign v2309c55 = hbusreq1 & v22ede16 | !hbusreq1 & v22f7241;
assign v230c5ad = stateG10_5_p & v22f61cc | !stateG10_5_p & v22fb3df;
assign v22f25a1 = hgrant3_p & v23fb699 | !hgrant3_p & v230b086;
assign v23fc260 = hbusreq3_p & v23fce15 | !hbusreq3_p & v84561b;
assign v22f910f = hgrant1_p & v845625 | !hgrant1_p & v23fb33a;
assign v22f23f6 = hlock3_p & v22f78c3 | !hlock3_p & v23065fc;
assign v23fc71a = hbusreq3_p & v22fb32a | !hbusreq3_p & v22eee99;
assign v23f1e1b = hmaster0_p & v231345a | !hmaster0_p & v230dce6;
assign v230207d = hbusreq0_p & v231124e | !hbusreq0_p & v22fb841;
assign v2302c91 = hbusreq3_p & v22f3c27 | !hbusreq3_p & v23fbf97;
assign v2300c56 = hbusreq3_p & v23f9758 | !hbusreq3_p & v84561b;
assign v23f51da = hgrant1_p & v23fa623 | !hgrant1_p & !v84561b;
assign v23040a8 = hmaster0_p & v23f54a0 | !hmaster0_p & v23fc785;
assign v22fa4a3 = hbusreq6_p & v23fa967 | !hbusreq6_p & v23fb957;
assign v22edcf1 = hbusreq1_p & v22fbeea | !hbusreq1_p & v23fc4c0;
assign v22f7713 = hgrant3_p & v230e882 | !hgrant3_p & v23f3c3b;
assign v23fc9a5 = hlock3_p & v2312b5a | !hlock3_p & v230197e;
assign v230070e = hbusreq3_p & v22fe920 | !hbusreq3_p & v23fb906;
assign v23f347b = hmaster0_p & v2307061 | !hmaster0_p & v23fc7f9;
assign v23f5f18 = hmaster2_p & v106ae19 | !hmaster2_p & !v23f5596;
assign v2302e9e = hgrant1_p & v84561b | !hgrant1_p & v22f7378;
assign v23fcb55 = hgrant1_p & v84561b | !hgrant1_p & v230941d;
assign v230ca57 = hmaster2_p & v22f17bb | !hmaster2_p & v22fc2bd;
assign v230e336 = hbusreq1_p & v230c342 | !hbusreq1_p & !v22ff457;
assign v23f7ce8 = hmaster2_p & v23fb90c | !hmaster2_p & v845620;
assign v23fbf1d = hbusreq1_p & v22faf60 | !hbusreq1_p & v22f6c1b;
assign v22ee457 = hbusreq5_p & v230b8cd | !hbusreq5_p & v22f4678;
assign v230446b = hbusreq6_p & v23fbe9d | !hbusreq6_p & v22f758c;
assign v23fccb5 = hgrant3_p & v84561b | !hgrant3_p & !v1aad45d;
assign v23f594f = hbusreq4_p & v23fc1aa | !hbusreq4_p & v23fb787;
assign v22fc7c2 = hbusreq1_p & v23f4d72 | !hbusreq1_p & v23f9a37;
assign v2302e73 = hmaster2_p & v2308d79 | !hmaster2_p & v23131e8;
assign v13afc19 = decide_p & v23007d9 | !decide_p & v2302c31;
assign v2307009 = hmaster2_p & v22f1ae7 | !hmaster2_p & v23fb175;
assign v23fc618 = hbusreq3_p & v23fc7a7 | !hbusreq3_p & v23117c1;
assign v23fc7f2 = hbusreq6_p & v23fce1b | !hbusreq6_p & !v230b77e;
assign v12cda0a = hmaster2_p & v2304ad5 | !hmaster2_p & v23f4808;
assign v23fbe0d = stateG10_5_p & v23fc5fe | !stateG10_5_p & v845620;
assign v23fc61d = hmaster0_p & v23f38a5 | !hmaster0_p & v22f0f36;
assign v15072de = hbusreq2 & v84564d | !hbusreq2 & v84561b;
assign v23f908f = hlock0_p & v84561b | !hlock0_p & v22f6f8f;
assign v2313189 = hbusreq4_p & v23fcafc | !hbusreq4_p & v22ed55a;
assign v191b1d9 = hmaster0_p & v22ebb82 | !hmaster0_p & v22f160c;
assign v23fc36e = hgrant0_p & v22fb00d | !hgrant0_p & v23fc8c3;
assign v23fb096 = hbusreq5 & v23fc530 | !hbusreq5 & !v84562a;
assign v22ec8d7 = hbusreq3_p & v230e860 | !hbusreq3_p & !v84561b;
assign v22f317b = hmaster2_p & v230945e | !hmaster2_p & v22ff732;
assign v22ebf90 = jx0_p & v23fbc95 | !jx0_p & v106a7d8;
assign v230cb9d = stateG2_p & v2302ca3 | !stateG2_p & !v22f349a;
assign v23fc169 = hmaster0_p & v23051fc | !hmaster0_p & v22f1fdb;
assign v23f437e = hlock6_p & v23fc4df | !hlock6_p & v2305933;
assign v23f1ec4 = hmaster2_p & v84561b | !hmaster2_p & !v845635;
assign v22f5568 = hbusreq3_p & v22fed5c | !hbusreq3_p & v23f3f40;
assign v231326a = hgrant5_p & v84561b | !hgrant5_p & v230c4bb;
assign v23f1fad = hmaster2_p & v23131e8 | !hmaster2_p & !v23fc017;
assign v22ecee2 = hbusreq2 & v230d630 | !hbusreq2 & !v84561b;
assign v23a2d0a = hready_p & v22fc837 | !hready_p & v845645;
assign v2312343 = stateG10_5_p & v230ba0a | !stateG10_5_p & !v23f908f;
assign v22fd2a3 = hmaster0_p & v2309e8e | !hmaster0_p & !v84561b;
assign v2393118 = hmaster2_p & v84561b | !hmaster2_p & v23f51e3;
assign v23fb980 = hbusreq5_p & v23930d2 | !hbusreq5_p & !v84561b;
assign v23fc8cf = hmaster1_p & v23fbff0 | !hmaster1_p & v230278d;
assign v23fa1f4 = hbusreq2 & v230f5a3 | !hbusreq2 & v84561b;
assign v23fc9cb = hbusreq5 & v2300c5a | !hbusreq5 & v84561b;
assign v22efc21 = hbusreq3 & v230a05f | !hbusreq3 & c16218;
assign v23f54ef = hlock0_p & v84561b | !hlock0_p & !v22f49c4;
assign v230b267 = hmaster2_p & v2306220 | !hmaster2_p & !v23fc017;
assign v15071da = stateA1_p & v84561b | !stateA1_p & !v23fa931;
assign v22ec37c = jx1_p & v23f651e | !jx1_p & v230095f;
assign v2393bcf = jx0_p & v23fcb8f | !jx0_p & v22f7289;
assign v230790b = hbusreq4 & v23fca10 | !hbusreq4 & v230f0de;
assign v23fcc84 = hmaster0_p & a1fbe9 | !hmaster0_p & v23f8689;
assign v22fc7e5 = hmaster0_p & v23fb045 | !hmaster0_p & v23fbb28;
assign v22efe1b = hbusreq3 & v23f232a | !hbusreq3 & !v22fde54;
assign v23f8913 = hmaster2_p & v22feae3 | !hmaster2_p & v23f8d76;
assign v230f151 = hmaster1_p & v22fa976 | !hmaster1_p & v15072a7;
assign v22f6d6e = hmaster0_p & v22fe869 | !hmaster0_p & v231147e;
assign v23fc4f9 = hgrant1_p & v12cd9f9 | !hgrant1_p & v22fba66;
assign v23f08a4 = hgrant1_p & v84561b | !hgrant1_p & v230f9e8;
assign v22f50ae = hmaster0_p & v23f8e04 | !hmaster0_p & v845625;
assign v22f7c32 = jx1_p & v230fe71 | !jx1_p & v22fc588;
assign v2302812 = hbusreq3 & v22f1c40 | !hbusreq3 & v22eebf5;
assign v9d0518 = hlock4_p & v22f52a0 | !hlock4_p & v23f60ba;
assign v23fceb5 = jx0_p & v2300b33 | !jx0_p & v23fc679;
assign v23fc9dc = hgrant3_p & v22eeb06 | !hgrant3_p & v230e8a8;
assign v23fcb94 = jx2_p & v23fc403 | !jx2_p & v23fc053;
assign v22fd8a4 = hbusreq3_p & v23f35ff | !hbusreq3_p & !v84561b;
assign v23039c8 = hbusreq6 & v22effdf | !hbusreq6 & v230829b;
assign v22f9078 = hgrant1_p & v84561b | !hgrant1_p & !v23f4761;
assign v22f18b4 = stateG10_5_p & v230f050 | !stateG10_5_p & !v2302e32;
assign v23fc4e0 = hmaster2_p & v84561b | !hmaster2_p & v23fc5f4;
assign v23f21e5 = hbusreq0 & v23fc48b | !hbusreq0 & v84561b;
assign v1506af9 = decide_p & v22ffc85 | !decide_p & v230fbe2;
assign v230c37d = hbusreq3_p & v23064ce | !hbusreq3_p & v23fc798;
assign v23fbe80 = hbusreq1_p & v230e4ef | !hbusreq1_p & v230ece0;
assign v22faf41 = hlock4_p & v22f4321 | !hlock4_p & v23f9c04;
assign v22eb3e3 = hgrant1_p & v22fcf7a | !hgrant1_p & v23fc59a;
assign v23f3ccf = hbusreq1_p & v22f7752 | !hbusreq1_p & !v84561b;
assign v23f5fc3 = hlock3_p & v8963c2 | !hlock3_p & v22f6e30;
assign v23139ef = hbusreq3_p & v230eafa | !hbusreq3_p & v22f7861;
assign v2393b99 = hmaster2_p & v23080ec | !hmaster2_p & v2309729;
assign v23fcbbb = hbusreq6_p & v23f6827 | !hbusreq6_p & a6c3d1;
assign v2301312 = hbusreq5 & v2313118 | !hbusreq5 & v23f1879;
assign v23f2353 = hmaster0_p & v191ad8e | !hmaster0_p & v23fb95f;
assign v23fba49 = hbusreq5_p & v23f200b | !hbusreq5_p & v2309c93;
assign v22f337b = hready & v230f6a7 | !hready & !v84561b;
assign v22eaf7a = locked_p & v22f03aa | !locked_p & v84561b;
assign v23fbff1 = jx0_p & v22fa99c | !jx0_p & v22f8c55;
assign v22f70d2 = hgrant1_p & v22f619f | !hgrant1_p & !v84561b;
assign v23f2c05 = hbusreq5_p & v23fc661 | !hbusreq5_p & !v84561b;
assign v2311831 = hgrant3_p & v23f9b49 | !hgrant3_p & v22f5125;
assign v22fd55f = hbusreq4 & v23f0dd1 | !hbusreq4 & v84561b;
assign v22efc04 = hmaster2_p & v230b125 | !hmaster2_p & v23fae9e;
assign v230b131 = hgrant3_p & v23f1643 | !hgrant3_p & v23f543d;
assign v22f036f = hmaster1_p & v1aae374 | !hmaster1_p & v2302348;
assign v22f031f = hbusreq3_p & v1e83f8d | !hbusreq3_p & v230697e;
assign v230fab4 = hlock5_p & v23f659c | !hlock5_p & v1b87690;
assign v22ebad7 = hbusreq0 & v22ef513 | !hbusreq0 & v84561b;
assign v22ede34 = hmaster2_p & v23fcfbb | !hmaster2_p & v84561b;
assign v150715d = hgrant5_p & v2309ab5 | !hgrant5_p & v22ec562;
assign bd1c32 = hgrant3_p & v84562e | !hgrant3_p & v23126f2;
assign v23fb5e3 = hbusreq0 & v22febe1 | !hbusreq0 & v84561b;
assign v22f5664 = hbusreq6 & v2307f77 | !hbusreq6 & v84561b;
assign v22fdd56 = hgrant3_p & v84562e | !hgrant3_p & v22ed067;
assign v22f24a3 = hbusreq6 & v191b1b9 | !hbusreq6 & v22fc22b;
assign v23f6f99 = hmaster2_p & v23fa2ec | !hmaster2_p & !v23fc9db;
assign v22f0e84 = jx1_p & v230f073 | !jx1_p & v230d282;
assign v22f81a7 = hbusreq4_p & v2302e7b | !hbusreq4_p & !v22f9cd9;
assign v230b19a = hmaster2_p & v2346b6a | !hmaster2_p & b10190;
assign v23fb879 = hmaster2_p & v22f1b4e | !hmaster2_p & v230a9eb;
assign v23086ef = hmaster2_p & v22f343b | !hmaster2_p & !v22f15fe;
assign v22f5c70 = hgrant3_p & v84561b | !hgrant3_p & v22fe60b;
assign v23fb845 = hbusreq6 & v23fb0c0 | !hbusreq6 & v84561b;
assign v22f5198 = hlock3_p & v22ec6e5 | !hlock3_p & v84561b;
assign v23f7795 = hgrant5_p & v2304299 | !hgrant5_p & !v22fdca9;
assign v22eea0f = hbusreq6_p & v22fab33 | !hbusreq6_p & v23fc616;
assign v22fc741 = hgrant1_p & v845626 | !hgrant1_p & v23f8536;
assign v22fd61b = hmaster0_p & v2308e0b | !hmaster0_p & v22fe181;
assign v230fb99 = hlock0_p & afc788 | !hlock0_p & v23fcabb;
assign v22ef242 = hmaster0_p & v22f97c3 | !hmaster0_p & !v106ae5a;
assign v23fbf0f = hlock3_p & v22ff2bf | !hlock3_p & v22f9374;
assign v23f1a1f = hlock6_p & v23111a4 | !hlock6_p & !v84561b;
assign v23fc1c9 = hlock2_p & v23f4bcd | !hlock2_p & v845620;
assign v22fa58f = hmaster2_p & v239383d | !hmaster2_p & !v12cc2ef;
assign v2313328 = jx2_p & v23f4a0f | !jx2_p & v22f43ec;
assign v23fc575 = hlock4_p & v22feb04 | !hlock4_p & !v230a0ad;
assign v22ff4e2 = hmaster2_p & v22f343b | !hmaster2_p & !v2301655;
assign v22f971f = hmaster2_p & v23fcb83 | !hmaster2_p & v23fc511;
assign v230c69b = hgrant1_p & v23f83ef | !hgrant1_p & v23f680b;
assign v23efe0a = hgrant0_p & v23133fa | !hgrant0_p & v23fc842;
assign v23fc3a4 = hbusreq3_p & v23fbcad | !hbusreq3_p & v84564d;
assign v22ede7f = hlock5_p & v230a9eb | !hlock5_p & !v12cd3f4;
assign v23fba66 = hmaster1_p & v23fcbf0 | !hmaster1_p & v23f1c0b;
assign v23fb672 = hmaster2_p & v22ff9d7 | !hmaster2_p & v84561b;
assign v23fce89 = hmaster0_p & v22fa0ec | !hmaster0_p & !v22ff21b;
assign v23fc5f8 = hbusreq3_p & v2392a3a | !hbusreq3_p & v22fe831;
assign v2304e0f = hmaster0_p & v23fc6a1 | !hmaster0_p & v230b38b;
assign v22efc28 = hmaster2_p & v22f7da7 | !hmaster2_p & v23fc741;
assign v230a735 = hbusreq3 & v23086ef | !hbusreq3 & !v22f4d37;
assign v22f7c44 = hbusreq3_p & v23f31a9 | !hbusreq3_p & v84561b;
assign v23f91d0 = hgrant3_p & v84562e | !hgrant3_p & v23fc275;
assign v191b1b9 = hgrant3_p & v22fb1bc | !hgrant3_p & v23f9ef5;
assign v2391fae = stateG10_5_p & v23fc3cb | !stateG10_5_p & a1fbc2;
assign v23f692f = hmaster2_p & v22fd696 | !hmaster2_p & v1507102;
assign v2392ef6 = hgrant3_p & v22efa0a | !hgrant3_p & v23fc194;
assign v2303147 = hbusreq1_p & v2301997 | !hbusreq1_p & v230ca7c;
assign v22f7a0c = hbusreq5_p & v230e07d | !hbusreq5_p & v22f3a6f;
assign v230e01b = hgrant3_p & v23fbe79 | !hgrant3_p & v23fc66d;
assign v23fb745 = hbusreq3 & v230fb76 | !hbusreq3 & v23f2d33;
assign v2301e20 = hbusreq0 & v13affaa | !hbusreq0 & v84564d;
assign v23fb8a8 = hlock1_p & v23fbadc | !hlock1_p & v845620;
assign c60af7 = hbusreq3 & v22f4f19 | !hbusreq3 & v84561b;
assign v230f161 = jx0_p & v2391e26 | !jx0_p & !v23f623e;
assign v230b011 = hbusreq5_p & v84564d | !hbusreq5_p & v23f7921;
assign v22fc5f0 = hlock0_p & v23082ec | !hlock0_p & v23f4b28;
assign v22fe343 = hgrant1_p & v84561b | !hgrant1_p & v230f755;
assign v23fcfa8 = hbusreq3_p & v23f5ae4 | !hbusreq3_p & !v23fcd8a;
assign v23f4a00 = hbusreq5 & v22fe421 | !hbusreq5 & v84561b;
assign v22fab02 = hmaster2_p & v23f2ec0 | !hmaster2_p & !v84561b;
assign v2302245 = hbusreq4_p & v2301292 | !hbusreq4_p & v22ec0d1;
assign v2310904 = locked_p & v84561b | !locked_p & !v23fb861;
assign v2391e8f = hbusreq3 & v230f538 | !hbusreq3 & v84564d;
assign v230e473 = hmaster2_p & v23fc89a | !hmaster2_p & v2306b2e;
assign v22fd6a4 = hbusreq1 & v22f6ac8 | !hbusreq1 & v84561b;
assign v23fc89b = hgrant3_p & v84561b | !hgrant3_p & !v22ff3e6;
assign v23fb66e = hbusreq4_p & v23f52b9 | !hbusreq4_p & v22fc399;
assign v23094ad = hbusreq0_p & v23126ae | !hbusreq0_p & v106af73;
assign v22f7e21 = hgrant3_p & v23f651a | !hgrant3_p & v23fcb99;
assign v22f2ed7 = hbusreq5_p & v84564d | !hbusreq5_p & v22f3643;
assign v22fea3e = hmaster2_p & v22f83cf | !hmaster2_p & v2391f2b;
assign v23fc106 = hmaster2_p & v2308110 | !hmaster2_p & !v12cc2ef;
assign v23fcebf = hmaster2_p & v23fcc70 | !hmaster2_p & a1fba6;
assign v23f3c86 = jx1_p & v23f651e | !jx1_p & v22f811e;
assign v2304856 = hbusreq6 & v22ef76f | !hbusreq6 & v84562d;
assign v230c0e9 = hbusreq2_p & v22fcf3e | !hbusreq2_p & !v23fa91a;
assign v2304fe7 = hgrant1_p & v845626 | !hgrant1_p & v23f133b;
assign v22f28aa = hgrant3_p & v23f9110 | !hgrant3_p & v23fc0c6;
assign v22eda36 = hlock2_p & v84561b | !hlock2_p & v13afe3a;
assign v23f3bc9 = hgrant3_p & v23125fb | !hgrant3_p & v2312f44;
assign v23f886a = hbusreq6_p & v2304d59 | !hbusreq6_p & v22fd079;
assign v22f0fb9 = hmaster2_p & v84564d | !hmaster2_p & !v2304ec7;
assign v230a117 = locked_p & v23081eb | !locked_p & v84561b;
assign v23fbe39 = hbusreq0_p & v22ebad7 | !hbusreq0_p & v84561b;
assign v2301abc = hbusreq0 & v2312bd0 | !hbusreq0 & v84561b;
assign v2302e47 = stateG2_p & v22f9369 | !stateG2_p & v23f8ecc;
assign v1507088 = hbusreq0_p & a1fc4e | !hbusreq0_p & !v22edaf2;
assign v22efc42 = hgrant5_p & v23fc2ba | !hgrant5_p & v230f050;
assign v2303329 = hgrant5_p & v22eaff1 | !hgrant5_p & !v22fb71d;
assign v9ad48f = hgrant3_p & v84562e | !hgrant3_p & v23f0872;
assign v2309bab = hmaster0_p & v23fcaa5 | !hmaster0_p & v23fcb3f;
assign v230a44f = hmaster2_p & v23ef8bb | !hmaster2_p & v23135fa;
assign v22f063d = hgrant3_p & v22f56c2 | !hgrant3_p & v23f4194;
assign v23fbcc0 = hbusreq5_p & v84564d | !hbusreq5_p & v23940ce;
assign v22ee581 = hlock2_p & v23f6411 | !hlock2_p & !v106ae19;
assign v23f596f = hbusreq5 & v22f0073 | !hbusreq5 & v15074fb;
assign v23fc378 = hmastlock_p & v1aad6c8 | !hmastlock_p & !v84561b;
assign v2306f4e = hmaster1_p & v231156b | !hmaster1_p & v84561b;
assign v230aec3 = jx2_p & v23fc403 | !jx2_p & v230f161;
assign v22f4bea = hbusreq3_p & v23fc5b6 | !hbusreq3_p & b7ab40;
assign v23fb8ee = stateG2_p & v84561b | !stateG2_p & v22faac8;
assign v23f76a5 = hbusreq4 & v22f05b9 | !hbusreq4 & !v84562a;
assign v2311ed7 = hbusreq5_p & v23fb67c | !hbusreq5_p & v230bdbb;
assign v23fc4a5 = hready & v23f7326 | !hready & v13afe3a;
assign v22f3294 = hburst0_p & v23fc116 | !hburst0_p & !v2309a51;
assign v230f654 = hready & v22fa2de | !hready & v230c899;
assign v2309f1a = hbusreq3_p & v22f695c | !hbusreq3_p & v13afe72;
assign v23f8ba7 = hmaster0_p & v23f8787 | !hmaster0_p & v23fbf68;
assign v23f0bbc = jx3_p & v84561b | !jx3_p & v23f6ef7;
assign v23fba70 = hbusreq0 & v22f60c6 | !hbusreq0 & v84561b;
assign v23fb9c7 = hbusreq4_p & v2302983 | !hbusreq4_p & v2311761;
assign v23f4bbd = hgrant5_p & v23f9d5f | !hgrant5_p & !v22fd973;
assign v230bb63 = hbusreq1 & v2306220 | !hbusreq1 & !v84561b;
assign v231171d = hbusreq5_p & v23f033c | !hbusreq5_p & !v22faee9;
assign v23fc85c = hmaster2_p & v22fcdf6 | !hmaster2_p & v1aae56f;
assign v23f4a2c = hgrant0_p & v22fbea4 | !hgrant0_p & !v84561b;
assign v22f05b4 = hbusreq4_p & v23139c9 | !hbusreq4_p & v22f3832;
assign v23053fb = hbusreq3_p & v22f4a68 | !hbusreq3_p & v23fd011;
assign v23fa397 = hbusreq5_p & v23fbbc9 | !hbusreq5_p & !v84561b;
assign v23f7698 = hbusreq3 & v22f1c40 | !hbusreq3 & v22f0fb9;
assign v23f215c = hbusreq6_p & v22f09b1 | !hbusreq6_p & v23fb947;
assign v23fcb8d = hlock3_p & v23fccbf | !hlock3_p & v84561b;
assign v22f7347 = hgrant3_p & v84561b | !hgrant3_p & v22f61b6;
assign v2305992 = hbusreq6_p & v2304e0f | !hbusreq6_p & v22ed7da;
assign v23fc1c2 = hmaster2_p & v22f23a1 | !hmaster2_p & v84561b;
assign v23faa52 = hlock5_p & v106ae1c | !hlock5_p & a1fbb6;
assign v85e5cf = hmaster1_p & v845625 | !hmaster1_p & v22f50ae;
assign v2310c54 = hbusreq4_p & v22f79c8 | !hbusreq4_p & !v84561b;
assign v2312ad7 = hgrant3_p & v23fc975 | !hgrant3_p & v230952f;
assign v23fc4b1 = hbusreq1_p & v2310826 | !hbusreq1_p & v84561b;
assign v22fbc04 = hmaster1_p & v22fd841 | !hmaster1_p & v22f41c4;
assign v22f2c72 = hbusreq3 & v2311629 | !hbusreq3 & v84561b;
assign v230b611 = hbusreq5_p & v2302a8c | !hbusreq5_p & v84561b;
assign v23fc7ef = hlock0_p & v23fbd1a | !hlock0_p & v22f1e0b;
assign v23fc947 = hlock5_p & v23f1f1e | !hlock5_p & v2309c93;
assign v2311675 = hmaster2_p & v2304ad5 | !hmaster2_p & v2312c77;
assign v22ed8b5 = hmaster2_p & v23056b1 | !hmaster2_p & v230f848;
assign v22ed725 = hbusreq6_p & v2312e39 | !hbusreq6_p & v22fd32a;
assign v22f0ac0 = hlock0_p & v2307836 | !hlock0_p & v22fce06;
assign v2308a75 = hbusreq6 & v2305031 | !hbusreq6 & !v22fa68b;
assign v23fc940 = hmaster0_p & v23fce46 | !hmaster0_p & v23f62a3;
assign v22f2eaf = hbusreq3_p & v22ee95f | !hbusreq3_p & !v84561b;
assign v22f8d38 = hmaster2_p & v22fa70c | !hmaster2_p & v2391d40;
assign v23fccc1 = hbusreq4 & v23f6acc | !hbusreq4 & !v84562d;
assign v2391b6c = hmaster2_p & v84561b | !hmaster2_p & v23114d2;
assign v23f6659 = hmaster2_p & v23fbdb0 | !hmaster2_p & v23003cc;
assign v230890f = hgrant6_p & v84563a | !hgrant6_p & v2311a24;
assign v23fcc9f = hmaster2_p & b9d013 | !hmaster2_p & v12cd3f4;
assign v23fb1c8 = hgrant0_p & v23fbcb2 | !hgrant0_p & !v2313a33;
assign v22eda0b = hbusreq3 & v23fc633 | !hbusreq3 & v84561b;
assign v23f0206 = hbusreq4 & v230180d | !hbusreq4 & v23f729b;
assign v23f5686 = hmaster1_p & v230edc0 | !hmaster1_p & v22ec531;
assign v238ae11 = hbusreq0_p & a1fbb6 | !hbusreq0_p & a1fba6;
assign v22f7176 = stateA1_p & v84561b | !stateA1_p & !v22ec1cb;
assign v2309520 = hbusreq4_p & v230b5cc | !hbusreq4_p & v84561b;
assign v230180d = hmaster2_p & v22ed59e | !hmaster2_p & !v23fbedc;
assign v11853ca = jx0_p & v23f51a6 | !jx0_p & v22f6986;
assign v23fb727 = hbusreq6 & v23fc30b | !hbusreq6 & v22f6ed4;
assign v23078ff = hmaster2_p & v22f6a1b | !hmaster2_p & !v22fcbbb;
assign b5e598 = hlock2_p & v84561b | !hlock2_p & !v23068a9;
assign v230ed85 = hmaster2_p & v23f8f25 | !hmaster2_p & v22f8aec;
assign v22f1dab = hgrant0_p & v1506ea6 | !hgrant0_p & v230aec0;
assign v22f3d79 = hgrant3_p & a1fbc2 | !hgrant3_p & v230fb4c;
assign v2312846 = hmaster0_p & v22f58c2 | !hmaster0_p & v23003f5;
assign v22eb682 = hbusreq5 & v23041c3 | !hbusreq5 & v84561b;
assign v22f5125 = hbusreq3_p & bd74f4 | !hbusreq3_p & v23fcff6;
assign v23f4d86 = hbusreq4_p & v23f1faa | !hbusreq4_p & v239158e;
assign v239302b = hbusreq5_p & v22eb32b | !hbusreq5_p & v22f4d68;
assign v2300cf1 = hmaster2_p & v23f5043 | !hmaster2_p & v2301e25;
assign v23fc588 = jx1_p & v23fbcf0 | !jx1_p & v84561b;
assign v2302094 = hgrant3_p & v84561b | !hgrant3_p & v150708b;
assign v23f54de = hbusreq3_p & v22f728a | !hbusreq3_p & v230ce98;
assign v23f7d43 = hmaster2_p & v84564d | !hmaster2_p & v2300de3;
assign v15074fb = hbusreq2_p & v23fa1f4 | !hbusreq2_p & v84561b;
assign v23fc25b = hbusreq6_p & v22eaec3 | !hbusreq6_p & v22f0dd3;
assign v23fc3eb = hbusreq3 & v23013a6 | !hbusreq3 & v84561b;
assign v23fc88f = hbusreq6_p & v2301484 | !hbusreq6_p & v22f6fa9;
assign v23058ae = hbusreq5_p & v230230d | !hbusreq5_p & v84561b;
assign v23fc914 = hlock0_p & v22f56d2 | !hlock0_p & !v2302e32;
assign v23fbfe9 = hmaster0_p & v22fe2a8 | !hmaster0_p & v22f5353;
assign v15071c7 = hmaster2_p & v230d30a | !hmaster2_p & v23100c8;
assign v23fb67c = hlock0_p & v23f6077 | !hlock0_p & v22edb22;
assign v22f6e47 = hbusreq5_p & v23fbe41 | !hbusreq5_p & bd9ec5;
assign v2302365 = hbusreq3_p & v23fa492 | !hbusreq3_p & v84561b;
assign v22f4507 = hlock6_p & v22eba1d | !hlock6_p & !v84561b;
assign v23fb144 = hbusreq4_p & v2308f89 | !hbusreq4_p & v23fbe6e;
assign v22f03a0 = hmaster2_p & v230d814 | !hmaster2_p & v2309550;
assign v12cd903 = hbusreq3_p & v23faaa0 | !hbusreq3_p & v230859e;
assign v22fda63 = jx1_p & v23fbc89 | !jx1_p & v23f4e90;
assign v22f91b6 = hbusreq3_p & v22f5576 | !hbusreq3_p & v84564d;
assign v23fcb60 = hmaster0_p & v22fcc89 | !hmaster0_p & v230017e;
assign v230432b = hmaster0_p & v2391670 | !hmaster0_p & v230f0de;
assign v2303972 = hgrant2_p & v84561b | !hgrant2_p & e1df2d;
assign v23fbfba = hbusreq3 & v22f3dc7 | !hbusreq3 & !v23f8e04;
assign v963922 = hmaster2_p & v23fb6e3 | !hmaster2_p & v1506ffd;
assign v23fcd56 = hlock1_p & v23f7014 | !hlock1_p & v84564d;
assign v23f3eed = hbusreq5 & v23fc19d | !hbusreq5 & v84561b;
assign v23fc2db = hgrant1_p & v22f55fa | !hgrant1_p & v23fc316;
assign v8fac11 = hbusreq6_p & v22efd39 | !hbusreq6_p & v84561b;
assign v22ee91d = hbusreq6 & v23fbe6f | !hbusreq6 & !v23120a3;
assign v23fcecc = hmaster2_p & v230d709 | !hmaster2_p & v23fc2db;
assign bd9ec5 = stateG10_5_p & v23fcb53 | !stateG10_5_p & v23fbe41;
assign v23f0288 = hbusreq3_p & v94e407 | !hbusreq3_p & v23f62a8;
assign v23fb200 = hmaster2_p & v22fe32b | !hmaster2_p & v2301cc6;
assign v23fce72 = hgrant5_p & v84561b | !hgrant5_p & !v23037d2;
assign v22edb22 = hbusreq0_p & v23f6077 | !hbusreq0_p & v845620;
assign v22fd6d8 = hbusreq5_p & v230e07d | !hbusreq5_p & v23fcf98;
assign f40d2d = hgrant1_p & v23f4267 | !hgrant1_p & v23fc44c;
assign v23f96aa = hmaster2_p & v230031f | !hmaster2_p & v23f87f4;
assign v2308a71 = hgrant1_p & v2311810 | !hgrant1_p & v2312577;
assign v990272 = hlock4_p & v23fcfba | !hlock4_p & v239407e;
assign v23f38b1 = hbusreq4_p & v23f711a | !hbusreq4_p & !v84561b;
assign v23fbf9d = hbusreq0 & v22f60c6 | !hbusreq0 & v84564d;
assign v23fc17c = hmaster0_p & v15071c7 | !hmaster0_p & v23fb937;
assign v22f39d3 = hmaster2_p & v23fc38f | !hmaster2_p & v2303679;
assign v22edfa7 = hmaster2_p & v22f11f6 | !hmaster2_p & v2301505;
assign v230b5b8 = stateG10_5_p & a678c9 | !stateG10_5_p & v22f0945;
assign v22fb941 = hmaster0_p & v230b8fb | !hmaster0_p & v2305aa9;
assign v191ae4a = hmaster2_p & ae7427 | !hmaster2_p & v22f23a1;
assign v23f2713 = hbusreq1 & v23fcb5b | !hbusreq1 & v2391bc1;
assign v23fc741 = hgrant1_p & v22f4163 | !hgrant1_p & v230cef0;
assign v23f5deb = hbusreq6_p & v22f7d00 | !hbusreq6_p & v23f4f2c;
assign v23f1b7a = hbusreq4_p & v23fbae0 | !hbusreq4_p & bd7ae5;
assign v230e78c = locked_p & v23fc53e | !locked_p & v84561b;
assign v230c55d = hgrant1_p & v84561b | !hgrant1_p & !v2391f87;
assign v22f6fb8 = hbusreq5_p & v23fc3cb | !hbusreq5_p & v2304883;
assign v22f5a08 = hgrant5_p & v22fe6c8 | !hgrant5_p & v23fbb8b;
assign v22ebb85 = hmaster2_p & v230913d | !hmaster2_p & !v84561b;
assign v230ce2b = hlock6_p & v23f6b18 | !hlock6_p & !v84561b;
assign v22f3aac = hmaster2_p & b50a75 | !hmaster2_p & v9c1abc;
assign v22f865d = hbusreq3_p & v2304fc6 | !hbusreq3_p & v22f83fb;
assign v23fb97c = hgrant3_p & v23fc139 | !hgrant3_p & !v23f67fe;
assign v22f3d00 = hbusreq1_p & v23faa23 | !hbusreq1_p & v84561b;
assign v230ec39 = hbusreq3_p & v23f7254 | !hbusreq3_p & v22f7da7;
assign v22f5243 = hbusreq5 & v230be24 | !hbusreq5 & b9c9ef;
assign v23fc6a0 = hgrant1_p & v231022d | !hgrant1_p & v23fc3fb;
assign v230cf9a = hgrant6_p & v2304da3 | !hgrant6_p & !v191abf8;
assign v191ae51 = hmaster2_p & b09503 | !hmaster2_p & v2311918;
assign v22f1681 = hbusreq2_p & v22fe46b | !hbusreq2_p & v845620;
assign v2310c98 = hlock6_p & v23f3c98 | !hlock6_p & v230f8f4;
assign v22fca3a = hbusreq4_p & v150744b | !hbusreq4_p & v22ed1d3;
assign v22f49ac = hbusreq5_p & v23f301a | !hbusreq5_p & v23fc811;
assign v23030ad = hmaster2_p & v230c8e9 | !hmaster2_p & v22ef062;
assign v230e71c = hbusreq2_p & v23fc250 | !hbusreq2_p & v84561b;
assign v23fbf87 = hlock5_p & v22f037a | !hlock5_p & !v84561b;
assign v23fc9eb = jx0_p & v23104db | !jx0_p & !v23fc628;
assign v22f7b83 = hbusreq1 & v23f9789 | !hbusreq1 & v22f0945;
assign v23082c9 = hmaster1_p & v23fbf13 | !hmaster1_p & v191b038;
assign v23fb384 = hbusreq6_p & v23f4160 | !hbusreq6_p & v2311011;
assign v22fb7a5 = hbusreq2 & v23f1207 | !hbusreq2 & f40cd3;
assign v2312d20 = hbusreq5 & v23fc9d2 | !hbusreq5 & v84561b;
assign v22ec8dc = hmaster0_p & v22ff30c | !hmaster0_p & v23fb954;
assign v22f852d = hgrant0_p & v23f20d7 | !hgrant0_p & v23f89db;
assign v22f5019 = hlock4_p & v22f87bf | !hlock4_p & v84561b;
assign a1b802 = hbusreq1 & v845620 | !hbusreq1 & v2303075;
assign v23047e5 = hbusreq3_p & v22f515e | !hbusreq3_p & v1aae12f;
assign v230ec1c = hmaster2_p & v23f3206 | !hmaster2_p & a6b8e0;
assign v23fc548 = jx0_p & v84561b | !jx0_p & !v23fbe1f;
assign fc8c53 = hmaster0_p & v2304a06 | !hmaster0_p & !v230e75b;
assign v23f94e5 = hbusreq5 & v22f442c | !hbusreq5 & !v84561b;
assign v22f065f = hbusreq3_p & da38c1 | !hbusreq3_p & v230052f;
assign v22f2e64 = stateG10_5_p & v22f4d04 | !stateG10_5_p & v22fe097;
assign v91ff8a = hmaster2_p & da38c1 | !hmaster2_p & v23f468c;
assign bd7a62 = hbusreq3 & b00aa0 | !hbusreq3 & v845625;
assign v23086b9 = hmaster2_p & v22fb77d | !hmaster2_p & v84561b;
assign v22fc13d = hbusreq1_p & v23f60ef | !hbusreq1_p & v22ef816;
assign v22ee4eb = hbusreq6_p & v23fcd42 | !hbusreq6_p & v230cfb5;
assign v230851f = hbusreq6 & v23f7cea | !hbusreq6 & v23fba11;
assign v2304118 = hlock3_p & a1ff0e | !hlock3_p & !v106ae19;
assign v23fc1db = hbusreq6_p & v2309459 | !hbusreq6_p & v23109c8;
assign v2312524 = hmaster1_p & v22f7fd1 | !hmaster1_p & v23f34d7;
assign v23f910c = hbusreq1 & v2305811 | !hbusreq1 & v84561b;
assign v21eabbd = hgrant2_p & v84561b | !hgrant2_p & v845629;
assign v239268e = hbusreq4_p & v2392697 | !hbusreq4_p & v231171e;
assign v23f4634 = hgrant5_p & v23fcfd6 | !hgrant5_p & v22fcf71;
assign v933ab1 = hmaster0_p & v22f87a1 | !hmaster0_p & !v230cdc1;
assign v191afb7 = hmaster0_p & v23f7039 | !hmaster0_p & !v23fc7a6;
assign v23fc44d = hbusreq4 & v2307c44 | !hbusreq4 & v230c4ae;
assign v1e840f2 = hmaster2_p & v23fbfce | !hmaster2_p & v23fc9d1;
assign v22fce2e = hbusreq6 & v22f99e3 | !hbusreq6 & v23002bf;
assign v845626 = hbusreq1 & v84561b | !hbusreq1 & !v84561b;
assign v22f31b9 = hmaster2_p & v2305b35 | !hmaster2_p & v230c2f4;
assign v23fade4 = hmaster2_p & v22f7b29 | !hmaster2_p & v2304deb;
assign v23108b7 = hlock0_p & v23fbaae | !hlock0_p & !a1fde3;
assign v23f316e = hgrant2_p & v23fc29c | !hgrant2_p & !v84561b;
assign b9d00f = hmastlock_p & v22f37ba | !hmastlock_p & v84561b;
assign v23fbfce = hbusreq1_p & v22fa70c | !hbusreq1_p & v22f78ee;
assign v2307309 = hgrant3_p & v2300f82 | !hgrant3_p & v23f5f18;
assign v22faa42 = jx0_p & v230ed07 | !jx0_p & !v23f64d3;
assign v22fcab7 = hbusreq6_p & v2302875 | !hbusreq6_p & v23f67fa;
assign b30f07 = hgrant5_p & v84561b | !hgrant5_p & v22f8fc0;
assign v2309057 = hmaster2_p & v23056b1 | !hmaster2_p & v106ae19;
assign v2382e8c = hmaster2_p & v23f6411 | !hmaster2_p & b5f51c;
assign v22ffea8 = hgrant3_p & v84561b | !hgrant3_p & v23f5c89;
assign v22ee75e = hgrant3_p & v23fc854 | !hgrant3_p & v22f865d;
assign v22ffcb8 = hbusreq1_p & v230bd05 | !hbusreq1_p & v23071f6;
assign v22f5583 = hlock0_p & v23fbb35 | !hlock0_p & v23f4b28;
assign v230e295 = hbusreq0_p & v22ed85a | !hbusreq0_p & v23fbdb0;
assign v230fe99 = hbusreq6 & v106af1c | !hbusreq6 & !v84561b;
assign v23fd01b = hlock1_p & v22f3a35 | !hlock1_p & !v106ae19;
assign v23f965d = hmaster0_p & v84564d | !hmaster0_p & v2302131;
assign v23131e8 = hmastlock_p & v23fba3a | !hmastlock_p & v84561b;
assign v22f73a3 = hmaster2_p & v23fc982 | !hmaster2_p & v23f76d0;
assign a1fbcb = hlock1_p & v23fcf96 | !hlock1_p & !v84561b;
assign v2304b35 = hbusreq1_p & bd7c9b | !hbusreq1_p & v84561b;
assign v22eb66f = hbusreq0_p & v23fc2fc | !hbusreq0_p & v84561b;
assign v23fcb0b = hgrant2_p & v84562a | !hgrant2_p & !v84561b;
assign v23f6f49 = hlock3_p & v2302365 | !hlock3_p & v23fb4a1;
assign v22ff120 = hgrant1_p & v230eb9b | !hgrant1_p & adb81d;
assign v23f88a9 = hmaster2_p & v84561b | !hmaster2_p & !v22f0add;
assign v23fa3b8 = hbusreq6 & v2312999 | !hbusreq6 & v84561b;
assign v23fca5c = hmaster0_p & v23f350b | !hmaster0_p & v22ecdde;
assign v22fbf38 = hgrant3_p & v84561b | !hgrant3_p & v23fbf07;
assign v22fe84a = hmaster0_p & v23fc3e8 | !hmaster0_p & v22f1d1f;
assign v23fc44c = hbusreq1_p & v2309b3e | !hbusreq1_p & v12cd920;
assign v230296a = hbusreq4_p & v22fdf70 | !hbusreq4_p & v23f2d60;
assign v2310047 = jx0_p & v23fbb85 | !jx0_p & v22f23e6;
assign v23126be = hgrant1_p & v23fce3b | !hgrant1_p & !v84561b;
assign v23fc11e = hbusreq2_p & v15072de | !hbusreq2_p & !v84562a;
assign v22f53e2 = hbusreq3_p & v23fc0e0 | !hbusreq3_p & v22fa857;
assign v23f9b49 = hlock3_p & v230a0d1 | !hlock3_p & !v23f7e3d;
assign v23fbeeb = hbusreq3_p & v845622 | !hbusreq3_p & v230fc56;
assign v22fe32b = hgrant1_p & v230f933 | !hgrant1_p & v22f94b6;
assign v22f5753 = hbusreq4 & v23fbff6 | !hbusreq4 & v22fd314;
assign v23efd4b = hbusreq6_p & v22fd48a | !hbusreq6_p & v2311e38;
assign v23fbf8d = hgrant3_p & v84561b | !hgrant3_p & v23fbdc1;
assign v23087d7 = hmaster2_p & v1aad5ad | !hmaster2_p & v84561b;
assign v2306eb5 = hbusreq3_p & v2307f3f | !hbusreq3_p & v84561b;
assign a9176f = hlock6_p & b59af9 | !hlock6_p & v23fc885;
assign v23fca56 = hbusreq1 & v23fc23d | !hbusreq1 & v84561b;
assign v23f20e8 = hmaster0_p & v23fc5dd | !hmaster0_p & v230d2a3;
assign v22f8420 = hmaster2_p & v230945e | !hmaster2_p & v22ee956;
assign v22fa27c = hbusreq6 & v23fc72d | !hbusreq6 & v84561b;
assign v15072a9 = hgrant1_p & v84561b | !hgrant1_p & v23fcdd7;
assign b13467 = hgrant5_p & v22f358f | !hgrant5_p & !v84561b;
assign v23fba81 = hlock3_p & v23fb41a | !hlock3_p & !v84561b;
assign v2310475 = hlock5_p & b62970 | !hlock5_p & v22f9567;
assign dab2cc = hbusreq6 & v23f6478 | !hbusreq6 & v84561b;
assign v230fd1c = hbusreq3_p & v23f3346 | !hbusreq3_p & v22f7ed8;
assign v22fbf28 = hbusreq3 & v191b041 | !hbusreq3 & v84561b;
assign v2313351 = hmaster2_p & v22fbd02 | !hmaster2_p & v845620;
assign v230e0d5 = hbusreq2 & v22ed878 | !hbusreq2 & v84561b;
assign v23fc0c1 = hmaster0_p & v2304189 | !hmaster0_p & v23fbdfc;
assign v2310291 = jx1_p & v22fa61c | !jx1_p & v22f1a0e;
assign v22febdb = hready_p & v23f960d | !hready_p & v23fc8ce;
assign v23f4e43 = hlock1_p & v22f037a | !hlock1_p & !v84561b;
assign v22f814a = hlock2_p & v191a876 | !hlock2_p & v84561b;
assign v23fb1a1 = hbusreq3_p & v230d134 | !hbusreq3_p & v23fb77d;
assign v230eb13 = hmastlock_p & v23f707f | !hmastlock_p & v84565f;
assign v23f8561 = hlock1_p & v22ff414 | !hlock1_p & !v84561b;
assign v23fbade = hlock0_p & v22ecee2 | !hlock0_p & v23fba4f;
assign v230e94e = hmaster1_p & v22ed725 | !hmaster1_p & v23fc2ff;
assign v23fc460 = hbusreq3_p & v22f069f | !hbusreq3_p & !v23fc6e5;
assign v230320e = hlock0_p & v2306d29 | !hlock0_p & v22f5e8c;
assign v22f90c3 = hbusreq3_p & v22f1754 | !hbusreq3_p & v84561b;
assign v23f06a5 = hmaster0_p & v23f6326 | !hmaster0_p & v23fc630;
assign v22f856d = hbusreq4_p & v23f62c2 | !hbusreq4_p & v23fcfce;
assign v23f5ab1 = busreq_p & a72160 | !busreq_p & v84561b;
assign v2301ad7 = hbusreq1 & v13afe3a | !hbusreq1 & !b00ad3;
assign v13afb01 = stateG10_5_p & v2305979 | !stateG10_5_p & !v23f39e5;
assign v230e628 = hlock6_p & v23f4d86 | !hlock6_p & v84561b;
assign v22f06fb = hgrant5_p & v84561b | !hgrant5_p & a1bfd6;
assign v1aad4fc = hbusreq5 & v13afe3a | !hbusreq5 & !b00ad3;
assign v22ef513 = hmastlock_p & v22ed458 | !hmastlock_p & !v84561b;
assign v2303a53 = hgrant3_p & a1fbc2 | !hgrant3_p & v2302353;
assign v23f6ace = jx1_p & v23fb196 | !jx1_p & v2305b5a;
assign fc8f95 = hmaster2_p & v2309dc4 | !hmaster2_p & v23fcdbe;
assign v22fea89 = hgrant0_p & v845622 | !hgrant0_p & v22fb727;
assign v22fe382 = hbusreq3_p & v22f6e30 | !hbusreq3_p & v23056bf;
assign v22ffc85 = hready_p & v230890f | !hready_p & !v230524c;
assign v23fb798 = hbusreq5 & v13afe3a | !hbusreq5 & v84561b;
assign v22f43ec = jx0_p & v23f9bcc | !jx0_p & !v22ecea2;
assign v2311668 = hgrant3_p & v22f2db6 | !hgrant3_p & !v84561b;
assign v23fa997 = hgrant5_p & v84561b | !hgrant5_p & v23058ae;
assign v22f2d35 = hbusreq3_p & v22edadc | !hbusreq3_p & v230361d;
assign v23f3ab0 = hmaster2_p & v22f954f | !hmaster2_p & a88394;
assign v2391c8a = hbusreq5_p & v230fec6 | !hbusreq5_p & v23f3e19;
assign v23fc1fa = hbusreq3_p & v23f1387 | !hbusreq3_p & !v84561b;
assign v2304299 = hbusreq5_p & v23f5cb3 | !hbusreq5_p & !v2301709;
assign v23fc5ea = jx0_p & v23049af | !jx0_p & v2301972;
assign v230cbde = stateG10_5_p & v230bc8b | !stateG10_5_p & v84564d;
assign v2309e57 = hbusreq3_p & v13afb18 | !hbusreq3_p & v2304bc1;
assign v23f21cf = hmaster2_p & v84561b | !hmaster2_p & !v22faa21;
assign v2305d15 = hbusreq5_p & v22fbf74 | !hbusreq5_p & v2302386;
assign a5a279 = hgrant5_p & v2311506 | !hgrant5_p & v22f41ee;
assign v23f2216 = hburst0_p & v84561b | !hburst0_p & v23fc8d7;
assign b00a55 = hmaster0_p & v2307fd0 | !hmaster0_p & v22fd048;
assign v230c469 = hbusreq5_p & v22f0945 | !hbusreq5_p & v84561b;
assign v23f40fd = hgrant3_p & v2311e03 | !hgrant3_p & v23fb672;
assign v230b23b = hbusreq5_p & v84564d | !hbusreq5_p & v230cbde;
assign v23fbe18 = hbusreq3_p & v23110a4 | !hbusreq3_p & v230cbf6;
assign v23f50dd = hbusreq4_p & v23fb86a | !hbusreq4_p & v22f9c34;
assign v22f0870 = hgrant1_p & v84561b | !hgrant1_p & v23022c5;
assign v230817b = hbusreq6_p & v22f6d6e | !hbusreq6_p & v22fae03;
assign v23fb1ca = hlock3_p & v2306d47 | !hlock3_p & v230a6ed;
assign v22f0210 = hmaster0_p & v22ffd0e | !hmaster0_p & v22f670f;
assign v22f7d5c = hmaster1_p & v23028fa | !hmaster1_p & v23115f8;
assign v22fca63 = hmaster1_p & v23f9bd1 | !hmaster1_p & v2393f3f;
assign v22ff66a = hmaster0_p & v23f7637 | !hmaster0_p & v23fb9e7;
assign v23fbce6 = hmaster2_p & v22f068b | !hmaster2_p & v22fe343;
assign v23fc69b = hmaster2_p & v22f337b | !hmaster2_p & v23f2be7;
assign v23fbbee = stateG10_5_p & v2302075 | !stateG10_5_p & !v84561b;
assign v23fc410 = hbusreq6 & v23f9aa8 | !hbusreq6 & v2310d04;
assign v230880f = hmaster2_p & v22ef403 | !hmaster2_p & v22f0593;
assign v23f193e = hgrant3_p & v84562e | !hgrant3_p & v23fbe95;
assign v2392254 = hgrant3_p & v230d4cc | !hgrant3_p & v23fc71a;
assign v23027f9 = hbusreq3_p & v23fcbdb | !hbusreq3_p & v230fb43;
assign v2391728 = hgrant5_p & v22ed48c | !hgrant5_p & v84561b;
assign v23fcabb = hbusreq0_p & afc788 | !hbusreq0_p & v845620;
assign v230e449 = hbusreq6_p & v2309ffa | !hbusreq6_p & v230d6b2;
assign v2303314 = hmaster0_p & v230d96b | !hmaster0_p & v23fbb4a;
assign b7b244 = hbusreq5_p & v2391d40 | !hbusreq5_p & v8d030a;
assign v23fbf5f = hbusreq5 & v23f6b25 | !hbusreq5 & v84561b;
assign v22fa2de = locked_p & v230a3ec | !locked_p & v84561b;
assign v22f20df = hbusreq3 & v23f5a39 | !hbusreq3 & !v84561b;
assign v23fcab0 = hbusreq0 & v84561b | !hbusreq0 & !v84564d;
assign v230beb6 = hbusreq2_p & v106ae4a | !hbusreq2_p & a1fba6;
assign v22f2bf1 = hbusreq6 & v2306405 | !hbusreq6 & !v84562a;
assign v23fc72d = hmaster2_p & v2312580 | !hmaster2_p & v84561b;
assign v23f8a5e = hlock4_p & v2301b38 | !hlock4_p & v84561b;
assign v23124aa = hbusreq3_p & v22fdbbe | !hbusreq3_p & v23fb550;
assign v22fa36f = hbusreq6 & v23f2873 | !hbusreq6 & v22f8ba5;
assign a507a6 = hbusreq4 & v22f7793 | !hbusreq4 & v84561b;
assign v230a25a = hgrant5_p & v22ffba8 | !hgrant5_p & v2393c3a;
assign v2307ff9 = hlock2_p & e1df2d | !hlock2_p & v84561b;
assign a1f79d = decide_p & v23f8fd7 | !decide_p & v230e312;
assign v230f9c2 = hmaster2_p & v1e84174 | !hmaster2_p & v230ce60;
assign v23fb4cf = hmaster2_p & v84561b | !hmaster2_p & !v23f7789;
assign v23fbe4d = hbusreq5_p & v84561b | !hbusreq5_p & !v230feb2;
assign v22f2ce7 = hmaster1_p & v230c155 | !hmaster1_p & v23fcf6a;
assign v23fb920 = locked_p & b9d00f | !locked_p & !v2309c8a;
assign v23ef951 = hbusreq3 & v22eefcf | !hbusreq3 & v23f4827;
assign v2391670 = hgrant3_p & v84562e | !hgrant3_p & v22fb9eb;
assign v2309c1f = hmaster2_p & v22f7da7 | !hmaster2_p & v84561b;
assign v23925af = hgrant0_p & v230fec6 | !hgrant0_p & !v22f1000;
assign v22f0aea = hbusreq3_p & v2393064 | !hbusreq3_p & v22f6719;
assign v23f7637 = hgrant3_p & v2308af4 | !hgrant3_p & v23f79a7;
assign v231363a = hbusreq3_p & v22fa851 | !hbusreq3_p & v84561b;
assign v22fd781 = hbusreq2 & v22f9911 | !hbusreq2 & v230f5a3;
assign v22f5e59 = hbusreq1_p & v23070c1 | !hbusreq1_p & !v22fa870;
assign v2308e85 = hbusreq1 & v2307150 | !hbusreq1 & v84561b;
assign v23f5d72 = hbusreq2_p & v2391a57 | !hbusreq2_p & !v84561b;
assign v230f8f4 = hmaster0_p & baa026 | !hmaster0_p & !v2305cac;
assign v230d4cc = hbusreq3_p & v23f558b | !hbusreq3_p & v22fe0b0;
assign v2307725 = hbusreq5 & v230446f | !hbusreq5 & !v84562a;
assign v23fc8ea = hgrant5_p & v23f520c | !hgrant5_p & !v12cda57;
assign v23fa823 = hmaster0_p & v84561b | !hmaster0_p & v22ffaef;
assign v23f6ec1 = hlock1_p & v230894d | !hlock1_p & v2304bc1;
assign v23f9f77 = hbusreq1_p & v22ffb2b | !hbusreq1_p & v84561b;
assign v23fc7d1 = hmaster2_p & b9d013 | !hmaster2_p & !v2304deb;
assign v22f595b = hmaster2_p & v23f2d28 | !hmaster2_p & v22f61b6;
assign v231160e = hgrant5_p & v23fb4fd | !hgrant5_p & v230f485;
assign v230c2c5 = hbusreq4_p & v230c439 | !hbusreq4_p & v23115f4;
assign v22fcad1 = hmaster2_p & fc8c68 | !hmaster2_p & !v84561b;
assign v230de82 = hbusreq6_p & v23fb701 | !hbusreq6_p & v23f36a3;
assign v22ed756 = hgrant3_p & v84562e | !hgrant3_p & v22f1f3f;
assign v22ebc28 = hbusreq4_p & v2311df1 | !hbusreq4_p & v23f1561;
assign v22efd4d = hmaster2_p & v22f7da7 | !hmaster2_p & v23fb5a1;
assign v23fbed5 = hgrant1_p & v845620 | !hgrant1_p & f40a9e;
assign v230ebff = hbusreq5 & v84561b | !hbusreq5 & !v22ef725;
assign v23f4b28 = hbusreq0_p & v23fbb35 | !hbusreq0_p & v84561b;
assign v23f0db6 = hmaster1_p & v22ef55f | !hmaster1_p & v23fccc5;
assign v1aaddfe = hbusreq6_p & a28a9e | !hbusreq6_p & v84561b;
assign v22f993e = hmaster2_p & v22fe5b1 | !hmaster2_p & v22f5037;
assign v2302c31 = hgrant6_p & v84561b | !hgrant6_p & !v845657;
assign v22ebc26 = hbusreq4_p & v22fe76b | !hbusreq4_p & v23fa2b8;
assign v23f40ab = hbusreq1 & v22f9911 | !hbusreq1 & v84561b;
assign v230a92e = hbusreq5_p & v2303fb9 | !hbusreq5_p & v84561b;
assign v23094a1 = hmaster1_p & v230b1a3 | !hmaster1_p & v2309ae3;
assign v22ee0d5 = hbusreq3_p & v23018a8 | !hbusreq3_p & v22ec3c3;
assign v9bd8c6 = hburst0 & v22f3294 | !hburst0 & v23fc116;
assign v23f7393 = hmaster0_p & v2391d2f | !hmaster0_p & v23fb6b5;
assign v23f3dcc = hmaster2_p & v106ae21 | !hmaster2_p & v2307150;
assign v23f5ef2 = hbusreq3 & v22f0945 | !hbusreq3 & v23f2d33;
assign v23fd05d = hmaster2_p & v23fa2ec | !hmaster2_p & v2301511;
assign v22ed933 = hmaster0_p & b9c985 | !hmaster0_p & !v22eb933;
assign v23fca78 = hbusreq3_p & v23f7d9f | !hbusreq3_p & v22ebd88;
assign e1e73c = hlock0_p & v23fb9b2 | !hlock0_p & !v84561b;
assign v2309939 = hlock0_p & v22f7928 | !hlock0_p & v22ec88f;
assign v23fbbf6 = hbusreq2_p & v2309a44 | !hbusreq2_p & v2313463;
assign v22ec64d = hbusreq6 & v23fcca1 | !hbusreq6 & v84561b;
assign v22f9f44 = stateG10_5_p & v22f05a9 | !stateG10_5_p & v22ec801;
assign v13afebe = hlock0_p & v22f1a26 | !hlock0_p & v23f3715;
assign v23fc303 = hbusreq2 & v22f1389 | !hbusreq2 & v84561b;
assign v23f37c6 = hbusreq2_p & v23f5043 | !hbusreq2_p & !v845620;
assign v22f995e = hgrant1_p & v23f6d19 | !hgrant1_p & v23111da;
assign v22ee4d5 = hbusreq3_p & v22ec060 | !hbusreq3_p & v845620;
assign v23928ae = hlock3_p & v22f6759 | !hlock3_p & v2307dfb;
assign v23f9fb5 = hmaster2_p & v84561b | !hmaster2_p & fc8e3a;
assign v23f940c = hbusreq1_p & v22ff45e | !hbusreq1_p & v84561b;
assign v22f2453 = hgrant0_p & v2307e48 | !hgrant0_p & v84561b;
assign v230996e = hmaster0_p & v23fcaa5 | !hmaster0_p & v23fbf8d;
assign v230cb0f = hbusreq3_p & bd7a67 | !hbusreq3_p & v230ed08;
assign v230e579 = hbusreq1 & v23f65b4 | !hbusreq1 & !v22ee7a7;
assign v23f51e3 = hgrant1_p & v84561b | !hgrant1_p & v22efb46;
assign v22ed928 = hmaster0_p & v1507157 | !hmaster0_p & !v96c563;
assign v22f049f = hbusreq5_p & v2311dcb | !hbusreq5_p & v2305799;
assign v2307e48 = locked_p & v23fb95d | !locked_p & v84561b;
assign v23f895d = hbusreq3_p & v23fc549 | !hbusreq3_p & v84561b;
assign v23fc209 = hbusreq5_p & v23f11a3 | !hbusreq5_p & v22ed1e8;
assign v22ee0c9 = hmaster1_p & v23fb5f1 | !hmaster1_p & !v2391e8e;
assign v22eb415 = hgrant1_p & v22ede4d | !hgrant1_p & v84561b;
assign v23f593d = hmaster0_p & v23107f0 | !hmaster0_p & v23f403e;
assign b159aa = hgrant2_p & v230219b | !hgrant2_p & v22f7f74;
assign v23fd050 = hbusreq2_p & v22fd86e | !hbusreq2_p & v84561b;
assign v2305866 = hmaster0_p & v2305bf5 | !hmaster0_p & v23f4a48;
assign b9c8ff = hmaster2_p & v23fcfb8 | !hmaster2_p & v22fc091;
assign v231339c = hbusreq0 & v23f8f21 | !hbusreq0 & !v23fbbd2;
assign v2391c72 = hbusreq5_p & v23fbd26 | !hbusreq5_p & !v23fbee6;
assign v22ec477 = hbusreq1_p & v106af73 | !hbusreq1_p & v191a879;
assign v22ed458 = stateG2_p & v84561b | !stateG2_p & !v230b364;
assign v22eea17 = hbusreq1 & v23f1207 | !hbusreq1 & v230b1ac;
assign v2308e0b = hgrant3_p & v84562e | !hgrant3_p & v23fc993;
assign v230a42d = stateG10_5_p & v23fc153 | !stateG10_5_p & v84562b;
assign v9932c2 = hlock5_p & v2313463 | !hlock5_p & !v84561b;
assign v23f07f9 = hbusreq3_p & v22f8477 | !hbusreq3_p & v2307e4c;
assign v85fc1a = hmaster1_p & v23fb724 | !hmaster1_p & v84562d;
assign v230d00c = hgrant3_p & v23fa94e | !hgrant3_p & v22f0b8a;
assign v23fc627 = hbusreq3_p & v2310e5d | !hbusreq3_p & !v84561b;
assign v22fd8fc = hbusreq1_p & v23fc39c | !hbusreq1_p & b30f07;
assign v231007d = hbusreq5_p & v22f0824 | !hbusreq5_p & v22f383e;
assign v22f84f8 = hbusreq6 & v22f4a40 | !hbusreq6 & v84561b;
assign v23fb70e = hbusreq6_p & v23fb139 | !hbusreq6_p & !v23f60ba;
assign v230f947 = hbusreq0 & v2303831 | !hbusreq0 & !v22f0860;
assign v23f06c9 = hbusreq6_p & v22f6e51 | !hbusreq6_p & v23fc296;
assign v23f6155 = hgrant5_p & v230edde | !hgrant5_p & v22ed984;
assign v22fd271 = hgrant5_p & v23fc512 | !hgrant5_p & v845635;
assign v2309ba2 = hbusreq5 & v23faf60 | !hbusreq5 & !v84561b;
assign v23107f5 = hbusreq6 & v22f3dc7 | !hbusreq6 & !v23f8e04;
assign v23fcea8 = hlock5_p & v845636 | !hlock5_p & !v84561b;
assign v2308af4 = hlock3_p & v23fbf12 | !hlock3_p & v2309c93;
assign v23fc904 = hlock0_p & v2306d29 | !hlock0_p & v22ef05d;
assign v1aae9a1 = hmaster2_p & v2302a4d | !hmaster2_p & !v22ffc69;
assign v23fb8c1 = hbusreq5_p & v23fb122 | !hbusreq5_p & v23f22a1;
assign v23fb0c9 = hgrant5_p & v84561b | !hgrant5_p & !v84564f;
assign v22f9894 = hbusreq0 & v22f337b | !hbusreq0 & v845620;
assign v90b913 = hbusreq1 & v23fc89a | !hbusreq1 & !v845622;
assign v22efeed = hgrant0_p & v22ffb9d | !hgrant0_p & !v23064ae;
assign v23fcc5e = hmaster1_p & v230695e | !hmaster1_p & v23fa3bb;
assign v230fb4c = hmaster2_p & v230313a | !hmaster2_p & v22fe204;
assign v2301567 = jx0_p & v23fba6a | !jx0_p & v231142b;
assign v23f626c = hmaster2_p & v22ed59e | !hmaster2_p & !v22f8bd0;
assign v23fa75a = hlock0_p & v230219b | !hlock0_p & v22f7f74;
assign v230afed = hgrant3_p & e1e258 | !hgrant3_p & v23fbeb5;
assign v23fc5ac = hbusreq6_p & v22f1744 | !hbusreq6_p & v23fb886;
assign v22fc37d = hmaster2_p & b9d013 | !hmaster2_p & v230f848;
assign v23fb0c0 = hmaster2_p & v2300827 | !hmaster2_p & v22ff5af;
assign v23fc58e = hgrant1_p & v84561b | !hgrant1_p & v23fbb89;
assign v2300f25 = hmaster2_p & v22ff043 | !hmaster2_p & v23fbedc;
assign v230a58e = hbusreq5_p & v230848d | !hbusreq5_p & v2310476;
assign v23fc362 = hgrant1_p & v106af73 | !hgrant1_p & v22f6d58;
assign v23057f1 = hmaster1_p & v230fd86 | !hmaster1_p & v191b085;
assign c173c8 = hmaster2_p & b6f86d | !hmaster2_p & v22f98fd;
assign v230dd15 = hgrant3_p & v22f8e29 | !hgrant3_p & v1e840d4;
assign v22eb38b = hmaster0_p & v2312a18 | !hmaster0_p & v94508c;
assign v87cfb8 = hbusreq0_p & v230446f | !hbusreq0_p & !v2301655;
assign v22f0d2b = hbusreq1_p & v23001a4 | !hbusreq1_p & v22f3b3c;
assign v23fc066 = hbusreq5 & v23f95e1 | !hbusreq5 & v22ecee2;
assign v23fbf49 = hgrant3_p & v23fbea6 | !hgrant3_p & v23008c7;
assign hmastlock = v17a2d5b;
assign v23fb18d = hmaster2_p & v23f80c1 | !hmaster2_p & v22fca28;
assign v23fc5d0 = hbusreq3 & v23fc4d0 | !hbusreq3 & v23051cf;
assign v22ee09a = hbusreq3_p & v22f7dbc | !hbusreq3_p & !v22f7ec9;
assign v23faede = hbusreq3_p & v22f2bab | !hbusreq3_p & v23fc162;
assign v22ed925 = hbusreq3_p & v23059ee | !hbusreq3_p & v23fc030;
assign v2312948 = hmaster2_p & v22ebbf1 | !hmaster2_p & v22ed10d;
assign v22ecba3 = hgrant1_p & v231128c | !hgrant1_p & v2310f46;
assign v22f383c = hgrant3_p & v23f5ace | !hgrant3_p & v22f4d97;
assign v23f8866 = hbusreq4_p & v23f1688 | !hbusreq4_p & v23fb604;
assign v22f1ca0 = locked_p & v230f776 | !locked_p & v84561b;
assign v22ffb6b = hgrant1_p & v845635 | !hgrant1_p & v22fd271;
assign v23049ad = hbusreq6 & v22f20b4 | !hbusreq6 & v84561b;
assign v22ed942 = hbusreq3_p & v22ec2a4 | !hbusreq3_p & v84561b;
assign v230b12a = stateG10_5_p & v22f6a0e | !stateG10_5_p & a1fbc2;
assign v22f39f4 = hgrant3_p & v106ae8b | !hgrant3_p & v23f60fb;
assign v23f450d = hgrant0_p & v84561b | !hgrant0_p & v23fb567;
assign v23026f7 = hmaster2_p & v84561b | !hmaster2_p & !v22ec753;
assign v23f301a = hlock0_p & v23f7789 | !hlock0_p & !v84561b;
assign b9c90c = hgrant3_p & v23fb937 | !hgrant3_p & v23f9ba6;
assign a5666b = hmaster2_p & v845661 | !hmaster2_p & v2304b4e;
assign v22f16bf = hmaster2_p & v23f55ea | !hmaster2_p & !v22fa870;
assign v10dbf78 = hready_p & v23f193c | !hready_p & v845643;
assign e1e250 = hgrant1_p & v22f65b7 | !hgrant1_p & v9ec6b5;
assign v23fc1ee = hbusreq1 & v22ed267 | !hbusreq1 & v84561b;
assign v22eb8ad = hmaster2_p & v97b973 | !hmaster2_p & !v23930d2;
assign v23f64e5 = hbusreq0_p & v23f51b1 | !hbusreq0_p & !b9d013;
assign v22f5fb4 = hbusreq3_p & v845627 | !hbusreq3_p & b50a75;
assign v230994d = hbusreq4_p & v23f8fd0 | !hbusreq4_p & v22f0284;
assign v2309fb1 = hbusreq1 & v230e916 | !hbusreq1 & v23f87f4;
assign v22ee9c4 = hbusreq2 & v13afe3a | !hbusreq2 & !fc8ab7;
assign v22fb00c = hmaster2_p & bc96dd | !hmaster2_p & v22f1d80;
assign v9bbf5d = hmaster2_p & v22f8b01 | !hmaster2_p & v23080ec;
assign v23fc7c0 = hlock3_p & v22f2718 | !hlock3_p & !v84561b;
assign v22eb12e = hbusreq4_p & v23039ea | !hbusreq4_p & v22f1d05;
assign v23fb926 = hbusreq6 & v23fcba1 | !hbusreq6 & v84561b;
assign v22fdad1 = hbusreq4_p & v22fb442 | !hbusreq4_p & v23fc5b3;
assign v2311d05 = hbusreq6_p & v230b0f2 | !hbusreq6_p & v2307eac;
assign v23f7370 = hgrant1_p & v84561b | !hgrant1_p & v2391f85;
assign v23058b0 = hbusreq6_p & v23fbdd2 | !hbusreq6_p & v23fa2b8;
assign v2305c24 = hbusreq1_p & v9526ac | !hbusreq1_p & a1fba6;
assign v23f6b0f = stateG10_5_p & v23f8176 | !stateG10_5_p & !v12cd3f4;
assign v2391bc1 = hbusreq2_p & v2309310 | !hbusreq2_p & v84561b;
assign v1aacf10 = decide_p & v2310537 | !decide_p & v84564d;
assign v230011a = hbusreq5 & v2312fc7 | !hbusreq5 & v84561b;
assign v23f1a83 = jx0_p & v23047dd | !jx0_p & v2312397;
assign v23080f9 = hbusreq4 & v23fcd7f | !hbusreq4 & v84561b;
assign v23fbae2 = hbusreq2 & v23f2a3d | !hbusreq2 & v84564d;
assign v23fca9c = hmaster2_p & v84561b | !hmaster2_p & !v23fc5cd;
assign v23f9307 = hlock3_p & v22fd6fb | !hlock3_p & v230833e;
assign aa26cc = hgrant3_p & v84561b | !hgrant3_p & v22f3bb0;
assign v22eccfc = hmaster2_p & a1fbb6 | !hmaster2_p & v2301a3f;
assign v22fe150 = hbusreq5_p & v23fb10d | !hbusreq5_p & v23f6e64;
assign v23fca40 = hgrant3_p & v23fc618 | !hgrant3_p & v2304fc6;
assign v23f8241 = hbusreq5_p & v23fc920 | !hbusreq5_p & !v23fcd05;
assign v230e7d4 = hbusreq1_p & v22ef403 | !hbusreq1_p & !v23f8490;
assign v22f324c = jx1_p & v85e5cf | !jx1_p & v23f805c;
assign v22ef9f7 = hgrant3_p & v23fc235 | !hgrant3_p & v22f7110;
assign v22f2e82 = hbusreq1_p & v23fc3ee | !hbusreq1_p & v22fdc74;
assign v1506aab = hbusreq6_p & v230e703 | !hbusreq6_p & v2392d0d;
assign v22f8271 = locked_p & v106ae1c | !locked_p & !v106ae19;
assign v9a6a67 = hlock1_p & v23f3ebd | !hlock1_p & v230ea4c;
assign v22f3839 = hgrant3_p & f405c6 | !hgrant3_p & v230b879;
assign v23f5a39 = hmaster2_p & v22f36ff | !hmaster2_p & !v22f3643;
assign v2309280 = hbusreq5_p & v22ec92f | !hbusreq5_p & !v84561b;
assign v23f1824 = hmaster0_p & v22eeb7a | !hmaster0_p & !v23f4edc;
assign v23f9db0 = hgrant3_p & v23fc430 | !hgrant3_p & v2307b9c;
assign v230b713 = hbusreq1_p & fc8e3a | !hbusreq1_p & !v84561b;
assign v230966c = hmaster0_p & v2300d5f | !hmaster0_p & v22f8ee3;
assign v1b87732 = hmaster0_p & v22eb5a9 | !hmaster0_p & v2309057;
assign v2393346 = hgrant1_p & v22f3738 | !hgrant1_p & v230ecac;
assign v2309305 = hmaster0_p & v23fc5d4 | !hmaster0_p & !v23fc28d;
assign v23fc33e = hmaster2_p & v84561b | !hmaster2_p & !v23f34d5;
assign v22ec2cb = hgrant2_p & v2310b8a | !hgrant2_p & v84561b;
assign v22fd029 = hgrant0_p & v84561b | !hgrant0_p & v230fe8e;
assign v22f64e0 = hbusreq0 & v23f65b4 | !hbusreq0 & !v22ee7a7;
assign v2300048 = hmaster2_p & v23fc393 | !hmaster2_p & !v106af73;
assign v23129fa = hgrant4_p & v23fb679 | !hgrant4_p & v23fbf48;
assign v23115f4 = hmaster0_p & v22f5992 | !hmaster0_p & v22ff92c;
assign v23f15c1 = hmaster2_p & v23f79d2 | !hmaster2_p & a1fbcb;
assign v230ba92 = hmaster0_p & v22f5b7c | !hmaster0_p & v22f9f47;
assign v8be441 = hbusreq1_p & v22f1ece | !hbusreq1_p & v230466d;
assign v23f3d14 = hlock0_p & v22ee9be | !hlock0_p & !v845622;
assign v23fc1b3 = hlock3_p & v12cde1b | !hlock3_p & v2305aea;
assign v230cb63 = hbusreq4 & v23fba11 | !hbusreq4 & v23fc223;
assign v22f9e08 = hbusreq4 & v2300de1 | !hbusreq4 & v84561b;
assign v8902b0 = hbusreq5_p & v23fcfbe | !hbusreq5_p & v845620;
assign v23fc92a = hgrant0_p & v23f1b3d | !hgrant0_p & v22ee8d8;
assign v23f47a1 = hmaster0_p & v230f072 | !hmaster0_p & v23fc3c2;
assign v22f7928 = hgrant2_p & v9526ac | !hgrant2_p & v2302149;
assign v2305a12 = hbusreq2_p & v2306d07 | !hbusreq2_p & v84561b;
assign v2312162 = hbusreq6_p & v230d66e | !hbusreq6_p & v84561b;
assign v230c910 = hgrant1_p & v845626 | !hgrant1_p & v2300b4f;
assign b00ad3 = hmastlock_p & v23f8e1f | !hmastlock_p & v84561b;
assign v23f3310 = hlock0_p & v23fbac1 | !hlock0_p & v23f5b39;
assign v23fb813 = hmaster0_p & v2307fcd | !hmaster0_p & v23060bb;
assign v23fc30a = hmaster0_p & v22ee394 | !hmaster0_p & v2303cda;
assign v23fbdf3 = jx0_p & v84561b | !jx0_p & v23117c5;
assign v23f50d9 = hmaster0_p & v22f4db6 | !hmaster0_p & !v22eb3bc;
assign v22fb841 = hgrant2_p & v84561b | !hgrant2_p & !v23001e2;
assign b6c104 = hgrant1_p & v84561b | !hgrant1_p & v22ed03d;
assign v23fcbc8 = hgrant5_p & v84561b | !hgrant5_p & v2308f80;
assign v23f6f4d = hlock5_p & v22f0105 | !hlock5_p & v191b096;
assign v2309d97 = hmaster2_p & v23fc98e | !hmaster2_p & v23fb966;
assign v230bafe = hbusreq1 & v22f8d74 | !hbusreq1 & v84561b;
assign v23faa5c = hmaster2_p & v22f15fe | !hmaster2_p & !v23fc530;
assign v23fb913 = hbusreq0_p & v22fa7f5 | !hbusreq0_p & v23fc1de;
assign v2304074 = hbusreq2_p & v9526ac | !hbusreq2_p & v23f972e;
assign v22f92a2 = hbusreq4 & v22f3d4b | !hbusreq4 & v2312f81;
assign v23fcc95 = hbusreq3 & v22fe573 | !hbusreq3 & v23fcc08;
assign bd7b44 = jx1_p & v1aae2e4 | !jx1_p & v23fcaae;
assign v22f0dc9 = hgrant3_p & v22f0aea | !hgrant3_p & v23fc820;
assign v23fcaaa = hburst1 & v22f3294 | !hburst1 & v23fc529;
assign v230e311 = hgrant0_p & v2310a7e | !hgrant0_p & v22eefab;
assign v23f16f6 = hburst0 & v22f3294 | !hburst0 & !v84561b;
assign v23012c6 = hbusreq5_p & v23fa2ec | !hbusreq5_p & v9ab66e;
assign v22f654f = hbusreq6 & v22f0c90 | !hbusreq6 & v84561b;
assign v23fcb9c = hgrant3_p & v22ff21b | !hgrant3_p & v22f7524;
assign v22fa56f = hlock1_p & v84561b | !hlock1_p & !fc8ab7;
assign v2309c99 = hmaster2_p & v23f9414 | !hmaster2_p & v2310d04;
assign v23fcb47 = hgrant5_p & v23f38ff | !hgrant5_p & v2391a89;
assign v22f800e = hmaster1_p & v23f7822 | !hmaster1_p & !v23f49cd;
assign v230f2d1 = hbusreq5 & v2301505 | !hbusreq5 & v84561b;
assign v23fb1a0 = hmaster2_p & v22eefd1 | !hmaster2_p & v23f0169;
assign v230ecac = hbusreq1_p & v230e6ea | !hbusreq1_p & v22ecced;
assign v23fcb7c = hmaster2_p & v23fcf70 | !hmaster2_p & !v84561b;
assign v22f9d79 = hlock6_p & v22f882c | !hlock6_p & v22f0dc0;
assign v23041ee = hmaster2_p & b9d02f | !hmaster2_p & v23fc7ee;
assign e1e34d = hmaster1_p & v239315b | !hmaster1_p & v23fba19;
assign v106af1c = hbusreq4 & v23f790a | !hbusreq4 & v230eaa1;
assign v23f67e2 = hbusreq3_p & v22fc99c | !hbusreq3_p & v23089c5;
assign v2301105 = hgrant3_p & v84561b | !hgrant3_p & !v230fd1c;
assign v22f1383 = hbusreq4_p & v2301292 | !hbusreq4_p & v23f515d;
assign v23fb4ba = hbusreq3_p & v23044cf | !hbusreq3_p & v23fc88c;
assign v23f6f5c = hbusreq0_p & v22fb09f | !hbusreq0_p & !v22fcf55;
assign v2303539 = hgrant1_p & v84561b | !hgrant1_p & !v23fb107;
assign v22f2564 = hgrant3_p & v84561b | !hgrant3_p & v22f8d0c;
assign v23f1109 = hgrant3_p & v2305a69 | !hgrant3_p & v23060ed;
assign v23f447e = hbusreq3_p & v22fb4ab | !hbusreq3_p & v23050c1;
assign v2305339 = jx2_p & v22f6534 | !jx2_p & v22fbbcc;
assign v22f8c55 = jx1_p & v22fa1ab | !jx1_p & a2cc4e;
assign v23f6d80 = hgrant1_p & v22f3d5a | !hgrant1_p & v22facd1;
assign v2304883 = stateG10_5_p & v22eb5cc | !stateG10_5_p & v23fc3cb;
assign v23001e2 = hbusreq2_p & v2305fe0 | !hbusreq2_p & v84564d;
assign v2392eb5 = hmaster1_p & v23fbf13 | !hmaster1_p & v106af28;
assign v23fbdf8 = jx2_p & v2301567 | !jx2_p & v2312e30;
assign v23fba18 = hmaster2_p & v845620 | !hmaster2_p & v23fc7ee;
assign v23fd00e = hbusreq4_p & bf150c | !hbusreq4_p & v22ec150;
assign v23fcd8d = hmaster2_p & v23fc0c9 | !hmaster2_p & v13afb18;
assign v230de18 = hbusreq5_p & v22eb332 | !hbusreq5_p & v84561b;
assign v23fbd04 = hbusreq4 & v230e54d | !hbusreq4 & v22fdfdd;
assign v22f3ed0 = hbusreq5_p & a1fbc2 | !hbusreq5_p & v22eb377;
assign v22ee6cb = hlock3_p & v87d84c | !hlock3_p & v22ec616;
assign v23f581f = hbusreq3_p & v23f1ccc | !hbusreq3_p & v23f4bfc;
assign a1fdf8 = hmaster0_p & v23fbf85 | !hmaster0_p & !v96c563;
assign v12cddb2 = hbusreq5 & v23f3d14 | !hbusreq5 & v84561b;
assign stateG10_2 = !v21ea5eb;
assign v23f7218 = hbusreq2_p & v23fc91f | !hbusreq2_p & v22ee59c;
assign v22f8312 = hbusreq4 & v22f28c4 | !hbusreq4 & v84561b;
assign v230e831 = hgrant3_p & v84561b | !hgrant3_p & v23f75e5;
assign v23f850a = hgrant5_p & v23111ee | !hgrant5_p & v22ecb9d;
assign v2300338 = hbusreq0_p & v106af4d | !hbusreq0_p & v23f2553;
assign v22fef36 = hgrant2_p & v22f8271 | !hgrant2_p & !v106ae19;
assign da38bd = hbusreq5 & v23fbf9d | !hbusreq5 & !v2309c70;
assign v23fcf69 = hgrant1_p & v23fb67c | !hgrant1_p & v230e897;
assign v22fbbcc = hgrant4_p & bd6575 | !hgrant4_p & v22f6db5;
assign v22fd7ee = hbusreq4 & v22eefd1 | !hbusreq4 & v84561b;
assign v23fbfb1 = hmaster1_p & v22fda35 | !hmaster1_p & v23117cd;
assign v23fc539 = hbusreq5_p & v23f3115 | !hbusreq5_p & v23faf60;
assign v22fb1f3 = hmaster2_p & c24eac | !hmaster2_p & bd9ab5;
assign v1aad5ad = hbusreq2_p & v22f88aa | !hbusreq2_p & v84561b;
assign v22faa40 = hgrant1_p & v22ee956 | !hgrant1_p & v22f4727;
assign v23fc8bc = hbusreq6_p & v23fbfd8 | !hbusreq6_p & v230764f;
assign v23f23e8 = stateG10_5_p & v22f9de9 | !stateG10_5_p & !v230baba;
assign v23fca6f = hbusreq4_p & v2303314 | !hbusreq4_p & v84561b;
assign v2301d76 = stateG2_p & v84561b | !stateG2_p & v23f4c9c;
assign v23063f8 = hgrant5_p & v22f05f3 | !hgrant5_p & v230b089;
assign v23135f8 = hmaster2_p & v23fca2a | !hmaster2_p & v84561b;
assign v2304d08 = hmaster0_p & v2303acd | !hmaster0_p & v23fc67b;
assign v22f197e = stateA1_p & v84561b | !stateA1_p & !v230177d;
assign v2302e80 = hbusreq0 & v22ff315 | !hbusreq0 & v845629;
assign v22fa371 = hgrant3_p & v22f6219 | !hgrant3_p & v23f7db2;
assign v22f61cc = hgrant0_p & v23fcbd3 | !hgrant0_p & v23045e7;
assign v23fb121 = hlock0_p & v22f3502 | !hlock0_p & v23fad76;
assign v22faa0e = hlock1_p & da38c1 | !hlock1_p & v84561b;
assign v23fc493 = hmaster2_p & v23f54ef | !hmaster2_p & v22fc8e5;
assign v22edf7b = hbusreq6_p & v22f7832 | !hbusreq6_p & !v84561b;
assign v1aad847 = hbusreq2_p & v23f6dc8 | !hbusreq2_p & !v84561b;
assign v2308be0 = hmaster1_p & v2307edb | !hmaster1_p & !v84561b;
assign v230f693 = hbusreq3_p & v1aad609 | !hbusreq3_p & v84561b;
assign v230f2d6 = hbusreq0 & v22f4e0b | !hbusreq0 & v230f5a3;
assign v23f9e84 = hmaster0_p & v2308967 | !hmaster0_p & !v2301c2e;
assign v22ffb12 = hgrant1_p & v845626 | !hgrant1_p & v22f14ed;
assign v23fc29c = hbusreq2_p & v23fc21d | !hbusreq2_p & v84564d;
assign v23fbe36 = jx0_p & v23fcabd | !jx0_p & v22ef3f8;
assign v2305847 = hbusreq6_p & v12cda8f | !hbusreq6_p & v2305498;
assign v23fcc67 = hbusreq3 & v230f370 | !hbusreq3 & v22f35f5;
assign v22f8b41 = hlock3_p & v23f2fd2 | !hlock3_p & v239288d;
assign a83396 = hbusreq3 & v22f4e64 | !hbusreq3 & v84561b;
assign v230ae19 = hgrant0_p & v84561b | !hgrant0_p & v23139aa;
assign v2305e79 = hmaster2_p & v22fc19c | !hmaster2_p & v22f03cf;
assign v2305148 = hgrant1_p & v12cd9f9 | !hgrant1_p & v22ec4ce;
assign v22f990d = hbusreq4_p & v23fbbeb | !hbusreq4_p & v231242d;
assign v22f18df = hgrant0_p & v84564d | !hgrant0_p & v2392e9d;
assign v231398c = hgrant3_p & v22ffa6e | !hgrant3_p & v23fc30d;
assign v868c84 = hmaster2_p & v22fc8e5 | !hmaster2_p & v2391950;
assign v22f067f = hbusreq5_p & v23f646e | !hbusreq5_p & v2307a0f;
assign v23f512e = hgrant2_p & v106af73 | !hgrant2_p & v191a879;
assign v22fecb6 = hbusreq3_p & v22ed83b | !hbusreq3_p & v23fcfcf;
assign v2301997 = hbusreq1 & bd74c0 | !hbusreq1 & v23fa2ec;
assign v23f51a4 = hgrant5_p & v84561b | !hgrant5_p & v23fc8eb;
assign v23fc8d7 = hburst1_p & v84561b | !hburst1_p & !v845649;
assign v862ce7 = hmaster1_p & v845631 | !hmaster1_p & v23f6a42;
assign v22ff1dd = hbusreq1_p & v2301509 | !hbusreq1_p & v84561b;
assign v2311a24 = jx2_p & v23f2a15 | !jx2_p & v22fcc70;
assign bd9916 = hready & v2302136 | !hready & v84564d;
assign v23fcbb6 = hbusreq1_p & v23f6ec1 | !hbusreq1_p & v2304bc1;
assign v22ff5ea = hmaster2_p & v84561b | !hmaster2_p & v23f4572;
assign v22ec2d6 = jx1_p & v231242a | !jx1_p & v230e991;
assign v230a56a = hmaster2_p & v230a035 | !hmaster2_p & !v84561b;
assign v22f915d = stateG10_5_p & v22ef683 | !stateG10_5_p & v845620;
assign v23f741d = hbusreq4_p & v23f3f38 | !hbusreq4_p & !v106a7a1;
assign v23f5f5f = hbusreq1_p & v22ffc07 | !hbusreq1_p & !v84561b;
assign v23fb08d = hmaster0_p & v23fb926 | !hmaster0_p & v22ec77a;
assign v22f75d4 = hbusreq1 & v23060d4 | !hbusreq1 & v23f87f4;
assign v23fb788 = hlock1_p & v230c116 | !hlock1_p & v191ae6e;
assign v22f1e46 = hbusreq3 & v22f5355 | !hbusreq3 & v84561b;
assign v23fa345 = hbusreq5_p & v2310475 | !hbusreq5_p & v84561b;
assign v23fbc75 = hburst0 & v23fc8a3 | !hburst0 & !v84561b;
assign v23f6ba0 = locked_p & v22ed56a | !locked_p & v84561b;
assign v23f8a99 = hgrant5_p & v23007a1 | !hgrant5_p & v22f3c3d;
assign v22f442c = hgrant0_p & v845622 | !hgrant0_p & v2302d85;
assign v2312057 = hlock1_p & v84561b | !hlock1_p & !v22ff6f9;
assign da38c9 = hgrant3_p & v22fe392 | !hgrant3_p & v23fbe1d;
assign v23102b2 = hgrant6_p & v84561b | !hgrant6_p & v22fd02d;
assign v22ff5c1 = jx0_p & v23f17ff | !jx0_p & v23f5a6d;
assign v23f3c84 = hmaster0_p & bd8ccb | !hmaster0_p & e1df54;
assign v2312acc = hgrant0_p & v23f5043 | !hgrant0_p & v23fbac1;
assign v22f0326 = hbusreq2_p & v2391c58 | !hbusreq2_p & v22ee59c;
assign v22ec09c = hbusreq1_p & v23fc355 | !hbusreq1_p & !v230345c;
assign v22ed5be = hmaster2_p & v23fa463 | !hmaster2_p & v84561b;
assign v23fbaa2 = hbusreq4 & v230aa94 | !hbusreq4 & v22eba71;
assign b61053 = hbusreq4_p & v2303a58 | !hbusreq4_p & v2305a91;
assign v22fe300 = hbusreq1 & v22f0add | !hbusreq1 & v84561b;
assign v23fcf25 = hbusreq2_p & v84561b | !hbusreq2_p & v22efdb1;
assign v22efae1 = hbusreq5 & v23f65b4 | !hbusreq5 & v84561b;
assign v1aad586 = hgrant0_p & v22f215c | !hgrant0_p & !v23fc7fb;
assign v230113d = hmaster2_p & v2309b7e | !hmaster2_p & !a39dae;
assign v23fc804 = hmaster2_p & v23fcb65 | !hmaster2_p & !v2391d17;
assign v23fc34f = hbusreq4 & v22fdcc7 | !hbusreq4 & v84561b;
assign v230524c = jx2_p & v23fd016 | !jx2_p & v22f509a;
assign v22ed495 = hgrant5_p & v23f494b | !hgrant5_p & v23fc8df;
assign v23fbb7e = hbusreq1_p & v22f1d8b | !hbusreq1_p & !v84561b;
assign v22f19dd = hmaster1_p & v23fbf8d | !hmaster1_p & v22fb8c0;
assign b52881 = hmaster0_p & v230eb9e | !hmaster0_p & v2310ab0;
assign v2312cb7 = hbusreq3 & v22f779f | !hbusreq3 & v23f9fb5;
assign v2303270 = hmaster2_p & v84561b | !hmaster2_p & v23f6729;
assign v22fdbbe = hbusreq3 & v2392258 | !hbusreq3 & !v2300479;
assign v23f052e = hgrant1_p & v84564d | !hgrant1_p & !v84561b;
assign v230c52a = hgrant5_p & b5e222 | !hgrant5_p & v23f40ba;
assign v22fd171 = hmaster2_p & v84561b | !hmaster2_p & v230cf0c;
assign v22fa195 = hbusreq2_p & v15072de | !hbusreq2_p & !v84561b;
assign v22eaa94 = hbusreq5_p & a1382d | !hbusreq5_p & v230bb30;
assign v23fb90f = hmaster2_p & v23fc716 | !hmaster2_p & v23fca72;
assign v23fc200 = stateG2_p & v84561b | !stateG2_p & v12cda44;
assign v22ee4ab = hmaster2_p & v2309c8a | !hmaster2_p & b9d013;
assign v9df685 = hmaster0_p & v22f7273 | !hmaster0_p & v2309440;
assign v2307836 = hbusreq0 & v22f0073 | !hbusreq0 & v15074fb;
assign v2313595 = hgrant3_p & v23fbd33 | !hgrant3_p & v230979d;
assign v2300f82 = hmaster2_p & v106ae19 | !hmaster2_p & !v22f3a35;
assign v22fb6f9 = hmaster2_p & v23fc925 | !hmaster2_p & v23fba9a;
assign v22ef1eb = hgrant3_p & v23fcb2d | !hgrant3_p & v2312925;
assign v2302370 = hmaster2_p & v23f32eb | !hmaster2_p & v84561b;
assign v88bc32 = hlock0_p & v22f9ef0 | !hlock0_p & v23934e0;
assign v23fcca4 = hbusreq0_p & v230af3a | !hbusreq0_p & v230b02b;
assign v22fb71d = hgrant0_p & v22ec303 | !hgrant0_p & !v84561b;
assign v22f42c9 = stateG10_5_p & v191b1f3 | !stateG10_5_p & !v22eb1f5;
assign v23f56c0 = hbusreq3_p & v23fb18e | !hbusreq3_p & v22f61d2;
assign v23f98f8 = hlock5_p & v84561b | !hlock5_p & !v23f820a;
assign v230b78b = hbusreq2 & v22f0d8d | !hbusreq2 & v84561b;
assign v13aff3b = hbusreq0 & v230e032 | !hbusreq0 & !v84561b;
assign v22ed984 = hgrant0_p & v84561b | !hgrant0_p & v230b161;
assign v22fc122 = hbusreq0 & v22f446e | !hbusreq0 & !v84561b;
assign v22f6af6 = hbusreq4_p & v22ede51 | !hbusreq4_p & v22fe1c8;
assign v23fcddb = hbusreq1_p & v230d2c7 | !hbusreq1_p & v23fb9a0;
assign v23fc1a7 = hbusreq2_p & a1fc4e | !hbusreq2_p & !v22edaf2;
assign v2393f17 = hbusreq5 & v230da4a | !hbusreq5 & !v23fc839;
assign v12cd4c5 = hmaster2_p & v23f45d2 | !hmaster2_p & v22fec8c;
assign v22fb759 = hbusreq3_p & v230b740 | !hbusreq3_p & v23fc114;
assign v22edcf4 = hmaster2_p & v22ffb12 | !hmaster2_p & v22fe346;
assign v22eafde = hmaster2_p & v191a86f | !hmaster2_p & v22eaaba;
assign v22f1153 = hmaster2_p & v84561b | !hmaster2_p & v23fa2b5;
assign v23087e9 = hmaster2_p & v22f9321 | !hmaster2_p & v23f6e68;
assign v2367a5a = hmaster0_p & e1d75b | !hmaster0_p & v23098d3;
assign v230f82f = jx2_p & fc8fcf | !jx2_p & v230387b;
assign v230545b = hmaster2_p & v23f14bc | !hmaster2_p & v23112ad;
assign v230bbb3 = hbusreq1_p & v23fc13a | !hbusreq1_p & !v84561b;
assign v2305f5e = hbusreq5_p & f40761 | !hbusreq5_p & v2303ce2;
assign v22f064a = hbusreq3_p & v85c335 | !hbusreq3_p & v22ee657;
assign v2308bcd = hgrant5_p & v22fd6d8 | !hgrant5_p & v22f71ca;
assign v23fd057 = hgrant5_p & f40c9d | !hgrant5_p & v2305522;
assign v23f0f9a = hgrant6_p & v230aec3 | !hgrant6_p & v231269d;
assign v2307d0e = hmaster2_p & v230b62c | !hmaster2_p & v22f0b62;
assign v2346b41 = hbusreq3_p & v22eed1b | !hbusreq3_p & v230a905;
assign v22ed4b0 = hbusreq4_p & v22f2e0c | !hbusreq4_p & v84561b;
assign v22ee47d = hmaster2_p & v23f4426 | !hmaster2_p & v23fc127;
assign v23f623e = jx3_p & v84561b | !jx3_p & !v8eb4b5;
assign v230f70d = hbusreq1 & v13afe3a | !hbusreq1 & !v22f9a51;
assign v230d32d = hbusreq0 & v2312ea7 | !hbusreq0 & v84561b;
assign v23f7d2e = hmaster2_p & v230b621 | !hmaster2_p & v8ef087;
assign v22fa3f5 = hbusreq6_p & v23fc8a2 | !hbusreq6_p & v231156b;
assign v22ffa6e = hlock3_p & v23f651a | !hlock3_p & !v84561b;
assign v23f3d7d = hready_p & v22f86fc | !hready_p & v23017b3;
assign v23f4808 = hgrant1_p & v84561b | !hgrant1_p & v22f3d00;
assign a1fcb8 = hgrant3_p & v23fc7a7 | !hgrant3_p & v12cd4be;
assign v230c872 = hbusreq3_p & v23fcb17 | !hbusreq3_p & v22f5437;
assign v22fb890 = hbusreq5 & v84564d | !hbusreq5 & v23fbb35;
assign v230889a = hmaster0_p & v23fae84 | !hmaster0_p & !v230a24c;
assign v23fcc49 = hmaster2_p & v22fe421 | !hmaster2_p & v84561b;
assign v22f419a = hbusreq1_p & v2308ae7 | !hbusreq1_p & bab0c9;
assign v23fc74c = hbusreq5_p & v22f5e18 | !hbusreq5_p & v84561b;
assign v230017e = hgrant3_p & b95000 | !hgrant3_p & v22f7d9a;
assign v2302868 = hbusreq0_p & v84562b | !hbusreq0_p & v23fbab2;
assign v22f8026 = hbusreq0 & v23f5043 | !hbusreq0 & v84561b;
assign v22ee956 = hbusreq2_p & a1fbc2 | !hbusreq2_p & v22eb377;
assign v22fd67c = hmaster0_p & v22feec8 | !hmaster0_p & v2302abd;
assign v22ecff8 = hlock0_p & v84561b | !hlock0_p & v23fbf08;
assign v845671 = stateG10_5_p & v84561b | !stateG10_5_p & !v84561b;
assign v23065d3 = hmaster0_p & v23fca4e | !hmaster0_p & v22f8cb9;
assign v22ee0ea = hmaster0_p & v23fcea2 | !hmaster0_p & v22ef5cd;
assign v23095fa = hlock2_p & fc8e3a | !hlock2_p & v84561b;
assign v22eec21 = hmaster2_p & v84561b | !hmaster2_p & v23fc4f5;
assign v23fca67 = hbusreq4_p & v23f6fe8 | !hbusreq4_p & v23021ec;
assign v23fb6ce = hbusreq5_p & v22ef983 | !hbusreq5_p & !v230262f;
assign v23fcfd6 = hbusreq5_p & v22fd8a6 | !hbusreq5_p & v23fc570;
assign v22f13ad = hbusreq5_p & v23f646e | !hbusreq5_p & v23fb55a;
assign v23fbefa = hbusreq0 & v2312f7e | !hbusreq0 & !v23022b1;
assign v8eb4b5 = jx1_p & v84561b | !jx1_p & !v84561b;
assign v230f453 = hbusreq5_p & v22ee956 | !hbusreq5_p & v23fc253;
assign v23045c3 = hgrant3_p & v23fb0c0 | !hgrant3_p & v23101b0;
assign ac37a1 = hready & v22f1ca0 | !hready & !v84561b;
assign v22f4d37 = hmaster2_p & v84562a | !hmaster2_p & v23f60ef;
assign v23fb537 = hmaster0_p & v2307816 | !hmaster0_p & v22ffffd;
assign v2302353 = hmaster2_p & v23101b1 | !hmaster2_p & v2311a3e;
assign v22eced4 = hburst1 & v22fdb21 | !hburst1 & af3c3f;
assign b0df38 = hbusreq1_p & v23fca36 | !hbusreq1_p & v22f7241;
assign v23f74b7 = hmaster0_p & v2304a06 | !hmaster0_p & v22eec2a;
assign v8a894a = hbusreq3 & v22f1762 | !hbusreq3 & v84561b;
assign v191ad69 = hbusreq5_p & v22ee0c4 | !hbusreq5_p & v2300290;
assign v23fcc22 = hbusreq5_p & v23fc153 | !hbusreq5_p & v23005e2;
assign v23fbabc = hmaster1_p & v230887b | !hmaster1_p & !v22f3f9f;
assign v230e979 = hbusreq3_p & v22f2c87 | !hbusreq3_p & v22eb74d;
assign v2311b20 = hgrant3_p & b00ac7 | !hgrant3_p & v230be96;
assign be86f6 = hmaster0_p & v23fcb8a | !hmaster0_p & v23fc9b7;
assign bd0733 = hbusreq6_p & v23f5e3d | !hbusreq6_p & v22ee681;
assign v23f1c0b = hbusreq6_p & e1e75d | !hbusreq6_p & !v84561b;
assign v23075a5 = hmaster2_p & v1506ad8 | !hmaster2_p & v230d814;
assign v22fa205 = hburst1_p & v22f53f3 | !hburst1_p & !v22f178d;
assign v22fed4f = hmaster0_p & v2300d0f | !hmaster0_p & v230b4b4;
assign v23fbe7b = hmaster0_p & v23fd051 | !hmaster0_p & v230e9d1;
assign v22fcdd3 = hbusreq3_p & v230c4c3 | !hbusreq3_p & v23fb143;
assign v2301c48 = hmaster0_p & v23fc34f | !hmaster0_p & v230c653;
assign v230e72d = hbusreq5 & v2306b2e | !hbusreq5 & !v845622;
assign v22f5734 = hbusreq1 & v230f5ee | !hbusreq1 & !v23067c1;
assign v23916d8 = jx1_p & v23f5686 | !jx1_p & v2301c10;
assign v22f5136 = hbusreq3_p & v23fb77d | !hbusreq3_p & v230a05f;
assign v230e800 = hbusreq4_p & a05106 | !hbusreq4_p & v230d532;
assign v2300479 = hmaster2_p & v84561b | !hmaster2_p & v22ee7a7;
assign v12cd63d = hmaster0_p & v23fb20f | !hmaster0_p & v22f6aa3;
assign v22ffaff = hbusreq5 & v23fb10d | !hbusreq5 & !v84561b;
assign v22f2123 = hmaster2_p & v84561b | !hmaster2_p & v22fbf74;
assign v1e84057 = hbusreq4 & v2307ec5 | !hbusreq4 & v2312be1;
assign v23f0958 = hmaster1_p & v230daec | !hmaster1_p & v84561b;
assign v22eb47c = hmaster1_p & v22fdd29 | !hmaster1_p & !v2311e9f;
assign v23fb115 = hmaster2_p & v22f5037 | !hmaster2_p & v23fb966;
assign v2310a5e = hlock0_p & e1df2d | !hlock0_p & v84561b;
assign v924a36 = hbusreq4_p & ad6e26 | !hbusreq4_p & v2301a99;
assign v22ff9c3 = hbusreq3_p & v23fcb3c | !hbusreq3_p & v23fcff6;
assign v11853d9 = decide_p & v230363f | !decide_p & v23fbe11;
assign v23fbf14 = hbusreq6_p & v23133b7 | !hbusreq6_p & !v84561b;
assign v230840f = hbusreq1 & v23fcf96 | !hbusreq1 & v84561b;
assign v2301da2 = hmaster0_p & b00aa6 | !hmaster0_p & v23070de;
assign v23f416b = hbusreq6_p & v22f16d8 | !hbusreq6_p & v23023aa;
assign v23f710c = jx1_p & v22fbb46 | !jx1_p & v23f55a4;
assign v22fd29a = stateG2_p & v23f6bf3 | !stateG2_p & !v22f349a;
assign v23fc192 = hbusreq3_p & v2300829 | !hbusreq3_p & v23f15ac;
assign v23fce57 = hgrant1_p & v1aae19c | !hgrant1_p & v9e8d9f;
assign v22f0f15 = hlock2_p & v84561b | !hlock2_p & !fc8e3a;
assign v22edd4c = hgrant4_p & v2393bcf | !hgrant4_p & v22ecab2;
assign v230e794 = hbusreq4_p & v22fe820 | !hbusreq4_p & v230e1bd;
assign v22ef062 = hbusreq1_p & v8a3511 | !hbusreq1_p & v84561b;
assign v22fa202 = hmaster0_p & v84561b | !hmaster0_p & !v845645;
assign b9d041 = hbusreq6 & v230c849 | !hbusreq6 & v84561b;
assign v22f1754 = hbusreq3 & v22edb60 | !hbusreq3 & v84561b;
assign v2305c54 = hbusreq3_p & v23fba12 | !hbusreq3_p & v22ed6e1;
assign v845645 = hmaster2_p & v84561b | !hmaster2_p & !v84561b;
assign v22f85a0 = hgrant1_p & v23fb6ff | !hgrant1_p & v22f3000;
assign v2309726 = hbusreq4 & v230c65f | !hbusreq4 & v2301e1a;
assign v23f2eb5 = hbusreq2_p & v22f46ab | !hbusreq2_p & v22ee59c;
assign v2308455 = hbusreq0 & v23128a1 | !hbusreq0 & v84561b;
assign v2306967 = jx1_p & v2306473 | !jx1_p & v2306f4e;
assign v22ec92b = hmaster0_p & v23130da | !hmaster0_p & v22ec350;
assign v23f535c = hmaster2_p & v23fcbcd | !hmaster2_p & v84561b;
assign v230dcd9 = hbusreq4_p & v2312d9c | !hbusreq4_p & v230aa5d;
assign v23fc0f0 = stateG10_5_p & v22f532c | !stateG10_5_p & !a1fba6;
assign v898be2 = hbusreq3_p & v1507157 | !hbusreq3_p & v230e2d4;
assign v22f03aa = hmastlock_p & v230cb9d | !hmastlock_p & !v84561b;
assign v230eb9e = hbusreq6 & v22fce0a | !hbusreq6 & v84561b;
assign v23f1812 = hmaster2_p & v22ee9be | !hmaster2_p & v84561b;
assign v23000a6 = hmaster2_p & v23915e9 | !hmaster2_p & v23126f2;
assign v2305b24 = hbusreq4_p & v23fc26a | !hbusreq4_p & v1aae277;
assign v23f446c = hgrant3_p & v84561b | !hgrant3_p & v22fec92;
assign v230607d = hmaster2_p & v23f5af5 | !hmaster2_p & v22f1b4e;
assign v230ae46 = hmaster0_p & v230d5a9 | !hmaster0_p & v22f0de0;
assign v23f9bcf = hmaster2_p & v22fca75 | !hmaster2_p & v22ed2e5;
assign v22f0362 = hburst1 & v22f80ca | !hburst1 & v191a90b;
assign v22fd48a = hmaster0_p & v23119a8 | !hmaster0_p & v84561b;
assign v23fa36c = hmaster0_p & v2304578 | !hmaster0_p & bd8af4;
assign v2307b64 = hmaster0_p & v239310f | !hmaster0_p & v23f2650;
assign v22f98fd = hbusreq2_p & v22fb7a5 | !hbusreq2_p & v845620;
assign v23fc82c = hgrant1_p & v22fe144 | !hgrant1_p & v23f6a76;
assign v23fb94d = stateG10_5_p & v22fe097 | !stateG10_5_p & !v2303e13;
assign v22fcbcd = hlock0_p & v2306d29 | !hlock0_p & !v191a86f;
assign v23fb5ba = hmaster2_p & v23fbaaa | !hmaster2_p & v23fb999;
assign v22f0a39 = hbusreq4_p & v2301c2a | !hbusreq4_p & v23fbf02;
assign v2300271 = hgrant1_p & v23f57a2 | !hgrant1_p & v22eef57;
assign v23049af = jx1_p & v1aae0dc | !jx1_p & v23f6954;
assign v230a035 = hgrant1_p & v23f6045 | !hgrant1_p & v8e4c22;
assign v22f5242 = hbusreq1_p & v2312057 | !hbusreq1_p & v23fb1aa;
assign v22f4cb3 = hmaster1_p & v22f3c10 | !hmaster1_p & v84561b;
assign v23f5e22 = hmaster2_p & v23f8465 | !hmaster2_p & v84561b;
assign v22fd002 = hgrant3_p & v2310ec8 | !hgrant3_p & e1e726;
assign v22ec8d1 = hmaster2_p & v23fbaaa | !hmaster2_p & v22faa40;
assign v2304b05 = hmaster2_p & v2310754 | !hmaster2_p & v230b0f5;
assign v23f6c16 = hbusreq6_p & v23fb704 | !hbusreq6_p & v23fc941;
assign v22eaff1 = hbusreq5_p & v84561b | !hbusreq5_p & !v22f0d4b;
assign v23061d7 = hbusreq1_p & v22fd72d | !hbusreq1_p & v84561b;
assign v230ccd6 = hmaster0_p & v84561b | !hmaster0_p & v23fc98c;
assign v22f6410 = hbusreq5_p & v22f0ddd | !hbusreq5_p & v22ec6e7;
assign b094ff = hlock0_p & v22fbea4 | !hlock0_p & !v84561b;
assign v1b87776 = hbusreq4_p & v2309b63 | !hbusreq4_p & v23fcc44;
assign v23f0bd2 = hlock1_p & v2312aec | !hlock1_p & v2304bc1;
assign v22ef05d = hbusreq0_p & v2306d29 | !hbusreq0_p & v23126ae;
assign v23fb175 = hgrant1_p & v230320e | !hgrant1_p & v23f2c8b;
assign v230ef09 = hgrant3_p & v84561b | !hgrant3_p & v23029ed;
assign v230fdf7 = hmaster0_p & v23078cb | !hmaster0_p & v23f3d0e;
assign v2306bd7 = hbusreq6_p & v22f8013 | !hbusreq6_p & v84561b;
assign v23fbab0 = hgrant1_p & v2301e25 | !hgrant1_p & v2312cdf;
assign v23fbace = hbusreq4_p & v23fc11b | !hbusreq4_p & v23065d3;
assign v230df5c = hgrant3_p & v23fc4c3 | !hgrant3_p & v23fbce0;
assign v230cd57 = hmaster2_p & a3cb61 | !hmaster2_p & v23f8f25;
assign v22eee6a = hbusreq3_p & v23fc54f | !hbusreq3_p & v23fca07;
assign v191b160 = hmaster0_p & b00aa6 | !hmaster0_p & v23f1160;
assign v231347a = hlock3_p & v23fc14b | !hlock3_p & v23111b2;
assign v23f10a4 = hbusreq1 & v22f03cf | !hbusreq1 & !v845622;
assign v2312d9c = hlock4_p & v22ed1b0 | !hlock4_p & v230aa5d;
assign v23fc2a5 = hbusreq5_p & v22f41ee | !hbusreq5_p & v23fcccd;
assign v1aad98e = hgrant5_p & v2392842 | !hgrant5_p & v22f5b27;
assign v231206c = stateG10_5_p & v23f4fa1 | !stateG10_5_p & v2393c3a;
assign v22f2965 = hbusreq6_p & v22f09b1 | !hbusreq6_p & !v84561b;
assign v2309a71 = hbusreq1_p & v23f9546 | !hbusreq1_p & v23f5b7b;
assign v22ec0d4 = stateG10_5_p & v23fbe4c | !stateG10_5_p & !v191a86f;
assign v22f3dc7 = hmaster2_p & v22fd74b | !hmaster2_p & v84561b;
assign v22fda32 = hlock0_p & v22f2db0 | !hlock0_p & v230f2dc;
assign v2300d6c = hbusreq2 & v869055 | !hbusreq2 & v84561b;
assign v23efb5a = hmaster2_p & v22fe497 | !hmaster2_p & v23fbb4b;
assign v23f83ef = hbusreq1_p & v22f1e96 | !hbusreq1_p & !v22f30fe;
assign v22f9340 = hbusreq6 & v23fc8f6 | !hbusreq6 & v84561b;
assign v22f5e91 = hbusreq1_p & v23fc143 | !hbusreq1_p & v84561b;
assign v22eaf16 = hmaster0_p & v2310895 | !hmaster0_p & v239315b;
assign v22ff789 = hlock4_p & v23f748c | !hlock4_p & v84562b;
assign v239310f = hbusreq6 & v2310d79 | !hbusreq6 & v84561b;
assign v23110a4 = hmaster2_p & v97b973 | !hmaster2_p & v230ea6d;
assign v22eefaf = hbusreq1_p & v23f7700 | !hbusreq1_p & v23f87f4;
assign v23fb107 = hgrant5_p & v22fd379 | !hgrant5_p & !v84561b;
assign v23f437d = hbusreq6_p & v230eed5 | !hbusreq6_p & v84561b;
assign v230557c = hbusreq6 & v23f5ede | !hbusreq6 & v84561b;
assign v22fa662 = stateG10_5_p & v23fb1d4 | !stateG10_5_p & !v23fba6b;
assign v239233a = hgrant3_p & v230cbc4 | !hgrant3_p & v22ee323;
assign a678c9 = hbusreq5 & v230fae0 | !hbusreq5 & v84561b;
assign v23fb540 = stateG10_5_p & v84561b | !stateG10_5_p & !v2313463;
assign v22f811e = hmaster1_p & v22eea0f | !hmaster1_p & !v230128b;
assign v22eec6e = hgrant1_p & v22f3643 | !hgrant1_p & v22fd699;
assign v230dbcc = jx1_p & v230049a | !jx1_p & v84561b;
assign v23fbda1 = hgrant1_p & v22f3d5a | !hgrant1_p & v22fd124;
assign v22fb87a = hmaster0_p & v22ee521 | !hmaster0_p & !v230638a;
assign v22f2e48 = hbusreq4 & v2310d79 | !hbusreq4 & v84561b;
assign v23fc631 = hmaster1_p & v230d849 | !hmaster1_p & v23fc4f4;
assign v230197e = hbusreq3_p & v23f1e3f | !hbusreq3_p & v84561b;
assign v22fc0ee = hbusreq3_p & v23fb4e8 | !hbusreq3_p & v22ecce6;
assign v230153c = hmaster2_p & v23f0699 | !hmaster2_p & !v84561b;
assign v23fc00a = hmaster0_p & v22ef823 | !hmaster0_p & !v23031f0;
assign v22ef9ff = hlock4_p & v2313230 | !hlock4_p & v23fc89d;
assign v230259f = hlock3_p & v23fc335 | !hlock3_p & v2308d20;
assign v953acf = hgrant1_p & v2300fb4 | !hgrant1_p & !v22f78b7;
assign v23fcf54 = hbusreq3_p & v2307aad | !hbusreq3_p & v9180fe;
assign v230a759 = hmaster2_p & v22fcdf6 | !hmaster2_p & v106ae21;
assign v22ebb7b = hgrant1_p & v22ff732 | !hgrant1_p & v23fa9df;
assign v22fd825 = hmaster2_p & v1e84174 | !hmaster2_p & v22fc10a;
assign v22ffea0 = hbusreq2 & v23f65b4 | !hbusreq2 & v84561b;
assign v22edee1 = hgrant0_p & v2309c14 | !hgrant0_p & v23fb4d1;
assign v22ebbf2 = hmaster0_p & v23fb8aa | !hmaster0_p & v23f5893;
assign v230493b = hburst1 & v22fdb21 | !hburst1 & v23f3c20;
assign v230b49b = hmaster2_p & v2310d04 | !hmaster2_p & v22f3618;
assign v1aadf2f = hmaster2_p & v22f8427 | !hmaster2_p & v230058a;
assign v230b27c = hbusreq1_p & v23fcfbe | !hbusreq1_p & v845620;
assign v23065ad = hlock0_p & v23126ae | !hlock0_p & v23094ad;
assign v23f4758 = hbusreq5_p & v22ef983 | !hbusreq5_p & !v22ebedc;
assign v23fbe6d = hlock3_p & v22f7b3e | !hlock3_p & !v84561b;
assign v23090fd = hbusreq6 & v23fc75c | !hbusreq6 & v23043b7;
assign v23f3715 = hbusreq0_p & v22f1a26 | !hbusreq0_p & !v230f8b2;
assign v230aa7a = hgrant3_p & v84562e | !hgrant3_p & v22fab50;
assign v2312231 = hgrant1_p & v22fdc30 | !hgrant1_p & v23fbbbd;
assign v1aad527 = hbusreq4_p & v22f8556 | !hbusreq4_p & v22fb653;
assign v23f95bd = hmaster0_p & v23f6ad0 | !hmaster0_p & !v23fc3da;
assign v2301d10 = hbusreq2_p & v845620 | !hbusreq2_p & v84561b;
assign v23fc630 = hbusreq6 & v23f44bd | !hbusreq6 & v845627;
assign v22f3c6b = hgrant1_p & v23fb5d1 | !hgrant1_p & v22f0332;
assign v2308d20 = hbusreq3 & v23fb8e4 | !hbusreq3 & v845627;
assign v23fc763 = hmaster1_p & v231108b | !hmaster1_p & v1507439;
assign v23fbcfc = hlock0_p & v84561b | !hlock0_p & v23fce98;
assign v22ecb08 = hgrant3_p & v84561b | !hgrant3_p & v23122cb;
assign v23fa903 = hmaster2_p & v845627 | !hmaster2_p & a1fbcb;
assign v23fc370 = hbusreq0_p & v22f8d2b | !hbusreq0_p & v23fcdcf;
assign v23f26fc = hlock3_p & v22f5ab0 | !hlock3_p & v23f53a0;
assign v22eb292 = hgrant0_p & v845647 | !hgrant0_p & !v230e71f;
assign v23fccf0 = hmaster0_p & v22f2aff | !hmaster0_p & !v96c563;
assign v22fc3c7 = hmaster0_p & v23fce64 | !hmaster0_p & v22f2f16;
assign v23fc820 = hmaster2_p & v23fcf7c | !hmaster2_p & v84561b;
assign v23fc5a4 = hbusreq1_p & v23004f1 | !hbusreq1_p & !v23f86f0;
assign v23f59dc = hbusreq4 & v23fc607 | !hbusreq4 & v22f5583;
assign v22f1b23 = hbusreq3 & v23fb4cd | !hbusreq3 & v84561b;
assign v230eb8e = hmaster1_p & v23fbf8d | !hmaster1_p & v23f51cc;
assign v23fcb2a = hmaster0_p & v23fbf6d | !hmaster0_p & v99a622;
assign v2311214 = hmaster2_p & v2309d55 | !hmaster2_p & v22fa700;
assign v22f20b4 = hgrant3_p & v23fb869 | !hgrant3_p & v23fc9a1;
assign v23fca94 = hmastlock_p & v22f4cca | !hmastlock_p & v84561b;
assign v23f9ef5 = hmaster2_p & v23fb1c1 | !hmaster2_p & v2309729;
assign v23f7c65 = hmaster1_p & v84561b | !hmaster1_p & v23010ae;
assign v22feb0d = hbusreq5_p & v23fc920 | !hbusreq5_p & !v23fcd52;
assign v23f6d65 = hmaster2_p & v23fbfb9 | !hmaster2_p & v23fbca3;
assign v23fc755 = hlock0_p & v84561b | !hlock0_p & v845621;
assign v230899e = hmaster0_p & v23026f7 | !hmaster0_p & v84561b;
assign v23fcc50 = hgrant0_p & bd7747 | !hgrant0_p & !v84561b;
assign v22f24ca = hgrant3_p & v2312919 | !hgrant3_p & v22f149c;
assign v22f6671 = hbusreq1_p & v22fc5fd | !hbusreq1_p & v22f316b;
assign v230aa2c = hgrant1_p & v84561b | !hgrant1_p & !v23fc680;
assign v22fe50f = hbusreq0_p & v22f037a | !hbusreq0_p & !v23f32eb;
assign v23fb649 = hgrant2_p & v22fb5b1 | !hgrant2_p & v84564d;
assign v23f5eb6 = hbusreq1_p & v2312f85 | !hbusreq1_p & v84561b;
assign v23fbeec = jx0_p & v23fb14d | !jx0_p & !v23fbb15;
assign v230ef38 = hmaster0_p & v22fc6ca | !hmaster0_p & v22edf29;
assign v230abf6 = hbusreq3_p & v84562b | !hbusreq3_p & v23fc746;
assign v22f9cd9 = hmaster0_p & v22fcdd3 | !hmaster0_p & v1aad4c6;
assign v23120b1 = hbusreq4_p & v23f2380 | !hbusreq4_p & v22f0de4;
assign v23f984b = stateG2_p & v84561b | !stateG2_p & v22ee959;
assign v23f6bf3 = hburst1 & v22ec1cb | !hburst1 & v23f2fe0;
assign v23fc79d = hlock3 & v23064ce | !hlock3 & v22ee1b8;
assign v23f1e1a = hgrant5_p & v23f8d64 | !hgrant5_p & v22eb16b;
assign v22f1ae9 = hlock3_p & v84561b | !hlock3_p & !v22f2eaf;
assign v23fbcce = hmaster2_p & v23fc7d5 | !hmaster2_p & v22f6741;
assign v2300246 = hgrant1_p & v84561b | !hgrant1_p & v22f5421;
assign v2310e10 = hlock1_p & v23f2be7 | !hlock1_p & !v84561b;
assign v23f9465 = hmaster0_p & v2310782 | !hmaster0_p & v191ae7d;
assign v23f11a3 = hlock0_p & v22f56d2 | !hlock0_p & v23fbc17;
assign v230b8ff = hbusreq1_p & v9526ac | !hbusreq1_p & v1506fe9;
assign v22ff469 = hbusreq5_p & v22f45ff | !hbusreq5_p & v84561b;
assign v23fc16b = hmaster2_p & v22fc10a | !hmaster2_p & v22fa105;
assign v230ece0 = hbusreq5_p & v230e4ef | !hbusreq5_p & v23015f8;
assign v1e84195 = hbusreq4_p & v22fd71a | !hbusreq4_p & v230089c;
assign v23fc4a4 = busreq_p & v21b35f9 | !busreq_p & v2300755;
assign v230792c = hmaster2_p & bd951f | !hmaster2_p & v23facc9;
assign b8cd18 = hbusreq5 & v22fb77d | !hbusreq5 & !v23108b7;
assign v22f60ce = hlock4_p & v23f9fc6 | !hlock4_p & v23fb975;
assign v22fbb7f = hbusreq4_p & v2391f9b | !hbusreq4_p & !v84561b;
assign v23f9f9d = hbusreq3 & a8a256 | !hbusreq3 & v84561b;
assign v23fc219 = stateG2_p & v84561b | !stateG2_p & v230a413;
assign v23fbd5c = hbusreq1 & v22f5037 | !hbusreq1 & v22f9927;
assign v230fa1a = hlock0_p & v230448f | !hlock0_p & v22fbe82;
assign v23fbeb3 = hbusreq5_p & v230360b | !hbusreq5_p & v13b0055;
assign v23f44b1 = hbusreq2_p & v2301933 | !hbusreq2_p & v23f5043;
assign v873a56 = hmaster1_p & v23f4fa9 | !hmaster1_p & v22eddfd;
assign v1e84b3d = hmaster0_p & v23fc282 | !hmaster0_p & !c20a75;
assign v230e32f = hmaster2_p & v2312c77 | !hmaster2_p & v22fc7e6;
assign v2301e50 = hbusreq1_p & v22f28d6 | !hbusreq1_p & v22f8c0b;
assign v231262f = hbusreq3_p & v1aadf2f | !hbusreq3_p & v22fbeb3;
assign v22ffc55 = hbusreq5_p & v230cd61 | !hbusreq5_p & v84561b;
assign v22ff36f = hbusreq4_p & v23fb99f | !hbusreq4_p & v23fb821;
assign v23111c0 = hmaster2_p & v84561b | !hmaster2_p & !v22f59e9;
assign v22faa39 = hmaster0_p & v23f9d9a | !hmaster0_p & !v2391a45;
assign v22f03cf = hlock0_p & v23f75aa | !hlock0_p & !v845622;
assign v22f94b6 = hgrant5_p & v23fcb0f | !hgrant5_p & v22f3324;
assign v2309459 = hmaster0_p & v23fbbc3 | !hmaster0_p & v23f97c6;
assign v2301e10 = hmaster2_p & v23f6b11 | !hmaster2_p & v23fba9a;
assign v230f9f1 = hmaster2_p & v230e13a | !hmaster2_p & v22f878c;
assign v22f6618 = hmaster1_p & v23f2c35 | !hmaster1_p & v22ecdc8;
assign v23f54be = start_p & v84561b | !start_p & !v845667;
assign v191ae6e = hgrant5_p & v22f05f3 | !hgrant5_p & v23efe0a;
assign v23f883a = hbusreq1_p & v23f1cd2 | !hbusreq1_p & v22fb5a3;
assign v22f3579 = hgrant3_p & v22f174d | !hgrant3_p & v230dfff;
assign v23fbcef = hbusreq2 & v1aae087 | !hbusreq2 & v84561b;
assign aa8bd6 = hlock0_p & v23fcd5d | !hlock0_p & v845620;
assign v23f7ba2 = hmaster1_p & v23031bc | !hmaster1_p & v23f886a;
assign v230b464 = hmaster0_p & v22f28aa | !hmaster0_p & v22f7713;
assign v22ffdf8 = hgrant3_p & v230b38b | !hgrant3_p & v23fcfdb;
assign v23f1f3f = hgrant4_p & v2302de2 | !hgrant4_p & v23131eb;
assign v23fbf6e = hgrant0_p & v84561b | !hgrant0_p & v1507056;
assign v23f7d57 = hgrant1_p & v22f6e0c | !hgrant1_p & v23fcac8;
assign v2309126 = stateG10_5_p & v12cc72f | !stateG10_5_p & !v2312392;
assign v22ed654 = jx1_p & v22f8acc | !jx1_p & v191acb4;
assign v230a3c9 = hlock6_p & v23f3bd2 | !hlock6_p & v845637;
assign v22fef14 = hmaster1_p & v23f38b1 | !hmaster1_p & v23fc8f3;
assign v22f5215 = hmaster0_p & v2310e4a | !hmaster0_p & !v84561b;
assign v23fc6d6 = hgrant5_p & v23fbeb3 | !hgrant5_p & v2391ada;
assign v23fcb62 = hbusreq6_p & v230c6f1 | !hbusreq6_p & bd772c;
assign v23fc8b3 = hbusreq1 & v2310da0 | !hbusreq1 & v84561b;
assign d49f32 = jx3_p & v873a56 | !jx3_p & v2393ecb;
assign v2300c47 = hbusreq5_p & v23126c6 | !hbusreq5_p & v23fceec;
assign v22f1e96 = hlock1_p & v23f1281 | !hlock1_p & v23f0c9a;
assign v22f2a2f = hmaster2_p & v2301655 | !hmaster2_p & !v84561b;
assign v2313367 = hbusreq3_p & v23fc21c | !hbusreq3_p & v22f2ffe;
assign v22fe51f = hbusreq5_p & v23f4b28 | !hbusreq5_p & v191ab91;
assign v2310253 = hbusreq3_p & v22ef65b | !hbusreq3_p & v84561b;
assign b84615 = hgrant2_p & v84561b | !hgrant2_p & !v230d23a;
assign v23915e9 = hgrant1_p & v845626 | !hgrant1_p & v22fe542;
assign v2302179 = hbusreq3_p & v23fc040 | !hbusreq3_p & v23fba9f;
assign v22f09c5 = hlock3_p & v23f482d | !hlock3_p & v231140b;
assign v2308277 = jx2_p & v23f4a0f | !jx2_p & v99005c;
assign v23101b0 = hmaster2_p & v22f08b7 | !hmaster2_p & v230de50;
assign v1128cd1 = decide_p & v22fd679 | !decide_p & v22ed287;
assign v22f0f7c = hmaster1_p & v2303fa1 | !hmaster1_p & v8f9141;
assign v23fbe82 = hgrant3_p & v84561b | !hgrant3_p & v2301de9;
assign v2392222 = hmaster0_p & v231024c | !hmaster0_p & v23f532f;
assign v22f9532 = jx0_p & v2312628 | !jx0_p & !v2302553;
assign v2308363 = hbusreq4 & v23fc27d | !hbusreq4 & v84561b;
assign v23049f8 = hbusreq3 & v23f60fb | !hbusreq3 & v22fe792;
assign v22fdda4 = hbusreq3_p & v230129b | !hbusreq3_p & v230052f;
assign v22ebfd7 = hbusreq1_p & v2305071 | !hbusreq1_p & !v84561b;
assign v2307edb = hbusreq6_p & v239154a | !hbusreq6_p & v23121aa;
assign v23f3c77 = hmaster2_p & v2308a71 | !hmaster2_p & v23fbaaa;
assign v22fc3b1 = busreq_p & v23036d1 | !busreq_p & v23f4e36;
assign v2306a0e = hmaster1_p & v23fbd1b | !hmaster1_p & v2301d4e;
assign v1aae29a = locked_p & v23fba7e | !locked_p & v13afe8f;
assign v2310c1a = jx1_p & v921155 | !jx1_p & v23f7c65;
assign v2306088 = hbusreq3_p & v2311af8 | !hbusreq3_p & v2312e4e;
assign v22f40e3 = hbusreq1 & v191ae42 | !hbusreq1 & v84561b;
assign v230dd35 = hmaster2_p & v230d9cf | !hmaster2_p & v23f5240;
assign v150742d = busreq_p & a1fbb6 | !busreq_p & v23f7ffb;
assign v12cd3aa = hmaster2_p & v23f6d80 | !hmaster2_p & v230bbce;
assign v23933b0 = hbusreq6_p & v23fcdb8 | !hbusreq6_p & v84561b;
assign v23f62fe = hgrant1_p & v23fb69d | !hgrant1_p & v2391f4b;
assign v23fb736 = jx0_p & v84561b | !jx0_p & v2305aee;
assign v23fcd47 = hmaster0_p & v84564d | !hmaster0_p & v23f2df5;
assign abf6b6 = hbusreq5 & v23f6836 | !hbusreq5 & v84561b;
assign v23074d2 = hbusreq4_p & v2310589 | !hbusreq4_p & v22f878c;
assign v22f18ad = hbusreq0 & v2312f7e | !hbusreq0 & v84561b;
assign v22edccd = jx1_p & v23fad54 | !jx1_p & v2306f4e;
assign v2311918 = hlock0_p & b09503 | !hlock0_p & v84561b;
assign v22fe421 = hbusreq2_p & v23fc91f | !hbusreq2_p & v84561b;
assign v23f0c9a = hbusreq1 & v22ffea0 | !hbusreq1 & !v22f4527;
assign e1dbd6 = hbusreq3 & v22fbf21 | !hbusreq3 & v22ef062;
assign v22f7d33 = hmaster0_p & v22fb465 | !hmaster0_p & v2313595;
assign v22ff3c6 = jx0_p & v22ebe5c | !jx0_p & v22fc68e;
assign v23fc96e = hgrant5_p & v23fbacc | !hgrant5_p & v22efda2;
assign v230fac9 = hmaster2_p & v23fb5d8 | !hmaster2_p & v84561b;
assign v22fa4f7 = hgrant4_p & v845635 | !hgrant4_p & v23fc7d4;
assign v2302ffc = hready_p & v230cf9a | !hready_p & !v23fcdca;
assign v23fc8f8 = hmaster2_p & v22fd0e6 | !hmaster2_p & v22fa105;
assign v22fc58a = hbusreq0_p & v191a86f | !hbusreq0_p & !v13afe8f;
assign v2310ec8 = hmaster2_p & v23fa2ec | !hmaster2_p & v22f4163;
assign v2305811 = hbusreq5_p & v22ed85a | !hbusreq5_p & v23fbdb0;
assign v23fc0b3 = hbusreq3_p & v23fbce4 | !hbusreq3_p & v84561b;
assign v23052a8 = hlock1_p & v23fb709 | !hlock1_p & v22f8fa4;
assign v1aada6e = hbusreq3_p & v2312cb7 | !hbusreq3_p & v84561b;
assign v23f55ea = hbusreq5_p & v191a876 | !hbusreq5_p & v191a879;
assign v12cd3bc = hlock1_p & v22fab6a | !hlock1_p & v22f4168;
assign v230b292 = hmaster2_p & v22f31b2 | !hmaster2_p & v230e916;
assign v230c9f0 = hlock3_p & v22f0719 | !hlock3_p & v22f83f2;
assign v22f1971 = hbusreq4_p & v84561b | !hbusreq4_p & v23fc83e;
assign v22f299f = hgrant0_p & v230b961 | !hgrant0_p & v23f3310;
assign v230bf72 = hgrant3_p & v84561b | !hgrant3_p & !v908162;
assign v2391d8a = jx3_p & v22f5d62 | !jx3_p & v84561b;
assign v22f3e2e = hgrant3_p & v84561b | !hgrant3_p & v23f69cd;
assign v230eef7 = hbusreq2 & v22f3643 | !hbusreq2 & v845620;
assign v23fc5b3 = hmaster0_p & v2308706 | !hmaster0_p & v23fbd8a;
assign v2301bb5 = hbusreq6_p & v1507437 | !hbusreq6_p & v191a909;
assign v23fb6b9 = jx3_p & v23fbf9a | !jx3_p & v23fbd50;
assign v2304a1e = hbusreq5 & v23fc7d5 | !hbusreq5 & v22f0add;
assign v22fdaa5 = hbusreq0 & v22ee7a7 | !hbusreq0 & !v84561b;
assign v12cda57 = hbusreq5_p & v2313618 | !hbusreq5_p & v23022f2;
assign v23fafaf = hgrant3_p & v84562e | !hgrant3_p & v2306e28;
assign v23fbd1a = hbusreq0 & v23fce71 | !hbusreq0 & v84561b;
assign v2309891 = locked_p & v2307460 | !locked_p & v84561b;
assign be4ff1 = hbusreq2_p & v2308a30 | !hbusreq2_p & v23fbc12;
assign v2309a1d = hmaster0_p & v23f6326 | !hmaster0_p & v23fbde1;
assign v23915cb = hbusreq4_p & v22ef44c | !hbusreq4_p & v1e840fd;
assign v22ff6ba = hbusreq4_p & v23fb4a3 | !hbusreq4_p & v22f0869;
assign v22ee68f = hmaster2_p & v23101b1 | !hmaster2_p & v22f7bb9;
assign v230fdc7 = stateG2_p & v2302ca3 | !stateG2_p & b9c92c;
assign e1e6ee = hbusreq4 & v22f5941 | !hbusreq4 & v23f2bc0;
assign v23f39fb = hbusreq3_p & v22fba9a | !hbusreq3_p & v23f4008;
assign v22f1b31 = hbusreq5 & v13affaa | !hbusreq5 & v84561b;
assign v23fb550 = hbusreq3 & v23fbcb1 | !hbusreq3 & !v23f7c8d;
assign v23fb236 = hmaster2_p & v22fbd02 | !hmaster2_p & v22fef20;
assign v22fcf55 = hbusreq0 & v1aae29a | !hbusreq0 & v23f8364;
assign v2393dd2 = hmaster0_p & v1b87752 | !hmaster0_p & v23074cd;
assign v22ebfa3 = hgrant5_p & v23fc788 | !hgrant5_p & !v2308aef;
assign v23fa577 = hgrant3_p & v2382e8c | !hgrant3_p & v23fc0a0;
assign v23f724a = hbusreq4_p & v22f48b7 | !hbusreq4_p & v23f33b2;
assign v23fc51f = hgrant0_p & v23f7961 | !hgrant0_p & !v84561b;
assign v8632f2 = hmaster1_p & v22ee413 | !hmaster1_p & v845629;
assign v22f22ec = hbusreq1_p & v22f0de9 | !hbusreq1_p & !v106ae19;
assign v230965a = hlock3_p & v13afe72 | !hlock3_p & v2309f1a;
assign v23fb1d6 = hmaster2_p & v230de18 | !hmaster2_p & v23fcd14;
assign v23fae22 = hmaster0_p & v22f38ab | !hmaster0_p & !e1e65a;
assign v2303bc3 = hbusreq1_p & v22ef21f | !hbusreq1_p & v84561b;
assign v23fb86a = hmaster0_p & v191aeb3 | !hmaster0_p & v230df5c;
assign v22ee7a7 = locked_p & v2308ae2 | !locked_p & v84561b;
assign v23fb4e1 = hbusreq5 & v22f36ff | !hbusreq5 & !v84561b;
assign v23f9b8d = hgrant1_p & v23035ba | !hgrant1_p & v22f9b5b;
assign v23fbc7f = hmaster0_p & v23101f4 | !hmaster0_p & v23fbd75;
assign v22f3bc9 = stateG10_5_p & v230eb8d | !stateG10_5_p & v845636;
assign v22f3d5a = hbusreq1_p & v22f7859 | !hbusreq1_p & v23fb5b4;
assign v23fb2f5 = hlock1_p & v84561b | !hlock1_p & v22f60c6;
assign v22fba03 = hgrant1_p & v22f0593 | !hgrant1_p & v2305055;
assign v23fc73b = jx1_p & v23f651e | !jx1_p & v23f5500;
assign v2391568 = hgrant3_p & v22f8e29 | !hgrant3_p & v23fbeb2;
assign hgrant6 = f4076d;
assign v22f8543 = hbusreq5_p & v2306414 | !hbusreq5_p & v84561b;
assign a1fda8 = hbusreq3 & v22edb43 | !hbusreq3 & v84561b;
assign v23105b1 = hmaster2_p & v230935d | !hmaster2_p & v9b93b3;
assign v2310969 = hmaster0_p & v23f3f24 | !hmaster0_p & v22eafde;
assign v2303516 = hgrant5_p & v22f13ad | !hgrant5_p & v22fbfe5;
assign v23fc3e1 = hbusreq4 & v23fb933 | !hbusreq4 & v2304899;
assign v22fb49a = hmaster1_p & v23fc438 | !hmaster1_p & v23fca67;
assign v9e3170 = hbusreq0 & v23fd050 | !hbusreq0 & v23124cc;
assign v22f165f = hbusreq6 & v2313144 | !hbusreq6 & v23077dc;
assign v22f5bca = hgrant5_p & v22f05f3 | !hgrant5_p & v230d8c2;
assign v22efb25 = hmaster2_p & v230ed27 | !hmaster2_p & v230dbc9;
assign v22ed7da = hmaster0_p & v23fc6a1 | !hmaster0_p & v22f6ae5;
assign v23fcb6c = hbusreq3 & bd7f18 | !hbusreq3 & !v22fb23d;
assign v22f9f68 = hbusreq4_p & v2305e00 | !hbusreq4_p & v2311e38;
assign v22fbadb = hbusreq2_p & fc8ab7 | !hbusreq2_p & b00ad3;
assign v23fc9f8 = hbusreq5_p & v22fd3f9 | !hbusreq5_p & v84561b;
assign v23fcb14 = hlock0_p & v23f75aa | !hlock0_p & !v84561b;
assign v2304f32 = hbusreq5 & v22f925b | !hbusreq5 & v84561b;
assign v2307b18 = hgrant2_p & v84561b | !hgrant2_p & v22ede4d;
assign v1e841ad = jx2_p & v230d1ff | !jx2_p & v230caee;
assign v23f2504 = hmaster2_p & v23101b1 | !hmaster2_p & v23f01f8;
assign v230fdb8 = hbusreq5_p & v23f08d9 | !hbusreq5_p & v23040f3;
assign v22ff315 = hbusreq2_p & v15070e0 | !hbusreq2_p & !v84561b;
assign v23fcb8a = hbusreq4 & v191b10f | !hbusreq4 & v84561b;
assign v22ef659 = hgrant0_p & v23065ad | !hgrant0_p & v230abf3;
assign v23f44bd = hmaster2_p & v23f79d2 | !hmaster2_p & v22f1faf;
assign v230d1a6 = hgrant0_p & v23f6411 | !hgrant0_p & v2303b9a;
assign v231022d = hbusreq1_p & v23f6ec1 | !hbusreq1_p & v23fc98a;
assign v22ed212 = hgrant3_p & v22f6ae5 | !hgrant3_p & v22ec8d1;
assign v2312d11 = hbusreq2_p & v230219b | !hbusreq2_p & v22f7f74;
assign v9ce77e = hbusreq6 & v22f6aa3 | !hbusreq6 & v23fb20f;
assign v2301e66 = hgrant1_p & v22ec9ce | !hgrant1_p & v23fbe09;
assign v22eefab = hbusreq2_p & v23fc7e5 | !hbusreq2_p & v84561b;
assign v23f6a5b = hmaster0_p & v23fcf87 | !hmaster0_p & v22edd3d;
assign v23f537c = hbusreq5_p & v2303b17 | !hbusreq5_p & v22f9d17;
assign v23fc680 = hgrant5_p & v2303245 | !hgrant5_p & !v84561b;
assign v1aad8ea = hbusreq4 & v230d8b2 | !hbusreq4 & v230c963;
assign v23f5af5 = locked_p & v150742d | !locked_p & !v2309c8a;
assign v22f8c6b = hbusreq6 & v22f3385 | !hbusreq6 & v22ed999;
assign v23fb4a4 = hburst1_p & v2309a51 | !hburst1_p & v84561b;
assign a89109 = hbusreq4_p & v2301937 | !hbusreq4_p & v22fc7e5;
assign v23fb978 = hbusreq2 & v23fc7d5 | !hbusreq2 & v9f4f45;
assign v23f6da6 = jx0_p & v23fca8a | !jx0_p & v84561b;
assign v22f1d80 = hbusreq1_p & v22f0cc4 | !hbusreq1_p & v84561b;
assign v22f1e8e = hmaster1_p & v22f5dc1 | !hmaster1_p & v22f8001;
assign v23fc7ad = hbusreq3_p & v230b0d6 | !hbusreq3_p & v230a735;
assign v23fc85b = hmaster0_p & v23fcdd1 | !hmaster0_p & !v230e9d1;
assign v23fc120 = hgrant1_p & v84561b | !hgrant1_p & v23fcbc8;
assign v191abed = hmaster1_p & v2311d05 | !hmaster1_p & v2305a52;
assign v22fb43e = hmaster0_p & v22feec8 | !hmaster0_p & !v22ffc90;
assign v2309add = hbusreq4_p & v23fbe14 | !hbusreq4_p & v2302d56;
assign v23fc1c8 = hgrant0_p & v22fc517 | !hgrant0_p & v22f302f;
assign v2393332 = hbusreq3_p & v23f8a29 | !hbusreq3_p & v22faf3a;
assign v22f866f = hlock1_p & v2308c50 | !hlock1_p & v23fc8a4;
assign v23f232d = hbusreq6 & v22eaeaf | !hbusreq6 & v84561b;
assign v230b5cc = hlock4_p & v23fc684 | !hlock4_p & v84561b;
assign v23f3cb8 = hbusreq2_p & v230536c | !hbusreq2_p & v84561b;
assign v23101ee = hbusreq2 & v23fc514 | !hbusreq2 & !v22f91c9;
assign v8c495d = hmaster0_p & v22f2abb | !hmaster0_p & v23fbe79;
assign v23063db = hgrant6_p & v84561b | !hgrant6_p & v22fcfee;
assign v2300d5f = hbusreq3_p & b00ac4 | !hbusreq3_p & v23f8a97;
assign v230b7c8 = hbusreq4_p & v22f83d7 | !hbusreq4_p & v23f4ff3;
assign v23f4c9c = hburst0_p & v22f178d | !hburst0_p & !v22fa205;
assign v2300934 = hbusreq5_p & v23fb4e1 | !hbusreq5_p & !v84561b;
assign v23fbb15 = jx3_p & v84561b | !jx3_p & v23f3c86;
assign v2307a21 = hmaster0_p & v23fbf17 | !hmaster0_p & v22f1166;
assign v230bd36 = hmaster2_p & v23fbf8b | !hmaster2_p & !bd7c3f;
assign v23fb51a = hmaster0_p & v23f7ad1 | !hmaster0_p & v23f39f2;
assign v12ce195 = hbusreq2 & v2312f7e | !hbusreq2 & !v22f91c9;
assign v22fe261 = jx1_p & v85e5cf | !jx1_p & !v230538a;
assign v23008e6 = hbusreq3 & v23fbddc | !hbusreq3 & v23f61ba;
assign v230564d = jx3_p & v22f9601 | !jx3_p & v22fab2d;
assign v22eb6e4 = hmaster0_p & v23fc0a3 | !hmaster0_p & v2303b0a;
assign v230f5b9 = hmaster2_p & v23fbaaa | !hmaster2_p & v22ebb7b;
assign v23fc58d = hbusreq3_p & v22fbef0 | !hbusreq3_p & v84561b;
assign v23f2cbb = hbusreq0 & v22f60c6 | !hbusreq0 & v230d7b7;
assign v23fc84e = hgrant1_p & v22fbf74 | !hgrant1_p & v22f9dd0;
assign v22f2ff1 = hmaster0_p & v23fbbbf | !hmaster0_p & v22f1acb;
assign v23f53e9 = hbusreq3_p & v230160e | !hbusreq3_p & v23fbb73;
assign v23fc640 = hlock4_p & v22ff114 | !hlock4_p & !v230a0ad;
assign v23f6cef = hbusreq1_p & v23faa16 | !hbusreq1_p & v2300936;
assign v23fbde0 = hbusreq1_p & v230e4ef | !hbusreq1_p & v22fcbac;
assign v22f0add = hready & v23fcb89 | !hready & v22f197e;
assign v22f9927 = hbusreq2 & v2306220 | !hbusreq2 & !v84561b;
assign v22f3be2 = hmaster2_p & v22fc10a | !hmaster2_p & v23fbab0;
assign v22f670f = hmaster2_p & v2310d04 | !hmaster2_p & v23f940c;
assign v23fbb1b = hmaster1_p & v23fcf15 | !hmaster1_p & !v2307a9e;
assign a1fd9c = hbusreq6 & v22f0d89 | !hbusreq6 & v22f0331;
assign v22eedcf = hbusreq0 & v845647 | !hbusreq0 & v84561b;
assign v23fb6d7 = hgrant3_p & v84561b | !hgrant3_p & v22f3feb;
assign v23fb9cb = hmaster0_p & v230b00c | !hmaster0_p & v22f6bae;
assign v22f1a26 = hready & v22edf54 | !hready & v84561b;
assign v230d6ca = hmaster2_p & v2300af8 | !hmaster2_p & v22f1c57;
assign v23fc943 = hgrant3_p & v84561b | !hgrant3_p & v22f154e;
assign v23fc19b = hmaster2_p & v22fef4f | !hmaster2_p & v191a86f;
assign v23f329a = hgrant3_p & v23f3856 | !hgrant3_p & !v84561b;
assign v2309b5d = hmaster0_p & v23fc15f | !hmaster0_p & v23f2daf;
assign v23fc039 = hbusreq3_p & v23126b1 | !hbusreq3_p & v23074aa;
assign v22ffd0e = hmaster2_p & v23f5eb6 | !hmaster2_p & v84561b;
assign v22f9ebc = hmaster2_p & v22f3643 | !hmaster2_p & !v22f36ff;
assign v2300687 = hmaster1_p & v23fc005 | !hmaster1_p & v23933b0;
assign v22fafd7 = hlock2_p & v22f79fb | !hlock2_p & v230333f;
assign v23f1225 = hmaster2_p & v191aa68 | !hmaster2_p & v2392d6d;
assign v22f66b0 = hgrant1_p & v23fc5a4 | !hgrant1_p & v22fe4be;
assign v23fc0eb = hgrant6_p & v845635 | !hgrant6_p & v230677d;
assign v23f730d = hbusreq5_p & v1e83f7c | !hbusreq5_p & v23fc8ef;
assign v22fe73f = hgrant0_p & v23fc3f7 | !hgrant0_p & v23f7218;
assign v23fc551 = stateG10_5_p & v22fe7f5 | !stateG10_5_p & !v23fccbe;
assign v23fcbcd = hbusreq2_p & v230bed2 | !hbusreq2_p & v84561b;
assign v23fcbe2 = hgrant3_p & v84561b | !hgrant3_p & v2306e8f;
assign v23fc086 = hmaster2_p & v23fbfd0 | !hmaster2_p & v23fc7ee;
assign v23fc020 = hmaster2_p & v1e83fd9 | !hmaster2_p & v22fee46;
assign v23fc001 = hbusreq3 & v23f9c5f | !hbusreq3 & v84561b;
assign v23fba71 = hlock6_p & v2308609 | !hlock6_p & v84561b;
assign v23f99ec = hbusreq6 & v84564d | !hbusreq6 & v23f87f4;
assign c08bce = jx3_p & v23004ba | !jx3_p & v12cd540;
assign v22ffdc5 = hbusreq3_p & v22f61f6 | !hbusreq3_p & v23fc35f;
assign v2307ee4 = hbusreq2_p & v230aded | !hbusreq2_p & a1fba6;
assign v230a8eb = jx0_p & v22f7083 | !jx0_p & !v23f623e;
assign v230cff8 = hbusreq6_p & v23115a7 | !hbusreq6_p & v2306bc5;
assign v23fb576 = hbusreq0_p & v2311a1d | !hbusreq0_p & v22fc2eb;
assign v23fb4d3 = hlock1_p & v230c0b2 | !hlock1_p & v845620;
assign v23f9945 = jx2_p & v23fc2f2 | !jx2_p & v23fb88f;
assign b7029b = hbusreq5_p & v23f4b28 | !hbusreq5_p & v23fcc7a;
assign v2309e9d = hmaster2_p & v84561b | !hmaster2_p & v23fcf96;
assign v230b4b4 = hgrant3_p & fc8fdb | !hgrant3_p & v230e2bb;
assign v23f5240 = hgrant1_p & b50a75 | !hgrant1_p & v84561b;
assign v230bdad = hgrant3_p & v84562e | !hgrant3_p & v22edcf4;
assign v23f2e61 = hbusreq5 & v22eda43 | !hbusreq5 & v84561b;
assign v22fc517 = hlock0_p & v22f1b4e | !hlock0_p & !v23081f5;
assign v22ef507 = hmaster2_p & v23fbf9d | !hmaster2_p & v84564d;
assign v23fbbc0 = hbusreq6_p & v23928f2 | !hbusreq6_p & v23fc841;
assign v2311645 = hbusreq4_p & v22f968e | !hbusreq4_p & v230ae46;
assign v23fa392 = hmaster2_p & v23f9789 | !hmaster2_p & v22f8543;
assign v230d23a = locked_p & v23fc2d2 | !locked_p & !v84561b;
assign v230e618 = hmaster2_p & v23fbb5f | !hmaster2_p & v84561b;
assign v23fbea4 = hmaster1_p & v230a742 | !hmaster1_p & v239300d;
assign v23fc3f5 = hgrant5_p & v22eb3ad | !hgrant5_p & v22f84ff;
assign v23046be = hbusreq3_p & v23f9f9d | !hbusreq3_p & v84561b;
assign v23fc8d2 = hgrant5_p & v23fc388 | !hgrant5_p & v22ef469;
assign v23075dd = hbusreq4 & v2307f2b | !hbusreq4 & !v845622;
assign v230430f = hlock4_p & v84564d | !hlock4_p & !v23f60ba;
assign v23f1391 = hbusreq3_p & v23fb5b7 | !hbusreq3_p & !v84561b;
assign v22ecced = hgrant5_p & v23fba0c | !hgrant5_p & v23fbd3e;
assign v230648e = jx1_p & v23f0958 | !jx1_p & v23f82dd;
assign v22fa05c = hbusreq5_p & v22ee889 | !hbusreq5_p & v22ee26d;
assign v23f1eac = hgrant4_p & v23f5109 | !hgrant4_p & v22eb95e;
assign v239281b = hbusreq3 & bd762f | !hbusreq3 & v23f3f59;
assign v23f15ba = hgrant6_p & v23fb732 | !hgrant6_p & !v23f5f62;
assign v23f592f = hmaster1_p & v22f8cb9 | !hmaster1_p & v23117d2;
assign v191ab29 = hmaster2_p & v84561b | !hmaster2_p & v22f925b;
assign v23fc78b = hgrant5_p & v230297f | !hgrant5_p & v22f3c3d;
assign v22ff916 = hgrant1_p & v230e1a3 | !hgrant1_p & v2307779;
assign v23f8ecc = stateA1_p & v22f0362 | !stateA1_p & v2306775;
assign v2312be0 = hbusreq6 & v23f72fe | !hbusreq6 & v84561b;
assign v22feae3 = hgrant1_p & v12cd6a1 | !hgrant1_p & v230e4ae;
assign v23f44e8 = hmaster1_p & v230bd1c | !hmaster1_p & !v22fdf28;
assign v22fa3df = hbusreq3 & v22fea98 | !hbusreq3 & v84561b;
assign v23fb796 = hbusreq1_p & v23930d2 | !hbusreq1_p & v23fb980;
assign v22ffc83 = jx1_p & v230c91d | !jx1_p & v23f6079;
assign v2342fc3 = hlock2_p & v230e032 | !hlock2_p & v23022b1;
assign bfce54 = hlock6_p & v22f07bb | !hlock6_p & v23fb544;
assign v23fc8ac = jx3_p & v84561b | !jx3_p & v23fc4eb;
assign v22f3699 = hmaster0_p & v22f7914 | !hmaster0_p & v230f0de;
assign v23133a7 = hbusreq5_p & v84561b | !hbusreq5_p & v23fcce3;
assign v96bd8b = hgrant5_p & v84561b | !hgrant5_p & !v23f8798;
assign v23fbcc3 = hmaster0_p & a1fe40 | !hmaster0_p & v23f74da;
assign v22f947f = hbusreq4_p & v23f8a5e | !hbusreq4_p & v84561b;
assign v2312cd5 = hlock3_p & v2307942 | !hlock3_p & v84561b;
assign v2309bda = hmaster1_p & v23f0b4e | !hmaster1_p & v22f45ac;
assign v98c729 = hgrant3_p & v84562e | !hgrant3_p & v22f07cd;
assign v191a965 = jx2_p & v23f4a0f | !jx2_p & v22f8c8b;
assign v22eff53 = hmaster0_p & v22f1963 | !hmaster0_p & v23fb91d;
assign v2312580 = hbusreq1_p & v22f2efc | !hbusreq1_p & v84561b;
assign v23015c7 = hmaster0_p & v23111c7 | !hmaster0_p & v22fd827;
assign v2302136 = locked_p & v84561b | !locked_p & v23fc90f;
assign v23fcdc0 = hbusreq0_p & b9d00f | !hbusreq0_p & v22eda7c;
assign v23fc7a1 = jx1_p & v84561b | !jx1_p & v1aae6b5;
assign v23fc738 = hmaster0_p & v23fc4a8 | !hmaster0_p & v23f74bc;
assign v23f7344 = hbusreq6_p & v2391d0b | !hbusreq6_p & v230a775;
assign v23fb604 = hmaster0_p & v23f9307 | !hmaster0_p & !v239387a;
assign v22f98ca = hmaster1_p & v23fc684 | !hmaster1_p & v84561b;
assign v22febf8 = jx1_p & v22f4442 | !jx1_p & v23fcb57;
assign v23f1432 = hbusreq3 & v2303da9 | !hbusreq3 & v22fa628;
assign v23fd045 = hbusreq0 & v84561b | !hbusreq0 & v23009f0;
assign v2306ee6 = hmaster2_p & v23f069d | !hmaster2_p & v230a51c;
assign v23fcccd = hgrant0_p & v230f63f | !hgrant0_p & !v22ee750;
assign v23fb8e4 = hmaster2_p & v845627 | !hmaster2_p & v22f1faf;
assign v22ec6a7 = hmaster1_p & v23f43db | !hmaster1_p & v23116cd;
assign v22fcf52 = hgrant3_p & v22ee657 | !hgrant3_p & v22f8e09;
assign v230814d = hbusreq3_p & v84562e | !hbusreq3_p & !v22ee657;
assign v23f669d = hlock4_p & v22eb856 | !hlock4_p & v23f33c7;
assign v23f732a = stateA1_p & v23fcb89 | !stateA1_p & !v23fc8a3;
assign v22f166c = hlock2_p & v845661 | !hlock2_p & !v84561b;
assign v230b313 = hgrant5_p & v23f809b | !hgrant5_p & a1bfd6;
assign v231140b = hbusreq3 & v23fcd7f | !hbusreq3 & v84561b;
assign v23fb8f3 = hlock3_p & v1aada6e | !hlock3_p & v84561b;
assign v22eea52 = hbusreq6_p & v230e1e4 | !hbusreq6_p & v23130d9;
assign v1e845a7 = hbusreq4 & v22fe675 | !hbusreq4 & v84561b;
assign v23fc56f = hgrant2_p & f40aac | !hgrant2_p & v23fbf26;
assign v230fb0a = hbusreq3 & v230545b | !hbusreq3 & v230ea57;
assign v22ee5fb = hmaster2_p & v84561b | !hmaster2_p & b6c104;
assign v23f5461 = hgrant3_p & v22f536a | !hgrant3_p & v23f3e42;
assign v23fcb57 = hmaster1_p & v239223a | !hmaster1_p & v23fb545;
assign v23fcc3d = hmaster2_p & v191a879 | !hmaster2_p & !v23fcc36;
assign v22eb404 = hgrant1_p & v23fbd89 | !hgrant1_p & !v84561b;
assign b910da = jx2_p & v22f30bb | !jx2_p & v23fc548;
assign v23fc567 = hlock6_p & v22ecbf0 | !hlock6_p & v22f748c;
assign v22fec30 = hgrant1_p & v23389c8 | !hgrant1_p & v2303d95;
assign v22f32b9 = hbusreq6 & v22ef507 | !hbusreq6 & !v22fa4ea;
assign v23085c5 = jx1_p & v86c49f | !jx1_p & v22f2a85;
assign v22fe0a8 = hmaster2_p & v1506ffd | !hmaster2_p & !a39dae;
assign v23f7efd = hready & v84561b | !hready & v22f60c6;
assign v23facc9 = hgrant1_p & v2300d2f | !hgrant1_p & v22f0d2b;
assign v2306fba = hmaster2_p & v22f7d5d | !hmaster2_p & v22f0e00;
assign v22f988a = hlock3_p & v23fcc0c | !hlock3_p & v2309c93;
assign v23fc6f7 = stateG10_5_p & v2313618 | !stateG10_5_p & e1dd6a;
assign v230fe82 = hgrant3_p & v22f6ae5 | !hgrant3_p & v23f62d5;
assign v23f1c14 = hbusreq3_p & v230607d | !hbusreq3_p & afffd9;
assign v2312ba0 = hmaster0_p & v22f8613 | !hmaster0_p & v22eaeaf;
assign v2304b49 = hmaster2_p & v106ae19 | !hmaster2_p & v230f848;
assign v2303b9a = hgrant2_p & v23f6411 | !hgrant2_p & !v106ae19;
assign v2393527 = hlock3_p & v23fbac3 | !hlock3_p & v1e840fa;
assign v22eb2fd = hbusreq6 & v22fc4a3 | !hbusreq6 & v2393742;
assign v23052dd = hmaster1_p & v23fc69f | !hmaster1_p & v23fd00e;
assign v230648c = hmaster2_p & c24eac | !hmaster2_p & v23f7d57;
assign v23135cc = hmaster2_p & v22f9c2f | !hmaster2_p & !v23109c3;
assign v2300aa8 = hbusreq4 & v23057ba | !hbusreq4 & v84561b;
assign v22f679a = hmaster2_p & v230f537 | !hmaster2_p & v84561b;
assign v22ed7a8 = locked_p & v230e58e | !locked_p & !v106ae19;
assign v230216e = hmaster2_p & v23f8f25 | !hmaster2_p & v23919f9;
assign v22eed68 = hgrant3_p & v2305d6f | !hgrant3_p & v230dcba;
assign a6a2f9 = hbusreq5_p & v22f3999 | !hbusreq5_p & v22fd2e2;
assign v2306292 = hbusreq3 & v22ec66d | !hbusreq3 & v2302f85;
assign v23f66ec = hbusreq3_p & v23fba45 | !hbusreq3_p & v2313131;
assign v2393abe = hgrant3_p & v23f5cd3 | !hgrant3_p & v22ff9d4;
assign v23060d4 = hbusreq5_p & v2305af1 | !hbusreq5_p & v84561b;
assign v22f5e57 = hgrant5_p & v22fa05c | !hgrant5_p & v23041c3;
assign v23fbe22 = hgrant1_p & v84564d | !hgrant1_p & v22eaaef;
assign v23f5057 = hbusreq3 & v23fb865 | !hbusreq3 & v84562a;
assign v23025ab = hlock2_p & v23f8364 | !hlock2_p & v84561b;
assign v2303c39 = hbusreq5 & v1aad518 | !hbusreq5 & v8d030a;
assign v17cf286 = decide_p & v230c771 | !decide_p & v23fb9d4;
assign v230d2a8 = hmastlock_p & v23f6d93 | !hmastlock_p & v84561b;
assign v22ed56a = start_p & v84561b | !start_p & !v845663;
assign v23f1bbf = hgrant1_p & v23fc904 | !hgrant1_p & v23fced8;
assign v2312696 = hbusreq5_p & v22fb17b | !hbusreq5_p & v84561b;
assign v23f24d1 = hgrant1_p & v845626 | !hgrant1_p & v22f923c;
assign v22fc61a = hgrant5_p & v22fb051 | !hgrant5_p & !v230848d;
assign v23fca43 = hmaster0_p & v22f4c34 | !hmaster0_p & b00ac7;
assign v1506fbf = hbusreq5 & v22ee0c4 | !hbusreq5 & v84561b;
assign v23f4154 = hbusreq1 & v23fc48b | !hbusreq1 & v84561b;
assign v23fc09c = hmaster0_p & v23fbf49 | !hmaster0_p & !v23fbe77;
assign v23008c7 = hmaster2_p & v12cd68e | !hmaster2_p & v22eb3e3;
assign a8b64b = hlock6_p & v23fcea0 | !hlock6_p & v84562b;
assign v23f9e4f = hbusreq5_p & v2308f46 | !hbusreq5_p & v84561b;
assign v191ad2f = hbusreq5_p & v22fe0c1 | !hbusreq5_p & v845623;
assign v22f1697 = hmaster2_p & v84561b | !hmaster2_p & v2309891;
assign v22fb427 = stateG2_p & v84561b | !stateG2_p & v912a31;
assign v23fb5f1 = hbusreq6_p & v23f6c7c | !hbusreq6_p & v22ec39f;
assign v23045fb = hbusreq1 & v23f8da8 | !hbusreq1 & v23f1d35;
assign v22ee0e1 = stateG2_p & v84561b | !stateG2_p & v22f39a1;
assign v2305507 = hmaster2_p & v23fcf69 | !hmaster2_p & v23919f9;
assign v1aad67e = hgrant3_p & v22f5088 | !hgrant3_p & !v84561b;
assign v231009b = hgrant2_p & v2309cb5 | !hgrant2_p & v23022b1;
assign v22ef270 = hbusreq6 & v230de81 | !hbusreq6 & v22fce8b;
assign v23f70cf = hbusreq3_p & v23fbb64 | !hbusreq3_p & v2309320;
assign v23f7688 = hbusreq3 & v2310051 | !hbusreq3 & aeff78;
assign v23fc957 = hgrant1_p & v845625 | !hgrant1_p & v23108a7;
assign v23fc0a4 = hbusreq3 & v22f05b9 | !hbusreq3 & !v84562a;
assign v22f79c8 = hlock4_p & v191abfa | !hlock4_p & !v84561b;
assign v22f63e8 = stateG2_p & v23023b3 | !stateG2_p & !v230ec21;
assign v23102f3 = hmaster0_p & v2306875 | !hmaster0_p & v23f3545;
assign v1e84184 = hbusreq5 & v23fcc10 | !hbusreq5 & v84561b;
assign v22fc963 = hmaster2_p & v23f3d14 | !hmaster2_p & v84561b;
assign v22f7ee5 = hbusreq6 & v23fca10 | !hbusreq6 & v230f0de;
assign v22ec335 = hbusreq0_p & v22eccee | !hbusreq0_p & !v845629;
assign v22fa6c0 = hbusreq6_p & v230339f | !hbusreq6_p & v23f5fe3;
assign v23fcd42 = hmaster0_p & v22f6629 | !hmaster0_p & !v23fa94e;
assign v23fba97 = hbusreq1 & v23f9789 | !hbusreq1 & v84561b;
assign v23faa39 = jx1_p & v22f19dd | !jx1_p & v22edf86;
assign v23fbadc = hbusreq1 & v230358b | !hbusreq1 & v22f8d74;
assign v22ef509 = hbusreq0 & v230882d | !hbusreq0 & !v84561b;
assign v22eb664 = hbusreq3_p & v22f2bab | !hbusreq3_p & v1aae9a1;
assign v23fafe3 = hbusreq6 & v23930d8 | !hbusreq6 & !v230efee;
assign v230960c = hgrant3_p & v84561b | !hgrant3_p & v22fb6db;
assign v23f89d9 = hbusreq6 & v22f2e9f | !hbusreq6 & v22f2623;
assign v23f6b11 = hgrant1_p & v845626 | !hgrant1_p & v23fb9b7;
assign v22ebc25 = hgrant3_p & v22f6c3a | !hgrant3_p & v230813c;
assign v23fb52f = hmaster0_p & v23f9737 | !hmaster0_p & v22fac35;
assign v23f78df = hbusreq4_p & v22f15ef | !hbusreq4_p & v23fc61d;
assign v22fdb4e = hmastlock_p & v12cd993 | !hmastlock_p & v84561b;
assign v23f85b5 = hmaster0_p & v22f4062 | !hmaster0_p & b00aa6;
assign v22feec8 = hmaster2_p & v22f54a4 | !hmaster2_p & v22f30df;
assign v230591e = hgrant3_p & v2303ae8 | !hgrant3_p & v8bbb53;
assign v23fc810 = hbusreq3 & v23fcfaa | !hbusreq3 & v22fdb5c;
assign v22ebce1 = hmaster2_p & v22f926d | !hmaster2_p & v13afb18;
assign v22fb6db = hmaster2_p & v22f9078 | !hmaster2_p & !v230f43d;
assign v23fbed7 = hbusreq4 & v230eb5a | !hbusreq4 & v22f061c;
assign v2302fbc = hbusreq3 & v23f363f | !hbusreq3 & v84561b;
assign v23016dc = hbusreq4_p & v230430f | !hbusreq4_p & !v23f60ba;
assign v2392258 = hmaster2_p & v23fba6b | !hmaster2_p & v23f65b4;
assign v230b089 = hgrant0_p & v22ff106 | !hgrant0_p & a476c2;
assign v22fb7bc = hbusreq2_p & v23f43af | !hbusreq2_p & v84564d;
assign v230f5ee = hbusreq5_p & v23fc530 | !hbusreq5_p & v23fc4f7;
assign v23f8180 = hmaster1_p & v22f4828 | !hmaster1_p & !v23f49cd;
assign v1aad5a0 = hbusreq1 & v23fc799 | !hbusreq1 & v22f7241;
assign v23fc46d = hmaster2_p & v2391d40 | !hmaster2_p & !v23f763f;
assign v23fc4a2 = hbusreq6_p & v23051a9 | !hbusreq6_p & v22f76b3;
assign v23fcd74 = hmaster2_p & b9d0d2 | !hmaster2_p & !v953acf;
assign v22f4339 = hmaster1_p & v23fc989 | !hmaster1_p & v22ee8ee;
assign v23f79a7 = hmaster2_p & v23fbda4 | !hmaster2_p & v2301e66;
assign v230aabf = hgrant4_p & v2303632 | !hgrant4_p & !v22f4bf5;
assign v23135ec = hbusreq4 & v22ecaeb | !hbusreq4 & v23fcaa5;
assign v22f39af = hlock5_p & v2301312 | !hlock5_p & v22f3692;
assign v230fec6 = hbusreq2_p & v84561b | !hbusreq2_p & !v106a782;
assign v23f6411 = locked_p & a1fbb6 | !locked_p & !v106ae19;
assign v2313618 = hgrant0_p & v22f5605 | !hgrant0_p & !v22f753d;
assign v23fc48f = hmaster2_p & v22ec9fa | !hmaster2_p & v84561b;
assign v23fcf2d = stateG10_5_p & v230828c | !stateG10_5_p & v230b8cd;
assign v23f4160 = hbusreq4_p & v2392ff9 | !hbusreq4_p & v99b664;
assign v2300070 = jx0_p & v230c213 | !jx0_p & c08bce;
assign v1aad703 = hbusreq4_p & v22eb0b3 | !hbusreq4_p & v23f62ee;
assign v23022d5 = hlock4_p & v2311b9e | !hlock4_p & !v23069b0;
assign v2303a32 = hmaster0_p & v23fcf87 | !hmaster0_p & v23fcf0e;
assign v23081eb = busreq_p & v22f4cca | !busreq_p & v23f4067;
assign v22fb95e = hgrant0_p & v191b187 | !hgrant0_p & !v84561b;
assign v23f2d1d = hbusreq3_p & v230e618 | !hbusreq3_p & v23f2b21;
assign v1aad6c8 = stateG2_p & v84561b | !stateG2_p & v22f7176;
assign v23fc063 = hmaster0_p & af7272 | !hmaster0_p & v22efc9e;
assign v22eefcf = hmaster2_p & v23fc742 | !hmaster2_p & v23fcb55;
assign v230727f = hbusreq3_p & v22ec1ae | !hbusreq3_p & v22fa934;
assign v22f11fe = hgrant1_p & v23f4491 | !hgrant1_p & v2300cb6;
assign v230cf2f = hmaster2_p & v2308d79 | !hmaster2_p & !v23fc514;
assign v23f89fd = hmaster0_p & v23f54f7 | !hmaster0_p & v23fc410;
assign v23fb477 = stateG2_p & v2302ca3 | !stateG2_p & !v23faacf;
assign v22edc8d = hlock0_p & v106ae1c | !hlock0_p & a1fbb6;
assign v2392fc4 = hbusreq6 & v22fc90d | !hbusreq6 & !v230df81;
assign v22f881b = hmaster2_p & v22ed878 | !hmaster2_p & v23fd050;
assign v230b6d9 = hmaster0_p & v84561b | !hmaster0_p & v23fd01f;
assign v2304764 = hmaster1_p & v84561b | !hmaster1_p & v22f9f68;
assign v2303674 = hbusreq3_p & v23f8bef | !hbusreq3_p & v84561b;
assign v22f35e8 = hlock0_p & v191aa68 | !hlock0_p & v230d24a;
assign v22f8dea = stateG10_5_p & v2305de3 | !stateG10_5_p & v23fb67c;
assign v23f8b2b = jx2_p & v23fc5ca | !jx2_p & v23fb50c;
assign v22f358f = hbusreq5_p & v2303046 | !hbusreq5_p & !v84561b;
assign v2309532 = hmaster1_p & v2311b7c | !hmaster1_p & v230a3b3;
assign v22f41ab = hmaster0_p & v231345a | !hmaster0_p & v23f5bf7;
assign v22ef255 = hmaster0_p & v22f6917 | !hmaster0_p & !v17a34ff;
assign v2308669 = hmaster0_p & v22f6e67 | !hmaster0_p & v230aa0b;
assign v23fb4ae = hbusreq5 & v2304ec7 | !hbusreq5 & !v84561b;
assign v22f7f74 = hmastlock_p & v23fc331 | !hmastlock_p & v84561b;
assign v23f2c35 = hbusreq6_p & v2304d08 | !hbusreq6_p & v23fce02;
assign v23fc517 = hgrant4_p & v23f6789 | !hgrant4_p & v23fc4ef;
assign v23f2862 = busreq_p & v106a7a0 | !busreq_p & v22ef0b3;
assign v15071c2 = hlock2_p & v13afe3a | !hlock2_p & !v84561b;
assign v23f8caa = hbusreq3_p & v23f9395 | !hbusreq3_p & v22f14bf;
assign v230b7c1 = hbusreq0 & v23fbb74 | !hbusreq0 & v84561b;
assign v22feb04 = hmaster0_p & v2312189 | !hmaster0_p & !v230fe87;
assign v23f69cd = hmaster2_p & v22f15b7 | !hmaster2_p & v23f7f8d;
assign bb324c = hmaster2_p & v84561b | !hmaster2_p & v23fb883;
assign v23fcae0 = hbusreq3 & v2304ccc | !hbusreq3 & v84561b;
assign v22f76b3 = hbusreq4_p & v23051a9 | !hbusreq4_p & v23fbd5b;
assign v2307b42 = hbusreq6_p & v230d91f | !hbusreq6_p & v22ff29c;
assign v23f614a = stateG10_5_p & v23fc338 | !stateG10_5_p & v84561b;
assign v22ffbb3 = hlock0_p & v23f6411 | !hlock0_p & v2309a78;
assign v23fc6c2 = hbusreq3 & v23f60fb | !hbusreq3 & !v84561b;
assign v23fbb74 = hmastlock_p & v22ec1cb | !hmastlock_p & v84561b;
assign v230deb1 = hmaster1_p & v23fb681 | !hmaster1_p & !v23f49cd;
assign v191b1ae = hmaster0_p & e1e6ee | !hmaster0_p & v2307d93;
assign v22eb2a2 = hbusreq1 & v23fc7b2 | !hbusreq1 & v22ff090;
assign v23fc3f3 = hmaster0_p & v23fbd48 | !hmaster0_p & !v230d00c;
assign v23fb583 = hmaster2_p & v23fba65 | !hmaster2_p & v230c727;
assign v23fb98b = hmaster1_p & v22ff244 | !hmaster1_p & v230fd1b;
assign v22f4626 = hbusreq3 & v22ee1b8 | !hbusreq3 & v23fc79d;
assign ab5bb8 = hlock2_p & fc8ab7 | !hlock2_p & v84561b;
assign b00aa0 = hmaster2_p & v22ff05e | !hmaster2_p & !v22f1d80;
assign v23050a2 = hbusreq3_p & v22f2429 | !hbusreq3_p & v23f76f4;
assign v1506f9f = hmaster2_p & v230d2c2 | !hmaster2_p & v22f17ca;
assign v23fb80e = stateG10_5_p & v23fc374 | !stateG10_5_p & v22fdc30;
assign v23fceb9 = hbusreq2_p & v2300d6c | !hbusreq2_p & v84561b;
assign v23fb12f = hbusreq3 & v23fc99a | !hbusreq3 & v230a70a;
assign v22eff6d = hbusreq5_p & v23fb619 | !hbusreq5_p & v84561b;
assign v23f51b1 = hgrant2_p & v23f76c2 | !hgrant2_p & !v106ae19;
assign v1507056 = hlock0_p & v2307b18 | !hlock0_p & v230083b;
assign v22fde54 = hmaster2_p & v845622 | !hmaster2_p & v23fc596;
assign v2308b9a = hmaster0_p & v22f368e | !hmaster0_p & v23fc2dc;
assign v2308bbe = hbusreq0_p & v1aae56f | !hbusreq0_p & v13affaa;
assign v191b17f = hgrant3_p & v84561b | !hgrant3_p & v23fcd5f;
assign v23f5bf7 = hgrant3_p & v84561b | !hgrant3_p & a04dcc;
assign v23fce08 = hmaster1_p & v23fb70e | !hmaster1_p & v22f7728;
assign v2310bf5 = hlock1_p & v1aae087 | !hlock1_p & !v84561b;
assign v2305dde = hmaster0_p & v230502a | !hmaster0_p & v23fba85;
assign v23fc9f3 = hbusreq1 & v23f45d2 | !hbusreq1 & v84561b;
assign v230e896 = hmaster1_p & v23f0dc7 | !hmaster1_p & a1fdd3;
assign v2311524 = hgrant3_p & v23fcab6 | !hgrant3_p & v22ef750;
assign v15070e0 = hbusreq2 & v15071c2 | !hbusreq2 & !v23095fa;
assign v2302149 = hbusreq2_p & v9526ac | !hbusreq2_p & a1fba6;
assign v230edb2 = hmaster0_p & v23035b0 | !hmaster0_p & v230e831;
assign v22fec56 = hbusreq3 & v230ca57 | !hbusreq3 & v22f5cf0;
assign v22f9dfb = hmaster2_p & v845620 | !hmaster2_p & v22f8cb7;
assign v2309aaa = stateG10_5_p & v22f6a93 | !stateG10_5_p & !v84561b;
assign v845661 = stateG2_p & v84561b | !stateG2_p & !v84561b;
assign f40764 = jx0_p & v22ffa07 | !jx0_p & v84561b;
assign v2309b7e = hbusreq1_p & v1506ffd | !hbusreq1_p & v22f3fec;
assign v22fcb45 = hmaster2_p & v23027bf | !hmaster2_p & v84561b;
assign v230e9ef = hmaster2_p & v1aae362 | !hmaster2_p & v84561b;
assign v23f0178 = hmaster2_p & v22efae1 | !hmaster2_p & v22eeb07;
assign v22f9add = hmaster2_p & v9d8aae | !hmaster2_p & v2306220;
assign v23fbbc9 = hlock5_p & v23fb798 | !hlock5_p & !v84561b;
assign v22fe9b7 = locked_p & v22fef4f | !locked_p & v23fba6b;
assign v1e84072 = hbusreq3_p & bc65c8 | !hbusreq3_p & v23f3ac9;
assign c16191 = hbusreq0 & v23fcbcd | !hbusreq0 & v23fbffc;
assign v23fcb09 = jx1_p & v2392eb5 | !jx1_p & v23082c9;
assign v2303376 = hbusreq0 & v23105cd | !hbusreq0 & v2312bd0;
assign v23fbfc9 = hlock1_p & v23fc7e6 | !hlock1_p & v845620;
assign v23122b0 = jx2_p & v22f6d51 | !jx2_p & a7e154;
assign v23fc55d = hbusreq5 & v23f450d | !hbusreq5 & v84561b;
assign v230075e = hbusreq5_p & v23126c6 | !hbusreq5_p & v22ee9be;
assign v23f660f = hgrant1_p & v12cc2ef | !hgrant1_p & v22f9b95;
assign v23fb483 = hgrant3_p & v84562e | !hgrant3_p & v22f8afa;
assign v23fb23b = hbusreq3_p & v22fd825 | !hbusreq3_p & v22f8463;
assign v23919d4 = hgrant5_p & v23fbc06 | !hgrant5_p & v2304339;
assign v23fc267 = hlock4_p & v22eaf66 | !hlock4_p & v2310969;
assign v22fa002 = hgrant0_p & v2393b93 | !hgrant0_p & v84561b;
assign v23f1861 = hbusreq5_p & v23f5c95 | !hbusreq5_p & !v23fc3a1;
assign v230b125 = hbusreq5_p & v23fc1d2 | !hbusreq5_p & !v84561b;
assign v17a2d5a = hready_p & v2309543 | !hready_p & v21eabbd;
assign v23fbd13 = hmaster0_p & v2303ebc | !hmaster0_p & v23f082a;
assign bd7747 = hlock0_p & v22f037a | !hlock0_p & !v84561b;
assign v23fd019 = hbusreq3_p & v23f60fb | !hbusreq3_p & v23fbd28;
assign v22f1a1b = hbusreq0_p & v22ed6ee | !hbusreq0_p & v84561b;
assign v22eb14c = jx1_p & v22fbaf1 | !jx1_p & !v22fbd0e;
assign v191ae6a = hbusreq2 & v22fc4d3 | !hbusreq2 & v2393116;
assign v23f6789 = jx0_p & v230c32e | !jx0_p & v22fc493;
assign v23fcc1f = hbusreq5_p & v23fcf1f | !hbusreq5_p & v845620;
assign v2391ada = hgrant0_p & v23fc22d | !hgrant0_p & !v22f69b7;
assign v2302d97 = hbusreq2_p & v2304910 | !hbusreq2_p & v84561b;
assign v23fbd71 = hmaster0_p & v23f2bb6 | !hmaster0_p & v22fee9e;
assign v230f549 = hmaster0_p & v2304a06 | !hmaster0_p & !v23025e4;
assign v22f8959 = hbusreq2_p & v23f43af | !hbusreq2_p & v23fbec8;
assign v23081e8 = hlock3_p & v23f4540 | !hlock3_p & v230664e;
assign v23fca59 = hlock6_p & v23fcb63 | !hlock6_p & v230994d;
assign v23fa524 = hburst0 & v23fb564 | !hburst0 & !v84561b;
assign v230f1a7 = hgrant2_p & v12cd523 | !hgrant2_p & !v150755e;
assign v23139c9 = hmaster0_p & v22f8cb9 | !hmaster0_p & v23f76fb;
assign v23fbaaa = hgrant1_p & v22eb377 | !hgrant1_p & v22f3b3c;
assign v2311374 = hbusreq5_p & v22f9927 | !hbusreq5_p & v23fb900;
assign v230ca71 = hready_p & v23f5558 | !hready_p & v23fbdc6;
assign v2304443 = hbusreq1_p & v23f4f34 | !hbusreq1_p & v84561b;
assign v23fba25 = hbusreq1_p & v23f79d2 | !hbusreq1_p & !v84561b;
assign v2313405 = hbusreq3_p & v2304669 | !hbusreq3_p & v84561b;
assign v22f8857 = hmaster2_p & v22ecba3 | !hmaster2_p & v23f3206;
assign v22fed78 = hmaster2_p & v84561b | !hmaster2_p & v23f5c95;
assign v231049c = hmaster2_p & v22f8aec | !hmaster2_p & v84561b;
assign v22f61bb = hmaster2_p & v230a92e | !hmaster2_p & v23f87f4;
assign v22fbdbc = hlock3_p & v23010b3 | !hlock3_p & v23fc753;
assign v22f779f = hmaster2_p & v84561b | !hmaster2_p & !v13afe3a;
assign a4c73f = jx2_p & v23fc403 | !jx2_p & bdab35;
assign v2306790 = hmaster0_p & v22eba1d | !hmaster0_p & v2307c3d;
assign v9aa6cf = hbusreq6_p & v231329e | !hbusreq6_p & !v84561b;
assign v22faf11 = hready_p & v1aad3bf | !hready_p & !v84561b;
assign v22fb77d = hbusreq0_p & v2305196 | !hbusreq0_p & v84561b;
assign v230d793 = stateG10_5_p & v22ef725 | !stateG10_5_p & !v230ebff;
assign v23f51ac = hmaster0_p & v23fcb9f | !hmaster0_p & v23fcb40;
assign v22f1e0b = hbusreq0_p & v23f50e0 | !hbusreq0_p & v84561b;
assign v23fb28e = hbusreq1 & v2306932 | !hbusreq1 & !v23f4722;
assign v23f5e84 = hmaster0_p & v2391d2f | !hmaster0_p & v23fcfc4;
assign v2304d7a = hlock3_p & v22eb75e | !hlock3_p & !v2312e04;
assign v23f5927 = hbusreq3_p & v22f0a19 | !hbusreq3_p & !v84561b;
assign v2305f49 = hmaster0_p & v23f88e6 | !hmaster0_p & v23f93b5;
assign v22fb2c5 = hbusreq3_p & v23fce4e | !hbusreq3_p & v84561b;
assign v23f6c84 = hgrant1_p & v12cc2f8 | !hgrant1_p & v23087b6;
assign v2303d9e = hbusreq6_p & v230a6c8 | !hbusreq6_p & !v23113f5;
assign v2306119 = hbusreq6_p & v23fce89 | !hbusreq6_p & v23fb9bf;
assign v230bf1e = hbusreq4_p & v22ed933 | !hbusreq4_p & v23fbf6b;
assign v106af28 = hbusreq6_p & v23fbc0c | !hbusreq6_p & v22f2ee3;
assign v23117cd = hmaster0_p & v22ff6c5 | !hmaster0_p & v23fbd19;
assign v22feb6b = hmaster2_p & v22f8b01 | !hmaster2_p & v22f5815;
assign v23f6949 = hmaster2_p & v106a782 | !hmaster2_p & v22f92fa;
assign v22f04eb = hmaster1_p & v22edd99 | !hmaster1_p & b00aa6;
assign v23fcc2a = hmaster0_p & v84564d | !hmaster0_p & v2302992;
assign v23f651a = hbusreq3_p & v84564d | !hbusreq3_p & !v84561b;
assign v23f15ac = hbusreq5_p & v23f4d58 | !hbusreq5_p & v84561b;
assign v23fc999 = hbusreq6 & v23fbce1 | !hbusreq6 & v23fca2f;
assign v23f9110 = hbusreq3_p & v23fc96d | !hbusreq3_p & v23fc85e;
assign v230d532 = hmaster0_p & v23fbaed | !hmaster0_p & v23fbbbe;
assign v22f5992 = hgrant3_p & v22f8e29 | !hgrant3_p & v23fbd34;
assign v231220c = hmaster1_p & v23fbf8d | !hmaster1_p & v22f88bb;
assign v23f9492 = hbusreq4 & v22ed400 | !hbusreq4 & v230f96f;
assign v22f26f5 = hbusreq3_p & v22f61f6 | !hbusreq3_p & v230bd36;
assign v22f14ed = hgrant5_p & v23fb24f | !hgrant5_p & v22ef945;
assign v22ef7a7 = jx0_p & v22f6d27 | !jx0_p & v2312bae;
assign v230c7f6 = hbusreq6_p & v23fc5f5 | !hbusreq6_p & v22fdaf3;
assign v23fc6a6 = hmaster1_p & v22fab7b | !hmaster1_p & v84561b;
assign v230fe54 = hbusreq6_p & v23fa3e0 | !hbusreq6_p & !v84561b;
assign v22ef757 = hbusreq6_p & v23f4f88 | !hbusreq6_p & v2312050;
assign v23f9ba6 = hmaster2_p & v23919f9 | !hmaster2_p & v84561b;
assign v23fa0aa = hgrant1_p & v22f3ed0 | !hgrant1_p & v22fc5ad;
assign v2391dd6 = hmaster1_p & v23fbb9e | !hmaster1_p & v22ed4b0;
assign v22ed881 = hbusreq3_p & v23fbbb9 | !hbusreq3_p & v23fb583;
assign v8f530a = hbusreq1_p & v84561b | !hbusreq1_p & v1aae087;
assign v1aad641 = hmaster2_p & v12cc2ef | !hmaster2_p & !v23f328e;
assign v22fc9bf = hgrant1_p & v22f7d5d | !hgrant1_p & !v23108aa;
assign v23fb1e3 = stateG10_5_p & v23fbed3 | !stateG10_5_p & v22ece03;
assign v23fc81c = stateG10_5_p & v23fc619 | !stateG10_5_p & v23fa2ec;
assign v22fa156 = hgrant1_p & v23f761c | !hgrant1_p & v22fcd7c;
assign v23fc0bf = hbusreq4_p & v22fdf3c | !hbusreq4_p & v22f125c;
assign v2300dcb = hmaster0_p & v22f2f3e | !hmaster0_p & v2302460;
assign v23f54f7 = hbusreq6 & v23fc48f | !hbusreq6 & v23fcc2e;
assign v23f4edc = hgrant3_p & v230200a | !hgrant3_p & v2391d99;
assign v23f8914 = hbusreq2 & v23131e8 | !hbusreq2 & v2306220;
assign v23fcb24 = hbusreq3 & v230dcf6 | !hbusreq3 & v84561b;
assign v23fb9c5 = hlock1_p & v22fc8e5 | !hlock1_p & v2309c93;
assign v2306f00 = stateG10_5_p & v22f6058 | !stateG10_5_p & v230aded;
assign v22fd2ac = hbusreq6 & v22edb40 | !hbusreq6 & v22efbd5;
assign v23fb931 = hgrant3_p & v230630c | !hgrant3_p & v239228f;
assign v22f2623 = hbusreq3_p & e1bfb3 | !hbusreq3_p & v230bd8f;
assign v22f9188 = hmaster1_p & v238aeb0 | !hmaster1_p & v23f1686;
assign v23f445f = hlock1_p & v845620 | !hlock1_p & !v84561b;
assign v23f93e7 = hmaster2_p & v22f17ca | !hmaster2_p & v23fc5ff;
assign v23f35ff = hmaster2_p & v1aadb8e | !hmaster2_p & v23fc346;
assign v23fced8 = hgrant5_p & v22f9049 | !hgrant5_p & !v1aad3ae;
assign v23fc2bc = hmaster0_p & v22ef848 | !hmaster0_p & v84561b;
assign v2301509 = hlock1_p & v23fb590 | !hlock1_p & v84564d;
assign v22f99e9 = hmaster2_p & v23fb1c6 | !hmaster2_p & v22ff732;
assign v230bdbb = stateG10_5_p & v22fbfaf | !stateG10_5_p & v23fb67c;
assign v23f7b32 = hgrant3_p & v84561b | !hgrant3_p & v23fc469;
assign v2312189 = hbusreq3_p & v23044cf | !hbusreq3_p & v23f41b9;
assign v2300c80 = hlock0_p & v2310104 | !hlock0_p & v2302868;
assign v22f8f49 = hlock4_p & v2309b80 | !hlock4_p & v23fa6eb;
assign v22f2d26 = hmaster2_p & v2304074 | !hmaster2_p & v22ff732;
assign v2305114 = hbusreq0_p & v23f6ba0 | !hbusreq0_p & v2309891;
assign v2312c13 = hgrant1_p & v22f7830 | !hgrant1_p & v2309943;
assign hmaster1 = v10dbf78;
assign v845621 = hbusreq0_p & v84561b | !hbusreq0_p & !v84561b;
assign v22fed24 = hgrant5_p & v230e851 | !hgrant5_p & !v231050f;
assign v23fc092 = hgrant3_p & v2310482 | !hgrant3_p & v23fcdde;
assign v22fee3b = hbusreq1_p & v230a355 | !hbusreq1_p & v84561b;
assign v8a6d1a = hmaster0_p & v22ef823 | !hmaster0_p & v22f346d;
assign v22f8c0b = hgrant5_p & v84561b | !hgrant5_p & !v22fb71d;
assign v2306a5d = hbusreq1 & v23f6836 | !hbusreq1 & v84564d;
assign v230ff42 = hbusreq5_p & v23fbb0b | !hbusreq5_p & !v23fbc20;
assign v230aca2 = hmaster2_p & v230b981 | !hmaster2_p & b60876;
assign v22fbe28 = hbusreq5_p & v845636 | !hbusreq5_p & !v84561b;
assign v23fb809 = hgrant5_p & v84561b | !hgrant5_p & v22ffa10;
assign v23fb1c5 = hlock3_p & v231363a | !hlock3_p & v1aad6a6;
assign v23f4f43 = hmaster0_p & v22f84f8 | !hmaster0_p & v22ec64d;
assign v22f5378 = jx0_p & v2308980 | !jx0_p & v22fcf35;
assign v2311b7c = hbusreq6_p & v2307eb9 | !hbusreq6_p & v23fb66f;
assign v23f6d19 = hbusreq1_p & v230f75a | !hbusreq1_p & !v2392077;
assign v23130b0 = hmaster2_p & v22f0add | !hmaster2_p & v230cbdd;
assign v230a573 = hbusreq3 & v903f7f | !hbusreq3 & v22ebe99;
assign v22fb417 = hbusreq4 & v23045ae | !hbusreq4 & v23fb922;
assign v2309bcf = hmaster1_p & v84561b | !hmaster1_p & !v22ed55a;
assign v23066df = hbusreq2_p & fc8ab7 | !hbusreq2_p & v22f9a51;
assign v23fb569 = hmaster0_p & v22ede34 | !hmaster0_p & !v23f5c60;
assign v22f98ad = hbusreq1 & v23fcac8 | !hbusreq1 & v84561b;
assign v23f7a8e = hmaster1_p & v22eddf2 | !hmaster1_p & v22f01b2;
assign v2307320 = hbusreq3 & v22f9f33 | !hbusreq3 & v84561b;
assign v2311c4d = hbusreq1_p & v22fe421 | !hbusreq1_p & v22fc8c8;
assign v2308a4c = hmastlock_p & v23069f2 | !hmastlock_p & v84561b;
assign v23fb4e8 = hmaster2_p & fc8ab7 | !hmaster2_p & v84561b;
assign v22f1d7b = jx2_p & v2309aca | !jx2_p & v22f65e3;
assign v23fb56e = hgrant2_p & v231086f | !hgrant2_p & !v2301d10;
assign v2311031 = hbusreq6_p & v22eb2ee | !hbusreq6_p & !fc8c53;
assign v22f50bf = hlock2_p & v2312ea7 | !hlock2_p & v230f654;
assign v22fdc20 = jx0_p & v2302a57 | !jx0_p & v23fa69e;
assign v22fb36e = hmaster2_p & v22f94ec | !hmaster2_p & v22fee3b;
assign v230810c = hgrant3_p & v23fb504 | !hgrant3_p & b194d1;
assign v23fc689 = hmaster0_p & bd8ccb | !hmaster0_p & v23f6bba;
assign v23128ab = hmaster2_p & v23fcac2 | !hmaster2_p & v1aad481;
assign v22ff414 = hbusreq5_p & v845620 | !hbusreq5_p & v22f79fd;
assign v23fcd03 = hbusreq3_p & v23fceb9 | !hbusreq3_p & v23fc746;
assign v23fcd90 = hlock3_p & v191ae90 | !hlock3_p & v230042c;
assign v23fc0c3 = hlock6_p & v2308aa9 | !hlock6_p & v23fb808;
assign v22f25fa = hbusreq4_p & v23f9bf9 | !hbusreq4_p & v23fb790;
assign v23107fc = hmaster2_p & v2310754 | !hmaster2_p & v191abc5;
assign v23fb9ac = hlock2_p & v230358b | !hlock2_p & v23f7efd;
assign a1382d = hlock5_p & v23fb942 | !hlock5_p & v2301f52;
assign v22f6bd4 = hmastlock_p & v23f2278 | !hmastlock_p & v84561b;
assign v22f5e36 = stateG10_5_p & v23f79a0 | !stateG10_5_p & v845636;
assign v23fbf58 = hmaster2_p & v84564d | !hmaster2_p & v2300c3d;
assign v22fac35 = hbusreq6 & v23f9c5f | !hbusreq6 & v84561b;
assign v22ee8dd = hmaster0_p & v23051cf | !hmaster0_p & v84561b;
assign v22f8aeb = hbusreq2 & v23fcc10 | !hbusreq2 & v230e547;
assign v22eb9b4 = hlock3_p & v230538c | !hlock3_p & !v1aad4c6;
assign v22f82ea = hmaster1_p & v239345a | !hmaster1_p & v22f0ceb;
assign v23fc254 = hgrant2_p & v84562a | !hgrant2_p & v23f5043;
assign v8f2065 = hlock5_p & v22fc8e5 | !hlock5_p & v2309c93;
assign v230170e = hmaster0_p & v23fc3aa | !hmaster0_p & v22f7fdd;
assign v23fb777 = hmaster0_p & v22f81ba | !hmaster0_p & !v22f6d19;
assign v23fbe27 = hmaster2_p & v2311a1d | !hmaster2_p & v84562b;
assign v230156d = hbusreq5_p & v8f2065 | !hbusreq5_p & v22f7dc7;
assign v22f958d = hgrant1_p & v230d56c | !hgrant1_p & v2308813;
assign v22fbb99 = hmaster0_p & v23fae84 | !hmaster0_p & v1aaddf4;
assign v2306473 = hmaster1_p & v23fa823 | !hmaster1_p & v84561b;
assign v23fb5b4 = hbusreq5_p & v84562b | !hbusreq5_p & v12cd4c6;
assign v230ca0f = hbusreq5_p & v191a86f | !hbusreq5_p & !v191a876;
assign v22ff483 = jx1_p & v23fc446 | !jx1_p & v23091d2;
assign v23fceb2 = hmaster2_p & v22f91c9 | !hmaster2_p & !v22f163a;
assign v23fcf4b = hmaster1_p & v2305797 | !hmaster1_p & v84561b;
assign v2310852 = hmaster0_p & v22f4ef0 | !hmaster0_p & v2300686;
assign v1e84038 = hmaster2_p & v23fc46b | !hmaster2_p & !v84561b;
assign v23f35a8 = hbusreq3_p & v22f878c | !hbusreq3_p & v22f511c;
assign v23f6d50 = hbusreq3_p & v22fc8e5 | !hbusreq3_p & v22f878c;
assign v22f5353 = hmaster2_p & v9526ac | !hmaster2_p & v2302149;
assign v230067a = hmaster2_p & v2313131 | !hmaster2_p & v2304d64;
assign v86d5f2 = hmaster0_p & v84561b | !hmaster0_p & !v23930d8;
assign v2308627 = hmaster2_p & b09503 | !hmaster2_p & b00ad2;
assign v23f2d28 = hgrant1_p & v84561b | !hgrant1_p & v2306597;
assign v23fccdb = hbusreq3_p & v23fd05d | !hbusreq3_p & v23fa2ec;
assign v23f40da = hbusreq3 & v230dc73 | !hbusreq3 & v2301319;
assign v230d854 = hmaster2_p & v23f8490 | !hmaster2_p & !v22f0593;
assign v8912cf = busreq_p & v22f8f91 | !busreq_p & v2308a4c;
assign v23fc32a = hmaster0_p & v23fc522 | !hmaster0_p & v22fb757;
assign v23fca34 = hbusreq6_p & v23086d9 | !hbusreq6_p & v23f60ba;
assign v2300ccc = hbusreq3 & v23fbae6 | !hbusreq3 & v845627;
assign v23fc5a9 = hbusreq5_p & v23fc2cc | !hbusreq5_p & v84561b;
assign v2307abc = hmaster0_p & v84561b | !hmaster0_p & v2308ecc;
assign v22f8c8b = hgrant4_p & v23f5201 | !hgrant4_p & v22faa42;
assign v22f2009 = hbusreq4 & v23f26fc | !hbusreq4 & v22ef39f;
assign v23fcfad = hlock3_p & v22fc893 | !hlock3_p & v845620;
assign v23fcf83 = hbusreq5_p & v2308e2e | !hbusreq5_p & v845620;
assign v23f8607 = hmaster2_p & v2306220 | !hmaster2_p & !v23027e9;
assign f405c6 = hbusreq3_p & v23028fc | !hbusreq3_p & da30fb;
assign v22f8d11 = stateG10_5_p & v22ee195 | !stateG10_5_p & v22fd767;
assign v230c12c = hbusreq4_p & v23fb92a | !hbusreq4_p & v84561b;
assign v230713e = hmaster0_p & v2311504 | !hmaster0_p & v1e845a7;
assign v22ed598 = hbusreq3 & v22f2a2f | !hbusreq3 & v1aad988;
assign v23fc6e0 = jx1_p & v23f05c0 | !jx1_p & v23f645e;
assign v22fee78 = hmaster2_p & a1f77b | !hmaster2_p & !v239383d;
assign v22fc6d7 = hlock0_p & v23084ce | !hlock0_p & v23fc18a;
assign v22f231d = hmaster2_p & v23f8da8 | !hmaster2_p & v845620;
assign v230b0f6 = hbusreq3_p & v23fc810 | !hbusreq3_p & v230282c;
assign v22f5c1b = hmaster2_p & v23fcf46 | !hmaster2_p & v23126ae;
assign v23fba43 = hbusreq6 & v22ed400 | !hbusreq6 & v23f9492;
assign v1aae8d3 = hbusreq4_p & v23022d5 | !hbusreq4_p & !v23069b0;
assign v2301c02 = hlock3_p & v84561b | !hlock3_p & v23fd025;
assign v23fc3a1 = stateG10_5_p & v230e8d0 | !stateG10_5_p & !v23f5c95;
assign v22fcdf6 = locked_p & v84561b | !locked_p & v8d360e;
assign v22ebe78 = hbusreq5_p & v23fcf46 | !hbusreq5_p & v23fb55a;
assign v230f554 = hbusreq5_p & v23fc315 | !hbusreq5_p & v22f9f44;
assign v23005e2 = hgrant0_p & v23fb97f | !hgrant0_p & v23fab8b;
assign v22f8839 = hmaster2_p & v84564d | !hmaster2_p & v2301e25;
assign v23fbf2a = stateG10_5_p & v84561b | !stateG10_5_p & v23fc5f4;
assign v23fb88f = hgrant4_p & v84561b | !hgrant4_p & !v22fbf19;
assign v230695e = hbusreq6_p & v22ec414 | !hbusreq6_p & v23f8866;
assign v2305a52 = hbusreq6_p & v22f8a0c | !hbusreq6_p & v22f5c1a;
assign v22f1796 = hgrant1_p & v22f3643 | !hgrant1_p & v2305ebc;
assign v2301511 = hbusreq2_p & v23fba1c | !hbusreq2_p & v84561b;
assign v230ea6d = hbusreq5 & v191a86f | !hbusreq5 & v84561b;
assign v22ed035 = hgrant1_p & v230fec6 | !hgrant1_p & v22f7100;
assign v23fb877 = hmaster0_p & v9ad48f | !hmaster0_p & v22f160c;
assign v23084ce = hbusreq0 & fc8e3a | !hbusreq0 & !v84561b;
assign v13afad9 = hlock5_p & b5f51c | !hlock5_p & !v106ae19;
assign v23fbfe4 = hbusreq5_p & v23fc660 | !hbusreq5_p & v845620;
assign v22ec0de = hbusreq3 & v23fca1c | !hbusreq3 & v84561b;
assign v22f8fa4 = hbusreq1 & v2303dcb | !hbusreq1 & v84561b;
assign v22ff1b0 = hbusreq1 & v22ff090 | !hbusreq1 & v84561b;
assign v23f2849 = hbusreq6_p & v23f8dba | !hbusreq6_p & v22fb7e2;
assign v2309eab = hbusreq3 & v22fd0f1 | !hbusreq3 & v845636;
assign v23fccb7 = hgrant3_p & v23fc975 | !hgrant3_p & v23fb5ba;
assign v23fbbb2 = hburst0_p & v23fc683 | !hburst0_p & !v22f3e8d;
assign v23fcb3f = hgrant3_p & v84561b | !hgrant3_p & v230fd50;
assign v2310075 = hgrant1_p & v84561b | !hgrant1_p & v23fcfbf;
assign v22fda61 = hmaster2_p & v22f6a6e | !hmaster2_p & v22f1895;
assign v22ff12b = hbusreq3 & v23f522c | !hbusreq3 & v84561b;
assign v23fc351 = hgrant3_p & v22ee09d | !hgrant3_p & v23fbadb;
assign bdf576 = hmaster2_p & v23fc89a | !hmaster2_p & !v22f98e3;
assign v230e514 = hbusreq1_p & v22f75d4 | !hbusreq1_p & v230464b;
assign v106a7bd = hgrant0_p & v84561b | !hgrant0_p & !v2306a6f;
assign v23f9452 = hbusreq3_p & v230d134 | !hbusreq3_p & v22efc21;
assign v22f6f0c = hmaster0_p & v23fad13 | !hmaster0_p & !v22ed12b;
assign v23fcced = hgrant1_p & v9526ac | !hgrant1_p & v22f0d2b;
assign v23fc658 = hbusreq5_p & v2303e60 | !hbusreq5_p & !v84561b;
assign v23fc8e4 = hmaster2_p & v106ae19 | !hmaster2_p & v12cd3f4;
assign v22f15e8 = hbusreq4 & c043dc | !hbusreq4 & !v845636;
assign v23f6bba = hgrant3_p & v23f6fa8 | !hgrant3_p & v23fb07c;
assign v23f9546 = hbusreq1 & v22fb0b7 | !hbusreq1 & v22f5583;
assign v23fb7d7 = hgrant3_p & v22ffad4 | !hgrant3_p & v22ef109;
assign v22f7b8b = hgrant1_p & v23fb820 | !hgrant1_p & !v2306b05;
assign v23117c5 = jx1_p & v84561b | !jx1_p & v22f82ea;
assign v239383d = hbusreq1_p & v23fbbf2 | !hbusreq1_p & v23f5a2e;
assign v23f4d1c = hbusreq5 & v22fcdf6 | !hbusreq5 & v84564d;
assign v23fca9e = hbusreq1_p & v2306b2e | !hbusreq1_p & !v23fbbf2;
assign v22ed1e8 = stateG10_5_p & v23fb8fc | !stateG10_5_p & v23f11a3;
assign v23f5f94 = hbusreq3_p & v22fc8d0 | !hbusreq3_p & v23017c7;
assign a1fcc9 = hgrant5_p & v22f8ccb | !hgrant5_p & v2393327;
assign v2306d47 = hbusreq3_p & v22fec56 | !hbusreq3_p & v230a6ed;
assign v23f1227 = hbusreq2_p & v22f4008 | !hbusreq2_p & v23fbaef;
assign v22f2703 = hbusreq5 & v23fc89a | !hbusreq5 & !v845622;
assign v230d65b = hmaster1_p & v84561b | !hmaster1_p & v23fa893;
assign v22f0546 = hbusreq3_p & v22f2c8b | !hbusreq3_p & v22efc04;
assign v22f9833 = hlock3_p & v22fd8a4 | !hlock3_p & !v84561b;
assign v230f974 = hmastlock_p & v22f0c5d | !hmastlock_p & v84561b;
assign v23fc21a = hgrant5_p & v230192f | !hgrant5_p & v22fea89;
assign v23041ab = hgrant3_p & v22f2db6 | !hgrant3_p & !v23f67fe;
assign v23f98ab = hbusreq1_p & a1fbc2 | !hbusreq1_p & v22eb377;
assign v22f6315 = hbusreq6 & v2300b80 | !hbusreq6 & !v23fb7d7;
assign v23fa1f9 = hmaster2_p & v1e84174 | !hmaster2_p & v84561b;
assign v22fbdcf = hbusreq6_p & v23fa95c | !hbusreq6_p & !v1b87732;
assign v23fce7e = hmaster2_p & v22fe5b1 | !hmaster2_p & v23fc98e;
assign v22eb60c = hmaster2_p & v22f5e91 | !hmaster2_p & v22ff1dd;
assign v22f94ec = hbusreq1_p & v22f1d8b | !hbusreq1_p & v84561b;
assign v191accc = hgrant2_p & v84562a | !hgrant2_p & !v230cff9;
assign v23fc847 = hbusreq5_p & v230320e | !hbusreq5_p & !v22ff404;
assign v23fba3d = hbusreq5_p & v23fc4a1 | !hbusreq5_p & v230573f;
assign v2308ee1 = stateG2_p & v2302ca3 | !stateG2_p & v2305e86;
assign v22eba40 = hmaster0_p & v22f56a5 | !hmaster0_p & v2312e4e;
assign v23fb592 = hgrant3_p & v230259f | !hgrant3_p & v22f1899;
assign v1aae277 = hmaster0_p & v2306fba | !hmaster0_p & v230749a;
assign v23f5aa7 = hgrant3_p & v23013a6 | !hgrant3_p & v22f3411;
assign v22f4bf4 = hbusreq5_p & v845636 | !hbusreq5_p & v23fd022;
assign v23096f8 = hbusreq6 & v22f16ef | !hbusreq6 & v230038a;
assign v23f4517 = hgrant2_p & v231241e | !hgrant2_p & v22f3b94;
assign v23f9fdc = hmaster2_p & v22fa7f7 | !hmaster2_p & v23f1e9c;
assign v23fc9d2 = hgrant0_p & v23133fa | !hgrant0_p & a476c2;
assign v23fc660 = hbusreq5 & c258f4 | !hbusreq5 & v845620;
assign v23fc3de = hmastlock_p & v22f8105 | !hmastlock_p & v84561b;
assign v22ffcbd = hlock6_p & v2301274 | !hlock6_p & v845623;
assign v23fbd69 = hbusreq3_p & v23fbb55 | !hbusreq3_p & v84561b;
assign v23040c7 = hlock6_p & v2300e95 | !hlock6_p & v12cd538;
assign v23113f5 = hbusreq4_p & v23f52f2 | !hbusreq4_p & v23fc0d4;
assign bd7b37 = hbusreq0 & v23fcd1b | !hbusreq0 & v84561b;
assign v23fc1d2 = hlock5_p & v230308e | !hlock5_p & !v84561b;
assign v2305e86 = hburst1 & v23fc8a3 | !hburst1 & v23fbc75;
assign v23fcdb0 = hbusreq4 & v23fb9fc | !hbusreq4 & !v23f06d7;
assign v23fca6c = hbusreq4 & v23fb9ca | !hbusreq4 & !v845622;
assign v12cd9e0 = jx1_p & v12cd5e1 | !jx1_p & v23091d2;
assign v23fc32b = stateG2_p & v84561b | !stateG2_p & v2312a9e;
assign v230e352 = hmaster0_p & v239310f | !hmaster0_p & v23fc3af;
assign v23efe71 = hmaster2_p & v23f60ef | !hmaster2_p & !v84561b;
assign v23094a3 = hgrant1_p & v23fb6ff | !hgrant1_p & v230d4c3;
assign v22f3bb0 = hmaster2_p & v84561b | !hmaster2_p & v22f2a4f;
assign v150708b = hmaster2_p & v23f5269 | !hmaster2_p & v23f7f8d;
assign v22ff043 = hbusreq1_p & v23f849c | !hbusreq1_p & v84561b;
assign v22f659a = hbusreq3_p & v22f61f6 | !hbusreq3_p & v23fbf45;
assign v22ed1d3 = hmaster0_p & af7272 | !hmaster0_p & v2308750;
assign v23f77d5 = hmaster2_p & v23f68d8 | !hmaster2_p & v84561b;
assign v22f694d = hbusreq6_p & v22f1b3b | !hbusreq6_p & v84561b;
assign v22fc5d8 = hbusreq3_p & v23fbcd0 | !hbusreq3_p & v2303a74;
assign v2310f5b = hbusreq1 & v23fbddb | !hbusreq1 & v84561b;
assign v22f3396 = hbusreq2_p & v22f1a26 | !hbusreq2_p & !v230f8b2;
assign fc8ab7 = hmastlock_p & v2302c4b | !hmastlock_p & v84561b;
assign v23f5140 = hgrant0_p & v84561b | !hgrant0_p & v23fc8a0;
assign v230d976 = stateG10_5_p & v22eb5cc | !stateG10_5_p & v22fd767;
assign v22fcd0c = hbusreq0_p & v22f1b63 | !hbusreq0_p & v84561b;
assign v22f0542 = stateG10_5_p & v23fcb5e | !stateG10_5_p & v84564d;
assign v23f7429 = hlock3_p & v84561b | !hlock3_p & !v22fc53d;
assign v2303558 = hlock1_p & v23f5cb3 | !hlock1_p & v23fbfb9;
assign v23f6396 = hmaster1_p & v239223a | !hmaster1_p & v23fb53c;
assign v2309783 = hbusreq3 & v23f2f8d | !hbusreq3 & !v845625;
assign v23088a4 = stateG10_5_p & v23fb1c8 | !stateG10_5_p & bdac8d;
assign v22f3b15 = hgrant3_p & v22f31b9 | !hgrant3_p & v23fcfae;
assign v22eef57 = hgrant5_p & v230c124 | !hgrant5_p & v22ef725;
assign v2312401 = hbusreq3_p & v2391d99 | !hbusreq3_p & v22fd150;
assign v22fdc30 = hbusreq2_p & v23126ae | !hbusreq2_p & v106af73;
assign v23fcd7c = hbusreq5_p & v22fd8a6 | !hbusreq5_p & v230b5b8;
assign v23fcab6 = hlock3_p & v23025ae | !hlock3_p & v84562b;
assign v23f3ebd = hbusreq1 & v2312696 | !hbusreq1 & !v23f2c05;
assign v230d5be = hgrant5_p & v23fc782 | !hgrant5_p & !v2300bb2;
assign v23fce9e = hbusreq3 & v23f6e78 | !hbusreq3 & v23f88a9;
assign v22fa771 = hgrant0_p & v84561b | !hgrant0_p & b84615;
assign v230d5aa = hgrant5_p & v230c469 | !hgrant5_p & f40d9e;
assign v22f07bb = hbusreq4_p & v23fcc6c | !hbusreq4_p & v22eafaa;
assign v23030ae = hbusreq3_p & v2393c38 | !hbusreq3_p & v84561b;
assign v22f4e48 = hbusreq4 & v22fcdd3 | !hbusreq4 & !v84561b;
assign v1e84028 = hmaster2_p & v84561b | !hmaster2_p & !v845647;
assign b533b5 = hmaster1_p & v23f2e65 | !hmaster1_p & v84561b;
assign v23f4a0f = jx0_p & v22fa655 | !jx0_p & !v23000a7;
assign v230cb9a = hbusreq1_p & v23fc838 | !hbusreq1_p & v84561b;
assign v23130ac = hlock1_p & v23f486d | !hlock1_p & v22eb06f;
assign v845647 = hmastlock_p & v84561b | !hmastlock_p & !v84561b;
assign v23fb14d = jx1_p & v85e5cf | !jx1_p & !v22efce1;
assign v2305400 = hgrant3_p & v2306c0c | !hgrant3_p & e1e7a3;
assign v23fc975 = hmaster2_p & v22eb377 | !hmaster2_p & v22ff732;
assign v23929d0 = hgrant1_p & f406c6 | !hgrant1_p & !v22ffcb8;
assign v22f7e37 = hgrant5_p & v23fca75 | !hgrant5_p & v239302b;
assign v23fbdec = hmaster2_p & v230de18 | !hmaster2_p & v22fb1bc;
assign v23faf72 = hbusreq4_p & v23fc459 | !hbusreq4_p & v22f9ab6;
assign v22f1874 = hgrant2_p & v230aded | !hgrant2_p & v9526ac;
assign bd7786 = hgrant0_p & v22ebc86 | !hgrant0_p & v22ee247;
assign v2311504 = hbusreq4 & v22f46d3 | !hbusreq4 & v84561b;
assign v23fc6f1 = hlock3_p & v22eecbb | !hlock3_p & !v22ed598;
assign af6dff = hgrant1_p & v22fcc32 | !hgrant1_p & v23fb6c6;
assign v2301c10 = hmaster1_p & v2307b42 | !hmaster1_p & v23fb66e;
assign v23fcf56 = hbusreq4_p & v22fd2e8 | !hbusreq4_p & v9df685;
assign v23fcff5 = hmaster0_p & v23fbb30 | !hmaster0_p & v23063b0;
assign v22f75b0 = hmaster0_p & v22f368e | !hmaster0_p & v22f2d26;
assign v23f6d92 = hbusreq3_p & v22f3092 | !hbusreq3_p & v84561b;
assign e1dcf6 = hbusreq5 & v22f9911 | !hbusreq5 & v230f5a3;
assign v230d8c2 = hbusreq5_p & v22eba12 | !hbusreq5_p & v22f18df;
assign v22f9414 = hbusreq4_p & v23fc1c4 | !hbusreq4_p & !v84561b;
assign v23121ff = hmaster0_p & v191ad8e | !hmaster0_p & v2309897;
assign v2392809 = hbusreq1_p & b2aff2 | !hbusreq1_p & v22f8ad4;
assign v2307b39 = hbusreq5_p & v22ed85a | !hbusreq5_p & v84564d;
assign v22fdfd9 = hmaster2_p & v23f24d1 | !hmaster2_p & v231025b;
assign v22eaf81 = hbusreq4 & v22ed85a | !hbusreq4 & v84561b;
assign v22f7524 = hmaster2_p & v22f954f | !hmaster2_p & v23fb188;
assign v22f0869 = hmaster0_p & v2306703 | !hmaster0_p & c24c97;
assign a15268 = hbusreq4_p & v22ee0ea | !hbusreq4_p & v22f0d28;
assign v2309c9d = hbusreq3_p & v23fad53 | !hbusreq3_p & v230f2ef;
assign v22fa0e4 = hlock3_p & v22eb41e | !hlock3_p & v22f8a7e;
assign v230658d = hgrant1_p & v230e7d4 | !hgrant1_p & v22fd8fc;
assign v9c1abc = hbusreq1_p & v23fc31a | !hbusreq1_p & v23f5526;
assign v22fc8e5 = hlock0_p & v84561b | !hlock0_p & v23fbb35;
assign v23f78a4 = hbusreq5_p & v23f6411 | !hbusreq5_p & !b9d013;
assign v2303a76 = hgrant1_p & a1fc74 | !hgrant1_p & v23f3c1b;
assign e1e1cb = stateG10_5_p & v23f40ba | !stateG10_5_p & v845636;
assign v22f04c8 = hbusreq3_p & v2311e03 | !hbusreq3_p & v22f1697;
assign bf8fe1 = hmastlock_p & v23fb8ee | !hmastlock_p & !v84561b;
assign v23fbe0b = hmaster2_p & v84561b | !hmaster2_p & v2310075;
assign v2310e53 = hmaster1_p & v22eb629 | !hmaster1_p & v22fe1e5;
assign v22ec531 = hbusreq4_p & v22efbaa | !hbusreq4_p & v84561b;
assign v22f4f14 = locked_p & v230fff1 | !locked_p & v84561b;
assign v2301565 = hbusreq4_p & v23fbea7 | !hbusreq4_p & v23fccd7;
assign v23fbffa = hbusreq3_p & v2312ec4 | !hbusreq3_p & v22f73a3;
assign v23051fd = hgrant5_p & v22f5a6c | !hgrant5_p & !v230ba0a;
assign v15071f7 = hbusreq6_p & v23fccf0 | !hbusreq6_p & v23fc76e;
assign v231029e = jx0_p & v23fced3 | !jx0_p & v84561b;
assign v22fd74b = hbusreq1_p & v22f70b0 | !hbusreq1_p & v84561b;
assign v230c025 = hbusreq5_p & v22f7ceb | !hbusreq5_p & v84561b;
assign v23f78c4 = hbusreq4 & v23fbcaa | !hbusreq4 & v22ee657;
assign v22f4bcc = hmaster0_p & v2312eaa | !hmaster0_p & v23fc281;
assign v23fcdf6 = hbusreq3_p & v22f4fb2 | !hbusreq3_p & v23fc3fd;
assign v22f9b95 = hbusreq1_p & v22f8c0b | !hbusreq1_p & bab0c9;
assign v22fa700 = hbusreq1_p & v84562a | !hbusreq1_p & v23067c1;
assign v23fc9b7 = hbusreq4 & v23008a6 | !hbusreq4 & v84561b;
assign v2305933 = hbusreq4_p & v23fc885 | !hbusreq4_p & v22eba40;
assign v22f8f8c = hmaster2_p & b79082 | !hmaster2_p & v84561b;
assign v23f76c2 = hbusreq2_p & v22ee581 | !hbusreq2_p & !v106ae19;
assign v22f2958 = stateA1_p & v84561b | !stateA1_p & !v230cfe2;
assign v22fc712 = hgrant0_p & v84561b | !hgrant0_p & v23fbe61;
assign v22fba3f = hbusreq1 & v23fc7d5 | !hbusreq1 & v22f0add;
assign v2309c14 = hlock0_p & v23fcb76 | !hlock0_p & v2310b6a;
assign v2300362 = hmaster2_p & v106af73 | !hmaster2_p & v230f63f;
assign v23fb9ea = hbusreq5 & v1e84012 | !hbusreq5 & v84561b;
assign v84565f = stateA1_p & v84561b | !stateA1_p & !v84561b;
assign v23f50ec = hlock1_p & v23002e0 | !hlock1_p & v22fe300;
assign v23fce54 = hbusreq3_p & v13afc0b | !hbusreq3_p & !v84561b;
assign v23f8062 = hmaster1_p & v23f5fb9 | !hmaster1_p & !v23f49cd;
assign v22ee495 = hbusreq5_p & a1fba6 | !hbusreq5_p & v22fb891;
assign v23077c2 = hbusreq5_p & v230d346 | !hbusreq5_p & v23f6575;
assign v23006ef = hlock3_p & v22f2e61 | !hlock3_p & !v84561b;
assign v22f99ee = hbusreq5 & v23f8a9d | !hbusreq5 & v84561b;
assign v22f925b = hbusreq2_p & v1aae56f | !hbusreq2_p & v13affaa;
assign v23fa9c5 = hgrant5_p & v22eaa94 | !hgrant5_p & v230bc0c;
assign v2304184 = hbusreq1 & v22fdb01 | !hbusreq1 & v84561b;
assign v2311b1e = hbusreq4_p & v2312846 | !hbusreq4_p & v22f8f64;
assign v23fba7c = hmaster2_p & v23f859a | !hmaster2_p & v23f9226;
assign v22ffe30 = hbusreq6 & v23fb115 | !hbusreq6 & v2306aef;
assign v22f661c = hbusreq1_p & v23fbc48 | !hbusreq1_p & v22ec41b;
assign v2308058 = hgrant5_p & v23fb98c | !hgrant5_p & !v22f6410;
assign v23fcc44 = hmaster0_p & v22ef377 | !hmaster0_p & !v96c563;
assign v23fcf9e = hmaster0_p & v23fb931 | !hmaster0_p & v22fd0fa;
assign v22fadb0 = hbusreq0_p & v230fc70 | !hbusreq0_p & v23fc2ee;
assign v2307d93 = hbusreq4 & v23fb145 | !hbusreq4 & v22f5fb4;
assign v22f4301 = hmaster2_p & v23f53bd | !hmaster2_p & v23933e8;
assign v230eafa = hbusreq3 & v23f15ac | !hbusreq3 & v84561b;
assign v2313463 = locked_p & v845661 | !locked_p & !v84561b;
assign v2305263 = hmaster0_p & v22f6066 | !hmaster0_p & v230d836;
assign v239160b = hgrant3_p & v23f581f | !hgrant3_p & v23f1ccc;
assign v22ff732 = hlock0_p & a1fbc2 | !hlock0_p & v22f8fe0;
assign v23f7b94 = hbusreq4_p & v2303e0d | !hbusreq4_p & v23fc013;
assign v2305d50 = hbusreq4 & v2304f11 | !hbusreq4 & v84561b;
assign v2307020 = hlock3_p & v230eac0 | !hlock3_p & v23fba73;
assign v23fab82 = hbusreq0 & v23fcb0b | !hbusreq0 & v84562a;
assign v22fb790 = hbusreq4_p & v23916ef | !hbusreq4_p & v84561b;
assign v23fb842 = jx2_p & v23f443d | !jx2_p & v230fe41;
assign v2311c98 = hbusreq3 & v23f53bd | !hbusreq3 & v23fba9a;
assign v10dbf63 = hlock6_p & v84564d | !hlock6_p & !v84561b;
assign v22f8917 = locked_p & v230ff13 | !locked_p & v23fba6b;
assign v23fa77d = hmaster2_p & v23f445f | !hmaster2_p & v230dbc9;
assign v22f0b8a = hmaster2_p & v22f954f | !hmaster2_p & v23934f0;
assign v22f4d28 = hmaster2_p & v2310e40 | !hmaster2_p & v23fccbe;
assign v22eb651 = hgrant3_p & v84561b | !hgrant3_p & v23fb77d;
assign v2310537 = hready_p & v22ebfcf | !hready_p & v22ec5e3;
assign v22f7d00 = hbusreq4_p & v23f7cec | !hbusreq4_p & v22fe84a;
assign v23fb6ed = hmaster2_p & v23f6bc1 | !hmaster2_p & v84561b;
assign v230bba4 = hbusreq3_p & v23fc5eb | !hbusreq3_p & v23f513d;
assign v23f31d6 = hbusreq4 & v23fc52d | !hbusreq4 & v23fa77d;
assign v22f9ef0 = hbusreq0 & v2303a7f | !hbusreq0 & v23f4462;
assign v23fc2d7 = hmaster2_p & v22fa8e6 | !hmaster2_p & b50a75;
assign v230b913 = hbusreq0 & v23fcf9b | !hbusreq0 & v84561b;
assign b9d0d2 = hgrant1_p & v22fd2ec | !hgrant1_p & !v23fb992;
assign v23fc583 = hbusreq5_p & v23fc243 | !hbusreq5_p & v84561b;
assign v23fc06c = hgrant1_p & v22edf62 | !hgrant1_p & !v230e598;
assign v231007b = hgrant1_p & v23fc904 | !hgrant1_p & v23f2a7c;
assign v23f2698 = hgrant3_p & v22fe9dc | !hgrant3_p & v23f73dd;
assign v2306298 = hbusreq5_p & v23f1a8d | !hbusreq5_p & v22f5ca6;
assign v2304d59 = hmaster0_p & v84561b | !hmaster0_p & v23fce31;
assign v22fe740 = hlock5_p & v2304a1e | !hlock5_p & !v84561b;
assign v23fc840 = hmaster0_p & v22f3e2e | !hmaster0_p & v23055c3;
assign v22f51b1 = hbusreq4_p & v23fce89 | !hbusreq4_p & v22f482d;
assign v22fb5b1 = hbusreq2_p & v22fd781 | !hbusreq2_p & !v22f39b0;
assign v23fbca4 = hbusreq5 & v22f60c6 | !hbusreq5 & v84561b;
assign v2310051 = hmaster2_p & v84561b | !hmaster2_p & v23fc4e8;
assign v22ef38d = hmaster1_p & v23fb7c8 | !hmaster1_p & !v23041ea;
assign v22f9734 = hbusreq4_p & v22f04bf | !hbusreq4_p & v84561b;
assign v2312c62 = hgrant3_p & v2305cac | !hgrant3_p & v22eeef8;
assign v23fb63e = hmaster0_p & v22f31b9 | !hmaster0_p & !v2303b1a;
assign v22ee4e7 = hlock4_p & v2307c15 | !hlock4_p & v23fcc7c;
assign v23fb993 = hbusreq5_p & v23fc3cb | !hbusreq5_p & v22f8d11;
assign v22f0051 = hbusreq5 & v22fa707 | !hbusreq5 & v84561b;
assign v22f87a1 = hbusreq6 & v23fb9ca | !hbusreq6 & !v845622;
assign v23fc98b = hmaster0_p & v23fc790 | !hmaster0_p & v23f89fc;
assign v2302bb2 = stateG10_5_p & v23f94e5 | !stateG10_5_p & v845636;
assign v23fb99f = hlock4_p & v230aa0c | !hlock4_p & v23fb821;
assign v23fc382 = hbusreq5 & v22f3c3d | !hbusreq5 & !v84561b;
assign v23fbc1b = hmaster0_p & v22f56a5 | !hmaster0_p & v23f1225;
assign v23f5ead = hlock1_p & v230bafe | !hlock1_p & v22ff1b0;
assign v23fc8ee = hbusreq0 & v13afe3a | !hbusreq0 & !fc8e3a;
assign v22f84a0 = hbusreq6 & v230d99c | !hbusreq6 & v23016d9;
assign v22eab03 = jx1_p & v231246b | !jx1_p & v23f8062;
assign v23fb218 = hbusreq5 & fc8e3a | !hbusreq5 & !v84561b;
assign v9bcad3 = hbusreq3 & v22fe285 | !hbusreq3 & v22fe2ae;
assign v22f6c46 = hmaster1_p & v231321e | !hmaster1_p & v23fb4a5;
assign v23fbf6c = hbusreq1_p & v22fc091 | !hbusreq1_p & v22f65d5;
assign v23fc0de = hbusreq5_p & v22eeb07 | !hbusreq5_p & v84561b;
assign v23fc364 = hlock4_p & v22f0f76 | !hlock4_p & v2308669;
assign v23fcc9a = hgrant1_p & v22f05a0 | !hgrant1_p & v22f6de3;
assign v23fbbbf = hbusreq4 & v22f9f88 | !hbusreq4 & v22eeece;
assign a6db07 = hgrant3_p & v84562e | !hgrant3_p & v22ef998;
assign v22f3730 = hbusreq6_p & v23fc4b7 | !hbusreq6_p & v22f79a5;
assign v23fbcd0 = hmaster2_p & v22f2998 | !hmaster2_p & v23fcced;
assign v22fbef0 = hbusreq3 & v23101b0 | !hbusreq3 & v84561b;
assign v2308c0b = hbusreq5_p & v23fc1fb | !hbusreq5_p & v2309963;
assign v2312d2c = jx3_p & v22f4339 | !jx3_p & v22f7f12;
assign v15071f0 = hbusreq5 & v23fc35a | !hbusreq5 & v2302d97;
assign v22ed4b7 = hbusreq3 & v230a65d | !hbusreq3 & v22ef062;
assign v23fc92f = hmaster2_p & v191a86f | !hmaster2_p & v22eb1f5;
assign v23fc2dd = hmastlock_p & v22f334e | !hmastlock_p & !v84565f;
assign v1aae2a8 = hbusreq5_p & v23062f0 | !hbusreq5_p & v84561b;
assign v230e2bd = jx1_p & v23f11ae | !jx1_p & v84561b;
assign v23f6e45 = hlock1_p & v23f8772 | !hlock1_p & v84562b;
assign v23fccc6 = hbusreq4_p & v22fca12 | !hbusreq4_p & v84561b;
assign v23fba16 = hbusreq6 & v22ebebe | !hbusreq6 & v84561b;
assign v22ec2e6 = hbusreq4 & v23fc72d | !hbusreq4 & v84561b;
assign v23f809b = hbusreq5_p & v84561b | !hbusreq5_p & v22fd3b1;
assign v23f087f = hbusreq5_p & v8f2065 | !hbusreq5_p & v23f1a43;
assign v23fb91d = hmaster2_p & v845627 | !hmaster2_p & v23fc511;
assign v23fbcb1 = hmaster2_p & v23fba6b | !hmaster2_p & !v230882d;
assign afffd9 = hmaster2_p & v23f5af5 | !hmaster2_p & v22ed7a8;
assign v230c995 = hgrant3_p & v23fb937 | !hgrant3_p & v230fae1;
assign v23fbf9b = hmaster1_p & v23fc754 | !hmaster1_p & v2302d12;
assign v23007a2 = hgrant2_p & v230c0e9 | !hgrant2_p & v13affaa;
assign v22f65b7 = hbusreq1_p & v23fb1ab | !hbusreq1_p & v84562b;
assign v22eb3fc = hmaster2_p & v22f1ae7 | !hmaster2_p & v23fc4a3;
assign v23fb6a6 = hbusreq1 & v1aadb8e | !hbusreq1 & v84561b;
assign v23f2380 = hmaster0_p & v22fcc78 | !hmaster0_p & v230afed;
assign v22eaf66 = hmaster0_p & v23f3f24 | !hmaster0_p & v22fde5c;
assign v23fc27d = hbusreq3_p & v23fcc91 | !hbusreq3_p & v22fc8c8;
assign v22ff613 = hbusreq5 & v23fcb5b | !hbusreq5 & v191aa95;
assign ae78a6 = hmaster2_p & v23faa16 | !hmaster2_p & v23fc04c;
assign v22fd02d = hgrant4_p & v84561b | !hgrant4_p & v2309410;
assign v23114a6 = locked_p & v22fd9be | !locked_p & !v84561b;
assign v23f0135 = hlock0_p & v230f4a8 | !hlock0_p & v22ee9be;
assign v22f0d5a = hbusreq3_p & v845622 | !hbusreq3_p & v22edff5;
assign v22f7004 = hgrant0_p & v23fc4f8 | !hgrant0_p & v2301b2d;
assign v230eafe = hbusreq1_p & v23fc047 | !hbusreq1_p & v22f1ae5;
assign e1df2d = locked_p & v23fca94 | !locked_p & v84561b;
assign v23fb073 = hmaster2_p & v23fccb2 | !hmaster2_p & v15070ca;
assign v23fbef9 = hbusreq1 & v2305ebc | !hbusreq1 & v84561b;
assign v23fc622 = hbusreq0_p & v23f5043 | !hbusreq0_p & v84564d;
assign v2392836 = hbusreq1_p & v22f4bb5 | !hbusreq1_p & v845620;
assign v230290f = hlock3_p & v22ee9bb | !hlock3_p & v23fce88;
assign v2301fe9 = hgrant5_p & v23f66a4 | !hgrant5_p & v23f36a5;
assign v1506a4c = hmaster2_p & v22f91c9 | !hmaster2_p & !v2392974;
assign v23fc9a4 = hgrant3_p & v84561b | !hgrant3_p & !v845651;
assign v230dfff = hmaster2_p & v23fc63b | !hmaster2_p & v1aae490;
assign v2393091 = hmaster0_p & v2305d50 | !hmaster0_p & v22fb44a;
assign v22f3b2e = hmaster0_p & a2e978 | !hmaster0_p & !v96c563;
assign v230b4d9 = hgrant5_p & v23080ab | !hgrant5_p & v230e191;
assign v22f1a0e = hmaster1_p & v22eb134 | !hmaster1_p & v84561b;
assign v22eb67a = hbusreq1_p & v22f3ad4 | !hbusreq1_p & v2313463;
assign v2302943 = hbusreq4_p & v22fa23d | !hbusreq4_p & bd8af4;
assign v22fa870 = hbusreq5_p & v2302e32 | !hbusreq5_p & v22eb1f5;
assign v2305252 = hmaster2_p & v2300c3d | !hmaster2_p & v84564d;
assign v2308ef0 = hbusreq6 & v22f961e | !hbusreq6 & v22f2ca2;
assign v23f51cc = hbusreq6_p & v22f2852 | !hbusreq6_p & v22f88bb;
assign a1fdb9 = hbusreq3_p & v23fb91d | !hbusreq3_p & v22f3aac;
assign v22f5e60 = hmastlock_p & v230c4a4 | !hmastlock_p & !v84561b;
assign v2302553 = jx3_p & v84561b | !jx3_p & v23fc73b;
assign v22f8fb2 = hburst1_p & v845649 | !hburst1_p & v84561b;
assign v22f2b34 = hmaster1_p & v22fd841 | !hmaster1_p & v23fc46c;
assign v2302048 = hbusreq2_p & v84561b | !hbusreq2_p & v22f1389;
assign v22ec1ef = hgrant3_p & v2301b00 | !hgrant3_p & v22f3add;
assign v23fc8a6 = hbusreq3_p & v2300d93 | !hbusreq3_p & v2308d80;
assign v230183d = hgrant4_p & v23934ed | !hgrant4_p & v23fceb5;
assign v9f4f45 = hlock2_p & v23f391e | !hlock2_p & v23fc739;
assign v23f38ff = hbusreq5_p & v23f847c | !hbusreq5_p & v22f2d51;
assign v2310589 = hlock4_p & v22fc8e5 | !hlock4_p & v2309c93;
assign v23f38b7 = hbusreq3_p & v22f243b | !hbusreq3_p & v22f5c1b;
assign v23f3958 = hlock6_p & v23fb813 | !hlock6_p & v2300b7b;
assign v1506ff4 = hmaster2_p & v84561b | !hmaster2_p & v22ed85a;
assign v23f89df = hgrant5_p & v22f9690 | !hgrant5_p & v12cc72f;
assign v23088ef = hbusreq3_p & v22ff0da | !hbusreq3_p & v1506a4c;
assign v23f17ff = hmaster1_p & v22edb96 | !hmaster1_p & v22f04b5;
assign v230e547 = hlock2_p & v22ff090 | !hlock2_p & v230abfb;
assign fc8f5a = hbusreq6_p & v22f216d | !hbusreq6_p & v23f427e;
assign v23f9bd1 = hbusreq6_p & v23f2353 | !hbusreq6_p & v231248c;
assign v230e54d = hmaster2_p & v22f5037 | !hmaster2_p & !v22fbeea;
assign v22ebddc = hgrant3_p & v84561b | !hgrant3_p & v23f552d;
assign v22ecc0d = stateG10_5_p & v22f217d | !stateG10_5_p & !v84561b;
assign v23102bf = hlock1_p & v1506f02 | !hlock1_p & v23f4e25;
assign v22f0a7b = jx3_p & v230eb8e | !jx3_p & v22f89c7;
assign v22ee4b6 = locked_p & v845661 | !locked_p & v106a782;
assign v23f4861 = hbusreq3_p & v2300d67 | !hbusreq3_p & v23f5ef2;
assign v230e322 = hbusreq3 & v22f99e0 | !hbusreq3 & v84561b;
assign v2310c7c = hbusreq2_p & v2309377 | !hbusreq2_p & !v23046f7;
assign v23f7a18 = hmaster2_p & v23fcf89 | !hmaster2_p & v230db4e;
assign v22f63e9 = hmaster0_p & v23fc0a3 | !hmaster0_p & v23f1495;
assign v23fc116 = start_p & v84561b | !start_p & !v22f476c;
assign v23f6ac2 = hmastlock_p & v230db9d | !hmastlock_p & v84561b;
assign v895ae7 = hgrant1_p & v23fb6ff | !hgrant1_p & v9347cd;
assign v2302f72 = hlock3_p & v23fb231 | !hlock3_p & v23fba62;
assign v23fcaec = hmaster0_p & v230502a | !hmaster0_p & v230a7c3;
assign v23fbf94 = hbusreq4 & v23fc56a | !hbusreq4 & v22f0331;
assign v23fb8e0 = hmaster2_p & v230358b | !hmaster2_p & v23fc48b;
assign v23fbd62 = hmaster0_p & v23f5868 | !hmaster0_p & v23fbcac;
assign v23fbcc8 = hbusreq3_p & v22f2bab | !hbusreq3_p & v23f2d31;
assign v23fc0ac = hmaster2_p & v2302a4d | !hmaster2_p & !v22f9980;
assign v230801c = hbusreq3_p & v22f1fca | !hbusreq3_p & v84561b;
assign v2312ebe = hlock4_p & v2393401 | !hlock4_p & v22eef1f;
assign v230ec4a = hbusreq3_p & v1aad988 | !hbusreq3_p & v230554d;
assign v2303e60 = hlock5_p & v22ff89d | !hlock5_p & !v84561b;
assign v23f37b9 = hmaster0_p & v23f439b | !hmaster0_p & v1aadcf6;
assign v23fbfd5 = hmaster2_p & v23fbc3f | !hmaster2_p & v22eb377;
assign v22fcfed = hbusreq3 & v23fbfc3 | !hbusreq3 & v23fc439;
assign v12cdab5 = hmaster2_p & v22f902d | !hmaster2_p & v22f7b29;
assign v22fd32a = hbusreq4_p & v22f6228 | !hbusreq4_p & v22f51ba;
assign v23068a9 = locked_p & v84565f | !locked_p & !v84561b;
assign v23f0bf1 = hgrant1_p & a07f9b | !hgrant1_p & v2392d4f;
assign v22f5c4c = hmaster0_p & v22fb10b | !hmaster0_p & !v23f8988;
assign v23f3206 = hgrant1_p & v2303d00 | !hgrant1_p & v22f214f;
assign v23fb724 = hmaster0_p & v23f2fb7 | !hmaster0_p & v84562d;
assign v230a434 = stateG3_0_p & v845665 | !stateG3_0_p & v84561b;
assign v22f5a27 = hbusreq4_p & v8bc4e1 | !hbusreq4_p & v22ec644;
assign v22ec87b = stateG2_p & v84561b | !stateG2_p & v23f54be;
assign v22f1133 = hlock0_p & v23efdd0 | !hlock0_p & v230818b;
assign v23f3d39 = hbusreq0_p & v23fc14e | !hbusreq0_p & !v22f6518;
assign v23fb964 = hbusreq4 & a20348 | !hbusreq4 & v22f8551;
assign v22f7ceb = hlock5_p & v84561b | !hlock5_p & !v23fb4ae;
assign v23f59e0 = hlock2_p & v22f8d74 | !hlock2_p & v845620;
assign v23f608b = hmaster0_p & v2302907 | !hmaster0_p & !v231089e;
assign v22fc091 = hbusreq0_p & v22ff38e | !hbusreq0_p & v84561b;
assign v23fc802 = hgrant3_p & v23fcd84 | !hgrant3_p & v23fc821;
assign v22ff90b = hgrant1_p & v84561b | !hgrant1_p & v22f74de;
assign v22fa6ae = hbusreq6_p & v22f6f2d | !hbusreq6_p & v191acb4;
assign v22fc723 = hgrant5_p & v84561b | !hgrant5_p & !v23fc51f;
assign v22f95a4 = hmaster0_p & v23fbcf8 | !hmaster0_p & v230b837;
assign v22f58c2 = hbusreq4 & v22fb554 | !hbusreq4 & v22f5583;
assign v23f9870 = hmaster2_p & v22f62ae | !hmaster2_p & v22f61b6;
assign v22ed48e = hmaster0_p & v2310782 | !hmaster0_p & v23928d0;
assign v23fcd4b = hbusreq3 & v230f370 | !hbusreq3 & v23070cf;
assign v230f087 = hgrant3_p & fc8fe6 | !hgrant3_p & v230da69;
assign v23fc7dd = hbusreq2_p & v22fe9b7 | !hbusreq2_p & v22f8917;
assign v23fb504 = hmaster2_p & v23f5043 | !hmaster2_p & v23fbb80;
assign v2308c4d = hgrant6_p & v191ac63 | !hgrant6_p & v1506fdd;
assign v23fc5ab = hmaster2_p & v23fbaaa | !hmaster2_p & v23fbddf;
assign v23f7fe8 = hmaster0_p & v22f6dee | !hmaster0_p & v22f1ab6;
assign v13afb18 = hbusreq5_p & v23fb0c2 | !hbusreq5_p & v84561b;
assign v23fbe1f = jx3_p & v85d975 | !jx3_p & !v84561b;
assign v23fa8d7 = hgrant5_p & v22eefc4 | !hgrant5_p & v22f533e;
assign v230e437 = jx1_p & v230efa2 | !jx1_p & v22ec6a7;
assign v2310037 = hbusreq6_p & v23fc0b9 | !hbusreq6_p & v12cd4da;
assign v2301216 = hmaster2_p & v22f94ec | !hmaster2_p & v23f9f77;
assign v23fbb0e = hgrant3_p & v845625 | !hgrant3_p & v17cf1d8;
assign v2309464 = hmaster2_p & v23fb6e3 | !hmaster2_p & !v22feb6e;
assign v23fcadf = hbusreq1 & v13afe8f | !hbusreq1 & v84561b;
assign v23fcafd = hbusreq3_p & v230067a | !hbusreq3_p & v2309130;
assign v22f8f5f = hmaster0_p & b00aa6 | !hmaster0_p & v23f446c;
assign v23f939f = hlock1_p & v230f70d | !hlock1_p & !v84561b;
assign v23fbb10 = hgrant2_p & v23fcf25 | !hgrant2_p & v22efdb1;
assign v22ff179 = hmaster2_p & v84564d | !hmaster2_p & !v23fb1a4;
assign v2312a18 = hbusreq6 & v23f8561 | !hbusreq6 & v84561b;
assign v2305f58 = hbusreq0_p & v23f51b1 | !hbusreq0_p & !v106ae19;
assign v22ffacb = hbusreq5_p & v23037b2 | !hbusreq5_p & !v84561b;
assign v230abc9 = hbusreq4_p & v2391fc6 | !hbusreq4_p & v23f397b;
assign v22ff9c5 = hbusreq3 & v845620 | !hbusreq3 & v23f7ce8;
assign v2308ae7 = hbusreq1 & v2306538 | !hbusreq1 & v22f8c0b;
assign v230ca62 = hmaster0_p & v23f3f24 | !hmaster0_p & !v22f324a;
assign v22efb8c = hbusreq6 & v22ee946 | !hbusreq6 & v23fc493;
assign v23faacb = hmaster2_p & a07f9b | !hmaster2_p & v22eb377;
assign v23fcba2 = hmaster0_p & v230b131 | !hmaster0_p & v23fb592;
assign v230cd87 = hmaster2_p & v1506ad8 | !hmaster2_p & v23fc094;
assign v23fc607 = hmaster2_p & v22f65d5 | !hmaster2_p & v22fc5f0;
assign v22fe985 = hbusreq4_p & v86a21a | !hbusreq4_p & v23fb0ab;
assign v22f53a0 = jx3_p & v23fcba6 | !jx3_p & !v230648e;
assign v2309033 = hgrant1_p & v22f4aa2 | !hgrant1_p & v22fc979;
assign v22eb0b3 = hmaster0_p & v84561b | !hmaster0_p & v22fed5c;
assign v23fa9d0 = hlock1_p & v22fe59c | !hlock1_p & !v84561b;
assign v2312f44 = hmaster2_p & v23fcc81 | !hmaster2_p & v22f742b;
assign v230571c = hbusreq1_p & v22f866f | !hbusreq1_p & !v23fccec;
assign v23fc84a = hmaster2_p & v23fa4bd | !hmaster2_p & v2303bc3;
assign v22ef2be = hbusreq3 & v23fb236 | !hbusreq3 & v2310238;
assign v22efa95 = hbusreq4_p & ad78c9 | !hbusreq4_p & v2302dca;
assign v23fc019 = hmaster2_p & v22fe497 | !hmaster2_p & v979b7c;
assign v1aaddcb = hlock6_p & v84561b | !hlock6_p & !v23fbb00;
assign bd9ab5 = hgrant1_p & v90af77 | !hgrant1_p & v9c12cb;
assign v23fce8b = stateG10_5_p & v23efed1 | !stateG10_5_p & !v23f96f7;
assign v23fcddd = hbusreq4_p & v933ab1 | !hbusreq4_p & v23fb7ea;
assign v22f68e5 = hmaster2_p & v2302a4d | !hmaster2_p & !v191a879;
assign v230be24 = hlock0_p & v22f15fe | !hlock0_p & v23fbd16;
assign ba1576 = hmaster2_p & v23f646e | !hmaster2_p & !v23f5cb3;
assign v23fbf16 = hbusreq6_p & v2305c7f | !hbusreq6_p & v23074d2;
assign v1aad4ef = hgrant3_p & v84561b | !hgrant3_p & v230a891;
assign v23fb2e9 = hmaster2_p & v22f7e4a | !hmaster2_p & v23f3dd3;
assign v23fc849 = stateG10_5_p & v239254b | !stateG10_5_p & v84562b;
assign v23f3a95 = hlock0_p & v230995b | !hlock0_p & v23fc1dc;
assign v22fc2bd = hlock0_p & v84561b | !hlock0_p & v22fe59a;
assign v15075a6 = hlock1_p & v22f3834 | !hlock1_p & fc8ab7;
assign v22f4168 = hbusreq1 & v2304009 | !hbusreq1 & v23fd021;
assign v23fcc09 = hbusreq2 & v22ee0c4 | !hbusreq2 & v845620;
assign v23f45d2 = hbusreq5_p & v85d110 | !hbusreq5_p & v22eefd1;
assign v22f8b43 = hbusreq1_p & v230df7b | !hbusreq1_p & b7427f;
assign v23f1a86 = hbusreq4 & v22ff18a | !hbusreq4 & v845627;
assign v191b038 = hbusreq6_p & v230e8a7 | !hbusreq6_p & v231005a;
assign v23fa511 = hmaster2_p & b9d013 | !hmaster2_p & !v22ffbb3;
assign v23fbbc7 = hbusreq2_p & v2307805 | !hbusreq2_p & !v84561b;
assign v22ffde1 = jx3_p & v22f43c9 | !jx3_p & v22f5033;
assign v23fce39 = jx1_p & v85e5cf | !jx1_p & !bd7535;
assign v22ec63d = hbusreq3_p & v22f8ad5 | !hbusreq3_p & v230859e;
assign v22f08f1 = jx0_p & v23f443c | !jx0_p & v22eec56;
assign v2307b25 = hbusreq6 & v22f60da | !hbusreq6 & !v84561b;
assign v22ff5af = hbusreq1_p & v23f5043 | !hbusreq1_p & v84564d;
assign v23fce77 = hmaster2_p & v23fcb5b | !hmaster2_p & v84561b;
assign v23fc02d = hmaster2_p & v22f6358 | !hmaster2_p & v22f66cf;
assign v23fc050 = hbusreq1 & v22ff414 | !hbusreq1 & v84561b;
assign v230bbf8 = hgrant3_p & v23fbad3 | !hgrant3_p & v22fb1f3;
assign v22f7914 = hgrant3_p & v84562e | !hgrant3_p & v23fc9e5;
assign v12cd6a2 = hlock3_p & v23fc898 | !hlock3_p & !v84561b;
assign v2305d2f = hgrant1_p & v84561b | !hgrant1_p & v23fce72;
assign v23f8324 = hbusreq4_p & v22fd2e8 | !hbusreq4_p & v23f4dc4;
assign v23f95c3 = hgrant3_p & v23006ef | !hgrant3_p & !v84561b;
assign v23f8e1f = stateG2_p & v84561b | !stateG2_p & v23f67dd;
assign v23fd015 = hlock3_p & v84561b | !hlock3_p & v22f5218;
assign b20f9d = hgrant6_p & v23f89f0 | !hgrant6_p & v23fcdbd;
assign v22f6963 = hbusreq4_p & v2391d0b | !hbusreq4_p & v230a775;
assign v22edcfc = hbusreq2 & c086a6 | !hbusreq2 & v84561b;
assign v230282c = hbusreq3 & v23fc864 | !hbusreq3 & !v230d7e4;
assign v23fc2a0 = hbusreq5_p & v84561b | !hbusreq5_p & v230474b;
assign v22f2590 = hbusreq0 & v2304ec7 | !hbusreq0 & !v84561b;
assign v230e7e4 = hmaster2_p & v23124cc | !hmaster2_p & v84561b;
assign v23fba29 = stateG2_p & v84561b | !stateG2_p & v22ef862;
assign v23f7c8d = hmaster2_p & v84561b | !hmaster2_p & v23f8364;
assign v23fb875 = hlock0_p & v9526ac | !hlock0_p & v238ae11;
assign v23fbaf0 = hbusreq5 & v13afe3a | !hbusreq5 & !fc8e3a;
assign v23f41ec = hbusreq4 & v22fea26 | !hbusreq4 & !v845625;
assign fc8fcf = hgrant4_p & v22fdc20 | !hgrant4_p & v22ec960;
assign v23fba03 = hgrant5_p & v22f7a0c | !hgrant5_p & v23fcc22;
assign v23112a4 = hbusreq3 & v23f5207 | !hbusreq3 & v2305507;
assign v2391655 = hmaster0_p & v2301be6 | !hmaster0_p & !v22fab21;
assign v2308b19 = hbusreq1 & v230e4ef | !hbusreq1 & v2391d40;
assign v2303efa = jx1_p & v191abed | !jx1_p & v22efd99;
assign v23fc822 = hbusreq4_p & v23fc97a | !hbusreq4_p & !v84561b;
assign v23fbda8 = hlock6_p & v23f1206 | !hlock6_p & !v106ae19;
assign v230333f = locked_p & v22ef27f | !locked_p & v84561b;
assign v23f34e1 = hbusreq4_p & v230c949 | !hbusreq4_p & v230adbf;
assign v23fce9c = hgrant5_p & v2311506 | !hgrant5_p & v22f1040;
assign v2309e12 = hmaster2_p & v23060d4 | !hmaster2_p & v23fb49a;
assign v23916d6 = hmastlock_p & v2308ee1 | !hmastlock_p & !v84561b;
assign v23fbb37 = hbusreq2_p & v2309515 | !hbusreq2_p & v84564d;
assign v22ed03d = hgrant5_p & v2391982 | !hgrant5_p & v22fa002;
assign v2312fc7 = hgrant0_p & v23f0135 | !hgrant0_p & v22fda30;
assign v23121aa = hmaster0_p & v23f38d5 | !hmaster0_p & !v2302370;
assign v239213c = hbusreq3 & v22f9657 | !hbusreq3 & v84561b;
assign v22f0acd = hgrant1_p & v2309a71 | !hgrant1_p & v2305e51;
assign v22f2ca2 = hlock3_p & v84562d | !hlock3_p & !v84561b;
assign v230c0b4 = hlock3_p & v22eeecc | !hlock3_p & v23f8c92;
assign ab2d7c = hmastlock_p & v22fccc4 | !hmastlock_p & v84561b;
assign v23019e9 = hmaster2_p & v23105cd | !hmaster2_p & v22f3643;
assign v23080ec = hgrant1_p & v23f87f4 | !hgrant1_p & b30f07;
assign v23fcd52 = stateG10_5_p & v23fc066 | !stateG10_5_p & v23f296d;
assign v230a688 = hmaster1_p & v22eec68 | !hmaster1_p & !v23fbc0d;
assign v2305606 = hmaster2_p & b9d049 | !hmaster2_p & !v84561b;
assign v22f5a56 = hbusreq1_p & v2301934 | !hbusreq1_p & v22f7241;
assign v22ed72b = hbusreq3_p & v22fc508 | !hbusreq3_p & v22ed5c8;
assign v2308b6b = stateG10_5_p & v22ff399 | !stateG10_5_p & v2311d9d;
assign c20101 = hmaster2_p & v23fc393 | !hmaster2_p & !v2306d29;
assign v2302022 = hgrant5_p & v84561b | !hgrant5_p & v22fd029;
assign v23fbbb9 = hmaster2_p & v23fba65 | !hmaster2_p & v22f954f;
assign v23f2bfa = hmaster2_p & v22ee9ac | !hmaster2_p & !v23fa345;
assign v22fc85f = hmaster0_p & v23fc5a0 | !hmaster0_p & v22fcdf7;
assign v22f2f33 = hbusreq5 & v23fd050 | !hbusreq5 & v23124cc;
assign v22f90bf = hbusreq5_p & v23f08e5 | !hbusreq5_p & v231206c;
assign v230fc8c = hbusreq5_p & v2306d29 | !hbusreq5_p & v23065ad;
assign v23fbf28 = hmaster0_p & v230ea9f | !hmaster0_p & v23fb699;
assign v23fc43d = hgrant3_p & v84561b | !hgrant3_p & v22fb769;
assign v23f01d5 = hbusreq6 & v2310ec5 | !hbusreq6 & v22f0d5a;
assign v23f80c9 = hbusreq3_p & v23f75e5 | !hbusreq3_p & v2300004;
assign v23fc18a = hbusreq0 & fc8ab7 | !hbusreq0 & !v84561b;
assign v23fc1bf = hbusreq5_p & v23fcbde | !hbusreq5_p & v2310558;
assign v23f552d = hmaster2_p & v22f1244 | !hmaster2_p & v22fc1df;
assign v22fb8d3 = hgrant2_p & v23fa2e7 | !hgrant2_p & !v106ae19;
assign v23fc923 = hbusreq5_p & v2304bd1 | !hbusreq5_p & v84561b;
assign v23f3915 = hmaster2_p & v230bd96 | !hmaster2_p & v23fc484;
assign v22efee2 = hbusreq1 & v106ae21 | !hbusreq1 & v84561b;
assign v23fb60e = hmaster2_p & v2312bd9 | !hmaster2_p & v23f51da;
assign v22ec562 = hbusreq5_p & v22f299f | !hbusreq5_p & v22f5974;
assign v23f8a06 = hbusreq1 & v8d360e | !hbusreq1 & !v84561b;
assign v22f1166 = hgrant3_p & v23fb97a | !hgrant3_p & v23fb0d9;
assign v22f7f2a = hgrant5_p & v22ec98c | !hgrant5_p & v84561b;
assign v2300cc2 = hmaster0_p & v23fbe2d | !hmaster0_p & v22fed78;
assign v22f4bdf = hmastlock_p & v23f2a1a | !hmastlock_p & v84561b;
assign v230b7fc = hbusreq3_p & v22f092f | !hbusreq3_p & v22f62ea;
assign v230aa96 = hmaster2_p & v22f31b2 | !hmaster2_p & v22f893a;
assign v23fbedb = hmaster2_p & v2300934 | !hmaster2_p & !v22fb1bc;
assign v23f7254 = hbusreq3 & v22efd4d | !hbusreq3 & v22f7195;
assign v2303c10 = hmaster2_p & v23fc58e | !hmaster2_p & v1aae09e;
assign f40d66 = hgrant1_p & v845625 | !hgrant1_p & v230d75a;
assign v23fbb95 = hbusreq1 & v23fbfd0 | !hbusreq1 & v23fce71;
assign v23fb8d1 = hmaster2_p & v22f954f | !hmaster2_p & v23fc4a3;
assign v2307a0f = stateG10_5_p & v22f7cab | !stateG10_5_p & !v10dbf64;
assign v230ab24 = hlock3_p & v12cd9b6 | !hlock3_p & v22ee024;
assign v23f443d = jx0_p & v23f52f3 | !jx0_p & v22f8f5c;
assign v23f8095 = hmaster1_p & v22fa823 | !hmaster1_p & v22f0a39;
assign v22f0b45 = stateG10_5_p & v22ed49b | !stateG10_5_p & v22fb706;
assign v23fc555 = hmaster2_p & v23fbaaa | !hmaster2_p & v23f01f8;
assign v23109e9 = hmastlock_p & v2306070 | !hmastlock_p & v84561b;
assign v230a44c = hbusreq5_p & v845620 | !hbusreq5_p & v22f915d;
assign v23fb8f4 = hlock4_p & v23117cd | !hlock4_p & !v23f216d;
assign v23f5dd2 = hbusreq4_p & v23f18a1 | !hbusreq4_p & v22fde04;
assign v23fce05 = hgrant3_p & v230d90f | !hgrant3_p & v2300774;
assign v22ef2c7 = hgrant5_p & v84561b | !hgrant5_p & v23f8b6b;
assign v22ed067 = hbusreq3_p & d962e3 | !hbusreq3_p & v22f6949;
assign v983a4e = hmaster1_p & v106a831 | !hmaster1_p & !v23f49cd;
assign v230913e = hgrant3_p & v22ee09a | !hgrant3_p & v23fcf38;
assign v2305b70 = hmaster2_p & v23f4da0 | !hmaster2_p & v230d3f5;
assign v22fcbbb = hgrant1_p & v2313463 | !hgrant1_p & !v230c2f4;
assign v2303481 = jx0_p & v84561b | !jx0_p & v23f24c0;
assign v22fe60b = hgrant1_p & v84561b | !hgrant1_p & v23f3051;
assign v22f1d1a = hbusreq3_p & v22f2bab | !hbusreq3_p & v23fc0ac;
assign v22fab50 = hmaster2_p & v23fc161 | !hmaster2_p & v23fba9a;
assign v22f72ff = hmaster0_p & v230ea9f | !hmaster0_p & v23079d8;
assign v23f04f2 = hmaster0_p & v23fbf1e | !hmaster0_p & v23f0e65;
assign v23fbf66 = hlock1_p & v106ae1c | !hlock1_p & a1fbb6;
assign v230ef5b = hbusreq1 & v230aef0 | !hbusreq1 & v845636;
assign v23111d5 = hlock3_p & v22f7659 | !hlock3_p & v23faaa0;
assign v22f1389 = locked_p & v84561b | !locked_p & v1aae087;
assign v23fb4a6 = stateG2_p & v2306d5c | !stateG2_p & !v23fbbf3;
assign v22fa77b = hmaster0_p & e1de6f | !hmaster0_p & v23fb554;
assign v12cde1b = hbusreq3_p & v22ec2a4 | !hbusreq3_p & v2305aea;
assign v22fde04 = hmaster0_p & v23f2bb6 | !hmaster0_p & v23fbf8e;
assign v22f5767 = hlock3_p & v23fc69b | !hlock3_p & !v84561b;
assign b9888a = hgrant2_p & v2310116 | !hgrant2_p & v2308a30;
assign v22fd6fb = hbusreq3_p & v22f2bab | !hbusreq3_p & v23117f5;
assign v23928cd = hbusreq2 & v22f337b | !hbusreq2 & v845620;
assign v2301f8c = hmaster0_p & v2307816 | !hmaster0_p & v22f6b3e;
assign v22f0b79 = hgrant1_p & v84561b | !hgrant1_p & v2303329;
assign v22fdbf7 = hgrant2_p & v23fb849 | !hgrant2_p & v22eb1f5;
assign v23073e6 = hbusreq6_p & v22f2851 | !hbusreq6_p & v2308dbf;
assign v23fb838 = hgrant1_p & v23fc127 | !hgrant1_p & v23fc8ea;
assign v2301797 = hgrant1_p & v23fcf74 | !hgrant1_p & v23fcd9f;
assign v22fda30 = hgrant2_p & v22fdf5b | !hgrant2_p & v230df15;
assign v22f0d89 = hlock3_p & v22fe74a | !hlock3_p & v23fcc99;
assign v2301884 = hbusreq1 & v230f5a3 | !hbusreq1 & v84561b;
assign v23fc4c3 = hmaster2_p & v23f6411 | !hmaster2_p & v22f3a35;
assign v2304dc4 = hmaster2_p & v2392ea0 | !hmaster2_p & v84564d;
assign v22fda85 = hmaster2_p & v84561b | !hmaster2_p & !v22f6741;
assign v9eaa59 = hbusreq3_p & v23fc19b | !hbusreq3_p & v22f5d84;
assign v23fd022 = stateG10_5_p & v2309ba2 | !stateG10_5_p & v845636;
assign v2306d26 = hbusreq3_p & v23107f9 | !hbusreq3_p & v22f231d;
assign v23f8976 = hbusreq3 & v23fca46 | !hbusreq3 & v84561b;
assign v230cc18 = hbusreq3_p & v22eb5a9 | !hbusreq3_p & v22ee4ab;
assign v23f4938 = stateG10_5_p & v191a973 | !stateG10_5_p & v1e83fd9;
assign v1e840b4 = hbusreq3_p & v23f58bb | !hbusreq3_p & v22fda61;
assign v23fc296 = hmaster0_p & v84561b | !hmaster0_p & v23fcb2b;
assign v22fbebb = hgrant3_p & v23fc975 | !hgrant3_p & v23fc5ab;
assign v23f1891 = hmaster2_p & v22fc564 | !hmaster2_p & !v12cc2ef;
assign v22fa6ab = hmaster2_p & v23fbf8b | !hmaster2_p & !v22f1ae7;
assign v230b6fc = jx3_p & b42c55 | !jx3_p & v23f710c;
assign v230ae4e = hmaster0_p & v23f756e | !hmaster0_p & v23fb810;
assign v2307816 = hbusreq4 & v23fc192 | !hbusreq4 & v84561b;
assign v23fcc8c = hgrant5_p & v22f39a8 | !hgrant5_p & v23fb4bd;
assign v22f46a6 = stateG10_5_p & v23fc612 | !stateG10_5_p & a07f9b;
assign v23f14ce = hmaster0_p & v230cc18 | !hmaster0_p & v22fc9cf;
assign v23fbe14 = hmaster0_p & v23f1afd | !hmaster0_p & v2312b99;
assign v22fcd06 = hgrant3_p & ad89b5 | !hgrant3_p & v22f52c3;
assign v23f23f1 = hbusreq5_p & v23fc853 | !hbusreq5_p & v23fc3c3;
assign bafb17 = hmaster2_p & v845622 | !hmaster2_p & v23fc3f2;
assign v23fc8ba = hbusreq3_p & v22f2bab | !hbusreq3_p & v230dc43;
assign v23003fc = hbusreq5_p & v845620 | !hbusreq5_p & v23fbe0d;
assign v230aef0 = hlock5_p & fc8f82 | !hlock5_p & v845636;
assign v230a407 = hbusreq6_p & v22f81a7 | !hbusreq6_p & v22f10a7;
assign v2392d45 = jx0_p & v23103f4 | !jx0_p & v84561b;
assign v23fc068 = hmaster2_p & v23fb1a4 | !hmaster2_p & !v2301e25;
assign b9ca3d = hlock5_p & v1b87673 | !hlock5_p & !v84561b;
assign v22f155f = hlock6_p & v230cffc | !hlock6_p & v22fe8a4;
assign v230d7b4 = hbusreq3 & v23fba11 | !hbusreq3 & v84561b;
assign v23fc7c7 = hmaster2_p & v10dbf64 | !hmaster2_p & v191a86f;
assign v22fc66c = hmaster2_p & a1fba6 | !hmaster2_p & v2304074;
assign v2301cf4 = hlock4_p & v22f5ea8 | !hlock4_p & !v84561b;
assign v23fc323 = hgrant3_p & v2301be6 | !hgrant3_p & v23fc58a;
assign v2310389 = hmaster2_p & v23112ad | !hmaster2_p & v22f61b6;
assign v23f1e9c = hbusreq1_p & v23fbf66 | !hbusreq1_p & a1fbb6;
assign v22fca1d = hmaster1_p & v23fc04e | !hmaster1_p & v84561b;
assign v22f217d = hgrant0_p & v84561b | !hgrant0_p & v845653;
assign v22ff0d7 = hbusreq5_p & v191ae28 | !hbusreq5_p & v84561b;
assign v23f3dd3 = hbusreq1_p & v22ffe51 | !hbusreq1_p & !v2307a62;
assign v2301d45 = hgrant5_p & v23fb3d1 | !hgrant5_p & v22f84ff;
assign v22f7dbc = hmaster2_p & v2306d29 | !hmaster2_p & v23fc904;
assign v23044f6 = hgrant3_p & v84562e | !hgrant3_p & v22f1713;
assign v22f89c7 = jx1_p & v22ec21e | !jx1_p & v231220c;
assign v2305a79 = hbusreq1_p & v230a25a | !hbusreq1_p & a1fe3e;
assign v230de50 = hgrant1_p & v23fb47e | !hgrant1_p & v2392809;
assign bd6575 = jx0_p & v977ddf | !jx0_p & v84561b;
assign a2cc4e = hmaster1_p & v2310317 | !hmaster1_p & v1aae9f4;
assign v23fcf99 = hbusreq4_p & v23f904c | !hbusreq4_p & v23fb965;
assign v23050ee = jx0_p & v23028ef | !jx0_p & v230539c;
assign v22f8bcf = hbusreq5 & v22ef513 | !hbusreq5 & v84561b;
assign v22ecbc3 = hbusreq3_p & v84562a | !hbusreq3_p & v2311214;
assign v2301eb1 = hlock1_p & v22f8f3d | !hlock1_p & v23fcaeb;
assign v23104a1 = jx1_p & v239162d | !jx1_p & v23f1908;
assign v23fa69c = hgrant1_p & v84561b | !hgrant1_p & v23fb89e;
assign v23f42ec = hbusreq6_p & v23fbf06 | !hbusreq6_p & !v22f639d;
assign v22ee660 = hbusreq2 & v23f1207 | !hbusreq2 & v22f42bd;
assign v2301934 = hbusreq1 & v22fbb54 | !hbusreq1 & v22f7241;
assign v22f3466 = hmaster0_p & v230814d | !hmaster0_p & v96c563;
assign v23fcbe9 = hmaster2_p & bdc4e2 | !hmaster2_p & v22f6358;
assign v23f3856 = hlock3_p & v22f3af7 | !hlock3_p & !v84561b;
assign v23fd040 = hgrant2_p & v84561b | !hgrant2_p & !v22eedf9;
assign v22fed40 = hmaster0_p & v23f3d38 | !hmaster0_p & a5666b;
assign v2392f02 = hlock3_p & v2300c56 | !hlock3_p & v22f5218;
assign v23fc1a1 = hmaster0_p & v23fccc1 | !hmaster0_p & !v22fb1d7;
assign v22f9b30 = hbusreq4_p & v990272 | !hbusreq4_p & v2392222;
assign v23082fe = hlock3_p & v230ad1e | !hlock3_p & v23f6843;
assign v22f8cb7 = hlock0_p & v845620 | !hlock0_p & v2302a2c;
assign v22f2195 = hgrant0_p & v2302c28 | !hgrant0_p & v230aec0;
assign v22ebb8e = hbusreq4 & v23916d5 | !hbusreq4 & v22f2ca2;
assign v230c3aa = hmaster0_p & v23f3915 | !hmaster0_p & v2312f4f;
assign v22f9eb0 = hmaster2_p & v22f411f | !hmaster2_p & v22f1244;
assign v23fc042 = hbusreq2_p & v23f404a | !hbusreq2_p & v845620;
assign v23f450b = hbusreq0 & v22fba61 | !hbusreq0 & v84561b;
assign v23fc1ec = hmaster0_p & v23fc3e8 | !hmaster0_p & v23fc7a7;
assign v230a775 = hmaster0_p & v84561b | !hmaster0_p & v2302370;
assign v23f19e4 = hbusreq1_p & v23fbf63 | !hbusreq1_p & f40a9e;
assign a1fe03 = hbusreq1 & v2392f6b | !hbusreq1 & !v84562a;
assign v191abf8 = jx2_p & v84561b | !jx2_p & v22f89d5;
assign v22fe2d5 = hlock3_p & v23f9452 | !hlock3_p & v23f35c7;
assign v23126b7 = hbusreq6_p & v22eee15 | !hbusreq6_p & v23088a9;
assign v22fa245 = hlock2_p & v22ebbea | !hlock2_p & !v230f5a3;
assign v2300bc5 = hgrant4_p & v230d65b | !hgrant4_p & v22f7d5c;
assign v22f5a2a = hbusreq5 & v2300de3 | !hbusreq5 & v84561b;
assign v84562b = hlock2_p & v84561b | !hlock2_p & !v84561b;
assign v230806a = hmaster2_p & v23fc71d | !hmaster2_p & v230910b;
assign v23fab11 = hlock3_p & v23fb62c | !hlock3_p & !v1e840fa;
assign v23fa967 = hmaster0_p & v23fc6a1 | !hmaster0_p & v230e857;
assign b60876 = hbusreq5_p & v230f9c8 | !hbusreq5_p & v84561b;
assign v23f63ab = hlock5_p & v22f448b | !hlock5_p & !v845636;
assign v22fea98 = hmaster2_p & v22fe421 | !hmaster2_p & v23f6b67;
assign v22fe963 = hbusreq0 & v2302e32 | !hbusreq0 & !v84561b;
assign v230f2dc = hbusreq0_p & v22f2db0 | !hbusreq0_p & v1aae98c;
assign v22efd62 = hbusreq0_p & v230a63b | !hbusreq0_p & v845629;
assign v23fcaad = hlock3_p & v22ed72b | !hlock3_p & v22ed5c8;
assign v23fc26c = hmaster0_p & v23faa0a | !hmaster0_p & v23fba16;
assign v22fe74a = hbusreq3_p & v23fc7b4 | !hbusreq3_p & v84561b;
assign v22ffc69 = hlock0_p & v191a876 | !hlock0_p & v2300474;
assign v23fb933 = hbusreq3_p & v2303fd8 | !hbusreq3_p & v84561b;
assign v23fbb48 = hmaster2_p & v22ff120 | !hmaster2_p & v23fc84e;
assign v23035f1 = hmaster2_p & v231171d | !hmaster2_p & v22f2883;
assign v2305bf5 = hbusreq6 & v22eaf81 | !hbusreq6 & v84561b;
assign v22f3c10 = hbusreq6_p & v23fc104 | !hbusreq6_p & v84561b;
assign v2306aef = hmaster2_p & v22f9927 | !hmaster2_p & v23fb966;
assign v2391b49 = hgrant2_p & v84561b | !hgrant2_p & !v230164e;
assign v23f7503 = hgrant3_p & v22f3643 | !hgrant3_p & v2393f95;
assign v2302f12 = jx1_p & v23129d7 | !jx1_p & v23fbad9;
assign v845651 = hgrant1_p & v84561b | !hgrant1_p & !v84561b;
assign v23fc24c = hlock4_p & v23fbca2 | !hlock4_p & !v84561b;
assign v23fc5d9 = hgrant1_p & v84561b | !hgrant1_p & v2308748;
assign v230c0e6 = hmaster2_p & v23fc89a | !hmaster2_p & !v23fbbf2;
assign v230a413 = stateA1_p & v22ef862 | !stateA1_p & !v863ce5;
assign v22fd9be = hmastlock_p & v23f732a | !hmastlock_p & v84561b;
assign v2308ae2 = stateA1_p & v84561b | !stateA1_p & v23f68bf;
assign v23fcd70 = hmaster2_p & v22fd696 | !hmaster2_p & v22f6671;
assign v22eb51e = hmaster2_p & v84564d | !hmaster2_p & v22f3643;
assign v23f5c2f = hmaster0_p & v230cc18 | !hmaster0_p & v23fcc9f;
assign v2306822 = hmaster1_p & v22ee93b | !hmaster1_p & !v22fe985;
assign v23fb69d = hbusreq1_p & v23fb591 | !hbusreq1_p & v22fdce0;
assign v23fbee2 = hbusreq3_p & v23f9870 | !hbusreq3_p & e1e353;
assign v22fdaf3 = hmaster0_p & v23fabb8 | !hmaster0_p & !v23075ce;
assign v23f4926 = hmaster2_p & v22fc2bd | !hmaster2_p & v84561b;
assign v23f1c12 = hgrant6_p & v23fb8f7 | !hgrant6_p & v230f82f;
assign v23fb811 = hgrant5_p & v22ef92c | !hgrant5_p & !v23fc9b9;
assign bdeff3 = hbusreq4 & v23fb8e4 | !hbusreq4 & v845627;
assign v23fbd53 = hbusreq1 & v191a86f | !hbusreq1 & v84561b;
assign v23fc387 = hmaster2_p & v23018c4 | !hmaster2_p & v15072a9;
assign v22fb706 = hgrant0_p & v23126ae | !hgrant0_p & v22f6a6b;
assign f405e4 = hmaster2_p & v84564d | !hmaster2_p & !v84561b;
assign v22edd3d = hbusreq4 & v191afef | !hbusreq4 & v230bbda;
assign v2309282 = hbusreq3_p & v23fce9e | !hbusreq3_p & v84561b;
assign v2307eb9 = hgrant3_p & v84561b | !hgrant3_p & v22ff90b;
assign v23fbe02 = hmaster2_p & v2306d29 | !hmaster2_p & v23070c1;
assign v23040af = hmastlock_p & v2301d2f | !hmastlock_p & v84561b;
assign e1de18 = hbusreq0 & v23fc514 | !hbusreq0 & !v22f91c9;
assign v23f361e = hbusreq3_p & v23fc46d | !hbusreq3_p & v23fc4fc;
assign v22f30bb = jx0_p & b7d0f1 | !jx0_p & v84561b;
assign v23038a2 = hbusreq5_p & v9526ac | !hbusreq5_p & v22fc1be;
assign v2311255 = locked_p & v84561b | !locked_p & v22f2718;
assign v22fc3ed = hready & v2304ec7 | !hready & v22f92f9;
assign v13aff5b = hbusreq0 & v2311255 | !hbusreq0 & v84561b;
assign v2301968 = hmaster0_p & v22f8613 | !hmaster0_p & v23fcc39;
assign v2304c86 = hmaster0_p & bd74ba | !hmaster0_p & v23fb9d6;
assign v230da9b = hbusreq4 & v22f3cc0 | !hbusreq4 & v23fc223;
assign v22f60c6 = locked_p & v22f37c1 | !locked_p & !v84561b;
assign v106af55 = hbusreq5_p & v23f19b4 | !hbusreq5_p & v2312020;
assign v23068bf = hgrant6_p & v2305ea5 | !hgrant6_p & v23f699c;
assign v22f481f = hbusreq5_p & v22fa345 | !hbusreq5_p & v22f549a;
assign v995fa2 = hgrant5_p & f40dab | !hgrant5_p & v23f3adc;
assign v22f108e = hgrant5_p & v23012c6 | !hgrant5_p & v9f009f;
assign v22fee59 = jx0_p & v22fed90 | !jx0_p & v22f8f70;
assign v22ebd72 = hgrant3_p & v84561b | !hgrant3_p & v23112ad;
assign v2300523 = hmaster2_p & v23fc38f | !hmaster2_p & v22fe940;
assign v23f00cf = stateG2_p & v84561b | !stateG2_p & !v2305aa1;
assign v9b1253 = hmaster1_p & v84561b | !hmaster1_p & v23efd4b;
assign v23fcea2 = hgrant3_p & v230965a | !hgrant3_p & baa026;
assign v2300d93 = hmaster2_p & v22f98e3 | !hmaster2_p & !v22f03cf;
assign v22fea26 = hbusreq3_p & v23f1b3c | !hbusreq3_p & v23fcc35;
assign v22ed805 = hbusreq3 & v23f97bb | !hbusreq3 & v84561b;
assign v22fa655 = jx1_p & v85fd50 | !jx1_p & v85fc1a;
assign v230e02e = hbusreq3_p & v84561b | !hbusreq3_p & v23124c5;
assign v2304ad5 = hgrant1_p & v84561b | !hgrant1_p & v23fc3ff;
assign v106af4d = hgrant2_p & v23fcbb5 | !hgrant2_p & !v191a86f;
assign v23fc11b = hmaster0_p & v22efd02 | !hmaster0_p & v22f8cb9;
assign v22eb3bc = hbusreq4 & a9da2d | !hbusreq4 & v230dd28;
assign v966100 = hbusreq4 & v23fca1c | !hbusreq4 & v84561b;
assign v23f36d3 = jx2_p & v191b107 | !jx2_p & v22faa4b;
assign v23fa6eb = hmaster0_p & v23f9fdc | !hmaster0_p & v230c97c;
assign v22f4163 = hlock0_p & v23fa2ec | !hlock0_p & v2312cf2;
assign v23f403e = hmaster2_p & v106ae1c | !hmaster2_p & v2301a3f;
assign v230dffa = hbusreq5 & v23fbfd0 | !hbusreq5 & v22f11f6;
assign v22fa987 = hbusreq4 & v22ee9be | !hbusreq4 & v23f1812;
assign v22fbf21 = hmaster2_p & v22f5e91 | !hmaster2_p & v2308765;
assign v230e7d6 = hmaster0_p & v23f600f | !hmaster0_p & v23fc284;
assign v23f54a0 = hbusreq4 & v22f640a | !hbusreq4 & !v84561b;
assign v23fb122 = hlock5_p & v23fc3c9 | !hlock5_p & v23f22a1;
assign v22f006c = hgrant6_p & v84561b | !hgrant6_p & v12cc315;
assign v2300962 = hbusreq2 & fc8ab7 | !hbusreq2 & !v84561b;
assign v2312050 = hmaster0_p & v22f25ae | !hmaster0_p & !v23037ac;
assign v23083c1 = hmaster2_p & v23fc7d5 | !hmaster2_p & v230cbdd;
assign v23f724e = hbusreq6_p & v23fba4a | !hbusreq6_p & !v23f5474;
assign v23fb7da = hlock3_p & v12cd534 | !hlock3_p & v22edf79;
assign v23001d6 = hgrant1_p & v230f9db | !hgrant1_p & v23fc545;
assign v23fc2a7 = hgrant0_p & v84561b | !hgrant0_p & !v2303a7f;
assign v23fcaa6 = hgrant5_p & v2304db3 | !hgrant5_p & v23f1f21;
assign v23fcd45 = hlock6_p & v22f6463 | !hlock6_p & v230b1ab;
assign v22eba1d = hbusreq6 & v84564d | !hbusreq6 & v23fa2ec;
assign v22ef983 = hlock5_p & v191aa68 | !hlock5_p & v191a86f;
assign v230c4ae = hmaster2_p & v2391d40 | !hmaster2_p & v22f1ae5;
assign v230c034 = hbusreq3_p & v2306690 | !hbusreq3_p & v230282c;
assign v23f5474 = hbusreq4_p & b3d617 | !hbusreq4_p & v22f18a3;
assign v22efceb = hbusreq4 & v23089f7 | !hbusreq4 & v22fb009;
assign v23f9193 = hmaster0_p & v191ab52 | !hmaster0_p & v23fca40;
assign v23057ba = hgrant3_p & v12cd6a2 | !hgrant3_p & v2306fb7;
assign v23fbe69 = hbusreq6_p & v230c322 | !hbusreq6_p & v23fc297;
assign v22fe370 = hbusreq3_p & v13afb6e | !hbusreq3_p & v2309783;
assign v23fcd0f = hgrant1_p & v23f7700 | !hgrant1_p & v23fc39c;
assign v2309b67 = hlock6_p & v2392122 | !hlock6_p & !v84561b;
assign v2305296 = hmaster2_p & v23fc957 | !hmaster2_p & v23fc6a0;
assign v23fc989 = hbusreq6_p & v23f38b1 | !hbusreq6_p & v22f4f0f;
assign v23f6acc = hbusreq3_p & v22f2c72 | !hbusreq3_p & v84561b;
assign v2311f99 = hmaster0_p & v84561b | !hmaster0_p & !v22ebb85;
assign v106a888 = hbusreq4 & v23067de | !hbusreq4 & v23f91bc;
assign v230c66e = hbusreq3_p & v230c2ff | !hbusreq3_p & v2309be5;
assign v239174f = hbusreq4 & v23fca46 | !hbusreq4 & v84561b;
assign v22fc493 = jx1_p & v84561b | !jx1_p & v23fc6b2;
assign v230e8a0 = hmaster2_p & v1aadac4 | !hmaster2_p & v84561b;
assign v22fd5fc = hbusreq6_p & v23f5b31 | !hbusreq6_p & v23fcf52;
assign v97f5b6 = hmaster2_p & v22f8c43 | !hmaster2_p & v22f61b6;
assign v23f2bb6 = hgrant3_p & v23fc473 | !hgrant3_p & v23fcd74;
assign v22f00eb = hmaster0_p & v23f7039 | !hmaster0_p & v230f760;
assign v23f18da = hbusreq3_p & v23fcdc1 | !hbusreq3_p & v22ed8fe;
assign v22ec7cf = hlock3_p & v22fc98d | !hlock3_p & v23fb93c;
assign v23000cf = hlock0_p & v22f13cb | !hlock0_p & v2392adb;
assign v230ecb1 = hbusreq6 & v23f85b6 | !hbusreq6 & !v84562d;
assign v22f9392 = hmaster0_p & v22eeb7a | !hmaster0_p & !v23fcb9c;
assign v23f7158 = hlock3_p & v84561b | !hlock3_p & v23fca55;
assign v23f3b81 = hbusreq6 & v22f45e9 | !hbusreq6 & v84561b;
assign aca9e4 = hbusreq5_p & v84564d | !hbusreq5_p & v84561b;
assign v2393501 = hbusreq1_p & v230b313 | !hbusreq1_p & v22f06fb;
assign v22fb151 = hgrant3_p & v84561b | !hgrant3_p & v23f35c2;
assign v23fa08a = jx1_p & b533b5 | !jx1_p & v22ec5ac;
assign aba695 = hmaster2_p & v2311810 | !hmaster2_p & v23fb1c6;
assign v230a3e2 = hmaster0_p & v23fc57e | !hmaster0_p & v22f3d18;
assign v23fbd33 = hlock3_p & v22ede9f | !hlock3_p & v22fd8c5;
assign v22ef292 = hmaster0_p & v230f18c | !hmaster0_p & v23f76fb;
assign v23fca4a = hbusreq4_p & v23039ea | !hbusreq4_p & v22f5521;
assign v2305498 = hbusreq4_p & v12cda8f | !hbusreq4_p & v230432b;
assign v22f0ea8 = hmaster0_p & v23f3c00 | !hmaster0_p & !v230a934;
assign v23fbdf1 = hgrant0_p & v845629 | !hgrant0_p & v21eabbd;
assign v23fd037 = hbusreq6 & v22ebce1 | !hbusreq6 & v23fcd8d;
assign v22eb8fb = jx0_p & v22fcf35 | !jx0_p & v2311cea;
assign v230e1f2 = hmaster2_p & v8d360e | !hmaster2_p & !v13afe8f;
assign v22f4619 = hmaster1_p & v22f8cb9 | !hmaster1_p & v2393142;
assign v23fbf36 = hmaster2_p & v22fc8e5 | !hmaster2_p & v84561b;
assign v23fbf74 = hbusreq6 & v2304452 | !hbusreq6 & v23fc9fb;
assign v23fc9f1 = hgrant2_p & v23fc9c6 | !hgrant2_p & !v23fb61f;
assign v22edf86 = hmaster1_p & v23fbf8d | !hmaster1_p & v230fe65;
assign v23f20a8 = hmaster0_p & v230f75b | !hmaster0_p & b00aa6;
assign v22f037f = hlock6_p & v22f320d | !hlock6_p & v23fcb90;
assign v2306bc5 = hbusreq4_p & v22f2ff1 | !hbusreq4_p & v22fcaa6;
assign v2312917 = hmaster2_p & v23fbfce | !hmaster2_p & v23fbde0;
assign v22f3840 = hgrant3_p & v22f8838 | !hgrant3_p & v22eeb27;
assign v230ac9e = hlock0_p & da38c1 | !hlock0_p & v23fce3d;
assign v22f25ae = hgrant3_p & v98d402 | !hgrant3_p & v22f26f5;
assign v23fc347 = hmaster2_p & v191a86f | !hmaster2_p & v22fa5a5;
assign v23f4cc1 = hmaster0_p & v22ef62d | !hmaster0_p & v230eab7;
assign b79082 = hgrant1_p & v845620 | !hgrant1_p & v23f7de2;
assign v23fb99d = hbusreq1_p & v15075a6 | !hbusreq1_p & !v84561b;
assign v22fa3fa = hbusreq6 & v22ff4af | !hbusreq6 & v22f5fb4;
assign v22ed6ee = hbusreq0 & v23fbac1 | !hbusreq0 & v84561b;
assign v22ed1b0 = hmaster0_p & v22f2009 | !hmaster0_p & v22fc92d;
assign v2309897 = hgrant3_p & v23fc6f1 | !hgrant3_p & v2311a27;
assign v22f0c75 = hmaster1_p & v2303ce3 | !hmaster1_p & v23fbd21;
assign v22fa6f5 = hmaster2_p & v23046f7 | !hmaster2_p & !v22eb5b3;
assign v23fc966 = hbusreq6_p & v23f1a1f | !hbusreq6_p & !v84561b;
assign v22f12fb = hbusreq3_p & v2300ab9 | !hbusreq3_p & c0aa95;
assign v23fc4d0 = hmaster2_p & v23fcf40 | !hmaster2_p & v2304402;
assign v22f56c2 = hlock3_p & v22f10d6 | !hlock3_p & v230e43d;
assign v23f66e6 = hbusreq1 & v23fcc8c | !hbusreq1 & v84561b;
assign v23f846c = hmaster0_p & v2393485 | !hmaster0_p & v22fe1c8;
assign v23fbd2e = hlock1_p & v2305fe0 | !hlock1_p & v84564d;
assign v22ecd9e = hmaster0_p & v22ed01c | !hmaster0_p & v23f15a7;
assign v230a744 = hlock3_p & v2303061 | !hlock3_p & !v23f9d0b;
assign v230ceb6 = hbusreq2_p & v23fc411 | !hbusreq2_p & a1fba6;
assign v230d529 = hbusreq0_p & v22edd64 | !hbusreq0_p & v84561b;
assign v23fbef7 = hbusreq0 & v23fcc10 | !hbusreq0 & v84561b;
assign v23f4edf = jx2_p & v23fba9c | !jx2_p & v2308ac3;
assign v23fc485 = hmaster2_p & v84561b | !hmaster2_p & !v2304b4e;
assign b3d617 = hmaster0_p & v2392d61 | !hmaster0_p & v23fcf5b;
assign v23f3a8b = hlock0_p & v23fc1c1 | !hlock0_p & v23fc4fb;
assign v1aad63a = hbusreq5_p & v22f898b | !hbusreq5_p & v23fb94d;
assign v230cb7a = hbusreq5_p & v239254b | !hbusreq5_p & v230c428;
assign v22f3000 = hgrant5_p & v23fc12b | !hgrant5_p & v23fc9d2;
assign v23fb4d1 = hgrant2_p & v23fb1b4 | !hgrant2_p & v23fb473;
assign v2309a44 = hlock2_p & v2313463 | !hlock2_p & !v84561b;
assign v23104c1 = hmaster1_p & v230a36f | !hmaster1_p & v22f88f9;
assign v2305833 = hgrant5_p & v84561b | !hgrant5_p & v8f4f78;
assign v22ef8a9 = hbusreq6 & v23f3c12 | !hbusreq6 & v23efe71;
assign bda6cc = hmaster0_p & v23fb9b6 | !hmaster0_p & !bd75f3;
assign v23f4267 = hbusreq1_p & v23fbeb0 | !hbusreq1_p & !v230f34c;
assign v13afbf0 = hbusreq4 & v23045c3 | !hbusreq4 & v84561b;
assign v23fc6b2 = hmaster1_p & v23050fb | !hmaster1_p & v22fc689;
assign v22f860b = hbusreq5_p & v2306b2e | !hbusreq5_p & !v23fbbf2;
assign v2308a8f = hmaster2_p & v84561b | !hmaster2_p & v23003cc;
assign v22f509a = jx0_p & v23fb8fb | !jx0_p & v23fbe85;
assign v22f43cf = hbusreq5_p & v2307e48 | !hbusreq5_p & v2304edd;
assign v22f78ef = hbusreq0 & v22fd3f7 | !hbusreq0 & v84561b;
assign v230ad1e = hbusreq3_p & v23fcae0 | !hbusreq3_p & v23f6843;
assign v23f3c98 = hmaster0_p & baa026 | !hmaster0_p & v22f5de1;
assign v13afad7 = hbusreq4 & v23fbb44 | !hbusreq4 & v84561b;
assign v23f3eda = hgrant3_p & v2304118 | !hgrant3_p & v22fbde2;
assign v22fd2ec = hbusreq1_p & v22f7d5d | !hbusreq1_p & !v22fccf1;
assign v23fcfce = hmaster0_p & v23f232d | !hmaster0_p & v23fbb9c;
assign v22f4a7a = stateG10_5_p & v12cd9c9 | !stateG10_5_p & !v106ae19;
assign v23fb97e = jx0_p & v22f28f7 | !jx0_p & v2304d26;
assign v22f457a = hbusreq6_p & v2311f22 | !hbusreq6_p & !v23fbb7b;
assign v22ebee0 = hbusreq0 & v23fc93e | !hbusreq0 & v84562a;
assign v23fc0a0 = hmaster2_p & v22f7b29 | !hmaster2_p & v22feafc;
assign v22fe907 = jx0_p & v22f5944 | !jx0_p & v22fe188;
assign v230278d = hbusreq4_p & v2300c06 | !hbusreq4_p & v23fd026;
assign v230b304 = hmaster2_p & v23031c2 | !hmaster2_p & v23f4da0;
assign v2312a98 = hlock4_p & v23fb52f | !hlock4_p & v23fcd47;
assign v22f78de = hgrant5_p & v23fb501 | !hgrant5_p & v23f81cf;
assign v22ffa1b = hmaster0_p & v2302514 | !hmaster0_p & v23f6650;
assign v23fb869 = hbusreq3_p & v23f344d | !hbusreq3_p & !v84561b;
assign v23fbdfd = hbusreq6 & v2308331 | !hbusreq6 & v23030ad;
assign v22f0dc0 = hmaster0_p & v23087bc | !hmaster0_p & v22ec4d6;
assign v230d6c1 = hbusreq0_p & v22f64e0 | !hbusreq0_p & !v23fb12a;
assign v9ab66e = stateG10_5_p & v9f009f | !stateG10_5_p & v23fa2ec;
assign v23fbdc6 = hgrant6_p & v22f82f1 | !hgrant6_p & v23fba4d;
assign v23faada = hmaster0_p & v23fbf3e | !hmaster0_p & v2304b49;
assign bd74f4 = hmaster2_p & v22f220a | !hmaster2_p & v23f8928;
assign v2307e4f = hbusreq0 & v23fbfd0 | !hbusreq0 & b9d02f;
assign v23fc340 = hmaster2_p & v23102d5 | !hmaster2_p & v22f0132;
assign v230b08b = hmaster2_p & v23f3d14 | !hmaster2_p & v1aad38a;
assign v95adb3 = hbusreq1_p & v23fca56 | !hbusreq1_p & v23015a7;
assign v22fc452 = hbusreq3_p & v22ee95f | !hbusreq3_p & !v23124c5;
assign v12cd538 = hmaster0_p & v23fcaad | !hmaster0_p & v230a4f1;
assign v23fc678 = hmaster1_p & v84561b | !hmaster1_p & v22fd48a;
assign v2300f96 = hbusreq1 & v84561b | !hbusreq1 & v845622;
assign bd7c9b = hbusreq1 & v8d360e | !hbusreq1 & v84561b;
assign v23fb1d7 = hready_p & v23f6013 | !hready_p & v23fbd8e;
assign v2307c9a = hbusreq4_p & v230b789 | !hbusreq4_p & v23fc05d;
assign v23fc04f = hmaster2_p & v84561b | !hmaster2_p & !v22ed7ba;
assign v2307779 = hbusreq1_p & v84561b | !hbusreq1_p & v23fa9c5;
assign v22f39b0 = hbusreq2 & v1aae29a | !hbusreq2 & v23f8364;
assign v23064ae = hlock0_p & v84561b | !hlock0_p & v230e40a;
assign v22ef109 = hmaster2_p & v23022b1 | !hmaster2_p & !v23fb9ad;
assign v23119a4 = hmaster1_p & v22fb1d6 | !hmaster1_p & v22f421a;
assign v23051eb = hbusreq3 & v230a56a | !hbusreq3 & v2312ef7;
assign v2312290 = hmaster0_p & v22f2281 | !hmaster0_p & v239315b;
assign v2306f3c = hmaster2_p & v230bdd0 | !hmaster2_p & v23fcb83;
assign v23fc1a2 = hbusreq3 & v2308a8f | !hbusreq3 & v84561b;
assign v230fa92 = hbusreq0 & v1aae087 | !hbusreq0 & v84561b;
assign v2310da2 = hbusreq5 & v22eb5b3 | !hbusreq5 & !v84561b;
assign v23fb849 = hbusreq2_p & v2309377 | !hbusreq2_p & !v22fd25c;
assign v22ec89f = hgrant1_p & v2307375 | !hgrant1_p & v22ff13f;
assign v22ed975 = hgrant3_p & v22f064a | !hgrant3_p & v23fa8c7;
assign v23f5dcc = hmaster2_p & v22eefd1 | !hmaster2_p & v84561b;
assign v23fba74 = hmaster2_p & v22fe920 | !hmaster2_p & v23f052e;
assign v23f2d60 = hmaster0_p & v22f4d74 | !hmaster0_p & v2392aaa;
assign v23fcf8a = hmaster2_p & v22f85a0 | !hmaster2_p & v22fa064;
assign v23fbc3a = hgrant3_p & v230f14b | !hgrant3_p & v2308d5a;
assign v22fb112 = hmaster0_p & v2308e08 | !hmaster0_p & v230b3a5;
assign jx2 = v123d721;
assign v23fcfd1 = jx1_p & v22f62e3 | !jx1_p & v23009d5;
assign v22fc6ca = hlock3_p & v22f4fb8 | !hlock3_p & v23fbe27;
assign v231188f = hbusreq6_p & v23fcea5 | !hbusreq6_p & v2391b52;
assign v23fba9b = stateG10_5_p & v22f316f | !stateG10_5_p & v106a782;
assign v23fc1ac = hmaster1_p & v84561b | !hmaster1_p & v23fc684;
assign v2301a7e = hmaster1_p & v23f1a2b | !hmaster1_p & !bc87ee;
assign v230c579 = hbusreq1_p & v23fbf59 | !hbusreq1_p & v84561b;
assign v230abfb = hready & v23fc491 | !hready & !v84561b;
assign v23fb2f7 = hbusreq1_p & v23f6411 | !hbusreq1_p & !b9d013;
assign v23f5c9b = hbusreq0_p & v230446f | !hbusreq0_p & !v23036ca;
assign v230a63b = hbusreq0 & a476c2 | !hbusreq0 & v84561b;
assign v2306f7b = hgrant5_p & v22f3ca0 | !hgrant5_p & v22feb95;
assign v2391a89 = hgrant0_p & v230bd6c | !hgrant0_p & v22f03ce;
assign v23fbf46 = hgrant5_p & v230b011 | !hgrant5_p & v23fd049;
assign v230d5a9 = hlock3_p & v230e02e | !hlock3_p & !v22fc452;
assign v2309294 = hmaster0_p & v23f29e9 | !hmaster0_p & v23f3321;
assign v23fc7ab = hbusreq3 & v22ebc9f | !hbusreq3 & v23fba9a;
assign v23fcb16 = jx1_p & a1fd70 | !jx1_p & v22f0c75;
assign v23f79a0 = hbusreq5 & v2301f92 | !hbusreq5 & !v84561b;
assign v2312009 = jx1_p & v2300e70 | !jx1_p & v23fc786;
assign v23fccd7 = hmaster0_p & v23fccc2 | !hmaster0_p & v84561b;
assign v22fa068 = stateG10_5_p & v23f1f3e | !stateG10_5_p & v84561b;
assign v22ec1a8 = hbusreq4_p & v23fcbd8 | !hbusreq4_p & v230713e;
assign v23f664b = hmaster0_p & v22f9cee | !hmaster0_p & v230be28;
assign v2303d8f = hbusreq0 & v23023c9 | !hbusreq0 & v845620;
assign v22ee0c4 = hready & v22ed8c2 | !hready & !v84561b;
assign v23fbe09 = hgrant5_p & v22ff890 | !hgrant5_p & v230b8cd;
assign v2312f81 = hmaster2_p & v23fa2ec | !hmaster2_p & v84561b;
assign v23f9680 = hgrant1_p & v22ec09c | !hgrant1_p & v230e2d8;
assign v2301b00 = hmaster2_p & v84564d | !hmaster2_p & v22fef02;
assign b00b0b = decide_p & v230812e | !decide_p & v230ca71;
assign v230144a = hlock6_p & v230ed77 | !hlock6_p & bd7530;
assign v2311fb5 = hmaster2_p & v1aae362 | !hmaster2_p & fc8ab7;
assign v22fcabb = hbusreq4_p & v2300995 | !hbusreq4_p & v23fc0d4;
assign v23fa1ad = hbusreq1_p & v2310f5b | !hbusreq1_p & v84561b;
assign v2308b02 = hmaster2_p & v22fa5fd | !hmaster2_p & v1aad38a;
assign v23f5ae3 = hlock6_p & v22eb4a6 | !hlock6_p & b208fd;
assign v23fc4b4 = hbusreq5_p & v22fa345 | !hbusreq5_p & v2392ed3;
assign v23f3955 = hgrant3_p & v2303415 | !hgrant3_p & v23fb8cb;
assign v2309598 = hbusreq0_p & v9526ac | !hbusreq0_p & v2304074;
assign v22ef55f = hbusreq6_p & v230b77c | !hbusreq6_p & !v84561b;
assign b0fc7a = hlock4_p & v2303822 | !hlock4_p & v22eff53;
assign v22f023b = hmaster2_p & v22f4cf3 | !hmaster2_p & !v13afe3a;
assign v23f111c = hbusreq1_p & v230cb59 | !hbusreq1_p & v84561b;
assign v23f5b7b = hbusreq1 & v2309b39 | !hbusreq1 & !v23fc614;
assign v22f9c2f = hgrant1_p & v17a34ff | !hgrant1_p & !v230dd9e;
assign v22f8db2 = stateA1_p & v2302ca3 | !stateA1_p & v23fba7e;
assign v23f917f = hmaster0_p & ae78a6 | !hmaster0_p & v2346b79;
assign v22f7aff = hbusreq5_p & v2306d29 | !hbusreq5_p & v23126ae;
assign v23fceb3 = hburst0_p & v23fc683 | !hburst0_p & !v230cb1f;
assign v23936a3 = hmaster2_p & v84561b | !hmaster2_p & !v23068a9;
assign v23fc941 = hbusreq4_p & bd7c6a | !hbusreq4_p & v22f3519;
assign v231138f = hbusreq4_p & v23fb670 | !hbusreq4_p & !v22edc69;
assign v23028f6 = hbusreq3_p & v2311e39 | !hbusreq3_p & v23fc99a;
assign v23fa825 = hmaster0_p & v22ed711 | !hmaster0_p & !bd74e7;
assign v22fba61 = hgrant2_p & v23f73a4 | !hgrant2_p & !v22f79fb;
assign v230c1dd = hgrant3_p & v23fbc82 | !hgrant3_p & !v84561b;
assign v86a21a = hmaster0_p & v230ad0f | !hmaster0_p & v23fc327;
assign v2307f3f = hbusreq3 & v23fc983 | !hbusreq3 & v23fcea3;
assign v22f7100 = hgrant5_p & v2391c8a | !hgrant5_p & v238b0d7;
assign v23064ce = hmaster2_p & v23fc48e | !hmaster2_p & v23101b1;
assign v22fec1c = hlock3_p & v23fbcca | !hlock3_p & v23fc18b;
assign v230828b = hlock0_p & v84562a | !hlock0_p & v230e551;
assign v230f072 = hbusreq4 & v231398c | !hbusreq4 & v22fe408;
assign v2307eac = hbusreq4_p & v22f8cb9 | !hbusreq4_p & v9ed019;
assign v23fbe2a = hgrant3_p & v23fb5a4 | !hgrant3_p & v22fbc47;
assign v23fb899 = hbusreq5 & v22fca61 | !hbusreq5 & v84561b;
assign v23fc91d = hmaster0_p & v84561b | !hmaster0_p & v22f8e0c;
assign v23fc8e6 = hmaster1_p & v22f8e53 | !hmaster1_p & !v23f49cd;
assign v23fb976 = hgrant3_p & v84561b | !hgrant3_p & v22f3c11;
assign v22fe3f6 = hgrant5_p & v23fc8a8 | !hgrant5_p & v84561b;
assign v22f092c = hgrant3_p & v84561b | !hgrant3_p & afb25b;
assign v23f8f25 = hgrant1_p & v23f4b28 | !hgrant1_p & v2312912;
assign v22fb8d6 = hbusreq1_p & v22f15fe | !hbusreq1_p & v2393ac5;
assign v23fb578 = hmaster2_p & v22f2718 | !hmaster2_p & v84561b;
assign v2307729 = hbusreq5_p & v23f4d1c | !hbusreq5_p & v23054ba;
assign v230db4e = hgrant1_p & v2300437 | !hgrant1_p & v22efc42;
assign v22f299d = hbusreq6_p & v239196f | !hbusreq6_p & v23fc46e;
assign v22f57ea = hmaster0_p & v22f9d92 | !hmaster0_p & !v22fd799;
assign v23fb44f = hbusreq1 & v230446f | !hbusreq1 & !v84562a;
assign v2306595 = stateG2_p & v84561b | !stateG2_p & !v845667;
assign v22f3be4 = hbusreq0 & v84564d | !hbusreq0 & !v84561b;
assign v22f7241 = hgrant5_p & v2304db3 | !hgrant5_p & v23f40ba;
assign v23fbe60 = hgrant1_p & v12cc2ef | !hgrant1_p & v230259a;
assign v23f6d9c = hbusreq1_p & v22f6385 | !hbusreq1_p & v22f6e29;
assign v22f5437 = hmaster2_p & v22f542d | !hmaster2_p & v22f26fc;
assign v23fbd16 = hbusreq2_p & v22f15fe | !hbusreq2_p & !v84561b;
assign a1f77b = hbusreq1_p & v23fc89a | !hbusreq1_p & v22f4587;
assign v2301482 = hbusreq5_p & v23f8c71 | !hbusreq5_p & v230fa13;
assign v2309dce = hmaster0_p & v23fb845 | !hmaster0_p & v2310ada;
assign v22f8985 = hbusreq3_p & v23f8607 | !hbusreq3_p & v22f1dc4;
assign v230e689 = hbusreq3 & v23f65eb | !hbusreq3 & v22fe19a;
assign v22ff30c = hgrant3_p & v230741d | !hgrant3_p & v2304f67;
assign v97808c = hbusreq5_p & v150745f | !hbusreq5_p & !v84561b;
assign v22f2286 = hbusreq3_p & v2302812 | !hbusreq3_p & !v84561b;
assign v2309573 = hbusreq6_p & v23101dc | !hbusreq6_p & v84561b;
assign v230385f = hmaster0_p & v2311a61 | !hmaster0_p & !v2392066;
assign v23fc151 = hlock2_p & v191aa68 | !hlock2_p & v191a86f;
assign v23f8e34 = hbusreq3_p & v2305bf7 | !hbusreq3_p & v23fcfcf;
assign v2392095 = hbusreq1_p & v2303f89 | !hbusreq1_p & v22fb5bd;
assign v230dbc9 = hbusreq1_p & v23102bf | !hbusreq1_p & v84561b;
assign v22eb657 = hmaster0_p & v23fce7f | !hmaster0_p & v84561b;
assign v22fd71a = hlock4_p & v23fb6b6 | !hlock4_p & v22eb01f;
assign v230e28d = hbusreq1_p & v12cda15 | !hbusreq1_p & v23fc98a;
assign v22fd6ad = hmaster1_p & v84561b | !hmaster1_p & v22fff51;
assign v22fb89a = hbusreq6 & v22ee0d5 | !hbusreq6 & !v22ff914;
assign v23fbab9 = hbusreq3_p & v22f5388 | !hbusreq3_p & !v84561b;
assign a6b8e0 = hgrant1_p & v231128c | !hgrant1_p & v231160e;
assign v22f0b50 = hmaster2_p & v230aa2c | !hmaster2_p & !v23fbd14;
assign v230f883 = hbusreq3_p & v230437d | !hbusreq3_p & v22f9ebc;
assign v2303c12 = hbusreq5_p & v845636 | !hbusreq5_p & v23f730c;
assign v23fb84f = hbusreq5_p & v23fc19d | !hbusreq5_p & v230ee28;
assign v23fbfca = hbusreq3_p & v230e8a0 | !hbusreq3_p & v960676;
assign v23fbaa7 = hbusreq5 & v22fc8c8 | !hbusreq5 & v84561b;
assign v2305b5a = hmaster1_p & v23fbf8d | !hmaster1_p & v23f7fcb;
assign v230cdfb = hbusreq1 & v2303831 | !hbusreq1 & !v22f0860;
assign v230af38 = hgrant1_p & v230e28d | !hgrant1_p & v23f883a;
assign v2302cce = hbusreq5_p & v23f68d8 | !hbusreq5_p & v22f42b0;
assign v23f5abd = hmaster2_p & v84561b | !hmaster2_p & v22ef5c2;
assign v23fc8a4 = hbusreq1 & v22efae1 | !hbusreq1 & !v23f75db;
assign v230b0c6 = stateG10_5_p & v22f4678 | !stateG10_5_p & v22f878c;
assign v230cfa5 = hlock6_p & v23f4f43 | !hlock6_p & v2313279;
assign v22f824f = hlock0_p & v22f8d80 | !hlock0_p & v22ee9be;
assign v23f4bab = jx0_p & e1d3f0 | !jx0_p & v22f4bcf;
assign v23934ed = jx0_p & v23fcfb1 | !jx0_p & v23f7b9b;
assign v23fce49 = hmaster2_p & v22f79fd | !hmaster2_p & v22f8cb7;
assign v23f7f77 = hbusreq1 & v23f3d14 | !hbusreq1 & v84561b;
assign v22ee024 = hbusreq3 & v2303c07 | !hbusreq3 & v84561b;
assign v22ff205 = jx1_p & v22ec6f1 | !jx1_p & v230892a;
assign v23f9c72 = hbusreq5 & bd74c0 | !hbusreq5 & v23fa2ec;
assign v2307a75 = hmastlock_p & v23fc200 | !hmastlock_p & v84561b;
assign v23055fd = hgrant1_p & v84561b | !hgrant1_p & !v23fbee9;
assign v230e1f3 = hgrant1_p & v84561b | !hgrant1_p & v22fe3f6;
assign v230448f = hbusreq0 & v2303dd7 | !hbusreq0 & v84561b;
assign v23051c4 = hgrant1_p & v845626 | !hgrant1_p & v2301d45;
assign v22f4eeb = hmaster2_p & v2301a75 | !hmaster2_p & v22f1585;
assign v2309b63 = hmaster0_p & v23fbdc0 | !hmaster0_p & !v96c563;
assign v230dd4d = jx0_p & v2303ce0 | !jx0_p & !v23f0bbc;
assign v23fbf00 = hmaster0_p & v23fb845 | !hmaster0_p & !v230786e;
assign e1e5c9 = hmaster1_p & v22f299d | !hmaster1_p & v23fcfe9;
assign v23fc75a = hbusreq6 & v84564d | !hbusreq6 & v22f5218;
assign v23fca3e = hbusreq1_p & v23fc904 | !hbusreq1_p & !v22eb5b3;
assign v23fc1f0 = hbusreq1 & v22f2ed7 | !hbusreq1 & v84561b;
assign v2304415 = hbusreq2 & v23f7d51 | !hbusreq2 & v84561b;
assign v22ff4aa = hmaster2_p & v1b87673 | !hmaster2_p & v22f5696;
assign v22f4284 = hmaster1_p & v22f1969 | !hmaster1_p & v230b5c7;
assign v191b096 = hbusreq5 & v23fd049 | !hbusreq5 & v84561b;
assign v2310e05 = hbusreq3_p & v22ee2b4 | !hbusreq3_p & add85b;
assign v2304fdd = hbusreq4 & v22ee7cf | !hbusreq4 & e1e5c7;
assign v23f7be0 = hmaster2_p & v84561b | !hmaster2_p & !v23fcba7;
assign v230d804 = hbusreq5_p & v2303b17 | !hbusreq5_p & v22f1ae5;
assign v23fd060 = hgrant1_p & a1fba6 | !hgrant1_p & v230f105;
assign v23fb3c7 = hbusreq1_p & v23fb49a | !hbusreq1_p & v230e8d3;
assign v23f4761 = hgrant5_p & v22f1ef6 | !hgrant5_p & !v84561b;
assign v22f443a = hmaster1_p & v191b0f9 | !hmaster1_p & !v22f8aa0;
assign v22ef945 = hgrant0_p & v845622 | !hgrant0_p & v23fcb0b;
assign v23fbab2 = hbusreq2_p & v230a6a7 | !hbusreq2_p & !v84561b;
assign v22f22b2 = hbusreq5_p & v23fc4f8 | !hbusreq5_p & v230f860;
assign v230193c = hmaster0_p & v2310d59 | !hmaster0_p & v230e97b;
assign v22f1e67 = hbusreq3 & v22ef6ce | !hbusreq3 & v230299b;
assign v2312283 = hbusreq2_p & v23fcf46 | !hbusreq2_p & !v23fba6b;
assign v230c93a = hbusreq1 & v22f79fd | !hbusreq1 & v84561b;
assign v22fb1bc = hbusreq5_p & v22fa48c | !hbusreq5_p & v84561b;
assign v2300cd4 = hmaster0_p & v2307061 | !hmaster0_p & v191ae51;
assign v22f6066 = hgrant3_p & v84561b | !hgrant3_p & v22f764d;
assign v23119b0 = hmaster1_p & v22f6fda | !hmaster1_p & v23fc4a2;
assign v22eec56 = jx1_p & v191acb4 | !jx1_p & v23fba1d;
assign v230a87b = hmaster0_p & v23fbdf6 | !hmaster0_p & !v2300362;
assign v2346bd3 = decide_p & v22faf11 | !decide_p & v23fcead;
assign v230a8b2 = hmaster2_p & v23fb565 | !hmaster2_p & v84561b;
assign v22f092f = hmaster2_p & v23fb67c | !hmaster2_p & v23f4b28;
assign v230a4f1 = hmaster2_p & v2304bc1 | !hmaster2_p & v22f2f44;
assign v8963c2 = hbusreq3_p & e1dbd6 | !hbusreq3_p & v22f6e30;
assign v23099c5 = hgrant5_p & v84561b | !hgrant5_p & v22ff469;
assign v2304f11 = hlock3_p & v23fbe5d | !hlock3_p & v23f90b2;
assign v2307aeb = hlock6_p & v22f4a16 | !hlock6_p & v924a36;
assign v231147e = hgrant3_p & v230b38b | !hgrant3_p & v22f2e7b;
assign v2313118 = hready & v84561b | !hready & v23f894b;
assign v22ef1f3 = hgrant3_p & v84562e | !hgrant3_p & v2301e10;
assign v22f6d61 = hgrant3_p & v84562e | !hgrant3_p & v23fccb0;
assign v23fc661 = hlock5_p & v230b504 | !hlock5_p & v2310a40;
assign v23fc58b = hlock3_p & v23f317c | !hlock3_p & !v22ec882;
assign e1dcf1 = hgrant5_p & v22f74f7 | !hgrant5_p & v997ca9;
assign v2308ddf = hbusreq4_p & v2309f3f | !hbusreq4_p & v22f053b;
assign v22f1acb = hbusreq4 & v230b292 | !hbusreq4 & v22f61bb;
assign v23f7968 = hgrant1_p & v22eeb03 | !hgrant1_p & v230b6a4;
assign v22ecc5a = hbusreq4 & v22fbd9a | !hbusreq4 & v845625;
assign v22f60dd = hmaster2_p & v22f3101 | !hmaster2_p & v22f8aba;
assign v23f99ae = hmaster2_p & v23f5be9 | !hmaster2_p & v84561b;
assign v23f3d0b = hbusreq3_p & v22f39d3 | !hbusreq3_p & v23fc957;
assign v2392534 = hbusreq5 & v191a86f | !hbusreq5 & !v84561b;
assign v23f83de = hmaster0_p & v230b8fb | !hmaster0_p & v22ee9d5;
assign v22f5f54 = hbusreq6_p & v23fcba2 | !hbusreq6_p & v239299c;
assign v23fb94b = hmaster0_p & v23fbf49 | !hmaster0_p & v22fedf7;
assign v22f1279 = hbusreq5_p & v23f5af5 | !hbusreq5_p & v23fbc4a;
assign bd5342 = hgrant2_p & v22f2f87 | !hgrant2_p & v2303f9a;
assign v23fbd3e = hbusreq5_p & v230ae19 | !hbusreq5_p & v22f18b1;
assign v23f6575 = hgrant0_p & v2309b0f | !hgrant0_p & v22f3b18;
assign v230d509 = hlock0_p & v2301e20 | !hlock0_p & !v22f6183;
assign v22f70a0 = hbusreq5 & v23f4254 | !hbusreq5 & v84561b;
assign v22eb1f5 = hbusreq2_p & v191a86f | !hbusreq2_p & !v191a879;
assign v230dde6 = hgrant3_p & v22ff67c | !hgrant3_p & v2309c1f;
assign v23fc094 = hgrant1_p & v23fbdef | !hgrant1_p & v23fb7e0;
assign v23fbe6a = hmaster2_p & v22f878c | !hmaster2_p & v12cc2ef;
assign v22fe573 = hmaster2_p & v23f3ccf | !hmaster2_p & v22ed59e;
assign v2303415 = hlock3_p & v230272d | !hlock3_p & v2302179;
assign v23fb1e5 = hgrant1_p & v22f5db6 | !hgrant1_p & !v23090fb;
assign v23fb4a0 = hbusreq3 & v230806a | !hbusreq3 & v23fcd6a;
assign b9c976 = hbusreq3_p & b09503 | !hbusreq3_p & v22f14bf;
assign v23056b2 = hmaster1_p & v23f06c9 | !hmaster1_p & v84561b;
assign v23fa95c = hlock6_p & v22ed7a4 | !hlock6_p & !v1b87732;
assign v22f799b = hbusreq3_p & v23faa5c | !hbusreq3_p & v22f1866;
assign v23f854f = hgrant0_p & v84561b | !hgrant0_p & v22ec2cb;
assign v22f6ba0 = hlock5_p & v22f8271 | !hlock5_p & !v23056b1;
assign v23fc633 = hmaster2_p & v22f8834 | !hmaster2_p & v84561b;
assign v23fc782 = hbusreq5_p & v23fc904 | !hbusreq5_p & !v22ff404;
assign v22fbe82 = hbusreq0_p & v22eefe2 | !hbusreq0_p & v84561b;
assign v22f6b45 = hbusreq1_p & v12cda15 | !hbusreq1_p & v2304bc1;
assign v23fc9a1 = hmaster2_p & v23fc4f9 | !hmaster2_p & v2306e35;
assign v2311476 = hbusreq6_p & v23fc0c3 | !hbusreq6_p & v23fb808;
assign v231065b = hlock4_p & v23fc32a | !hlock4_p & v23f5446;
assign v8b7fb1 = hlock2_p & v845647 | !hlock2_p & !v84561b;
assign v23064ca = hbusreq3 & v22f3be2 | !hbusreq3 & v84561b;
assign v22f4db6 = hbusreq4 & v22f3dc7 | !hbusreq4 & !v23f8e04;
assign v23fc5bf = hlock4_p & v22f606c | !hlock4_p & v23f15e7;
assign v2305660 = hbusreq4_p & v2307dae | !hbusreq4_p & v2308f5d;
assign v22fc88a = hbusreq3_p & v22efa0a | !hbusreq3_p & !v23fc8e4;
assign v22f6d82 = hbusreq3_p & v23fb2d6 | !hbusreq3_p & !v23108db;
assign v230468d = hmaster2_p & v23fc38f | !hmaster2_p & v22f61ac;
assign v23079d8 = hmaster2_p & v22f3618 | !hmaster2_p & v2303b6a;
assign v23f1908 = hmaster1_p & v230f0de | !hmaster1_p & v23fbd21;
assign v22f696f = hbusreq4_p & v23fcccb | !hbusreq4_p & v23fa66e;
assign v22fcf71 = hgrant0_p & v22f824f | !hgrant0_p & v23fb912;
assign v23f43d6 = hbusreq3_p & v22ffe44 | !hbusreq3_p & v22f2f26;
assign v9f5c3c = hmaster2_p & v22f7b47 | !hmaster2_p & v23fc741;
assign v22f73fb = hbusreq6 & v2302783 | !hbusreq6 & !v23fbeeb;
assign v8a7512 = hgrant1_p & v84561b | !hgrant1_p & v23f7898;
assign v230f9b8 = hmaster2_p & v2312231 | !hmaster2_p & v23f8036;
assign v2305e00 = hmaster0_p & v2393abe | !hmaster0_p & v84561b;
assign v230d82a = jx0_p & v2300e6b | !jx0_p & v22fdb07;
assign v23f835c = hbusreq0_p & v84561b | !hbusreq0_p & v230eb9b;
assign v22fb081 = hbusreq3_p & v23fce4e | !hbusreq3_p & v23fc957;
assign v23fcedf = hbusreq3_p & v22f227e | !hbusreq3_p & v23fcbe9;
assign v22f0b56 = hmaster2_p & v22f0add | !hmaster2_p & v22f6741;
assign v230ca7c = hbusreq1 & v2302071 | !hbusreq1 & !v230af81;
assign v23f9370 = hgrant1_p & v230e514 | !hgrant1_p & !v191ad4f;
assign v23fbf3f = hbusreq4 & v23fbe18 | !hbusreq4 & !v150718d;
assign v239300d = hbusreq6_p & v230cfa5 | !hbusreq6_p & v84561b;
assign v22efe2f = hbusreq4 & v22fa9ce | !hbusreq4 & v84561b;
assign v2309ff9 = hlock1_p & v2392d97 | !hlock1_p & v23f66e6;
assign v23fc027 = hmaster2_p & v84561b | !hmaster2_p & v230471d;
assign v23f729b = hmaster2_p & v22ef46e | !hmaster2_p & !v23fbedc;
assign v22f4ace = hbusreq0 & bd9916 | !hbusreq0 & v84561b;
assign v23fc190 = hgrant5_p & v22f05f3 | !hgrant5_p & fc8f72;
assign v23f33b2 = hmaster0_p & v230b8fb | !hmaster0_p & v2302e1b;
assign v22f8001 = hbusreq6_p & v2303b2a | !hbusreq6_p & bf9ce3;
assign v22f2d10 = hmaster0_p & v22ecb5c | !hmaster0_p & v2301392;
assign v23f60d2 = hbusreq3_p & v23fc19b | !hbusreq3_p & v1aae9a1;
assign v2304253 = jx0_p & v23fcc4e | !jx0_p & v22f161f;
assign v23fcd1e = hbusreq5 & v2304009 | !hbusreq5 & v23fb966;
assign v23f49cd = hmaster0_p & v2309499 | !hmaster0_p & v23f9714;
assign v1e841b6 = decide_p & v23fb1d7 | !decide_p & v23fbc7b;
assign v2310a35 = hlock5_p & v22fe627 | !hlock5_p & !v84561b;
assign v230b1ac = hready & v84561b | !hready & !v2302c4b;
assign v22f9cd7 = hbusreq5 & v22fe097 | !hbusreq5 & v84561b;
assign v230a562 = hgrant1_p & v23f4491 | !hgrant1_p & v23fcd33;
assign v2301a75 = hbusreq1_p & v23fcd56 | !hbusreq1_p & v84561b;
assign v23efb3a = hmaster0_p & v23fbffa | !hmaster0_p & !v22eede3;
assign v22f853d = hbusreq3_p & v84561b | !hbusreq3_p & v2305abd;
assign v230c95c = hmaster2_p & v845627 | !hmaster2_p & v2303bc3;
assign v23fc38f = hgrant1_p & v23fb6ff | !hgrant1_p & v2312351;
assign v23fca4b = hmaster0_p & v2300d5f | !hmaster0_p & v23fba06;
assign v22f779a = jx1_p & v12cd570 | !jx1_p & v2300ce0;
assign v22fb2f7 = hlock5_p & v22f8062 | !hlock5_p & v23fc9cb;
assign v2306f2e = hbusreq3 & v23f5dcc | !hbusreq3 & v84561b;
assign v23fb691 = hbusreq5 & v23fc619 | !hbusreq5 & v9f009f;
assign v22fb589 = hmaster2_p & v2312c13 | !hmaster2_p & v22fe497;
assign v22f0a19 = hbusreq3 & v84564d | !hbusreq3 & v2302131;
assign v230129b = hmaster2_p & da38c1 | !hmaster2_p & v84561b;
assign v22f83f2 = hbusreq3_p & v230c749 | !hbusreq3_p & v84561b;
assign v23fbe5d = hbusreq3_p & v23f9319 | !hbusreq3_p & v84561b;
assign v2312f4f = hmaster2_p & v191a86f | !hmaster2_p & v22f35e8;
assign v22efcd6 = hlock0_p & v23f69ba | !hlock0_p & v84561b;
assign v23fbd75 = hbusreq6 & v22fdbd2 | !hbusreq6 & v230988d;
assign v230466d = hbusreq5_p & v22f1ece | !hbusreq5_p & !v84561b;
assign v23fcfe9 = hbusreq4_p & v22efcee | !hbusreq4_p & v23fc0c7;
assign v23fbc0c = hmaster0_p & v84561b | !hmaster0_p & v22f2c87;
assign v23fca7e = hbusreq3_p & v22f6a3a | !hbusreq3_p & v23fba18;
assign bdac8b = jx1_p & v23071f4 | !jx1_p & v22efbe2;
assign v23fce65 = stateG2_p & v84561b | !stateG2_p & !v23f2216;
assign v22ec29a = locked_p & v22fef4f | !locked_p & v10dbf64;
assign v231354e = hmaster2_p & v22f426a | !hmaster2_p & v23fb9fe;
assign v23fca1b = hmaster0_p & v22f81ba | !hmaster0_p & !v23fc20d;
assign v23fbe7f = hbusreq3_p & v22f909b | !hbusreq3_p & v23f660f;
assign v2304922 = hbusreq1_p & v22f2db0 | !hbusreq1_p & v1aae98c;
assign v239254b = hgrant0_p & v22fe0f9 | !hgrant0_p & v23fceb9;
assign v23fbe91 = hbusreq3 & v2308c76 | !hbusreq3 & v84561b;
assign v22ff0de = hbusreq4_p & v2302e7b | !hbusreq4_p & !v23fc061;
assign v22ed645 = hbusreq4_p & v22f525a | !hbusreq4_p & v23f20e8;
assign v23f5ae4 = hbusreq3 & v23fbe1c | !hbusreq3 & v23f87f4;
assign v22f7303 = hmaster0_p & v22f5b7c | !hmaster0_p & v22f09c4;
assign v23110b9 = hbusreq0 & v22f60c6 | !hbusreq0 & !v2391a57;
assign v8ebd5d = hbusreq5 & v22fe73f | !hbusreq5 & v84561b;
assign v22ed42c = hgrant6_p & v2304744 | !hgrant6_p & v231353a;
assign v23fced3 = jx1_p & v85e5cf | !jx1_p & v84561b;
assign v1e840fd = hmaster0_p & v23fca89 | !hmaster0_p & !v23fb201;
assign v230629d = hmaster0_p & v2312680 | !hmaster0_p & v22eb952;
assign v230c439 = hmaster0_p & v23fb6d7 | !hmaster0_p & v23f5382;
assign v23fc6c0 = hgrant1_p & v230031f | !hgrant1_p & v22f2a60;
assign v22f979e = hbusreq6_p & v2312248 | !hbusreq6_p & v23fc04e;
assign v23fb95d = hmastlock_p & v23f7326 | !hmastlock_p & v84561b;
assign v230b91d = hgrant2_p & v23f5af5 | !hgrant2_p & v2308a30;
assign v23faf60 = hgrant0_p & v845622 | !hgrant0_p & v23fc1e3;
assign v23f6fa8 = hmaster2_p & v22fdc30 | !hmaster2_p & v23fccbe;
assign v22ebe20 = hmaster0_p & v22f97c3 | !hmaster0_p & v23fbc9f;
assign v2303e13 = hbusreq5 & v191a876 | !hbusreq5 & v84561b;
assign v22f8593 = hbusreq1_p & v22fead6 | !hbusreq1_p & v23f909e;
assign v22fbb8a = hgrant2_p & v23066df | !hgrant2_p & fc8ab7;
assign v23013f8 = hbusreq4_p & v22f41c4 | !hbusreq4_p & v230fe6b;
assign v2303513 = hbusreq4 & v22ee8bf | !hbusreq4 & v23fc51e;
assign v2306854 = jx2_p & v191b1a1 | !jx2_p & v23f7073;
assign v23fb0ce = hgrant1_p & a1fba6 | !hgrant1_p & v23fcba5;
assign v230cdc1 = hbusreq6 & v2300d93 | !hbusreq6 & v23f3297;
assign v230b77e = hmaster0_p & v22fcdd3 | !hmaster0_p & !v23fc541;
assign v23fcfb7 = hgrant5_p & v23fca15 | !hgrant5_p & v22fe73f;
assign v23f9ca2 = hgrant2_p & v23fb9ff | !hgrant2_p & !v84561b;
assign v22ffc31 = hbusreq4_p & v2306d2c | !hbusreq4_p & v23f347b;
assign v22fa69c = hbusreq4_p & v22f8556 | !hbusreq4_p & v22f35fd;
assign v230f760 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v23f11a3;
assign v230a36f = hbusreq6_p & v230a5f5 | !hbusreq6_p & v22f53b1;
assign v23fc753 = hbusreq3_p & v22ed5c8 | !hbusreq3_p & v231051e;
assign v1aadb8e = locked_p & v22f334e | !locked_p & v13afe8f;
assign v1aad518 = hlock0_p & v230e4ef | !hlock0_p & v84561b;
assign v23fcb9a = hgrant5_p & v22f6cc8 | !hgrant5_p & v23fc2a5;
assign v22ece0e = hmaster0_p & v22f4c34 | !hmaster0_p & v23fbdec;
assign v23fc6af = hmaster0_p & v2310319 | !hmaster0_p & v22fec34;
assign v23039fa = hbusreq4_p & v9ae938 | !hbusreq4_p & v22fc4af;
assign v23fce06 = hbusreq4_p & v1e84b3d | !hbusreq4_p & v22fb062;
assign v2302da4 = hgrant3_p & v22f3628 | !hgrant3_p & v230c3f5;
assign v22f4bb5 = hlock1_p & v22f5d87 | !hlock1_p & v845620;
assign a0de1c = hbusreq3 & v22f7e19 | !hbusreq3 & v84561b;
assign v2306e27 = hbusreq5_p & v230320e | !hbusreq5_p & !v23012e5;
assign fc88ba = hmaster2_p & v22f9911 | !hmaster2_p & v23fb9c2;
assign v22eaf27 = jx0_p & v22ec240 | !jx0_p & v23fb13c;
assign v22ef78e = hmaster1_p & v230499e | !hmaster1_p & v230ea78;
assign v23fcad4 = hbusreq0 & v84561b | !hbusreq0 & fc8ab7;
assign b9c9d4 = hbusreq3 & v1aad31f | !hbusreq3 & v84561b;
assign v2301d23 = hlock1_p & v23f2b14 | !hlock1_p & v2309c93;
assign v23f717f = hgrant1_p & b50a75 | !hgrant1_p & v23108a7;
assign v23fc2ba = hbusreq5_p & v22f56d2 | !hbusreq5_p & v22f18b4;
assign v2307fd0 = hgrant3_p & v13afe72 | !hgrant3_p & baa026;
assign v230042c = hbusreq3_p & v2304be0 | !hbusreq3_p & !v84561b;
assign v23056e9 = hgrant2_p & v22fdc30 | !hgrant2_p & v22f9980;
assign v23fc9ef = hgrant5_p & v23fc583 | !hgrant5_p & v23fc356;
assign v22ec6f1 = hmaster1_p & v23103f8 | !hmaster1_p & v23fccd3;
assign v22f6dee = hgrant3_p & baf3e5 | !hgrant3_p & v23f447e;
assign v23fa2eb = hbusreq3 & v22fbd9a | !hbusreq3 & v845625;
assign v22f099c = hbusreq2 & v23fb9ac | !hbusreq2 & v23f59e0;
assign v23007a4 = hlock1_p & v23f5af5 | !hlock1_p & !v2309c8a;
assign v230aa17 = hgrant3_p & v84561b | !hgrant3_p & v22fba6d;
assign v230d25c = hbusreq5_p & v22f34d8 | !hbusreq5_p & !v84561b;
assign v22fca75 = hbusreq5_p & v22fd311 | !hbusreq5_p & !v84561b;
assign v22fc19c = hbusreq0 & v23f65b4 | !hbusreq0 & v84561b;
assign v23fbd7e = hbusreq3_p & v22ff21b | !hbusreq3_p & !v23fc92f;
assign v2311559 = hmaster2_p & v2311810 | !hmaster2_p & a1fbc2;
assign v2300503 = hbusreq4 & v23053fb | !hbusreq4 & v84561b;
assign f40c9d = hbusreq5_p & v22f3a35 | !hbusreq5_p & v22ebd62;
assign v23fb544 = hbusreq4_p & v9cf5cf | !hbusreq4_p & v22ff80d;
assign v23fc3f1 = hgrant1_p & v23fbc94 | !hgrant1_p & v84561b;
assign v22f595f = hlock0_p & v1506a9e | !hlock0_p & !v230e40a;
assign v22ed4ea = hmaster1_p & v23073e6 | !hmaster1_p & v231396f;
assign v22fea74 = hmaster2_p & v23f3206 | !hmaster2_p & v85f4fd;
assign v23f7ea0 = hbusreq5 & v22f98e3 | !hbusreq5 & v23fc3f2;
assign v23f5be9 = hlock0_p & v84561b | !hlock0_p & v23fba70;
assign v22fa594 = hbusreq5 & v22fc5f0 | !hbusreq5 & v22f5583;
assign v22f2653 = stateG10_5_p & v23fcffa | !stateG10_5_p & v22ee956;
assign v230aba5 = hbusreq5_p & v230f63f | !hbusreq5_p & v22f42c9;
assign v230eac0 = hbusreq3_p & v23fc5e9 | !hbusreq3_p & v23fba73;
assign v22f0768 = hlock6_p & v2309add | !hlock6_p & v22f990d;
assign v22fbc05 = hbusreq1 & v22ed6c5 | !hbusreq1 & v84564d;
assign v2306220 = hmastlock_p & v230fdc7 | !hmastlock_p & v84561b;
assign v230cd1c = hmaster1_p & v22f8f5f | !hmaster1_p & v23f85b5;
assign v22ec71a = hgrant1_p & v230abce | !hgrant1_p & v22fdb01;
assign v23027b1 = hbusreq6 & v22f7fcc | !hbusreq6 & v22f1a8f;
assign v22ee03c = hbusreq3 & v230f863 | !hbusreq3 & v84561b;
assign v22ed346 = hgrant2_p & v106a782 | !hgrant2_p & v23f354c;
assign c0aa95 = hmaster2_p & v23fcb55 | !hmaster2_p & v2310754;
assign v2309d55 = hbusreq1_p & v84562a | !hbusreq1_p & v230af81;
assign v22f46d3 = hbusreq3_p & v230d291 | !hbusreq3_p & bd9c35;
assign v1e840d4 = hbusreq3_p & v15072a9 | !hbusreq3_p & v23fcdbe;
assign v191aa89 = hgrant1_p & v22f54a4 | !hgrant1_p & v23f1e1a;
assign v23fcfb1 = jx1_p & v23f5d39 | !jx1_p & v23070ef;
assign v23f99bc = hgrant3_p & v23fba39 | !hgrant3_p & v2302a77;
assign v23fb732 = jx2_p & v23fc7b5 | !jx2_p & v84561b;
assign v230c155 = hbusreq6_p & v2309856 | !hbusreq6_p & v23f18fc;
assign v23fc511 = hbusreq1_p & v23fc31a | !hbusreq1_p & v84561b;
assign v23f496d = hlock6_p & a0f5d5 | !hlock6_p & v22fabad;
assign v23f368a = hbusreq1_p & v22f2f44 | !hbusreq1_p & v23f6038;
assign v2311e58 = hgrant4_p & v23fbeec | !hgrant4_p & v22eef3b;
assign v22f950e = hbusreq5_p & v845636 | !hbusreq5_p & v23fb5d0;
assign v23f9a5b = hbusreq3_p & v23f5ae4 | !hbusreq3_p & !v2309eab;
assign v23f46d8 = hlock4_p & v23fcf44 | !hlock4_p & v22f7b49;
assign v23f2df5 = hbusreq6 & v23fbcad | !hbusreq6 & !v230e860;
assign v22fead6 = hbusreq1 & v22fda32 | !hbusreq1 & v23fa2ec;
assign v2308748 = hgrant5_p & v23f65b6 | !hgrant5_p & v84561b;
assign v22f97e9 = stateG2_p & v84561b | !stateG2_p & v23f71c9;
assign v22fe7b0 = hmaster2_p & v23fba9a | !hmaster2_p & v231025b;
assign v230a84b = hbusreq3_p & v22f575a | !hbusreq3_p & v23f56bc;
assign v23fc49c = hbusreq4_p & v23fbbaa | !hbusreq4_p & !v84561b;
assign v22f903f = hmaster2_p & v23fc9d1 | !hmaster2_p & v23f328e;
assign v23fb1a6 = hgrant2_p & v12cd523 | !hgrant2_p & !v1aae98c;
assign v2392898 = hlock4_p & v23fbf0a | !hlock4_p & v23fd038;
assign v22f7fc1 = hbusreq6_p & v2306cca | !hbusreq6_p & !v84561b;
assign v23fac6d = hbusreq3_p & v22ed598 | !hbusreq3_p & v22f0dc3;
assign v22eca65 = hgrant3_p & v23035ba | !hgrant3_p & v23fb90f;
assign v23fb0f3 = hmaster0_p & v23f48a1 | !hmaster0_p & v22fc5a9;
assign v1507157 = hbusreq3 & v2305a94 | !hbusreq3 & v23fbd9c;
assign v23f67fe = hbusreq3_p & v22f1e46 | !hbusreq3_p & v84561b;
assign v23f1f36 = hlock6_p & v84561b | !hlock6_p & v23f6532;
assign v22f3832 = hmaster0_p & v22f8cb9 | !hmaster0_p & v23fcaf6;
assign v22fdf70 = hlock4_p & v2310bd4 | !hlock4_p & v23f2d60;
assign v23059d8 = hbusreq0 & v22f2718 | !hbusreq0 & v84561b;
assign v23fbced = jx1_p & v2301a7e | !jx1_p & v22ef38d;
assign v22f4e77 = hbusreq1 & v22fd699 | !hbusreq1 & v2305ebc;
assign v23fbaac = hbusreq1_p & v23f2b6d | !hbusreq1_p & v22f878c;
assign v22f9dab = hmaster0_p & v22fc903 | !hmaster0_p & v23fbc3a;
assign v230786e = hbusreq6 & v22f0545 | !hbusreq6 & !v84561b;
assign v22f6056 = stateG10_5_p & v22ec6e7 | !stateG10_5_p & !v2393f17;
assign v230025c = hbusreq4_p & v23fbbeb | !hbusreq4_p & bda6cc;
assign v23fcb64 = hgrant3_p & v22f8309 | !hgrant3_p & v22f8093;
assign v2306d07 = hbusreq2 & v22f1a26 | !hbusreq2 & v84561b;
assign v230f6d0 = hgrant6_p & v230a9ca | !hgrant6_p & v2312dfa;
assign af7272 = hmaster2_p & v22f86f3 | !hmaster2_p & v23f3d47;
assign v23928d0 = hbusreq6 & v23f31d6 | !hbusreq6 & v12ce0d0;
assign v23f4462 = hgrant2_p & v22f8f0b | !hgrant2_p & !v84561b;
assign v22f7e16 = hready & v22fc63c | !hready & !v84561b;
assign v23fc4f4 = hbusreq6_p & v23fca59 | !hbusreq6_p & v230994d;
assign v22f5eee = locked_p & v2306667 | !locked_p & v84561b;
assign v230ab2e = hlock3_p & v23f35ff | !hlock3_p & !v84561b;
assign v2304910 = hbusreq2 & v22f0f15 | !hbusreq2 & v84561b;
assign v2309dc4 = hgrant1_p & v12cc2ef | !hgrant1_p & v22f419a;
assign v22ff7d0 = hbusreq0 & v84561b | !hbusreq0 & v2304ec7;
assign v2310c6d = hbusreq5_p & v230aef0 | !hbusreq5_p & !v84561b;
assign v23125fb = hlock3_p & v22fc8e1 | !hlock3_p & !v106ae19;
assign v23fbf2c = hbusreq1_p & v230a951 | !hbusreq1_p & !v230ef5b;
assign v22fca4e = hgrant0_p & v84561b | !hgrant0_p & v23039be;
assign v22ef683 = hgrant0_p & v845620 | !hgrant0_p & v23fcdd5;
assign v230a579 = hbusreq3 & bdf576 | !hbusreq3 & !bafb17;
assign v22ee59c = hbusreq2 & v845620 | !hbusreq2 & v84561b;
assign v2303e0d = hmaster0_p & v23fcb64 | !hmaster0_p & v22ebc60;
assign v22eb771 = hbusreq5_p & v23fc5f4 | !hbusreq5_p & v23fbf2a;
assign v22ef2b4 = hmaster2_p & v23fb7fc | !hmaster2_p & v22f389b;
assign v23fb652 = hbusreq4_p & v23f4b8f | !hbusreq4_p & v22fe4f6;
assign v230d9d9 = hbusreq5_p & v23f9c72 | !hbusreq5_p & v2308b6b;
assign b0fe84 = hbusreq3_p & v2300487 | !hbusreq3_p & v23fbc83;
assign v2302d56 = hmaster0_p & v23f1afd | !hmaster0_p & v23fcfa5;
assign bd74c0 = hbusreq2_p & v23fcd73 | !hbusreq2_p & v84561b;
assign v23f9c5f = hmaster2_p & v84561b | !hmaster2_p & v2302048;
assign v22f1cb7 = hbusreq1_p & v23fcd39 | !hbusreq1_p & v845620;
assign bd7a67 = hbusreq3 & v22ee0d6 | !hbusreq3 & v2312f81;
assign v22f8387 = hgrant5_p & v230f453 | !hgrant5_p & v22ecf87;
assign v23fb1c1 = hgrant1_p & v22fb1bc | !hgrant1_p & v23fbacf;
assign v23fcaff = hmaster2_p & v2391b6f | !hmaster2_p & v230c69b;
assign v23fc006 = hbusreq4_p & v23fcec4 | !hbusreq4_p & v23fc83e;
assign v23f7031 = hbusreq5_p & v23f988f | !hbusreq5_p & v2311891;
assign bda69e = hmaster2_p & v22f26fc | !hmaster2_p & v23f8d76;
assign v23fb9f8 = hbusreq5_p & v23fcf91 | !hbusreq5_p & v230186e;
assign v230d04a = stateG2_p & v84561b | !stateG2_p & a1ff27;
assign v1aad4b2 = hbusreq5 & v22f84ff | !hbusreq5 & !v84561b;
assign v23fbd11 = hmaster0_p & v2392254 | !hmaster0_p & v230f27a;
assign v22f0284 = hmaster0_p & v22eec11 | !hmaster0_p & v23f3b81;
assign v230efb1 = stateA1_p & v84561b | !stateA1_p & v845649;
assign v23fc3e8 = hmaster2_p & v22f7aff | !hmaster2_p & v23fc757;
assign v8bbb53 = hmaster2_p & v23fb1c1 | !hmaster2_p & v22f5815;
assign a84b89 = hlock0_p & v230f2d6 | !hlock0_p & !v84561b;
assign v230f03c = hmaster0_p & v22f8e29 | !hmaster0_p & v23105aa;
assign v230236f = hbusreq6_p & v23fbf7f | !hbusreq6_p & v23f8e1c;
assign v23934f3 = hmaster2_p & v22f4d20 | !hmaster2_p & v23f717f;
assign v239353f = hbusreq3 & v2305f8e | !hbusreq3 & !v845622;
assign v2307480 = hbusreq4_p & v22eb701 | !hbusreq4_p & v2367a5a;
assign v23fce3a = hmaster2_p & v22f13e3 | !hmaster2_p & v23f4c8c;
assign v22eed1b = hmaster2_p & v23fbe41 | !hmaster2_p & v22f037a;
assign v23fb196 = hmaster1_p & v22eb15f | !hmaster1_p & v22ee36e;
assign v2305345 = hmaster2_p & v22f61b6 | !hmaster2_p & v2311be9;
assign v22ff463 = hbusreq5_p & v2306d29 | !hbusreq5_p & v22ec0d4;
assign v23fc88b = hmaster2_p & v22f6358 | !hmaster2_p & v84561b;
assign v22ee957 = hmaster2_p & v22fc8c8 | !hmaster2_p & v23fcb5b;
assign v23fbff6 = hmaster2_p & v2312f7e | !hmaster2_p & v22fdc17;
assign v2306d36 = hgrant4_p & v84561b | !hgrant4_p & v23f3ab8;
assign v23060e3 = hmaster2_p & v22fc13d | !hmaster2_p & v22fa700;
assign v22f88bb = hgrant3_p & v84561b | !hgrant3_p & v2313131;
assign v230d2a3 = hbusreq6 & v23f82e4 | !hbusreq6 & v23fcaab;
assign v23fc31a = hlock1_p & v84561b | !hlock1_p & v23f301a;
assign v2300edd = hburst1 & v22f3294 | !hburst1 & v23f16f6;
assign v22f1ee5 = hready & v23fb95d | !hready & v22f197e;
assign v22f33e0 = hmaster2_p & v23112ad | !hmaster2_p & v22ec894;
assign v22f03ec = hbusreq6_p & v22f9d79 | !hbusreq6_p & v22fa65d;
assign v2307dfb = hbusreq3_p & v23fc19b | !hbusreq3_p & v23f6db4;
assign v23fc438 = hbusreq6_p & v23f1a4c | !hbusreq6_p & v22ff650;
assign v23f0699 = hbusreq0_p & v23fca48 | !hbusreq0_p & v845622;
assign v22fa474 = hbusreq1 & v106ae21 | !hbusreq1 & v84564d;
assign v22eebf5 = hmaster2_p & v84564d | !hmaster2_p & !v2391a57;
assign v2304db3 = hbusreq5_p & v845636 | !hbusreq5_p & bd7bf6;
assign v23f3545 = hmaster2_p & v84561b | !hmaster2_p & v23f468c;
assign bd8367 = hbusreq3_p & v22f2d7c | !hbusreq3_p & v22fede6;
assign v13aff51 = hlock3_p & v2309e9d | !hlock3_p & !v84561b;
assign v230590b = hgrant1_p & v84561b | !hgrant1_p & v23f7f0d;
assign v23f645e = hbusreq6_p & v84564d | !hbusreq6_p & v22f4f0f;
assign v22f8477 = hmaster2_p & v23fc63b | !hmaster2_p & v22f61b6;
assign v230bc8b = hgrant0_p & v84564d | !hgrant0_p & v23fc926;
assign v23f7a5f = hbusreq0 & v2302048 | !hbusreq0 & v84561b;
assign v230de87 = hmaster0_p & v230a9a3 | !hmaster0_p & v230d45f;
assign v22ec644 = hmaster0_p & v22ec77a | !hmaster0_p & v23fb924;
assign v22f1b18 = hgrant3_p & d49f2b | !hgrant3_p & v23fbca1;
assign v23fbc95 = jx1_p & v23f3d09 | !jx1_p & v22fc481;
assign v23fbb85 = jx1_p & v22f5429 | !jx1_p & v22f2b34;
assign v12cd9f9 = hbusreq1_p & v84564d | !hbusreq1_p & !v84561b;
assign v23fcedd = hgrant0_p & v23133fa | !hgrant0_p & v22f446e;
assign v22f4f19 = hmaster2_p & v22fd0e6 | !hmaster2_p & v22ee8f3;
assign v2309e8e = hmaster2_p & v23084c9 | !hmaster2_p & !v84561b;
assign v22f5944 = jx1_p & v23fc08c | !jx1_p & v230b9f3;
assign v230b95f = hbusreq5_p & v22f5fa1 | !hbusreq5_p & v230a42d;
assign v23fb481 = locked_p & v23fbfaf | !locked_p & v23fc8be;
assign v2311491 = hgrant4_p & v230a8eb | !hgrant4_p & v22fb31a;
assign v22f94c1 = jx1_p & v85e5cf | !jx1_p & f406a3;
assign v9122cc = hgrant3_p & v84561b | !hgrant3_p & !v23fb5cf;
assign v15071ed = hlock4_p & v23f5e84 | !hlock4_p & v23f7393;
assign v230254a = stateG10_5_p & v22ed49b | !stateG10_5_p & v23fbc42;
assign v17a34ea = hbusreq1_p & v230b09e | !hbusreq1_p & v84561b;
assign v2300359 = jx1_p & v23049cc | !jx1_p & v230892a;
assign v230d64e = hbusreq1_p & v23fcc8e | !hbusreq1_p & v2305128;
assign v22fd655 = hlock0_p & v2308455 | !hlock0_p & v22f1e0b;
assign v22ebb82 = hgrant3_p & v84562e | !hgrant3_p & v2301c57;
assign v23fcd05 = stateG10_5_p & v22edeb5 | !stateG10_5_p & v22fc430;
assign hmaster0 = !v214cf31;
assign v2312248 = hmaster0_p & v230f6e9 | !hmaster0_p & v84561b;
assign v22efc9e = hmaster2_p & v2306d29 | !hmaster2_p & v22fe426;
assign v22ec60b = hbusreq6_p & v8958ff | !hbusreq6_p & v23fcbaf;
assign v230ad0e = hmaster1_p & v23f96b7 | !hmaster1_p & v23f4168;
assign v22fd311 = hbusreq5 & v23fc514 | !hbusreq5 & !v22f91c9;
assign v23fc1c6 = hmaster2_p & v13afb18 | !hmaster2_p & v230c025;
assign v22f6629 = hbusreq3_p & c20101 | !hbusreq3_p & v23f3e38;
assign v2391d2f = hgrant3_p & v84561b | !hgrant3_p & v230545b;
assign bda6a0 = hbusreq0 & v2392ea0 | !hbusreq0 & v23f2ecd;
assign v23fca8a = jx1_p & v84561b | !jx1_p & v230ed31;
assign v23f0652 = hlock0_p & v230af3a | !hlock0_p & v23fcca4;
assign v2312dc5 = hbusreq4_p & v23f8f18 | !hbusreq4_p & v22f884c;
assign v22fe4ea = hgrant3_p & v230290f | !hgrant3_p & v23f7a18;
assign v23f522c = hmaster2_p & v84564d | !hmaster2_p & v84561b;
assign v23044e1 = hmaster0_p & v230ed7d | !hmaster0_p & v2312a93;
assign v22fa6b2 = hmaster2_p & v84561b | !hmaster2_p & !v230cbdd;
assign v2305d89 = hbusreq3_p & v2308d5a | !hbusreq3_p & v22fa5f9;
assign v23fcf17 = hbusreq3_p & v23fbca0 | !hbusreq3_p & v230e9ef;
assign v2308dd1 = hlock3_p & v23fc873 | !hlock3_p & v23fcf9c;
assign a1fd70 = hmaster1_p & v23fc16f | !hmaster1_p & v23fba19;
assign v23fca10 = hgrant3_p & v84562e | !hgrant3_p & v231025b;
assign v23fc3cb = hgrant0_p & a1fbc2 | !hgrant0_p & v22eed66;
assign v23f4ab8 = hbusreq0 & v23fc842 | !hbusreq0 & v84561b;
assign v23fc04e = hmaster0_p & v23fba11 | !hmaster0_p & v84561b;
assign v23fb47c = hbusreq0 & v23f6b25 | !hbusreq0 & v84561b;
assign v22f55fa = hbusreq1_p & v230916d | !hbusreq1_p & v22ee9be;
assign v22fb0ac = hbusreq4_p & v23f1824 | !hbusreq4_p & v23f165d;
assign v22f87bf = hmaster0_p & v84561b | !hmaster0_p & !v22fc90d;
assign v22fc2eb = hbusreq2_p & v23fce8d | !hbusreq2_p & !v84561b;
assign v2303d00 = hbusreq1_p & v230e6ba | !hbusreq1_p & v23fba97;
assign v22fd079 = hbusreq4_p & v2304d59 | !hbusreq4_p & v23fc888;
assign v22facbb = hbusreq5_p & v230e07d | !hbusreq5_p & v23f9f68;
assign v23fb8e5 = hgrant3_p & v84561b | !hgrant3_p & v2391b6c;
assign v22ec9b2 = hbusreq3_p & v22f909b | !hbusreq3_p & v22f61b6;
assign v23fc5cd = hbusreq1_p & v22f7ad6 | !hbusreq1_p & !v84561b;
assign v23fb1c3 = hbusreq4 & v23fbe4f | !hbusreq4 & v84561b;
assign v85d110 = hlock0_p & v22f8d80 | !hlock0_p & v1507161;
assign a1fe52 = hbusreq5_p & v22ffbb3 | !hbusreq5_p & v2304a64;
assign v23fc366 = hbusreq4 & v22fc8fb | !hbusreq4 & v84561b;
assign v22ee60e = hbusreq6_p & v23fbd11 | !hbusreq6_p & v23f965c;
assign v23fcbab = hbusreq5_p & v23fcf46 | !hbusreq5_p & v9bf2ce;
assign v23fb5a4 = hmaster2_p & v2301511 | !hmaster2_p & v2309c28;
assign v23fcb0f = hbusreq5_p & v23fba98 | !hbusreq5_p & v2312e57;
assign v23060bb = hbusreq6 & v22f8ed1 | !hbusreq6 & v23fcd6c;
assign v230681b = hbusreq3 & v2300dab | !hbusreq3 & !v22f7e7a;
assign v23fb1b5 = hgrant3_p & v84561b | !hgrant3_p & v23fb073;
assign v22f2a4f = hgrant1_p & v84561b | !hgrant1_p & v23f35d5;
assign v23f7564 = hmaster0_p & v23fcf07 | !hmaster0_p & !v22ef8a9;
assign v23fb8f1 = hbusreq4 & v230bf9f | !hbusreq4 & v84561b;
assign f4066f = hmaster2_p & v22f958d | !hmaster2_p & v2313564;
assign v23034e5 = hbusreq3_p & v230930b | !hbusreq3_p & v84561b;
assign v2303d65 = hbusreq3_p & v84571e | !hbusreq3_p & v84561b;
assign b79a15 = jx0_p & v22f65c9 | !jx0_p & v23085c5;
assign v23f2704 = hbusreq3 & v23efbfd | !hbusreq3 & v23f5eba;
assign v22ffe44 = hmaster2_p & v22f64b2 | !hmaster2_p & v22fe497;
assign v2303051 = hbusreq4_p & v22edc14 | !hbusreq4_p & v22ff259;
assign v23f4694 = locked_p & v84561b | !locked_p & !v22f532c;
assign v2303bee = hbusreq3_p & v22f5405 | !hbusreq3_p & v23fc4f8;
assign v22f4a16 = hbusreq4_p & v2311756 | !hbusreq4_p & v230cb53;
assign v22fc531 = hbusreq4_p & v2307081 | !hbusreq4_p & v23fb946;
assign v23fc920 = hbusreq5 & v23fa63b | !hbusreq5 & !v23f3978;
assign v22f814e = hbusreq6_p & v22fb87a | !hbusreq6_p & v22f7d67;
assign v22fefde = hbusreq6_p & v2311b9e | !hbusreq6_p & v23fcb75;
assign v23fba09 = hbusreq5 & v23f34d4 | !hbusreq5 & v84561b;
assign v2306bb2 = hgrant0_p & b094ff | !hgrant0_p & !v84561b;
assign v23fb657 = hbusreq4_p & v23fcec4 | !hbusreq4_p & v84561b;
assign v230cc70 = jx1_p & v23fc8b8 | !jx1_p & v22fca1d;
assign v23074c9 = hbusreq3 & v12cd4c5 | !hbusreq3 & v84561b;
assign v230f099 = hgrant3_p & v17a34ff | !hgrant3_p & v22f5204;
assign v23fc522 = hbusreq6 & v2300503 | !hbusreq6 & v84561b;
assign v23f3bcb = hbusreq3_p & adc67b | !hbusreq3_p & v2304f67;
assign v23fc0e7 = hbusreq6_p & a9176f | !hbusreq6_p & v23007de;
assign v22f5355 = hmaster2_p & v22ec71a | !hmaster2_p & bd9ab5;
assign v2307750 = hbusreq2 & v22fafaa | !hbusreq2 & v84561b;
assign v15070f7 = hbusreq5 & v22fa002 | !hbusreq5 & v84561b;
assign v22fb7e2 = hbusreq4_p & v22ff789 | !hbusreq4_p & v922c74;
assign v22fb744 = hbusreq3 & v22f2cf1 | !hbusreq3 & v23fbd0d;
assign v22f4e9f = hmaster0_p & v22ed9a9 | !hmaster0_p & v23fcb3b;
assign v22fa707 = hgrant0_p & v22f3643 | !hgrant0_p & v23fcd1b;
assign v22f9690 = hbusreq5_p & bbc337 | !hbusreq5_p & v2309126;
assign v230b3a5 = hgrant5_p & v84561b | !hgrant5_p & v845635;
assign v22ebd80 = hready_p & v22ee913 | !hready_p & v845647;
assign v23111c7 = hgrant3_p & v22f4016 | !hgrant3_p & !v2303634;
assign v23f98a9 = hlock4_p & v23fb63e | !hlock4_p & v23fc3ac;
assign v22fda8c = hgrant3_p & v22fee58 | !hgrant3_p & v230788d;
assign v845663 = stateG3_0_p & v84561b | !stateG3_0_p & !v84561b;
assign bd785e = decide_p & v22fb638 | !decide_p & bd76c5;
assign v23f8a89 = hmaster0_p & v23007c9 | !hmaster0_p & v22f8eb8;
assign v23f6849 = hbusreq3_p & v230ed6b | !hbusreq3_p & v84561b;
assign v22f17ca = hbusreq1_p & v238c168 | !hbusreq1_p & v84561b;
assign v2302c68 = hbusreq3_p & v23fb04e | !hbusreq3_p & v23fc0e4;
assign v22ff914 = hbusreq3_p & v84562a | !hbusreq3_p & v2309d55;
assign v22f0c5f = hmaster1_p & v23f416b | !hmaster1_p & v9a3d0c;
assign v230a092 = hmaster0_p & v23fbf3e | !hmaster0_p & v22ed8b5;
assign v22ee2bb = hbusreq0 & v22f68fe | !hbusreq0 & v84561b;
assign v23fcc90 = hgrant3_p & v23f32db | !hgrant3_p & v22f5355;
assign v23129c2 = hbusreq4_p & da310c | !hbusreq4_p & v230629d;
assign v23fb5cf = hmaster2_p & v22fe920 | !hmaster2_p & v230d533;
assign v2302783 = hbusreq3_p & v2307f2b | !hbusreq3_p & v23025d8;
assign v22f09fe = hgrant3_p & v230b199 | !hgrant3_p & bd8367;
assign v2300995 = hmaster0_p & v23fb7c3 | !hmaster0_p & v23f39e6;
assign v22fdaa1 = hlock2_p & v22f8d74 | !hlock2_p & v23fb581;
assign v2312ec4 = hmaster2_p & v23f1228 | !hmaster2_p & v230f046;
assign v23fa600 = hmaster2_p & v2303539 | !hmaster2_p & !v22f70d2;
assign v2307419 = hgrant3_p & v84561b | !hgrant3_p & v84562d;
assign jx3 = !b910da;
assign v22f14ff = hgrant3_p & v84562e | !hgrant3_p & v2311a34;
assign v23915d8 = hbusreq1 & v230a3af | !hbusreq1 & v22f8ad4;
assign v22edff5 = hmaster2_p & v230fc56 | !hmaster2_p & !v12cc2ef;
assign v2303fec = hbusreq4 & v23f70cf | !hbusreq4 & v23fbeeb;
assign v22f4bca = stateG10_5_p & v84561b | !stateG10_5_p & v23f1ca8;
assign v1aae222 = hgrant3_p & v22f8f56 | !hgrant3_p & v22eb3fc;
assign v2308e64 = hmaster2_p & v22ffc69 | !hmaster2_p & !v2309871;
assign v23f0a0b = stateG10_5_p & v23f1d8b | !stateG10_5_p & v22fd25c;
assign v23f5fe3 = hmaster0_p & v2312f45 | !hmaster0_p & v23fac09;
assign v22f2852 = hlock6_p & v191a8f7 | !hlock6_p & v230996e;
assign v23fc335 = hbusreq3_p & v22ed4b7 | !hbusreq3_p & v2308d20;
assign bd7c1c = hbusreq1_p & b3865a | !hbusreq1_p & !v106ae19;
assign v22ece6c = hbusreq1 & v22eb742 | !hbusreq1 & v84561b;
assign v22f8c84 = hbusreq6_p & v2307add | !hbusreq6_p & v22f4ba1;
assign v2392f25 = hbusreq4 & v23f74bf | !hbusreq4 & v22f5fb4;
assign bd74e7 = hmaster2_p & v23f4426 | !hmaster2_p & v23070c1;
assign v22fef4f = busreq_p & v22fb4e3 | !busreq_p & !v22f7f74;
assign v22f6894 = hbusreq3_p & v2300523 | !hbusreq3_p & v22f9124;
assign v230d45f = hmaster2_p & v23f6bc1 | !hmaster2_p & v22f0824;
assign v22f9c37 = hgrant1_p & v84561b | !hgrant1_p & !v23f36f9;
assign v22f1585 = hbusreq1_p & v23fb2f5 | !hbusreq1_p & v84561b;
assign v2392ea0 = hbusreq2_p & v22ef772 | !hbusreq2_p & v84564d;
assign v22f3e8d = hburst1_p & v230cb1f | !hburst1_p & v84561b;
assign v23fbb4e = hlock0_p & v84564d | !hlock0_p & !v23fcab0;
assign v8b4671 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v9b93b3;
assign v2305aea = hbusreq3 & v23fcf96 | !hbusreq3 & v84561b;
assign v22fde18 = hbusreq4 & v22ee9be | !hbusreq4 & v2301a42;
assign v22f7efa = hlock2_p & v23fba6b | !hlock2_p & !v84561b;
assign v22ee6e8 = hmaster2_p & v22f0b79 | !hmaster2_p & v22f61b6;
assign v22f561a = hlock1_p & v2393f41 | !hlock1_p & addc42;
assign v2304672 = hgrant5_p & v2311ed7 | !hgrant5_p & v22fbfaf;
assign v23f08e5 = hgrant0_p & v230f5d0 | !hgrant0_p & !v230f1a7;
assign v230ad60 = hbusreq4_p & v23fb9d9 | !hbusreq4_p & v84561b;
assign v22f36a0 = hbusreq3 & v23fbe4f | !hbusreq3 & v84561b;
assign v23f4b56 = stateG2_p & v84561b | !stateG2_p & v23f906a;
assign v23fd01e = hgrant3_p & v23f37bf | !hgrant3_p & v230c3f5;
assign v21ea5eb = decide_p & v17a2d5a | !decide_p & v2309543;
assign v23f6b25 = locked_p & v2312fc4 | !locked_p & !v84561b;
assign v23ef95f = jx0_p & v84561b | !jx0_p & v2391d8a;
assign v23f79a9 = hbusreq2_p & v106ae69 | !hbusreq2_p & v84561b;
assign v22f54a4 = hbusreq5_p & v2301511 | !hbusreq5_p & v23fa2ec;
assign v23f748c = hmaster0_p & v23fceb9 | !hmaster0_p & v22fa631;
assign v23083e6 = hbusreq5_p & v1e84012 | !hbusreq5_p & v22ef542;
assign v22f163a = hbusreq2_p & v23101ee | !hbusreq2_p & !v84561b;
assign v23fbce1 = hbusreq4 & v22f7a20 | !hbusreq4 & v84561b;
assign v2311b96 = hbusreq6_p & v23fc52e | !hbusreq6_p & v22efa95;
assign v23095b3 = hbusreq1 & v23fc96e | !hbusreq1 & v84561b;
assign v22edf4f = hbusreq3 & v191ab29 | !hbusreq3 & v2302131;
assign v2308bfc = hmaster0_p & v22f1962 | !hmaster0_p & b00aa6;
assign v22f257b = hmaster1_p & v22eb397 | !hmaster1_p & v1e8408c;
assign v23fcb5b = hbusreq2_p & v22eb334 | !hbusreq2_p & v84561b;
assign v22fc63c = locked_p & v84561b | !locked_p & v23f8134;
assign v22f9a75 = hmaster0_p & v23fc89e | !hmaster0_p & v22f03c8;
assign v23117f5 = hmaster2_p & v2302a4d | !hmaster2_p & !v23f55ea;
assign v2312d0e = hbusreq3_p & v22fb589 | !hbusreq3_p & v2310256;
assign v22f19f7 = hgrant1_p & v84561b | !hgrant1_p & v23fbadd;
assign v1e8404d = hmaster2_p & v845661 | !hmaster2_p & v22f92fa;
assign v1aad571 = hbusreq1_p & v23fc17b | !hbusreq1_p & v84561b;
assign v2311da7 = hbusreq4_p & v23fb818 | !hbusreq4_p & v2312cb9;
assign v22f89d5 = hgrant4_p & v23ef95f | !hgrant4_p & v23fb736;
assign v2303c9d = hmaster2_p & v22fef4f | !hmaster2_p & !v23f55ea;
assign v230c104 = hbusreq0 & v1aad5ad | !hbusreq0 & v2312775;
assign v23fcc36 = hlock0_p & v191a86f | !hlock0_p & v23fce86;
assign v23113b5 = hmaster2_p & v23fcba3 | !hmaster2_p & v191abc5;
assign v23faa0a = hbusreq6 & v230a67e | !hbusreq6 & v84561b;
assign v23f9b8f = hlock6_p & v2302efc | !hlock6_p & !v84561b;
assign v23f8787 = hbusreq4 & v22f0b0d | !hbusreq4 & v230bdad;
assign v2305abd = hmaster2_p & v230f9db | !hmaster2_p & v12cc2ef;
assign v22effdf = hmaster2_p & v23f58e5 | !hmaster2_p & v2304990;
assign v23fc0d0 = hmaster2_p & v84561b | !hmaster2_p & v22f2430;
assign v106a81a = hbusreq1_p & v106ae4a | !hbusreq1_p & v2304cc4;
assign v22f53f3 = start_p & v84561b | !start_p & !v230f4d3;
assign v2300437 = hbusreq1_p & v22f56d2 | !hbusreq1_p & !v2302e32;
assign v23fce25 = hmaster0_p & v2309c9d | !hmaster0_p & !v22f6315;
assign v231055e = hbusreq5_p & v23f6f4d | !hbusreq5_p & v84561b;
assign v22fee33 = hlock4_p & v84561b | !hlock4_p & !v84563a;
assign v23127b3 = hbusreq1_p & v22f8c2f | !hbusreq1_p & v231271d;
assign v23fc519 = hgrant5_p & v84561b | !hgrant5_p & !v2306bb2;
assign v23fb4cb = hlock1_p & v84564d | !hlock1_p & !v84561b;
assign v2311c0b = hgrant3_p & v22f8e29 | !hgrant3_p & v22ffcbf;
assign v23fba99 = hmaster2_p & v84561b | !hmaster2_p & !v845622;
assign v22f7ed8 = hmaster2_p & v23f052e | !hmaster2_p & v23f51da;
assign v22edbc3 = hmaster1_p & v23fc891 | !hmaster1_p & !v23f49cd;
assign v22fe44f = hmaster2_p & v84561b | !hmaster2_p & !v23fb9ad;
assign v8d1fa5 = hgrant3_p & v23f16dc | !hgrant3_p & v23f61e5;
assign v230eb9b = locked_p & v84561b | !locked_p & !v106a782;
assign v2312020 = hgrant0_p & v84561b | !hgrant0_p & !v106ae25;
assign v22f695c = hmaster2_p & v106a782 | !hmaster2_p & !v84561b;
assign v23f2eff = hmaster0_p & v23f58bb | !hmaster0_p & !v23fba12;
assign v230f485 = hbusreq5_p & v22f0faf | !hbusreq5_p & v84561b;
assign v2303fa0 = hbusreq6 & v230c0da | !hbusreq6 & v84561b;
assign v2301d40 = stateG10_5_p & v23fc384 | !stateG10_5_p & v845636;
assign v23efbfd = hmaster2_p & v2311255 | !hmaster2_p & v84561b;
assign v22ef62d = hbusreq3_p & v23faa78 | !hbusreq3_p & v23f87f4;
assign v2307ed4 = hbusreq2_p & v23f1a8d | !hbusreq2_p & v23fcb69;
assign v23fc19e = hmaster0_p & v2302f72 | !hmaster0_p & v22f98e7;
assign v23fc45d = jx3_p & b6f226 | !jx3_p & v23fbe6c;
assign v22f789c = hmaster2_p & v22f5db6 | !hmaster2_p & v23fbfc0;
assign v22f6e30 = hbusreq3 & v2307206 | !hbusreq3 & v845627;
assign v2300fb4 = hbusreq1_p & v2303558 | !hbusreq1_p & !v22fd25c;
assign v23f34b8 = hmaster0_p & v2392e6c | !hmaster0_p & v2304dc2;
assign v13aff46 = hbusreq3 & v22f6a3a | !hbusreq3 & v84561b;
assign b3772b = hbusreq6 & v23fb483 | !hbusreq6 & v230aa7a;
assign v23021e1 = hburst1_p & v84561b | !hburst1_p & v22f53f3;
assign v22ebbde = hbusreq6_p & v230de87 | !hbusreq6_p & v22f7d04;
assign v23f3940 = hbusreq5_p & v22eb32b | !hbusreq5_p & v84561b;
assign v2302f60 = hlock6_p & v23f460c | !hlock6_p & v22fa77b;
assign v23f4eb4 = hgrant0_p & v23fcf92 | !hgrant0_p & !v23fb1a6;
assign v23fc63a = jx0_p & aa51ef | !jx0_p & v22fef21;
assign v22ed8c4 = hbusreq3_p & v22f2eba | !hbusreq3_p & v230fb43;
assign v23fc529 = hburst0 & v22f3294 | !hburst0 & !v2309a51;
assign v2301319 = hbusreq1_p & v845636 | !hbusreq1_p & v22fbe28;
assign v23fb924 = hbusreq6 & v845620 | !hbusreq6 & v23f65f3;
assign v23fa14e = hmaster0_p & v22eafd6 | !hmaster0_p & !v22f39b4;
assign v230ae06 = hbusreq1_p & v23fcef5 | !hbusreq1_p & v22f92f8;
assign v22efeb6 = hbusreq6 & v2301800 | !hbusreq6 & !v95ca80;
assign v23016d9 = hbusreq4 & v22f9bed | !hbusreq4 & v22fe81e;
assign v22eee34 = hgrant1_p & v23000e2 | !hgrant1_p & !v22fac2f;
assign v230f256 = hgrant5_p & fc9434 | !hgrant5_p & v84561b;
assign v23fbce0 = hmaster2_p & v22f7b29 | !hmaster2_p & v23f5596;
assign v15072cc = hgrant3_p & v23fc020 | !hgrant3_p & v22f5471;
assign v22fab7b = hbusreq6_p & v23fbe56 | !hbusreq6_p & v84561b;
assign v22f8d58 = hgrant3_p & v84562d | !hgrant3_p & v2300142;
assign v22ec20d = hgrant3_p & v22f8be5 | !hgrant3_p & v22f61b1;
assign v23fc139 = hbusreq3 & v84564d | !hbusreq3 & v84561b;
assign v23f5dfe = hmaster0_p & v23f38b7 | !hmaster0_p & v23fb661;
assign v23fcccb = hmaster0_p & v23111d5 | !hmaster0_p & v230c95c;
assign v23fb4fd = hbusreq5_p & v23fc818 | !hbusreq5_p & v84561b;
assign v84563e = hburst0 & v84561b | !hburst0 & !v84561b;
assign v23fb479 = hmaster2_p & v22feb0d | !hmaster2_p & v23fb4c7;
assign v23fbd0e = hbusreq1_p & v230320e | !hbusreq1_p & !v23fcc36;
assign v23f77a4 = hmaster1_p & v230b9fc | !hmaster1_p & !v23f5deb;
assign v23fb4b6 = hbusreq0_p & v2307582 | !hbusreq0_p & v23fc9f1;
assign v22ff1b9 = hlock6_p & b15ae7 | !hlock6_p & v2301135;
assign v22f1c40 = hmaster2_p & v84564d | !hmaster2_p & v22f60c6;
assign v230c322 = hmaster0_p & v230b7fc | !hmaster0_p & v23fbf5d;
assign v23fc7c4 = hbusreq1_p & v106a782 | !hbusreq1_p & v23fbf92;
assign v23fc040 = hbusreq3 & v239214a | !hbusreq3 & v230e966;
assign v22f8209 = hbusreq2_p & v22efa3b | !hbusreq2_p & !v84561b;
assign v230ec04 = hgrant3_p & v84561b | !hgrant3_p & !v23f052e;
assign v1b8769e = hgrant5_p & v22f4d65 | !hgrant5_p & !v23060a6;
assign v106a8b9 = decide_p & v23f8263 | !decide_p & v22febdb;
assign v22f7063 = jx0_p & v22ed30e | !jx0_p & v22eb69b;
assign v22ed8fe = hmaster2_p & v22ecbbd | !hmaster2_p & v22eeb19;
assign v23fb9ec = hgrant3_p & v22f88ee | !hgrant3_p & v22f2d7c;
assign v22fdca9 = hbusreq5_p & v23fcf91 | !hbusreq5_p & v23fc745;
assign v22fd136 = hgrant2_p & v23fc1a7 | !hgrant2_p & v2302e32;
assign v23fac04 = stateG10_5_p & v230df30 | !stateG10_5_p & v23f8093;
assign v2307c2a = hmaster2_p & v22fe5b1 | !hmaster2_p & v2311072;
assign v23fce52 = hgrant3_p & v84561b | !hgrant3_p & v22f90a5;
assign v106ae69 = hbusreq2 & v23f1f6f | !hbusreq2 & v84561b;
assign v23f931e = hbusreq1_p & v84561b | !hbusreq1_p & v230eb9b;
assign v22f1cbc = hbusreq1 & v2312f7e | !hbusreq1 & !v23022b1;
assign v23034a4 = hmaster0_p & v22ef823 | !hmaster0_p & v23fc851;
assign v22edd9f = hbusreq6_p & v22f4ae7 | !hbusreq6_p & !v84561b;
assign v2308b33 = hmaster2_p & v23f0bf1 | !hmaster2_p & v23101b1;
assign v22f21f6 = hlock3_p & v22ec63d | !hlock3_p & v12cd903;
assign v23fcc11 = hgrant3_p & v2305cac | !hgrant3_p & v230f47e;
assign v23fb942 = hbusreq5 & v22f1389 | !hbusreq5 & v84561b;
assign d49f4d = decide_p & v2305b67 | !decide_p & v2306798;
assign c24eac = hgrant1_p & v230d64e | !hgrant1_p & b50bc7;
assign v22f4b6d = jx1_p & v84561b | !jx1_p & v1507a21;
assign v23f6954 = hmaster1_p & v2302c0e | !hmaster1_p & v23f65cd;
assign v22f97f5 = jx3_p & v230892a | !jx3_p & v2300359;
assign v23f4ccb = hlock5_p & v23127fb | !hlock5_p & v2300a5a;
assign v23fbba0 = hbusreq4_p & v22f446b | !hbusreq4_p & v23fc1ec;
assign v239346f = hgrant1_p & v22ff732 | !hgrant1_p & v22eb5dd;
assign v23fcc42 = hmaster2_p & v23fc393 | !hmaster2_p & !v23f4426;
assign v23fbc43 = hbusreq1_p & v23f4758 | !hbusreq1_p & v22f6a6e;
assign v23fb661 = hmaster2_p & v2310e40 | !hmaster2_p & v22f56d2;
assign v22f691e = hmastlock_p & v23fbab3 | !hmastlock_p & v84561b;
assign e1e722 = hbusreq3 & v23fb236 | !hbusreq3 & v23f3f73;
assign v23f817b = hbusreq3_p & v22fc4a3 | !hbusreq3_p & v22ec326;
assign v22f575a = hbusreq3 & v22eb60c | !hbusreq3 & v22ef062;
assign v22f4ba1 = hbusreq4_p & v23fc24c | !hbusreq4_p & !v84561b;
assign v23fc114 = hbusreq3 & v230bd81 | !hbusreq3 & v191aec6;
assign v2301e1a = hmaster2_p & v23f1879 | !hmaster2_p & v84561b;
assign v23f9682 = hgrant1_p & v230faec | !hgrant1_p & v22f518e;
assign v22ef040 = hmaster1_p & v2305819 | !hmaster1_p & v23130f6;
assign v230038a = hmaster2_p & v22ef062 | !hmaster2_p & v84561b;
assign v230d32a = hmaster1_p & v23fc97f | !hmaster1_p & !v22fd15a;
assign v845649 = start_p & v84561b | !start_p & !v84561b;
assign v23fc838 = hbusreq1 & v2312f7e | !hbusreq1 & v84561b;
assign v23041a1 = hbusreq5_p & v23035ba | !hbusreq5_p & v2391a43;
assign v23f475e = hbusreq6_p & v22f9392 | !hbusreq6_p & v23f165d;
assign v22ebdbc = hbusreq5_p & v22f2db0 | !hbusreq5_p & v1aae98c;
assign v23f7714 = hbusreq4_p & v23051a9 | !hbusreq4_p & v23fb66d;
assign v2312aec = hbusreq1 & v23fcaf0 | !hbusreq1 & v230f010;
assign v22f17ed = hbusreq3_p & v23075a5 | !hbusreq3_p & v230cd87;
assign v230fc56 = hbusreq1_p & v845622 | !hbusreq1_p & v23fc614;
assign v2393c38 = hbusreq3 & v23fc881 | !hbusreq3 & v84561b;
assign v22f46ab = hbusreq2 & v230cff9 | !hbusreq2 & v84561b;
assign v22fc92d = hbusreq4 & v22f954a | !hbusreq4 & v23fd015;
assign v22f4809 = hlock3_p & v230b0f6 | !hlock3_p & v230c034;
assign v23fca08 = hmaster2_p & v84561b | !hmaster2_p & !v22f1ae5;
assign v23fb9fc = hbusreq3_p & v23fa3b6 | !hbusreq3_p & v84561b;
assign v23fb6bd = hbusreq6_p & v23f4cc1 | !hbusreq6_p & v230fe9b;
assign v22fe367 = hbusreq0_p & v23fc2fc | !hbusreq0_p & v845629;
assign v23f34d5 = hbusreq1_p & v23fc9b6 | !hbusreq1_p & !v84561b;
assign v23fc7d6 = hmaster0_p & v84564d | !hmaster0_p & v23fc3a4;
assign v22fb386 = stateG3_0_p & v845665 | !stateG3_0_p & !v84561b;
assign v23f49b3 = hbusreq5_p & v230aded | !hbusreq5_p & v2306f00;
assign v23f2f8d = hmaster2_p & bc96dd | !hmaster2_p & v2307b06;
assign v106ae19 = hmastlock_p & v23f906a | !hmastlock_p & !v84561b;
assign v9ee8a4 = stateG10_5_p & v84561b | !stateG10_5_p & e1df2d;
assign v23001a4 = hgrant5_p & v22f3754 | !hgrant5_p & v23fc3cb;
assign v23fc142 = hbusreq4_p & v22f4bcc | !hbusreq4_p & v23fc04e;
assign v22f0218 = hgrant1_p & v22f3d5a | !hgrant1_p & v22f2319;
assign v23f2602 = hbusreq3_p & v23f4a02 | !hbusreq3_p & v23fc232;
assign v23fc384 = hbusreq5 & v22ff33b | !hbusreq5 & !v84561b;
assign v22fdd6b = hmaster1_p & v230193c | !hmaster1_p & v230e97b;
assign v231142b = jx1_p & v230aa9b | !jx1_p & v2393c3f;
assign v22fb2dc = hlock4_p & bfde5b | !hlock4_p & v2311928;
assign v22f149c = hbusreq3_p & v22f4626 | !hbusreq3_p & v230c132;
assign v22f19ce = hmaster2_p & v1506ffd | !hmaster2_p & !v23fa345;
assign v13afeef = stateG10_5_p & v22f288e | !stateG10_5_p & v22ee956;
assign v22f9403 = hbusreq3_p & v23fc8a5 | !hbusreq3_p & v84561b;
assign v2308a42 = hbusreq0 & v23fb2e5 | !hbusreq0 & v84561b;
assign v22f6e56 = hgrant3_p & v23f2e5d | !hgrant3_p & v23fb4e8;
assign v22f8440 = hmaster2_p & v2304421 | !hmaster2_p & v22eb415;
assign v2392d61 = hmaster2_p & v22fccf1 | !hmaster2_p & v23f4201;
assign v23fbd46 = hmaster0_p & v22eeb7a | !hmaster0_p & !v23fc67b;
assign v2303f9a = hbusreq2_p & v84564d | !hbusreq2_p & !v84561b;
assign v23f85b0 = hmaster0_p & v23fcf94 | !hmaster0_p & v23fbdfd;
assign v22ffb10 = hgrant1_p & v84561b | !hgrant1_p & v23fc215;
assign v230f933 = hbusreq1_p & v22f8da3 | !hbusreq1_p & b7427f;
assign v23fd017 = hbusreq1_p & v230704c | !hbusreq1_p & b7427f;
assign v2305a69 = hbusreq3_p & v22f8be5 | !hbusreq3_p & !v23fcf5b;
assign v23fc5fe = hgrant0_p & v845620 | !hgrant0_p & v23017f0;
assign v23fc02e = hmaster0_p & ae78a6 | !hmaster0_p & v1507317;
assign v2391545 = hbusreq2_p & v23fbb70 | !hbusreq2_p & !v84561b;
assign v230bdd9 = hbusreq5_p & v22f5fa1 | !hbusreq5_p & v22f3a6f;
assign v22fe497 = hgrant1_p & bd7c1c | !hgrant1_p & v23f595d;
assign v23fc898 = hbusreq3_p & v23132cd | !hbusreq3_p & !v84561b;
assign v22f2b59 = jx3_p & v84561b | !jx3_p & v22ec37c;
assign v230383e = hlock5_p & v23f37ba | !hlock5_p & !v84561b;
assign v2303350 = hlock5_p & v23fbca4 | !hlock5_p & !v84561b;
assign v22fdfdd = hmaster2_p & v22f9927 | !hmaster2_p & !v22fbeea;
assign v98d402 = hbusreq3_p & v23f4f13 | !hbusreq3_p & v2393769;
assign v23fcaa1 = stateG2_p & v84561b | !stateG2_p & !v23fc249;
assign v23097f5 = hbusreq4_p & v23f29f5 | !hbusreq4_p & v23fc738;
assign v22f954a = hlock3_p & v22f1f78 | !hlock3_p & v22f5218;
assign v23fc681 = hbusreq0 & v2301e25 | !hbusreq0 & v84561b;
assign v22fbd9a = hmaster2_p & v22ff05e | !hmaster2_p & !v2307b06;
assign v22f2281 = hgrant3_p & v84562e | !hgrant3_p & v22f407c;
assign v22fa976 = hbusreq6_p & a8b64b | !hbusreq6_p & v2308b24;
assign v22f214f = hgrant5_p & v84561b | !hgrant5_p & v23fc9aa;
assign v22f61b6 = hgrant1_p & v84561b | !hgrant1_p & v22f8c0b;
assign v22fda6e = hmaster2_p & v84561b | !hmaster2_p & !v84562a;
assign v230df15 = hbusreq2 & v2310d74 | !hbusreq2 & v84561b;
assign v230faec = hbusreq1_p & v99d709 | !hbusreq1_p & !v84561b;
assign v22f9f88 = hmaster2_p & v84561b | !hmaster2_p & v23fb3c7;
assign v22f971b = hlock3_p & v22fe62a | !hlock3_p & v84562b;
assign v2310222 = hbusreq3_p & v23fc3e8 | !hbusreq3_p & !v22ec354;
assign abf9f6 = hmaster0_p & v23f537e | !hmaster0_p & v230ecb1;
assign v23fbffc = hbusreq2_p & v23fcd88 | !hbusreq2_p & v84561b;
assign v22fd008 = hgrant1_p & v845626 | !hgrant1_p & a37ffd;
assign v2302514 = hgrant3_p & v230f330 | !hgrant3_p & v22fa5a0;
assign v22f609b = hlock1_p & v23052c9 | !hlock1_p & v230e579;
assign v2313339 = hbusreq5_p & v230d1a6 | !hbusreq5_p & !v23fc463;
assign v22fc351 = hbusreq3 & v22eec6e | !hbusreq3 & v23f9d8e;
assign v23f25c8 = hbusreq1 & v22eefd1 | !hbusreq1 & v84561b;
assign v22f5037 = hbusreq2 & v23131e8 | !hbusreq2 & !v84561b;
assign v22fcc70 = hgrant4_p & v845632 | !hgrant4_p & v22fef4c;
assign v22f9838 = hlock0_p & v23f4ae1 | !hlock0_p & v22f6735;
assign f40d2a = hbusreq2 & v23fccfe | !hbusreq2 & v84561b;
assign v22f2e69 = hmaster2_p & v230d56c | !hmaster2_p & v2308818;
assign v13afed6 = jx1_p & v23fc3fe | !jx1_p & v22fafef;
assign v23930d2 = hlock5_p & v22f7885 | !hlock5_p & v845636;
assign b194d1 = hmaster2_p & v22fc10a | !hmaster2_p & v230971e;
assign v231254f = hmaster0_p & v23fc75d | !hmaster0_p & v22f853d;
assign v22ee889 = hbusreq5 & v23f6836 | !hbusreq5 & v84564d;
assign v2310b8a = hbusreq2_p & v2307e48 | !hbusreq2_p & v2309891;
assign v23f1b3c = hmaster2_p & v2304b35 | !hmaster2_p & bc96dd;
assign v22eedf9 = hbusreq2_p & v84562a | !hbusreq2_p & !v84561b;
assign v22f207c = hmaster0_p & v23fc002 | !hmaster0_p & v23fc048;
assign v2304bcb = hgrant3_p & v845635 | !hgrant3_p & v230bf51;
assign v22f36da = hbusreq3_p & v23fba7c | !hbusreq3_p & da38ba;
assign v23035c1 = hbusreq3_p & v22ee47d | !hbusreq3_p & v23fbfaa;
assign v23f43af = hbusreq2 & v1aae56f | !hbusreq2 & v84564d;
assign v230891d = hbusreq3_p & v23ef951 | !hbusreq3_p & v22ef663;
assign v230118f = hbusreq3 & v2306838 | !hbusreq3 & v868c84;
assign v17cf1d8 = hgrant1_p & v84561b | !hgrant1_p & v845625;
assign v23f307c = hgrant5_p & v84561b | !hgrant5_p & v23fc454;
assign v230ad74 = hbusreq6_p & v23fce1b | !hbusreq6_p & !fc8c53;
assign v230feae = hbusreq1_p & v22f3f15 | !hbusreq1_p & !v23faaef;
assign v22eaee8 = hmaster2_p & v191aa89 | !hmaster2_p & v2392d9f;
assign v23062f0 = hlock5_p & v23f2e61 | !hlock5_p & v230b04e;
assign v23fb522 = jx1_p & v85fd50 | !jx1_p & !v85fc1a;
assign v23f16fd = hlock0_p & v23fb66a | !hlock0_p & v23f7ffc;
assign v23fba1c = hbusreq2 & v23f5043 | !hbusreq2 & v84561b;
assign v2300cb6 = hgrant5_p & v23f84b2 | !hgrant5_p & v23f81cf;
assign v22ff1d8 = hbusreq4 & v22ee0d5 | !hbusreq4 & !v22ff914;
assign v1aae1af = hmaster1_p & v23fc25b | !hmaster1_p & v22fd49d;
assign v23fc880 = hbusreq3_p & v23f052e | !hbusreq3_p & v23fb906;
assign v23f4c32 = hbusreq5_p & v23f5af5 | !hbusreq5_p & v23f46ba;
assign v23024e8 = hmaster0_p & v22ed491 | !hmaster0_p & v23fc723;
assign v23015c2 = hmaster2_p & v845620 | !hmaster2_p & v23fbf24;
assign v23f64dd = hmaster0_p & v231347a | !hmaster0_p & v230def2;
assign v1aad34c = hbusreq6 & v84564d | !hbusreq6 & v23fbb35;
assign v230052f = hmaster2_p & v22f0126 | !hmaster2_p & v84561b;
assign v22eaec3 = hmaster0_p & v2310d59 | !hmaster0_p & v1aad67e;
assign v23fcb6f = hmaster2_p & v23101b1 | !hmaster2_p & v23fbddf;
assign v230875c = hbusreq5_p & v23f15ec | !hbusreq5_p & v2303ee8;
assign v231271d = hbusreq1 & v230ea6d | !hbusreq1 & !v845636;
assign v22ff890 = hbusreq5_p & v8f2065 | !hbusreq5_p & v8bb259;
assign v1506fe9 = hbusreq5_p & v9526ac | !hbusreq5_p & v23f972e;
assign v2303f89 = hbusreq1 & v23fcd4a | !hbusreq1 & v22f108e;
assign v231128c = hbusreq1_p & v22ed121 | !hbusreq1_p & v23fb625;
assign v22f6a1b = hgrant1_p & v2305b35 | !hgrant1_p & !v23f73d7;
assign v23fb625 = hbusreq1 & v22f0945 | !hbusreq1 & v84561b;
assign v23f6623 = hmaster1_p & v22f8e56 | !hmaster1_p & v2306bd7;
assign v23f8c22 = hbusreq1 & a68bda | !hbusreq1 & v84561b;
assign v23f849c = hbusreq1 & v22ef513 | !hbusreq1 & v84561b;
assign v2301652 = hbusreq3_p & v23015c2 | !hbusreq3_p & a7482d;
assign v23fbdf6 = hbusreq3_p & c20101 | !hbusreq3_p & v2300048;
assign v22fe59a = hbusreq0 & v13afe3a | !hbusreq0 & v84561b;
assign v23fb9aa = hgrant6_p & a4c73f | !hgrant6_p & v2305f67;
assign v23fbdb0 = hready & v22fc63c | !hready & v84564d;
assign v22fbb46 = hmaster1_p & v230236f | !hmaster1_p & v22ec2c0;
assign v23f5046 = hbusreq6 & v22f5941 | !hbusreq6 & v23f2bc0;
assign v22f7ce8 = jx1_p & v2391dd6 | !jx1_p & v23f9dd8;
assign v22f68fe = hgrant2_p & v2303f9a | !hgrant2_p & !v230333f;
assign v2310a9f = hbusreq1 & v22f60c6 | !hbusreq1 & !v2304ec7;
assign v2307d7f = hbusreq3 & v230b267 | !hbusreq3 & !v84561b;
assign v23fcd0d = hgrant3_p & v230a2c6 | !hgrant3_p & v23efb5a;
assign v23fbbbd = hgrant5_p & v23f5d36 | !hgrant5_p & v23fc374;
assign v23fca17 = hmaster1_p & v23fa893 | !hmaster1_p & v84561b;
assign v22f5815 = hgrant1_p & v23fcd14 | !hgrant1_p & v2305833;
assign v22ee73b = hbusreq5_p & v84561b | !hbusreq5_p & v230eb9b;
assign v2301b70 = hbusreq3_p & v23f62d5 | !hbusreq3_p & v23fb52d;
assign v22f92b8 = hbusreq5 & v2302075 | !hbusreq5 & v84561b;
assign v230c73d = hbusreq3_p & v84561b | !hbusreq3_p & !v23f41c2;
assign v85b90c = hbusreq4_p & a48bb0 | !hbusreq4_p & v2301f5d;
assign v23f95e1 = hbusreq2 & v22f3959 | !hbusreq2 & !v84561b;
assign v23fbd08 = hbusreq6_p & v22f9414 | !hbusreq6_p & v22ecd3a;
assign v22ef39f = hlock3_p & v84561b | !hlock3_p & v23f53a0;
assign v23f9a36 = jx1_p & v22ebe70 | !jx1_p & v23fcb57;
assign v22ee24a = hlock6_p & v22fed40 | !hlock6_p & v23f6c8f;
assign v231086f = hbusreq2_p & v2309cfe | !hbusreq2_p & !v22fc3ed;
assign v22f4e1f = stateG10_5_p & v23f81cf | !stateG10_5_p & v22ee9be;
assign v23fc12b = hbusreq5_p & v12cc317 | !hbusreq5_p & v23095d8;
assign v23f7b85 = hmaster0_p & v23fb132 | !hmaster0_p & !v23fcbe2;
assign v239383b = stateG10_5_p & v23fbd42 | !stateG10_5_p & v23fb8fa;
assign v23fa950 = hmaster0_p & e1de6f | !hmaster0_p & v22f9552;
assign a1fd35 = stateG2_p & v84561b | !stateG2_p & v23fcb5d;
assign v23fc7fe = hmaster1_p & v23f05e3 | !hmaster1_p & v2303507;
assign v22fef6a = hmaster0_p & v22fbdbc | !hmaster0_p & v22f3262;
assign v23fcf44 = hmaster0_p & v22f2009 | !hmaster0_p & v23fc08e;
assign v2311a61 = hbusreq3_p & v23fb553 | !hbusreq3_p & v23fba11;
assign v12cd2e3 = hmaster2_p & v84561b | !hmaster2_p & !v2310bdf;
assign ad89b5 = hmaster2_p & v23f87f4 | !hmaster2_p & v22f0593;
assign v23fc95a = hmaster2_p & v2310d04 | !hmaster2_p & v23f3997;
assign v23f47e3 = hmaster2_p & v2313255 | !hmaster2_p & v84561b;
assign v2310a63 = hbusreq5 & v22f0add | !hbusreq5 & v84561b;
assign v23fbc53 = hbusreq6 & v22f8ec8 | !hbusreq6 & v84561b;
assign v23fb172 = hbusreq2_p & v2300d6c | !hbusreq2_p & !v84561b;
assign v23fc095 = jx0_p & v22ffed0 | !jx0_p & v23fcb01;
assign v22ed12b = hbusreq4 & v22f799b | !hbusreq4 & v23f925b;
assign v2392c72 = hbusreq1_p & v1aae56f | !hbusreq1_p & v106ae21;
assign v22f9183 = hgrant3_p & v23088ef | !hgrant3_p & v22ff0da;
assign v23092cd = hbusreq4 & v23fbcbf | !hbusreq4 & v84561b;
assign v230c4ea = hmaster2_p & v23fcf69 | !hmaster2_p & v23fc716;
assign v230c398 = hmaster0_p & v1aae22e | !hmaster0_p & v22ec7e8;
assign v23fcf5c = hgrant2_p & a1fba6 | !hgrant2_p & v22f80b8;
assign v230aa0b = hlock3_p & v23053bd | !hlock3_p & !v23f1726;
assign v2308aef = hbusreq5_p & v15071d8 | !hbusreq5_p & v23efed1;
assign v230ab7a = hmaster1_p & v22fa8d7 | !hmaster1_p & !v23f6710;
assign v22f7919 = busreq_p & v84561b | !busreq_p & v23fbda6;
assign v22f9dd0 = hgrant5_p & v2305d15 | !hgrant5_p & v22ec61a;
assign v230164e = locked_p & v84561b | !locked_p & !v22f1691;
assign v230a905 = hmaster2_p & v23fbe41 | !hmaster2_p & !v23f32eb;
assign v2310900 = stateG10_5_p & v22f45a5 | !stateG10_5_p & v2303c39;
assign v2309475 = hbusreq1_p & v191a86f | !hbusreq1_p & !v191a879;
assign v23f7ae7 = hlock1_p & v22f12c8 | !hlock1_p & v23fc341;
assign v23fb9d3 = hbusreq4_p & v22f60ce | !hbusreq4_p & v230e80e;
assign v23f6d39 = hlock1_p & b9d00f | !hlock1_p & a1fbb6;
assign v2311268 = stateG10_5_p & v2310476 | !stateG10_5_p & !v23064ae;
assign v23fce6b = hbusreq1_p & v84561b | !hbusreq1_p & v23fc646;
assign v22f6953 = jx1_p & v23f651e | !jx1_p & v22eb47c;
assign v90af77 = hbusreq1_p & v22f115b | !hbusreq1_p & v239208c;
assign v23fb045 = hgrant3_p & v23fc0d8 | !hgrant3_p & v23f447e;
assign v23f96d1 = hmaster1_p & v2310406 | !hmaster1_p & v22ffdc3;
assign v1506a9c = hbusreq1 & v23fc0de | !hbusreq1 & !v22fbe28;
assign v23f580c = hbusreq1_p & v23fc432 | !hbusreq1_p & v84561b;
assign v23fc798 = hmaster2_p & v23fc48e | !hmaster2_p & v23fbaaa;
assign v23fb1fc = hmaster2_p & v23051c4 | !hmaster2_p & v23f53bd;
assign v22f065b = hgrant3_p & v23fc75d | !hgrant3_p & v23f80c9;
assign v2303075 = hbusreq5 & v845620 | !hbusreq5 & v22ee9be;
assign v230c0b2 = hbusreq1 & v23fd050 | !hbusreq1 & v23124cc;
assign v23f2c65 = hbusreq3_p & v22f6b7d | !hbusreq3_p & v230a226;
assign v23fbbd2 = hmastlock_p & v2308ae2 | !hmastlock_p & v84561b;
assign v23fd013 = jx1_p & v85e5cf | !jx1_p & v23fcf04;
assign v23fb82a = hbusreq3_p & v22eb02e | !hbusreq3_p & v22f0e99;
assign v22ff58f = hbusreq5_p & v22ecf87 | !hbusreq5_p & v22f288e;
assign v23fcffa = hgrant0_p & v22ee956 | !hgrant0_p & v23f72ff;
assign v22f264a = hbusreq5 & v2312acc | !hbusreq5 & v84561b;
assign v230156f = hmaster2_p & v22ed6c5 | !hmaster2_p & v22f9911;
assign v22f19a0 = hbusreq1_p & v2301a7d | !hbusreq1_p & !v84561b;
assign v22f10cc = hbusreq1_p & v23fbfe2 | !hbusreq1_p & v84561b;
assign v2302a58 = hmaster0_p & v23f9887 | !hmaster0_p & v23fc9d8;
assign v22fdc74 = hgrant5_p & v239367b | !hgrant5_p & !v230a58e;
assign v23fced1 = hmaster2_p & v22ec745 | !hmaster2_p & !v22f383b;
assign v23fcf4d = hgrant3_p & v23fbe79 | !hgrant3_p & v23f412d;
assign v23031c2 = hgrant1_p & v22f1cb7 | !hgrant1_p & v23f19e4;
assign v22ed236 = hmaster2_p & v22f5110 | !hmaster2_p & v23fb636;
assign v23fbcf0 = hmaster1_p & v2302fbf | !hmaster1_p & v22f3e5b;
assign v22f5941 = hbusreq3_p & v230fb9e | !hbusreq3_p & v22eaf73;
assign v22f2005 = hgrant3_p & v2308d63 | !hgrant3_p & v22f9f67;
assign v22f4b44 = hbusreq4 & v22ecb49 | !hbusreq4 & v230fac9;
assign v23f94bc = hbusreq5_p & v23fcd29 | !hbusreq5_p & v23fcccf;
assign v22f14d1 = hbusreq6_p & v22fe2b6 | !hbusreq6_p & v23f9dba;
assign v22f5a29 = hbusreq5_p & v22ee956 | !hbusreq5_p & v22f2653;
assign v12cd9b6 = hbusreq3_p & v2305ee5 | !hbusreq3_p & v22ee024;
assign v23fce3f = hgrant5_p & v2306cae | !hgrant5_p & v23925af;
assign v23f9150 = hbusreq3_p & v230fe87 | !hbusreq3_p & v106ae19;
assign v230fe87 = hmaster2_p & v106ae19 | !hmaster2_p & !b5f51c;
assign v23fc35e = hmaster0_p & v2306656 | !hmaster0_p & v23fcbe2;
assign v12cd5dd = hbusreq1_p & v23091e0 | !hbusreq1_p & !v106ae19;
assign v2307704 = hbusreq3 & v23fb578 | !hbusreq3 & v23936a3;
assign v23fc7e9 = hbusreq5 & v230b780 | !hbusreq5 & !v22fc6d7;
assign v23f482d = hbusreq3_p & v2305c78 | !hbusreq3_p & v231140b;
assign v23088db = hbusreq4 & v84561b | !hbusreq4 & !v23fba11;
assign v22f0e4e = hmaster2_p & a1fbb6 | !hmaster2_p & v230ceb6;
assign v23fc047 = hlock1_p & v230f82b | !hlock1_p & v23fba0b;
assign v22f3879 = hmaster0_p & v22ee394 | !hmaster0_p & v2304cd0;
assign v22f1d05 = hmaster0_p & v22f709c | !hmaster0_p & v191abd1;
assign v2309c93 = hlock0_p & v84561b | !hlock0_p & !v845622;
assign v22ebca0 = hgrant1_p & v845626 | !hgrant1_p & v23fcaa6;
assign v22f57e9 = hmaster2_p & v2309c8a | !hmaster2_p & v23f86f0;
assign hmaster2 = v23a2d0a;
assign v23fccb2 = hgrant1_p & v84561b | !hgrant1_p & v1aad4d7;
assign v22f6ac3 = hgrant0_p & v231151a | !hgrant0_p & !v84561b;
assign v22efda2 = hbusreq5_p & v23fc732 | !hbusreq5_p & v12cc72f;
assign v23f5dab = hlock0_p & v23f95e1 | !hlock0_p & v230c58d;
assign v23fc232 = hmaster2_p & v23131e8 | !hmaster2_p & !v2392974;
assign v23fbc6b = hmaster2_p & v845636 | !hmaster2_p & v23f75db;
assign v23059e1 = hbusreq3_p & v2303edc | !hbusreq3_p & v84561b;
assign v91c376 = hgrant1_p & v84561b | !hgrant1_p & v23f3b1d;
assign v2300382 = hgrant3_p & v84561b | !hgrant3_p & v23f9870;
assign v23fcfc4 = hbusreq4 & v23fc136 | !hbusreq4 & v23fb6b5;
assign v23fc613 = hlock4_p & v22fcea3 | !hlock4_p & v23fc9d6;
assign v2308c31 = hbusreq5_p & v23f90c4 | !hbusreq5_p & v23fb1e3;
assign v22fca12 = hlock4_p & v231008b | !hlock4_p & v84561b;
assign v17a34f9 = hbusreq5_p & v84562b | !hbusreq5_p & v23fb562;
assign v230af39 = hbusreq6_p & v230f069 | !hbusreq6_p & v23f6fe7;
assign v22eb359 = hgrant3_p & v84561b | !hgrant3_p & v23fa837;
assign v23041c1 = stateG10_5_p & v230e191 | !stateG10_5_p & v22ee956;
assign v23fcb67 = hmaster2_p & v230ea6d | !hmaster2_p & v22eeb07;
assign v22ff70d = hbusreq6 & v84564d | !hbusreq6 & v2300791;
assign v2310b15 = hbusreq4_p & v23fc613 | !hbusreq4_p & v23f2eff;
assign v23125e2 = hmaster1_p & v23fc4ce | !hmaster1_p & v84561b;
assign v22f4d61 = hmaster2_p & v23930d2 | !hmaster2_p & !v22eeb07;
assign v22fa1a2 = hmaster2_p & v23fc514 | !hmaster2_p & v2310bdf;
assign v23fc937 = hmaster0_p & v23f1a86 | !hmaster0_p & v23f561c;
assign v2303226 = hbusreq3_p & v22fb428 | !hbusreq3_p & !v23f5057;
assign v230d58c = hmaster2_p & a1fba6 | !hmaster2_p & v2302149;
assign v8fb6b6 = hmaster0_p & v230cc18 | !hmaster0_p & v23fc8e4;
assign v23f71c9 = stateA1_p & v22f3294 | !stateA1_p & !v84561b;
assign v2309aa0 = stateG10_5_p & v230e311 | !stateG10_5_p & v84562b;
assign v23f1f3e = hgrant0_p & v84561b | !hgrant0_p & v1aad4fb;
assign v22f1691 = busreq_p & v2305b74 | !busreq_p & !v230105a;
assign v23111da = hbusreq1_p & v23fc3dd | !hbusreq1_p & v22fd762;
assign bd74cf = hbusreq4 & v23fb483 | !hbusreq4 & v230aa7a;
assign bd7adc = hmaster2_p & v22f0218 | !hmaster2_p & v23fc203;
assign v23fc6ce = hbusreq3_p & v2306f5b | !hbusreq3_p & v22f848f;
assign v22f8cce = hbusreq6 & v22f6277 | !hbusreq6 & v23f91bc;
assign v23f3dc2 = stateG10_5_p & bd7786 | !stateG10_5_p & v2309c28;
assign v2308aec = hmaster2_p & v22f3643 | !hmaster2_p & v84564d;
assign v22f2805 = hbusreq3_p & v22fb589 | !hbusreq3_p & v230c521;
assign v22ec88f = hbusreq0_p & v22f7928 | !hbusreq0_p & v23fb57d;
assign v23127ef = hlock0_p & v23fcf46 | !hlock0_p & !v23fba6b;
assign v230829b = hmaster2_p & v230ef0b | !hmaster2_p & v2310d04;
assign v22f20c0 = hmaster2_p & v22ed0d9 | !hmaster2_p & v22fbe6a;
assign v2311f53 = stateG2_p & v84561b | !stateG2_p & v22f8088;
assign v23069b0 = hmaster0_p & v23fae84 | !hmaster0_p & v22f68f1;
assign v23fc5e9 = hbusreq3 & v22eefd1 | !hbusreq3 & v84561b;
assign v22ed8c2 = busreq_p & v23fbdcc | !busreq_p & v230efb1;
assign v23fba45 = hbusreq3 & v1aadb61 | !hbusreq3 & v2304a45;
assign v23fb8bf = hbusreq0_p & v191a86f | !hbusreq0_p & !v191a876;
assign v23f2f42 = hbusreq5_p & v23fc3cb | !hbusreq5_p & v230d976;
assign v22f7832 = hlock6_p & v22eba97 | !hlock6_p & v23f4900;
assign b15a69 = hgrant5_p & v23f4268 | !hgrant5_p & v22f69cc;
assign v230e817 = hmaster2_p & v84561b | !hmaster2_p & v23f68d8;
assign v22f135c = hbusreq1_p & v23fc8d3 | !hbusreq1_p & v23fc6b1;
assign v22eedac = hmaster2_p & e1df2d | !hmaster2_p & v84561b;
assign v22ff3d1 = hmaster2_p & v23f3ccf | !hmaster2_p & !v230cb9a;
assign v23fc32d = hmaster2_p & v23fcdc9 | !hmaster2_p & !v22fb8d6;
assign v23fc997 = hbusreq5_p & v2312acc | !hbusreq5_p & v23fcb5e;
assign v230de91 = hbusreq1_p & v22f1cbc | !hbusreq1_p & !v2307a62;
assign v84561b = 1;
assign v23fb5d8 = hlock0_p & v22ec992 | !hlock0_p & v230d529;
assign v22f25e0 = hmaster0_p & v2303bee | !hmaster0_p & v22ff67c;
assign v22fe62e = hbusreq6_p & v9ae0d1 | !hbusreq6_p & v23fc48a;
assign v22f8834 = locked_p & ab2d7c | !locked_p & v84561b;
assign v22fc508 = hbusreq3 & v22fa6a4 | !hbusreq3 & v22fad24;
assign v22f0e6b = hmaster2_p & v22eec6e | !hmaster2_p & v23f8ca4;
assign v15071d8 = hgrant0_p & v22ec303 | !hgrant0_p & !v2310af0;
assign v23fb598 = hbusreq5 & v845647 | !hbusreq5 & v84561b;
assign v23f1a2b = hbusreq6_p & v22eaf2a | !hbusreq6_p & v22f5c2b;
assign v22f9d19 = hmaster2_p & v22f1244 | !hmaster2_p & v230a574;
assign v23fcbdb = hbusreq3 & v2393420 | !hbusreq3 & v2307c2a;
assign v22ed35b = hbusreq6_p & bfce54 | !hbusreq6_p & v23f5cd7;
assign v2304e9c = stateG10_5_p & v230cf1a | !stateG10_5_p & !v106ae19;
assign v23fcf7a = hmaster2_p & v2304fae | !hmaster2_p & v23fcf89;
assign v23fbb39 = hbusreq3 & v22fb22e | !hbusreq3 & v2310d04;
assign v23fc92c = hgrant3_p & af7272 | !hgrant3_p & v2311a4a;
assign v22f1324 = hmaster0_p & v23fbf17 | !hmaster0_p & v2305400;
assign v1e8439a = hlock4_p & v23fcb75 | !hlock4_p & !v22f334c;
assign v150755e = hbusreq2_p & v22faef8 | !hbusreq2_p & v84561b;
assign v22fd69b = hgrant1_p & v23f68d8 | !hgrant1_p & v84561b;
assign v22ecbf0 = hmaster0_p & v23fc671 | !hmaster0_p & v2310b27;
assign v22fb7ef = hbusreq6 & v2304f11 | !hbusreq6 & v84561b;
assign v22fd0fb = hgrant6_p & v230754a | !hgrant6_p & v23f8848;
assign v2392867 = hmaster1_p & v22fd841 | !hmaster1_p & v23f7f35;
assign v23fa155 = hbusreq5_p & v23fa2ec | !hbusreq5_p & v23fc81c;
assign v2310d6a = hgrant1_p & v845626 | !hgrant1_p & v23f4d72;
assign v230a934 = hmaster2_p & v191a876 | !hmaster2_p & !v22ecc15;
assign v230f31f = hmaster0_p & v22f7ad4 | !hmaster0_p & !v23fcc9e;
assign e1dea8 = hbusreq6 & v23fbf8d | !hbusreq6 & v22f88bb;
assign v22ec9fa = hbusreq1_p & b425f1 | !hbusreq1_p & v84561b;
assign bd94fd = hbusreq4_p & v22f5019 | !hbusreq4_p & v84561b;
assign v230eeb6 = hmaster2_p & v2304b5d | !hmaster2_p & v23fbe1b;
assign v23fb083 = hbusreq6 & v23f6470 | !hbusreq6 & v23fa2ec;
assign v22ebccd = hbusreq3 & v23fb8c7 | !hbusreq3 & v12cd900;
assign v230a67e = hlock3_p & v2306d26 | !hlock3_p & v22f231d;
assign v23fc13a = hlock1_p & v2310a9f | !hlock1_p & !v84561b;
assign v22f3f9f = hbusreq4_p & v23fcb0d | !hbusreq4_p & v230b82e;
assign v23fbbb0 = hbusreq5 & v1aae98c | !hbusreq5 & v23fa2ec;
assign v23fbb30 = hbusreq6 & v22ebd72 | !hbusreq6 & v22ef9d0;
assign v22eb4a6 = hmaster0_p & v84561b | !hmaster0_p & v23642d5;
assign v23fb900 = hlock0_p & v22f9927 | !hlock0_p & v22ffc44;
assign v22f0bb6 = hbusreq4_p & v2304082 | !hbusreq4_p & b1e9fa;
assign v23005ea = hgrant3_p & b95000 | !hgrant3_p & v23fb487;
assign v23f8d64 = hbusreq5_p & v2305a12 | !hbusreq5_p & v22f39a5;
assign v23f6f06 = hbusreq4_p & v23096e7 | !hbusreq4_p & v22fc56c;
assign v22f7cbf = hbusreq4 & v22f8e1b | !hbusreq4 & da38c9;
assign v23fb188 = hgrant1_p & v22f56d2 | !hgrant1_p & v23fce9c;
assign v2313255 = hgrant1_p & v84561b | !hgrant1_p & v23061d7;
assign v230841a = hmastlock_p & v23fc0fd | !hmastlock_p & !v84561b;
assign v22f3068 = hlock6_p & v230ff52 | !hlock6_p & d97946;
assign v22ec012 = hmaster1_p & v230c1e1 | !hmaster1_p & v22f9b30;
assign v2303811 = hmaster2_p & v23fc98e | !hmaster2_p & !v22edcf1;
assign a8e3ee = hbusreq3 & v23f9507 | !hbusreq3 & !v84561b;
assign v2300aab = hbusreq1_p & v22fa7b8 | !hbusreq1_p & v84561b;
assign v23fc879 = hbusreq1 & v22f8ad4 | !hbusreq1 & v84561b;
assign v2304b4e = hbusreq2_p & v22f166c | !hbusreq2_p & v106a782;
assign v230e6ea = hgrant5_p & v22ff4c3 | !hgrant5_p & v230ae19;
assign v22fe46b = hbusreq2 & v23fb9ac | !hbusreq2 & v230561d;
assign v22f1b63 = hbusreq0 & v23fc01c | !hbusreq0 & v84561b;
assign v22f92ec = hbusreq0 & v23023c9 | !hbusreq0 & v84561b;
assign v23fcd6e = hbusreq6_p & v22fdb73 | !hbusreq6_p & v22f68c3;
assign v191a879 = hmastlock_p & v2310c2b | !hmastlock_p & v84561b;
assign v22fa70c = hbusreq0_p & v23fc976 | !hbusreq0_p & !v84561b;
assign v22f69eb = hlock1_p & v1b87673 | !hlock1_p & !v84561b;
assign v230e1bd = hmaster0_p & v23fb479 | !hmaster0_p & !v23fbd04;
assign a28a9e = hbusreq4_p & v23fb95a | !hbusreq4_p & v230f31f;
assign v22f76ae = hgrant1_p & v84561b | !hgrant1_p & v23fb811;
assign v1507a21 = hmaster1_p & v22f95e4 | !hmaster1_p & v23f6325;
assign v23fbea2 = hgrant3_p & v22f670f | !hgrant3_p & v23107fc;
assign v23fc5c5 = hgrant6_p & v23006c2 | !hgrant6_p & v1aadd09;
assign v2310c61 = hmaster1_p & v84561b | !hmaster1_p & !v2303102;
assign v23fc284 = hgrant3_p & v8c875e | !hgrant3_p & v230bf27;
assign v23fb59e = hbusreq0_p & v22f78ef | !hbusreq0_p & v84561b;
assign v22fe948 = stateG10_5_p & v22f70a0 | !stateG10_5_p & v23fc526;
assign v22f76c6 = hgrant3_p & b0fe84 | !hgrant3_p & v22f3dab;
assign v230a2ae = hmaster2_p & v22fe96a | !hmaster2_p & v23fc82c;
assign v23f7fb6 = hbusreq6 & v1aad8ea | !hbusreq6 & v84561b;
assign v23fc2cc = hlock5_p & b09503 | !hlock5_p & v84561b;
assign v230aa54 = hbusreq5 & v2301e25 | !hbusreq5 & v84561b;
assign v22f1f71 = hmaster2_p & v22f037a | !hmaster2_p & !v84561b;
assign v22fe009 = hbusreq0 & v230446f | !hbusreq0 & !v84562a;
assign v22f5d49 = hbusreq5 & v22ed6c5 | !hbusreq5 & v84561b;
assign v230fc36 = hlock3_p & v22ed942 | !hlock3_p & v22f5218;
assign v22eafea = hready & v84561b | !hready & !v23fbdfe;
assign v22ee1d1 = hbusreq3 & v22f993e | !hbusreq3 & v23f111b;
assign v23060ed = hmaster2_p & v23f8928 | !hmaster2_p & v22f249f;
assign v23fc34a = hmaster1_p & v23f957f | !hmaster1_p & v22f638b;
assign v2311d16 = hmaster1_p & v23fb936 | !hmaster1_p & v23fba52;
assign v22f61f6 = hmaster2_p & v23fbf8b | !hmaster2_p & !v22f954f;
assign v231329e = hlock6_p & v23f5b67 | !hlock6_p & !v84561b;
assign decide = !v2391935;
assign v231032d = hgrant0_p & v84561b | !hgrant0_p & v22f8603;
assign v2391cf3 = hbusreq4_p & v15071ed | !hbusreq4_p & v22f7347;
assign v22f6183 = hbusreq0 & v191a876 | !hbusreq0 & v84561b;
assign v22ee0c0 = hgrant3_p & v84561b | !hgrant3_p & !v22f20c0;
assign v22f7152 = hlock4_p & v22f5efe | !hlock4_p & v22fa502;
assign v23f39e6 = hmaster2_p & v191a86f | !hmaster2_p & v23fcc36;
assign v23f14e1 = hbusreq6 & v230c4e8 | !hbusreq6 & v230f0de;
assign v231192e = stateG10_5_p & v23f5140 | !stateG10_5_p & v23035ba;
assign v22eb2ee = hlock6_p & v23fbe9d | !hlock6_p & !v23f74b7;
assign v85fd50 = hmaster1_p & v845635 | !hmaster1_p & !v23f4ab4;
assign v2303cd6 = hbusreq3_p & v23fb60a | !hbusreq3_p & v1aadf44;
assign v23fbc83 = hbusreq3 & v2312888 | !hbusreq3 & v84561b;
assign v23f9758 = hbusreq3 & v231243e | !hbusreq3 & v84561b;
assign v23fbff9 = hmaster0_p & v2305bf5 | !hmaster0_p & v23f4c5b;
assign v23f47e1 = hgrant3_p & b23404 | !hgrant3_p & v23fc88b;
assign v22f8f0b = hbusreq2_p & v23fcbba | !hbusreq2_p & !v84561b;
assign v191b041 = hmaster2_p & v22feae3 | !hmaster2_p & v23f3b1e;
assign v230aa1f = hlock0_p & v23099de | !hlock0_p & v22f0fd7;
assign v22f7b29 = hgrant1_p & v23f6411 | !hgrant1_p & v22f0de9;
assign v22fba38 = hlock3_p & v23fc026 | !hlock3_p & v22f580d;
assign v22f0380 = hbusreq5_p & v845636 | !hbusreq5_p & v23043b8;
assign v230c24b = hgrant4_p & v2392d45 | !hgrant4_p & v23100d2;
assign v22ff6e8 = hbusreq0_p & v106af4d | !hbusreq0_p & v2303d1d;
assign v23f7fcb = hmaster0_p & v230f904 | !hmaster0_p & v22fbf38;
assign a1fee6 = hbusreq2 & v23117af | !hbusreq2 & v84564d;
assign v2392d14 = hbusreq1_p & v23f7b1d | !hbusreq1_p & v84561b;
assign v2307758 = hgrant1_p & v17a34ff | !hgrant1_p & e1dcf1;
assign v230e598 = hgrant5_p & v23077e6 | !hgrant5_p & !v23fc923;
assign v23fbad9 = hmaster1_p & v22f082c | !hmaster1_p & v23f6f06;
assign v22f2c30 = hlock0_p & v22f8d80 | !hlock0_p & !v845622;
assign v230842d = hbusreq4_p & v22eb52b | !hbusreq4_p & v23fce78;
assign v23f6721 = hlock0_p & v22fbea4 | !hlock0_p & !v22ff7d0;
assign v22f3789 = hbusreq0_p & v230f947 | !hbusreq0_p & !v22f1fec;
assign bd7f79 = hbusreq6 & v23fccd8 | !hbusreq6 & !v845636;
assign v23fb62b = hmaster2_p & v106ae19 | !hmaster2_p & !v23fcc9a;
assign v22f3692 = hbusreq5 & v2313118 | !hbusreq5 & v845620;
assign v23fd008 = hbusreq3_p & v23fbe91 | !hbusreq3_p & v84561b;
assign v2301178 = hbusreq1_p & v23f4f34 | !hbusreq1_p & v23f7796;
assign v22ff1f8 = hbusreq6 & v84564d | !hbusreq6 & v23055f4;
assign v23f4855 = hgrant1_p & v94e4a6 | !hgrant1_p & v22f08d0;
assign v23fc619 = hgrant0_p & v23fa2ec | !hgrant0_p & v23fd040;
assign v230cdc7 = hbusreq4_p & v22fdf70 | !hbusreq4_p & v23f3af2;
assign v23f71d5 = hbusreq5_p & v23fcf1f | !hbusreq5_p & v23fbdea;
assign v22f6e51 = hmaster0_p & v84561b | !hmaster0_p & v23fc722;
assign v1506ad8 = hgrant1_p & v22f67ef | !hgrant1_p & v23fc0bc;
assign v23929a6 = hbusreq5_p & v23f6bc1 | !hbusreq5_p & v23f92d5;
assign v23fc36b = hmaster0_p & v919672 | !hmaster0_p & !v2308e64;
assign v23fce64 = hgrant3_p & v22f368e | !hgrant3_p & v22ef648;
assign v22f7484 = hmaster2_p & v22f9880 | !hmaster2_p & !v22edcf1;
assign v22faa4d = hbusreq3 & v23f1032 | !hbusreq3 & b50a75;
assign v23fc26e = hbusreq5_p & v845629 | !hbusreq5_p & v23faaac;
assign v2308b2f = hmaster2_p & v23fcf83 | !hmaster2_p & v23fbe96;
assign v22fe74e = stateG10_5_p & v1aad4b2 | !stateG10_5_p & v845636;
assign v23fcc72 = hbusreq1_p & v15074eb | !hbusreq1_p & !v84561b;
assign v230cd17 = hlock4_p & v22ec5f2 | !hlock4_p & v84561b;
assign v22f4d20 = hgrant1_p & v845625 | !hgrant1_p & v2301178;
assign v23f5983 = hbusreq6_p & v1e84195 | !hbusreq6_p & v23faf72;
assign v23fc7e6 = hbusreq1 & v23fbfd0 | !hbusreq1 & v22f11f6;
assign v22f2d51 = stateG10_5_p & v2391a89 | !stateG10_5_p & v230af72;
assign v230f370 = hmaster2_p & v845620 | !hmaster2_p & v23f1207;
assign b23404 = hlock3_p & v230d6b6 | !hlock3_p & v230a226;
assign v2392a0d = hbusreq5_p & v22ff399 | !hbusreq5_p & v23f6890;
assign v23fc207 = stateG10_5_p & v22ef659 | !stateG10_5_p & v23065ad;
assign v23fb66d = hmaster0_p & v23934b5 | !hmaster0_p & v2304048;
assign v2311ed4 = hbusreq1_p & v23fca2a | !hbusreq1_p & !v23fc84b;
assign v22f3628 = hmaster2_p & v84561b | !hmaster2_p & v22ede4d;
assign v23fb2ea = hbusreq1_p & v22f5f7e | !hbusreq1_p & v230c93a;
assign v22f5471 = hmaster2_p & v23fbcfb | !hmaster2_p & v23101b1;
assign v23fc374 = hgrant0_p & v22fdc30 | !hgrant0_p & v23056e9;
assign v23f397b = hmaster0_p & v2300d5f | !hmaster0_p & v23f0588;
assign v22eb3aa = stateG2_p & v84561b | !stateG2_p & v23f2216;
assign v23fceb6 = hgrant1_p & v23fcda9 | !hgrant1_p & v23099c5;
assign v23f2837 = hbusreq3_p & v230f7ce | !hbusreq3_p & v230b8fe;
assign v22ed121 = hbusreq1 & v23f15ac | !hbusreq1 & v84561b;
assign v23fc7d5 = hready & v23f7326 | !hready & v22fab99;
assign v23107b6 = hbusreq1_p & v230f75a | !hbusreq1_p & !v22f2624;
assign v23f7f35 = hbusreq4_p & v22f41c4 | !hbusreq4_p & v22f75b0;
assign v230720b = hlock4_p & v230020c | !hlock4_p & v23102f3;
assign v23001d0 = hmaster0_p & v22fbd15 | !hmaster0_p & v23130c9;
assign v23fc9c8 = hgrant5_p & v23f23f1 | !hgrant5_p & v23fc19d;
assign v22f6d51 = jx0_p & v23047dd | !jx0_p & v22f7988;
assign bebe64 = jx2_p & v22ff294 | !jx2_p & v22fd030;
assign v23f3f40 = hmaster2_p & v12cc2ef | !hmaster2_p & !v22f3f2d;
assign v2302d1f = hlock0_p & v23f51b1 | !hlock0_p & v2305f58;
assign v22ff294 = hgrant4_p & v23fc9f2 | !hgrant4_p & v22f7b24;
assign v23f6858 = hbusreq5_p & v22f2957 | !hbusreq5_p & !v84561b;
assign v23fd002 = hgrant4_p & v1506a7a | !hgrant4_p & v230ea67;
assign v23f8ddb = hbusreq3 & v23f3d14 | !hbusreq3 & v84561b;
assign v22f0098 = hbusreq2_p & v23fb920 | !hbusreq2_p & v23fbc12;
assign v22ee3c9 = hbusreq6_p & v22f6c01 | !hbusreq6_p & v23fc49c;
assign v23fae84 = hbusreq3_p & v22f666d | !hbusreq3_p & v23f606c;
assign v23fc199 = hbusreq2 & v8d360e | !hbusreq2 & !v84561b;
assign v23f72ff = hgrant2_p & v2307ed4 | !hgrant2_p & v23fb5e8;
assign v22fd0cd = hgrant0_p & v23fbeaa | !hgrant0_p & v22ebf1f;
assign v23fa492 = hbusreq3 & v23fc01a | !hbusreq3 & v84561b;
assign v23fcebe = hmaster1_p & v23f8fc1 | !hmaster1_p & v23f5dd2;
assign v23fc416 = hbusreq1 & v13afe3a | !hbusreq1 & !v22fbb8a;
assign v23fb545 = hmaster0_p & v23126e2 | !hmaster0_p & v239223a;
assign v23fc3fe = hmaster1_p & v23fca5a | !hmaster1_p & v23fb673;
assign v23018c4 = hgrant1_p & v84561b | !hgrant1_p & v22f2db9;
assign v2309ae3 = hbusreq6_p & v230296a | !hbusreq6_p & v230cdc7;
assign v23fbb3c = stateG10_5_p & v23fc9d2 | !stateG10_5_p & v84564d;
assign v23fbfa0 = hbusreq6_p & v2309599 | !hbusreq6_p & v23f8db0;
assign v2303a62 = hmaster2_p & v8d360e | !hmaster2_p & v191a86f;
assign v230879e = hbusreq1_p & v2393739 | !hbusreq1_p & v84561b;
assign v22ee9d5 = hmaster2_p & v23065ad | !hmaster2_p & v230320e;
assign v22efbaa = hmaster0_p & v23fb1c3 | !hmaster0_p & a507a6;
assign v23fba11 = hmaster2_p & v845620 | !hmaster2_p & v84561b;
assign v23fb0ba = hlock2_p & v22f1b4e | !hlock2_p & !v23056b1;
assign v845623 = hlock0_p & v84561b | !hlock0_p & !v84561b;
assign v23115bd = hbusreq5_p & v84561b | !hbusreq5_p & v22f067b;
assign v22f0bb4 = hgrant1_p & v2312c3c | !hgrant1_p & v22f214f;
assign v23fa031 = jx1_p & v23f3768 | !jx1_p & v22fcf35;
assign v23fc6cc = hmaster2_p & v23f7ab7 | !hmaster2_p & v23f3997;
assign v23fbf1e = hgrant3_p & v84562e | !hgrant3_p & v22eb0b1;
assign v23040a5 = hmaster0_p & v22ffea8 | !hmaster0_p & e1e1ba;
assign v23062fe = hbusreq0_p & v23f1a8d | !hbusreq0_p & v23fcb69;
assign v23fb66f = hbusreq4_p & v2307eb9 | !hbusreq4_p & v230e71d;
assign v2308880 = hgrant1_p & v23fb498 | !hgrant1_p & v22f3e93;
assign v23fc5f4 = locked_p & da38c1 | !locked_p & v84561b;
assign v23fbf92 = hgrant5_p & v22f2730 | !hgrant5_p & v23fc6b3;
assign v2309d29 = hgrant2_p & v84561b | !hgrant2_p & v2302e76;
assign v23fa2c3 = hmaster0_p & v84561b | !hmaster0_p & v23fc263;
assign v22f2c87 = hmaster2_p & v84561b | !hmaster2_p & !v230d804;
assign v230d61c = hbusreq5_p & v22ee956 | !hbusreq5_p & v13afeef;
assign v23129e8 = hgrant3_p & v22faba5 | !hgrant3_p & v12cd3a7;
assign v22eedd0 = hbusreq5_p & a1fbc2 | !hbusreq5_p & v230b12a;
assign v22ee34a = hgrant2_p & v2310c7c | !hgrant2_p & v2302e32;
assign v2392803 = hlock2_p & v1b87673 | !hlock2_p & !v84561b;
assign v23fc3d4 = hbusreq1_p & v9526ac | !hbusreq1_p & v2304074;
assign v23fc2c8 = hgrant5_p & v230a774 | !hgrant5_p & v22f7ec4;
assign v23061de = hbusreq4_p & v22ee4e7 | !hbusreq4_p & v23fcc7c;
assign v23faa11 = jx1_p & v23017a9 | !jx1_p & v22fad67;
assign v2304060 = hmaster2_p & v23fc105 | !hmaster2_p & b50a75;
assign v23fc843 = stateG10_5_p & v23fbc07 | !stateG10_5_p & v84561b;
assign v23f3499 = jx3_p & v23056b2 | !jx3_p & v23fc855;
assign v22ee7cf = hmaster2_p & v23fcb5b | !hmaster2_p & v23f6b67;
assign v22eaed2 = hmaster0_p & v84561b | !hmaster0_p & !v2392fc4;
assign v23fbd64 = hbusreq3_p & v230e322 | !hbusreq3_p & v84561b;
assign v23f5868 = hgrant3_p & v22ffa6e | !hgrant3_p & v22ee2b4;
assign v13afeb1 = hbusreq6 & c043dc | !hbusreq6 & !v845636;
assign v23f5bf3 = hbusreq1_p & v23f2a7c | !hbusreq1_p & v23f2c8b;
assign v23068cd = hbusreq4 & v23f5a39 | !hbusreq4 & !v84561b;
assign b00ac7 = hmaster2_p & v23f87f4 | !hmaster2_p & v22fb1bc;
assign v23f8fc1 = hbusreq6_p & v22ebe13 | !hbusreq6_p & v23fbfb6;
assign v2303c5b = hmaster0_p & v22f7c44 | !hmaster0_p & !v230acb5;
assign v23fb599 = hlock6_p & v23f7086 | !hlock6_p & v23fcff5;
assign v22f151d = hbusreq6_p & v230ccaf | !hbusreq6_p & !v22f0bb6;
assign v23fc854 = hbusreq3_p & v23fc7a7 | !hbusreq3_p & v23fcc3d;
assign v23f5f4d = hmaster0_p & v22fea3f | !hmaster0_p & !v23031f0;
assign v22ef2c3 = hmastlock_p & v2301d76 | !hmastlock_p & v84561b;
assign v23fc5f5 = hmaster0_p & v230bb92 | !hmaster0_p & v230dcf9;
assign v230af81 = hbusreq5_p & v84562a | !hbusreq5_p & v2392fa3;
assign v22fe1ad = hbusreq3_p & v23fcd4b | !hbusreq3_p & v22ff9c5;
assign v22fa8e8 = hbusreq4_p & v23fcb1b | !hbusreq4_p & v23fb569;
assign v23f9e87 = hbusreq4_p & v15071ed | !hbusreq4_p & v22f6aa3;
assign v23fbc0d = hbusreq4_p & v22fb941 | !hbusreq4_p & v23f83de;
assign v2306126 = hmaster0_p & v84561b | !hmaster0_p & !v22ee345;
assign b6f226 = hmaster1_p & v23fcc89 | !hmaster1_p & v23f5deb;
assign v23fb473 = hbusreq2_p & v2302c08 | !hbusreq2_p & v22ee59c;
assign v22f243b = hmaster2_p & v23fcf46 | !hmaster2_p & v2306d29;
assign v23135a4 = hmaster2_p & v23f4d0d | !hmaster2_p & v84561b;
assign v22f19cb = hlock3_p & v23f7206 | !hlock3_p & !v84561b;
assign v23031c5 = hgrant3_p & v2308d63 | !hgrant3_p & v230b6e3;
assign v22f83fd = hmaster0_p & v22f2de3 | !hmaster0_p & v22fd522;
assign v22ef094 = hlock6_p & v23fb078 | !hlock6_p & v22fee33;
assign v23fb6c7 = hlock3_p & v2392537 | !hlock3_p & v22fe382;
assign v230e8d3 = hbusreq5_p & v22ec5f6 | !hbusreq5_p & v84561b;
assign v231228e = hlock0_p & v191a86f | !hlock0_p & v22fc58a;
assign v23fb5b9 = hmaster0_p & v2303acd | !hmaster0_p & v23fcb9c;
assign a090d5 = jx3_p & v23fcf10 | !jx3_p & v12cd9e0;
assign v23f5470 = hbusreq6_p & v23fcd45 | !hbusreq6_p & v23fbccc;
assign v23fbe00 = hbusreq5_p & v22f7cab | !hbusreq5_p & v230f222;
assign v23035a3 = stateG10_5_p & v23040f3 | !stateG10_5_p & !v230f34c;
assign v23fcc81 = hgrant1_p & v12cd5dd | !hgrant1_p & v22fa2dd;
assign v23fc687 = hmaster0_p & v22f4c34 | !hmaster0_p & !v23fbedb;
assign v23fcf4c = hbusreq6_p & v22fc0ec | !hbusreq6_p & v23fc067;
assign v22f5b73 = hbusreq0_p & adf3a3 | !hbusreq0_p & !v84561b;
assign v22f1aae = hgrant0_p & v22f56d2 | !hgrant0_p & !v22fd136;
assign v230933a = hgrant6_p & v23fc523 | !hgrant6_p & v23f1eac;
assign b7427f = hbusreq1 & v845620 | !hbusreq1 & v84561b;
assign v22f0faf = hlock5_p & a678c9 | !hlock5_p & v23fc55d;
assign v23fc6a3 = hbusreq3_p & v239281b | !hbusreq3_p & v23f3f59;
assign be29ff = hgrant3_p & v84561b | !hgrant3_p & v22f62ae;
assign v22f08d0 = hgrant5_p & v22f1a02 | !hgrant5_p & v22f0e5e;
assign v22fe315 = hbusreq6_p & v191b160 | !hbusreq6_p & v2392d8a;
assign v22f1e02 = locked_p & v12cd9cd | !locked_p & !v84561b;
assign v22feafc = hgrant1_p & b5f51c | !hgrant1_p & v2306f7b;
assign v2391cf8 = hmaster1_p & v230440f | !hmaster1_p & !v23ef987;
assign v22ef5c2 = hgrant1_p & v23fb6ff | !hgrant1_p & v191ae6e;
assign v230aeb3 = hbusreq1_p & v230d804 | !hbusreq1_p & v23f537c;
assign v238c168 = hbusreq1 & v1aae56f | !hbusreq1 & v84561b;
assign v2301a42 = hbusreq3_p & v23f1812 | !hbusreq3_p & v22ee9be;
assign v23f147c = hbusreq6_p & v22f41c4 | !hbusreq6_p & v22fd445;
assign v23fb998 = jx3_p & v22ef0a0 | !jx3_p & v23f53c1;
assign v2312bd9 = hgrant1_p & v84564d | !hgrant1_p & !v23fa1ad;
assign v23f8134 = hmastlock_p & v23083ed | !hmastlock_p & v84561b;
assign v23fca4e = hgrant3_p & v84561b | !hgrant3_p & !v2312f1b;
assign v2307add = hlock6_p & v22ff134 | !hlock6_p & v23fc24c;
assign v23fc726 = hbusreq1 & v9347cd | !hbusreq1 & v84561b;
assign v22fe6f8 = hbusreq6_p & v23139c9 | !hbusreq6_p & v22f05b4;
assign v22ecbbd = hgrant1_p & v230e28d | !hgrant1_p & v23fc3fb;
assign v23fc86a = hlock6_p & v23fc7d9 | !hlock6_p & !v22fcabb;
assign v230b68a = hmaster2_p & v230c727 | !hmaster2_p & v23f1bbf;
assign v23fbb64 = hmaster2_p & v23fbbf2 | !hmaster2_p & !v22f03cf;
assign v22f0755 = hbusreq1_p & v2306a5d | !hbusreq1_p & v23fcd0e;
assign v22f9ca3 = hmaster0_p & v23f8895 | !hmaster0_p & v96c563;
assign a2e978 = hgrant3_p & v22ee657 | !hgrant3_p & v22fb744;
assign v22f230d = hmaster1_p & v22f7f3f | !hmaster1_p & v22f7d00;
assign v2309c52 = hgrant1_p & v84561b | !hgrant1_p & v23f3724;
assign v23fb98f = hgrant0_p & v230a9eb | !hgrant0_p & v22fdaa0;
assign v22eda3a = hmaster2_p & v22f9911 | !hmaster2_p & v23f6836;
assign v22f4062 = hgrant3_p & v84561b | !hgrant3_p & v2309b33;
assign v23f3472 = hlock1 & v22fa682 | !hlock1 & v23f8deb;
assign v230f846 = hbusreq1_p & v23f9546 | !hbusreq1_p & v22fb8f1;
assign v22fa823 = hbusreq6_p & v23fbe7b | !hbusreq6_p & v22f2bc2;
assign v2311aad = hbusreq1 & v22f337b | !hbusreq1 & v845620;
assign v22f81ba = hbusreq3_p & c20101 | !hbusreq3_p & v23fbd56;
assign v2308b2e = hmaster2_p & v23fba9a | !hmaster2_p & v23f53bd;
assign v23f2d8c = hlock0_p & v230153d | !hlock0_p & v992f98;
assign v22fcc0d = hgrant0_p & v22ffb9d | !hgrant0_p & !v23fb682;
assign v22ece21 = jx0_p & v23057a4 | !jx0_p & v23fb998;
assign v23fa3bb = hbusreq4_p & v22ef144 | !hbusreq4_p & v22f57ea;
assign v23fb9c4 = hbusreq4_p & v230c398 | !hbusreq4_p & v23fc98b;
assign v23f8c92 = hbusreq3_p & v22f7319 | !hbusreq3_p & v84561b;
assign v22f4abc = hbusreq4 & v23fc8f6 | !hbusreq4 & v22eed0b;
assign v22ef99b = hgrant3_p & v84561b | !hgrant3_p & v230b9b4;
assign v191ace8 = hbusreq1 & v1aad481 | !hbusreq1 & v23fc7ef;
assign v230e37a = hmaster2_p & v22f19f7 | !hmaster2_p & v15070ca;
assign v12cd900 = hmaster2_p & v23fb565 | !hmaster2_p & !v23f5d72;
assign v22f2eba = hbusreq3 & b63b0c | !hbusreq3 & v22fc7b7;
assign v230a890 = hbusreq1_p & v2311a1d | !hbusreq1_p & v230c805;
assign v23fcfed = hmaster1_p & v22f47c6 | !hmaster1_p & v2312885;
assign v22f6ad2 = hbusreq1_p & v239174c | !hbusreq1_p & v230840f;
assign v908162 = hbusreq3_p & v22f7ed8 | !hbusreq3_p & v23122cf;
assign v23fbcbf = hmaster2_p & v22ff090 | !hmaster2_p & v84561b;
assign v22f639a = hmaster2_p & v22f337b | !hmaster2_p & v23f7123;
assign v231005a = hbusreq4_p & v230e8a7 | !hbusreq4_p & v23fd032;
assign v22f25ed = hmaster1_p & v23fbd08 | !hmaster1_p & !v2309d0b;
assign v22fc903 = hgrant3_p & v23060ff | !hgrant3_p & v22fa86d;
assign v230fa21 = hbusreq3_p & v2303bfd | !hbusreq3_p & v23fc0a4;
assign v230411f = stateG10_5_p & v23045ac | !stateG10_5_p & !v2309c8a;
assign v94e4a6 = hbusreq1_p & v22eeb03 | !hbusreq1_p & !v2311d0c;
assign v191b1a1 = hgrant4_p & v23fbdf3 | !hgrant4_p & v23fc63a;
assign v23115a7 = hbusreq4_p & v22f2ff1 | !hbusreq4_p & v22fdc16;
assign v12ce0d0 = hbusreq4 & v23fc52d | !hbusreq4 & v22efb25;
assign v23fc7e5 = hbusreq2 & v23fc443 | !hbusreq2 & v84561b;
assign v23fa1e3 = hgrant5_p & v2302f2c | !hgrant5_p & v22ee457;
assign v23f9044 = hbusreq1_p & v23f00ec | !hbusreq1_p & v23fa1e3;
assign v23fcbb2 = hgrant0_p & v23f68d8 | !hgrant0_p & v84561b;
assign v22fd666 = hmaster0_p & v22ede0b | !hmaster0_p & v2300aa8;
assign v22faa26 = hbusreq3_p & v23f0eec | !hbusreq3_p & v23f1225;
assign v23f56c3 = hbusreq3 & v22eaf73 | !hbusreq3 & v22f9160;
assign v230d99c = hbusreq4 & v2305bbb | !hbusreq4 & v23fb3a3;
assign v23f8895 = hbusreq3 & v84561b | !hbusreq3 & v845645;
assign v22f0ddd = hgrant0_p & v22ec303 | !hgrant0_p & !v23024b6;
assign v22eeaaf = stateA1_p & v23fc8d7 | !stateA1_p & !v84561b;
assign v22f6c1b = hgrant5_p & v84561b | !hgrant5_p & v84564f;
assign v22ebebe = hmaster2_p & v84561b | !hmaster2_p & v2301505;
assign b9c9cc = hmaster2_p & v23f3d14 | !hmaster2_p & v22ee9be;
assign v13b0055 = stateG10_5_p & v2391ada | !stateG10_5_p & v23fb096;
assign v22fb3f4 = hgrant3_p & v84561b | !hgrant3_p & v23faa19;
assign v23fcff1 = hgrant2_p & v845620 | !hgrant2_p & !v23f4e3d;
assign v22f99e3 = hmaster2_p & v22fc091 | !hmaster2_p & v84561b;
assign v23f68d8 = locked_p & b09503 | !locked_p & v84561b;
assign v23fc220 = hbusreq1 & v2307150 | !hbusreq1 & v84564d;
assign v23fb828 = hmaster0_p & v23f2810 | !hmaster0_p & v22f8cce;
assign v2310682 = hgrant1_p & v845625 | !hgrant1_p & v23fbbc2;
assign v22f3754 = hbusreq5_p & a1fbc2 | !hbusreq5_p & v2391fae;
assign v2305024 = hmaster2_p & v22fc96c | !hmaster2_p & v84561b;
assign v231114e = hbusreq0_p & v23fd045 | !hbusreq0_p & v230a8ea;
assign v2311967 = hmaster2_p & v2304bc1 | !hmaster2_p & v23112d5;
assign v8819d8 = hmaster2_p & v23082bc | !hmaster2_p & v2392ece;
assign v22fefa1 = hmaster0_p & v2307949 | !hmaster0_p & v230557c;
assign v230173a = hbusreq5_p & v23fc4f8 | !hbusreq5_p & v23fb6c2;
assign v23074dd = hmaster0_p & v23fc437 | !hmaster0_p & v23fcfd9;
assign v23f8466 = hmaster2_p & v106ae43 | !hmaster2_p & !v84561b;
assign v2308f5d = hmaster0_p & v23f72e4 | !hmaster0_p & f40c98;
assign v23f2c89 = hlock0_p & v22ef509 | !hlock0_p & v84561b;
assign v22f1a02 = hbusreq5_p & v23fcf46 | !hbusreq5_p & v2307a0f;
assign v23fc176 = hmaster2_p & v23113a4 | !hmaster2_p & v22fce73;
assign v22f0074 = hmaster1_p & v230723b | !hmaster1_p & v231324d;
assign v22f1037 = hgrant0_p & v23fc393 | !hgrant0_p & v230bf92;
assign v23fc4b2 = hlock5 & v22f20d3 | !hlock5 & v2304e69;
assign v22fd150 = hmaster2_p & v23fc362 | !hmaster2_p & v23f8036;
assign v23f2dbb = hbusreq4_p & v22fcef4 | !hbusreq4_p & v845637;
assign v22f32df = hbusreq6_p & v22ff0de | !hbusreq6_p & v22f0635;
assign v23fc0b9 = hmaster0_p & b3772b | !hmaster0_p & v22f7ee5;
assign v23f4194 = hbusreq3_p & v239228f | !hbusreq3_p & v12cd3aa;
assign v22f53b1 = hbusreq4_p & v22faf41 | !hbusreq4_p & v23f9c04;
assign v23f987b = hbusreq5 & v23052cc | !hbusreq5 & v84561b;
assign v191b0f9 = hbusreq6_p & v22ef9aa | !hbusreq6_p & v23fc081;
assign v22ecf87 = hgrant0_p & v22ee956 | !hgrant0_p & v22f7928;
assign v23f0a6b = hbusreq3_p & v22fa631 | !hbusreq3_p & v22ffdd1;
assign v230094d = hbusreq5 & v23fc23d | !hbusreq5 & v84561b;
assign v1b87890 = decide_p & v23fbd8c | !decide_p & v23f9f71;
assign v23f7b1d = hbusreq1 & b2aff2 | !hbusreq1 & v84561b;
assign v22f061c = hlock3_p & v23fcf17 | !hlock3_p & v230e9ef;
assign v23fb821 = hmaster0_p & v22fa101 | !hmaster0_p & v2311967;
assign v22f7159 = hbusreq0_p & v845620 | !hbusreq0_p & v22f9894;
assign v23fc885 = hmaster0_p & v23928ae | !hmaster0_p & v2311af8;
assign v23fcc7a = stateG10_5_p & v230fa13 | !stateG10_5_p & v23f4b28;
assign v86df86 = hmaster2_p & v23129e0 | !hmaster2_p & v2301797;
assign v23fb11d = hlock2_p & v22ede4d | !hlock2_p & v84561b;
assign f40618 = jx2_p & v84561b | !jx2_p & f40764;
assign v22ffab6 = hgrant3_p & v84561b | !hgrant3_p & v22f28e6;
assign v23fb673 = hbusreq6_p & v22ff36f | !hbusreq6_p & v22f6176;
assign v22eff0e = hburst1_p & v2309a51 | !hburst1_p & !v845649;
assign v22f41c0 = hbusreq3_p & v23fbea6 | !hbusreq3_p & !v23fbf3e;
assign v22fafa5 = hmaster2_p & bd7c3f | !hmaster2_p & v230c2b1;
assign v22fbc73 = hbusreq3_p & v230e54d | !hbusreq3_p & v22f7484;
assign v23f6a8a = hbusreq2_p & v22fef4f | !hbusreq2_p & v23fc393;
assign v23930d8 = hbusreq3_p & v23fbe89 | !hbusreq3_p & v23fc5de;
assign v22ef663 = hbusreq3 & v23f4fbf | !hbusreq3 & v230b304;
assign v22f04bf = hmaster0_p & v22f2e48 | !hmaster0_p & v22fd55f;
assign v22f1744 = hbusreq4_p & v22fd364 | !hbusreq4_p & v23fbe9d;
assign v23fc7ba = hbusreq1_p & v23046b5 | !hbusreq1_p & v23fbf93;
assign v22fce1f = hbusreq4_p & v23fb545 | !hbusreq4_p & v239223a;
assign v23fc605 = hbusreq5_p & v23f24c5 | !hbusreq5_p & v22f4e1f;
assign v23fbb9e = hbusreq6_p & v23fcd35 | !hbusreq6_p & v23f240c;
assign v23f6b67 = hlock0_p & v22fe421 | !hlock0_p & v23007b3;
assign v22f5eae = hmaster0_p & v2303e9a | !hmaster0_p & v22f4855;
assign v2305b34 = hbusreq3_p & v23fbdb9 | !hbusreq3_p & !v84561b;
assign v23fb3d1 = hbusreq5_p & v845636 | !hbusreq5_p & v23f31d3;
assign v22fbfe3 = hmaster0_p & b9c985 | !hmaster0_p & v22f85c0;
assign v23fc44e = hbusreq6 & v230e01b | !hbusreq6 & v23fcf4d;
assign v22f7d67 = hmaster0_p & v22ee521 | !hmaster0_p & !v1aae222;
assign v22ebc38 = hgrant4_p & v845632 | !hgrant4_p & v22eaf27;
assign v230677d = hgrant4_p & v845635 | !hgrant4_p & v22f2a85;
assign v2309ab5 = hbusreq5_p & v23fbb80 | !hbusreq5_p & v22ed1f3;
assign v23039be = hgrant2_p & v2308225 | !hgrant2_p & v84561b;
assign v22fb5da = hgrant1_p & v84561b | !hgrant1_p & !v22fe552;
assign v22ff18a = hbusreq3_p & v23070c0 | !hbusreq3_p & v22f2095;
assign v23f1686 = hbusreq4_p & v2301a5f | !hbusreq4_p & v23fbeaf;
assign v22f94ea = hbusreq1_p & v230bd05 | !hbusreq1_p & v2393417;
assign v23f5bdc = hburst0 & v23fa931 | !hburst0 & !v84561b;
assign v2306f84 = hbusreq1_p & v23052a8 | !hbusreq1_p & v84561b;
assign v2308e08 = hmaster2_p & v22fd271 | !hmaster2_p & v230b3a5;
assign v22f320d = hbusreq4_p & v230c3d2 | !hbusreq4_p & v23f18f2;
assign v23fc140 = hbusreq6_p & v2307a72 | !hbusreq6_p & v23fc44a;
assign bd74ba = hgrant3_p & v22f2ca2 | !hgrant3_p & v22f6265;
assign v23fc8a3 = hburst0_p & v22f178d | !hburst0_p & !v22f53f3;
assign v23f6ad0 = hbusreq3_p & v230c4c3 | !hbusreq3_p & v22eec47;
assign v1aad5c9 = hgrant5_p & v23fb159 | !hgrant5_p & !v22eb292;
assign v2302c0e = hbusreq6_p & v23fbc7f | !hbusreq6_p & v23f50f8;
assign v23fbfcf = stateG10_5_p & c258f4 | !stateG10_5_p & v22f3643;
assign v22f42d3 = hmaster0_p & v22f368e | !hmaster0_p & v23fc884;
assign v23f9a04 = hgrant1_p & v84561b | !hgrant1_p & !b13467;
assign v22fc8e1 = hbusreq3_p & v22ff6c5 | !hbusreq3_p & !v106ae19;
assign v23fc349 = hmaster0_p & v23fb526 | !hmaster0_p & v22ee75e;
assign v23fb13c = jx3_p & v1aae124 | !jx3_p & v22ef35b;
assign v23fc905 = hmaster2_p & v84561b | !hmaster2_p & v84562a;
assign v22fcb9d = hmaster1_p & v22fd841 | !hmaster1_p & v22fd445;
assign v2306597 = hbusreq1_p & v22ed614 | !hbusreq1_p & v22f8c0b;
assign v22f0719 = hbusreq3_p & v2310ff6 | !hbusreq3_p & v84561b;
assign v2303bfd = hbusreq3 & v23f6470 | !hbusreq3 & v23fa2ec;
assign v23fc78e = hbusreq1_p & v230bd05 | !hbusreq1_p & v22f6d58;
assign v22fc6e6 = hmaster2_p & v230b125 | !hmaster2_p & !v84561b;
assign v22fa766 = hbusreq5 & v23f81cf | !hbusreq5 & v84561b;
assign v2303ce3 = hmaster0_p & v23044f6 | !hmaster0_p & v230f0de;
assign v230bd81 = hmaster2_p & v23fb6e3 | !hmaster2_p & v2309b7e;
assign v22ee06a = hgrant1_p & v23113e8 | !hgrant1_p & v22f8694;
assign v23f7ab7 = hbusreq1_p & v23fc252 | !hbusreq1_p & v84561b;
assign v22fba9a = hmaster2_p & v22f12e5 | !hmaster2_p & v23fb7fc;
assign v22ec299 = hgrant5_p & v84561b | !hgrant5_p & v2311d12;
assign v23fc27a = hbusreq4_p & v23f29f5 | !hbusreq4_p & v22f4810;
assign v23fb6bb = hgrant1_p & v84561b | !hgrant1_p & !v23fbfe0;
assign v23078cb = hbusreq6 & v2308b14 | !hbusreq6 & v84561b;
assign v23fbb70 = hbusreq2 & v2310ad7 | !hbusreq2 & v22f3de9;
assign v23faca5 = hbusreq0 & v22ff315 | !hbusreq0 & v84561b;
assign v2302b3e = hbusreq3_p & v23fcbed | !hbusreq3_p & v23fbc96;
assign v231151a = hlock0_p & v23fba70 | !hlock0_p & !v84561b;
assign v23fc42e = hmaster1_p & v22f14d1 | !hmaster1_p & v1aad4b7;
assign v23f2d37 = hbusreq3_p & v22fa86d | !hbusreq3_p & v2305296;
assign v22f5d15 = hbusreq5_p & v845647 | !hbusreq5_p & !v22ff0d2;
assign v2303cda = hbusreq4 & v22fe5f9 | !hbusreq4 & v23f87f4;
assign v22f6a0e = hgrant0_p & v22fee46 | !hgrant0_p & v22eed66;
assign v230a9ca = hmaster1_p & v191ac87 | !hmaster1_p & v84561b;
assign v2307f77 = hbusreq3_p & v230e115 | !hbusreq3_p & v23fc340;
assign v2310e40 = locked_p & v230d2a8 | !locked_p & v191a879;
assign v23f7aea = hmaster2_p & bd7c3f | !hmaster2_p & v23fb838;
assign v2309a10 = hmaster2_p & a1fd0b | !hmaster2_p & v84564d;
assign v2301e9c = hbusreq1_p & v23f4e43 | !hbusreq1_p & !v84561b;
assign v23fbf44 = hlock1_p & v23fca56 | !hlock1_p & v23fa623;
assign v22f367c = hmaster2_p & v230882d | !hmaster2_p & !v22eb5b3;
assign v22f1f9f = hlock4_p & v1aae99f | !hlock4_p & !v23052b7;
assign v22fab33 = hmaster0_p & v23fcab7 | !hmaster0_p & !v22f2123;
assign v23f3c1b = hbusreq1_p & v2300387 | !hbusreq1_p & v22fd762;
assign v2304cc4 = hbusreq5_p & v106ae4a | !hbusreq5_p & v22f8cd8;
assign v22f2ece = hbusreq4 & v22ec354 | !hbusreq4 & !v84561b;
assign v23f1726 = hbusreq3_p & v2306bed | !hbusreq3_p & !v84561b;
assign v230cae4 = hbusreq3_p & v22f19ce | !hbusreq3_p & v2310a05;
assign v22f407c = hbusreq3_p & v2312ae4 | !hbusreq3_p & v1507045;
assign v2393420 = hmaster2_p & v22fe5b1 | !hmaster2_p & !v23fa63b;
assign v230197f = hbusreq4_p & v22f4089 | !hbusreq4_p & v22ee057;
assign v230363f = hready_p & v23fbe11 | !hready_p & v2307419;
assign v22fe37c = hbusreq5_p & v22f98e3 | !hbusreq5_p & v23f2c89;
assign v106aead = hbusreq1 & v23fc46b | !hbusreq1 & !v23fc4f5;
assign v23fc671 = hbusreq6 & v22fb554 | !hbusreq6 & v22f5583;
assign v22f5edf = hbusreq3 & v230b930 | !hbusreq3 & !v845645;
assign v23fc5c4 = stateG10_5_p & v22f7004 | !stateG10_5_p & !v2312259;
assign v2303650 = jx0_p & v23047dd | !jx0_p & v23f196c;
assign v22f939d = hbusreq3_p & v230ccc4 | !hbusreq3_p & !v22fd907;
assign v23fcec3 = stateG10_5_p & v230a941 | !stateG10_5_p & v84561b;
assign v23fcb75 = hmaster0_p & v22f2f3e | !hmaster0_p & bd74e7;
assign v23fb9ef = hgrant3_p & v22ee9d5 | !hgrant3_p & v2307009;
assign v1506a62 = hlock6_p & v23fcfda | !hlock6_p & v22f8824;
assign v22f2759 = stateA1_p & v22fb386 | !stateA1_p & v23fc8a3;
assign v17a2d5b = decide_p & v22ebd80 | !decide_p & v22f19c3;
assign v23fbfd0 = hready & v23fb95d | !hready & v13afe3a;
assign v23fba0a = hbusreq6_p & v1506a62 | !hbusreq6_p & v84561b;
assign v22f444f = hbusreq6 & v23018ac | !hbusreq6 & v22f38db;
assign be9b63 = hgrant1_p & v22ff732 | !hgrant1_p & v230d921;
assign v22f2ffe = hmaster2_p & v23fbed5 | !hmaster2_p & v84561b;
assign v22f43c9 = hmaster1_p & v2311919 | !hmaster1_p & v84561b;
assign v22faa66 = hmaster2_p & v845620 | !hmaster2_p & v23fc023;
assign v2302225 = hlock0_p & v84561b | !hlock0_p & v23faca5;
assign v106ae8b = hbusreq3_p & v23f60fb | !hbusreq3_p & v230b739;
assign v23f4096 = stateG2_p & v84561b | !stateG2_p & v23fc8a3;
assign v23006e9 = hgrant5_p & v22ed148 | !hgrant5_p & v23920d8;
assign v23fbf06 = hlock6_p & v22f1744 | !hlock6_p & !v23fc4e2;
assign v22f48b7 = hmaster0_p & v230b8fb | !hmaster0_p & !v23130d6;
assign v23029bb = hlock3_p & v23fc2df | !hlock3_p & v22f03a7;
assign v2306494 = hbusreq1 & v22f925b | !hbusreq1 & v84564d;
assign v23fc53b = hmaster2_p & v230031f | !hmaster2_p & v22fb1bc;
assign v230cbdd = hbusreq0 & v23fc7d5 | !hbusreq0 & v22f0add;
assign v23fcffb = hmaster2_p & v23f80c1 | !hmaster2_p & v23f024e;
assign v1aadc9e = hmaster0_p & v23fb1ca | !hmaster0_p & v22f8f2b;
assign v22ee499 = hgrant3_p & v84562e | !hgrant3_p & v23fb1fc;
assign v230278e = stateG10_5_p & v22f322a | !stateG10_5_p & v84561b;
assign v23f7605 = stateG2_p & v22f9369 | !stateG2_p & b8656c;
assign v22fa4df = hbusreq4 & v23064ad | !hbusreq4 & v239233a;
assign v23fcf62 = hlock6_p & v22f5272 | !hlock6_p & !v23094c7;
assign v23f1925 = jx0_p & v22fca43 | !jx0_p & v23fbf90;
assign v23f7ff2 = hbusreq4_p & v23fc6af | !hbusreq4_p & v22f1683;
assign v22f9e5b = hbusreq0 & v23105cd | !hbusreq0 & !v230e6ee;
assign v2307946 = hbusreq0_p & v23fbb3e | !hbusreq0_p & v84561b;
assign v23fa8c8 = hmaster2_p & v23fc84b | !hmaster2_p & !v22f0824;
assign v23efdcb = hmaster2_p & v2306932 | !hmaster2_p & v23f763f;
assign v2306da6 = hmaster0_p & v2300d5f | !hmaster0_p & v22f6ae5;
assign ae0418 = hmaster2_p & v23105cd | !hmaster2_p & v22fef02;
assign v22fa415 = hmaster2_p & v23f8da8 | !hmaster2_p & v23fce71;
assign v22fbb33 = hbusreq3_p & bd74e7 | !hbusreq3_p & v22f16bf;
assign v23f6d6c = hbusreq1_p & v23fc879 | !hbusreq1_p & v84561b;
assign v230554d = hmaster2_p & v2309d55 | !hmaster2_p & !v84561b;
assign v22fe820 = hmaster0_p & v23fb479 | !hmaster0_p & v23f8013;
assign v23fcf87 = hgrant3_p & v22f82cd | !hgrant3_p & v23fc2c6;
assign v22f3b00 = hmaster2_p & v23f9a04 | !hmaster2_p & v2312ad2;
assign v22ef530 = jx2_p & v22f26d2 | !jx2_p & v23fc6dd;
assign v22f3add = hmaster2_p & v22fd0e6 | !hmaster2_p & v23f8ca4;
assign v22f0445 = hbusreq4_p & v2308a1b | !hbusreq4_p & v22ec6c7;
assign v23fccf5 = hmaster2_p & v22f9a51 | !hmaster2_p & !v1aad847;
assign v22f69cc = hgrant2_p & v84561b | !hgrant2_p & v2301511;
assign v23fc733 = hlock5_p & v2305fe0 | !hlock5_p & v84564d;
assign v2308506 = hmaster1_p & v84561b | !hmaster1_p & v23039af;
assign v22ef100 = hbusreq6_p & v22f2214 | !hbusreq6_p & v2303051;
assign v22f4114 = hbusreq1_p & v23fcea8 | !hbusreq1_p & v23fc98a;
assign v22fcaa6 = hmaster0_p & v23fc7b9 | !hmaster0_p & !v23fcf51;
assign v23faa78 = hmaster2_p & v23f87f4 | !hmaster2_p & v23f7700;
assign v23fcfd3 = hbusreq3 & v22f16ef | !hbusreq3 & v230038a;
assign v23f6aab = jx1_p & v2309532 | !jx1_p & v2301e40;
assign v230d8af = hmaster2_p & a1fbc2 | !hmaster2_p & v22ff732;
assign v230bb2a = hbusreq5_p & v22f8271 | !hbusreq5_p & !v2312839;
assign v23f925b = hbusreq3_p & v2301a04 | !hbusreq3_p & v23060e3;
assign v23fc6f3 = hbusreq2_p & v22f1b4e | !hbusreq2_p & v22ed7a8;
assign v23effbc = hbusreq0_p & b9888a | !hbusreq0_p & v22ffb52;
assign v23132db = hmaster0_p & v22ec354 | !hmaster0_p & v22efe81;
assign v23088b3 = hbusreq2_p & fc8e3a | !hbusreq2_p & !v84561b;
assign v23fa63b = hbusreq2_p & v23fcfcd | !hbusreq2_p & v84561b;
assign v23f839a = hlock6_p & v23045fa | !hlock6_p & b52881;
assign v23fcd0c = hgrant1_p & v2313463 | !hgrant1_p & !v23fcb10;
assign v23fb155 = hgrant1_p & v23f5af5 | !hgrant1_p & v23fbe8b;
assign v2393ecb = jx1_p & v23fc42e | !jx1_p & v230e94e;
assign v22f3af7 = hbusreq3_p & v22ed8a3 | !hbusreq3_p & !v84561b;
assign b9d061 = hgrant1_p & v12cd6a1 | !hgrant1_p & v23f4634;
assign v2306c0c = hlock3_p & v23f9a5b | !hlock3_p & !v2309eab;
assign v23fa3a4 = hgrant0_p & v2303b76 | !hgrant0_p & v23f0652;
assign v23fbbf9 = hmaster2_p & v84561b | !hmaster2_p & !v22f92fa;
assign v22eaaba = hbusreq1_p & v23f3a16 | !hbusreq1_p & v2309871;
assign v23fc6b6 = hbusreq3_p & v23fc5d0 | !hbusreq3_p & v23fc2d7;
assign v15070d3 = hlock0_p & v23fba79 | !hlock0_p & v22f0470;
assign v23f8747 = hgrant2_p & v2310904 | !hgrant2_p & !v23fb861;
assign v2308dcf = hbusreq6 & v84564d | !hbusreq6 & v22f23a1;
assign v230b8fb = hmaster2_p & v230fc8c | !hmaster2_p & v2301ef1;
assign v22f5fa1 = hlock5_p & v22f6397 | !hlock5_p & v84562b;
assign v22fcf3e = hbusreq2 & v13affaa | !hbusreq2 & v84564d;
assign v22eeb06 = hmaster2_p & v23f87f4 | !hmaster2_p & v23fcda9;
assign v23fc17f = hmaster0_p & v22fb10b | !hmaster0_p & !v230da3e;
assign a04d83 = hbusreq4 & v22fbf21 | !hbusreq4 & v22ef062;
assign v23fb143 = hmaster2_p & v23fba6b | !hmaster2_p & !v191a876;
assign v22fec34 = hgrant3_p & v2305aa9 | !hgrant3_p & v23074aa;
assign v23fc745 = stateG10_5_p & v22ed49b | !stateG10_5_p & v22ef659;
assign v22fd25c = locked_p & v2310c2b | !locked_p & v191a879;
assign v22ff13f = hgrant5_p & v23fb8e3 | !hgrant5_p & v230c03a;
assign v2300ab9 = hmaster2_p & v23fcb55 | !hmaster2_p & v23fcba3;
assign v22ef2aa = hbusreq3 & v22eefcf | !hbusreq3 & v23f36c8;
assign v23f12fa = hbusreq5 & v2306932 | !hbusreq5 & !aa6574;
assign v23f1ccc = hmaster2_p & v231171d | !hmaster2_p & v230de91;
assign v23f9c45 = hgrant1_p & v23f794b | !hgrant1_p & bc5d21;
assign da38b9 = hbusreq0_p & b09503 | !hbusreq0_p & v230a180;
assign v230f2ef = hmaster2_p & v2308d79 | !hmaster2_p & v84561b;
assign v1aadac4 = hgrant1_p & v23f794b | !hgrant1_p & v9ec6b5;
assign v23f3ab8 = jx0_p & v22eea15 | !jx0_p & v2309410;
assign v22ec978 = hmaster0_p & v23135ec | !hmaster0_p & v23fcb3f;
assign v23f6969 = hburst0 & v84561b | !hburst0 & !v23fc8d7;
assign v23fc2b1 = hmaster2_p & v22ffb10 | !hmaster2_p & v84561b;
assign v22ed148 = hbusreq5_p & v23fbaa7 | !hbusreq5_p & v22f53df;
assign v23f4e3d = hbusreq2_p & v22ff123 | !hbusreq2_p & !v845620;
assign v13afe72 = hmaster2_p & v106a782 | !hmaster2_p & v2313463;
assign v23f7b0a = hmaster0_p & v23fc585 | !hmaster0_p & v230774f;
assign v239196f = hmaster0_p & v23fb4ba | !hmaster0_p & v23fb879;
assign v23f8798 = hgrant0_p & v23fcce5 | !hgrant0_p & !v84561b;
assign v23fb80a = stateG10_5_p & v230df30 | !stateG10_5_p & v230bc0c;
assign v22f839c = hmaster0_p & v23fa8d8 | !hmaster0_p & v23f5ba9;
assign v23012e5 = stateG10_5_p & v23022f2 | !stateG10_5_p & !v230320e;
assign v23053bd = hbusreq3_p & v23fc867 | !hbusreq3_p & v84561b;
assign v231345a = hgrant3_p & v84561b | !hgrant3_p & v22f969f;
assign v23fc740 = hbusreq6_p & v22f5272 | !hbusreq6_p & v2308a2f;
assign v23fb1ab = hlock1_p & v23fbae8 | !hlock1_p & v84562b;
assign v22fdd92 = hmaster0_p & v22f654f | !hmaster0_p & v2304432;
assign v23fc790 = hbusreq4 & v22fc0a4 | !hbusreq4 & !v84562a;
assign v23fc624 = hbusreq4 & v23fc8d8 | !hbusreq4 & v23f2bb9;
assign v23fc2fe = hgrant3_p & v230e185 | !hgrant3_p & v23038dd;
assign v22f26d2 = hgrant4_p & v23fbff1 | !hgrant4_p & v23fc5ea;
assign v23113a4 = hbusreq5_p & v84561b | !hbusreq5_p & v22f1389;
assign v23fca5d = hlock1_p & v23f7014 | !hlock1_p & v22ee50f;
assign v23f223a = hbusreq6_p & v2391fc6 | !hbusreq6_p & v230966c;
assign v23934d5 = hbusreq3 & v2312999 | !hbusreq3 & v84561b;
assign v22eec5f = hbusreq5_p & v84561b | !hbusreq5_p & !v22ecc0d;
assign v23f4a48 = hbusreq6 & v15071a6 | !hbusreq6 & v84561b;
assign v22ffea6 = hbusreq3 & v2310389 | !hbusreq3 & v22f61b6;
assign v22f9980 = hbusreq2_p & v191a876 | !hbusreq2_p & v191a879;
assign v23f6865 = hgrant5_p & v230d4f1 | !hgrant5_p & v23f94bc;
assign v2303ebc = hbusreq4 & v2312999 | !hbusreq4 & v84561b;
assign v23fcb1f = hbusreq5_p & v2309c28 | !hbusreq5_p & v23f3dc2;
assign v845641 = hmaster0_p & v84561b | !hmaster0_p & !v84561b;
assign v22f3e94 = hbusreq0 & v22f343b | !hbusreq0 & !v84562a;
assign v2306b0a = hmaster0_p & v22f9403 | !hmaster0_p & !v23fbab9;
assign bfb87c = hmaster2_p & a3cb61 | !hmaster2_p & v23fc716;
assign v23fb5ec = hmaster2_p & v23130a1 | !hmaster2_p & !v22fb272;
assign v22f4e3c = start_p & v84561b | !start_p & v2308b8e;
assign v22f8a0c = hbusreq4_p & a8ec08 | !hbusreq4_p & ad78c9;
assign v22fd6c8 = hmaster2_p & v84562b | !hmaster2_p & v84561b;
assign v22ed1c4 = hbusreq6_p & v230ce2b | !hbusreq6_p & !v84561b;
assign v23fce79 = hlock0_p & v84561b | !hlock0_p & !c16bc3;
assign v8b5388 = hgrant2_p & v84561b | !hgrant2_p & v2307e48;
assign v22ed751 = hbusreq1 & v23fcc10 | !hbusreq1 & v22ff090;
assign v230a241 = hbusreq4_p & v23f8ba7 | !hbusreq4_p & v230f0de;
assign v22eab01 = hbusreq2 & v22fa245 | !hbusreq2 & !v84561b;
assign v230a77a = hmaster1_p & v84561b | !hmaster1_p & !v22f847c;
assign v23f2b6d = hlock1_p & v23f68c1 | !hlock1_p & v2309c93;
assign v8da3ef = hgrant3_p & v22fbd88 | !hgrant3_p & v23f5f94;
assign v23f75db = hlock5_p & v23fca37 | !hlock5_p & v845636;
assign v231072a = hmaster2_p & v2308a71 | !hmaster2_p & v23101b1;
assign v845631 = hbusreq4_p & v84561b | !hbusreq4_p & !v84561b;
assign v22edd64 = hbusreq0 & v22ff090 | !hbusreq0 & v84561b;
assign v23fb0ab = hmaster0_p & v230ad0f | !hmaster0_p & v23fc092;
assign v2304283 = hgrant1_p & a1fba6 | !hgrant1_p & v22fa682;
assign v23084fa = hbusreq3 & v22f3b24 | !hbusreq3 & v84561b;
assign v23fb3f3 = hbusreq4_p & v23f73af | !hbusreq4_p & !v84561b;
assign v23f2daf = hbusreq6 & v22fa0e4 | !hbusreq6 & v84561b;
assign v23104db = jx1_p & v2308f7f | !jx1_p & v23f7456;
assign v87d737 = hbusreq6 & v230af06 | !hbusreq6 & v23fd015;
assign v230ec4b = hgrant6_p & v84561b | !hgrant6_p & v23fcb61;
assign v2300420 = hmaster0_p & v23f78c4 | !hmaster0_p & !v96c563;
assign v2308b8e = stateG3_0_p & v84561b | !stateG3_0_p & !v845665;
assign v23f646e = locked_p & v84561b | !locked_p & !v10dbf64;
assign v23f4254 = hgrant0_p & v23fca61 | !hgrant0_p & v230d2d1;
assign v2305568 = hbusreq1 & v23fc519 | !hbusreq1 & v230f755;
assign v23fcc94 = hmaster1_p & v230e0c0 | !hmaster1_p & v23f42a6;
assign v22ec74f = hmaster1_p & v23f38b1 | !hmaster1_p & v2310c54;
assign v230089c = hgrant3_p & v22f2ca2 | !hgrant3_p & v84561b;
assign v230916d = hlock1_p & v2312526 | !hlock1_p & v23f32a6;
assign v22f62a9 = hbusreq4_p & v22f7347 | !hbusreq4_p & v22f6aa3;
assign v2305bf7 = hbusreq3 & v23f9424 | !hbusreq3 & v23109e5;
assign v22efd33 = hbusreq3 & v23019e9 | !hbusreq3 & v84561b;
assign v22fca36 = hlock3_p & v22f6f5c | !hlock3_p & v23fb81d;
assign v23fc067 = hbusreq4_p & v2392898 | !hbusreq4_p & !v22f3466;
assign v22f6053 = hmaster0_p & b00aa6 | !hmaster0_p & v22ef4de;
assign v23120a3 = hmaster2_p & v23f3978 | !hmaster2_p & v23fb966;
assign v23fc2f3 = hburst0 & v84561b | !hburst0 & !v23fb564;
assign v22f6f5c = hbusreq3_p & v23fa175 | !hbusreq3_p & v84561b;
assign v23083ed = stateG2_p & v22ec1cb | !stateG2_p & v2301d2f;
assign v22ec1c3 = hgrant5_p & v22f65c0 | !hgrant5_p & v239254b;
assign v2304a2d = hlock3_p & v23fcdd8 | !hlock3_p & v2311d6b;
assign v2303634 = hbusreq3_p & v22fba9a | !hbusreq3_p & v23fbcae;
assign v23fbec5 = hmaster2_p & v23fcac2 | !hmaster2_p & v23f3d14;
assign v23927e4 = hbusreq4_p & v22ed335 | !hbusreq4_p & v23fc17c;
assign v23fbda6 = hmastlock_p & v23f8486 | !hmastlock_p & !v84565f;
assign v230580d = hbusreq5_p & v23f5ce0 | !hbusreq5_p & v84561b;
assign v22fd8e1 = hbusreq1_p & v23015be | !hbusreq1_p & v23ef93c;
assign v23fcf45 = jx0_p & v23fcc1e | !jx0_p & !v23f8f24;
assign v230fd1b = hbusreq6_p & v2307aeb | !hbusreq6_p & a1fe5a;
assign v22ec1ae = hmaster2_p & v23fb67c | !hmaster2_p & v23fbeb0;
assign v22ff0ef = hbusreq4_p & v22efe01 | !hbusreq4_p & v23fc349;
assign v23f35c2 = hmaster2_p & v84561b | !hmaster2_p & v94701c;
assign v230a571 = jx0_p & v2307c17 | !jx0_p & v22febf8;
assign v23fc839 = hlock0_p & v845622 | !hlock0_p & v84561b;
assign v2305cac = hmaster2_p & v84561b | !hmaster2_p & v230fec6;
assign v22f0dd3 = hbusreq4_p & v23fc3ca | !hbusreq4_p & v2311668;
assign v23fcdaa = stateA1_p & v84561b | !stateA1_p & !v23fbbb2;
assign v22f9cee = hgrant3_p & v23fbbcb | !hgrant3_p & v23066e8;
assign v23f5907 = hbusreq1_p & v2308d09 | !hbusreq1_p & !v191a876;
assign v23fcaef = hmaster2_p & v23f1a1c | !hmaster2_p & !v2307b06;
assign v230a6ed = hmaster2_p & v22f17bb | !hmaster2_p & v2309c93;
assign v230eb18 = hbusreq5_p & v2303e06 | !hbusreq5_p & v84561b;
assign v22fa7b8 = hlock1_p & b09503 | !hlock1_p & v84561b;
assign v23fcc97 = hmaster1_p & a03e3a | !hmaster1_p & v22f5120;
assign v230ff65 = hmaster0_p & v22f368e | !hmaster0_p & v22f99e9;
assign v2308a2f = hmaster0_p & v230f133 | !hmaster0_p & v1aad535;
assign v230536c = hbusreq2 & v23f5a88 | !hbusreq2 & v84561b;
assign v230d82c = hgrant5_p & v84561b | !hgrant5_p & v23f854f;
assign v22ec686 = hbusreq1_p & v22eb6fc | !hbusreq1_p & v23108aa;
assign v23f4ab4 = hmaster0_p & v23f1ec4 | !hmaster0_p & !v845635;
assign v23fc5c7 = stateG10_5_p & v23f6380 | !stateG10_5_p & v23f4eb4;
assign v230104e = hbusreq1_p & v22fd6a4 | !hbusreq1_p & v84561b;
assign v23f3346 = hmaster2_p & v22fe920 | !hmaster2_p & v22fda59;
assign bd74a3 = hbusreq4_p & v22eaf16 | !hbusreq4_p & v2312290;
assign v2309b80 = hmaster0_p & v23f9fdc | !hmaster0_p & v2310c11;
assign v2312e80 = hbusreq3 & v191b1ba | !hbusreq3 & v22fef65;
assign v22eaafa = hmaster2_p & v23f8da8 | !hmaster2_p & v23fbfd0;
assign v230d5ca = hbusreq4_p & v23fb92f | !hbusreq4_p & v23100e9;
assign v23fbd9b = hlock1_p & v23fc744 | !hlock1_p & v2310c62;
assign v23fc2bf = hbusreq1 & v191a876 | !hbusreq1 & v84561b;
assign v2392d52 = hbusreq5 & v23fc48b | !hbusreq5 & v84561b;
assign v23fc25a = hbusreq6 & v23fbab4 | !hbusreq6 & v84561b;
assign v23fc8ce = hgrant6_p & v23fcd13 | !hgrant6_p & v23f6dfb;
assign v22edb13 = hbusreq5_p & v23126ae | !hbusreq5_p & v2308b98;
assign v23fc7c6 = hlock1_p & b7427f | !hlock1_p & !v84561b;
assign v23f65c8 = hmaster2_p & v230080a | !hmaster2_p & v22f0678;
assign v13aff86 = hmaster2_p & v23fbf8b | !hmaster2_p & !v2312231;
assign v22f96f1 = hbusreq3_p & v23f4dd0 | !hbusreq3_p & v84561b;
assign v2304e69 = hgrant0_p & a1fba6 | !hgrant0_p & v22f19a1;
assign v22fe992 = hlock0_p & v2303978 | !hlock0_p & v84561b;
assign v23f62a3 = hgrant3_p & v22ffa6e | !hgrant3_p & v230468d;
assign v22f2efc = hlock1_p & v23f910c | !hlock1_p & v23f93ee;
assign v22fe165 = hbusreq2 & v2310d44 | !hbusreq2 & !v84561b;
assign v2301cc6 = hgrant1_p & v23f22d2 | !hgrant1_p & v23f2768;
assign v23fca46 = hmaster2_p & v2310a55 | !hmaster2_p & v23f4a07;
assign v230a644 = hmaster2_p & v22fc9bf | !hmaster2_p & !v23929d0;
assign v230e9a6 = stateG10_5_p & v2300c5a | !stateG10_5_p & !v84561b;
assign v22f118f = jx2_p & v23fcaa7 | !jx2_p & v23129fa;
assign v23f58d2 = hlock2_p & v22ebbea | !hlock2_p & v22ee7a7;
assign v22f0af2 = hbusreq1_p & v230a951 | !hbusreq1_p & !v23f4b35;
assign v22f0974 = hmaster0_p & v2305d50 | !hmaster0_p & v22ece29;
assign v239387a = hmaster2_p & v23f55ea | !hmaster2_p & !v22fa5a5;
assign v23fc7a6 = hmaster2_p & v2306d29 | !hmaster2_p & v23f11a3;
assign v22ec616 = hbusreq3_p & v230681b | !hbusreq3_p & v230e874;
assign v230708b = hbusreq5_p & a33e98 | !hbusreq5_p & v845620;
assign af3c3f = hburst0 & v22fdb21 | !hburst0 & !v23f2216;
assign v23fd033 = hbusreq1_p & v23f4426 | !hbusreq1_p & v23f55ea;
assign v22ee524 = hbusreq4_p & v23fc827 | !hbusreq4_p & v22f1498;
assign v2309751 = hmaster0_p & v22ef62d | !hmaster0_p & !v230d854;
assign v2392e6c = hbusreq6 & v230b236 | !hbusreq6 & v84562f;
assign v862ae0 = hlock0_p & v2305fe0 | !hlock0_p & v84564d;
assign v22f0860 = hbusreq2 & v23fbbd2 | !hbusreq2 & !v84561b;
assign v23fbd51 = hmaster1_p & v22f7fc1 | !hmaster1_p & v23fbc46;
assign v23fc5a0 = hgrant3_p & v22efef6 | !hgrant3_p & v23fcb36;
assign v22ee750 = hgrant2_p & v2307ff5 | !hgrant2_p & v22eb1f5;
assign v22f21bd = hmaster2_p & v23fba25 | !hmaster2_p & v23f471a;
assign v23fb487 = hmaster2_p & v84561b | !hmaster2_p & v2307c5d;
assign v23f03d2 = hbusreq3_p & v2311d04 | !hbusreq3_p & v23fb667;
assign v22f380e = hgrant2_p & v2307e48 | !hgrant2_p & v84561b;
assign v2303831 = hbusreq2 & v23f8f21 | !hbusreq2 & v84561b;
assign v23916c0 = hgrant5_p & v22eedd0 | !hgrant5_p & v22f6a0e;
assign v23091d2 = hmaster1_p & v22ef354 | !hmaster1_p & v23128f3;
assign v22f4f0f = hbusreq4_p & v84564d | !hbusreq4_p & !v84561b;
assign v230a226 = hbusreq3 & v845620 | !hbusreq3 & v84561b;
assign v230a671 = hlock0_p & v84561b | !hlock0_p & !v23fc18a;
assign v23fcab1 = hgrant3_p & v23f1c14 | !hgrant3_p & v23f292d;
assign v22f2639 = hlock0_p & v845622 | !hlock0_p & v22fadb0;
assign v23099de = hbusreq0 & v22fca61 | !hbusreq0 & v84561b;
assign v23002d1 = hmaster2_p & a1fbb6 | !hmaster2_p & v22f4f42;
assign bf150c = hmaster0_p & v22f368e | !hmaster0_p & v230d8af;
assign v22f12c8 = hbusreq1 & v230a753 | !hbusreq1 & v22f64de;
assign v23fc6be = hbusreq6_p & v230f8f4 | !hbusreq6_p & v23fb8c9;
assign v22fe924 = hbusreq3_p & v23934d5 | !hbusreq3_p & v1aad323;
assign v23fc411 = hlock2_p & b9d00f | !hlock2_p & a1fbb6;
assign v23fb58e = hbusreq4 & v2308a7d | !hbusreq4 & v23f1391;
assign v23fc23a = hbusreq3_p & v23f8895 | !hbusreq3_p & v23f3a5b;
assign v22f7d4e = hlock0_p & v22ecc15 | !hlock0_p & v23fca2d;
assign v23fcb5d = stateA1_p & v84561b | !stateA1_p & !v2306775;
assign v23f6fe7 = hbusreq4_p & v23fc2da | !hbusreq4_p & fc894d;
assign v22ec0f7 = hbusreq3_p & v22f679a | !hbusreq3_p & v230c499;
assign v22ed7ba = hbusreq1_p & v2307a6d | !hbusreq1_p & !v84561b;
assign v23f0eec = hmaster2_p & v191aa68 | !hmaster2_p & v22ecc15;
assign v9c8a7f = hbusreq3 & v23fc6ef | !hbusreq3 & v23fbec5;
assign v22eb5b3 = hlock0_p & v191a86f | !hlock0_p & v23fb8bf;
assign v23fb8fb = jx1_p & v23089cd | !jx1_p & !v22ede66;
assign v23f7de2 = hgrant5_p & v23003fc | !hgrant5_p & v23fc5fe;
assign fc894d = hmaster0_p & v2307fee | !hmaster0_p & v23fc4e7;
assign v23f8d36 = hmaster0_p & v22f4ef0 | !hmaster0_p & v2393495;
assign v23f79f6 = hgrant1_p & v22f8593 | !hgrant1_p & v23fc6d6;
assign v22fa502 = hmaster0_p & v2302831 | !hmaster0_p & v23f353e;
assign v22f4998 = hgrant1_p & v84561b | !hgrant1_p & v22f8da5;
assign v23fb1c0 = hmaster0_p & v230d25d | !hmaster0_p & v23f7997;
assign v22f53d4 = hlock1_p & v23f2713 | !hlock1_p & v845620;
assign v90eab4 = hmaster0_p & v22f368e | !hmaster0_p & v22f317b;
assign v23f96b7 = hbusreq6_p & v2303e0d | !hbusreq6_p & v23f7b94;
assign v2392cce = hmaster0_p & v23fc50a | !hmaster0_p & !v23fc00b;
assign v22edc69 = hmaster0_p & v23fb7c3 | !hmaster0_p & !v2309d23;
assign v22eef3f = hlock3_p & v917514 | !hlock3_p & v9eaa59;
assign v22ef4f0 = hmaster2_p & v23fcc3c | !hmaster2_p & v23f9dd1;
assign v23026db = stateG2_p & v84561b | !stateG2_p & v15071da;
assign v191ae28 = hlock5_p & v22fd6ba | !hlock5_p & v230b04e;
assign v23fa8aa = hbusreq2_p & v22f5037 | !hbusreq2_p & !v84561b;
assign v23fb7fc = hgrant1_p & v84564d | !hgrant1_p & !v22fe495;
assign v23fc02b = hmaster2_p & v23fc514 | !hmaster2_p & v22f163a;
assign b0fad6 = hlock4 & v22feb5c | !hlock4 & v22f24ca;
assign v23fbd91 = hgrant6_p & v2306cad | !hgrant6_p & v1e841ad;
assign v230ed07 = jx1_p & v85e5cf | !jx1_p & !v2307479;
assign v22f1682 = hbusreq0_p & v22f1b4e | !hbusreq0_p & v22ed7a8;
assign v230e115 = hmaster2_p & v23102d5 | !hmaster2_p & v22f94ec;
assign v23f6a95 = hgrant3_p & v84561b | !hgrant3_p & v22f483c;
assign v13afe8f = hmastlock_p & v23fb564 | !hmastlock_p & v84561b;
assign v23fc008 = hbusreq6 & v23fc192 | !hbusreq6 & v84561b;
assign v22f0538 = hmaster2_p & v23fb8a2 | !hmaster2_p & v22f3aa1;
assign v230e40c = hmaster0_p & v2306fba | !hmaster0_p & v22ee47d;
assign v23fc56a = hlock3_p & v2306837 | !hlock3_p & v22f71ee;
assign v2309515 = hbusreq2 & v106ae21 | !hbusreq2 & v84564d;
assign v2305b58 = hbusreq3 & v22edfa7 | !hbusreq3 & v84561b;
assign v23f8884 = hgrant5_p & v2308c0b | !hgrant5_p & v22f33d3;
assign v22f5120 = hbusreq6_p & v23fcf9e | !hbusreq6_p & v2392fa6;
assign v2302844 = hmaster0_p & v23f8a43 | !hmaster0_p & v2392f25;
assign v23fbc9c = hmaster0_p & v23fa3b8 | !hmaster0_p & v23fb5a7;
assign v22fc745 = hlock5_p & v15071f0 | !hlock5_p & v84562b;
assign v22f0d28 = hmaster0_p & v22fd152 | !hmaster0_p & v22ef5cd;
assign v23f9a3a = hbusreq6_p & v2302b81 | !hbusreq6_p & v22f0fcd;
assign v23025d8 = hmaster2_p & v2311606 | !hmaster2_p & v22ffff6;
assign v23fcdd7 = hbusreq1_p & v2306538 | !hbusreq1_p & v22f8c0b;
assign v23f5b67 = hmaster0_p & v1aad34c | !hmaster0_p & v22f32b9;
assign v230ef5e = hbusreq5_p & v22f985c | !hbusreq5_p & v845620;
assign v22ebd1b = hbusreq6 & v22eb60c | !hbusreq6 & v22ef062;
assign v23f0cce = hmaster2_p & v13afe3a | !hmaster2_p & v23f34d4;
assign v23fb527 = hbusreq5_p & v97b973 | !hbusreq5_p & v84561b;
assign v23fb7ea = hmaster0_p & v22eb22e | !hmaster0_p & !a1fd0e;
assign v230b30c = jx0_p & v2306967 | !jx0_p & v2387c0f;
assign v23fbb77 = hmaster0_p & v23fcea2 | !hmaster0_p & !v23fcc11;
assign v23f7e43 = hbusreq2_p & v22f47b0 | !hbusreq2_p & v84561b;
assign v23fc3ee = hgrant5_p & v84561b | !hgrant5_p & !v230848d;
assign v22fc67e = hmaster0_p & v2301be6 | !hmaster0_p & v22f2849;
assign v23fc94d = hmaster0_p & v2306593 | !hmaster0_p & v22f6ae5;
assign v2302a57 = jx1_p & v23132e5 | !jx1_p & v23108bb;
assign v23fce31 = hmaster2_p & v84561b | !hmaster2_p & !v23fbc48;
assign v23fcab4 = hmaster1_p & v23fcb62 | !hmaster1_p & v22ef962;
assign v22ef751 = hbusreq2_p & v22f3643 | !hbusreq2_p & !v84561b;
assign v22fa9be = hbusreq0 & v23fbfd0 | !hbusreq0 & v84561b;
assign v22f8291 = hmaster1_p & v22fcab7 | !hmaster1_p & v23f594f;
assign v23fc982 = hbusreq1_p & v23f1228 | !hbusreq1_p & v22eb05f;
assign v23fbcad = hmaster2_p & v22f60c6 | !hmaster2_p & v84564d;
assign v23fbeae = hbusreq4_p & v23f7fe8 | !hbusreq4_p & v23125ab;
assign v23f0ba3 = hbusreq3 & v23efb4d | !hbusreq3 & v22f54cb;
assign v23f3e19 = stateG10_5_p & v238b0d7 | !stateG10_5_p & v230fec6;
assign v23086c5 = hgrant5_p & v84561b | !hgrant5_p & v2393900;
assign v1507437 = hmaster0_p & v23f3955 | !hmaster0_p & v230389f;
assign v23fb936 = hbusreq6_p & v22fbfe3 | !hbusreq6_p & v230bf1e;
assign v23f2324 = hbusreq5 & v23fbfd0 | !hbusreq5 & v23fce71;
assign v230a2c7 = hgrant1_p & v23fbaac | !hgrant1_p & v23f50bb;
assign v23fcb0e = hbusreq6_p & v9bcd2e | !hbusreq6_p & v23008a1;
assign v23094c7 = hmaster0_p & v23f6ad0 | !hmaster0_p & v23fbe50;
assign v23fc815 = hgrant3_p & v230d8af | !hgrant3_p & v23f2504;
assign v2308be5 = hlock0_p & v23f7218 | !hlock0_p & v2308d66;
assign v22fdd65 = hbusreq3_p & v23fc7ab | !hbusreq3_p & v23fba9a;
assign v2306e8f = hmaster2_p & v84561b | !hmaster2_p & v23f745f;
assign v22f05f3 = hbusreq5_p & v22f004e | !hbusreq5_p & !v84561b;
assign v23f5218 = hbusreq5_p & v2301655 | !hbusreq5_p & v23f366d;
assign v2303978 = hbusreq0 & v23f7218 | !hbusreq0 & v84561b;
assign v230c727 = hgrant1_p & v23126ae | !hgrant1_p & v22f79be;
assign v1aadb95 = hgrant2_p & a1fba6 | !hgrant2_p & v9526ac;
assign e1deb1 = hmaster0_p & v23f4338 | !hmaster0_p & v23fc0a5;
assign v23f5500 = hmaster1_p & v23f3c98 | !hmaster1_p & !v22fd15a;
assign v22f3a11 = hgrant0_p & v845622 | !hgrant0_p & v191accc;
assign e1e659 = hmaster2_p & v22f995e | !hmaster2_p & v22ee06a;
assign v23fba62 = hbusreq3_p & v230a6ed | !hbusreq3_p & v230f9f1;
assign v22fca64 = hlock4_p & v22fbbd0 | !hlock4_p & v23f273b;
assign v23fcbb0 = hlock6_p & v23fc684 | !hlock6_p & v84561b;
assign v2310a40 = hbusreq5 & v23022b1 | !hbusreq5 & !v84561b;
assign f40a8f = hbusreq3_p & v2303bfd | !hbusreq3_p & v22fb592;
assign a20348 = hgrant3_p & v84562e | !hgrant3_p & v2308b2e;
assign v23fcff6 = hmaster2_p & v22f220a | !hmaster2_p & v23129e0;
assign v23fc706 = stateG10_5_p & v84561b | !stateG10_5_p & !v106a782;
assign v23f1ca8 = hgrant0_p & v230eb9b | !hgrant0_p & v23fa8bb;
assign v230313a = hgrant1_p & a1fbc2 | !hgrant1_p & v23f8825;
assign v23fccc2 = hbusreq6 & v23fba11 | !hbusreq6 & v230cb63;
assign v23fc4dd = jx1_p & v2312524 | !jx1_p & v84561b;
assign v230774f = hbusreq4 & v12cd4f6 | !hbusreq4 & v23fa392;
assign v230e50f = jx0_p & v23fc588 | !jx0_p & v22f1154;
assign v2391d99 = hmaster2_p & v230c727 | !hmaster2_p & a88394;
assign v23f8a36 = hgrant5_p & v84561b | !hgrant5_p & v230db01;
assign v231024c = hbusreq4 & v23f8561 | !hbusreq4 & v84561b;
assign v230c499 = hmaster2_p & b10190 | !hmaster2_p & v23fc957;
assign v22f0945 = hbusreq5 & v845620 | !hbusreq5 & v84561b;
assign v23fbf0e = hmaster2_p & v23f4808 | !hmaster2_p & v23fbfa7;
assign v23fc6d3 = hbusreq1 & v2302048 | !hbusreq1 & v84561b;
assign v22f9b6f = hmaster2_p & v84561b | !hmaster2_p & !v22f49ac;
assign v23fcb1a = hgrant1_p & v84561b | !hgrant1_p & v23fcdd9;
assign v2302907 = hbusreq6 & v23f4fa4 | !hbusreq6 & !v22ff914;
assign v2309310 = hbusreq2 & v22f50bf | !hbusreq2 & v84561b;
assign v23fc778 = hlock1_p & v23fc823 | !hlock1_p & !v84561b;
assign v22f549a = stateG10_5_p & v230d16b | !stateG10_5_p & v2392534;
assign v23f9fc1 = hbusreq5_p & v2391a57 | !hbusreq5_p & !v84561b;
assign v23011cb = locked_p & v23efa52 | !locked_p & v84561b;
assign v22f115b = hbusreq1 & v23fb9c2 | !hbusreq1 & v84564d;
assign v23fc14e = hbusreq0 & v22ffea0 | !hbusreq0 & !v22f4527;
assign v23fc46b = hbusreq5_p & v13afe3a | !hbusreq5_p & v845647;
assign v22eb6ca = hmaster0_p & v22ef62d | !hmaster0_p & v230880f;
assign v23fc514 = hmastlock_p & a1fd35 | !hmastlock_p & !v84561b;
assign v23fbadb = hmaster2_p & v23f5fb5 | !hmaster2_p & v84561b;
assign v22f3091 = hbusreq3_p & v22f3628 | !hbusreq3_p & v84561b;
assign v2308d9e = hbusreq4 & v2301044 | !hbusreq4 & !v23fbeeb;
assign v95ca19 = hbusreq6_p & v23fba71 | !hbusreq6_p & v84561b;
assign v12cd4c6 = hlock0_p & v84562b | !hlock0_p & v23fbab2;
assign v23121b5 = hbusreq5 & v23f4ca0 | !hbusreq5 & v84561b;
assign v230ed7d = hbusreq4 & v23fca95 | !hbusreq4 & v23fc034;
assign v22fe58b = hlock3_p & v23f4861 | !hlock3_p & v23fb9a7;
assign v1506f02 = hbusreq1 & v23f8a9d | !hbusreq1 & v84561b;
assign v230b08d = hgrant3_p & v84561b | !hgrant3_p & bd761f;
assign c17224 = jx1_p & v2308fb4 | !jx1_p & v1aae5da;
assign v22f00b6 = hbusreq6_p & v231170f | !hbusreq6_p & !v230889a;
assign v23fbc40 = hbusreq3 & v84561b | !hbusreq3 & v23051cf;
assign v23fc47e = hbusreq2_p & v23fcc09 | !hbusreq2_p & v845620;
assign v23faf8a = hgrant0_p & v2312f3c | !hgrant0_p & v23f0652;
assign v230df44 = hmaster2_p & v22f7808 | !hmaster2_p & v2309729;
assign v22f2e61 = hbusreq3_p & v22ebccd | !hbusreq3_p & !v84561b;
assign v23fa175 = hbusreq3 & v23fccd6 | !hbusreq3 & v84561b;
assign v22edaad = hbusreq5_p & v22f39af | !hbusreq5_p & v22f1bec;
assign v22feb39 = jx1_p & v23125e2 | !jx1_p & v23fce7a;
assign bfba4f = jx0_p & v23fbced | !jx0_p & v2307ab6;
assign v23f9f89 = hmaster2_p & v2312990 | !hmaster2_p & v84561b;
assign v2305c74 = hmaster1_p & v23fbec3 | !hmaster1_p & v23f3166;
assign v23114d2 = hgrant1_p & v84561b | !hgrant1_p & v22ef769;
assign v230efa0 = jx0_p & v230ba49 | !jx0_p & v23fc917;
assign v230502a = hlock3_p & v23fbbf0 | !hlock3_p & v2302d3c;
assign v23f6077 = hbusreq0 & v22f3643 | !hbusreq0 & v845620;
assign v22f6ee2 = hlock1_p & v230a9eb | !hlock1_p & !v12cd3f4;
assign v15072b7 = hmaster2_p & v23fcd0f | !hmaster2_p & v22fba03;
assign v22eb58b = hmaster0_p & v23fceb8 | !hmaster0_p & v22fa080;
assign v2302e76 = hbusreq2_p & v22ede4d | !hbusreq2_p & v84561b;
assign v22fffa6 = hbusreq6 & v22fccd1 | !hbusreq6 & v22f9bc8;
assign v22eebd6 = hlock4_p & v22ebe20 | !hlock4_p & v22ef242;
assign v23fc8eb = hgrant0_p & v84561b | !hgrant0_p & v23fcff1;
assign v230a6a7 = hbusreq2 & v84562b | !hbusreq2 & !v84561b;
assign v2393723 = hlock0_p & v23f1e72 | !hlock0_p & v845620;
assign v22f923c = hgrant5_p & v22fb403 | !hgrant5_p & v22f3a11;
assign v230daec = hbusreq6_p & v23131fd | !hbusreq6_p & v84561b;
assign b355fd = hmaster0_p & v191b037 | !hmaster0_p & v23f99ec;
assign v23f55fb = hlock6_p & v22fe816 | !hlock6_p & v22ff400;
assign v22ff9d9 = hbusreq5_p & v230f63f | !hbusreq5_p & v22f9c42;
assign v230360b = hbusreq5 & v22fda32 | !hbusreq5 & v23fa2ec;
assign v23fc8b8 = hmaster1_p & v23fbe69 | !hmaster1_p & v230d5ca;
assign v2392897 = stateG2_p & v2302ca3 | !stateG2_p & v22ef867;
assign v22eb856 = hmaster0_p & v230eeb6 | !hmaster0_p & v22fb6df;
assign v2307a27 = hbusreq0 & v22ed6c5 | !hbusreq0 & v84564d;
assign v22f8d74 = hready & v22f5eee | !hready & v22febb1;
assign v22fa4b4 = hbusreq5 & v1aae362 | !hbusreq5 & !v84561b;
assign v84562d = hbusreq3_p & v84561b | !hbusreq3_p & !v84561b;
assign v1aad5ee = hmaster0_p & v23f48a1 | !hmaster0_p & v2391e5e;
assign v22f53c0 = hgrant1_p & v230f9db | !hgrant1_p & v22f2e82;
assign v23fb1b9 = hbusreq3 & v230a83f | !hbusreq3 & v84561b;
assign v23f7e3d = hbusreq3_p & v23f8efa | !hbusreq3_p & v23f57c1;
assign v23f00ec = hgrant5_p & v12cda32 | !hgrant5_p & v22efa67;
assign v2312ef7 = hmaster2_p & v230a035 | !hmaster2_p & v84561b;
assign v23fcb02 = hlock6_p & v23f58a6 | !hlock6_p & v22fdd61;
assign v22f1a8f = hlock6 & v22feb5c | !hlock6 & v22f7fcc;
assign v23117c1 = hmaster2_p & v191a876 | !hmaster2_p & !v22eb5b3;
assign v23f022d = hbusreq2_p & v22fe165 | !hbusreq2_p & !v84561b;
assign v22f35fa = hlock0_p & v2307e4f | !hlock0_p & v845620;
assign v230f27a = hgrant3_p & v230b38b | !hgrant3_p & v230074c;
assign v23071cd = hmaster2_p & v22ed85a | !hmaster2_p & v23003cc;
assign v23fc153 = hgrant0_p & v2310a7e | !hgrant0_p & v23fceb9;
assign v23fb0d9 = hmaster2_p & v2392ece | !hmaster2_p & v22f7b8b;
assign v23fc478 = hbusreq6 & v23f15ac | !hbusreq6 & v84561b;
assign v1b876be = hbusreq4 & v22f2e92 | !hbusreq4 & v22fd1a7;
assign v230d4f1 = hbusreq5_p & v23126ae | !hbusreq5_p & v23fc004;
assign v23fc336 = hbusreq5_p & v23065ad | !hbusreq5_p & v23fc207;
assign v23fbe38 = hlock6_p & v22f0cf9 | !hlock6_p & v23fb657;
assign v23fbb55 = hbusreq3 & v22fb1f3 | !hbusreq3 & v84561b;
assign v23fc1c1 = hgrant2_p & v2310116 | !hgrant2_p & v23fb920;
assign v23919c0 = hmaster2_p & v91c376 | !hmaster2_p & v22fd69b;
assign v230c480 = hmaster2_p & v23102d5 | !hmaster2_p & v13afc17;
assign v22fe5f9 = hmaster2_p & v23fb49a | !hmaster2_p & v22f893a;
assign v23f93b5 = hbusreq6 & v23fc546 | !hbusreq6 & v84561b;
assign v2306b9f = hmaster2_p & v23fb796 | !hmaster2_p & !v23fbf53;
assign v22f8943 = hbusreq5_p & v23fc393 | !hbusreq5_p & v230354e;
assign v22f764d = hmaster2_p & v23f40d6 | !hmaster2_p & v23109fb;
assign v22fa646 = hbusreq3_p & v84561b | !hbusreq3_p & v23fc957;
assign v230ab72 = hbusreq4 & v23fc068 | !hbusreq4 & !v84561b;
assign v2310c62 = hbusreq1 & v23fcc10 | !hbusreq1 & v84561b;
assign v23fc75d = hbusreq3_p & v84561b | !hbusreq3_p & v230f9db;
assign v23fc43e = hlock3_p & ba4552 | !hlock3_p & v230a226;
assign v23f30cf = hmaster2_p & v1506fbf | !hmaster2_p & v84561b;
assign v22f6f8f = hbusreq0_p & v84561b | !hbusreq0_p & !v106a782;
assign v22ecc3f = hbusreq0_p & v2306d29 | !hbusreq0_p & v22fdc30;
assign v22fef02 = hlock0_p & v84564d | !hlock0_p & v23fcc5a;
assign v2392f11 = hbusreq3 & v1506ff4 | !hbusreq3 & v84561b;
assign v22fd532 = hbusreq6_p & v22f11cc | !hbusreq6_p & v2310934;
assign v231050f = hbusreq5_p & v22f3999 | !hbusreq5_p & e1beab;
assign v23030e8 = hgrant0_p & v84561b | !hgrant0_p & v22f3813;
assign v23f4cb5 = hlock1_p & v23fbb95 | !hlock1_p & v845620;
assign v23fbb83 = hmaster0_p & v892c49 | !hmaster0_p & v23fc293;
assign v23fc3da = hbusreq3_p & v23fc541 | !hbusreq3_p & v230e75b;
assign v23f15e7 = hmaster0_p & v1aae2a5 | !hmaster0_p & v22f4abc;
assign v23fca89 = hbusreq6 & v23f73dd | !hbusreq6 & v84561b;
assign v22fd794 = hbusreq0_p & v23fd040 | !hbusreq0_p & v2301b2d;
assign v22f04b5 = hbusreq4_p & v22ff3c3 | !hbusreq4_p & v22ec8dc;
assign v23fcfbb = hbusreq1_p & v23fc1f0 | !hbusreq1_p & v84561b;
assign v230251b = hmaster2_p & v845620 | !hmaster2_p & v230984f;
assign v2310bdf = hlock0_p & v22fe19b | !hlock0_p & !v84561b;
assign v230efe0 = hgrant3_p & v22ffa6e | !hgrant3_p & v22f39d3;
assign v23fb4bd = hgrant0_p & v22eaafd | !hgrant0_p & v230158e;
assign v230dcf6 = hmaster2_p & v191a86f | !hmaster2_p & v191ae42;
assign v22fef21 = jx1_p & v230e534 | !jx1_p & v22fca63;
assign v23fcf51 = hbusreq4 & v23fc6ce | !hbusreq4 & v22f2623;
assign v22eb6ba = hgrant1_p & v22f95c8 | !hgrant1_p & v23fc96e;
assign v23127ee = hgrant3_p & v84562d | !hgrant3_p & v22f5136;
assign v2310256 = hmaster2_p & v2312c13 | !hmaster2_p & !b9d013;
assign v23fbf73 = jx0_p & v22f4b6d | !jx0_p & v84561b;
assign v22f8e09 = hbusreq3 & v22ef350 | !hbusreq3 & v22fd6c0;
assign v191a909 = hmaster0_p & v23f3955 | !hmaster0_p & v230379f;
assign v23f4cfb = hmaster2_p & v23f9226 | !hmaster2_p & v22efa93;
assign v8fafbf = hbusreq6 & v2305e79 | !hbusreq6 & !v22eb3e5;
assign v230bb30 = stateG10_5_p & v230bc0c | !stateG10_5_p & v2301f52;
assign v191abfa = hmaster0_p & v84564d | !hmaster0_p & v2305252;
assign v22ff3c3 = hmaster0_p & v22ff30c | !hmaster0_p & v22fec34;
assign v22ef44c = hmaster0_p & v23fca89 | !hmaster0_p & v2301adf;
assign v2304b1d = hmaster2_p & v23fc2ce | !hmaster2_p & !v106ae19;
assign bd8ccb = hgrant3_p & v22f789c | !hgrant3_p & a0b7a3;
assign b1e9fa = hmaster0_p & v23fc3aa | !hmaster0_p & !v23fc372;
assign v230c3d2 = hmaster0_p & v23f3b8f | !hmaster0_p & v2312be0;
assign v23122fa = hmaster0_p & v23fcd2a | !hmaster0_p & !v23008f3;
assign v22ed8bc = hbusreq3_p & v23f6769 | !hbusreq3_p & v84561b;
assign v23fc74f = hbusreq5_p & v106af73 | !hbusreq5_p & v23fc004;
assign v23fcfb4 = hmaster2_p & v1aae98c | !hmaster2_p & v22fda32;
assign v23f5066 = hbusreq3_p & v230200a | !hbusreq3_p & v2300362;
assign f40761 = hlock5_p & v22ffbb3 | !hlock5_p & !v230f848;
assign v22f9b0c = hbusreq3_p & a83396 | !hbusreq3_p & v84561b;
assign v23027c2 = hbusreq1 & v22fc723 | !hbusreq1 & v22fe657;
assign v2302608 = jx1_p & v22ed4ea | !jx1_p & v23f8095;
assign v22ebbf1 = hgrant1_p & v12cd6a1 | !hgrant1_p & v23fc9c8;
assign v23fb5d1 = hbusreq1_p & v22fead6 | !hbusreq1_p & v22f5734;
assign v23fc65d = hmaster2_p & v191aa68 | !hmaster2_p & v22f35e8;
assign v22eddfd = hbusreq6_p & v23fc2ff | !hbusreq6_p & v1aad4b7;
assign v2312a52 = hgrant3_p & v84562d | !hgrant3_p & v22fe2d5;
assign v23f619d = hmaster0_p & v230cea0 | !hmaster0_p & v1e84190;
assign v1aae9dc = jx0_p & v1aae6ba | !jx0_p & v230e991;
assign v23017b3 = hmaster1_p & v2306291 | !hmaster1_p & v23fcc82;
assign v22ee884 = hlock1_p & v23fb743 | !hlock1_p & v22f7b83;
assign v12cd632 = hlock6_p & v22f1d08 | !hlock6_p & v22f968e;
assign v2309b0f = hlock0_p & v23f5af5 | !hlock0_p & !v2309c8a;
assign v230e651 = hbusreq5 & v22ebbea | !hbusreq5 & !v84561b;
assign v2304e51 = hbusreq4_p & v230ae14 | !hbusreq4_p & v2312ba0;
assign v23081f5 = hbusreq0_p & v23056b1 | !hbusreq0_p & v23f86f0;
assign v2304924 = hmaster2_p & v23035d7 | !hmaster2_p & v23f0d46;
assign v23f525c = hgrant3_p & v230b199 | !hgrant3_p & v22f2d7c;
assign v13afc0b = hbusreq3 & v23fc089 | !hbusreq3 & v23fbf0b;
assign v22f8b01 = hgrant1_p & v23f87f4 | !hgrant1_p & v23fa997;
assign v22ef0b4 = hmaster2_p & v22f1244 | !hmaster2_p & v2310fcd;
assign e1e78b = hgrant4_p & v84561b | !hgrant4_p & v845631;
assign v23fc612 = hgrant0_p & a07f9b | !hgrant0_p & v23fcf8f;
assign v2303f7c = hbusreq3 & v23f9aa8 | !hbusreq3 & v2310d04;
assign v22f9b00 = hbusreq3_p & v23fba07 | !hbusreq3_p & v84561b;
assign v2393739 = hlock1_p & v22ede4d | !hlock1_p & v84561b;
assign v150745f = hlock5_p & v22f621f | !hlock5_p & v845636;
assign v22f6955 = hgrant4_p & v23f1925 | !hgrant4_p & v230d82a;
assign v23119a8 = hmaster2_p & v84561b | !hmaster2_p & !v23f0865;
assign v22fe346 = hgrant1_p & v845626 | !hgrant1_p & v23f8a99;
assign v2302b93 = hmaster0_p & v22ec354 | !hmaster0_p & !v22fa6f5;
assign v23fc757 = hbusreq1_p & v2306d29 | !hbusreq1_p & v23126ae;
assign v2308225 = hbusreq2_p & v23fb11d | !hbusreq2_p & v84561b;
assign v23f7499 = hgrant0_p & v84561b | !hgrant0_p & v22f49e4;
assign v230ad5b = hgrant2_p & v2312283 | !hgrant2_p & !v23fc7dd;
assign bd7476 = hbusreq5_p & v230446f | !hbusreq5_p & !v23f366d;
assign v23fce9a = hlock3_p & v23fca78 | !hlock3_p & v23fcfe4;
assign v23fc9e5 = hbusreq3_p & v23fccb0 | !hbusreq3_p & v1506add;
assign v22ede6c = hbusreq3_p & v22fc963 | !hbusreq3_p & v230e635;
assign v23f9319 = hbusreq3 & v23056bc | !hbusreq3 & v84561b;
assign v23f1263 = hgrant3_p & v230727f | !hgrant3_p & v23fbe3a;
assign c16602 = hmaster1_p & v23fbf16 | !hmaster1_p & v23f2041;
assign v22f6721 = hbusreq3_p & v230dfff | !hbusreq3_p & e1e659;
assign v230646f = hbusreq3_p & v230d0a3 | !hbusreq3_p & v84561b;
assign v23fb93c = hbusreq3_p & v230fb0a | !hbusreq3_p & v23f660f;
assign v23f6532 = hmaster0_p & v231398c | !hmaster0_p & v230efe0;
assign a07f9b = locked_p & v23fcad0 | !locked_p & a1fba6;
assign e1de6f = hbusreq6 & v2310d2f | !hbusreq6 & v84562f;
assign v22f7728 = hbusreq6_p & v10dbf63 | !hbusreq6_p & !v84561b;
assign v2306660 = hmaster2_p & v22ed7a8 | !hmaster2_p & v230a9eb;
assign v23fc781 = hmaster1_p & v230bdd4 | !hmaster1_p & v84561b;
assign v23126b8 = hmaster2_p & v22fc8c8 | !hmaster2_p & v84561b;
assign v2391a43 = stateG10_5_p & v22f96f2 | !stateG10_5_p & v23035ba;
assign v23f13f3 = hbusreq3_p & v2307701 | !hbusreq3_p & v23f9a56;
assign v22ff9d4 = hmaster2_p & v84561b | !hmaster2_p & !v23f9dd1;
assign v22f6611 = hmaster2_p & b9d049 | !hmaster2_p & v84561b;
assign v23fb8c0 = stateA1_p & v23fceb3 | !stateA1_p & v23fbbb2;
assign v23fbe15 = hbusreq4 & v23fbdf9 | !hbusreq4 & v84561b;
assign v22fc5d2 = hmaster2_p & v191aa68 | !hmaster2_p & v23041e2;
assign v23fc081 = hmaster0_p & v23081e8 | !hmaster0_p & v2308e49;
assign v23fccfd = jx0_p & v22eb015 | !jx0_p & v2303efa;
assign v22f2e41 = hmaster2_p & v9d8aae | !hmaster2_p & v23131e8;
assign v991952 = hmaster2_p & v22ebca0 | !hmaster2_p & v23fb624;
assign v23133be = hbusreq4_p & v230cd17 | !hbusreq4_p & v84561b;
assign v23fa966 = hmaster1_p & v23f5983 | !hmaster1_p & v2311f82;
assign v23f8692 = hmaster0_p & v23fbf3f | !hmaster0_p & !v22f1b30;
assign v22fa88a = hbusreq5_p & v84561b | !hbusreq5_p & v23f614a;
assign b15ae7 = hmaster0_p & v22f1d6c | !hmaster0_p & v23076e7;
assign v22f160c = hgrant3_p & v84562e | !hgrant3_p & v23fb624;
assign aa6574 = hbusreq0 & v23fbbd2 | !hbusreq0 & !v84561b;
assign v23f699c = hgrant4_p & v23055b0 | !hgrant4_p & v23119a4;
assign v23fc6ef = hmaster2_p & v23fcac2 | !hmaster2_p & v22ee9be;
assign v23fc16f = hbusreq6_p & v22eaf16 | !hbusreq6_p & bd74a3;
assign v13aff30 = hbusreq5 & v230d16b | !hbusreq5 & v84561b;
assign v230e2d4 = hbusreq3 & v22ed533 | !hbusreq3 & v23f9f89;
assign v23f363f = hmaster2_p & v22f1a26 | !hmaster2_p & v2301e25;
assign v22f3fec = hbusreq5_p & v1506ffd | !hbusreq5_p & !v84561b;
assign v22f36ba = hlock0_p & v2307a27 | !hlock0_p & v2301aab;
assign v23f97c6 = hgrant3_p & v22fe370 | !hgrant3_p & !v22f9801;
assign v23085df = stateG2_p & v23fc331 | !stateG2_p & v22ff64f;
assign v23f7ffc = hbusreq0_p & v22f8d2b | !hbusreq0_p & v22eddb2;
assign a72160 = hmastlock_p & v22fb427 | !hmastlock_p & v84561b;
assign v23fb5d6 = hgrant1_p & v84561b | !hgrant1_p & v23f307c;
assign v2301505 = hbusreq2_p & v23fced7 | !hbusreq2_p & v845620;
assign v23004ba = hmaster1_p & v22f2965 | !hmaster1_p & bee61a;
assign v2305af1 = hlock5_p & v22f5d49 | !hlock5_p & bbc337;
assign v230f105 = hgrant5_p & v22ee495 | !hgrant5_p & v22fa20a;
assign v230ef73 = hbusreq3_p & v2300362 | !hbusreq3_p & v23025e4;
assign v23087e8 = hbusreq3 & v23fbb5a | !hbusreq3 & v845622;
assign v2301135 = hmaster0_p & v23fbad4 | !hmaster0_p & v22ef7a5;
assign v23fbe8f = hbusreq6_p & v22f5d45 | !hbusreq6_p & v23fc76e;
assign v2308d51 = hgrant1_p & v84561b | !hgrant1_p & v23fcddb;
assign v23f69ba = hbusreq0 & v191a876 | !hbusreq0 & !v84561b;
assign v230e4c7 = hmaster1_p & v22fa6c0 | !hmaster1_p & v2307c9a;
assign v2312ebb = hmaster0_p & v23fc3aa | !hmaster0_p & !v23068f2;
assign v23fccd4 = hbusreq3 & v22eef66 | !hbusreq3 & !v23f089b;
assign bd762f = hmaster2_p & v22f1244 | !hmaster2_p & v23fafc5;
assign v23052c9 = hbusreq1 & v22f9911 | !hbusreq1 & !v22ebbea;
assign v22fc9cf = hmaster2_p & v23056b1 | !hmaster2_p & v12cd3f4;
assign v191ae7d = hbusreq4 & v22efa5e | !hbusreq4 & v22fc23d;
assign v23fc9bf = hbusreq4 & v23fbb99 | !hbusreq4 & v23fbfcb;
assign v230ae3f = hmaster2_p & v84561b | !hmaster2_p & !v12cc2ef;
assign v23fb102 = hbusreq3_p & v230c4ae | !hbusreq3_p & v22f903f;
assign v23fca0a = hbusreq5 & v22f65d5 | !hbusreq5 & v22f5583;
assign b9c969 = hbusreq5_p & v22f17bb | !hbusreq5_p & v23fce79;
assign v22faa1f = hburst0_p & v84561b | !hburst0_p & v23fb77e;
assign v22fc10a = hgrant1_p & v23f5043 | !hgrant1_p & b2aff2;
assign v23fbe63 = hmaster0_p & v23fcec5 | !hmaster0_p & v23115e2;
assign v2304faf = hmaster2_p & v23fc2d2 | !hmaster2_p & !v84561b;
assign v2309b3a = stateG10_5_p & v22f3e40 | !stateG10_5_p & v845636;
assign v2304189 = hgrant3_p & v22fe58b | !hgrant3_p & v22eb99d;
assign v23fcf21 = hbusreq3 & v23f8466 | !hbusreq3 & v84561b;
assign v23f439a = hbusreq3_p & v22f62ae | !hbusreq3_p & v22f53c0;
assign v23f97de = hbusreq1 & v23fb1a4 | !hbusreq1 & !v84561b;
assign v22f91a6 = hmaster0_p & v22ef4f0 | !hmaster0_p & v23f0cce;
assign v230f795 = hmaster2_p & v2313476 | !hmaster2_p & v845620;
assign v230fe41 = jx0_p & v230b3d2 | !jx0_p & v22fbbd2;
assign v22eba12 = hgrant0_p & v84564d | !hgrant0_p & a476c2;
assign v23f4e25 = hbusreq1 & v23f2d8c | !hbusreq1 & v84561b;
assign v23f340b = hbusreq0 & v23f1f6f | !hbusreq0 & v84561b;
assign v23ef95a = hgrant3_p & v84561b | !hgrant3_p & v23f6849;
assign v2304d26 = jx1_p & v22f1e8e | !jx1_p & v2313429;
assign v23fa0a3 = hgrant3_p & v22f2ca2 | !hgrant3_p & v2301bcb;
assign v22f7758 = hgrant3_p & v23fc43e | !hgrant3_p & v2303270;
assign v23fc8a1 = hmaster1_p & v22fff51 | !hmaster1_p & v84561b;
assign v22fa105 = hgrant1_p & v23fbb80 | !hgrant1_p & v22f6246;
assign v22f85f2 = jx0_p & v23fb1e0 | !jx0_p & v22fd693;
assign v1aaddf4 = hmaster2_p & v23fbfb9 | !hmaster2_p & v22fa870;
assign v22eb3c2 = hbusreq5 & v22f8cb7 | !hbusreq5 & v84561b;
assign v22ec992 = hbusreq0 & v22eda43 | !hbusreq0 & v84561b;
assign v2301073 = hgrant3_p & v23fbf5d | !hgrant3_p & v22ecc3b;
assign v2391e26 = jx1_p & v85e5cf | !jx1_p & v23fb9c9;
assign v2304f67 = hmaster2_p & v22fc9bf | !hmaster2_p & !v22f7879;
assign v23fc390 = hmaster0_p & v22fc8e5 | !hmaster0_p & v23f99ae;
assign v23f40d1 = hbusreq1 & v22f8834 | !hbusreq1 & v84561b;
assign v23f7e8f = hbusreq6 & v23fc369 | !hbusreq6 & v84561b;
assign v2308c76 = hmaster2_p & v22ec71a | !hmaster2_p & v23f7d57;
assign v22fb9ad = hmaster0_p & v2308967 | !hmaster0_p & v23fb1d6;
assign v23fce66 = stateG10_5_p & v2310251 | !stateG10_5_p & v23f7ea0;
assign v22fd83a = hbusreq6_p & v2302245 | !hbusreq6_p & v22f1383;
assign v23067c3 = hmaster0_p & v23066bf | !hmaster0_p & !v23fc9be;
assign v8c875e = hlock3_p & v230d235 | !hlock3_p & !v23fac6d;
assign v22f0b62 = hgrant1_p & v22f8271 | !hgrant1_p & v22f22ec;
assign v23fb1e0 = jx1_p & v22f9554 | !jx1_p & v983a4e;
assign v2307e2c = hbusreq5 & v22ef945 | !hbusreq5 & !v84561b;
assign f40a94 = hgrant5_p & v22f47fe | !hgrant5_p & v23fb993;
assign v22fccbd = hbusreq6 & v23fbb5a | !hbusreq6 & v845622;
assign v22f8f1e = hbusreq3_p & v23fc19b | !hbusreq3_p & v23f2d31;
assign v230391b = hbusreq3 & v230bf9f | !hbusreq3 & v84561b;
assign v15075f0 = jx0_p & v22ed654 | !jx0_p & v230564d;
assign v22fb068 = hbusreq4 & v230e0d6 | !hbusreq4 & v22f9bc8;
assign v2311af8 = hmaster2_p & v191a86f | !hmaster2_p & v22ecc15;
assign v12cd69f = hbusreq2_p & v23fce71 | !hbusreq2_p & b9d02f;
assign v22fa628 = hmaster2_p & v8912cf | !hmaster2_p & v23022b1;
assign v22f52d4 = hbusreq3_p & v23fb138 | !hbusreq3_p & v22fe2ae;
assign v106ae4a = hmastlock_p & v23fba29 | !hmastlock_p & v84561b;
assign v23fb9fe = hbusreq1_p & v22f69eb | !hbusreq1_p & !v84561b;
assign v230a891 = hlock3_p & v22f4a20 | !hlock3_p & v2306de4;
assign v23f9593 = hbusreq1 & v2301e25 | !hbusreq1 & v84561b;
assign v2304568 = hmaster1_p & v84561b | !hmaster1_p & v2309520;
assign v23fcfaa = hmaster2_p & v23060d4 | !hmaster2_p & v22f31b2;
assign v22ede9f = hbusreq3_p & v23f63dc | !hbusreq3_p & v22fd8c5;
assign v2307c3d = hbusreq6 & v2304dc4 | !hbusreq6 & v23fb0ee;
assign v231101b = hbusreq3_p & v23fbac0 | !hbusreq3_p & v23f5948;
assign v23fc5b7 = hmaster1_p & v84561b | !hmaster1_p & v23f88a1;
assign v2307aad = hmaster2_p & v84561b | !hmaster2_p & v23f8a9d;
assign v22ebfcb = hbusreq4 & v22f3cc0 | !hbusreq4 & v23fba11;
assign v22fb877 = hbusreq2_p & v22f1a26 | !hbusreq2_p & !v23fb1a4;
assign v23110f1 = hgrant3_p & v84561b | !hgrant3_p & v230c79d;
assign v23090a6 = hmaster0_p & v87d737 | !hmaster0_p & da3103;
assign v2303b0a = hbusreq4 & v13aff51 | !hbusreq4 & !v22f5198;
assign v23fcaf6 = hgrant3_p & v84561b | !hgrant3_p & !v23fbf31;
assign v230ff13 = busreq_p & v23f707f | !busreq_p & !v23085df;
assign v2310fcd = hgrant1_p & v84561b | !hgrant1_p & v23fcdce;
assign v230d513 = hbusreq6 & v23fbe89 | !hbusreq6 & !v23fc2b4;
assign v23f62ee = hmaster0_p & v22f8e29 | !hmaster0_p & v22f5568;
assign v150736d = hgrant5_p & v230875c | !hgrant5_p & v23f5d6f;
assign v23fbdb1 = hlock3_p & v23fbd64 | !hlock3_p & v22f5218;
assign v23fc0b7 = hmaster1_p & v84561b | !hmaster1_p & v22f6963;
assign v2308e3c = hgrant2_p & v23fc882 | !hgrant2_p & !v12cd3f4;
assign v22f968e = hmaster0_p & v22f1ae9 | !hmaster0_p & v22f2fe1;
assign v22ecce6 = hmaster2_p & v22f9a51 | !hmaster2_p & v84561b;
assign da30f9 = hbusreq5_p & v230e100 | !hbusreq5_p & v23fbb8a;
assign v23f2199 = hmaster0_p & v23fba92 | !hmaster0_p & v2391568;
assign v23fb709 = hbusreq1 & v230e4ae | !hbusreq1 & v84561b;
assign v2305a09 = hbusreq3_p & v2308aec | !hbusreq3_p & v22f3643;
assign v23063de = jx1_p & v22f4cb3 | !jx1_p & v23f82dd;
assign v23037d3 = hlock6_p & v230ef38 | !hlock6_p & v2312d71;
assign v23f7822 = hbusreq4_p & v2300420 | !hbusreq4_p & v23fc76e;
assign v22fc7b7 = hmaster2_p & v22fe5b1 | !hmaster2_p & v22f0860;
assign v23fbbc5 = hlock4_p & v8920c5 | !hlock4_p & v22eb970;
assign v23fcb10 = hbusreq1_p & v84561b | !hbusreq1_p & adb81d;
assign v22fb2b4 = hbusreq1_p & v2303329 | !hbusreq1_p & bab0c9;
assign v230e568 = jx1_p & v2300e92 | !jx1_p & v23f60dc;
assign v2310f77 = hgrant3_p & v84562e | !hgrant3_p & v22f4301;
assign v22ffff6 = hbusreq1_p & v2306b2e | !hbusreq1_p & !v23f5a2e;
assign v23f37ba = hbusreq5 & v22f60c6 | !hbusreq5 & !v2304ec7;
assign v23f8c1f = hbusreq6 & v23fbe89 | !hbusreq6 & !v2303cfd;
assign v23fbe7e = hbusreq0 & v13afe8f | !hbusreq0 & v84561b;
assign v23f9904 = hburst1 & v22f3294 | !hburst1 & v230204f;
assign v23fb0ee = hmaster2_p & v23f2ecd | !hmaster2_p & v84561b;
assign v22f8639 = jx0_p & v23f7c5a | !jx0_p & v23123a3;
assign v22fbfaf = hgrant0_p & v230fb99 | !hgrant0_p & v22f76f0;
assign v23130dd = hmaster2_p & a1fba6 | !hmaster2_p & v230ceb6;
assign v23fb4e5 = hgrant3_p & v22eb9b4 | !hgrant3_p & v230160e;
assign a6c3d1 = hbusreq4_p & v23f6827 | !hbusreq4_p & v23fb323;
assign v22edb43 = hmaster2_p & v22ff414 | !hmaster2_p & v22ee772;
assign v2305bb2 = hlock1_p & v84561b | !hlock1_p & !v2391a57;
assign ae3590 = hmaster0_p & v23fba1a | !hmaster0_p & v191b17f;
assign v23f62f2 = hbusreq4_p & b1d009 | !hbusreq4_p & v22eaeaf;
assign v23f6478 = hmaster2_p & v22f0132 | !hmaster2_p & v23f9f77;
assign v23f6ef7 = jx1_p & v23f651e | !jx1_p & v230d32a;
assign v22f79fb = locked_p & v23f2862 | !locked_p & !v23fba6b;
assign v2304477 = hbusreq3_p & b5b985 | !hbusreq3_p & v84561b;
assign v22fe542 = hbusreq1_p & v2309c55 | !hbusreq1_p & v23fba3e;
assign v23fb574 = hbusreq1 & v1507134 | !hbusreq1 & !aa6574;
assign b9d0a0 = hbusreq3 & v2301e43 | !hbusreq3 & v84564d;
assign v22faee9 = stateG10_5_p & v23fc8f9 | !stateG10_5_p & v2308b7c;
assign v22f2f16 = hgrant3_p & v23fc975 | !hgrant3_p & v230a1c7;
assign v845633 = hlock4_p & v84561b | !hlock4_p & !v84561b;
assign v230c15a = hmaster2_p & v2304ec7 | !hmaster2_p & !v84564d;
assign v23f7ed6 = hbusreq6_p & v23f0489 | !hbusreq6_p & v84561b;
assign v22ffa4c = hgrant3_p & v84561b | !hgrant3_p & v22fb30f;
assign v2303943 = hbusreq5_p & v22f1a26 | !hbusreq5_p & v23f22f9;
assign v23fcabe = hlock4_p & v23fc92d | !hlock4_p & v22f0ad8;
assign v23f4872 = hbusreq0_p & v22f264f | !hbusreq0_p & v23ef9c4;
assign v106a7a3 = hbusreq5_p & v23f987b | !hbusreq5_p & v84561b;
assign v22f7659 = hbusreq3_p & v22f8ad5 | !hbusreq3_p & v23faaa0;
assign v23fc750 = hmaster2_p & v2310e81 | !hmaster2_p & v23fc362;
assign v23f179d = hbusreq3_p & v22ef2aa | !hbusreq3_p & v2311bc4;
assign v23022d0 = hgrant3_p & v84561b | !hgrant3_p & v23f7853;
assign v23fb4be = hgrant1_p & v23fbe41 | !hgrant1_p & v22eb6dd;
assign v22fcf7a = hbusreq1_p & v22f1b4e | !hbusreq1_p & v22ed7a8;
assign v22ef65b = hbusreq3 & v23f832b | !hbusreq3 & v84561b;
assign v23109c3 = hgrant1_p & v845647 | !hgrant1_p & !e1dcf1;
assign v22f7ad4 = hbusreq6 & v23fbe4f | !hbusreq6 & v84561b;
assign ba569c = hbusreq5 & v2306bb2 | !hbusreq5 & v22fb71d;
assign v106a7d6 = stateA1_p & v22f79de | !stateA1_p & v23f9904;
assign v22f53df = stateG10_5_p & v230b756 | !stateG10_5_p & v22f0945;
assign v23fb6b6 = hmaster0_p & v23f20d0 | !hmaster0_p & v2310197;
assign v23f682a = hbusreq3 & v22fe0ef | !hbusreq3 & v84561b;
assign v23fceec = hbusreq5 & v22ee9be | !hbusreq5 & v23f3d14;
assign v23fba0f = hmaster2_p & v84561b | !hmaster2_p & v22f0bb4;
assign v23fba4a = hlock6_p & bc87ee | !hlock6_p & !v23f5474;
assign v12cc317 = hlock5_p & v22eec14 | !hlock5_p & !v84561b;
assign v22f9601 = hmaster1_p & v23f7cbe | !hmaster1_p & v22fa6ae;
assign v22ff94b = hbusreq3_p & v23110a4 | !hbusreq3_p & v23f47b3;
assign v23fc21c = hbusreq3 & v230e85f | !hbusreq3 & v22f2ffe;
assign v23fc8f9 = hbusreq5 & v22f3959 | !hbusreq5 & v230d630;
assign v22ecaeb = hgrant3_p & v84561b | !hgrant3_p & v1aadb61;
assign v22fba66 = hgrant5_p & v22f2f19 | !hgrant5_p & v2300c5a;
assign v23f8d76 = hgrant1_p & f405d5 | !hgrant1_p & v22ed267;
assign v22ef816 = hbusreq5_p & v23f60ef | !hbusreq5_p & b9c9ef;
assign v23fbd3a = jx1_p & v22f7b24 | !jx1_p & v22eb95e;
assign v22f46b1 = hbusreq6 & fc88ba | !hbusreq6 & v230a83f;
assign v230104a = hbusreq1_p & v2391a57 | !hbusreq1_p & !v84561b;
assign v22ee323 = hmaster2_p & v8a7512 | !hmaster2_p & v84561b;
assign v23fcac2 = hlock0_p & v23fb5e3 | !hlock0_p & !v845622;
assign v22eb6fc = hgrant5_p & v2304299 | !hgrant5_p & !v2391a62;
assign v23f35c4 = hbusreq2 & v22f79fd | !hbusreq2 & v84561b;
assign v22eba97 = hmaster0_p & v22eb6ab | !hmaster0_p & v23fca63;
assign v23f924a = hmaster2_p & v1507529 | !hmaster2_p & v2310682;
assign v230446f = hbusreq2 & v191a86f | !hbusreq2 & v84561b;
assign v23fc178 = stateG10_5_p & v84561b | !stateG10_5_p & !v84564d;
assign v23f88d9 = hmaster0_p & v23fce64 | !hmaster0_p & v1507446;
assign v2304048 = hgrant3_p & v84562d | !hgrant3_p & v22fa646;
assign v2393b5a = hbusreq5_p & v2300b96 | !hbusreq5_p & v23064ae;
assign v23fbe2d = hmaster2_p & v22ee73b | !hmaster2_p & v23f931e;
assign bc2a58 = hbusreq1 & v22fb77d | !hbusreq1 & !v23108b7;
assign v23fc91f = hbusreq2 & v22ed85a | !hbusreq2 & v84561b;
assign v23f9283 = hmaster0_p & v2302514 | !hmaster0_p & v2307b93;
assign v22ed8a3 = hbusreq3 & v84564d | !hbusreq3 & v230a8b2;
assign v230fa04 = hbusreq6 & v23f14ef | !hbusreq6 & v22f9280;
assign v23f7961 = hlock0_p & v23f2cbb | !hlock0_p & !v84561b;
assign v230b9b4 = hmaster2_p & v84561b | !hmaster2_p & v23126fc;
assign v23fc765 = hgrant1_p & v22f2ed7 | !hgrant1_p & v23fc26f;
assign v2309465 = hbusreq3_p & v23fcf65 | !hbusreq3_p & v22fa055;
assign v230979f = hgrant0_p & v84561b | !hgrant0_p & !v23f4462;
assign v23fb12a = hbusreq0 & v230882d | !hbusreq0 & v23f8364;
assign v22fe6c8 = hbusreq5_p & v2392d52 | !hbusreq5_p & v239383b;
assign v23f4e1c = hbusreq3_p & v23f1e4f | !hbusreq3_p & v84561b;
assign v2304937 = hlock0_p & v94dcdf | !hlock0_p & !v23efdd4;
assign v23fc01c = hgrant2_p & v2306fa2 | !hgrant2_p & !v2301d10;
assign v23fcb0a = hbusreq1 & v23fbfd0 | !hbusreq1 & b9d02f;
assign v23fbe06 = hmaster1_p & v2301bb5 | !hmaster1_p & v23120b1;
assign v230b789 = hmaster0_p & v2301b52 | !hmaster0_p & v23fbb42;
assign v22fa309 = hmaster1_p & v23f215c | !hmaster1_p & v94f831;
assign v22efa0f = hgrant3_p & v23fab26 | !hgrant3_p & !v22ef2b4;
assign v22f1e91 = hbusreq1_p & v23fb1ab | !hbusreq1_p & v23fb5b4;
assign v23fb231 = hbusreq3_p & v22fec56 | !hbusreq3_p & v230f9f1;
assign v22ee057 = hmaster0_p & v2312a52 | !hmaster0_p & v22f8d58;
assign v23fbafc = hmaster2_p & v23fcf69 | !hmaster2_p & v23f9b8d;
assign v23fbe79 = hmaster2_p & v2310d04 | !hmaster2_p & v2309cdc;
assign v23f476a = hmaster2_p & v22eeb03 | !hmaster2_p & v2306d29;
assign v2301484 = hmaster0_p & v22f6d61 | !hmaster0_p & v230f0de;
assign v23fca7d = hgrant2_p & v845620 | !hgrant2_p & !v23f5043;
assign v2309066 = hbusreq0 & v230913d | !hbusreq0 & !v22f8ac3;
assign v231248c = hbusreq4_p & v23121ff | !hbusreq4_p & v230e7d6;
assign v2311246 = hmaster0_p & v23fc002 | !hmaster0_p & v23fc07e;
assign v23fcc0c = hbusreq3_p & v23fbf36 | !hbusreq3_p & v2309c93;
assign v12cd4f6 = hmaster2_p & v22f0945 | !hmaster2_p & v22f8543;
assign v230ba0a = hgrant0_p & v2313463 | !hgrant0_p & !v23f908f;
assign v23125a8 = hmaster0_p & v2306fba | !hmaster0_p & v22f8be5;
assign v23f3bde = hlock4_p & v22fa5f1 | !hlock4_p & !v23f38f8;
assign v2308fc5 = hbusreq5_p & v22faefb | !hbusreq5_p & !v22f1d46;
assign v2303c9e = hbusreq5 & v84561b | !hbusreq5 & !v23fc732;
assign v23fc851 = hmaster2_p & v191aa68 | !hmaster2_p & v22f7d4e;
assign v23fbcba = hgrant3_p & v84561b | !hgrant3_p & v8d83bb;
assign v12cd995 = hburst1_p & v230371b | !hburst1_p & v84561b;
assign b9ca52 = decide_p & v23fb189 | !decide_p & v23f1a76;
assign v22f3b08 = hgrant3_p & v2308967 | !hgrant3_p & f40c96;
assign v2305fbf = hbusreq3_p & v23fcf5d | !hbusreq3_p & v84561b;
assign v22fbda1 = hgrant2_p & v84562a | !hgrant2_p & v2310fde;
assign v2302983 = hmaster0_p & f40ab9 | !hmaster0_p & v23fb97c;
assign v23fcdbd = jx2_p & v22eccde | !jx2_p & v22edd4c;
assign v230ad18 = hmaster0_p & v2300d5f | !hmaster0_p & v230fb96;
assign v22fe59c = hbusreq1 & v23fc4a5 | !hbusreq1 & v22f0add;
assign v22f8bd0 = hbusreq1_p & v22f30be | !hbusreq1_p & v84561b;
assign v23f90bc = hmaster2_p & v845647 | !hmaster2_p & !v22fafe4;
assign v22f3519 = hmaster0_p & v2312196 | !hmaster0_p & v23fc76a;
assign v22ebc57 = hgrant3_p & v84561b | !hgrant3_p & v22fb5da;
assign v23fc948 = hbusreq4 & v1507157 | !hbusreq4 & v22ee657;
assign v22f07d3 = hbusreq3_p & v22ec882 | !hbusreq3_p & v22f57e9;
assign v230cfe6 = hbusreq1 & v22fcdf6 | !hbusreq1 & v84561b;
assign v13afbf5 = hmastlock_p & v22f2759 | !hmastlock_p & !v84561b;
assign v22fa821 = hbusreq2 & v845620 | !hbusreq2 & !v84561b;
assign v12cc6e0 = hmaster2_p & v84561b | !hmaster2_p & v23fc198;
assign v23fcfba = hmaster0_p & v22ec2e6 | !hmaster0_p & v22fb068;
assign v230f347 = hgrant1_p & v23fb6ff | !hgrant1_p & v2307788;
assign v23043b7 = hbusreq4 & v230a67e | !hbusreq4 & v23f2b69;
assign v1aae98c = hbusreq2_p & v23fb104 | !hbusreq2_p & v84561b;
assign v23f8979 = hbusreq2_p & v23fc303 | !hbusreq2_p & v84561b;
assign v230d02b = hmaster0_p & v230ea9f | !hmaster0_p & v106af01;
assign v23034f8 = hlock3_p & v23fce7d | !hlock3_p & !v84561b;
assign v22f409f = hgrant5_p & v23fbe4d | !hgrant5_p & !v230b20b;
assign v23fbe8e = hmaster2_p & v23f9e4f | !hmaster2_p & v23f15ac;
assign v23fbad3 = hbusreq3_p & v2391e8f | !hbusreq3_p & v230f4e5;
assign v23fbfb5 = hmaster2_p & v84561b | !hmaster2_p & !v22fec81;
assign v22f8613 = hbusreq4 & v22ee4d5 | !hbusreq4 & v84561b;
assign v230471d = hgrant1_p & v84561b | !hgrant1_p & v23124e2;
assign v22f1faf = hlock1_p & v23fc346 | !hlock1_p & !v84561b;
assign v23f3b8f = hbusreq6 & v23fc234 | !hbusreq6 & v84561b;
assign v23f328e = hbusreq1_p & v22f1ae5 | !hbusreq1_p & v23f53e4;
assign v2309d23 = hmaster2_p & v22fd25c | !hmaster2_p & !v23fcc36;
assign v22f7d93 = jx1_p & v22ec74f | !jx1_p & v22ff727;
assign v23fb553 = hbusreq3 & v2311d38 | !hbusreq3 & v23fba11;
assign v230361d = hmaster2_p & b10190 | !hmaster2_p & v2393346;
assign v23f6cdb = hmaster2_p & v191aa68 | !hmaster2_p & v22fa5a5;
assign b3cfb7 = hbusreq6 & v23f67e2 | !hbusreq6 & v23fa2ec;
assign v22ef575 = hgrant3_p & v23fbf0f | !hgrant3_p & v2313041;
assign v23fc683 = start_p & v84561b | !start_p & v230a434;
assign v22eec2a = hmaster2_p & v23fbfb9 | !hmaster2_p & v22eb1f5;
assign v230064b = hbusreq3_p & v23fb77d | !hbusreq3_p & c16218;
assign v2307e4c = hmaster2_p & v22f995e | !hmaster2_p & v23f660f;
assign v22fa5fd = hbusreq1_p & v23f3d14 | !hbusreq1_p & v2310a55;
assign v23fbbf3 = stateA1_p & v84561b | !stateA1_p & !v22f4e3c;
assign v2307d4e = hgrant1_p & v23fc102 | !hgrant1_p & v2301fe9;
assign v2302d68 = jx0_p & v22f07fc | !jx0_p & !v23f623e;
assign v231363b = hbusreq6 & v22ec191 | !hbusreq6 & v2306873;
assign v22ef0fe = hbusreq2 & v2313118 | !hbusreq2 & v84561b;
assign v23fcd38 = hgrant5_p & v231164b | !hgrant5_p & v23f4254;
assign v23f80cc = hbusreq3 & v23f52c1 | !hbusreq3 & v22fae48;
assign v23f1221 = jx3_p & v23f2af5 | !jx3_p & v22fb631;
assign v230b09e = hlock1_p & v84561b | !hlock1_p & v2312351;
assign v22f1491 = hmaster2_p & v2307758 | !hmaster2_p & v22fb74c;
assign v23fb21a = hmaster0_p & v22fa27c | !hmaster0_p & v2309ce6;
assign v23fc0da = hlock0_p & v2308fe7 | !hlock0_p & !v22fc997;
assign v23f97bb = hmaster2_p & v2305811 | !hmaster2_p & v1507071;
assign v23077dc = hmaster2_p & v22fabd2 | !hmaster2_p & v2310108;
assign v230b8fe = hmaster2_p & v191a86f | !hmaster2_p & v2309871;
assign v23fd035 = hgrant3_p & v23074c0 | !hgrant3_p & v2303e03;
assign v23f8c7b = hgrant5_p & v23038a2 | !hgrant5_p & v23fb993;
assign v231086d = hbusreq5 & v23f5043 | !hbusreq5 & v84561b;
assign v2300985 = hbusreq4 & v2302783 | !hbusreq4 & !v23fbeeb;
assign v23fb73e = hbusreq6_p & v23fcf56 | !hbusreq6_p & v23f8324;
assign v23f789c = hmaster2_p & v22f2db0 | !hmaster2_p & v22fda32;
assign v23063fa = hgrant6_p & v2302ba4 | !hgrant6_p & v2303220;
assign v22fdd29 = hmaster0_p & v23fcab7 | !hmaster0_p & v23077ec;
assign v23fb043 = hbusreq4 & v230a65d | !hbusreq4 & v22ef062;
assign v23fbe1b = hbusreq1_p & v23fb4d3 | !hbusreq1_p & v845620;
assign v23093e2 = hbusreq4 & v23083c1 | !hbusreq4 & v23130b0;
assign v1aad9cb = hlock6_p & v23fcb96 | !hlock6_p & v23024e8;
assign v22fb0cb = hmaster2_p & v22eeb03 | !hmaster2_p & v2310e40;
assign v230a71c = hbusreq3_p & v230e262 | !hbusreq3_p & v230a226;
assign v22f73a9 = hbusreq4_p & v23fcb60 | !hbusreq4_p & v23fc7cb;
assign v23fc2ae = hbusreq3_p & v22f42a5 | !hbusreq3_p & v23f56bc;
assign v23fa9dd = stateG10_5_p & v22fddc8 | !stateG10_5_p & !v230e72d;
assign v22f7fdd = hbusreq3_p & v22efe81 | !hbusreq3_p & v22f91ef;
assign v22f3643 = hready & v84564d | !hready & !v84561b;
assign v97b973 = hlock5_p & v23f420e | !hlock5_p & !v845636;
assign v22f7f52 = hmastlock_p & v22faeec | !hmastlock_p & v84561b;
assign v22fd2e2 = stateG10_5_p & v23fb82c | !stateG10_5_p & v22fcc0d;
assign v22fcf04 = hmaster0_p & v23fbad4 | !hmaster0_p & v23f82b3;
assign v230bdd4 = hbusreq4_p & v23fa2c3 | !hbusreq4_p & v231156b;
assign v230444c = hbusreq4_p & v23116b7 | !hbusreq4_p & v23fc04e;
assign v2303cfd = hmaster2_p & v22fc6d7 | !hmaster2_p & v84561b;
assign v23fcb38 = hmastlock_p & v23085df | !hmastlock_p & v84561b;
assign v23919bb = hbusreq1_p & v230cb59 | !hbusreq1_p & v23f7796;
assign v23fca37 = hbusreq5 & v22ee7a7 | !hbusreq5 & !v84561b;
assign v2311c16 = hlock3_p & v23020a2 | !hlock3_p & v2305b2e;
assign v22f6124 = hbusreq3_p & v22ed805 | !hbusreq3_p & a1fda8;
assign v22ff0d2 = stateG10_5_p & v997ca9 | !stateG10_5_p & !v845647;
assign v2302b2c = hbusreq3_p & v22f695c | !hbusreq3_p & v23fbc97;
assign v230d8b2 = hmaster2_p & v22f4e0b | !hmaster2_p & v84564d;
assign v23fc19c = hgrant0_p & v845623 | !hgrant0_p & v23fc686;
assign v22ff83d = hmaster2_p & v23fb155 | !hmaster2_p & v22f7b29;
assign v230e13a = hbusreq1_p & v22f17bb | !hbusreq1_p & b9c969;
assign v23fcbe8 = hmaster2_p & v23f86f0 | !hmaster2_p & v230f848;
assign v23fc1bb = hbusreq5 & v22fef02 | !hbusreq5 & v84561b;
assign v22f803b = hmaster1_p & v22f4af5 | !hmaster1_p & v2310cbb;
assign v23f9d8e = hmaster2_p & v22eec6e | !hmaster2_p & v22f1796;
assign v22f4d65 = hbusreq5_p & v84561b | !hbusreq5_p & !v230a580;
assign v22fe605 = jx0_p & v22f6bba | !jx0_p & v23104a1;
assign v23fc4fb = hbusreq0_p & v23fc1c1 | !hbusreq0_p & v23fc564;
assign v22fa945 = hbusreq5_p & v84561b | !hbusreq5_p & v23fcec3;
assign v13afef6 = hbusreq4_p & v22f9dab | !hbusreq4_p & v22f752e;
assign v23f8383 = hbusreq5 & v22f15fe | !hbusreq5 & v23f60ef;
assign v23fba73 = hbusreq3 & v22ee9be | !hbusreq3 & v84561b;
assign v230abb0 = hmaster2_p & v2310e40 | !hmaster2_p & v230f63f;
assign v2310d2f = hlock3_p & v22feb47 | !hlock3_p & !v84561b;
assign v23fb47e = hbusreq1_p & v22f1a26 | !hbusreq1_p & !v23fb1a4;
assign v22f438c = hmaster2_p & v2313463 | !hmaster2_p & !v23f5c95;
assign v23f820a = hbusreq5 & v2391a57 | !hbusreq5 & !v84561b;
assign v23fcb89 = start_p & v84561b | !start_p & !v22fb386;
assign v22eedbb = hmaster0_p & v22f878c | !hmaster0_p & v23f35a8;
assign v23fc3cd = hmaster0_p & v2308967 | !hmaster0_p & v2303ae8;
assign v230fa13 = hgrant0_p & v84561b | !hgrant0_p & v23fc949;
assign v22ffb9d = hlock0_p & v23fbb35 | !hlock0_p & v84561b;
assign v2310303 = hlock1_p & v22ffbb3 | !hlock1_p & !v230f848;
assign v22f7ec4 = hbusreq5_p & v23fc3cb | !hbusreq5_p & v23fc2e8;
assign v23fbdbe = hmaster2_p & v84564d | !hmaster2_p & v23f5043;
assign v22ece0d = hbusreq5_p & v23fbc5a | !hbusreq5_p & v22f4d68;
assign v230f9c8 = hlock5_p & v230f2d1 | !hlock5_p & v22f0d22;
assign v230efee = hbusreq3_p & v2393d28 | !hbusreq3_p & !v845645;
assign v23fa931 = hburst0_p & v22f178d | !hburst0_p & !v23fc17d;
assign v22f6ae5 = hmaster2_p & v22eb377 | !hmaster2_p & v22ee956;
assign v230eb5a = hlock3_p & v22f4eab | !hlock3_p & v230cfc7;
assign v22f3aa1 = hgrant1_p & v22f6b45 | !hgrant1_p & v230580d;
assign v2307517 = hmaster2_p & v23fc716 | !hmaster2_p & v84561b;
assign v22ef542 = stateG10_5_p & v1e84012 | !stateG10_5_p & v22eed5b;
assign v23f9666 = hmaster2_p & v84561b | !hmaster2_p & v230b713;
assign v23f3c28 = hbusreq3_p & v23fc38f | !hbusreq3_p & v22efce2;
assign v23f763f = hlock0_p & b572e8 | !hlock0_p & v22f2481;
assign bd8af4 = hbusreq3_p & v23fcea8 | !hbusreq3_p & v22f4114;
assign v23117af = locked_p & v84561b | !locked_p & !v22f7f74;
assign v23fcea0 = hmaster0_p & v23fceb9 | !hmaster0_p & v22f4d77;
assign v2393485 = hgrant3_p & v845635 | !hgrant3_p & v22f4bea;
assign v23f5a6d = jx3_p & v22f4284 | !jx3_p & v22eb6e2;
assign v230bb69 = hgrant3_p & v2303226 | !hgrant3_p & v22f728a;
assign v23f4fa1 = hgrant0_p & v23fc0da | !hgrant0_p & !v22f7d41;
assign v230c2f4 = hbusreq1_p & v84561b | !hbusreq1_p & !v106a782;
assign v230f7ce = hmaster2_p & v191a86f | !hmaster2_p & v23f3a16;
assign v22ec41b = hbusreq5_p & v23fbc48 | !hbusreq5_p & v230b573;
assign v23f8328 = hbusreq6_p & v2308bfc | !hbusreq6_p & v23f20a8;
assign v23fbd50 = jx1_p & v23f592f | !jx1_p & v22ef78e;
assign v230e40a = hbusreq0_p & v84561b | !hbusreq0_p & v845629;
assign v2391f87 = hgrant5_p & v23fbe7a | !hgrant5_p & !v84561b;
assign v23fbd76 = hbusreq1 & v231228e | !hbusreq1 & !v84561b;
assign v23fbf61 = hgrant3_p & v8cded5 | !hgrant3_p & v23f4cfb;
assign v23f5019 = hbusreq3_p & v23f558b | !hbusreq3_p & v23fd02c;
assign v2307205 = hgrant5_p & v22fb68b | !hgrant5_p & v2392a0d;
assign v23f149d = hbusreq3 & v23fcb67 | !hbusreq3 & !v845636;
assign v23fc356 = hbusreq5_p & v22edbe0 | !hbusreq5_p & v84561b;
assign v2393327 = hbusreq5_p & v230d1a6 | !hbusreq5_p & !v23fbde8;
assign v230056c = hmaster0_p & a1fbc2 | !hmaster0_p & v230f08b;
assign v22f95ec = hmaster0_p & v2307d30 | !hmaster0_p & v12cd66d;
assign v2306c5e = hgrant5_p & v84561b | !hgrant5_p & v106a7bd;
assign v2305b67 = hready_p & v22fa63e | !hready_p & v2312282;
assign v22eb16b = hbusreq5_p & v22f69cc | !hbusreq5_p & v9f009f;
assign f4064b = hmaster0_p & v1aae2a5 | !hmaster0_p & v2309b75;
assign v23f3e44 = hlock6_p & v22edec8 | !hlock6_p & v22f839c;
assign v23f5a02 = hmaster2_p & v23fcba3 | !hmaster2_p & v23fc164;
assign v23f193c = hgrant6_p & v84561b | !hgrant6_p & !v22f1d7b;
assign v12cd51b = hmaster0_p & v23fce0b | !hmaster0_p & v22f4858;
assign v2305748 = hbusreq1 & v22fc19c | !hbusreq1 & !v23fc596;
assign v23fc7b5 = jx0_p & v84561b | !jx0_p & v23faa93;
assign v23fcf65 = hmaster2_p & v845647 | !hmaster2_p & !v2310da0;
assign v2305c2e = hbusreq0 & v23f1207 | !hbusreq0 & b6f86d;
assign v23f9226 = hgrant1_p & v84561b | !hgrant1_p & v17a34ea;
assign v23f680b = hbusreq1_p & v23fb6c6 | !hbusreq1_p & v230a25a;
assign v1b87672 = hbusreq4 & v22fdf30 | !hbusreq4 & !v84561b;
assign v2305b74 = hmastlock_p & v23fcaa1 | !hmastlock_p & !v84561b;
assign v22f9d17 = hlock0_p & v22eedcf | !hlock0_p & v84561b;
assign v23fcefc = hmaster0_p & v23f95c3 | !hmaster0_p & v23f329a;
assign a1fdd3 = hbusreq6_p & v23fb818 | !hbusreq6_p & v2311da7;
assign v23fc15d = jx0_p & v2310c1a | !jx0_p & v23fca35;
assign v2302b44 = hbusreq5 & v23fcc10 | !hbusreq5 & v22ff090;
assign v22f02bd = hmaster0_p & v84561b | !hmaster0_p & b9d0ca;
assign v22f7808 = hgrant1_p & v22fb1bc | !hgrant1_p & v22ec299;
assign v22f8ad4 = hgrant5_p & v22eca17 | !hgrant5_p & v23fcb5e;
assign v2308e2e = hlock5_p & v23f2324 | !hlock5_p & v845620;
assign v230b837 = hgrant3_p & v230d8af | !hgrant3_p & v230ebb1;
assign v84563f = hburst1_p & v84561b | !hburst1_p & !v84561b;
assign v230592c = jx0_p & v23fc6e0 | !jx0_p & v2312d2c;
assign v2301450 = hmaster0_p & v22ed309 | !hmaster0_p & v23075ba;
assign v2304d0c = hmaster1_p & v23115b1 | !hmaster1_p & !v230c94b;
assign v22eb6dd = hgrant5_p & v22f6e47 | !hgrant5_p & v23fcb53;
assign v23fcc25 = hmaster1_p & v22f313c | !hmaster1_p & v22fd169;
assign v23fc71b = hbusreq1_p & v23f97de | !hbusreq1_p & !v84561b;
assign v22fcc05 = hgrant3_p & v23fbf5d | !hgrant3_p & v23f9631;
assign v22f04d8 = hgrant1_p & v84561b | !hgrant1_p & v2301e50;
assign v23ef89d = hgrant5_p & v2391b32 | !hgrant5_p & !v22f4f1e;
assign v23f8263 = hready_p & v22f6f7e | !hready_p & v2313328;
assign v22f95c8 = hbusreq1_p & v23f93ee | !hbusreq1_p & !v84561b;
assign v22f9acf = hlock0_p & v22f8271 | !hlock0_p & !v23056b1;
assign v22f01c1 = hgrant1_p & v22ee956 | !hgrant1_p & v23f243b;
assign v230b4d4 = hmaster2_p & v22f36ff | !hmaster2_p & !v22fef02;
assign v23fcf89 = hgrant1_p & v191b18a | !hgrant1_p & v22ed741;
assign v22f83cf = hgrant1_p & v23f4491 | !hgrant1_p & v23f6155;
assign v230538a = hmaster1_p & v1506eb2 | !hmaster1_p & a1fbc2;
assign v23f425f = hmaster2_p & v23f8928 | !hmaster2_p & v22ee0db;
assign v2305141 = hmaster1_p & v230ad74 | !hmaster1_p & v23fc087;
assign v23fb4a9 = hmaster1_p & v23f6c16 | !hmaster1_p & v22ffc31;
assign v22efd70 = hbusreq6 & v23f91e7 | !hbusreq6 & v230bdd6;
assign v23f32db = hbusreq3_p & v23f9a46 | !hbusreq3_p & !v22ee03c;
assign v23f2d39 = hbusreq3_p & v12cda11 | !hbusreq3_p & v23fa215;
assign v23f4f1e = hgrant1_p & v84561b | !hgrant1_p & v23fc4b1;
assign v23086ec = hmaster0_p & v22eb2fd | !hmaster0_p & !v84561b;
assign v2309c79 = hlock6_p & v84561b | !hlock6_p & v230089c;
assign v22f15fd = hbusreq2_p & v23fbc55 | !hbusreq2_p & v23fc739;
assign v22f288e = hgrant0_p & v22ee956 | !hgrant0_p & v23fb57d;
assign v22f3385 = hmaster2_p & v845620 | !hmaster2_p & v2310108;
assign v23fc89e = hbusreq6 & v2307f2b | !hbusreq6 & !v845622;
assign v23fc4a8 = hmaster2_p & v23fba49 | !hmaster2_p & v230d4d9;
assign v23f4900 = hmaster0_p & v230ac1b | !hmaster0_p & !v2312268;
assign v23fb5e9 = hgrant3_p & v23f817b | !hgrant3_p & v22fc4a3;
assign jx1 = b9ca52;
assign v23fc3f6 = jx0_p & v22ffffa | !jx0_p & v23fcd6d;
assign v2308ba7 = hbusreq4 & b00aa6 | !hbusreq4 & v22f1962;
assign v23052b7 = hmaster0_p & v23f54a0 | !hmaster0_p & !v95aaca;
assign bd8ac4 = hmaster0_p & v23f38b7 | !hmaster0_p & v230200a;
assign v23fc99a = hmaster2_p & v22ed878 | !hmaster2_p & v845620;
assign v23fac09 = hgrant3_p & v22f6ae5 | !hgrant3_p & v2301b70;
assign v22f0b0d = hgrant3_p & v84562e | !hgrant3_p & v23fbbf8;
assign v23fc523 = hmaster1_p & v22f6e51 | !hmaster1_p & v84561b;
assign v22f7078 = hburst1 & v84561b | !hburst1 & v23f6969;
assign v23fcaae = hmaster1_p & v23fc740 | !hmaster1_p & v23041ea;
assign v23fb99b = hbusreq1 & v22fd699 | !hbusreq1 & v845620;
assign v22ff2bf = hbusreq3_p & v2306292 | !hbusreq3_p & v230a579;
assign fc8c68 = hgrant1_p & v23fbe41 | !hgrant1_p & v106ae74;
assign v230de93 = hgrant5_p & v84561b | !hgrant5_p & v22feecb;
assign v2307f27 = stateG10_5_p & v84561b | !stateG10_5_p & v22ede4d;
assign v23f52f3 = jx1_p & v23fcc5e | !jx1_p & v23fc776;
assign v23f7f8d = hgrant1_p & v84561b | !hgrant1_p & v22f06fb;
assign v22f9445 = hmaster2_p & v23112ad | !hmaster2_p & v2311be9;
assign v23fcc24 = hbusreq1_p & v230a5e6 | !hbusreq1_p & v23fc126;
assign v23fc0cd = jx1_p & v2301b06 | !jx1_p & v23fcf4b;
assign v22ebe5c = jx1_p & v23f79e9 | !jx1_p & v84561b;
assign v230b20b = hbusreq5_p & v22f679f | !hbusreq5_p & v22efeed;
assign v23fc453 = hbusreq1 & v22f60c6 | !hbusreq1 & !v2391a57;
assign v23f2d6c = hmaster1_p & v84561b | !hmaster1_p & v23f0b27;
assign b72216 = hgrant3_p & v22f971b | !hgrant3_p & v230e8a0;
assign v22f8cee = hbusreq4_p & v22f1125 | !hbusreq4_p & v84561b;
assign v22ef46e = hbusreq1_p & v230bb63 | !hbusreq1_p & !v84561b;
assign v23fad76 = hbusreq0_p & v22f3502 | !hbusreq0_p & v230ad5b;
assign v2301adf = hbusreq6 & v23f6646 | !hbusreq6 & v84561b;
assign v23fcd69 = hgrant3_p & v84561b | !hgrant3_p & v23fc4ca;
assign stateG10_3 = !v11853d9;
assign v22ed999 = hbusreq4 & v191b1ba | !hbusreq4 & v2312e80;
assign v22f4407 = hbusreq1_p & v23fca5d | !hbusreq1_p & v22ee50f;
assign v2346b90 = jx1_p & v22f9188 | !jx1_p & v22fca1d;
assign v230418f = jx1_p & v2392394 | !jx1_p & v23f7c5a;
assign v22fb9eb = hbusreq3_p & v22ebc9f | !hbusreq3_p & v22fb6f9;
assign v23fbbf0 = hbusreq3_p & v23fb4a0 | !hbusreq3_p & v2302d3c;
assign v22ff399 = hgrant0_p & v2302779 | !hgrant0_p & !v22f12cd;
assign v23fb8e7 = hgrant5_p & v2307ff1 | !hgrant5_p & !v84561b;
assign v23fbea0 = hbusreq6_p & v22f85c2 | !hbusreq6_p & v2392cce;
assign v23fd025 = hbusreq3_p & v23f682a | !hbusreq3_p & v84561b;
assign v2307949 = hbusreq6 & v22f3cc0 | !hbusreq6 & v23fc223;
assign v22fccf1 = hbusreq5_p & v191a86f | !hbusreq5_p & !v191a879;
assign v23fc32f = hlock4_p & v2307cdf | !hlock4_p & v23f60e8;
assign v23fb704 = hlock6_p & v23f28de | !hlock6_p & bd7c6a;
assign v230ae1e = hgrant5_p & v230156d | !hgrant5_p & v23fc99f;
assign v2310430 = hgrant5_p & v22edaad | !hgrant5_p & v84561b;
assign v22f6ba1 = busreq_p & v106a782 | !busreq_p & !v84561b;
assign v23f47ae = hmaster1_p & v2309573 | !hmaster1_p & v23f7ed6;
assign v23fbb41 = hbusreq1 & v23fa9c5 | !hbusreq1 & v84561b;
assign v230e07d = hlock5_p & v23fceb9 | !hlock5_p & v84562b;
assign v22ee92e = hbusreq0 & v22f925b | !hbusreq0 & v84564d;
assign v191aec6 = hmaster2_p & v23fb6e3 | !hmaster2_p & v8be441;
assign v2392a17 = hbusreq5 & v2312f7e | !hbusreq5 & !v231009b;
assign v2302d3c = hbusreq3 & v22fe34f | !hbusreq3 & v22f803d;
assign v22ee09d = hmaster2_p & v84561b | !hmaster2_p & !v2305fe0;
assign v23fc5d4 = hlock3_p & v22ed07d | !hlock3_p & v2304faf;
assign v22f3101 = hbusreq5_p & v2308a0c | !hbusreq5_p & v845620;
assign v12cd931 = stateG10_5_p & v22eb5cc | !stateG10_5_p & v22fee46;
assign v2307b93 = hgrant3_p & v22f6ae5 | !hgrant3_p & v22eea08;
assign v23fbd6c = jx1_p & v2307ffd | !jx1_p & v230e1e0;
assign v230439f = hbusreq5_p & v845620 | !hbusreq5_p & v23919ec;
assign v23fcb43 = hbusreq6 & v23fb1c5 | !hbusreq6 & !v23fb593;
assign v23f4f34 = hlock1_p & v23f84cc | !hlock1_p & v22f3000;
assign v23f0234 = hbusreq6 & v13aff51 | !hbusreq6 & v84562f;
assign v23fc497 = hmaster2_p & v22f79fd | !hmaster2_p & v23f7123;
assign v230bdd0 = hbusreq1_p & v2312057 | !hbusreq1_p & v84561b;
assign v22f854f = hmaster2_p & v23fba6b | !hmaster2_p & v23fbfb9;
assign v12cdba9 = hmaster2_p & v2308d79 | !hmaster2_p & v23022b1;
assign v23fc2ca = hbusreq5_p & v23fc338 | !hbusreq5_p & v23f1f3e;
assign v23f3c00 = hlock3_p & v23faede | !hlock3_p & v23fcec8;
assign v191b04d = hbusreq5_p & v23fbe4c | !hbusreq5_p & v23f5fcd;
assign v23071be = hmaster1_p & v22fcc62 | !hmaster1_p & v22f58e8;
assign v2311b78 = hmaster2_p & v23f9b8d | !hmaster2_p & v84561b;
assign v230199e = hbusreq3_p & v22ec0de | !hbusreq3_p & v230a226;
assign v230c876 = hlock0_p & v2312067 | !hlock0_p & !v84561b;
assign v230b5c7 = hbusreq6_p & v23fb144 | !hbusreq6_p & v22f04b5;
assign v230b756 = hbusreq5 & v23920d8 | !hbusreq5 & v84561b;
assign v22ee918 = hbusreq3 & v23efbfd | !hbusreq3 & v84561b;
assign v23fc2fd = hbusreq0 & v23fc55f | !hbusreq0 & v84561b;
assign v2311c26 = hbusreq3_p & v22fbf28 | !hbusreq3_p & v84561b;
assign v23fbfaa = hmaster2_p & v23f55ea | !hmaster2_p & !v23fbca3;
assign v23fb947 = hbusreq4_p & v230089c | !hbusreq4_p & v22f9ab6;
assign v997ca9 = hgrant0_p & v17a34ff | !hgrant0_p & v230e71f;
assign v22eaaa7 = hmaster0_p & v22f9d92 | !hmaster0_p & v2302c67;
assign v23fcdb1 = hmaster1_p & v2302e98 | !hmaster1_p & v22fcd49;
assign v23f805c = hmaster1_p & v23fcca7 | !hmaster1_p & v23f741d;
assign v23fc572 = hbusreq1_p & v22fbb07 | !hbusreq1_p & v1506a9c;
assign v2302e87 = stateG10_5_p & v23f36a5 | !stateG10_5_p & !v84561b;
assign v230c771 = hready_p & v23fb9d4 | !hready_p & v17cf1d8;
assign v84562f = hlock3_p & v84561b | !hlock3_p & !v84561b;
assign v2302c42 = jx0_p & v22ec2d6 | !jx0_p & v230e991;
assign v23f85a9 = hbusreq4 & v230429d | !hbusreq4 & v23f90b2;
assign v23916d5 = hlock3_p & v22eb57a | !hlock3_p & !v84561b;
assign v23fcf35 = hgrant3_p & v84562e | !hgrant3_p & v991952;
assign v2305cf5 = hmaster2_p & v23fc38f | !hmaster2_p & v22ef5c2;
assign v22ec2e9 = hmaster1_p & v22f3b2e | !hmaster1_p & !v23f49cd;
assign v22eccde = hgrant4_p & c242c8 | !hgrant4_p & v23fcca2;
assign v23fc301 = hgrant3_p & v23050a2 | !hgrant3_p & v22fdc37;
assign v231242a = hgrant3_p & v84561b | !hgrant3_p & !v22fbe6a;
assign v9d1fa2 = hbusreq6 & v22f4fb2 | !hbusreq6 & v22ee657;
assign v230a4ef = hbusreq3_p & v23f74bc | !hbusreq3_p & v23fbe6a;
assign v22fc979 = hgrant5_p & v230a989 | !hgrant5_p & v230fdb8;
assign v23fcc70 = hbusreq1_p & b9d00f | !hbusreq1_p & v22ef56f;
assign v23fbb0b = hbusreq5 & v23fcfb8 | !hbusreq5 & v22f5583;
assign v22f1b3b = hlock6_p & v2391d0b | !hlock6_p & v84561b;
assign v22fabaf = jx3_p & v23fc60e | !jx3_p & v230e880;
assign v94778a = hmaster0_p & v230d6ca | !hmaster0_p & v22eff51;
assign v22f6b3e = hbusreq4 & v23045f5 | !hbusreq4 & v84561b;
assign v23fc7f5 = hgrant0_p & v22f878c | !hgrant0_p & v22f2639;
assign v2303ee8 = stateG10_5_p & v23f5d6f | !stateG10_5_p & v2306c80;
assign v23045fa = hmaster0_p & v23fc808 | !hmaster0_p & v22ede8c;
assign v23f4e36 = hmastlock_p & v2392897 | !hmastlock_p & v84561b;
assign v23fb9d0 = hmaster2_p & v22f954f | !hmaster2_p & v23f8036;
assign v23fcc2e = hmaster2_p & v2310d04 | !hmaster2_p & v84561b;
assign v23f1cdf = jx0_p & v22ff483 | !jx0_p & a090d5;
assign v23fcca1 = hgrant3_p & v230a71c | !hgrant3_p & v2310731;
assign v2301992 = hmaster0_p & v23fbed7 | !hmaster0_p & !v22efeb6;
assign v2311ed2 = hmaster0_p & v23fb7c3 | !hmaster0_p & v22f91ef;
assign v230219b = locked_p & v84561b | !locked_p & v22f7f74;
assign v23fca1c = hmaster2_p & v22ed65e | !hmaster2_p & v2311c4d;
assign v2301937 = hmaster0_p & v22f6dee | !hmaster0_p & v230fe82;
assign v22efb8e = hlock3_p & v22f2286 | !hlock3_p & !v84561b;
assign v231196d = hlock3_p & v23fb095 | !hlock3_p & fc8f81;
assign v2309aca = hgrant4_p & v84561b | !hgrant4_p & !v2302c42;
assign v23fc30d = hmaster2_p & v22f85a0 | !hmaster2_p & v22f9089;
assign v22eddf2 = hbusreq6_p & v23037d3 | !hbusreq6_p & v23fb5d7;
assign v23fc926 = hgrant2_p & v84564d | !hgrant2_p & !v84561b;
assign v22ffffd = hbusreq4 & v23f15ac | !hbusreq4 & v84561b;
assign v22ee43f = hmaster0_p & v22f3ac3 | !hmaster0_p & v22f6edc;
assign v8d07e3 = hmaster1_p & v22f160c | !hmaster1_p & v23fb877;
assign v230d235 = hbusreq3_p & v23fc083 | !hbusreq3_p & !v22f0dc3;
assign v23fcee2 = hbusreq2 & v23f0fd1 | !hbusreq2 & v9526ac;
assign v23f4ad7 = jx2_p & v23fc9eb | !jx2_p & v22ef7a7;
assign v23fcaf1 = hbusreq1_p & v23fbedf | !hbusreq1_p & v84561b;
assign v23fc361 = hbusreq1 & v22f3643 | !hbusreq1 & v84561b;
assign v23fc932 = hbusreq6 & v230f0de | !hbusreq6 & v230aa7a;
assign v23fb90a = hbusreq3 & v231025b | !hbusreq3 & v23fba9a;
assign v22f1d96 = hmaster2_p & v2308d79 | !hmaster2_p & v2306220;
assign v23f173d = hmaster0_p & v230b7fc | !hmaster0_p & !v2303115;
assign v22f1a14 = hgrant3_p & v23fc58b | !hgrant3_p & v23f43d6;
assign v230334d = hbusreq4_p & v23fc364 | !hbusreq4_p & v2308669;
assign v23fb9c9 = hmaster1_p & v23fd010 | !hmaster1_p & v231304d;
assign v23040f3 = hbusreq5 & v23f5140 | !hbusreq5 & v23fcfcc;
assign v22f8f3d = hbusreq1 & v2301505 | !hbusreq1 & v84561b;
assign v23fbc64 = hbusreq6_p & v23097f5 | !hbusreq6_p & v23fc27a;
assign v106a831 = hmaster0_p & v22ed975 | !hmaster0_p & !v96c563;
assign v23f8da8 = hready & v2300755 | !hready & !v84561b;
assign v22febe1 = hready & v21b35f9 | !hready & !v84561b;
assign v23013a6 = hmaster2_p & v84564d | !hmaster2_p & v23fbb80;
assign v22ecfe0 = hbusreq2 & v22f3643 | !hbusreq2 & v84561b;
assign v22f5fb8 = hgrant0_p & v230f480 | !hgrant0_p & !v23f908f;
assign v23fbedd = hmaster1_p & v84561b | !hmaster1_p & v22f947f;
assign v12cd9cd = hmastlock_p & v2309263 | !hmastlock_p & !v84561b;
assign v23934e0 = hbusreq0 & v23fbb1c | !hbusreq0 & v23f4462;
assign v23f2873 = hmaster2_p & v1aae29a | !hmaster2_p & !v191ae42;
assign v23fc4d3 = hgrant1_p & v845635 | !hgrant1_p & v231258e;
assign v23f53c1 = jx1_p & v23fc8e6 | !jx1_p & v22fcf35;
assign v2310d59 = hgrant3_p & v22efb8e | !hgrant3_p & !v84561b;
assign v23f243b = hgrant5_p & v230d61c | !hgrant5_p & v22ff58f;
assign v23fc51c = hgrant1_p & v230935d | !hgrant1_p & v23123b4;
assign v23fbb99 = hbusreq3_p & v2308955 | !hbusreq3_p & v23fc106;
assign v23fbf83 = hgrant6_p & v23fbdf8 | !hgrant6_p & v23fcf6b;
assign v23f4928 = hmaster1_p & v84561b | !hmaster1_p & v2306b99;
assign v230f046 = hbusreq1_p & v22eece2 | !hbusreq1_p & !v2308b19;
assign v23fb9d9 = hmaster0_p & v23f7af2 | !hmaster0_p & v22f46b1;
assign v230a02b = hmaster0_p & v2303e9a | !hmaster0_p & v22ffdf8;
assign v230f911 = hbusreq3_p & v23fcf21 | !hbusreq3_p & !v84562e;
assign v23fc87a = hmaster0_p & a25b7d | !hmaster0_p & v23fc4c2;
assign v2304aae = hmaster0_p & v22f56a5 | !hmaster0_p & v2306088;
assign v2309dca = hbusreq4 & v2306f5b | !hbusreq4 & e1bfb3;
assign v23fc22f = hbusreq6 & b06cee | !hbusreq6 & !v84561b;
assign v23fcec1 = hbusreq3_p & v23fcb24 | !hbusreq3_p & v84561b;
assign bc5d21 = hgrant5_p & v23fbe81 | !hgrant5_p & v230e311;
assign v23fc2e0 = hbusreq0 & v23fb1a4 | !hbusreq0 & !v84561b;
assign v23087f2 = hbusreq1 & v22f518e | !hbusreq1 & v84561b;
assign v23fcdcb = hmaster1_p & v23fc88f | !hmaster1_p & v23fbd21;
assign v2302c88 = hbusreq3_p & v230b49b | !hbusreq3_p & v22ff257;
assign v23135fa = hgrant1_p & v23fb6ff | !hgrant1_p & v23f880f;
assign v22fde5c = hmaster2_p & v191aa68 | !hmaster2_p & v22eaaba;
assign v8f8537 = hbusreq1 & v22fe421 | !hbusreq1 & v84561b;
assign v23f7114 = stateG2_p & v84561b | !stateG2_p & v23fb0ea;
assign v23fcf92 = hlock0_p & v2306b74 | !hlock0_p & !v239379c;
assign v2306bfb = hbusreq3_p & v2305aa9 | !hbusreq3_p & !v23f39e6;
assign v23f616b = hbusreq1 & v2312f7e | !hbusreq1 & !v22f91c9;
assign v23fb8c7 = hmaster2_p & v84564d | !hmaster2_p & a1fd0b;
assign v23fba85 = hbusreq6 & v23fc41e | !hbusreq6 & v230aca2;
assign v23f0db7 = hbusreq4 & v23036a1 | !hbusreq4 & v84561b;
assign v22fafef = hmaster1_p & v2312301 | !hmaster1_p & v22fd83a;
assign v230702c = hbusreq6_p & v239174b | !hbusreq6_p & v2311da1;
assign v239288d = hbusreq3 & v23fba94 | !hbusreq3 & v84561b;
assign v230ced0 = hmaster2_p & v23f6cef | !hmaster2_p & v22f7e59;
assign v230ce60 = hgrant1_p & v22f3643 | !hgrant1_p & v23fb952;
assign v231182b = hmaster0_p & v2301190 | !hmaster0_p & v23f5fd9;
assign v22f4bc7 = hmaster0_p & v2308967 | !hmaster0_p & v22f8838;
assign v23f6588 = hbusreq3 & v23128ab | !hbusreq3 & v2300df6;
assign fc907f = hbusreq3_p & v22f5e97 | !hbusreq3_p & v239353f;
assign v22f79a5 = hbusreq4_p & v23fce02 | !hbusreq4_p & v23f664b;
assign v2307d30 = hgrant3_p & v23fba81 | !hgrant3_p & !v84561b;
assign a8d315 = hlock5_p & v84561b | !hlock5_p & v23fbca4;
assign b1e86b = hbusreq6 & v230be4a | !hbusreq6 & v23f38c4;
assign v2303d87 = hmaster0_p & v84561b | !hmaster0_p & !v22eb3fd;
assign v23fc297 = hmaster0_p & v230b7fc | !hmaster0_p & v23035ba;
assign v2303b6a = hbusreq1_p & v23f9593 | !hbusreq1_p & v84561b;
assign v23fc39d = hbusreq4_p & v2300834 | !hbusreq4_p & v23084cc;
assign v22ee959 = stateA1_p & v84561b | !stateA1_p & v23fca93;
assign v22ee3e8 = hgrant4_p & v84561b | !hgrant4_p & !v230abf9;
assign v23fb76c = hready_p & v23098ce | !hready_p & v23102b2;
assign v22fb31a = jx0_p & v22ee9d2 | !jx0_p & !v23f623e;
assign v23036c1 = hgrant1_p & v84561b | !hgrant1_p & v22f349c;
assign v22fbd02 = hlock1_p & v23f8da8 | !hlock1_p & !v84561b;
assign v22efce2 = hmaster2_p & v23fc38f | !hmaster2_p & v23ef8bb;
assign v23f1609 = jx1_p & v23fc747 | !jx1_p & !v2393efc;
assign v845625 = hbusreq1_p & v84561b | !hbusreq1_p & !v84561b;
assign v2300d1d = hbusreq5 & v23fcedd | !hbusreq5 & v84561b;
assign v23fa215 = hmaster2_p & v2367a45 | !hmaster2_p & v9442ad;
assign v23fbf68 = hbusreq4 & v2310f77 | !hbusreq4 & a6db07;
assign v23064e4 = hbusreq1 & v23022b1 | !hbusreq1 & !v84561b;
assign v23fb489 = hbusreq5_p & a1fba6 | !hbusreq5_p & v230972f;
assign v22f4f40 = hbusreq5 & v230358b | !hbusreq5 & v22f8d74;
assign v22ec92f = hlock5_p & bbc337 | !hlock5_p & !v23fc9cb;
assign v22f01c5 = hbusreq1_p & v23046b5 | !hbusreq1_p & v22f5039;
assign v22f3f2d = hbusreq1_p & v23fc047 | !hbusreq1_p & v23f53e4;
assign v230848d = hgrant0_p & v9bc7cb | !hgrant0_p & !v84561b;
assign v230df7b = hbusreq1 & v23f6b67 | !hbusreq1 & v84561b;
assign v230ef1c = hlock1_p & v23f841d | !hlock1_p & !v84561b;
assign v23fcb31 = hbusreq3 & v2305d92 | !hbusreq3 & v84561b;
assign v22fbfe5 = hgrant0_p & v23f646e | !hgrant0_p & v2300d51;
assign v23fce4e = hbusreq3 & v23f004a | !hbusreq3 & v84561b;
assign v23fcc31 = hbusreq5 & v22f60c6 | !hbusreq5 & v84564d;
assign v23f2bbf = hmaster2_p & v230031f | !hmaster2_p & !v2300934;
assign v22ed1b5 = hmaster2_p & v23f7700 | !hmaster2_p & v23fcda9;
assign v191afde = hbusreq4_p & v2391a4f | !hbusreq4_p & v22f6f0c;
assign v23085b7 = hmaster1_p & v23f4be7 | !hmaster1_p & !v23fcf99;
assign v23f7933 = hbusreq4 & v23fb4cd | !hbusreq4 & !v230c15a;
assign v191ab30 = hbusreq1_p & v2309943 | !hbusreq1_p & v23f8017;
assign v23f6a42 = hbusreq4_p & v22fa202 | !hbusreq4_p & !v84561b;
assign b16326 = hgrant0_p & v22f878c | !hgrant0_p & v22fb5f7;
assign v23f1afd = hbusreq6 & v22f9f88 | !hbusreq6 & v22eeece;
assign v22ff50f = hbusreq3_p & v23112a4 | !hbusreq3_p & acdb9d;
assign v23f7ef4 = hlock6_p & v230fe14 | !hlock6_p & v8bc4e1;
assign v22fe260 = stateG10_5_p & v22f533e | !stateG10_5_p & v23fcf46;
assign v2300c5a = hgrant0_p & v23133fa | !hgrant0_p & v22f68fe;
assign v231016f = hmaster1_p & v84561b | !hmaster1_p & v23133be;
assign v230c65f = hmaster2_p & v22f8d74 | !hmaster2_p & v84561b;
assign v1507009 = hgrant1_p & v230aaa7 | !hgrant1_p & v22f4593;
assign v23fcd9b = hbusreq6_p & v230b93b | !hbusreq6_p & !v23fcae1;
assign v2307c15 = hmaster0_p & v231354e | !hmaster0_p & v2306d22;
assign v23f4c8c = hbusreq1_p & v230446f | !hbusreq1_p & !v23f5218;
assign v23125fd = hbusreq1 & v2393ac5 | !hbusreq1 & v22ef816;
assign v12cda11 = hmaster2_p & v2310bf5 | !hmaster2_p & a1fbcb;
assign v22fd79d = hbusreq3 & v2309eb8 | !hbusreq3 & !v84561b;
assign v230fbb3 = hmaster1_p & v15074d0 | !hmaster1_p & !v22f1d85;
assign v22fd152 = hgrant3_p & v230965a | !hgrant3_p & b84511;
assign ac10e3 = hbusreq4_p & v23074dd | !hbusreq4_p & v22ed0f0;
assign v22f1040 = hbusreq5_p & v22f41ee | !hbusreq5_p & v23fc636;
assign v23f5cfd = hbusreq5_p & v9526ac | !hbusreq5_p & v22f8986;
assign v22f771b = hbusreq4_p & v23fbe99 | !hbusreq4_p & v22f0ea8;
assign v23f3f36 = hbusreq6_p & v22faa39 | !hbusreq6_p & v23037b3;
assign v23fc808 = hbusreq6 & v22ef9f7 | !hbusreq6 & v84561b;
assign v2393d28 = hbusreq3 & v23fb89b | !hbusreq3 & !v845645;
assign v23fb8d7 = jx0_p & v23f1609 | !jx0_p & !v23f8299;
assign v23fb25c = hbusreq0_p & v23fc2fd | !hbusreq0_p & v845629;
assign v22fede6 = hmaster2_p & v2304962 | !hmaster2_p & v84561b;
assign v23fcf6a = hbusreq4_p & v22fba10 | !hbusreq4_p & v22f42d3;
assign v22ef9df = hbusreq5 & v230eb8d | !hbusreq5 & !v84561b;
assign v23fc2b8 = hmaster2_p & v84561b | !hmaster2_p & v23f9682;
assign v22eec0e = hgrant1_p & v22f6b45 | !hgrant1_p & v23f1cd2;
assign v98151e = hmaster0_p & v23fcbd0 | !hmaster0_p & v23fba6c;
assign v22f8be5 = hmaster2_p & v2306d29 | !hmaster2_p & v23fc127;
assign v23f7073 = hgrant4_p & v84561b | !hgrant4_p & v23fc3f6;
assign v23fcbd3 = hlock0_p & v22f4ace | !hlock0_p & v230b913;
assign v23fbf27 = hgrant3_p & v23fc95a | !hgrant3_p & v2304b05;
assign v1aadd09 = jx2_p & v23fc403 | !jx2_p & v23065d6;
assign v23f2298 = jx1_p & v22f09a2 | !jx1_p & v23f029a;
assign v22fd747 = hbusreq0 & v23fa8aa | !hbusreq0 & v22ffc44;
assign v23fc60b = hmaster2_p & v23fc4f8 | !hmaster2_p & v22f4163;
assign v191aeb3 = hgrant3_p & v22ff6c5 | !hgrant3_p & v2307d0e;
assign v230e4da = hgrant3_p & v23fc4e0 | !hgrant3_p & v1aad8c1;
assign v230f63f = hbusreq2_p & v2306d29 | !hbusreq2_p & v106af73;
assign v230306f = hgrant3_p & v2301bdf | !hgrant3_p & v22fc4a3;
assign v230dacd = hbusreq3 & bda69e | !hbusreq3 & v84561b;
assign v23efa39 = hmaster2_p & v106a782 | !hmaster2_p & v845661;
assign v23f8a97 = hmaster2_p & a1fba6 | !hmaster2_p & v22eb377;
assign a48bb0 = hmaster0_p & v22f9403 | !hmaster0_p & v2305a37;
assign v23f2a25 = hmaster0_p & v22f4989 | !hmaster0_p & v22fa768;
assign v23fc17b = hlock1_p & v22ece6c | !hlock1_p & v23fc726;
assign v22f4af1 = hbusreq4 & v23046be | !hbusreq4 & v23f91bc;
assign v23f7aa3 = hbusreq0_p & v22ed85a | !hbusreq0_p & v84564d;
assign v22f959d = hbusreq6 & v23f7423 | !hbusreq6 & v230875f;
assign v892c49 = hbusreq6 & v22fcf46 | !hbusreq6 & v84561b;
assign v23fc0bc = hgrant5_p & v22f049f | !hgrant5_p & v22eb2f1;
assign v230e897 = hgrant5_p & v23fc7d7 | !hgrant5_p & v2305de3;
assign v2302dd1 = hburst1 & v23fc8a3 | !hburst1 & v22fa5b4;
assign v230b2a1 = hgrant4_p & v84561b | !hgrant4_p & !v845655;
assign v230aedf = hbusreq6 & v23f2d39 | !hbusreq6 & v22f5fb4;
assign v22fe9e0 = hmastlock_p & v23f4096 | !hmastlock_p & !v84561b;
assign v22f4bcf = jx3_p & v22ee2eb | !jx3_p & v23fb8fd;
assign v106a7a0 = hmastlock_p & v22f91f3 | !hmastlock_p & !v84561b;
assign v23f54ac = hgrant2_p & v845629 | !hgrant2_p & !v84561b;
assign v12cc2ef = hbusreq1_p & v84561b | !hbusreq1_p & v23f5526;
assign v23fb63c = hbusreq3_p & v2308b2f | !hbusreq3_p & v230ca2b;
assign v23fd02c = hmaster2_p & a1fba6 | !hmaster2_p & v1506fe9;
assign v23fb9c2 = hbusreq2_p & v1aae56f | !hbusreq2_p & v106ae21;
assign v2306944 = hbusreq4 & v23fb8e0 | !hbusreq4 & v23fa2f1;
assign v22f6265 = hlock3_p & v22f9b00 | !hlock3_p & v23f6d92;
assign v230297f = hbusreq5_p & v845636 | !hbusreq5_p & v23fbe9a;
assign v23f4d0d = hbusreq5_p & v22f6c36 | !hbusreq5_p & !v84561b;
assign v22f05a0 = hbusreq1_p & v23f688e | !hbusreq1_p & !v106ae19;
assign c1f7e4 = hbusreq6 & v23fbe18 | !hbusreq6 & !v150718d;
assign v22eef9f = hgrant3_p & v22f8b41 | !hgrant3_p & v191b041;
assign v23f8274 = hbusreq5 & v84561b | !hbusreq5 & !v23f6bf0;
assign v2311302 = hbusreq3_p & v230a919 | !hbusreq3_p & v23fb12f;
assign v23fbc71 = hgrant4_p & v84561b | !hgrant4_p & v22f1841;
assign v23fba52 = hbusreq4_p & v22fe56f | !hbusreq4_p & v23006a1;
assign v23f3115 = hgrant0_p & v845622 | !hgrant0_p & v23fc93e;
assign v23fb7b2 = hgrant3_p & v23f5066 | !hgrant3_p & v2312401;
assign v2300d0f = hgrant3_p & v2301f9a | !hgrant3_p & v230dd35;
assign v23fcc8f = hbusreq4_p & v23fa460 | !hbusreq4_p & v23fc04e;
assign v23fc891 = hbusreq4_p & v22f908b | !hbusreq4_p & v23fc76e;
assign v22f5d73 = hlock3_p & v23facd7 | !hlock3_p & v23f441d;
assign v23f7d9f = hbusreq3 & v23f55ae | !hbusreq3 & v8c25df;
assign v23fca14 = hlock6_p & v9b33d9 | !hlock6_p & v23fcef8;
assign v22f0e2f = hmaster2_p & v23fb6e3 | !hmaster2_p & v22ee9ac;
assign v230875f = hgrant3_p & v2309cdc | !hgrant3_p & v2305b70;
assign v23fb671 = hmaster2_p & v22f9911 | !hmaster2_p & v2307150;
assign v22f30df = hbusreq1_p & v2301511 | !hbusreq1_p & v23fa2ec;
assign v23fc99f = hbusreq5_p & v230b59f | !hbusreq5_p & v23fc19c;
assign v23f7b33 = hbusreq1 & v23fa63b | !hbusreq1 & !v2311072;
assign v22eb701 = hmaster0_p & e1d75b | !hmaster0_p & v22ffab6;
assign bab0c9 = hgrant5_p & v23fbe4d | !hgrant5_p & !v23f9773;
assign v23fb699 = hmaster2_p & v2310d04 | !hmaster2_p & v2303b6a;
assign v23fc4e8 = hbusreq1_p & v230ea6d | !hbusreq1_p & !v2310c6d;
assign v22fafa3 = hbusreq1_p & v22f4864 | !hbusreq1_p & v84561b;
assign v22eea63 = hbusreq5 & v22fc091 | !hbusreq5 & v22f5583;
assign v22f248e = hmaster0_p & v23027b1 | !hmaster0_p & v22f7fed;
assign v22f7861 = hbusreq3 & v22f0945 | !hbusreq3 & v84561b;
assign v23fc4b0 = hlock3_p & v22ed942 | !hlock3_p & v23fbd38;
assign v23112ad = hgrant1_p & v84561b | !hgrant1_p & v2306538;
assign v2307ab9 = hbusreq1_p & b50bc7 | !hbusreq1_p & v22fdb01;
assign v230664e = hbusreq3_p & v22f3196 | !hbusreq3_p & !v84561b;
assign b00a78 = hbusreq1_p & v22ef21f | !hbusreq1_p & v23133a7;
assign f40628 = hbusreq3 & v22fab02 | !hbusreq3 & v23079bc;
assign v2304c8b = hbusreq6_p & v230e9be | !hbusreq6_p & v22ec77a;
assign v22f9faa = hmaster2_p & v106a782 | !hmaster2_p & !v22ed035;
assign v22f04ac = hmaster0_p & v22ed9a9 | !hmaster0_p & v22ec20d;
assign v23f4963 = hbusreq2 & v13afe3a | !hbusreq2 & !v84561b;
assign v23fb818 = hmaster0_p & v2301105 | !hmaster0_p & v2312b9e;
assign v231261b = hbusreq4 & v22f8012 | !hbusreq4 & v22eaee7;
assign v23076e7 = hbusreq6 & v2307578 | !hbusreq6 & v22ebbab;
assign v22f5b7c = hbusreq4 & v22f0c90 | !hbusreq4 & v84561b;
assign v2307ab6 = jx1_p & v23f44e8 | !jx1_p & v230fbb3;
assign v230df19 = hgrant5_p & v230e7e3 | !hgrant5_p & v22f08be;
assign v22fba0e = hlock3_p & v22f6dfa | !hlock3_p & !v22f68f1;
assign v23fcf5e = hbusreq3_p & v230f578 | !hbusreq3_p & v22f8626;
assign v22ffba8 = hbusreq5_p & v23fbbb0 | !hbusreq5_p & v23f43cf;
assign v23fcd6d = jx3_p & v22fdb97 | !jx3_p & v230960d;
assign v23026ed = hgrant5_p & v23111c2 | !hgrant5_p & v23fc5a3;
assign v22f7e80 = hlock0_p & v84564d | !hlock0_p & v2301f3a;
assign v22fe22a = hbusreq3 & v230d90f | !hbusreq3 & v84561b;
assign v23fbd93 = hbusreq5_p & v23f5043 | !hbusreq5_p & v23fcb5c;
assign v23fc2f1 = hmaster0_p & v23fc802 | !hmaster0_p & v23f1109;
assign v23fad53 = hbusreq3 & v230cf2f | !hbusreq3 & v12cdba9;
assign v22f0cf9 = hbusreq4_p & v2302c02 | !hbusreq4_p & v84561b;
assign v23022c5 = hgrant5_p & v84561b | !hgrant5_p & v22f2817;
assign v22ec894 = hgrant1_p & v84561b | !hgrant1_p & v23fc519;
assign v22f235b = stateG2_p & v23023b3 | !stateG2_p & !v23fcb5d;
assign v2312cf2 = hbusreq0_p & v23fa2ec | !hbusreq0_p & v23fc4f8;
assign v23fb91a = hbusreq6_p & v23fc567 | !hbusreq6_p & v23fcddd;
assign v22f7f12 = jx1_p & v22fef14 | !jx1_p & v23f645e;
assign v22f0fe4 = hmaster2_p & v230c55d | !hmaster2_p & v22fb5da;
assign c0084f = hmaster2_p & v22fca28 | !hmaster2_p & v23f9682;
assign v23fab9b = hgrant5_p & v230bdd9 | !hgrant5_p & v23fcc22;
assign a8a256 = hmaster2_p & v106ae21 | !hmaster2_p & v23fb9c2;
assign v2393142 = hbusreq6_p & v23fc11b | !hbusreq6_p & v23fbace;
assign v23f76dc = hbusreq4 & v22fcf52 | !hbusreq4 & v22ee657;
assign v22fc7c1 = stateG10_5_p & v23fbc42 | !stateG10_5_p & v106af73;
assign v2308db0 = hmaster0_p & v23fc89b | !hmaster0_p & v2312b9e;
assign v23fc696 = hbusreq3_p & v22f483c | !hbusreq3_p & v23fba34;
assign v2391ab6 = hburst0_p & v84561b | !hburst0_p & v23021e1;
assign v230201b = hbusreq4_p & v23028be | !hbusreq4_p & v23f7950;
assign b5f51c = hbusreq2_p & v23f6411 | !hbusreq2_p & !v106ae19;
assign v23060a6 = hgrant0_p & v23fbb4e | !hgrant0_p & !v84561b;
assign v22faa24 = stateG10_5_p & v22ed127 | !stateG10_5_p & v845636;
assign v22efc50 = hgrant0_p & v2301e25 | !hgrant0_p & v23f280c;
assign v23fbfcb = hbusreq3_p & v23fc3f2 | !hbusreq3_p & v23f1891;
assign v23fcd9e = hbusreq1 & v22f2db0 | !hbusreq1 & v23fa2ec;
assign v23f20d0 = hbusreq4 & v23fbb98 | !hbusreq4 & v84561b;
assign a7b623 = hbusreq3_p & v23010f6 | !hbusreq3_p & v23f8f1d;
assign v23fb242 = hbusreq4_p & v230ec04 | !hbusreq4_p & v9ed019;
assign v23fc161 = hgrant1_p & v845626 | !hgrant1_p & v230c52a;
assign bc65c8 = hbusreq3 & v230eca1 | !hbusreq3 & v23f87f4;
assign v230caee = hgrant4_p & v22f5378 | !hgrant4_p & v22ece21;
assign v23f3073 = hmaster0_p & v22ffd0e | !hmaster0_p & v2391fb2;
assign v22ed741 = hgrant5_p & v23f47ca | !hgrant5_p & v23fcd29;
assign v230709c = hbusreq3 & v23018f2 | !hbusreq3 & v84561b;
assign v230eed2 = hmaster0_p & v22f636a | !hmaster0_p & v2301c02;
assign v22f1ef1 = hmaster2_p & v22f1796 | !hmaster2_p & v22ee8f3;
assign v230aa94 = hbusreq3_p & v23018f1 | !hbusreq3_p & v84561b;
assign v23fb8a0 = hgrant1_p & v230b8ff | !hgrant1_p & v22f0d2b;
assign v23f8486 = stateG2_p & v2306d5c | !stateG2_p & v2301d2f;
assign v230ecb6 = hbusreq4_p & v23f3501 | !hbusreq4_p & v22ebbf2;
assign v22f29e5 = hbusreq3_p & v23051f6 | !hbusreq3_p & v23f97a7;
assign v23fcf04 = hmaster1_p & v23fcb0e | !hmaster1_p & v2308d06;
assign v22f2e7b = hmaster2_p & v23101b1 | !hmaster2_p & v23f8e6b;
assign v22fe392 = hmaster2_p & v2309cdc | !hmaster2_p & v23f3997;
assign v2310b6a = hbusreq0 & v22f79fd | !hbusreq0 & v84561b;
assign v22fed5c = hmaster2_p & v84561b | !hmaster2_p & !v230eafe;
assign v23f0d8a = hgrant3_p & v22ecaf6 | !hgrant3_p & v23f77b1;
assign v22f0332 = hbusreq1_p & v23fc6d6 | !hbusreq1_p & v23faece;
assign v23fccb0 = hmaster2_p & v2310d6a | !hmaster2_p & v23fba9a;
assign v23fb139 = hlock6_p & v84564d | !hlock6_p & !v23f60ba;
assign v22fab30 = hgrant1_p & v22f035c | !hgrant1_p & v2305a79;
assign v23fce5f = hbusreq3_p & v230dcba | !hbusreq3_p & v22fb29c;
assign v2310c26 = hbusreq3 & v23fc0c6 | !hbusreq3 & v84561b;
assign v22ff090 = hready & v23fc491 | !hready & v230c899;
assign v23ef9c4 = hgrant2_p & v22ed898 | !hgrant2_p & v23fbb37;
assign v22fe657 = hgrant5_p & v84561b | !hgrant5_p & !v22f6ac3;
assign a54167 = jx0_p & v23fce39 | !jx0_p & !v22f2b59;
assign v23f92d5 = stateG10_5_p & v23f8c71 | !stateG10_5_p & v23f6bc1;
assign v23f1f21 = hbusreq5_p & v22f051d | !hbusreq5_p & v23f40ba;
assign v22f313c = hmaster0_p & v22f4266 | !hmaster0_p & v23f193e;
assign v22fd796 = hbusreq6_p & v23fbfe9 | !hbusreq6_p & v231096b;
assign v23fb9bf = hmaster0_p & v22fa0ec | !hmaster0_p & !v230200a;
assign v22f23a1 = hbusreq1_p & v84564d | !hbusreq1_p & v84561b;
assign v22ec702 = hbusreq6 & v22ffa4c | !hbusreq6 & v22f7347;
assign v2393f52 = hgrant0_p & v22f0ac0 | !hgrant0_p & !v22f69b7;
assign v23fcf71 = hgrant5_p & v22f481f | !hgrant5_p & v230d16b;
assign v23fbf0b = hmaster2_p & v84561b | !hmaster2_p & v22ff090;
assign v22f6a6e = hbusreq5_p & v22ef983 | !hbusreq5_p & !v22fcd0f;
assign v23fc458 = hgrant3_p & v84561b | !hgrant3_p & !v22f7ed8;
assign v22f7dc7 = stateG10_5_p & b16326 | !stateG10_5_p & v22f878c;
assign v22f3c27 = hmaster2_p & v22f1ece | !hmaster2_p & !v23fa345;
assign v23fc105 = hbusreq1_p & v230928c | !hbusreq1_p & v845635;
assign v23fb8de = jx0_p & v22fc365 | !jx0_p & v22f0a7b;
assign v23f2bb9 = hmaster2_p & v2312025 | !hmaster2_p & a39dae;
assign v23fbb4b = hgrant1_p & v231350d | !hgrant1_p & v22fd50f;
assign v23018f1 = hbusreq3 & v23fb671 | !hbusreq3 & v84561b;
assign v1aae385 = hmaster2_p & v22f0860 | !hmaster2_p & v23fb966;
assign v230887b = hbusreq6_p & v23fc3f3 | !hbusreq6_p & v23fbfb2;
assign v230be9e = hbusreq6_p & v22faa19 | !hbusreq6_p & v23fc94d;
assign v23068f2 = hbusreq3_p & v22fa6f5 | !hbusreq3_p & v2309d23;
assign v2305aa1 = hburst0_p & v84561b | !hburst0_p & !v845649;
assign v2306667 = hmastlock_p & v22f39a1 | !hmastlock_p & v84561b;
assign v22f9049 = hbusreq5_p & v23fc904 | !hbusreq5_p & !v2307646;
assign v22f536a = hlock3_p & v2312053 | !hlock3_p & bd9dce;
assign v2306e3c = hmaster0_p & v23fb73d | !hmaster0_p & v22f444f;
assign v22fc6b9 = hbusreq3_p & v22f0a24 | !hbusreq3_p & v23fcc3d;
assign v22f4b91 = hbusreq6 & v22fb00c | !hbusreq6 & !v845625;
assign v23f8e93 = hbusreq5 & v23f2c89 | !hbusreq5 & v22f7929;
assign v23f5d6f = hgrant0_p & v23fc4fd | !hgrant0_p & v23fbcfc;
assign a1fe5a = hbusreq4_p & ad6e26 | !hbusreq4_p & v23f608b;
assign v22f517c = hmaster0_p & v23fc761 | !hmaster0_p & !v22ee91d;
assign v2308cec = hmaster2_p & v23036c1 | !hmaster2_p & v2303cc1;
assign v23f38d5 = hmaster2_p & v23fbe41 | !hmaster2_p & !v84561b;
assign v2303e23 = hmaster2_p & v84561b | !hmaster2_p & v23f1879;
assign v23fcd0a = hgrant1_p & v84561b | !hgrant1_p & v22f8629;
assign v23934cb = hmaster1_p & v22ef255 | !hmaster1_p & !v22f288d;
assign v230bf27 = hbusreq3_p & v2311a27 | !hbusreq3_p & v22f97fe;
assign v22fdc16 = hmaster0_p & v22f15e8 | !hmaster0_p & !v2309dca;
assign v23fc870 = hgrant1_p & v84561b | !hgrant1_p & v1b8769e;
assign v23fb910 = hlock3_p & v22faef4 | !hlock3_p & v22fb759;
assign v230287e = hbusreq0 & v23fbfd0 | !hbusreq0 & v22f11f6;
assign v2312a9e = start_p & v84561b | !start_p & !v845665;
assign v2310538 = hgrant3_p & v84564d | !hgrant3_p & !v84561b;
assign v22f37c1 = hmastlock_p & v22ebffc | !hmastlock_p & v84561b;
assign v230adbf = hmaster0_p & v22f6169 | !hmaster0_p & v23f781b;
assign v230ac1b = hbusreq6 & v23f9ae7 | !hbusreq6 & !v84561b;
assign v22f8afa = hmaster2_p & v230c910 | !hmaster2_p & v231025b;
assign v230dfa0 = hmaster0_p & v2392d61 | !hmaster0_p & !v22f45d7;
assign v23fc281 = hbusreq4 & v23019e9 | !hbusreq4 & v84561b;
assign v230b781 = hbusreq6 & v22f0102 | !hbusreq6 & v84561b;
assign v23f56b1 = hbusreq4_p & v84561b | !hbusreq4_p & v231254f;
assign v22ee274 = jx2_p & v23056b2 | !jx2_p & v230e3d1;
assign v2306785 = hlock0_p & v13aff5b | !hlock0_p & v23059d8;
assign v23fa875 = hbusreq1_p & v23fc40f | !hbusreq1_p & v2393b5a;
assign v22f3206 = hmaster2_p & a07f9b | !hmaster2_p & v23fcb69;
assign v23f082a = hbusreq4 & v23fbe8e | !hbusreq4 & v230fce3;
assign v23fa2d6 = hmaster2_p & v22ef513 | !hmaster2_p & v23fc017;
assign v23fc7e3 = hmaster2_p & a1fba6 | !hmaster2_p & v22f4f42;
assign v23fbbc2 = hbusreq1_p & v23126de | !hbusreq1_p & v23f7796;
assign v230a989 = hbusreq5_p & v2306609 | !hbusreq5_p & v23035a3;
assign v22ebeb2 = hgrant3_p & v230727f | !hgrant3_p & v22ff50f;
assign v22f7c2b = hmaster0_p & v22f9d92 | !hmaster0_p & v22f7022;
assign v22f3a6f = stateG10_5_p & v23005e2 | !stateG10_5_p & v12cd4c6;
assign v22f06fc = hbusreq0_p & v23fc93e | !hbusreq0_p & v22fbda1;
assign v231210f = hbusreq4_p & v230f0de | !hbusreq4_p & v22edbd4;
assign v22f49e4 = hgrant2_p & v84561b | !hgrant2_p & v23fc5f4;
assign v2304578 = hbusreq3_p & v23fcea8 | !hbusreq3_p & !v23f946b;
assign v22ed01d = hlock3_p & v22ef026 | !hlock3_p & v23fbd38;
assign v2312eaa = hbusreq4 & v2305a09 | !hbusreq4 & v23fba11;
assign v230d6b6 = hbusreq3_p & v2306844 | !hbusreq3_p & v230a226;
assign v22f244d = hmaster1_p & v23f6042 | !hmaster1_p & v23fb9d3;
assign v22fcc78 = hgrant3_p & v22fcea7 | !hgrant3_p & v23fcecc;
assign v23049d7 = hbusreq3_p & v23070c0 | !hbusreq3_p & v23fb22d;
assign v230fd1d = hlock3_p & v22fbb33 | !hlock3_p & v22f16bf;
assign v22ec77a = hbusreq6 & v845620 | !hbusreq6 & v84561b;
assign v22fe62b = hbusreq5_p & v22fef4f | !hbusreq5_p & a1fe27;
assign v23642d5 = hbusreq6 & v22f9b6f | !hbusreq6 & v23fca08;
assign v23fa5d4 = hbusreq3 & v22f023b | !hbusreq3 & v23fca20;
assign v2309be5 = hmaster2_p & v23fa2ec | !hmaster2_p & !v22ec921;
assign v23fafca = hbusreq3 & v23fb9c6 | !hbusreq3 & v2311214;
assign v22ee10b = hbusreq3_p & v22edf4f | !hbusreq3_p & v23fbcc4;
assign v23fc4f8 = hbusreq2_p & v230eef7 | !hbusreq2_p & v845620;
assign v22fb802 = hgrant3_p & v84561b | !hgrant3_p & v22f0b42;
assign v230dcba = hmaster2_p & v2391b88 | !hmaster2_p & v23f9680;
assign v23fbf54 = hbusreq6_p & v2391fc6 | !hbusreq6_p & v230abc9;
assign v23fce10 = hbusreq3 & v23fc8f8 | !hbusreq3 & v84561b;
assign v84563a = hbusreq6 & v84561b | !hbusreq6 & !v84561b;
assign v23017ee = hbusreq1_p & v23f0bd2 | !hbusreq1_p & v2304bc1;
assign v230717d = jx0_p & v23fc42e | !jx0_p & d49f32;
assign v23f2f5d = hbusreq3_p & v2310c26 | !hbusreq3_p & v84561b;
assign v23084c2 = stateG10_5_p & v2310da0 | !stateG10_5_p & v2303393;
assign v22ec326 = hmaster2_p & v22f6cec | !hmaster2_p & !v84561b;
assign v23fb636 = hbusreq1_p & v23fa9d0 | !hbusreq1_p & !v84561b;
assign v22ff114 = hmaster0_p & v2312189 | !hmaster0_p & v2382e8c;
assign v230538c = hbusreq3_p & v22ff21b | !hbusreq3_p & !v1aad4c6;
assign v23f2f40 = hbusreq4_p & v2308bfc | !hbusreq4_p & v22f2e20;
assign v23f7db2 = hmaster2_p & v22ec89f | !hmaster2_p & v22f66cf;
assign a4e378 = hbusreq3_p & v22f3982 | !hbusreq3_p & v84561b;
assign v22f4855 = hgrant3_p & v22f6ae5 | !hgrant3_p & v230dcef;
assign v22fb40c = jx1_p & v230a688 | !jx1_p & v23fc5ce;
assign v22f446e = hgrant2_p & v22f2f87 | !hgrant2_p & !v2304ec7;
assign v22f0360 = hgrant0_p & v84561b | !hgrant0_p & !v23f9ca2;
assign bd7bf6 = stateG10_5_p & v23fc85a | !stateG10_5_p & v845636;
assign v23f1e3f = hbusreq3 & v22f6741 | !hbusreq3 & v84561b;
assign v230a3ec = hmastlock_p & v22ee0e1 | !hmastlock_p & v84561b;
assign v23fc95c = hgrant3_p & v84561b | !hgrant3_p & v23fc027;
assign v23fbc7d = stateG2_p & v84561b | !stateG2_p & !v23fcdc4;
assign v23f9ee2 = hgrant5_p & v84561b | !hgrant5_p & v22f517e;
assign v23fcdce = hgrant5_p & v84561b | !hgrant5_p & v23f19b4;
assign v2303ce2 = stateG10_5_p & v23fc1c8 | !stateG10_5_p & !v230f848;
assign da38ba = hmaster2_p & v23fc796 | !hmaster2_p & v1507529;
assign v231141f = hbusreq3_p & v23fce31 | !hbusreq3_p & v22fd41b;
assign v22fad0f = hbusreq6 & v22ec890 | !hbusreq6 & v22eca65;
assign v22f8c01 = hmaster0_p & v23f38b7 | !hmaster0_p & v22ff21b;
assign v22ef9db = hbusreq3_p & v2304f4c | !hbusreq3_p & !v2304b49;
assign adb81d = hgrant5_p & v231200e | !hgrant5_p & v23f1ca8;
assign v22f5820 = hready & abfa28 | !hready & !v84561b;
assign v230f375 = hbusreq3_p & v23fcbdb | !hbusreq3_p & v22ee1d1;
assign v22f3550 = hgrant3_p & v22eb51e | !hgrant3_p & v23fbcd4;
assign v1aad46b = hbusreq3 & v2305a2a | !hbusreq3 & v84561b;
assign v230df30 = hgrant0_p & v22fa654 | !hgrant0_p & v22f8e10;
assign v23fb52d = hmaster2_p & v23fbaaa | !hmaster2_p & v15070fa;
assign v22fea3f = hlock3_p & v22eb664 | !hlock3_p & v23f60d2;
assign v2304421 = hgrant1_p & v84561b | !hgrant1_p & v22f7f2a;
assign v22f01b6 = hbusreq6_p & v1aae8d3 | !hbusreq6_p & v22f9396;
assign v23f8089 = hbusreq2 & v15071c2 | !hbusreq2 & !ab5bb8;
assign v22ef377 = hbusreq3_p & v23fbdc0 | !hbusreq3_p & f40628;
assign v23fc4df = hbusreq4_p & b59af9 | !hbusreq4_p & v23fbc1b;
assign v2308235 = hbusreq1 & v22eef57 | !hbusreq1 & v84561b;
assign v23fba3e = hgrant5_p & v2392842 | !hgrant5_p & v22fa711;
assign v214cf31 = hready_p & v230ec4b | !hready_p & !v845641;
assign v22f8499 = jx3_p & v2391cf8 | !jx3_p & v230cc50;
assign v22f178d = start_p & v84561b | !start_p & v230f4d3;
assign v22f1ece = hbusreq5 & v2306220 | !hbusreq5 & !v84561b;
assign v23fcce5 = hlock0_p & v22f037a | !hlock0_p & v22fe50f;
assign v22f7b24 = hmaster1_p & a878fd | !hmaster1_p & v2301f50;
assign v22ef217 = hgrant1_p & v17a34ff | !hgrant1_p & v1aad5c9;
assign v22f5e18 = hlock5_p & e1df2d | !hlock5_p & v84561b;
assign v1aae9e2 = hgrant5_p & v2306298 | !hgrant5_p & v23f2f42;
assign v22f8093 = hmaster2_p & v2313059 | !hmaster2_p & v230f537;
assign v22f3d18 = hbusreq4 & v22fd002 | !hbusreq4 & v22f13d8;
assign v23fbff0 = hbusreq6_p & v230ec2b | !hbusreq6_p & v22f7d33;
assign v22f848f = hmaster2_p & v23fb796 | !hmaster2_p & !v22f5b4b;
assign v2303f50 = hlock3_p & v2311094 | !hlock3_p & v22ec9b2;
assign v23f0b4e = hbusreq6_p & v230178e | !hbusreq6_p & v230521a;
assign bd94ed = hbusreq0_p & v84561b | !hbusreq0_p & !v2313463;
assign v22ee8d8 = hlock0_p & v22f264f | !hlock0_p & v23f4872;
assign v22f30be = hbusreq1 & v23027e9 | !hbusreq1 & v84561b;
assign v22ff9d7 = hgrant1_p & v84561b | !hgrant1_p & v22f62dc;
assign v23fc9dd = hbusreq1_p & v23fa623 | !hbusreq1_p & !v84561b;
assign v22ff0da = hmaster2_p & v23022b1 | !hmaster2_p & !v23027e9;
assign v2308815 = hmaster2_p & v1e83fd9 | !hmaster2_p & a1fbc2;
assign v22f263c = hmaster2_p & v23919f9 | !hmaster2_p & v22f6b4c;
assign v230cc50 = hmaster1_p & v23f7b85 | !hmaster1_p & !v23ef987;
assign v22ebd62 = stateG10_5_p & v2305522 | !stateG10_5_p & v22f3a35;
assign v23fcb87 = hlock3_p & v191a964 | !hlock3_p & v23fced0;
assign v22f1172 = jx1_p & v23fbb25 | !jx1_p & v23fbf9b;
assign v23f2b69 = hlock3_p & v22fe1ad | !hlock3_p & v22ff9c5;
assign v23fba13 = hbusreq0 & v2312f7e | !hbusreq0 & !v22f91c9;
assign v2301f50 = hmaster0_p & v22f725a | !hmaster0_p & v23fc943;
assign v23010f6 = hbusreq3 & v22f99e3 | !hbusreq3 & v23002bf;
assign v23fc5ba = hbusreq2_p & v22f9497 | !hbusreq2_p & !v845620;
assign v23fb136 = stateG2_p & v84561b | !stateG2_p & v2310c2b;
assign v230df28 = hbusreq4 & v23faa5c | !hbusreq4 & v2301a04;
assign v22fb88d = hbusreq6 & v845620 | !hbusreq6 & v23fba11;
assign v2303046 = hlock5_p & da38bd | !hlock5_p & !v84561b;
assign v23f4572 = hgrant1_p & v84561b | !hgrant1_p & v22f06ac;
assign v2312a3d = hbusreq3 & v23fbdc1 | !hbusreq3 & v2313131;
assign v23fbe0a = hlock5_p & v23fb8a7 | !hlock5_p & e1dcf4;
assign v230d66e = hlock6_p & v2309192 | !hlock6_p & v230a58f;
assign v2310482 = hmaster2_p & v230eb9b | !hmaster2_p & v23f5c95;
assign v23f4f2c = hbusreq4_p & e1c7f2 | !hbusreq4_p & v22fc2d0;
assign v22ee281 = hbusreq5_p & v84561b | !hbusreq5_p & v1aae087;
assign v23fca23 = hgrant5_p & v2307dbf | !hgrant5_p & v23fb0cd;
assign v23fc380 = hbusreq6_p & v23f496d | !hbusreq6_p & v22fabad;
assign e1e7a3 = hmaster2_p & v23fc921 | !hmaster2_p & v22f7b8b;
assign v22f8ccb = hbusreq5_p & v22f1b4e | !hbusreq5_p & !v22f3483;
assign v23f9714 = hbusreq4 & v23fb5b3 | !hbusreq4 & !v23fba99;
assign v23001c7 = hlock1_p & v84561b | !hlock1_p & v13afe3a;
assign v23fb62d = hbusreq4 & v23127ee | !hbusreq4 & v2303c5a;
assign v22f48ce = hbusreq3_p & v23fc3eb | !hbusreq3_p & v84561b;
assign v22ec20e = hlock4_p & v2391d0b | !hlock4_p & v84561b;
assign v23fcd7a = hbusreq3_p & v22f88ee | !hbusreq3_p & v84561b;
assign v23fb099 = hmaster2_p & v22ecba3 | !hmaster2_p & fc8c3f;
assign v22fe204 = hgrant1_p & v22fee46 | !hgrant1_p & v23001a4;
assign v84565b = hgrant6_p & v84561b | !hgrant6_p & !v84561b;
assign v23fcd13 = jx2_p & v23f4a0f | !jx2_p & v22fa4c3;
assign v23f1561 = hmaster0_p & v2311be2 | !hmaster0_p & !v2303598;
assign v2391c55 = hlock4_p & v230fdf7 | !hlock4_p & !v84561b;
assign v22fa86d = hmaster2_p & v84561b | !hmaster2_p & v22ebe03;
assign v23f48a1 = hbusreq6 & v22ee4d5 | !hbusreq6 & v84561b;
assign v22fd298 = hbusreq3_p & v23fb18e | !hbusreq3_p & v230c6c0;
assign v23fc0c2 = hbusreq5_p & v23f08e5 | !hbusreq5_p & v23fc5c7;
assign v22f2e9f = hbusreq3_p & v22f4d61 | !hbusreq3_p & v2306b9f;
assign v23f8036 = hgrant1_p & v230f63f | !hgrant1_p & v23f480d;
assign v239158d = hbusreq6_p & v23f5d1a | !hbusreq6_p & v2300dcb;
assign da38c1 = hmastlock_p & v23f61f7 | !hmastlock_p & v84561b;
assign v1aad535 = hbusreq3_p & v23fb661 | !hbusreq3_p & v230abb0;
assign v230c03a = hgrant0_p & v230bae0 | !hgrant0_p & v84561b;
assign v2313247 = hgrant1_p & v230031f | !hgrant1_p & v23057e6;
assign v22fb465 = hgrant3_p & v23fc318 | !hgrant3_p & v23113d2;
assign v230c041 = stateG2_p & v84561b | !stateG2_p & !v22f197e;
assign v23f8ade = hbusreq5 & v231228e | !hbusreq5 & !v84561b;
assign v1506add = hmaster2_p & v88c9bf | !hmaster2_p & v23fba9a;
assign v23fccaf = hmaster0_p & v23fcdd1 | !hmaster0_p & !v23fb7b2;
assign v22fce66 = hbusreq2_p & v2300711 | !hbusreq2_p & !v84561b;
assign v23fb5b7 = hbusreq3 & v22f8ba5 | !hbusreq3 & !v84561b;
assign v22ecd54 = hmaster2_p & a1fba6 | !hmaster2_p & v23f972e;
assign v230eca1 = hmaster2_p & v23fb49a | !hmaster2_p & v230e916;
assign v23139e3 = hmaster2_p & v23105b6 | !hmaster2_p & v22f8549;
assign v230da2f = hmaster2_p & v23f052e | !hmaster2_p & v22eb404;
assign e1e726 = hmaster2_p & v23fb5a1 | !hmaster2_p & v23fc741;
assign v22f619f = hbusreq1_p & v23fbd2e | !hbusreq1_p & v84564d;
assign v23fbea7 = hmaster0_p & v23f78a3 | !hmaster0_p & v23fc999;
assign v22f4627 = hlock3_p & v23fc67f | !hlock3_p & v2300bb5;
assign v23fc3ca = hgrant3_p & v23fc139 | !hgrant3_p & !v84561b;
assign v230741d = hmaster2_p & v22f7d5d | !hmaster2_p & v23f3d47;
assign v23fb98d = hburst1 & v84561b | !hburst1 & v2391f3b;
assign v23069f2 = stateG2_p & v23fcfa4 | !stateG2_p & v23f1316;
assign v22fdf30 = hmaster2_p & v84561b | !hmaster2_p & v2302e32;
assign v22f1427 = hbusreq1_p & v23fb85c | !hbusreq1_p & v23089ec;
assign v23fcbca = hbusreq1_p & v2309cb0 | !hbusreq1_p & v84561b;
assign v2393de1 = hgrant3_p & v23fcbc9 | !hgrant3_p & v23fbfca;
assign v23f4bcd = hready & v84561b | !hready & !v22fe9e0;
assign v23f558b = hmaster2_p & a1fba6 | !hmaster2_p & v9526ac;
assign v23fce88 = hmaster2_p & v191a876 | !hmaster2_p & !v2302e32;
assign v23fbbcf = stateG10_5_p & v230a9f0 | !stateG10_5_p & a1fba6;
assign v1aae206 = hbusreq3_p & v230391b | !hbusreq3_p & !v84561b;
assign v23f3adc = hgrant0_p & v22fc05f | !hgrant0_p & v23fb648;
assign v22ed8e2 = hlock6_p & v23f593d | !hlock6_p & v23038ea;
assign v23096af = jx1_p & v2304d0c | !jx1_p & v23fcc83;
assign v22f8d0c = hmaster2_p & v230e1f3 | !hmaster2_p & v22fd283;
assign v2393bce = hlock2_p & v22ed85a | !hlock2_p & v84561b;
assign v230c0b8 = hgrant1_p & v845620 | !hgrant1_p & v93dace;
assign v23fbe4c = hgrant0_p & v22fcbcd | !hgrant0_p & v106af4d;
assign v23046fe = hgrant6_p & v23fc8a1 | !hgrant6_p & v22f5f72;
assign v23fca4f = hbusreq0 & v23105cd | !hbusreq0 & v84561b;
assign v22eeb03 = hbusreq5_p & v23fcf46 | !hbusreq5_p & v23f646e;
assign v22f621f = hbusreq5 & v23f8364 | !hbusreq5 & !v84561b;
assign v2306c16 = hgrant5_p & v84561b | !hgrant5_p & v22fca4e;
assign v2303598 = hgrant3_p & v2393392 | !hgrant3_p & v23fb62b;
assign v230bae0 = hlock0_p & v22efd4a | !hlock0_p & v22ee9be;
assign v23f6250 = hlock1_p & v23fbc1d | !hlock1_p & v22f5f1c;
assign v2391bb7 = hlock0_p & v84561b | !hlock0_p & v230a63b;
assign v22fa48c = hbusreq5 & v22f3643 | !hbusreq5 & v84561b;
assign v979b7c = hgrant1_p & v22eec8b | !hgrant1_p & v2309c2c;
assign v22ed92a = jx2_p & v23fce16 | !jx2_p & v22fa4f7;
assign v22f0de0 = hlock3_p & v230c73d | !hlock3_p & !v22ff6a8;
assign v1507439 = hbusreq4_p & v22f95a4 | !hbusreq4_p & v23f69e4;
assign v23fcaa5 = hgrant3_p & v84561b | !hgrant3_p & v23f704d;
assign v230d5af = hbusreq6_p & v22fc531 | !hbusreq6_p & v230585c;
assign v1507317 = hmaster2_p & v23fc35a | !hmaster2_p & v22fc5fd;
assign v23084c9 = hbusreq5_p & v230154b | !hbusreq5_p & !v84561b;
assign v2300e95 = hmaster0_p & v23fcaad | !hmaster0_p & v22efd70;
assign v2307dbf = hbusreq5_p & v23fc828 | !hbusreq5_p & v23fac04;
assign v23fbc97 = hmaster2_p & v106a782 | !hmaster2_p & !v22ff120;
assign v22fb07c = hbusreq5 & v23fbb80 | !hbusreq5 & v84561b;
assign v845636 = hbusreq5 & v84561b | !hbusreq5 & !v84561b;
assign v23fb095 = hbusreq3_p & v2305d6e | !hbusreq3_p & v22faa4d;
assign v2307e0c = hmaster2_p & v23fbc3f | !hmaster2_p & a1fbc2;
assign v22feee5 = hlock1_p & v22f2822 | !hlock1_p & v845620;
assign v22ef962 = hbusreq4_p & v22ef9ff | !hbusreq4_p & v23fc36b;
assign v22f5898 = jx3_p & v22ed220 | !jx3_p & v23fbd3a;
assign v230beed = hbusreq1 & v1aae29a | !hbusreq1 & !v84561b;
assign v230754e = jx1_p & v23f7c5a | !jx1_p & v231228f;
assign v23060ff = hlock3_p & v191ac40 | !hlock3_p & v2304bc1;
assign v2306837 = hbusreq3_p & v23fb074 | !hbusreq3_p & v84561b;
assign v23fc617 = hmaster1_p & v23fc35e | !hmaster1_p & v23ef987;
assign v23fcc83 = hmaster1_p & v2303fa7 | !hmaster1_p & !v23f84f9;
assign v23fc7b2 = hready & v22fbf54 | !hready & v2307a75;
assign v150718d = hbusreq3_p & v845636 | !hbusreq3_p & v2301319;
assign v191a8e5 = hbusreq6 & v22f7347 | !hbusreq6 & v23fcfd2;
assign v22f6e67 = hlock3_p & v23f8a41 | !hlock3_p & v230f693;
assign v230e2f9 = hgrant2_p & v23fcf46 | !hgrant2_p & !v22fe9b7;
assign v23fc35a = hbusreq2_p & a1fcc3 | !hbusreq2_p & v84561b;
assign v22fbc63 = hbusreq5_p & v23fa3a4 | !hbusreq5_p & v23f4cd4;
assign v1507071 = hbusreq1_p & v22ed85a | !hbusreq1_p & v23fbdb0;
assign v230ac29 = hbusreq5 & v22f654e | !hbusreq5 & v2300a72;
assign v2391eaa = hgrant5_p & b7029b | !hgrant5_p & v230fa13;
assign v230df81 = hmaster2_p & v23fb99d | !hmaster2_p & v84561b;
assign v23f98d2 = hgrant6_p & v23facb5 | !hgrant6_p & v230d7e2;
assign v23fc0e0 = hbusreq3 & v22f83e8 | !hbusreq3 & v23f4ed3;
assign v23039c0 = hmaster2_p & v84561b | !hmaster2_p & v23fc637;
assign v22f1f92 = hmaster2_p & v2310e40 | !hmaster2_p & v23f11a3;
assign v2302251 = hmaster2_p & v2306d29 | !hmaster2_p & v23fccbe;
assign v23fc5de = hmaster2_p & v845647 | !hmaster2_p & !v84561b;
assign v23efc03 = hbusreq5 & v2306932 | !hbusreq5 & !v23f4722;
assign v191b0e4 = hbusreq0 & v2312f7e | !hbusreq0 & !v231009b;
assign v23fbe95 = hbusreq3_p & v23fb90a | !hbusreq3_p & v23fba9a;
assign v2312e50 = hmaster2_p & v230358b | !hmaster2_p & v22ed85a;
assign v23f8e6b = hgrant1_p & v22ee956 | !hgrant1_p & v230b4d9;
assign v2311e38 = hmaster0_p & v23fc4d1 | !hmaster0_p & v84561b;
assign v23f2d33 = hmaster2_p & v84561b | !hmaster2_p & v22f0945;
assign v23f6326 = hbusreq6 & v22ff18a | !hbusreq6 & v845627;
assign v23fb865 = hmaster2_p & v2301655 | !hmaster2_p & !v23fc530;
assign v2302ea0 = hgrant0_p & v84561b | !hgrant0_p & f40d81;
assign v230f70f = hbusreq3_p & v23fc7b7 | !hbusreq3_p & c173c8;
assign v22ed53e = hmaster1_p & v23f7344 | !hmaster1_p & v84561b;
assign v23fc446 = hmaster1_p & v12cc310 | !hmaster1_p & v23f1cf2;
assign v23fcf82 = hbusreq3_p & v22f61f6 | !hbusreq3_p & v22fa9de;
assign v23fcf14 = hmaster1_p & v22fa3f5 | !hmaster1_p & v84561b;
assign v22eec14 = hbusreq5 & v22f60c6 | !hbusreq5 & !v2391a57;
assign v230ecba = hmaster1_p & v23fc2ab | !hmaster1_p & v230a534;
assign v22ef469 = hgrant0_p & v23fb1c6 | !hgrant0_p & v230aec0;
assign v23fbfbb = hlock3_p & v23fbe24 | !hlock3_p & v23f9395;
assign v8958ff = hmaster0_p & v23fb82a | !hmaster0_p & v23fc20d;
assign v22f77e4 = hbusreq1 & v97b973 | !hbusreq1 & !v845636;
assign v23fb790 = hmaster0_p & v23fc323 | !hmaster0_p & v23fc9dc;
assign v22ee2eb = hmaster1_p & v23f475e | !hmaster1_p & !v230b5c7;
assign v23389c8 = hbusreq1_p & v22f609b | !hbusreq1_p & !v23f0734;
assign v22efc2a = hlock0_p & v230f63f | !hlock0_p & !v22eb1f5;
assign v23fc147 = hmaster2_p & v22ef46e | !hmaster2_p & !v22f8bd0;
assign v2300881 = hbusreq5_p & v22fdabc | !hbusreq5_p & v22f4d68;
assign v22ef772 = hbusreq2 & v22f60c6 | !hbusreq2 & v84564d;
assign v22f2158 = hbusreq3_p & v22fe22a | !hbusreq3_p & v84561b;
assign v23f05c0 = hmaster1_p & v23f38b1 | !hmaster1_p & v23fb3f3;
assign v22fe098 = hmaster0_p & f40ab9 | !hmaster0_p & v230b4c5;
assign v23fce7f = hlock3_p & v22ec96a | !hlock3_p & v84561b;
assign v23fbb50 = hlock3_p & v2306eb5 | !hlock3_p & v84561b;
assign v2311729 = hgrant5_p & v84561b | !hgrant5_p & v23fc2a7;
assign v23fbf90 = jx3_p & v23fce61 | !jx3_p & v23f87e4;
assign v22fab99 = stateG2_p & v84561b | !stateG2_p & !v22f3294;
assign v1b8771f = hbusreq4 & v2307f77 | !hbusreq4 & v84561b;
assign v22f0d07 = hgrant2_p & v23f5af5 | !hgrant2_p & v23fb920;
assign v23f75e5 = hmaster2_p & v22f62ae | !hmaster2_p & v23fcd0a;
assign v22fbdb1 = hmaster1_p & v23058b0 | !hmaster1_p & !v23f84dc;
assign v23fc261 = hbusreq3_p & v23fc664 | !hbusreq3_p & v23f660f;
assign v23f6c8f = hmaster0_p & v23f3d38 | !hmaster0_p & !v23fc485;
assign v22f638b = hbusreq4_p & v23fb94b | !hbusreq4_p & v23fc09c;
assign v23fc15b = hmaster0_p & v23f41ec | !hmaster0_p & !v22ecc5a;
assign v230387b = hgrant4_p & v239298e | !hgrant4_p & v22ff5c1;
assign v2310ab0 = hbusreq6 & v22fb373 | !hbusreq6 & v84561b;
assign v2312be7 = stateG2_p & v84561b | !stateG2_p & !v22f5fa8;
assign v23fc1fb = hlock5_p & e1dcf6 | !hlock5_p & v2392cdd;
assign v23fb0d0 = hmaster2_p & v23f4b28 | !hmaster2_p & v22f0824;
assign v23115ff = hgrant1_p & v106a782 | !hgrant1_p & v23fc7c4;
assign v23fc476 = hbusreq3_p & v2303a62 | !hbusreq3_p & v230e1f2;
assign v23fc772 = hbusreq5_p & v22f037a | !hbusreq5_p & !v23fb4f0;
assign b06cee = hmaster2_p & v84561b | !hmaster2_p & v231228e;
assign v191b186 = hgrant3_p & v23fcf54 | !hgrant3_p & v2307aad;
assign v230cbf6 = hmaster2_p & v23facc2 | !hmaster2_p & !v23fbf32;
assign v23f8edc = hmaster2_p & v22eefd1 | !hmaster2_p & v85d110;
assign v23fba94 = hmaster2_p & v845620 | !hmaster2_p & v23f2be7;
assign v22f6759 = hbusreq3_p & v22f2bab | !hbusreq3_p & v23f6db4;
assign v23fca70 = hgrant1_p & v84561b | !hgrant1_p & v22fe657;
assign v231185e = hmaster1_p & v231242a | !hmaster1_p & v23fc970;
assign v22faf3a = hmaster2_p & v23f9414 | !hmaster2_p & !v23f5f5f;
assign v2303acd = hgrant3_p & v22fd298 | !hgrant3_p & v22ed881;
assign v23fcbba = hbusreq2 & v22ec658 | !hbusreq2 & v84562b;
assign v22fd762 = hgrant5_p & v23fc37d | !hgrant5_p & !v23fc6ed;
assign v23fc6a1 = hbusreq3_p & v2311559 | !hbusreq3_p & v23fcd28;
assign v23fc338 = hgrant0_p & v84561b | !hgrant0_p & v231124e;
assign v23f906a = stateA1_p & v84561b | !stateA1_p & !v23f54be;
assign b10190 = hgrant1_p & v22f3738 | !hgrant1_p & v23f50bb;
assign v23fd011 = hmaster2_p & v23fc23d | !hmaster2_p & v23fbdb0;
assign v22f0ceb = hbusreq6_p & v2312be4 | !hbusreq6_p & v191afde;
assign v23f6283 = hlock3_p & v23f1ad7 | !hlock3_p & v23fc25e;
assign v23f46b3 = hgrant3_p & v2302c68 | !hgrant3_p & v23f54f3;
assign v22ed631 = hbusreq6_p & v22f3eed | !hbusreq6_p & v23fa825;
assign v23fbfcd = hmaster0_p & v23fb1ca | !hmaster0_p & b1e86b;
assign v22fac26 = hbusreq1_p & v23f7ae7 | !hbusreq1_p & v22f64de;
assign v23fc2ab = hbusreq6_p & v22ebe86 | !hbusreq6_p & v84561b;
assign v2306656 = hgrant3_p & v22ecb28 | !hgrant3_p & v23f5e22;
assign v231243e = hmaster2_p & v22f1389 | !hmaster2_p & v2302048;
assign v23f96f7 = hbusreq5 & v23fcb14 | !hbusreq5 & !v23fc839;
assign v22f34c1 = hmaster2_p & v23f1207 | !hmaster2_p & v23fbf24;
assign v23f2553 = hgrant2_p & v23fcd8e | !hgrant2_p & v191a876;
assign v23fcd4f = hmaster2_p & v230a51c | !hmaster2_p & v22f249f;
assign v23fb4c7 = hbusreq1_p & v230da35 | !hbusreq1_p & !v23fbd5c;
assign v230062b = hbusreq3 & v230db5e | !hbusreq3 & v22ef0ab;
assign v23fc331 = stateA1_p & v84561b | !stateA1_p & v22ec1cb;
assign v23fb9ad = hbusreq2_p & v230248b | !hbusreq2_p & !v84561b;
assign v1aad4fb = hlock0_p & v231124e | !hlock0_p & v230207d;
assign v22f9ac5 = hmaster2_p & v23fb1c6 | !hmaster2_p & v22ee956;
assign v23009d5 = hmaster1_p & v2306119 | !hmaster1_p & !v22f7d00;
assign v23fce02 = hmaster0_p & v2303acd | !hmaster0_p & v23f4edc;
assign v22ffcb0 = hlock6_p & v23fc75a | !hlock6_p & !v84561b;
assign v22f42bd = hlock2_p & v230b1ac | !hlock2_p & v845620;
assign v23fbe0e = hmaster2_p & v2391b46 | !hmaster2_p & v23f7ef3;
assign v23fcb61 = hgrant4_p & v84561b | !hgrant4_p & !v22f5c70;
assign v22ec5f2 = hmaster0_p & v84561b | !hmaster0_p & !v23fc5de;
assign v22f2f04 = hbusreq2_p & v17a34e6 | !hbusreq2_p & !v84561b;
assign v23f5767 = jx0_p & v22f5d5e | !jx0_p & v22f7c32;
assign v230aa0d = hgrant5_p & v22f8943 | !hgrant5_p & v22f1037;
assign v22f3272 = hbusreq4 & v23fb58b | !hbusreq4 & v12cc2ff;
assign v23fc57e = hgrant3_p & v22f2e69 | !hgrant3_p & f4066f;
assign v22f1895 = hbusreq1_p & v2308d09 | !hbusreq1_p & !v191a879;
assign v23fccbf = hbusreq3_p & v23f70c6 | !hbusreq3_p & v84561b;
assign v2306873 = hbusreq4 & v22ec191 | !hbusreq4 & v8da3ef;
assign v23102b0 = hlock3_p & v23fbfee | !hlock3_p & v230bead;
assign v23fbac1 = hgrant2_p & v23f5043 | !hgrant2_p & v23f37c6;
assign v2306d9e = hbusreq5 & v22fab80 | !hbusreq5 & !v84561b;
assign v23f4e90 = hmaster1_p & bd0733 | !hmaster1_p & !v230ecb6;
assign v2312b5a = hbusreq3_p & v13aff46 | !hbusreq3_p & v84561b;
assign v22fb773 = hmaster2_p & v22f954f | !hmaster2_p & v230c2b1;
assign v22ff0be = hmaster2_p & v23fcb83 | !hmaster2_p & v2303bc3;
assign v22fb1d6 = hmaster0_p & v23fc351 | !hmaster0_p & v23f710b;
assign v23f7a6d = jx2_p & v23f4a0f | !jx2_p & v230dd4d;
assign v23f50e0 = hbusreq0 & v22f0add | !hbusreq0 & v84561b;
assign v22ed48a = busreq_p & v23f7ffb | !busreq_p & a1fba6;
assign v23fba6b = busreq_p & v191a86f | !busreq_p & !v2309295;
assign v106a782 = hmastlock_p & v845661 | !hmastlock_p & !v84561b;
assign v2312dc1 = hgrant1_p & v84561b | !hgrant1_p & v22fc61a;
assign v23fc1dc = hbusreq0 & v191ae42 | !hbusreq0 & !v84561b;
assign v2392fd0 = hgrant5_p & c25c58 | !hgrant5_p & v23fc9d2;
assign v22fe01a = hmaster0_p & v22f25e6 | !hmaster0_p & v22f56ce;
assign v23f5d5f = hbusreq1_p & v150745f | !hbusreq1_p & v97808c;
assign v23f8bef = hbusreq3 & v932767 | !hbusreq3 & v84561b;
assign v23fc856 = hbusreq1_p & v2307e48 | !hbusreq1_p & v2309891;
assign v230dc43 = hmaster2_p & v22fef4f | !hmaster2_p & !v191a879;
assign v2302f2c = hbusreq5_p & v23fc947 | !hbusreq5_p & v230b0c6;
assign v22f954f = hgrant1_p & v2306d29 | !hgrant1_p & v230bd05;
assign v2305031 = hmaster2_p & v22ffea0 | !hmaster2_p & v84561b;
assign v23fc545 = hbusreq1_p & v22f8629 | !hbusreq1_p & v23f4bbd;
assign v23f3e68 = hbusreq4_p & v2308db0 | !hbusreq4_p & v23fbb53;
assign v23fa21b = hbusreq3_p & v23fbdc1 | !hbusreq3_p & v2313131;
assign v23fbbbe = hbusreq4 & v2306b35 | !hbusreq4 & v84561b;
assign v230fcf6 = hgrant3_p & v23f06ee | !hgrant3_p & v23fc972;
assign v22ec354 = hmaster2_p & v230ca0f | !hmaster2_p & v23fc963;
assign v22f4e2e = hgrant1_p & v84561b | !hgrant1_p & v23058da;
assign v23f1325 = hmaster2_p & v22ffacb | !hmaster2_p & !v84561b;
assign v23fc469 = hlock3_p & v230646f | !hlock3_p & v23059e1;
assign v22f4587 = hbusreq5_p & v23fc89a | !hbusreq5_p & v230da4a;
assign v2303dd7 = hgrant2_p & v22f1681 | !hgrant2_p & v23fc042;
assign v23fc994 = hlock4_p & v230345b | !hlock4_p & v22fd666;
assign v22ed65e = hbusreq5_p & v22fe421 | !hbusreq5_p & v22fc8c8;
assign v23fc76a = hmaster2_p & v84561b | !hmaster2_p & b00ad2;
assign v22f8463 = hmaster2_p & v1e84174 | !hmaster2_p & v22fd0e6;
assign v23fcd84 = hbusreq3_p & v2306fba | !hbusreq3_p & !v2392d61;
assign v2312c3c = hbusreq1_p & v22ee884 | !hbusreq1_p & v22f0945;
assign v12cd540 = jx1_p & v23017a9 | !jx1_p & v23fba66;
assign v23f0d46 = hgrant1_p & v22f6ad2 | !hgrant1_p & v150736d;
assign v22fe4bb = hlock2_p & v106ae1c | !hlock2_p & a1fbb6;
assign v22f893a = hbusreq5_p & v22f19cc | !hbusreq5_p & v84561b;
assign v9bc7cb = hlock0_p & v1506a9e | !hlock0_p & !v84561b;
assign v23f883c = hmaster2_p & v23fcc10 | !hmaster2_p & v2300de3;
assign v2312351 = hgrant5_p & v22f05f3 | !hgrant5_p & v23fc9d2;
assign v2310af0 = hlock0_p & v23fbfd9 | !hlock0_p & v22eb66f;
assign v2393f08 = hbusreq5_p & v22fdabc | !hbusreq5_p & !v84561b;
assign v22fc1df = hgrant1_p & v84561b | !hgrant1_p & v23fb809;
assign v22f4864 = hbusreq1 & v22f6246 | !hbusreq1 & v84561b;
assign v2313134 = hbusreq6_p & v23f9a8e | !hbusreq6_p & v84561b;
assign v23fbbef = hmaster0_p & v23078cb | !hmaster0_p & v22fb74f;
assign v9bcd2e = hmaster0_p & v23fb4ba | !hmaster0_p & v22efa0a;
assign v22fed4e = hburst1_p & v2309a51 | !hburst1_p & !v23fc116;
assign v23fc853 = hlock5_p & v22f4f40 | !hlock5_p & v845620;
assign v22fbf54 = hmastlock_p & v23f984b | !hmastlock_p & v84561b;
assign v230f573 = hgrant5_p & v230bb2a | !hgrant5_p & v2313339;
assign v23020a2 = hbusreq3_p & v23fbf36 | !hbusreq3_p & v22f511c;
assign v22f6372 = stateG10_5_p & v2311891 | !stateG10_5_p & !v22f36ff;
assign v22fffe4 = hmaster2_p & v23fce71 | !hmaster2_p & v2301505;
assign v2309569 = hbusreq3_p & v22f2eba | !hbusreq3_p & v22ee1d1;
assign v22ffc90 = hmaster2_p & v22ec921 | !hmaster2_p & !v2309c28;
assign v22fe19b = hbusreq0 & v23fc514 | !hbusreq0 & !v23022b1;
assign v22ef21f = hlock1_p & v84561b | !hlock1_p & v2304009;
assign v2309499 = hmaster2_p & v845636 | !hmaster2_p & v845626;
assign v22ec08f = hgrant1_p & f406c6 | !hgrant1_p & !v22f4638;
assign v23036a1 = hgrant3_p & v2300de1 | !hgrant3_p & v22fc908;
assign v22efafa = hmaster0_p & v22ebb5c | !hmaster0_p & a1fdb9;
assign v22f18f3 = hmaster2_p & v22f791d | !hmaster2_p & v23fb7d1;
assign v23f6650 = hgrant3_p & v230b38b | !hgrant3_p & v23f0b47;
assign v22f7da7 = hgrant1_p & v23fc4f8 | !hgrant1_p & v22fb5bd;
assign v2301306 = hbusreq4 & v191b186 | !hbusreq4 & v2311dc5;
assign v23fbc42 = hgrant0_p & v106af73 | !hgrant0_p & v23f512e;
assign v22f4a68 = hmaster2_p & v23fc23d | !hmaster2_p & v22ed85a;
assign v23008a1 = hmaster0_p & v23fb4ba | !hmaster0_p & !v22faba5;
assign v2310271 = hgrant1_p & v22eb67a | !hgrant1_p & !v230c2f4;
assign bfde5b = hmaster0_p & v966100 | !hmaster0_p & v2304fdd;
assign v23031eb = hbusreq1 & v23f5218 | !hbusreq1 & v230af81;
assign v23fb9cf = hgrant1_p & v230a9eb | !hgrant1_p & v23f770f;
assign v22f4a4f = hmaster2_p & v22f39e3 | !hmaster2_p & !v22eee34;
assign v9e764b = hbusreq0_p & v2301511 | !hbusreq0_p & v23fa2ec;
assign v22f985c = hlock5_p & v22f0128 | !hlock5_p & v845620;
assign v23f84f8 = hmaster0_p & v23fb910 | !hmaster0_p & v23fbdf5;
assign v22f6d0b = jx1_p & v23055c3 | !jx1_p & v2309410;
assign v22f8f34 = hbusreq6 & v230d2d8 | !hbusreq6 & v84561b;
assign v230a574 = hgrant1_p & v84561b | !hgrant1_p & v23f6e9c;
assign v22fa99c = jx1_p & v23fc3c7 | !jx1_p & v231160c;
assign v22eeea9 = hmaster2_p & v84561b | !hmaster2_p & v23fc120;
assign v22f975b = hmaster2_p & v22fcdf6 | !hmaster2_p & v84561b;
assign v2310d79 = hgrant3_p & v23fbe4f | !hgrant3_p & v23fc881;
assign v23ef93c = hbusreq1 & v2306b2e | !hbusreq1 & !v845622;
assign b16aac = hlock0_p & v84561b | !hlock0_p & !v23084ce;
assign v23fbd41 = hbusreq1 & v230d7b7 | !hbusreq1 & v84561b;
assign v23fc33a = hmaster0_p & v23fc15f | !hmaster0_p & v23f79ba;
assign v22f737d = hmaster0_p & v22f49ff | !hmaster0_p & v230cd34;
assign v22ed6bc = hbusreq0 & v23fb912 | !hbusreq0 & v84561b;
assign v2304ea9 = hbusreq3_p & v8a894a | !hbusreq3_p & v84561b;
assign v1e83fd9 = locked_p & v22ed48a | !locked_p & a1fba6;
assign v230e23c = hbusreq5_p & v23f763f | !hbusreq5_p & v22f4e7f;
assign v23fb856 = hmaster2_p & v23fd050 | !hmaster2_p & v23fb7d1;
assign v23f6079 = hmaster1_p & v23fb64a | !hmaster1_p & !v22f0a39;
assign v23f0e65 = hgrant3_p & v84562e | !hgrant3_p & v22fe775;
assign v230a580 = stateG10_5_p & v23060a6 | !stateG10_5_p & !v84561b;
assign v23fa1cd = hmaster1_p & v1aadb45 | !hmaster1_p & v22f6403;
assign v2393417 = hgrant5_p & v23fc336 | !hgrant5_p & v22ef659;
assign v23fcdd1 = hgrant3_p & v98d402 | !hgrant3_p & v22f659a;
assign v23fa4ca = hbusreq5_p & v191a86f | !hbusreq5_p & !v13afe8f;
assign v23fb456 = hmaster0_p & v23f38d5 | !hmaster0_p & !v84561b;
assign v23013b5 = hbusreq4_p & v23f3bde | !hbusreq4_p & !v23f38f8;
assign v2306cca = hlock6_p & v84561b | !hlock6_p & v22f4ecf;
assign v23f632e = hmaster0_p & v22f31b9 | !hmaster0_p & !v2308d63;
assign v23fcc9e = hbusreq6 & v230b4d4 | !hbusreq6 & !v84561b;
assign v23022b1 = hmastlock_p & v230b364 | !hmastlock_p & v84561b;
assign v22f5e45 = hbusreq1 & v22fcbac | !hbusreq1 & b7b244;
assign v22f64b2 = hgrant1_p & v22f7830 | !hgrant1_p & v230a9d5;
assign v106ae25 = hlock0_p & v22f9ef0 | !hlock0_p & v230d680;
assign v23f6b2f = hbusreq3_p & v23f0ba3 | !hbusreq3_p & v2393742;
assign v23fc587 = hgrant3_p & v23f120d | !hgrant3_p & v2305d89;
assign v230327d = hmaster1_p & v22f397b | !hmaster1_p & v23064bf;
assign v13afb04 = hbusreq4 & bf7e60 | !hbusreq4 & v84562f;
assign v22ed10d = hgrant1_p & v2392836 | !hgrant1_p & v230e4ae;
assign v2302dc1 = jx1_p & v230ad0e | !jx1_p & v23119b0;
assign v22ed674 = hbusreq4_p & v23fcc45 | !hbusreq4_p & v22ee665;
assign v22efb46 = hgrant5_p & v84561b | !hgrant5_p & v22f0ecb;
assign v22fecf3 = hbusreq3_p & a8e3ee | !hbusreq3_p & v230ae3f;
assign v23f2856 = hmaster0_p & v23f439b | !hmaster0_p & v23fc2c1;
assign c086a6 = hlock2_p & v23fce71 | !hlock2_p & v22f1ee5;
assign v23f8a9d = hlock0_p & v230ae24 | !hlock0_p & v845620;
assign v22fcc62 = hbusreq6_p & v17a3514 | !hbusreq6_p & v230b4f9;
assign v2303154 = hbusreq3_p & v22fe852 | !hbusreq3_p & v84561b;
assign v22fabad = hbusreq4_p & v22fdd92 | !hbusreq4_p & v230c0dd;
assign v12cc2ff = hbusreq3_p & v22f28df | !hbusreq3_p & v22fe22b;
assign v2304b8d = hlock3_p & v22f90c3 | !hlock3_p & v2312c3f;
assign v22fc835 = stateG10_5_p & v22f6058 | !stateG10_5_p & a1fba6;
assign v22fb147 = hmaster0_p & v23f2698 | !hmaster0_p & v23f1eb7;
assign v22fb28f = hbusreq3 & v1e84183 | !hbusreq3 & v23fbf55;
assign v23f2e5d = hbusreq3_p & v23fb4e8 | !hbusreq3_p & v23022c3;
assign v2305f67 = jx2_p & v23fc403 | !jx2_p & v2311491;
assign b5b985 = hbusreq3 & v2305194 | !hbusreq3 & v84561b;
assign v23f6658 = hgrant5_p & v84561b | !hgrant5_p & v2312ccb;
assign v22f1d6c = hbusreq6 & v23f26fc | !hbusreq6 & v22ef39f;
assign v230105a = hmastlock_p & v22f2d05 | !hmastlock_p & v84561b;
assign v22f90af = hbusreq6 & v2311ef7 | !hbusreq6 & v23fa9b8;
assign v23111b2 = hbusreq3_p & v2305bf7 | !hbusreq3_p & v23091ef;
assign v230429d = hbusreq3_p & v22f7ad5 | !hbusreq3_p & v84561b;
assign v23fc93e = hgrant2_p & v84562a | !hgrant2_p & v84561b;
assign v23fc197 = hbusreq3_p & v239214a | !hbusreq3_p & v22ee9be;
assign v23f9081 = hmaster2_p & v22fe497 | !hmaster2_p & v23026c8;
assign v191b215 = decide_p & v230b516 | !decide_p & v23fbff5;
assign v22f07cd = hbusreq3_p & v23fba9a | !hbusreq3_p & v22f6949;
assign v23108cb = hbusreq6_p & v23fbda8 | !hbusreq6_p & !v106ae19;
assign v23090fb = hgrant5_p & v2304299 | !hgrant5_p & !v23fb9f8;
assign v23fc2da = hlock4_p & v22fa49d | !hlock4_p & v22eb6e4;
assign v23fb5ee = hgrant3_p & v230b38b | !hgrant3_p & v87c96d;
assign v1aad39a = hbusreq3_p & v23fb5f6 | !hbusreq3_p & v23fbc86;
assign v23efb4d = hmaster2_p & v23fc7ce | !hmaster2_p & !v84561b;
assign v22edeb5 = hbusreq5 & v23f5dab | !hbusreq5 & v23fbade;
assign v23fc136 = hgrant3_p & v84561b | !hgrant3_p & v2305345;
assign v230f331 = hbusreq1_p & v23fbdac | !hbusreq1_p & v2391eaa;
assign v23fbc19 = jx0_p & v23fc9f2 | !jx0_p & bd770f;
assign v15071a6 = hbusreq4 & v2312e50 | !hbusreq4 & v22f0646;
assign v22fa616 = hmaster1_p & v23fcb78 | !hmaster1_p & v230ce9d;
assign v2310558 = stateG10_5_p & v22fb4a1 | !stateG10_5_p & v230aef9;
assign v22ebf32 = hlock4_p & v23f77c5 | !hlock4_p & v23fca5c;
assign v23fc08e = hbusreq4 & v2392f02 | !hbusreq4 & v23fd015;
assign v2391aa0 = hgrant2_p & v84561b | !hgrant2_p & !v23fc556;
assign v23f6afa = hbusreq2_p & v22f037a | !hbusreq2_p & !v23f32eb;
assign v23f606c = hmaster2_p & v2311d0c | !hmaster2_p & !v23f55ea;
assign v23f7094 = hbusreq5 & v23f6e64 | !hbusreq5 & !v84561b;
assign v230ce9d = hmaster0_p & v23f5ac2 | !hmaster0_p & v22f5317;
assign v23fc125 = hlock0_p & v23fcb58 | !hlock0_p & !v230b7c1;
assign v23f5429 = hmaster1_p & v23fc29b | !hmaster1_p & v22f151d;
assign v22f7efd = hgrant5_p & v230b95f | !hgrant5_p & v23fc153;
assign v22fc020 = hbusreq3 & v230c963 | !hbusreq3 & v84561b;
assign v22ff259 = hmaster0_p & v23107f5 | !hmaster0_p & !v2304abd;
assign v22f5e97 = hbusreq3 & v23f9fa4 | !hbusreq3 & v22f5583;
assign v23f7796 = hgrant5_p & v845635 | !hgrant5_p & v22f6090;
assign v239342f = hgrant1_p & v23fca3e | !hgrant1_p & v2392229;
assign v230ce52 = hlock3_p & v22fc88a | !hlock3_p & !v23fc8e4;
assign v23fc1e1 = hbusreq3 & v23f8607 | !hbusreq3 & !v84561b;
assign v230f82b = hbusreq1 & v23f301a | !hbusreq1 & v22fede1;
assign v2300bb2 = hbusreq5_p & v2308356 | !hbusreq5_p & v1aad586;
assign v230aaa7 = hbusreq1_p & v22f1e96 | !hbusreq1_p & !v23125fd;
assign v23fbee9 = hgrant5_p & v23f4cf7 | !hgrant5_p & !v84561b;
assign v23efce3 = hbusreq3_p & v2306728 | !hbusreq3_p & !v84561b;
assign v22f49c4 = hbusreq0 & v2391a57 | !hbusreq0 & !v84561b;
assign v23fa2b8 = hmaster0_p & v23fbdf6 | !hmaster0_p & !v230abb0;
assign v2300cbb = hlock1_p & v23fc1ee | !hlock1_p & v23087f2;
assign v22fc9ad = hbusreq3 & v23fbf58 | !hbusreq3 & v22ff4eb;
assign v23fc17d = hburst1_p & v22f53f3 | !hburst1_p & v84561b;
assign v2304193 = hmaster1_p & v23067cd | !hmaster1_p & !v22ecdc8;
assign v23fbcc2 = hlock6_p & v23fbfcd | !hlock6_p & v1aadc9e;
assign v23036d1 = hmastlock_p & v2300c4a | !hmastlock_p & v84561b;
assign v23f3b1d = hgrant5_p & v2302cce | !hgrant5_p & v84561b;
assign v845643 = hmaster1_p & v84561b | !hmaster1_p & !v84561b;
assign v23fc72c = hmaster0_p & v23fb7b4 | !hmaster0_p & v23fb043;
assign v22f37de = hgrant3_p & v2311748 | !hgrant3_p & v22f4d97;
assign v22fd907 = hmaster2_p & v2311d0c | !hmaster2_p & !v22fae6e;
assign v22f542d = hgrant1_p & v95adb3 | !hgrant1_p & v23fcd38;
assign v2303707 = hgrant5_p & v23fc847 | !hgrant5_p & !v1aad586;
assign v23fc647 = jx3_p & v23f6ec6 | !jx3_p & v22fcf35;
assign v23fc41e = hmaster2_p & v230910b | !hmaster2_p & b60876;
assign v22f7144 = hmaster2_p & v1aad481 | !hmaster2_p & v84561b;
assign v23fc23c = hmaster0_p & v9ce77e | !hmaster0_p & v22f6aa3;
assign v9ad58e = hbusreq3 & v2302e73 | !hbusreq3 & v22f1d96;
assign v22f791d = hbusreq2_p & v230ca2e | !hbusreq2_p & v84561b;
assign v23007a1 = hbusreq5_p & v845636 | !hbusreq5_p & v22ecaef;
assign v23f87ea = hbusreq0 & v22ed6c5 | !hbusreq0 & v84561b;
assign v22f6c3a = hbusreq3_p & v22f2188 | !hbusreq3_p & v230a66b;
assign v22f03c1 = hbusreq6 & b08eee | !hbusreq6 & v84561b;
assign bd74ad = hbusreq1_p & v23112d5 | !hbusreq1_p & v191ad2f;
assign v230bff5 = hbusreq6 & v23fcf88 | !hbusreq6 & v23002bf;
assign v230b740 = hbusreq3 & v2309464 | !hbusreq3 & v22f0e2f;
assign v13affaa = locked_p & v84561b | !locked_p & !v191a876;
assign v23fcf7c = hgrant1_p & v84561b | !hgrant1_p & v23fcbca;
assign f406a3 = hmaster1_p & v230e449 | !hmaster1_p & v23fd00e;
assign v2311ec3 = hbusreq0_p & v23f5cb3 | !hbusreq0_p & !v2310e40;
assign v23fc7cb = hmaster0_p & v22fcc89 | !hmaster0_p & !v23031c5;
assign v2392d8a = hbusreq4_p & v191b160 | !hbusreq4_p & v22f70bd;
assign v22fa2dd = hgrant5_p & v1e84124 | !hgrant5_p & v22fbe99;
assign v2304899 = hbusreq3_p & v22fb3ef | !hbusreq3_p & v84561b;
assign v22ed7b6 = hbusreq3_p & v23131a6 | !hbusreq3_p & v84561b;
assign v22fa4ea = hmaster2_p & v2309c70 | !hmaster2_p & !v23fbb35;
assign v230a7c3 = hbusreq6 & v23fc7c8 | !hbusreq6 & v2392b3d;
assign v2307c44 = hmaster2_p & v230e4ef | !hmaster2_p & v22f1ae5;
assign v2308164 = hmaster0_p & v22f91f1 | !hmaster0_p & v23f6a95;
assign v22ebc9f = hmaster2_p & v231025b | !hmaster2_p & v23fba9a;
assign v23fbe77 = hgrant3_p & v23fa511 | !hgrant3_p & v23fc7d1;
assign v23fb928 = hlock5_p & bbc337 | !hlock5_p & !v22f92b8;
assign v23f73d7 = hgrant5_p & v22ee7e0 | !hgrant5_p & !v22fa16b;
assign v22eb377 = locked_p & v84561b | !locked_p & a1fba6;
assign v230404f = stateG10_5_p & v22f4f1e | !stateG10_5_p & !v84561b;
assign v22fc908 = hmaster2_p & v84561b | !hmaster2_p & v22fa105;
assign v23f6bc1 = hbusreq0_p & v22f8026 | !hbusreq0_p & v84561b;
assign v2310a41 = hbusreq5_p & v22fa594 | !hbusreq5_p & !v13afb01;
assign v2308fe7 = hbusreq0 & v230e71c | !hbusreq0 & v23fa2ec;
assign v22f14bf = hmaster2_p & v22edd3f | !hmaster2_p & v84561b;
assign v22f7ef7 = hmaster2_p & v23fcfa6 | !hmaster2_p & !v845627;
assign v23fc5eb = hbusreq3 & v23fbb64 | !hbusreq3 & v845622;
assign v2305a2a = hmaster2_p & v85d110 | !hmaster2_p & v84561b;
assign v2310f61 = hgrant3_p & v9a4fb4 | !hgrant3_p & v23fc77b;
assign f40ab9 = hgrant3_p & v23fc139 | !hgrant3_p & !v2303154;
assign v23fc6f5 = hgrant6_p & v23fba0d | !hgrant6_p & v23f9945;
assign v230aded = locked_p & v23f5ab1 | !locked_p & a1fba6;
assign v2392d97 = hbusreq1 & v23fcd38 | !hbusreq1 & v84561b;
assign v23f5558 = hgrant6_p & v22f98ca | !hgrant6_p & v22fec16;
assign v23f7b86 = hmaster2_p & v22f8b01 | !hmaster2_p & v23fcd0f;
assign stateG3_1 = !b00b0b;
assign v23fc6ca = hbusreq1_p & v2304184 | !hbusreq1_p & v84561b;
assign v2311b32 = hbusreq4_p & v2393031 | !hbusreq4_p & v191a905;
assign v22eeb19 = hgrant1_p & v230e28d | !hgrant1_p & v230ae06;
assign v191ad8e = hgrant3_p & v23f3e81 | !hgrant3_p & v22f29e5;
assign e1e65a = hgrant3_p & v230fe87 | !hgrant3_p & v23f1c0f;
assign v22f5b4b = hbusreq1_p & v23f63ab | !hbusreq1_p & v1e8413d;
assign v22ee0d6 = hmaster2_p & v22f2db0 | !hmaster2_p & v84561b;
assign ad78c9 = hmaster0_p & v23fc458 | !hmaster0_p & v230ec04;
assign v22eaee7 = hlock3_p & v2311302 | !hlock3_p & v23fb12f;
assign v23f76fb = hgrant3_p & v84561b | !hgrant3_p & !v23fba74;
assign v23089f7 = hmaster2_p & v23fbfd0 | !hmaster2_p & v230984f;
assign v2309889 = hgrant3_p & v22ffa6e | !hgrant3_p & v2305cf5;
assign v22f341f = hmaster2_p & v23fc84b | !hmaster2_p & !v84561b;
assign v2312dfa = hgrant4_p & v2304568 | !hgrant4_p & v23f1133;
assign v22f2319 = hbusreq1_p & v9ec6b5 | !hbusreq1_p & v23fba03;
assign v23f859a = hgrant1_p & v84561b | !hgrant1_p & v1aad571;
assign v22f0f76 = hmaster0_p & v22f6e67 | !hmaster0_p & v23fc038;
assign b8656c = stateA1_p & v22f0362 | !stateA1_p & v22eced4;
assign v22fd032 = hmaster0_p & v15071c7 | !hmaster0_p & !v22f341f;
assign v23f1e80 = hbusreq3 & v230156f | !hbusreq3 & v22f372e;
assign v23f2650 = hbusreq6 & v23fb31d | !hbusreq6 & v84561b;
assign v23f2df7 = hlock6_p & v2302a58 | !hlock6_p & v23fb1c0;
assign v22fb74f = hbusreq6 & v23f35ff | !hbusreq6 & v84561b;
assign v23131af = hmaster2_p & v1507529 | !hmaster2_p & v22f910f;
assign v23f6b18 = hmaster0_p & v22ff1f8 | !hmaster0_p & v22f4642;
assign v23fcb68 = hbusreq3_p & e1cfe5 | !hbusreq3_p & !v84561b;
assign v22f9c34 = hmaster0_p & v191aeb3 | !hmaster0_p & !v2307309;
assign v230272d = hbusreq3_p & v2301f5c | !hbusreq3_p & v23fba9f;
assign v22fc7e6 = hgrant1_p & v84561b | !hgrant1_p & v22f10cc;
assign v23fc834 = hmaster0_p & v23049ad | !hmaster0_p & v22f9b46;
assign v23f0cbe = hbusreq3_p & bd766b | !hbusreq3_p & v22f2b52;
assign v2310476 = hgrant0_p & v22f595f | !hgrant0_p & !v23064ae;
assign v23fc121 = hmaster2_p & v23fbf32 | !hmaster2_p & !v23fbf53;
assign v22fd314 = hmaster2_p & v22ef513 | !hmaster2_p & v22fdc17;
assign v23f7c5a = hmaster1_p & v2311031 | !hmaster1_p & v23067c9;
assign e1e7b0 = hgrant1_p & v84561b | !hgrant1_p & v22ef2c7;
assign v23100c8 = hbusreq1_p & v23f6bc1 | !hbusreq1_p & v23f4b28;
assign v23fc2c6 = hmaster2_p & v2309033 | !hmaster2_p & f40d2d;
assign v1506ec2 = hbusreq4_p & v23fcc45 | !hbusreq4_p & v22ed12a;
assign v23076ca = hmaster1_p & v22f979e | !hmaster1_p & v84561b;
assign v22f03a7 = hbusreq3_p & v2306690 | !hbusreq3_p & v230e19d;
assign v845665 = stateG3_1_p & v84561b | !stateG3_1_p & !v84561b;
assign hgrant4 = !v13afc19;
assign v22fa5a6 = hbusreq4_p & v22ebf32 | !hbusreq4_p & v23f8124;
assign v230ea57 = hmaster2_p & v23fc870 | !hmaster2_p & v22f068b;
assign v230ac33 = hbusreq1 & v845647 | !hbusreq1 & v84561b;
assign v23fbda4 = hgrant1_p & v22ecd97 | !hgrant1_p & v23f00ec;
assign v23fbec3 = hbusreq6_p & v23f55fb | !hbusreq6_p & v2308ddf;
assign v22f867e = hbusreq4_p & v84561b | !hbusreq4_p & v22f20a2;
assign v230e966 = hmaster2_p & v84561b | !hmaster2_p & v22ee9be;
assign v23133fe = hmaster0_p & v23fcdd1 | !hmaster0_p & !v2391a45;
assign v2308e49 = hbusreq6 & v2306540 | !hbusreq6 & v23fcd90;
assign v23f965c = hmaster0_p & v2392254 | !hmaster0_p & v22ed212;
assign v23fbedf = hbusreq1 & v9c12cb | !hbusreq1 & v84561b;
assign v2301044 = hbusreq3_p & v230e473 | !hbusreq3_p & v22fee78;
assign v2393769 = hmaster2_p & v23fc393 | !hmaster2_p & !v2310e40;
assign v22fc05f = hlock0_p & v23f7a5f | !hlock0_p & v22edb0c;
assign v23f2e42 = hgrant1_p & v845626 | !hgrant1_p & v23031b6;
assign v2392ece = hgrant1_p & v23127b3 | !hgrant1_p & !v23fbaf3;
assign v23fcd49 = hmaster2_p & v22eb303 | !hmaster2_p & v230a2c7;
assign v22f909b = hbusreq3 & v22f33e0 | !hbusreq3 & v23fbce6;
assign v2303b2a = hlock6_p & v22f8cee | !hlock6_p & bf9ce3;
assign v22f9023 = hmaster2_p & v23082bc | !hmaster2_p & v23fc921;
assign v230f1c8 = hbusreq3_p & v23fc498 | !hbusreq3_p & !v84561b;
assign v231241e = hbusreq2_p & v23fbae2 | !hbusreq2_p & !v23f1cd5;
assign v2309d0b = hbusreq4_p & v23fc449 | !hbusreq4_p & v84561b;
assign v22f931f = hbusreq0_p & v2303376 | !hbusreq0_p & !v22f36ff;
assign v22f6358 = hgrant1_p & v23fd017 | !hgrant1_p & v23006e9;
assign v22fe2b6 = hmaster0_p & v2311831 | !hmaster0_p & v22ed5c5;
assign v23fc7a4 = stateG10_5_p & v230f222 | !stateG10_5_p & !v10dbf64;
assign v22eb498 = hbusreq3_p & v23fcf38 | !hbusreq3_p & c0e31a;
assign v23fafc5 = hgrant1_p & v84561b | !hgrant1_p & v230a753;
assign v23003a8 = hmastlock_p & v23fb477 | !hmastlock_p & !v84561b;
assign v22ed267 = hgrant5_p & v23fcefd | !hgrant5_p & v23fc1a3;
assign v23f2c8b = hgrant5_p & v2306e27 | !hgrant5_p & !v23022f2;
assign v22f9cb4 = hburst1_p & v84561b | !hburst1_p & v845649;
assign v22f4eab = hbusreq3_p & v23fa5d4 | !hbusreq3_p & v230cfc7;
assign v2311f22 = hlock6_p & v9e23c0 | !hlock6_p & v2309248;
assign v23fcead = hready_p & v23068bf | !hready_p & !v84561b;
assign v22f03a2 = hbusreq3 & v230b4d4 | !hbusreq3 & !v84561b;
assign v22f8309 = hlock3_p & v22f3189 | !hlock3_p & v2309c93;
assign v239315b = hgrant3_p & v84562e | !hgrant3_p & v22ffe8d;
assign v2311be2 = hgrant3_p & v23fc58b | !hgrant3_p & v2311826;
assign v1aadcf6 = hgrant3_p & v84564d | !hgrant3_p & !v23fd008;
assign v23fbc3f = hbusreq5_p & v230aded | !hbusreq5_p & a1fba6;
assign v22f23e7 = hbusreq1_p & v22f7378 | !hbusreq1_p & v231326a;
assign v22f6385 = hgrant5_p & v22f067f | !hgrant5_p & v22f7cab;
assign v23f6890 = hgrant0_p & v230942e | !hgrant0_p & !v22f12cd;
assign v23fbce4 = hbusreq3 & v2300cf1 | !hbusreq3 & v84561b;
assign bf9ce3 = hlock4_p & v22f58a9 | !hlock4_p & !v845632;
assign v23fb145 = hbusreq3_p & v23f15c1 | !hbusreq3_p & v22f5afa;
assign v23f60fb = hmaster2_p & v84561b | !hmaster2_p & !v2304009;
assign v22f5ea8 = hmaster0_p & v84564d | !hmaster0_p & v23fbcad;
assign v22ef4ce = hgrant0_p & v2309b0f | !hgrant0_p & v23fc1c1;
assign v23fbdac = hgrant5_p & v23929a6 | !hgrant5_p & v23f8c71;
assign v23f8ca8 = hgrant3_p & v22fc0ee | !hgrant3_p & v23fb4e8;
assign v23f5cb3 = locked_p & v23fc378 | !locked_p & v191a86f;
assign v23041a6 = hlock6_p & v23fcfe9 | !hlock6_p & !v23f3922;
assign v230f480 = hlock0_p & v2313463 | !hlock0_p & !bd94ed;
assign v23efe7d = hmaster1_p & v22f6053 | !hmaster1_p & v2308bfc;
assign v9a4fb4 = hlock3_p & v23fcfa8 | !hlock3_p & !v23fc0f8;
assign v22f6cec = hbusreq5_p & v23f3a07 | !hbusreq5_p & !v84561b;
assign v230e086 = hbusreq4_p & v23faa94 | !hbusreq4_p & v2306b0a;
assign v23fbe96 = hbusreq1_p & v23f4cb5 | !hbusreq1_p & v845620;
assign v2307ff1 = hbusreq5_p & v2303350 | !hbusreq5_p & !v84561b;
assign v22f8ba5 = hmaster2_p & v23f8364 | !hmaster2_p & v84561b;
assign v1aae374 = hbusreq6_p & v23fbeae | !hbusreq6_p & a89109;
assign v2301ef1 = hbusreq1_p & v2306d29 | !hbusreq1_p & v23065ad;
assign v23f4540 = hbusreq3_p & v22f5edf | !hbusreq3_p & !v84561b;
assign a1ff39 = hgrant5_p & v23fc2a0 | !hgrant5_p & v230474b;
assign v8ce364 = hlock0_p & v2308a42 | !hlock0_p & v23fb25c;
assign v23fcdc1 = hmaster2_p & v22f3aa1 | !hmaster2_p & v23059b0;
assign v23041c3 = hgrant0_p & v22fc11b | !hgrant0_p & v230679a;
assign v22fb17b = hbusreq5 & v2312f7e | !hbusreq5 & v84561b;
assign v230cdf2 = hmaster2_p & fc8c3f | !hmaster2_p & v85f4fd;
assign v230c440 = hmaster0_p & v23f48a1 | !hmaster0_p & v22fb88d;
assign v2301f92 = hgrant0_p & v845622 | !hgrant0_p & v23fc254;
assign v2310895 = hgrant3_p & v84562e | !hgrant3_p & v2312ae4;
assign v230e6ad = stateA1_p & v84561b | !stateA1_p & v22ed56a;
assign v23f3c2a = hbusreq1_p & v1aada71 | !hbusreq1_p & !v23056b1;
assign v22f451b = hmaster0_p & v2312a18 | !hmaster0_p & v22f28eb;
assign v22ee44f = hbusreq1 & v1aae98c | !hbusreq1 & v23fa2ec;
assign v22fc99c = hmaster2_p & bd74c0 | !hmaster2_p & v22f2db0;
assign v23f5787 = stateG10_5_p & v2393775 | !stateG10_5_p & v22f0945;
assign v22f4ecf = hbusreq4_p & v230184a | !hbusreq4_p & !v84561b;
assign v22f484b = hmaster0_p & v23fc804 | !hmaster0_p & v2305483;
assign v22f475e = hmaster2_p & v23fc7c6 | !hmaster2_p & v84561b;
assign v2306538 = hgrant5_p & v84561b | !hgrant5_p & !v2306b33;
assign v22ebe52 = hbusreq6_p & v23fc965 | !hbusreq6_p & v23fbd92;
assign v22fe6b3 = hbusreq5_p & v84561b | !hbusreq5_p & !v23fb8ae;
assign v22f9e3d = hbusreq5_p & v23fccbe | !hbusreq5_p & !v23fc551;
assign v22f9793 = hmaster1_p & v230e7d2 | !hmaster1_p & v1506aab;
assign v22fe627 = hbusreq5 & v22f60c6 | !hbusreq5 & v230d7b7;
assign v22eaea8 = hmaster2_p & v23f62fe | !hmaster2_p & v22f995e;
assign v2309b75 = hbusreq4 & v23fce9d | !hbusreq4 & v22eed0b;
assign v239208c = hbusreq1 & v191ae42 | !hbusreq1 & !v84561b;
assign v230af0f = hmaster0_p & v23f0776 | !hmaster0_p & !v96c563;
assign v22f6e70 = hbusreq5 & v23fa3a4 | !hbusreq5 & v84561b;
assign v23fc56c = hmaster0_p & v23f85a9 | !hmaster0_p & v22f4af1;
assign v13afb6e = hbusreq3 & v1aadad9 | !hbusreq3 & v2310d04;
assign v23fb4a3 = hmaster0_p & v22ef575 | !hmaster0_p & v22f3579;
assign v23f7b9e = hbusreq4_p & v2311027 | !hbusreq4_p & v22eedbb;
assign v22fb727 = hlock0_p & v23fbb84 | !hlock0_p & v23025aa;
assign v23fc07d = hready & v230164e | !hready & v84561b;
assign v2308955 = hmaster2_p & v22f98e3 | !hmaster2_p & !v84561b;
assign v2301f9a = hlock3_p & v23fb84a | !hlock3_p & v23f8345;
assign v230fc1f = hmaster2_p & v23f7ab7 | !hmaster2_p & v2309cdc;
assign v23fcf74 = hbusreq1_p & v230f63f | !hbusreq1_p & !v22eb1f5;
assign v23fca1e = stateG10_5_p & v22ee195 | !stateG10_5_p & v23f972e;
assign b9eb75 = hbusreq5_p & v845636 | !hbusreq5_p & v22f5e36;
assign v23f6adf = hmaster1_p & v23fbf8d | !hmaster1_p & v23fcf60;
assign v23fba0d = jx2_p & v23f6da6 | !jx2_p & v84561b;
assign v22f4ef0 = hbusreq4 & v22f0567 | !hbusreq4 & v2310d04;
assign v22f5768 = jx3_p & v22fb3c8 | !jx3_p & !v22eb14c;
assign v22f8c43 = hgrant1_p & v22fd8e1 | !hgrant1_p & v2300387;
assign v23f486d = hbusreq1 & v2312f7e | !hbusreq1 & !v230e032;
assign v22f6cc8 = hbusreq5_p & v22f56d2 | !hbusreq5_p & v22f9c42;
assign v23f6380 = hgrant0_p & v230a9a0 | !hgrant0_p & !v22f7d41;
assign v23f89b6 = jx1_p & v1507118 | !jx1_p & v84561b;
assign v2301b06 = hmaster1_p & v23fbba6 | !hmaster1_p & v84561b;
assign v23925a8 = hgrant3_p & v230aa99 | !hgrant3_p & v22f0538;
assign v2307eee = hbusreq5 & v1aad481 | !hbusreq5 & v23fc7ef;
assign v23fc946 = hbusreq6_p & v22fa5f1 | !hbusreq6_p & v23fc01f;
assign v23fcac8 = hgrant5_p & v22eea67 | !hgrant5_p & v23fc92a;
assign v23fbeb0 = hbusreq0_p & v23fca4f | !hbusreq0_p & v84561b;
assign v23fc59e = hgrant4_p & v84562d | !hgrant4_p & v2307419;
assign v22f10a7 = hbusreq4_p & v23f420c | !hbusreq4_p & !v23faade;
assign v230f3e5 = hbusreq3_p & v23fbe27 | !hbusreq3_p & v22fa857;
assign v2308a60 = hmaster0_p & v22ee0c0 | !hmaster0_p & v231242a;
assign v23f14ef = hmaster2_p & v23f0169 | !hmaster2_p & v22eefd1;
assign v23fcda1 = hgrant2_p & v2313463 | !hgrant2_p & !v230fec6;
assign v22f3999 = hgrant0_p & v22ec303 | !hgrant0_p & !v23f0ded;
assign v23f57c1 = hmaster2_p & v10dbf64 | !hmaster2_p & !v22fd25c;
assign v2307ec5 = hgrant3_p & v84561b | !hgrant3_p & bd762f;
assign v22fc22b = hgrant3_p & v22fb1bc | !hgrant3_p & v230df44;
assign v2301a7d = hbusreq1 & v23fc514 | !hbusreq1 & !v23022b1;
assign v23f24c5 = hlock5_p & v23f1515 | !hlock5_p & v22f2a76;
assign v12cd993 = stateG2_p & v84561b | !stateG2_p & v2305aa1;
assign v1aadb61 = hmaster2_p & v23055fd | !hmaster2_p & v23fbdc1;
assign v23f5948 = hmaster2_p & v23f660f | !hmaster2_p & v230080a;
assign v22fc90d = hmaster2_p & v23fc93b | !hmaster2_p & !v84561b;
assign v2300791 = hmaster2_p & v23fbb35 | !hmaster2_p & v84561b;
assign b9d038 = hbusreq6 & v23f7158 | !hbusreq6 & v23fc9e4;
assign v23fc8d3 = hgrant5_p & v22f05f3 | !hgrant5_p & !v84561b;
assign v23fba78 = hbusreq3_p & v23fbdbe | !hbusreq3_p & v84564d;
assign v2300e70 = hmaster1_p & v230817b | !hmaster1_p & v23f8d91;
assign v22eb6c8 = jx2_p & v23059c5 | !jx2_p & v22ec763;
assign v23128a1 = hready & v1aae294 | !hready & !v22f3294;
assign v23031f0 = hmaster2_p & v22ffc69 | !hmaster2_p & !v22f7d4e;
assign v230704c = hbusreq1 & v22fc8c8 | !hbusreq1 & v84561b;
assign v230cfba = hbusreq5_p & v22fd8a6 | !hbusreq5_p & v22f4faf;
assign v23fba9f = hbusreq3 & v22ee9be | !hbusreq3 & v230e966;
assign v2306fdd = hmaster2_p & v230708b | !hmaster2_p & v22ecdfe;
assign v23f200b = hlock5_p & v22edfb7 | !hlock5_p & v2309c93;
assign v22f3b33 = hbusreq1 & v13affaa | !hbusreq1 & v84564d;
assign v23f01d2 = hbusreq0 & v23fcc10 | !hbusreq0 & v22ff090;
assign v2308d83 = hmaster0_p & v2304189 | !hmaster0_p & v23fc6a2;
assign v22f37e5 = hbusreq4_p & v2307abc | !hbusreq4_p & v22f02bd;
assign v2300487 = hbusreq3 & v2301216 | !hbusreq3 & v84561b;
assign v22fef4c = jx0_p & bdac8b | !jx0_p & v22fd411;
assign v23022b3 = hbusreq1_p & v230de92 | !hbusreq1_p & v84561b;
assign v23f9c7b = hmaster1_p & v22ebd0b | !hmaster1_p & v2311476;
assign v106a7a1 = hmaster0_p & v23fbf3e | !hmaster0_p & v23fcbe8;
assign v230186e = stateG10_5_p & v22ed49b | !stateG10_5_p & v23fc374;
assign v23042b7 = hmaster2_p & v23fb8be | !hmaster2_p & v2387c09;
assign v23109e5 = hmaster2_p & v22fa70c | !hmaster2_p & aa6574;
assign v2300c5c = hbusreq5_p & v22f56d2 | !hbusreq5_p & v22f42c9;
assign v23fcd66 = hmaster2_p & v106ae4a | !hmaster2_p & a1fbb6;
assign v23fc473 = hbusreq3_p & v230741d | !hbusreq3_p & !v23fb7c3;
assign v23f682c = hmaster0_p & v22ed491 | !hmaster0_p & v22f6aa1;
assign v22eefe2 = hbusreq0 & v23fb567 | !hbusreq0 & v84561b;
assign v22fbde2 = hmaster2_p & v22fe497 | !hmaster2_p & v23fcc9a;
assign v2303d2e = hlock5_p & b9d00f | !hlock5_p & a1fbb6;
assign v230a3b3 = hbusreq6_p & v9ae938 | !hbusreq6_p & v23039fa;
assign v23fcb35 = stateG10_5_p & v84564f | !stateG10_5_p & !v84561b;
assign v23fcd22 = hbusreq5_p & a07f9b | !hbusreq5_p & v22f46a6;
assign v23fc225 = hbusreq5_p & v22faefb | !hbusreq5_p & !v23f0a0b;
assign v230f0c6 = hbusreq4_p & v22f878c | !hbusreq4_p & v22eedbb;
assign v2305799 = stateG10_5_p & v22eb2f1 | !stateG10_5_p & v22fd713;
assign v22f8e4d = hbusreq6 & v2307c0c | !hbusreq6 & v845636;
assign v22f2a1b = hmaster1_p & v22ee60e | !hmaster1_p & v2313504;
assign v23f537e = hbusreq6 & v23fb9fc | !hbusreq6 & !v84562d;
assign v23fc5b0 = stateG10_5_p & v23f6890 | !stateG10_5_p & v22f58f9;
assign v23f790a = hmaster2_p & v23131e8 | !hmaster2_p & !v22fdc17;
assign v23fc0fc = hlock2_p & v84564d | !hlock2_p & v230333f;
assign v23fa590 = hbusreq6_p & v8c495d | !hbusreq6_p & v23fc7e8;
assign v23f2768 = hbusreq1_p & v22ff13f | !hbusreq1_p & v23006e9;
assign v22f5421 = hbusreq1_p & v22ef2c7 | !hbusreq1_p & v23f6658;
assign v2311899 = hgrant5_p & v84561b | !hgrant5_p & v22f2453;
assign v1e84183 = hmaster2_p & v22ed85a | !hmaster2_p & v230358b;
assign v22f6fda = hbusreq6_p & v230089c | !hbusreq6_p & v23fb947;
assign v230928c = hlock1_p & v84561b | !hlock1_p & v23fc658;
assign v23fad33 = hgrant3_p & v22f7dbc | !hgrant3_p & v23fc0ab;
assign v22f8f5c = jx1_p & v22f0074 | !jx1_p & v22f257b;
assign v22f517e = hgrant0_p & v23fc907 | !hgrant0_p & v84561b;
assign e1beab = stateG10_5_p & v2310251 | !stateG10_5_p & v23fb1d1;
assign v22fd827 = hgrant3_p & v23fb17e | !hgrant3_p & !v231262f;
assign v23f6042 = hbusreq6_p & v22ee24a | !hbusreq6_p & v23f723b;
assign v22f68f1 = hmaster2_p & v191a86f | !hmaster2_p & v22fa870;
assign v230813c = hbusreq3_p & v22eea9a | !hbusreq3_p & v2303461;
assign b9ff2b = hmaster2_p & v23fc1ce | !hmaster2_p & v23fba9a;
assign v23fc84b = hbusreq0_p & v23fc2e0 | !hbusreq0_p & !v84561b;
assign v2393775 = hbusreq5 & v230c03a | !hbusreq5 & v84561b;
assign v23f4f9f = hmaster2_p & v2303831 | !hmaster2_p & !v23fb966;
assign v23f4ce2 = hbusreq3 & c043dc | !hbusreq3 & !v845636;
assign v23fcf63 = hmaster2_p & v9526ac | !hmaster2_p & v22ff732;
assign v22fd6c0 = hmaster2_p & v2309c52 | !hmaster2_p & v84561b;
assign v23fba7e = hburst1 & v23fb564 | !hburst1 & v23fa524;
assign v2310fb9 = hmaster0_p & v23f7039 | !hmaster0_p & !v22f1f92;
assign v22f6d06 = hlock0_p & v2303b9a | !hlock0_p & v22ec7a2;
assign v2309a51 = start_p & v84561b | !start_p & v22f476c;
assign v230caac = hbusreq4_p & v2308ced | !hbusreq4_p & v84561b;
assign v22f1a04 = hbusreq1_p & a5a279 | !hbusreq1_p & v23f480d;
assign v22ec763 = hgrant4_p & v230efa0 | !hgrant4_p & v2300070;
assign v22ff79d = hbusreq4_p & v23fb9bf | !hbusreq4_p & v230a87b;
assign v2300c4a = stateG2_p & v2302ca3 | !stateG2_p & !v84561b;
assign v23f37bf = hlock3_p & v22f3091 | !hlock3_p & v84561b;
assign v2305258 = hlock0_p & v23fbfd9 | !hlock0_p & v22fe367;
assign v23fcd96 = hlock5_p & v23fd055 | !hlock5_p & !v84561b;
assign v22f7ad6 = hlock1_p & v23f85d7 | !hlock1_p & !v84561b;
assign v2393f1a = hmaster2_p & v22f2718 | !hmaster2_p & v1aadb8e;
assign v2307b4c = stateG10_5_p & v23fcb53 | !stateG10_5_p & v23fb481;
assign v23fc0c7 = hmaster0_p & v23fbea6 | !hmaster0_p & !v23fa511;
assign v23fc9cf = hbusreq6 & v23fcf96 | !hbusreq6 & v84561b;
assign v12cd570 = hmaster1_p & v2309e42 | !hmaster1_p & v230e97b;
assign v22f0105 = hbusreq5 & v2391a89 | !hbusreq5 & v84561b;
assign v23fb71f = hbusreq2 & v2312f7e | !hbusreq2 & !v22ef3e8;
assign v23fc038 = hbusreq4 & v22ef0c8 | !hbusreq4 & v22fca36;
assign v23f79e9 = hmaster1_p & ad06d5 | !hmaster1_p & v22f448e;
assign v22efa0a = hmaster2_p & v23f6411 | !hmaster2_p & v230a9eb;
assign v22ed48c = hbusreq5_p & v22fd145 | !hbusreq5_p & v84561b;
assign v22efc7f = hbusreq4 & v23925e9 | !hbusreq4 & v84561b;
assign a8ec08 = hmaster0_p & v230f18c | !hmaster0_p & v23fccb5;
assign v2392cdd = hbusreq5 & v22f9911 | !hbusreq5 & !v22ee7a7;
assign v2306e0e = hmaster0_p & v22f81ba | !hmaster0_p & v22f4ef7;
assign v22efcee = hmaster0_p & v23fbea6 | !hmaster0_p & v2304f4c;
assign v22ff45e = hbusreq1 & v23fbb80 | !hbusreq1 & v84561b;
assign v230cfc7 = hmaster2_p & v22f4cf3 | !hmaster2_p & v84561b;
assign v23faa94 = hmaster0_p & v22f9403 | !hmaster0_p & v230801c;
assign v22f51ba = hmaster0_p & v23f9db0 | !hmaster0_p & v22fe4ea;
assign v1e84170 = hbusreq4 & v22ef0de | !hbusreq4 & v230ec4a;
assign v22f743b = hlock3_p & v23f66ec | !hlock3_p & v2305719;
assign v12ce4ac = hmaster2_p & v23fc23d | !hmaster2_p & v230358b;
assign v230984f = hbusreq5_p & v23f8a9d | !hbusreq5_p & v23fb52e;
assign v230d674 = hbusreq4 & v2308955 | !hbusreq4 & v23fc3f2;
assign v23f08af = hbusreq3_p & v22f3c11 | !hbusreq3_p & v23f65c8;
assign v23fc85e = hbusreq3 & v22f60da | !hbusreq3 & !v84561b;
assign v22f2939 = hready_p & v23fc6f5 | !hready_p & v23fbb27;
assign v230b52c = hbusreq5_p & v2391ada | !hbusreq5_p & v2393f52;
assign v230e262 = hbusreq3 & v22ed85a | !hbusreq3 & v84561b;
assign v23fc596 = hlock0_p & v22fdaa5 | !hlock0_p & v845622;
assign v230c4e8 = hgrant3_p & v84562e | !hgrant3_p & v22fdfd9;
assign fc8e3a = hmastlock_p & v22f3294 | !hmastlock_p & v84561b;
assign v23067cd = hbusreq6_p & v23fbd46 | !hbusreq6_p & v23f1824;
assign v230128b = hmaster0_p & v23fbe2d | !hmaster0_p & !v22f438c;
assign v2302992 = hmaster2_p & v23fb793 | !hmaster2_p & v84564d;
assign v22ecaf6 = hlock3_p & v23fcd03 | !hlock3_p & v230abf6;
assign v22f91a8 = hlock3_p & v22ee10b | !hlock3_p & v23fbcc4;
assign v23fc01a = hmaster2_p & v23fbfd0 | !hmaster2_p & v2301505;
assign v23fcc68 = hbusreq4_p & v2308164 | !hbusreq4_p & v23fcb2a;
assign v23fb562 = hlock0_p & v84562b | !hlock0_p & v2302868;
assign v22f3324 = hbusreq5_p & v230c03a | !hbusreq5_p & v23920d8;
assign v2310104 = hbusreq0 & v23fc35a | !hbusreq0 & v2302d97;
assign v2303632 = jx0_p & v22f7d93 | !jx0_p & v2309094;
assign v22ed907 = hgrant3_p & v230eab7 | !hgrant3_p & v15072b7;
assign v23037f2 = hmaster1_p & v23fc0e7 | !hmaster1_p & v2312b57;
assign v23fc8a8 = hbusreq5_p & e1df2d | !hbusreq5_p & v9ee8a4;
assign bd7c3f = hgrant1_p & v23f4426 | !hgrant1_p & v23071f6;
assign v230b504 = hbusreq5 & v230e032 | !hbusreq5 & !v84561b;
assign v2313111 = hmaster0_p & v23fccdb | !hmaster0_p & v2312f81;
assign v23f8a0e = hgrant5_p & v23f087f | !hgrant5_p & v230b59f;
assign v23fcd5c = hgrant3_p & v23f651a | !hgrant3_p & !v84561b;
assign v23f8f21 = hmastlock_p & v22fb157 | !hmastlock_p & v84565f;
assign v2313394 = hbusreq6 & v2304ec9 | !hbusreq6 & !v23f2bfa;
assign v22f902d = hgrant1_p & v23f5af5 | !hgrant1_p & v23089b2;
assign v23fc252 = hbusreq1 & v23105cd | !hbusreq1 & v84561b;
assign v23094f0 = hgrant3_p & v106af01 | !hgrant3_p & v23f5a02;
assign v22eaf83 = hbusreq4_p & v22f8686 | !hbusreq4_p & !v2312ebb;
assign v22f037a = locked_p & v1b87673 | !locked_p & !v84561b;
assign v230b23c = hmaster2_p & v22fe740 | !hmaster2_p & v22f2363;
assign v23f53d0 = hlock3_p & v22f9e59 | !hlock3_p & v2306de4;
assign v23fbf32 = hbusreq1_p & v230aef0 | !hbusreq1_p & v2310c6d;
assign v230fe15 = hbusreq4 & v23fc528 | !hbusreq4 & v23faab2;
assign v23fb109 = hlock0_p & v23f21e5 | !hlock0_p & v23f617e;
assign v23fc8df = hgrant0_p & v9526ac | !hgrant0_p & v230aec0;
assign v12cd534 = hbusreq3_p & v23fba07 | !hbusreq3_p & v23fc957;
assign v23fb8b8 = hlock4_p & v8958ff | !hlock4_p & !v23fc061;
assign v23f960d = hgrant6_p & v23106c2 | !hgrant6_p & v191a965;
assign v2391f3c = hmaster2_p & v23fd060 | !hmaster2_p & v23101b1;
assign v23fbf3e = hmaster2_p & v22ff457 | !hmaster2_p & v23f807d;
assign a7dd55 = hbusreq4 & v23f2843 | !hbusreq4 & v22f4627;
assign v1506ea6 = hlock0_p & v23f1a8d | !hlock0_p & v23062fe;
assign v23fc969 = hbusreq0 & v22ed878 | !hbusreq0 & v230e0d5;
assign v22fc23d = hmaster2_p & v23022b3 | !hmaster2_p & v230dbc9;
assign v23fc79a = hbusreq4_p & v2312164 | !hbusreq4_p & v23f507b;
assign v23f2a5b = hmaster2_p & v23fa463 | !hmaster2_p & !v84561b;
assign v230b9f3 = hmaster1_p & v22f9b3f | !hmaster1_p & v23f04f2;
assign v191b037 = hbusreq6 & v84564d | !hbusreq6 & v22eeece;
assign v22f316f = hgrant0_p & v106a782 | !hgrant0_p & v2306d37;
assign v23fcbf3 = hbusreq3_p & v23fbbb9 | !hbusreq3_p & v23fc750;
assign v230f6e9 = hbusreq6 & v84561b | !hbusreq6 & v23fba11;
assign v23fcab8 = hmaster0_p & b3cfb7 | !hmaster0_p & v22ef270;
assign v230b11a = hbusreq4_p & v23038ea | !hbusreq4_p & v23f810b;
assign v23fcf49 = hlock1_p & v23f8e52 | !hlock1_p & !v84561b;
assign v22ff5bd = hbusreq4 & v1506ff4 | !hbusreq4 & v84561b;
assign v2312885 = hmaster0_p & v23f91d0 | !hmaster0_p & v22f47c6;
assign v23fc742 = hgrant1_p & v22f1cb7 | !hgrant1_p & v22fcf5b;
assign v23f5fcd = stateG10_5_p & v23f1d8b | !stateG10_5_p & v23fcccf;
assign v22f0698 = hbusreq6 & v23fcfb4 | !hbusreq6 & v23fa2ec;
assign v22fbeb3 = hmaster2_p & v230b621 | !hmaster2_p & v22f015d;
assign v22fa65d = hbusreq4_p & v230b5ad | !hbusreq4_p & v2311196;
assign v23fb95a = hmaster0_p & v22f7ad4 | !hmaster0_p & v23f0978;
assign v2302d9a = hgrant1_p & v845629 | !hgrant1_p & v23fb5a2;
assign v23fc053 = jx0_p & v22fb406 | !jx0_p & !v23f623e;
assign v23fb5c4 = hbusreq5_p & v23fb691 | !hbusreq5_p & v22f7004;
assign v230c437 = hgrant3_p & v2312f81 | !hgrant3_p & v22fdc80;
assign v23fb201 = hbusreq6 & v12cd2e3 | !hbusreq6 & !v84561b;
assign v22ec0d1 = hmaster0_p & v22f636a | !hmaster0_p & v23f7429;
assign v230d96b = hbusreq4 & v23fba78 | !hbusreq4 & v84561b;
assign v23fc722 = hmaster2_p & v2307e48 | !hmaster2_p & v84561b;
assign v22ec5e3 = jx2_p & v22f2835 | !jx2_p & v23f1cdf;
assign v23f6db4 = hmaster2_p & v22fef4f | !hmaster2_p & !v191a876;
assign v23fc70c = hbusreq5_p & v22fd8a6 | !hbusreq5_p & v23043af;
assign v22fae48 = hmaster2_p & v2310d04 | !hmaster2_p & v230ef0b;
assign v2306514 = hbusreq1 & v22fcdf6 | !hbusreq1 & v84564d;
assign v2304987 = hgrant3_p & v23f37bf | !hgrant3_p & v22fcabc;
assign v23fc57c = hmaster1_p & v22f5f54 | !hmaster1_p & v22ef9ea;
assign v23f7921 = stateG10_5_p & v23fd049 | !stateG10_5_p & !v84561b;
assign v22fa11e = hmaster0_p & v1b87752 | !hmaster0_p & v230fe15;
assign v23065db = hmaster0_p & v84564d | !hmaster0_p & v2309a10;
assign v23facab = hbusreq3 & da3886 | !hbusreq3 & v84561b;
assign v22f43d7 = hbusreq4_p & v22f8864 | !hbusreq4_p & v23f84f8;
assign v22f220a = hgrant1_p & v23f79b4 | !hgrant1_p & v22f6385;
assign v23f972e = locked_p & v9526ac | !locked_p & a1fbb6;
assign v2311e62 = hbusreq0_p & v23f3a55 | !hbusreq0_p & v23007a2;
assign v23fbc8c = locked_p & v13afbf5 | !locked_p & v84561b;
assign v22f05a9 = hbusreq5 & v2346b8a | !hbusreq5 & v84561b;
assign v23fc083 = hbusreq3 & v22f3d4b | !hbusreq3 & v2312f81;
assign v23f5acd = hbusreq5_p & v23f6a11 | !hbusreq5_p & !v84561b;
assign v2392fa6 = hbusreq4_p & v23fcf9e | !hbusreq4_p & v23fc5c6;
assign v22efdfe = hbusreq3 & v23fbb44 | !hbusreq3 & v84561b;
assign v23fb9a7 = hbusreq3_p & v23fb745 | !hbusreq3_p & v23f5ef2;
assign v22ec5ac = hmaster1_p & v23fc2bc | !hmaster1_p & v84561b;
assign v2308be7 = hbusreq4_p & v230c81f | !hbusreq4_p & v23fbc65;
assign v23fb58b = hbusreq3_p & v22fe0a8 | !hbusreq3_p & v230113d;
assign v23084cf = hbusreq5 & v22ed984 | !hbusreq5 & v84561b;
assign v23027bf = hgrant1_p & v84561b | !hgrant1_p & a1ff39;
assign v230345c = hbusreq1 & v22f98e3 | !hbusreq1 & v23fc3f2;
assign v22fcdf7 = hgrant3_p & v230fd1d | !hgrant3_p & v22f33c4;
assign v23fbe7a = hbusreq5_p & v22fff6e | !hbusreq5_p & !v84561b;
assign stateA1 = !v191b215;
assign v23fca50 = hlock3_p & v22f3cf2 | !hlock3_p & v230e43d;
assign v230fae1 = hmaster2_p & v23f8f25 | !hmaster2_p & v84561b;
assign v22eee15 = hbusreq4_p & v230193c | !hbusreq4_p & v23fc3ca;
assign v22efbe2 = hmaster1_p & v2305847 | !hmaster1_p & v23fbd21;
assign v23f7561 = hmaster2_p & v23fc71b | !hmaster2_p & !v2303b6a;
assign v1e83f8d = hmaster2_p & v106ae4a | !hmaster2_p & v106ae1c;
assign fc8c9b = decide_p & v22f2939 | !decide_p & v22eda04;
assign v22fdba7 = hmaster0_p & v23f90b2 | !hmaster0_p & v23f936e;
assign v23facc2 = hbusreq1_p & v97b973 | !hbusreq1_p & v23fb527;
assign v2310bd4 = hmaster0_p & v22f4d74 | !hmaster0_p & v23f58f9;
assign v22f7c09 = hbusreq5_p & v23fbaa7 | !hbusreq5_p & v22f5109;
assign v12cd66d = hgrant3_p & v23fbe6d | !hgrant3_p & !v84561b;
assign v23f592d = hgrant3_p & v230c20b | !hgrant3_p & v23fcedf;
assign v2300e6b = jx1_p & v22f2a1b | !jx1_p & v23fc786;
assign v2306c80 = hbusreq5 & v23fcf96 | !hbusreq5 & v84561b;
assign v23fc54f = hbusreq3 & v22febaf | !hbusreq3 & v2306e5a;
assign v23f5b39 = hbusreq0_p & v23fbac1 | !hbusreq0_p & v2308848;
assign v23fbfc0 = hbusreq1_p & v2306d29 | !hbusreq1_p & v22fdc30;
assign b9c8dc = hlock2_p & v23fce71 | !hlock2_p & v845620;
assign v23086d9 = hlock6_p & v22f52a0 | !hlock6_p & v23f60ba;
assign v23f196c = jx3_p & v23047dd | !jx3_p & v1aae37a;
assign bd7c53 = stateG10_5_p & v22eb292 | !stateG10_5_p & !v17a34ff;
assign v22f58a9 = hmaster0_p & v23f8d53 | !hmaster0_p & v23fbc53;
assign v23fb999 = hgrant1_p & v22ff732 | !hgrant1_p & v23fb53b;
assign v22febb1 = hmastlock_p & v12cda44 | !hmastlock_p & v84561b;
assign v23f5fdb = hbusreq3 & v23118f7 | !hbusreq3 & !v84561b;
assign v23fbf63 = hbusreq1 & v22fd699 | !hbusreq1 & f40a9e;
assign v2312faa = hmaster0_p & v23fc8ad | !hmaster0_p & !v22fa36f;
assign v2393e5c = start_p & v84561b | !start_p & v1e83f7f;
assign v2304258 = hready_p & v23063fa | !hready_p & v2300f19;
assign v2304990 = hbusreq1_p & v22f8f27 | !hbusreq1_p & v84561b;
assign v23fc443 = hlock2_p & v84561b | !hlock2_p & !v2304ec7;
assign v91ba6f = stateG10_5_p & v22ef9df | !stateG10_5_p & v845636;
assign v23fcfb2 = hbusreq6 & v22f4e48 | !hbusreq6 & v84561b;
assign v2310251 = hgrant0_p & v22ec303 | !hgrant0_p & !v2393364;
assign v22f47c6 = hgrant3_p & v84562e | !hgrant3_p & v2312186;
assign v23fba92 = hgrant3_p & v22f8e29 | !hgrant3_p & v22ec7cf;
assign v22f9f33 = hmaster2_p & v22f0add | !hmaster2_p & v230c876;
assign v2393efc = hmaster1_p & v84561b | !hmaster1_p & !v2305741;
assign v230e040 = hbusreq3 & v2305cf5 | !hbusreq3 & v84561b;
assign v22f92fa = hlock0_p & v845661 | !hlock0_p & !v22f6f8f;
assign v23fcd1b = hgrant2_p & v22f3643 | !hgrant2_p & v22ef751;
assign v23fca2f = hbusreq4 & v22f3550 | !hbusreq4 & v84561b;
assign v23fbb81 = hmaster1_p & v22ec60b | !hmaster1_p & v23f4f2c;
assign v23116b7 = hmaster0_p & v2392f52 | !hmaster0_p & v84561b;
assign v23f9c66 = hgrant4_p & v23f2d6c | !hgrant4_p & v230b18b;
assign v2313370 = hgrant1_p & v12cc2ef | !hgrant1_p & v22f118a;
assign v22fc9cd = hbusreq6_p & v2308d83 | !hbusreq6_p & v23fc0c1;
assign v23fced0 = hbusreq3_p & v23f8345 | !hbusreq3_p & v23f56c3;
assign v23fb14b = hmaster2_p & v23fcd0f | !hmaster2_p & v23fceb6;
assign v22f4ef7 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v230f63f;
assign v22ff0a6 = hbusreq5_p & v22fb2f7 | !hbusreq5_p & v84561b;
assign v22f8e2f = hmaster2_p & v23fc7b2 | !hmaster2_p & v84561b;
assign v22f6a3a = hmaster2_p & v845620 | !hmaster2_p & v2301505;
assign v22fc4d8 = hbusreq2_p & v22f343b | !hbusreq2_p & v84561b;
assign v230d3f5 = hgrant1_p & v84561b | !hgrant1_p & v23fbcbb;
assign v22f4e0b = locked_p & v22f7f52 | !locked_p & !v84561b;
assign v23fb77e = hburst1_p & v84561b | !hburst1_p & v2309a51;
assign v2312025 = hbusreq5_p & v22f8bcf | !hbusreq5_p & v84561b;
assign v23fca5a = hbusreq6_p & v23040c7 | !hbusreq6_p & v230128e;
assign v23fbacb = hbusreq5_p & v23fc8df | !hbusreq5_p & v22ef469;
assign v23f39f2 = hbusreq6 & v23fc7db | !hbusreq6 & v84561b;
assign v2301709 = stateG10_5_p & v22ed49b | !stateG10_5_p & v2310e40;
assign v23032db = hmaster0_p & v191b212 | !hmaster0_p & v86374c;
assign v23fbd28 = hmaster2_p & v84561b | !hmaster2_p & !v1aad847;
assign v23fc77d = hbusreq4 & v22ee499 | !hbusreq4 & v22eb1a8;
assign v2303f04 = hbusreq3_p & v23fc19b | !hbusreq3_p & v91b2de;
assign v22f9b5b = hgrant5_p & v13afaae | !hgrant5_p & v23f5140;
assign v2312dd2 = hmaster2_p & v84561b | !hmaster2_p & v23fc346;
assign v1e83f7f = stateG3_2_p & v22f476c | !stateG3_2_p & v84561b;
assign v230a7a5 = hbusreq3_p & v2303199 | !hbusreq3_p & v2306fdd;
assign v22f6518 = hbusreq0 & v22f15fe | !hbusreq0 & v23f60ef;
assign v2392974 = hbusreq2_p & v12ce195 | !hbusreq2_p & !v23f8914;
assign v23ef4b1 = hmaster2_p & v84561b | !hmaster2_p & v22f69c6;
assign v22f0953 = hmaster2_p & v23fbe60 | !hmaster2_p & v23f660f;
assign v23f89f6 = hgrant1_p & v12cd9f9 | !hgrant1_p & v23fbf46;
assign v22fe144 = hbusreq1_p & v23fb8a8 | !hbusreq1_p & v2311aad;
assign v23fc342 = jx1_p & v23f9c7b | !jx1_p & v84561b;
assign v230bb21 = hbusreq1_p & v22ec1c3 | !hbusreq1_p & v23f8970;
assign v23fcf40 = hbusreq5_p & v23faee6 | !hbusreq5_p & !v84561b;
assign v23efec0 = hbusreq4_p & v22fc67e | !hbusreq4_p & v2391655;
assign v23f6114 = hmaster0_p & v22fa27c | !hmaster0_p & dab2cc;
assign v230de81 = hmaster2_p & v22f0073 | !hmaster2_p & v84561b;
assign v23fce60 = hbusreq6_p & v22ed928 | !hbusreq6_p & v2306b06;
assign v22f125c = hmaster0_p & v22ff1d8 | !hmaster0_p & !v1e84170;
assign v23fc907 = hlock0_p & v2307e48 | !hlock0_p & v2305114;
assign v2311011 = hbusreq4_p & v2392ff9 | !hbusreq4_p & v23fbc61;
assign v23f3501 = hmaster0_p & v23fb8aa | !hmaster0_p & !v230d664;
assign v23fbf84 = hbusreq4_p & v23fbe99 | !hbusreq4_p & v22f65dd;
assign v23f4008 = hmaster2_p & v22f12e5 | !hmaster2_p & v22f8427;
assign v2312236 = hbusreq3_p & v23fc4c3 | !hbusreq3_p & !v106ae19;
assign v2391e5e = hbusreq6 & v845620 | !hbusreq6 & v23fb0bb;
assign fc8f81 = hbusreq3_p & v2307224 | !hbusreq3_p & v22faa4d;
assign v2301972 = jx1_p & v22ec2ba | !jx1_p & v2311c65;
assign v230b0d6 = hbusreq3 & v23fc8d1 | !hbusreq3 & v23f6f99;
assign v2306875 = hmaster2_p & v191b147 | !hmaster2_p & v2313549;
assign v22ecab8 = hmaster2_p & v23115ff | !hmaster2_p & v106a782;
assign v23f741e = hgrant6_p & v22ed53e | !hgrant6_p & v22f3a91;
assign v1aae1de = hbusreq4_p & v22f9a75 | !hbusreq4_p & v2311470;
assign v22faf4e = hmaster2_p & v84561b | !hmaster2_p & v23f32eb;
assign v22f2f3e = hbusreq3_p & v23f476a | !hbusreq3_p & v23fbf37;
assign v231359f = hmaster0_p & v2311a61 | !hmaster0_p & v2305fbf;
assign v23fb938 = hgrant3_p & v23fca7e | !hgrant3_p & v22f6a3a;
assign v23fcdfa = hmaster0_p & v23fceb9 | !hmaster0_p & v2307de6;
assign v2301190 = hbusreq6 & v2308b2f | !hbusreq6 & v84561b;
assign v22fe1c8 = hgrant3_p & v845635 | !hgrant3_p & b7ab40;
assign v2391a45 = hgrant3_p & v23fc20d | !hgrant3_p & v23fb9d0;
assign v2393031 = hmaster0_p & v22f4fb2 | !hmaster0_p & !v96c563;
assign v22fd8a6 = hbusreq5 & v22ed85a | !hbusreq5 & v84561b;
assign v23fc0a6 = hbusreq3_p & v23fbce3 | !hbusreq3_p & v23fba11;
assign v23fcf9c = hbusreq3_p & v22efe1b | !hbusreq3_p & v23fcb6c;
assign v239171e = hlock0_p & v22f03b8 | !hlock0_p & v22f1412;
assign v2311756 = hmaster0_p & v23fb083 | !hmaster0_p & v23f23fb;
assign v13b0013 = hbusreq0_p & v22ee2bb | !hbusreq0_p & v845629;
assign v22f6fba = hmaster1_p & v23f534c | !hmaster1_p & fc8f5a;
assign v22f18b5 = hmaster2_p & v22f902d | !hmaster2_p & !v106ae19;
assign v22fda59 = hgrant1_p & v22f24f8 | !hgrant1_p & !v84561b;
assign v23f282d = hbusreq4_p & v22ee920 | !hbusreq4_p & v23f917f;
assign v23fc786 = hmaster1_p & v22f5cd9 | !hmaster1_p & v23fc39d;
assign v23fc009 = hbusreq6_p & v23fb9c1 | !hbusreq6_p & v230f0de;
assign v2309270 = hmaster2_p & v23f1a8d | !hmaster2_p & v22ee956;
assign v23067c9 = hbusreq6_p & v23fc86a | !hbusreq6_p & !v22fcabb;
assign v23fc6b0 = hlock1_p & v23fc416 | !hlock1_p & !v84561b;
assign v23f1a76 = hready_p & v23fc5c5 | !hready_p & v23fb9aa;
assign v23fc6ed = hbusreq5_p & v23fb1d1 | !hbusreq5_p & v22fcc0d;
assign v13affe0 = hbusreq2_p & v2304415 | !hbusreq2_p & v23f1cd5;
assign v230c213 = jx1_p & v22f3a1f | !jx1_p & v23fba66;
assign v23fce75 = hmaster2_p & v23fb155 | !hmaster2_p & !b9d013;
assign v23fc4fd = hlock0_p & v84561b | !hlock0_p & v231114e;
assign v22fa736 = hmaster2_p & v84561b | !hmaster2_p & !v22f163a;
assign v12cc310 = hbusreq6_p & v23fc270 | !hbusreq6_p & v22f696f;
assign v23fb89c = hgrant3_p & v23f558b | !hgrant3_p & v23f447e;
assign v23f89f0 = jx2_p & v23fb97e | !jx2_p & fc88bb;
assign v22efa49 = hbusreq5_p & v230e07d | !hbusreq5_p & v230a42d;
assign v22eb993 = hgrant4_p & v230e50f | !hgrant4_p & v2304253;
assign v23fbe6e = hmaster0_p & v23fcbfb | !hmaster0_p & v23f56de;
assign v22f129b = hbusreq1_p & v2305a12 | !hbusreq1_p & !v22ec921;
assign v22f86f3 = hbusreq1_p & v22f7aff | !hbusreq1_p & v22f7d5d;
assign v2304fae = hgrant1_p & v22f9df1 | !hgrant1_p & v23f75e9;
assign v22fd196 = hmaster2_p & v22f2a94 | !hmaster2_p & v23129e0;
assign v23fbe6f = hmaster2_p & v23fa63b | !hmaster2_p & !v23fb966;
assign v22f2095 = hmaster2_p & v230665f | !hmaster2_p & v2310bf5;
assign v23f6d75 = jx1_p & v23f3ed0 | !jx1_p & v84561b;
assign v22f8c8d = hmaster0_p & v23fbdf6 | !hmaster0_p & v22f4ef7;
assign v230def2 = hbusreq6 & v23fb5f6 | !hbusreq6 & v23fc46d;
assign v2302cfa = hbusreq3_p & v23f7e51 | !hbusreq3_p & !v84561b;
assign v230716c = hmaster0_p & v230124d | !hmaster0_p & v22f4b44;
assign v23f2e65 = hmaster0_p & v23fcb8d | !hmaster0_p & v84561b;
assign v2301d2f = stateA1_p & v23fb564 | !stateA1_p & v84561b;
assign v23f76f4 = hbusreq3 & v2306405 | !hbusreq3 & !v84562a;
assign v23fcd6a = hmaster2_p & v23fc71d | !hmaster2_p & v230b981;
assign v23fbbc3 = hgrant3_p & v22f4016 | !hgrant3_p & !v23f39fb;
assign v230065b = hgrant3_p & v2309465 | !hgrant3_p & v23fcf65;
assign v23fc6c4 = hgrant1_p & v22f3643 | !hgrant1_p & v23f17e2;
assign v22eb1a8 = hgrant3_p & v84562e | !hgrant3_p & v22f69aa;
assign v23f4426 = hbusreq5_p & v23126ae | !hbusreq5_p & v106af73;
assign v22fd0f1 = hmaster2_p & v230aef0 | !hmaster2_p & !v22eeb07;
assign v2304574 = hbusreq1 & v1e8413d | !hbusreq1 & !v22fbe28;
assign v23082bc = hgrant1_p & v23f8357 | !hgrant1_p & !v191ad4f;
assign v1507102 = hbusreq1_p & v84561b | !hbusreq1_p & v23133a7;
assign v23fc716 = hgrant1_p & v23035ba | !hgrant1_p & v22f9f27;
assign v2303fe4 = hmaster2_p & v84561b | !hmaster2_p & v2300de3;
assign v2311748 = hbusreq3_p & v22f4d97 | !hbusreq3_p & v23f21cf;
assign v22f74f7 = hbusreq5_p & v17a34ff | !hbusreq5_p & v8a0e71;
assign v23f677f = hmaster0_p & v22f38ab | !hmaster0_p & v23fa577;
assign v22f79be = hgrant5_p & v22edb13 | !hgrant5_p & v22fb706;
assign v23fc6ac = hbusreq0 & v22f9911 | !hbusreq0 & v230f5a3;
assign v230f790 = hgrant3_p & v22f2bb8 | !hgrant3_p & v22f2d35;
assign v191aed3 = hmaster2_p & v231026b | !hmaster2_p & v2392c72;
assign v8e4c22 = hbusreq1_p & v2310812 | !hbusreq1_p & v84561b;
assign v23f4be7 = hbusreq6_p & v23fbb77 | !hbusreq6_p & a15268;
assign v23fb8bd = jx3_p & v23f6623 | !jx3_p & v2310291;
assign v22f3b8c = hbusreq6 & v230cbdd | !hbusreq6 & v84561b;
assign v22f9d92 = hmaster2_p & v22f6a6e | !hmaster2_p & v22eb840;
assign v1aae37a = jx1_p & v23013d7 | !jx1_p & v23047dd;
assign v22eef66 = hmaster2_p & v2304b35 | !hmaster2_p & !v23f1a1c;
assign v2306b05 = hgrant5_p & v23f36f1 | !hgrant5_p & !v231055e;
assign v2393742 = hmaster2_p & v22ec745 | !hmaster2_p & !v84561b;
assign v23fc48e = hgrant1_p & v2307ee4 | !hgrant1_p & v22fa682;
assign v879c1f = hbusreq3_p & v23fce10 | !hbusreq3_p & v84561b;
assign v23f98d4 = hbusreq3_p & v2307c44 | !hbusreq3_p & v23fb93f;
assign v230cf1d = hlock6_p & v22f517c | !hlock6_p & v2304b2a;
assign v23106e3 = hmaster2_p & v23101b1 | !hmaster2_p & v22f122e;
assign v23fb9a0 = hgrant5_p & v23fc21b | !hgrant5_p & v23fc2ca;
assign v22fd767 = hgrant0_p & v22eb377 | !hgrant0_p & v22f94a7;
assign v2307a6d = hlock1_p & v2301ad7 | !hlock1_p & !v84561b;
assign v23fbe81 = hbusreq5_p & v230e07d | !hbusreq5_p & v2309aa0;
assign v22f331e = hbusreq1_p & v22f1393 | !hbusreq1_p & v22f5bca;
assign v22f3027 = hlock3_p & v230f4d0 | !hlock3_p & !v230bba4;
assign v23fb567 = hbusreq2 & v23fc7b2 | !hbusreq2 & v22ef8af;
assign v230fb96 = hmaster2_p & v1506fe9 | !hmaster2_p & v22ee956;
assign v2305979 = hgrant0_p & v23fbcb2 | !hgrant0_p & !v2310af0;
assign v23fbeaa = hbusreq0_p & v22ee9be | !hbusreq0_p & v84561b;
assign v22f4a20 = hbusreq3_p & v23fce7b | !hbusreq3_p & v84561b;
assign v22f9f27 = hgrant5_p & v23062f8 | !hgrant5_p & v23fcfcc;
assign v23fb90c = hbusreq0 & v845620 | !hbusreq0 & v22eafea;
assign v23fcdf8 = hmaster1_p & v23fb90b | !hmaster1_p & v84561b;
assign v2310bf7 = stateA1_p & v23fc8a3 | !stateA1_p & !v84561b;
assign v22ff129 = hbusreq3 & v22f1ef1 | !hbusreq3 & v84561b;
assign e1cfe5 = hbusreq3 & v22fda85 | !hbusreq3 & !v84561b;
assign v191ad4f = hgrant5_p & v2309280 | !hgrant5_p & !v22ff0a6;
assign v23fc315 = hbusreq5 & v22eefd1 | !hbusreq5 & v84561b;
assign v22fad24 = hmaster2_p & v23fc40f | !hmaster2_p & v230f010;
assign v23f1879 = hready & v84561b | !hready & v22febb1;
assign v23fbddf = hgrant1_p & v22ff732 | !hgrant1_p & v22ed495;
assign v2310641 = hbusreq3_p & v23fb865 | !hbusreq3_p & v23fb9c6;
assign v23fbf3b = hmaster0_p & v23fc566 | !hmaster0_p & v22f065b;
assign v23f2a15 = hgrant4_p & v845632 | !hgrant4_p & v22fe907;
assign v230acb5 = hbusreq4 & v23fc1fa | !hbusreq4 & v23f3fb6;
assign v22f5de1 = hmaster2_p & v2313463 | !hmaster2_p & !v230fec6;
assign v191ae90 = hbusreq3_p & v23fc1e1 | !hbusreq3_p & !v84561b;
assign v230a05f = hmaster2_p & v23fc957 | !hmaster2_p & v23f717f;
assign v2309c07 = hgrant1_p & v2309c28 | !hgrant1_p & v23fc19a;
assign v23072f3 = hmaster0_p & v84561b | !hmaster0_p & v230330d;
assign v1aada71 = hlock1_p & v22f8271 | !hlock1_p & !v23056b1;
assign v2301edd = hbusreq1 & v231171d | !hbusreq1 & v84561b;
assign v22fa9de = hmaster2_p & v23fbf8b | !hmaster2_p & !v230c727;
assign v191a876 = hmastlock_p & v23fb136 | !hmastlock_p & v84561b;
assign v2300621 = hbusreq5_p & v84561b | !hbusreq5_p & v23f450d;
assign v230ce72 = hmaster0_p & v23fbea6 | !hmaster0_p & v22fcb7b;
assign v2309a8c = hbusreq4_p & v22fcf04 | !hbusreq4_p & v230f0d2;
assign v2307572 = hmaster0_p & v23f90b2 | !hmaster0_p & v22ed7b6;
assign v2303ba8 = hbusreq3 & v23fa903 | !hbusreq3 & v845627;
assign v23fc9fb = hbusreq4 & v22f0b56 | !hbusreq4 & v84561b;
assign v2307d70 = hgrant4_p & v845625 | !hgrant4_p & v23fbb0e;
assign v23fb50c = jx0_p & v22fb214 | !jx0_p & v22f5768;
assign v2308d60 = hbusreq4_p & v22f2592 | !hbusreq4_p & !v230dfa0;
assign v23f22d2 = hbusreq1_p & v22f53d4 | !hbusreq1_p & v845620;
assign v23fbe7c = jx1_p & v23f651e | !jx1_p & v23085b7;
assign v22fa61c = hmaster1_p & v23fc9e8 | !hmaster1_p & v22f836e;
assign v23fcf94 = hbusreq6 & v23f0288 | !hbusreq6 & v22ef062;
assign v2302c28 = hlock0_p & v9526ac | !hlock0_p & v2309598;
assign v23fc900 = hbusreq2 & v22f9911 | !hbusreq2 & !v23f58d2;
assign v22eb99d = hbusreq3_p & v22f8857 | !hbusreq3_p & v23fb099;
assign v22f8686 = hlock4_p & v23f3501 | !hlock4_p & !v230170e;
assign v22ef76f = hbusreq3_p & v22fd79d | !hbusreq3_p & !v84561b;
assign v22ff4eb = hmaster2_p & aca9e4 | !hmaster2_p & !v23f9fc1;
assign v23f5526 = hbusreq5_p & v84561b | !hbusreq5_p & v845623;
assign v22ed55a = hmaster0_p & v2393742 | !hmaster0_p & !v84561b;
assign v23f66a8 = hbusreq1_p & v23fbef9 | !hbusreq1_p & v84561b;
assign v23fc30b = hgrant3_p & v84561b | !hgrant3_p & v23f1703;
assign v23fbc37 = hbusreq4 & v23f2f8d | !hbusreq4 & !v845625;
assign v2308ac3 = jx0_p & v2303253 | !jx0_p & v23fc31c;
assign v22faf49 = hmaster1_p & v94116b | !hmaster1_p & v230e94c;
assign v23fb498 = hbusreq1_p & v2301997 | !hbusreq1_p & v230fc03;
assign v22f6741 = hbusreq2 & v23fc7d5 | !hbusreq2 & v23f391e;
assign v2305eb1 = hmaster0_p & v23f3915 | !hmaster0_p & !v230c83a;
assign v23101dc = hmaster0_p & v23fbcde | !hmaster0_p & v22ff2c4;
assign v23f424b = hmaster2_p & v106a782 | !hmaster2_p & !v22ed000;
assign v2392d6f = hbusreq0_p & v22f1a26 | !hbusreq0_p & !v23fb1a4;
assign c098a9 = jx1_p & v23071be | !jx1_p & v23f83d7;
assign v23070ef = hmaster1_p & v22f9d07 | !hmaster1_p & v22eaf83;
assign v22faa86 = hbusreq4 & v22fbc73 | !hbusreq4 & v23f740f;
assign v1aad38a = hlock0_p & v22f825a | !hlock0_p & v22f1376;
assign v23fcbc3 = hmaster2_p & v23101b1 | !hmaster2_p & be9b63;
assign v22ecdde = hbusreq4 & v23fa903 | !hbusreq4 & !v22f7ef7;
assign v22ed493 = hlock0_p & v23f7789 | !hlock0_p & !v23fcad4;
assign v22edaf2 = locked_p & v230d2a8 | !locked_p & v22f7f74;
assign v22efd4a = hbusreq0 & v22fe421 | !hbusreq0 & v84561b;
assign v22ff33b = hgrant0_p & v845622 | !hgrant0_p & v23fab20;
assign v23fc22d = hlock0_p & v2307836 | !hlock0_p & v23f3d39;
assign v23fb0c2 = hlock5_p & v84561b | !hlock5_p & bbc337;
assign e1e70f = hmaster2_p & v22fc13d | !hmaster2_p & !v84561b;
assign v23fc564 = hgrant2_p & v2310116 | !hgrant2_p & v22f0098;
assign v23f43cf = stateG10_5_p & v2393c3a | !stateG10_5_p & !v21b0f6a;
assign v230b00c = hgrant3_p & v22ffa6e | !hgrant3_p & v2310e05;
assign v22fb4a6 = hbusreq4_p & v23fc32f | !hbusreq4_p & v23f60e8;
assign v23fb919 = hbusreq3_p & v22fb379 | !hbusreq3_p & v2303ba8;
assign v2304a64 = stateG10_5_p & v22f277f | !stateG10_5_p & v22ffbb3;
assign v23fc525 = hgrant3_p & v23fc75d | !hgrant3_p & v23f439a;
assign v23fc570 = stateG10_5_p & v2311089 | !stateG10_5_p & v22f0945;
assign v2306cad = jx2_p & v22fcf35 | !jx2_p & v23fbfa5;
assign v23fb53c = hmaster0_p & v22ecb08 | !hmaster0_p & v239223a;
assign v23fc7db = hmaster2_p & v84561b | !hmaster2_p & v23f3ca5;
assign v23fcc99 = hbusreq3_p & v239213c | !hbusreq3_p & v84561b;
assign v23fc246 = hlock0_p & bda6a0 | !hlock0_p & !v230e40a;
assign v23fbca2 = hmaster0_p & v22f755a | !hmaster0_p & v23fc9cf;
assign v231256b = hgrant3_p & v230d8af | !hgrant3_p & v22f802b;
assign v23fa623 = hbusreq1 & v84564d | !hbusreq1 & v84561b;
assign v23fbde8 = stateG10_5_p & v22f532c | !stateG10_5_p & b9d013;
assign v2312cf9 = hlock3_p & v230ef73 | !hlock3_p & v23025e4;
assign v230ae14 = hlock4_p & v23fb537 | !hlock4_p & v2312ba0;
assign v2312053 = hbusreq3_p & v230118f | !hbusreq3_p & v22f878c;
assign e1e72e = hbusreq6_p & v22ffcbd | !hbusreq6_p & v22f878c;
assign v230941d = hbusreq1_p & v22fd549 | !hbusreq1_p & v84561b;
assign v22eb6ab = hbusreq6 & v23fce9a | !hbusreq6 & !v84561b;
assign v23fb8aa = hbusreq3_p & v23fc3e8 | !hbusreq3_p & v230741d;
assign v230c20b = hlock3_p & v23fc5f8 | !hlock3_p & v22fe831;
assign v22f1498 = hmaster0_p & v2304a2d | !hmaster0_p & !v96c563;
assign v2303388 = hbusreq5_p & v84561b | !hbusreq5_p & v23fc843;
assign v23f649a = hbusreq6_p & v22ff1b9 | !hbusreq6_p & v2309a8c;
assign v23066bf = hlock3_p & v22f1d1a | !hlock3_p & v22ec855;
assign v22eda04 = hgrant6_p & v84561b | !hgrant6_p & v230b2a1;
assign v22f9527 = busreq_p & v2300c4a | !busreq_p & v22ef867;
assign v230bf92 = hgrant2_p & v23fc393 | !hgrant2_p & v22f2903;
assign v230d75a = hbusreq1_p & v84561b | !hbusreq1_p & v23133b3;
assign v23f6130 = hbusreq5_p & v106af73 | !hbusreq5_p & v22fc7c1;
assign v2310eb0 = hgrant3_p & v22f23f6 | !hgrant3_p & v23f2d37;
assign v106ae1c = hmastlock_p & v22ef862 | !hmastlock_p & v84561b;
assign v23fc48b = hbusreq2_p & v22ed85a | !hbusreq2_p & v23fbdb0;
assign v22f878c = hlock0_p & v845622 | !hlock0_p & !v84561b;
assign v230b739 = hmaster2_p & v84561b | !hmaster2_p & !v22fce66;
assign v23f0ded = hlock0_p & v230e606 | !hlock0_p & v2300597;
assign v2393635 = hbusreq6 & v22f19ce | !hbusreq6 & v22f3c27;
assign v13afa38 = hgrant0_p & v23127ef | !hgrant0_p & v22f3502;
assign v22fda35 = hbusreq6_p & v22ff114 | !hbusreq6_p & v22feb04;
assign v22f7e19 = hmaster2_p & v1aae087 | !hmaster2_p & v23fc346;
assign v23fcf60 = hmaster0_p & v230b08d | !hmaster0_p & v22fb802;
assign v23fc0f5 = hmastlock_p & v1e8408b | !hmastlock_p & v84561b;
assign v2310ab6 = hmaster2_p & v84561b | !hmaster2_p & v23fc03f;
assign v2307403 = jx1_p & v230ab7a | !jx1_p & !v23f9812;
assign v23f5276 = hbusreq5_p & v2303e1a | !hbusreq5_p & v22f012b;
assign v230d7e4 = hmaster2_p & v2301319 | !hmaster2_p & v23f5d5f;
assign v23059b0 = hgrant1_p & v22f6b45 | !hgrant1_p & v23fcef5;
assign v2301271 = hmaster2_p & v23fa63b | !hmaster2_p & v22fbeea;
assign v22f48a5 = hbusreq1 & v22f1e02 | !hbusreq1 & !v84561b;
assign v23f58ed = hmaster1_p & v23f99bb | !hmaster1_p & v84561b;
assign v23f3a16 = hlock0_p & v191aa68 | !hlock0_p & v23fb8bf;
assign b8c90d = hbusreq1 & v22fbbb8 | !hbusreq1 & v2311374;
assign v23fb4d8 = hbusreq5 & v13afe3a | !hbusreq5 & !v22fbb8a;
assign v239174b = hmaster0_p & v23fcf35 | !hmaster0_p & v22f160c;
assign v22f15ef = hmaster0_p & v23f38a5 | !hmaster0_p & v22fa371;
assign v22ec414 = hlock6_p & v22fd559 | !hlock6_p & v231253d;
assign v23fbd21 = hmaster0_p & v230aa7a | !hmaster0_p & v230f0de;
assign v22f6870 = hbusreq3 & v23111c0 | !hbusreq3 & v943604;
assign v22ec1b1 = hmaster0_p & v22f2c8a | !hmaster0_p & v23f781b;
assign v23f8093 = hbusreq5 & v1aadb8e | !hbusreq5 & v84561b;
assign v231045a = hbusreq4_p & v23fc267 | !hbusreq4_p & v230ca62;
assign v230c649 = hbusreq5 & v22ecb9d | !hbusreq5 & v84561b;
assign v230080a = hgrant1_p & v12cc2ef | !hgrant1_p & v230b9ad;
assign v22fd048 = hgrant3_p & v22f52a4 | !hgrant3_p & v22f9faa;
assign v22f5272 = hmaster0_p & v230f133 | !hmaster0_p & !v23045dc;
assign v12cd552 = hmaster0_p & v23fc68e | !hmaster0_p & v22ebb8e;
assign v22f3c9a = hbusreq5_p & v23fa720 | !hbusreq5_p & !v84561b;
assign v2307805 = hbusreq2 & v2310ad7 | !hbusreq2 & !v23fc669;
assign v230bf69 = stateA1_p & v84561b | !stateA1_p & !v23fb564;
assign v2302c4b = stateG2_p & v84561b | !stateG2_p & v22f3294;
assign v230074c = hmaster2_p & v23101b1 | !hmaster2_p & v22faa40;
assign v2301cee = hmaster2_p & v23fba9a | !hmaster2_p & v22fe346;
assign v22efbd5 = hbusreq3_p & v230b08b | !hbusreq3_p & v2308b02;
assign v2304913 = hmaster0_p & v23fc1ab | !hmaster0_p & v22eb359;
assign v23006c2 = jx2_p & v23fc403 | !jx2_p & v23fc8d9;
assign v22ec66d = hmaster2_p & v23fcfb8 | !hmaster2_p & v22fb77d;
assign v2309c2c = hgrant5_p & v12ce9b8 | !hgrant5_p & v12cd9c9;
assign v2301bdf = hbusreq3_p & v22fc4a3 | !hbusreq3_p & v22fc6e6;
assign v23fcffd = hbusreq6_p & v23fbd62 | !hbusreq6_p & v23f9a4d;
assign v2311a27 = hmaster2_p & v22fc80c | !hmaster2_p & v230e3a0;
assign v2310d74 = hlock2_p & ac37a1 | !hlock2_p & !v84561b;
assign bd76c5 = hready_p & v23063db | !hready_p & v22f006c;
assign v22f836e = hbusreq4_p & v2303a32 | !hbusreq4_p & v23f6a5b;
assign e1dcf4 = hbusreq5 & v230415a | !hbusreq5 & v230979f;
assign v2302c45 = hbusreq4_p & v23f7564 | !hbusreq4_p & v230560c;
assign v22eec02 = hbusreq5 & v2392ea0 | !hbusreq5 & v23f2ecd;
assign v85f4fd = hgrant1_p & v231128c | !hgrant1_p & v23fc9ef;
assign v23f999c = hbusreq0_p & v84561b | !hbusreq0_p & v23f8747;
assign v23fc68e = hbusreq4 & v22f961e | !hbusreq4 & v22f2ca2;
assign v22fd7ea = hgrant5_p & v23f9a06 | !hgrant5_p & v230a9f0;
assign v230bd8f = hmaster2_p & v23f5d5f | !hmaster2_p & v2301319;
assign v22fe2dc = hmaster2_p & v230bdd0 | !hmaster2_p & v23fa4bd;
assign v22f1244 = hgrant1_p & v84561b | !hgrant1_p & v22eeb7d;
assign v23100e9 = hmaster0_p & v22f82cd | !hmaster0_p & !v22feac9;
assign v23fba08 = hgrant0_p & v845620 | !hgrant0_p & v23fca7d;
assign v238b0d7 = hgrant0_p & v230fec6 | !hgrant0_p & !v23fcda1;
assign v23fcfd9 = hbusreq6 & v1aada96 | !hbusreq6 & v84561b;
assign v86e576 = hgrant3_p & v230d8af | !hgrant3_p & v23fcb6f;
assign v23fcaf8 = hmaster1_p & v84561b | !hmaster1_p & v230381a;
assign c24c97 = hgrant3_p & v22f3027 | !hgrant3_p & v22f6721;
assign v23fabb8 = hbusreq6 & v23f6acc | !hbusreq6 & !v23f06d7;
assign v230031f = hbusreq5_p & v23fb825 | !hbusreq5_p & v845620;
assign bcc479 = hbusreq4_p & v22ff66a | !hbusreq4_p & v23f8d5a;
assign v23f23bf = hmaster1_p & v23fa590 | !hmaster1_p & v22fa8e8;
assign v2309094 = jx1_p & v23f645e | !jx1_p & v22fdb25;
assign v22eec47 = hmaster2_p & v10dbf64 | !hmaster2_p & !v191a879;
assign v2307c17 = jx1_p & v239223a | !jx1_p & v23f6396;
assign bd74b6 = hbusreq6_p & v22ed291 | !hbusreq6_p & v22fb0ac;
assign v23f761c = hbusreq1_p & v23f619e | !hbusreq1_p & !v84561b;
assign v23131eb = hmaster1_p & v23fc9c2 | !hmaster1_p & v23fcffd;
assign v22f9f2f = hbusreq6_p & a9176f | !hbusreq6_p & v22f771b;
assign d49f20 = hbusreq2 & v22f2718 | !hbusreq2 & v84561b;
assign v106af01 = hmaster2_p & v22ebb79 | !hmaster2_p & v2303b6a;
assign v23fa882 = hmaster2_p & v22ede4d | !hmaster2_p & v84561b;
assign v23fc577 = stateG10_5_p & v84564f | !stateG10_5_p & v84561b;
assign v22fe723 = hbusreq6_p & v22ece0e | !hbusreq6_p & v23fc687;
assign v23065d6 = hgrant4_p & v23fb5c0 | !hgrant4_p & v2302d68;
assign v23fc821 = hmaster2_p & b9d0d2 | !hmaster2_p & !v2307852;
assign v23fc9c2 = hbusreq6_p & v23fc940 | !hbusreq6_p & v23fbe94;
assign v23919f9 = hgrant1_p & v23f4b28 | !hgrant1_p & v2391eaa;
assign v22f2db6 = hbusreq3_p & v23fc139 | !hbusreq3_p & !v84561b;
assign v230a3af = hgrant5_p & v230b23b | !hgrant5_p & v230bc8b;
assign v106af57 = hgrant0_p & v23f5af5 | !hgrant0_p & v22f0d07;
assign v2311e03 = hmaster2_p & v84561b | !hmaster2_p & v2307e48;
assign v2310197 = hbusreq4 & v23fc846 | !hbusreq4 & v84561b;
assign v22ef481 = jx1_p & v23fa966 | !jx1_p & v23fcc97;
assign v231246b = hmaster1_p & v23fcf4c | !hmaster1_p & !v23f49cd;
assign v230158e = hgrant2_p & v22fa195 | !hgrant2_p & !v84561b;
assign v2300290 = hlock0_p & v22ee0c4 | !hlock0_p & v23fc47e;
assign v22ef3e8 = hlock2_p & v230e032 | !hlock2_p & v23fbbd2;
assign v231051e = hmaster2_p & v23fa875 | !hmaster2_p & v22f4114;
assign v22f96e9 = hlock0_p & v2311a1d | !hlock0_p & v23fb576;
assign v22f2aa4 = hbusreq0 & v22feb47 | !hbusreq0 & v84561b;
assign v22fc569 = hlock2_p & v230882d | !hlock2_p & v84561b;
assign v2300387 = hgrant5_p & v2368b8a | !hgrant5_p & !v22f3999;
assign v2392077 = hbusreq1 & v23f5a2e | !hbusreq1 & v23fc614;
assign v22f0678 = hgrant1_p & v12cc2ef | !hgrant1_p & v22f6187;
assign v23fcee9 = hgrant0_p & v84561b | !hgrant0_p & v22fca2f;
assign v22fc9cb = hbusreq3_p & v22f8e08 | !hbusreq3_p & v23fbfba;
assign v23107f0 = hlock3_p & v23f2578 | !hlock3_p & v23fcd66;
assign v22f8ed1 = hmaster2_p & v1aad481 | !hmaster2_p & v1aad38a;
assign v22ff066 = hgrant0_p & v23fce0d | !hgrant0_p & v84561b;
assign v23130a1 = hgrant1_p & v230fc8c | !hgrant1_p & !v23f7795;
assign v22fbf19 = jx0_p & v23fc3b9 | !jx0_p & v2313637;
assign v23f50f8 = hmaster0_p & v23101f4 | !hmaster0_p & v23fb727;
assign v23f9424 = hmaster2_p & v22fa70c | !hmaster2_p & !v1507134;
assign v23fb4b1 = stateG10_5_p & v22f8107 | !stateG10_5_p & v22f9de9;
assign v230af11 = hmaster0_p & v23fbdf6 | !hmaster0_p & v23045dc;
assign v230b5ad = hmaster0_p & v23087bc | !hmaster0_p & !v23fbdc2;
assign v2310385 = hbusreq4 & v23f7503 | !hbusreq4 & v84561b;
assign v23f82bb = hmaster2_p & v2301fc9 | !hmaster2_p & !v23f87f4;
assign v22f4f42 = hlock0_p & b9d00f | !hlock0_p & v238ae11;
assign v2312edb = hbusreq6_p & v2307abc | !hbusreq6_p & v22f37e5;
assign v23fc637 = hgrant1_p & v84561b | !hgrant1_p & v22f6607;
assign v2308ef6 = jx1_p & v23f651e | !jx1_p & v23fc32e;
assign v23fca45 = jx1_p & v230cc12 | !jx1_p & v230f151;
assign v23f58e1 = hgrant3_p & v231196d | !hgrant3_p & v22f36da;
assign v23fc673 = hmaster0_p & v230ada5 | !hmaster0_p & v22f8f34;
assign v23f4af5 = hbusreq5_p & v22fb706 | !hbusreq5_p & v23fbc42;
assign v23fbaf3 = hgrant5_p & v23efc12 | !hgrant5_p & !v230eb18;
assign v2310b47 = hmaster0_p & v230cc18 | !hmaster0_p & v23f7659;
assign v22f6ac8 = hgrant5_p & v22f8b0a | !hgrant5_p & v23fa3a4;
assign v22fcea7 = hbusreq3_p & v23074c9 | !hbusreq3_p & v23f8976;
assign v22fb157 = stateA1_p & v84561b | !stateA1_p & !v23fba7e;
assign v2312e02 = hbusreq1_p & v230de18 | !hbusreq1_p & !v2300934;
assign v23fc97a = hlock4_p & v23fc7d6 | !hlock4_p & !v84561b;
assign v22ff404 = stateG10_5_p & v1aad586 | !stateG10_5_p & v23fcc36;
assign v23f8c71 = hgrant0_p & v84561b | !hgrant0_p & v22f1a1b;
assign v23f38a5 = hgrant3_p & v230199e | !hgrant3_p & v23fb200;
assign v22f8626 = hmaster2_p & v2312f7e | !hmaster2_p & v2392974;
assign v23fbb5a = hmaster2_p & v23fbbf2 | !hmaster2_p & !v84561b;
assign v23fbbf2 = hlock0_p & v23f69ba | !hlock0_p & v845622;
assign v22f3ca0 = hbusreq5_p & b5f51c | !hbusreq5_p & e1e73a;
assign v2391935 = decide_p & v230884d | !decide_p & v2304258;
assign v230a51c = hgrant1_p & v23fd033 | !hgrant1_p & v23f6865;
assign v230997b = hbusreq1_p & v2306514 | !hbusreq1_p & v23f8a06;
assign v23fc430 = hlock3_p & v23107cf | !hlock3_p & !v230627c;
assign v23933e8 = hgrant1_p & v845626 | !hgrant1_p & v23fc799;
assign v23fbd38 = hbusreq3_p & v23fbcad | !hbusreq3_p & v84561b;
assign v2311568 = hgrant3_p & v84561b | !hgrant3_p & v22f33e0;
assign v23fceb0 = hbusreq5_p & v23fc4a1 | !hbusreq5_p & v22f5515;
assign v22f07d5 = hmaster2_p & v22f8427 | !hmaster2_p & v22f389b;
assign v22ede8c = hbusreq6 & v22f7758 | !hbusreq6 & v84561b;
assign v23fbdfc = hgrant3_p & v22ec0d9 | !hgrant3_p & v23fc709;
assign v23f4cdc = hlock0_p & v22f9d69 | !hlock0_p & !v23fbe7e;
assign v23f1f1e = hbusreq5 & v23f5be9 | !hbusreq5 & v23f54ef;
assign v2392066 = hbusreq3_p & v22f20df | !hbusreq3_p & !v84561b;
assign v23fbc28 = hmaster1_p & v22eb657 | !hmaster1_p & v84561b;
assign v1aad421 = hlock3_p & v23fbd7e | !hlock3_p & !v92eb35;
assign v230c805 = hbusreq5_p & v2311a1d | !hbusreq5_p & v22f96e9;
assign v22f25c6 = hbusreq2_p & v23fbafd | !hbusreq2_p & v84561b;
assign addc42 = hgrant5_p & v23fcfdf | !hgrant5_p & !v84561b;
assign v23f3bd2 = hmaster0_p & v13afb18 | !hmaster0_p & v23fd037;
assign v2305a1c = hbusreq5 & v23fc1a3 | !hbusreq5 & v84561b;
assign v230fc70 = hbusreq0 & a476c2 | !hbusreq0 & !v84561b;
assign v1e8408c = hbusreq4_p & v230f257 | !hbusreq4_p & v2305eb1;
assign v22ee9ac = hbusreq5 & v23fbbd2 | !hbusreq5 & !v84561b;
assign v23037b2 = hlock5_p & v23fc7e9 | !hlock5_p & !v84561b;
assign v230c70b = hbusreq1_p & v230ea6d | !hbusreq1_p & !v230aef0;
assign v23fc19a = hgrant5_p & v23fcb1f | !hgrant5_p & bd7786;
assign v22eb49d = hbusreq3_p & v23fcb6f | !hbusreq3_p & v23f2504;
assign v23f3e42 = hbusreq3_p & v22f8093 | !hbusreq3_p & v230b19a;
assign v22fe920 = hgrant1_p & v23fb6ff | !hgrant1_p & !v84561b;
assign v22ee62f = hbusreq3_p & v22f128d | !hbusreq3_p & !v23087e8;
assign v23006f8 = hgrant3_p & v23fc460 | !hgrant3_p & v23fb8ec;
assign v23fba39 = hbusreq3_p & v2306f2e | !hbusreq3_p & v23fba73;
assign v22fc997 = hbusreq0 & v22fe165 | !hbusreq0 & v84562a;
assign v230c616 = hmaster0_p & v23fb923 | !hmaster0_p & v22f7cbf;
assign v22ff29c = hmaster0_p & v2303bee | !hmaster0_p & !v23f8a70;
assign v230d90f = hmaster2_p & v22f3643 | !hmaster2_p & v22fef02;
assign v23fbbe7 = hgrant1_p & v22f7830 | !hgrant1_p & v191ab30;
assign v23938ff = hbusreq1 & v230910b | !hbusreq1 & v230b981;
assign bd9e8b = hbusreq1 & v22f0945 | !hbusreq1 & v23f9789;
assign v23f8a49 = hmaster0_p & v22f56a5 | !hmaster0_p & v22faa26;
assign v23fbdc1 = hgrant1_p & v84561b | !hgrant1_p & !v23fc8d3;
assign v22f1000 = hgrant2_p & v23fbbf6 | !hgrant2_p & !v230fec6;
assign v2392d9f = hgrant1_p & v22f129b | !hgrant1_p & v23fcd30;
assign v17a34f8 = hbusreq2_p & v22ef0fe | !hbusreq2_p & v22ee59c;
assign v22f5d84 = hmaster2_p & v22fef4f | !hmaster2_p & !v22f9980;
assign v23054d5 = hmaster0_p & v230b7fc | !hmaster0_p & v23099fc;
assign v191a973 = hgrant0_p & v1e83fd9 | !hgrant0_p & v23f8395;
assign v23139c3 = hbusreq3_p & v230e2bb | !hbusreq3_p & v23f924a;
assign hgrant0 = !bd785e;
assign v23006a1 = hmaster0_p & v23fc23e | !hmaster0_p & !v8d1fa5;
assign v230b161 = hlock0_p & v22ed6bc | !hlock0_p & a51d7a;
assign v230bed2 = hbusreq2 & v23105cd | !hbusreq2 & v84561b;
assign v23fcd73 = hbusreq2 & v22f0785 | !hbusreq2 & v84561b;
assign v23fbc6d = hbusreq3 & v84564d | !hbusreq3 & aca9e4;
assign v230fb9e = hlock1_p & v22ee281 | !hlock1_p & !v84561b;
assign v23faacf = stateA1_p & v84561b | !stateA1_p & !v2305e86;
assign v230522c = hgrant5_p & v230173a | !hgrant5_p & v2312336;
assign v22fb5bd = hgrant5_p & v22f22b2 | !hgrant5_p & v22f7004;
assign v230824c = hmaster0_p & v23fbe74 | !hmaster0_p & v2312007;
assign v2306e1a = hbusreq5_p & v22f3643 | !hbusreq5_p & v22fd2f5;
assign v23f134a = hgrant5_p & v84561b | !hgrant5_p & v23f4e99;
assign v22f0128 = hbusreq5 & v23fbfd0 | !hbusreq5 & b9d02f;
assign e1d3f0 = jx1_p & v23fbabc | !jx1_p & v2304193;
assign v230da3e = hgrant3_p & v22f2123 | !hgrant3_p & v22fb27b;
assign v22f580d = hbusreq3_p & v23fc19b | !hbusreq3_p & v2303c9d;
assign v23f302c = hbusreq6 & v2302992 | !hbusreq6 & v191ae4a;
assign v23fbd19 = hmaster2_p & v22f8271 | !hmaster2_p & v22f3a35;
assign v23113e8 = hbusreq1_p & v23fc561 | !hbusreq1_p & v23fc1fe;
assign v230a0d1 = hbusreq3_p & ba1576 | !hbusreq3_p & !v23f57c1;
assign v23f3ac9 = hbusreq3 & v23fccd8 | !hbusreq3 & !v845636;
assign v22f0295 = hbusreq1_p & v22fd7ea | !hbusreq1_p & v22fa682;
assign v23009cc = hgrant2_p & v84561b | !hgrant2_p & v9526ac;
assign v23fbae0 = hmaster0_p & v84564d | !hmaster0_p & v23fcfab;
assign v22fbb07 = hbusreq1 & v22f893a | !hbusreq1 & v23f87f4;
assign v230e8a8 = hmaster2_p & v23080ec | !hmaster2_p & v23fceb6;
assign v230c117 = hbusreq6 & v1b87672 | !hbusreq6 & v84561b;
assign v23fbe66 = hmaster2_p & v22fb8d6 | !hmaster2_p & !v84561b;
assign v23fc747 = hmaster1_p & v23f07c2 | !hmaster1_p & v23fcd6e;
assign v23127ff = hgrant1_p & v845626 | !hgrant1_p & v23fcfbc;
assign v22ee394 = hbusreq4 & v22f6844 | !hbusreq4 & v23f87f4;
assign v2300b6b = hlock1_p & v23fcb0a | !hlock1_p & v845620;
assign v23fcba6 = hmaster1_p & v22edf7b | !hmaster1_p & !v2313134;
assign bd9dce = hbusreq3_p & v2309c93 | !hbusreq3_p & v22f878c;
assign v9d8aae = busreq_p & v23f273d | !busreq_p & v23fc63e;
assign v23f41c2 = hmaster2_p & v84561b | !hmaster2_p & !v1507102;
assign v22f5d89 = hbusreq6_p & v22f21d0 | !hbusreq6_p & v22fea77;
assign v230c899 = hmastlock_p & v15071da | !hmastlock_p & v84561b;
assign v22f4a1f = hbusreq3_p & v23f35ea | !hbusreq3_p & v22f61b6;
assign v92eb35 = hbusreq3_p & v1aad4c6 | !hbusreq3_p & v23fc92f;
assign v2308b24 = hbusreq4_p & v84562b | !hbusreq4_p & v922c74;
assign v2302244 = hmaster0_p & v23f58e1 | !hmaster0_p & v22eedcd;
assign v23f7992 = hburst0_p & v22f4e3c | !hburst0_p & v23119e0;
assign v22fb511 = hbusreq3_p & v23135ca | !hbusreq3_p & v84561b;
assign v22ec502 = hmaster0_p & v15071c7 | !hmaster0_p & v23135f8;
assign v23fcbed = hbusreq3 & v230d291 | !hbusreq3 & v22f3f32;
assign v23f7af2 = hbusreq6 & v22f95c1 | !hbusreq6 & v84564d;
assign v23fbe1d = hmaster2_p & v23f4da0 | !hmaster2_p & v230b0f5;
assign v22ff4bc = hbusreq4_p & v23fbcd2 | !hbusreq4_p & v23051a9;
assign v1aad988 = hmaster2_p & v84562a | !hmaster2_p & !v84561b;
assign v2308c3d = hbusreq3 & b06cee | !hbusreq3 & !v84561b;
assign v23f9ae7 = hbusreq3_p & v23f1432 | !hbusreq3_p & v22f9db5;
assign stateG10_4 = !v1128cd1;
assign v22f8d8e = hbusreq1 & v22ee9be | !hbusreq1 & v84561b;
assign v23f32a6 = hbusreq1 & v23f3d14 | !hbusreq1 & v22ee9be;
assign v919ce6 = hready & v230bf6d | !hready & !v84561b;
assign v231124e = hgrant2_p & v84561b | !hgrant2_p & !v2305fe0;
assign v23fc002 = hmaster2_p & v230efeb | !hmaster2_p & v2305c24;
assign v230ad15 = hbusreq6 & v23fc27d | !hbusreq6 & v84561b;
assign v22fd3c7 = hgrant4_p & v2303650 | !hgrant4_p & v23fbe36;
assign v230fc03 = hbusreq1 & v22f343b | !hbusreq1 & !v84562a;
assign v23fc8f6 = hlock3_p & v22f9dfb | !hlock3_p & !v84561b;
assign v2308a91 = hgrant3_p & v2312f81 | !hgrant3_p & v191a912;
assign v22f2879 = hbusreq0 & v2301b2d | !hbusreq0 & v2312637;
assign v23fce1b = hlock6_p & v22fd364 | !hlock6_p & !v23f6c83;
assign v22fd387 = hbusreq0 & v13afe3a | !hbusreq0 & !v22f9a51;
assign v869055 = hlock2_p & v84561b | !hlock2_p & v84564d;
assign v23fd03b = hgrant0_p & v23f5af5 | !hgrant0_p & v230b91d;
assign v23fc20d = hmaster2_p & v2306d29 | !hmaster2_p & v230f63f;
assign v23fcccf = hgrant0_p & v22f66bc | !hgrant0_p & v2303d1d;
assign v23fbab4 = hmaster2_p & v22fc8c8 | !hmaster2_p & v23f6b67;
assign v2391f85 = hbusreq1_p & v230a2bb | !hbusreq1_p & v22eeb7d;
assign v230ed77 = hbusreq4_p & v23f9fc8 | !hbusreq4_p & v2312d33;
assign v22fb3c1 = hbusreq5 & v23f3115 | !hbusreq5 & v23f40ba;
assign v230192f = hbusreq5_p & v845636 | !hbusreq5_p & v22ed6ac;
assign v1aad69f = hbusreq6 & v23f1263 | !hbusreq6 & v22fd1ba;
assign v23108bb = hmaster1_p & v23fc946 | !hmaster1_p & v230ecb6;
assign v23010ae = hmaster0_p & v2309c45 | !hmaster0_p & v84561b;
assign v22f8acc = hmaster1_p & v23fc065 | !hmaster1_p & v22f1efd;
assign v191aa98 = jx0_p & v2303a2d | !jx0_p & v22feb39;
assign v2391fc6 = hmaster0_p & v2300d5f | !hmaster0_p & v230e857;
assign v22ef3d4 = hbusreq5_p & v23fcf91 | !hbusreq5_p & v230254a;
assign v22f324f = hmaster2_p & v23fb5a1 | !hmaster2_p & v23f0329;
assign v22f2884 = hbusreq0 & v2313118 | !hbusreq0 & v23f1879;
assign v22f368e = hmaster2_p & v22f3ed0 | !hmaster2_p & v23f98ab;
assign v23fbf10 = hbusreq1_p & v2303558 | !hbusreq1_p & !v22fae6e;
assign v23007de = hbusreq4_p & v2302e0f | !hbusreq4_p & v22f65dd;
assign v22ede66 = hmaster1_p & v22f831d | !hmaster1_p & v23f49cd;
assign v230bdd6 = hmaster2_p & v22ffc55 | !hmaster2_p & v22f2f44;
assign v22efd39 = hlock6_p & v22fff51 | !hlock6_p & v84561b;
assign v23fba4f = hbusreq2_p & v22ecee2 | !hbusreq2_p & !v84561b;
assign v23031bc = hbusreq6_p & v84561b | !hbusreq6_p & v23fc42c;
assign v22ef725 = hgrant0_p & v23f87b7 | !hgrant0_p & v230faaf;
assign v23fc51e = hgrant3_p & v22efb8e | !hgrant3_p & d79b38;
assign v23fb619 = hlock5_p & v22f9cd7 | !hlock5_p & v230d379;
assign v922c74 = hmaster0_p & v230e43d | !hmaster0_p & v22eb338;
assign v23fc061 = hmaster0_p & v2304a06 | !hmaster0_p & v23fc92f;
assign v22eb970 = hmaster0_p & v84564d | !hmaster0_p & v230bb9f;
assign v2309317 = hmaster0_p & v22ff6c5 | !hmaster0_p & !v2300f82;
assign v22f39e3 = hgrant1_p & v23120a5 | !hgrant1_p & !v23fb8da;
assign v23f598e = hgrant3_p & v84561b | !hgrant3_p & !v22eb8ae;
assign v230d7b7 = locked_p & v2307a75 | !locked_p & !v84561b;
assign v22fdb5c = hmaster2_p & v23f87f4 | !hmaster2_p & !v23fcf77;
assign v2301bcb = hlock3_p & v2310253 | !hlock3_p & v230105d;
assign v230e8d0 = hgrant0_p & v2313463 | !hgrant0_p & !v23f0162;
assign v22fc32c = hmaster2_p & v2310e81 | !hmaster2_p & v22f954f;
assign v2300a72 = hbusreq0 & v230d630 | !hbusreq0 & !v84561b;
assign v22f511c = hmaster2_p & v22f878c | !hmaster2_p & !v84561b;
assign v2307c0c = hmaster2_p & v230aef0 | !hmaster2_p & !v23f63ab;
assign a88394 = hgrant1_p & v22f56d2 | !hgrant1_p & a5a279;
assign v1506fdd = jx2_p & v230183d | !jx2_p & v935301;
assign v22f3586 = hmaster0_p & v23f9e9f | !hmaster0_p & v2310f61;
assign v2391665 = hgrant3_p & v23f651a | !hgrant3_p & v23fc6bd;
assign v22eeb4b = hbusreq4_p & v23fbcc3 | !hbusreq4_p & v84561b;
assign v2311629 = hmaster2_p & v8d360e | !hmaster2_p & v84561b;
assign v2312e04 = hbusreq3_p & v230c15a | !hbusreq3_p & !v84561b;
assign v2392fbd = hbusreq5_p & v23f908f | !hbusreq5_p & !v23f47d5;
assign v23f1e5c = hmaster0_p & v22f789c | !hmaster0_p & v2302251;
assign v23fcea3 = hmaster2_p & v84561b | !hmaster2_p & v23088b3;
assign v22f3b24 = hmaster2_p & v1e84174 | !hmaster2_p & v22ee8f3;
assign v23fc71d = hlock5_p & v230ec10 | !hlock5_p & !v845636;
assign v22ee681 = hmaster0_p & v23fbdf6 | !hmaster0_p & !v23f5066;
assign b8a8d7 = hbusreq1_p & v12cd3bc | !hbusreq1_p & v23fb966;
assign v2305a26 = hbusreq3_p & v23f6588 | !hbusreq3_p & v9c8a7f;
assign v22ff80d = hmaster0_p & v23f96b0 | !hmaster0_p & v22ef079;
assign v23fcbd8 = hlock4_p & v22f0c6d | !hlock4_p & v230713e;
assign v23f44d0 = hmaster2_p & v23fcdb4 | !hmaster2_p & v22ef062;
assign v22eeff5 = hbusreq3_p & v22ff538 | !hbusreq3_p & v22f61b6;
assign v230f857 = hmaster0_p & v2393909 | !hmaster0_p & v230a510;
assign v23f420e = hbusreq5 & v23fba6b | !hbusreq5 & v84561b;
assign v22f52c1 = hlock2_p & b09503 | !hlock2_p & v84561b;
assign v23fce6f = hmaster1_p & a1fd78 | !hmaster1_p & !v2311eb3;
assign v23fbb25 = hmaster1_p & v22fe723 | !hmaster1_p & v23fbe4b;
assign v23f2d31 = hmaster2_p & v22fef4f | !hmaster2_p & !v22f4986;
assign v22fb379 = hbusreq3 & v22ec2c4 | !hbusreq3 & v22ef062;
assign v9bf2ce = stateG10_5_p & v13afa38 | !stateG10_5_p & !v23fba6b;
assign v22f6c36 = hlock5_p & v23fb218 | !hlock5_p & v23fbe12;
assign v23fbb1c = hgrant2_p & v23fb3cf | !hgrant2_p & !v84561b;
assign v23f420c = hlock4_p & bd8ac4 | !hlock4_p & !v23faade;
assign v23fba34 = hmaster2_p & v23fcdbe | !hmaster2_p & v2313370;
assign v845620 = hready & v84561b | !hready & !v84561b;
assign v22f6534 = hgrant4_p & v84561b | !hgrant4_p & v23fccfd;
assign v22efe6e = hgrant3_p & v23fb0d0 | !hgrant3_p & v22f263c;
assign v23fc628 = jx1_p & v22f25ed | !jx1_p & !v23f89f4;
assign v23fc621 = hmaster0_p & v2301f63 | !hmaster0_p & v23110f1;
assign v23fb883 = hgrant1_p & v84561b | !hgrant1_p & v23fcb44;
assign v23fc2dc = hbusreq3_p & v23fcf63 | !hbusreq3_p & v22eb563;
assign v23fcbdc = hgrant3_p & v84562e | !hgrant3_p & v22ebc9f;
assign v23f3b00 = stateG10_5_p & v2393f52 | !stateG10_5_p & v23fbd03;
assign v22f8483 = hbusreq3_p & v22f2bab | !hbusreq3_p & v91b2de;
assign v2312e39 = hmaster0_p & v22ebe46 | !hmaster0_p & v23fb4e5;
assign v23046d0 = hbusreq1_p & v22f561a | !hbusreq1_p & v23fc6b1;
assign v1aae5da = hmaster1_p & v23fbfa0 | !hmaster1_p & v23f4961;
assign v23f2be7 = hbusreq2_p & v845620 | !hbusreq2_p & v22f79fd;
assign v22fdaa0 = hgrant2_p & v23fc6f3 | !hgrant2_p & !v12cd3f4;
assign v23fce22 = hgrant2_p & v22fbadb | !hgrant2_p & fc8ab7;
assign v2302ba4 = jx2_p & v23fbaf6 | !jx2_p & v22ff3c6;
assign v23fbf9c = hgrant5_p & v23fcec2 | !hgrant5_p & !v22fa16b;
assign v23fcb1b = hmaster0_p & v22ede34 | !hmaster0_p & v23fc6cc;
assign v23f85b6 = hbusreq3_p & v23040c8 | !hbusreq3_p & v84561b;
assign v22f9f01 = hbusreq6_p & v22ff09a | !hbusreq6_p & v2304e51;
assign v22ed07d = hbusreq3_p & v23fa4cb | !hbusreq3_p & v2304faf;
assign v230a4b6 = hbusreq1_p & v23f87f4 | !hbusreq1_p & v22fb1bc;
assign ba4552 = hbusreq3_p & v2392f11 | !hbusreq3_p & v230a226;
assign v22ff257 = hmaster2_p & v2310d04 | !hmaster2_p & !v23fc71b;
assign v23fc2ea = stateG10_5_p & v84561b | !stateG10_5_p & !v2305fe0;
assign v23fc2d8 = jx0_p & v22fa299 | !jx0_p & v22fabaf;
assign v23fcb5a = hbusreq3_p & v22ff129 | !hbusreq3_p & v84561b;
assign v239407e = hmaster0_p & v231024c | !hmaster0_p & v22efa8c;
assign v22f802b = hmaster2_p & v23101b1 | !hmaster2_p & v22ebb7b;
assign v943604 = hmaster2_p & v84561b | !hmaster2_p & !v22fede1;
assign v23f1133 = hmaster1_p & v23fcbbb | !hmaster1_p & v2305263;
assign v23fc0f3 = hlock5_p & v22f3a35 | !hlock5_p & !v106ae19;
assign v22ec334 = hlock1_p & v23f40d1 | !hlock1_p & v22f60c6;
assign v22f09c4 = hbusreq4 & v845620 | !hbusreq4 & v23fba11;
assign v22f5696 = hbusreq2_p & v2392803 | !hbusreq2_p & !v84561b;
assign v22f28df = hmaster2_p & v22f1ece | !hmaster2_p & !a39dae;
assign v230f4a8 = hbusreq0 & v22fc8c8 | !hbusreq0 & v84561b;
assign v230c2b1 = hgrant1_p & v23070c1 | !hgrant1_p & v23fcb9a;
assign v22f45e9 = hlock3_p & v23fce49 | !hlock3_p & !v84561b;
assign v230d836 = hgrant3_p & v84561b | !hgrant3_p & v22eeea9;
assign v230fd86 = hbusreq6_p & v22ffa1b | !hbusreq6_p & v23f9283;
assign v23fb217 = hbusreq5_p & v23fc853 | !hbusreq5_p & v230c5ad;
assign v23fcd88 = hbusreq2 & v2312bd0 | !hbusreq2 & v84561b;
assign v22f16ef = hmaster2_p & v23f91a5 | !hmaster2_p & v84561b;
assign v23f3768 = hmaster1_p & v22f1f55 | !hmaster1_p & !v23f49cd;
assign v22fdb01 = hgrant5_p & v22ee269 | !hgrant5_p & v22f9de9;
assign v230a83f = hmaster2_p & v230f5a3 | !hmaster2_p & v84564d;
assign v87eb7a = hbusreq4_p & v23fc87a | !hbusreq4_p & v22f7997;
assign v22ef607 = hmaster0_p & v2302da4 | !hmaster0_p & v23fb9a3;
assign v23113d2 = hbusreq3_p & v2311675 | !hbusreq3_p & v12cda0a;
assign v23139aa = hlock0_p & v84561b | !hlock0_p & v23f4ab8;
assign v22fff51 = hmaster0_p & v84561b | !hmaster0_p & v22eedac;
assign v23023c9 = hgrant2_p & v22f3643 | !hgrant2_p & !v84561b;
assign v22f154e = hmaster2_p & v84561b | !hmaster2_p & v22feb20;
assign v2300071 = hbusreq5_p & v22fd8a6 | !hbusreq5_p & v84561b;
assign v23fc521 = hbusreq4 & v23fcec1 | !hbusreq4 & !v84562d;
assign v230088c = hlock2_p & v84564d | !hlock2_p & !v84564d;
assign v23f90c4 = hbusreq5 & v23fb9c2 | !hbusreq5 & v84564d;
assign v23fb584 = hbusreq1 & v23fa997 | !hbusreq1 & b30f07;
assign v23075ba = hgrant3_p & v84561b | !hgrant3_p & v15072a9;
assign v23fb7b4 = hbusreq4 & v23f0288 | !hbusreq4 & v22ef062;
assign v22f9089 = hgrant1_p & v230bbb3 | !hgrant1_p & v2312351;
assign v22ebc3c = hbusreq5_p & v2311810 | !hbusreq5_p & v22f04a6;
assign v230c233 = hbusreq1_p & v23f8a0e | !hbusreq1_p & v230ae1e;
assign v23fb4af = hmaster0_p & v23fc585 | !hmaster0_p & v23fb96b;
assign v22f59e9 = hlock0_p & v23f9545 | !hlock0_p & !v84561b;
assign v23fcb90 = hbusreq4_p & v23fb635 | !hbusreq4_p & !v84563a;
assign v22fae6e = hbusreq5_p & v23046f7 | !hbusreq5_p & v22fd25c;
assign v13afc17 = hbusreq1_p & v23fbd9b | !hbusreq1_p & v84561b;
assign v22f1c57 = hbusreq1_p & v23f6d39 | !hbusreq1_p & a1fba6;
assign v23fbc94 = hlock1_p & v22eb2a2 | !hlock1_p & !v84561b;
assign v22f118a = hbusreq1_p & v22f28d6 | !hbusreq1_p & bab0c9;
assign v230ea9f = hbusreq3_p & v23f73ba | !hbusreq3_p & v2310d04;
assign v22f5f1c = hbusreq1 & v23fb8c1 | !hbusreq1 & v84561b;
assign v22efa3b = hbusreq2 & v22f4e0b | !hbusreq2 & v230f5a3;
assign v22f898b = hbusreq5 & v13affaa | !hbusreq5 & v84564d;
assign v12cd54c = hbusreq1 & v23131e8 | !hbusreq1 & !v84561b;
assign v2312b99 = hbusreq6 & v230eca1 | !hbusreq6 & v23f87f4;
assign v22fadf8 = hbusreq3_p & v22f595b | !hbusreq3_p & v22f0953;
assign v23f3f46 = hlock5_p & v845661 | !hlock5_p & !v84561b;
assign v23fb4d4 = hbusreq0_p & v2303d8f | !hbusreq0_p & v845620;
assign v23052a2 = jx0_p & v23fce12 | !jx0_p & v23fb8bd;
assign v2301d4e = hbusreq4_p & v12cda51 | !hbusreq4_p & v22ee36d;
assign v23fb9b7 = hbusreq1_p & v23fcbe3 | !hbusreq1_p & v22f7241;
assign v23f9e9f = hgrant3_p & v22f4809 | !hgrant3_p & v230ae4f;
assign v22fe428 = hlock1_p & v23f1d35 | !hlock1_p & !v845622;
assign v23919ec = stateG10_5_p & v23fba08 | !stateG10_5_p & v845620;
assign v22f4d69 = hbusreq5 & v2307150 | !hbusreq5 & v84564d;
assign v22fc80c = hgrant1_p & v23fbb8d | !hgrant1_p & v230a25a;
assign v22fa711 = hbusreq5_p & v23f40ba | !hbusreq5_p & v22f442c;
assign v191ac63 = jx2_p & v2303554 | !jx2_p & v22f8639;
assign v23fb5a7 = hbusreq6 & v23045f5 | !hbusreq6 & v84561b;
assign v22eb74d = hmaster2_p & v12cc2ef | !hmaster2_p & !v230aeb3;
assign v22ec6e7 = hgrant0_p & v22ffb9d | !hgrant0_p & !v2300c97;
assign a878fd = hmaster0_p & v23f0aec | !hmaster0_p & v22ef3d1;
assign v239162d = hmaster1_p & v22fb011 | !hmaster1_p & v2300c23;
assign v23fc921 = hgrant1_p & v23fbf2c | !hgrant1_p & !v191aada;
assign v23f9d9a = hgrant3_p & v98d402 | !hgrant3_p & v22fa73a;
assign v23089b2 = hgrant5_p & v23f4c32 | !hgrant5_p & v23fd03b;
assign v23fb482 = hbusreq6_p & v22f037f | !hbusreq6_p & v84561b;
assign v23f61f7 = stateG2_p & v84561b | !stateG2_p & bd3bb2;
assign v23fb7c3 = hmaster2_p & v22fccf1 | !hmaster2_p & v2309475;
assign v2310a05 = hmaster2_p & v2309b7e | !hmaster2_p & !v23fa345;
assign v23fb8e3 = hbusreq5_p & v23f4a00 | !hbusreq5_p & v23f5787;
assign v22f4cca = stateG2_p & v84561b | !stateG2_p & v22f4e3c;
assign v23fcbaf = hmaster0_p & v23fb82a | !hmaster0_p & v2300362;
assign v23fb476 = stateG2_p & v84561b | !stateG2_p & v230e6ad;
assign v22f216d = hmaster0_p & v23fcfd2 | !hmaster0_p & v22f7347;
assign v22f931d = hlock0_p & v22f5037 | !hlock0_p & v23fa8aa;
assign v2310934 = hbusreq4_p & v22f3879 | !hbusreq4_p & v23f8692;
assign v230d3c2 = hmaster2_p & v84561b | !hmaster2_p & v2301e25;
assign v23009f0 = locked_p & v23f68bf | !locked_p & v84561b;
assign v23fb925 = hbusreq3 & v22f9f88 | !hbusreq3 & v22eeece;
assign v23f0588 = hmaster2_p & v23f972e | !hmaster2_p & v22ee956;
assign v23fd06a = hgrant0_p & v23fb97f | !hgrant0_p & v2308e98;
assign v2302fbf = hbusreq6_p & v230d02b | !hbusreq6_p & v23fbf28;
assign v230d282 = hmaster1_p & v22f25c5 | !hmaster1_p & v2307480;
assign v22fe81e = hgrant3_p & v230f70f | !hgrant3_p & v23fc7b7;
assign v2309ca8 = hbusreq3_p & v22fd0f1 | !hbusreq3_p & v23fc121;
assign v23fce3b = hbusreq1_p & v22f037a | !hbusreq1_p & !v23f32eb;
assign v23fce4c = hgrant1_p & v23f794b | !hgrant1_p & v22ec1c3;
assign v23fc9b9 = hgrant0_p & v84564d | !hgrant0_p & !v84561b;
assign v22eeb7a = hgrant3_p & v98d402 | !hgrant3_p & v23fcf82;
assign v22fc8fb = hgrant3_p & v1aae206 | !hgrant3_p & v1aad31f;
assign v23fa893 = hmaster0_p & v84561b | !hmaster0_p & v22f7e09;
assign v22ee0db = hgrant1_p & v22f5e59 | !hgrant1_p & v938878;
assign v23fcc3c = hbusreq5_p & v22f76c2 | !hbusreq5_p & !v84561b;
assign v23fbe4f = hmaster2_p & v22f2ed7 | !hmaster2_p & v22fbeb1;
assign v230f863 = hmaster2_p & v13afe8f | !hmaster2_p & !v191ae42;
assign v23fc90b = hmaster1_p & v22f3730 | !hmaster1_p & v106a7d3;
assign v23fb8a7 = hbusreq5 & v23fc2a7 | !hbusreq5 & v230979f;
assign v22ee9d2 = jx1_p & v85e5cf | !jx1_p & v23057f1;
assign a1fbc2 = locked_p & v84561b | !locked_p & a1fbb6;
assign v22ee26d = stateG10_5_p & v23041c3 | !stateG10_5_p & v2310da2;
assign v23f75aa = hbusreq0 & v2302e32 | !hbusreq0 & v84561b;
assign v22efe01 = hmaster0_p & v23fb526 | !hmaster0_p & v22f6d45;
assign v23fcb01 = jx3_p & v22ef3fe | !jx3_p & v230cc70;
assign v23f77b1 = hbusreq3_p & v23f5cfe | !hbusreq3_p & bd7adc;
assign v23fc5ce = hmaster1_p & v230997a | !hmaster1_p & !v23fbba0;
assign v230b3d2 = jx1_p & v23fcc1c | !jx1_p & aacd54;
assign v2310aee = hgrant3_p & v23082fe | !hgrant3_p & v2305d92;
assign v23fcd7f = hmaster2_p & v23f445f | !hmaster2_p & v2310e10;
assign v2304339 = hbusreq5_p & v22fea89 | !hbusreq5_p & v22ff33b;
assign v230b38b = hmaster2_p & a1fbc2 | !hmaster2_p & v22ee956;
assign v23fc268 = hgrant3_p & v22ed1b5 | !hgrant3_p & v23fb14b;
assign v22f3a35 = hlock0_p & v23f6411 | !hlock0_p & v230377f;
assign v22eb5a9 = hmaster2_p & v2309c8a | !hmaster2_p & v106ae19;
assign v23007d9 = hready_p & v23f15ba | !hready_p & v23f4ad7;
assign v230723b = hbusreq6_p & v23f437e | !hbusreq6_p & v23fbf84;
assign v22fe08f = hmaster0_p & v84562e | !hmaster0_p & v96c563;
assign v230932e = stateG2_p & v84561b | !stateG2_p & !v15071da;
assign v2301e8c = hmaster0_p & v22f25e6 | !hmaster0_p & v230ae9d;
assign v23fc23d = hready & v8e28ac | !hready & v84564d;
assign v22f3de9 = hlock2_p & v230d7b7 | !hlock2_p & !v84561b;
assign v22eb05f = hbusreq5_p & v22f6f2b | !hbusreq5_p & !v2310900;
assign v230573f = stateG10_5_p & v23f6575 | !stateG10_5_p & !v2309c8a;
assign v230dcef = hmaster2_p & v23fbaaa | !hmaster2_p & v22f01c1;
assign v1aae296 = hbusreq4_p & v2304e28 | !hbusreq4_p & v230f03c;
assign v22f2c8a = hgrant3_p & v22f368e | !hgrant3_p & v23042b7;
assign v22feca2 = hmaster1_p & v22fe1c8 | !hmaster1_p & v22f0b75;
assign v230f691 = hbusreq3 & v22fa58f | !hbusreq3 & v22edff5;
assign v23f7789 = hbusreq0 & v13afe3a | !hbusreq0 & !fc8ab7;
assign v22f1376 = hbusreq0_p & v230d1de | !hbusreq0_p & v84561b;
assign v2391b88 = hgrant1_p & v230f846 | !hgrant1_p & v22fed24;
assign v22ff192 = hmaster0_p & v22ffd0e | !hmaster0_p & v23f3f65;
assign v2309b39 = hbusreq5_p & v2306b2e | !hbusreq5_p & !v22efcd6;
assign v23fb701 = hlock6_p & v23f8a49 | !hlock6_p & v2304aae;
assign v2310c2b = stateA1_p & v84561b | !stateA1_p & v23fb564;
assign v22ecf16 = hmaster0_p & v2302177 | !hmaster0_p & v22ebce1;
assign v22f2114 = hmaster2_p & v2391f2b | !hmaster2_p & v230a562;
assign v2305838 = hlock1_p & v2305792 | !hlock1_p & v230abb1;
assign v23fc98a = hbusreq5_p & v23fcea8 | !hbusreq5_p & !v84561b;
assign v22f2363 = hlock1_p & v22fba3f | !hlock1_p & !v84561b;
assign v22ed2f0 = hgrant0_p & v17a34ff | !hgrant0_p & !v845647;
assign v22f7d5d = hbusreq5_p & v2306d29 | !hbusreq5_p & v106af73;
assign v230bf6d = locked_p & v22ebf47 | !locked_p & v84561b;
assign v22fc4af = hmaster0_p & v23106ba | !hmaster0_p & v191ae7e;
assign v22f9c73 = locked_p & v230ff13 | !locked_p & v10dbf64;
assign v230f6a7 = locked_p & v23083ed | !locked_p & v23040af;
assign v23fc5fb = hbusreq6 & v23f5dcc | !hbusreq6 & v84561b;
assign v22f78b7 = hbusreq1_p & v23fba24 | !hbusreq1_p & v231343f;
assign v22ebb5c = hbusreq3_p & v22f1963 | !hbusreq3_p & v2304060;
assign v22f6bba = jx1_p & v8d07e3 | !jx1_p & v23fcc25;
assign v22f6e0c = hbusreq1_p & v23fc220 | !hbusreq1_p & v23fbd76;
assign v22f515e = hbusreq3 & v22f8ad3 | !hbusreq3 & v22f5583;
assign v22f6844 = hbusreq3_p & v2309e12 | !hbusreq3_p & v22f0393;
assign v23fc818 = hlock5_p & v84561b | !hlock5_p & v23fc55d;
assign v2311c5d = hgrant5_p & v22f05f3 | !hgrant5_p & v22f4bec;
assign v23f855f = hbusreq3_p & v22fb428 | !hbusreq3_p & !v23fafca;
assign v22f1dec = hmaster1_p & v2312ea4 | !hmaster1_p & v230af39;
assign v12cc30c = hmaster2_p & v22f2b78 | !hmaster2_p & v22f7da7;
assign v2302933 = hlock0_p & v23f7218 | !hlock0_p & v22fcceb;
assign v22fccc4 = stateG2_p & v84561b | !stateG2_p & !v2310bf7;
assign v2302aac = hmaster2_p & v23fc112 | !hmaster2_p & !v84561b;
assign v22fe95c = hbusreq5 & v22fb77d | !hbusreq5 & !v23fc596;
assign v2303e1a = hlock5_p & v23f6411 | !hlock5_p & !v106ae19;
assign v23f1a43 = stateG10_5_p & v230b59f | !stateG10_5_p & v2309c93;
assign v23f3d09 = hmaster1_p & v23fbf14 | !hmaster1_p & v230fe54;
assign v23f4b35 = hbusreq1 & v2310c6d | !hbusreq1 & v22fbe28;
assign v23f7086 = hmaster0_p & v23fc5bc | !hmaster0_p & v22ec702;
assign v22ec1f4 = hmaster2_p & v22f878c | !hmaster2_p & v23fca52;
assign v23f354c = hbusreq2_p & v106a782 | !hbusreq2_p & v22ee4b6;
assign v23fcd24 = hmaster2_p & v191a879 | !hmaster2_p & !v2392d6d;
assign v22fe831 = hbusreq3 & v845620 | !hbusreq3 & v22fe2ae;
assign v2308e63 = busreq_p & v230d70b | !busreq_p & v23fca58;
assign v845667 = stateG3_2_p & v84561b | !stateG3_2_p & !v84561b;
assign v22f6e29 = hgrant5_p & v239253c | !hgrant5_p & v23fbe00;
assign v22eb665 = hbusreq3 & v23f6739 | !hbusreq3 & v23fbf0b;
assign v1e84b3e = hbusreq6_p & v23fc6f0 | !hbusreq6_p & v23fcaec;
assign v22f6b7d = hbusreq3 & v23fbab4 | !hbusreq3 & v84561b;
assign v23f232a = hmaster2_p & v23fc89a | !hmaster2_p & v22fc19c;
assign v22fa1af = hbusreq2 & v13afe8f | !hbusreq2 & v84561b;
assign v230960d = jx1_p & v22fc690 | !jx1_p & v23efe7d;
assign v23070c1 = hbusreq5_p & v22f56d2 | !hbusreq5_p & v230f63f;
assign v22f5fe4 = hbusreq4_p & v2308a1b | !hbusreq4_p & v23f28a1;
assign v22f2851 = hmaster0_p & v2306d08 | !hmaster0_p & v22feb8b;
assign v22f8ac3 = hbusreq2_p & v2300962 | !hbusreq2_p & !v84561b;
assign v23f039f = hbusreq2_p & v23f60ef | !hbusreq2_p & !v84561b;
assign v22f07e0 = hmaster1_p & v22f814e | !hmaster1_p & !v23f7ff2;
assign v231185d = hbusreq3_p & v2305782 | !hbusreq3_p & v22ff179;
assign v8ea3a5 = hmaster2_p & v23035ba | !hmaster2_p & v84561b;
assign v2306d08 = hgrant3_p & v22eb899 | !hgrant3_p & v23f13f3;
assign v230930b = hbusreq3 & v22eb51e | !hbusreq3 & v84561b;
assign v22f8b9c = stateG10_5_p & v22fa766 | !stateG10_5_p & v12cddb2;
assign v2304082 = hmaster0_p & v23fc3aa | !hmaster0_p & v22f8a46;
assign v22ed4e1 = hmaster2_p & v22f1a26 | !hmaster2_p & v23fbb80;
assign b0d6e5 = hbusreq1 & a1fd0b | !hbusreq1 & !v23f5d72;
assign v230a753 = hgrant5_p & v84561b | !hgrant5_p & v23fc632;
assign v230b961 = hlock0_p & v22f1a26 | !hlock0_p & v2392d6f;
assign v23fd04d = hbusreq4_p & v23f05ee | !hbusreq4_p & v23fc23c;
assign v23fc7ee = hbusreq2_p & v191ae6a | !hbusreq2_p & v845620;
assign v23efe10 = stateG2_p & v2302ca3 | !stateG2_p & v23f8ecc;
assign v23fbdb7 = hbusreq5_p & v845636 | !hbusreq5_p & v22faa24;
assign v23119e3 = hmaster2_p & fc8ab7 | !hmaster2_p & !v2304009;
assign v23efdd0 = hbusreq0 & v1aae56f | !hbusreq0 & v84564d;
assign v23fc46e = hmaster0_p & v23fb4ba | !hmaster0_p & v2306660;
assign v23fced7 = hbusreq2 & v22fc4d3 | !hbusreq2 & b9c8dc;
assign v23fcd6b = hmaster2_p & v22fca28 | !hmaster2_p & v2300271;
assign v2392833 = hbusreq5 & v22f79fd | !hbusreq5 & v84561b;
assign v23fb1c6 = hlock0_p & v9526ac | !hlock0_p & v23fcae8;
assign v2304332 = hbusreq4 & v2305f8e | !hbusreq4 & !v845622;
assign v2303679 = hgrant1_p & v23fb6ff | !hgrant1_p & v23063f8;
assign v22febde = hmaster0_p & v23fbe74 | !hmaster0_p & v23ef95a;
assign v230650d = stateG2_p & v84561b | !stateG2_p & v22f5fa8;
assign v230f1d9 = hmaster1_p & v1aae2c1 | !hmaster1_p & v22ffaf3;
assign v23fc93b = hbusreq1_p & v13afe3a | !hbusreq1_p & v845647;
assign v22ebb15 = hbusreq6_p & v23f6591 | !hbusreq6_p & v231359f;
assign v2307224 = hbusreq3 & v23070c0 | !hbusreq3 & v23fc1bc;
assign v23fc826 = hmaster0_p & v87d737 | !hmaster0_p & v23fcb9d;
assign v2304ec9 = hmaster2_p & v22feb6e | !hmaster2_p & v23fa345;
assign v22ed0f0 = hmaster0_p & v23fc437 | !hmaster0_p & v23001a6;
assign v23047dd = hbusreq6_p & v84561b | !hbusreq6_p & v230a1fa;
assign v2391d17 = hbusreq1_p & v230ac33 | !hbusreq1_p & !v84561b;
assign v23fb9c6 = hmaster2_p & v23fcf70 | !hmaster2_p & !v22ec782;
assign v23f18f2 = hmaster0_p & v23fcfb2 | !hmaster0_p & v230c117;
assign v23ef8bb = hgrant1_p & v23fb6ff | !hgrant1_p & v22eaaef;
assign v23098ce = hgrant6_p & v84561b | !hgrant6_p & v22f2d88;
assign v23fcb63 = hbusreq4_p & v2309b5d | !hbusreq4_p & v23fc33a;
assign v23f65cd = hbusreq4_p & v2393dd2 | !hbusreq4_p & v22fa11e;
assign v22ec078 = jx1_p & v85e5cf | !jx1_p & !v23fcc94;
assign v9585ce = hlock0_p & v22f343b | !hlock0_p & v22fc4d8;
assign v2312cdf = hgrant5_p & v23111c2 | !hgrant5_p & v23052cc;
assign v23f5893 = hbusreq3_p & v22f1d1f | !hbusreq3_p & v2302e1b;
assign v23051f6 = hmaster2_p & v2308880 | !hmaster2_p & af6dff;
assign v23f61e5 = hmaster2_p & b9d013 | !hmaster2_p & !v23fbb4b;
assign v22fcd0f = stateG10_5_p & v22f7f74 | !stateG10_5_p & v191a879;
assign v22f1d1f = hmaster2_p & v2310e40 | !hmaster2_p & v23fc904;
assign v2309790 = hbusreq3_p & v23f5fdb | !hbusreq3_p & !v84561b;
assign v230065d = hgrant5_p & v23041a1 | !hgrant5_p & v22f96f2;
assign v23fbe8b = hgrant5_p & v22f1279 | !hgrant5_p & v106af57;
assign v230420d = hlock3_p & v22f90d2 | !hlock3_p & !v84561b;
assign v22f8e56 = hbusreq6_p & v22fefa1 | !hbusreq6_p & v22eb134;
assign v22fd549 = hbusreq1 & v230a3af | !hbusreq1 & v84561b;
assign v23f111f = hbusreq6_p & v23fcdda | !hbusreq6_p & v23fb819;
assign v22fbd15 = hbusreq6 & v22fdcc7 | !hbusreq6 & v84561b;
assign v9ed9e1 = hmaster0_p & v22f8cb9 | !hmaster0_p & v23fccb5;
assign v23091e0 = hlock1_p & v23f6653 | !hlock1_p & !v106ae19;
assign v992f98 = hbusreq0 & v845620 | !hbusreq0 & !v84561b;
assign v23fcd91 = hbusreq4_p & v22f07ac | !hbusreq4_p & v84561b;
assign v23fb957 = hmaster0_p & v23fc6a1 | !hmaster0_p & v22f9ac5;
assign v23f8e04 = hmaster2_p & v845625 | !hmaster2_p & !v84561b;
assign v230204f = hburst0 & v22f3294 | !hburst0 & !v22faa1f;
assign v22f8107 = hgrant0_p & v23fc125 | !hgrant0_p & v23f4517;
assign v2308f80 = hgrant0_p & v230dc56 | !hgrant0_p & v84561b;
assign v23fc8ad = hbusreq6 & v23fc476 | !hbusreq6 & !v84561b;
assign v230313e = hmaster1_p & v22ee4eb | !hmaster1_p & !v22fca3a;
assign v230d9cf = hgrant1_p & v84561b | !hgrant1_p & v2304443;
assign v22f6a93 = hgrant0_p & v862ae0 | !hgrant0_p & !v84561b;
assign v230db9d = stateA1_p & v84561b | !stateA1_p & !v2302dd1;
assign v2300b4f = hgrant5_p & v22f950e | !hgrant5_p & v23f3115;
assign v230bf9f = hmaster2_p & v2307b39 | !hmaster2_p & v23fb6a4;
assign v23fb8fa = hbusreq5 & v23f2be7 | !hbusreq5 & v84561b;
assign v2304c4c = hgrant5_p & v23fc24a | !hgrant5_p & v2301482;
assign v230b1db = hbusreq5 & v22f1a26 | !hbusreq5 & v84561b;
assign v2312be1 = hgrant3_p & v84561b | !hgrant3_p & v23fcd63;
assign v23fc39c = hgrant5_p & v84561b | !hgrant5_p & v23f3fca;
assign v17a3514 = hbusreq4_p & v22ebd72 | !hbusreq4_p & v22f7347;
assign v23fc7a7 = hmaster2_p & v23126ae | !hmaster2_p & v23fc904;
assign v23f441d = hbusreq3_p & v9bcad3 | !hbusreq3_p & v23fbe76;
assign v23f60ef = hbusreq2 & v23025ab | !hbusreq2 & !v84561b;
assign v23fba61 = hgrant0_p & a1fba6 | !hgrant0_p & v23fb83c;
assign v23fce12 = jx1_p & v23065ee | !jx1_p & v84561b;
assign v2305050 = hbusreq5_p & v22f2c2c | !hbusreq5_p & v22efeed;
assign v23fba6a = jx1_p & v1aad346 | !jx1_p & v23052dd;
assign v22f636a = hlock3_p & v22ecc58 | !hlock3_p & v230685f;
assign v22f1b4e = locked_p & b9d00f | !locked_p & !v106ae19;
assign v23fbd0d = hmaster2_p & v23fb98a | !hmaster2_p & v84561b;
assign v22eef3b = jx0_p & v22ec078 | !jx0_p & !v23fc8ac;
assign v23fcf0e = hbusreq4 & v230c995 | !hbusreq4 & b9c90c;
assign v23075ce = hbusreq6 & v230d2b0 | !hbusreq6 & v23f1391;
assign v23f30b2 = hmaster2_p & v84561b | !hmaster2_p & v23f8d76;
assign b9c985 = hgrant3_p & v23fd00d | !hgrant3_p & v2312d0e;
assign v22fa4c3 = jx0_p & v22fe261 | !jx0_p & !v22ee7ee;
assign v2304c95 = hmaster1_p & ae3590 | !hmaster1_p & v23021d9;
assign v23fb1b4 = hbusreq2_p & v23fb9dc | !hbusreq2_p & v23f35c4;
assign v23fc5e5 = hlock4_p & v2393091 | !hlock4_p & v23f3e77;
assign v23f5f07 = hbusreq2_p & v22f46ab | !hbusreq2_p & !v84562a;
assign v22ec6c7 = hmaster0_p & v2301ac0 | !hmaster0_p & v2312679;
assign v22eb5cc = hgrant0_p & v23f4694 | !hgrant0_p & v22fd106;
assign ae1a21 = hmaster0_p & v23f40fd | !hmaster0_p & v23fc95c;
assign v22f8c2f = hbusreq1 & v23fb49a | !hbusreq1 & v23f87f4;
assign v22f26fc = hgrant1_p & v23fb2ea | !hgrant1_p & v2304ee5;
assign v22f8aea = hgrant3_p & v22efef6 | !hgrant3_p & v23f0cbe;
assign a04dcc = hlock3_p & v22f603b | !hlock3_p & v2313405;
assign v23043b8 = stateG10_5_p & v2306d9e | !stateG10_5_p & v845636;
assign v2303fb9 = hlock5_p & v23fb899 | !hlock5_p & v23fbf5f;
assign v23f4e63 = hgrant3_p & v2304919 | !hgrant3_p & v230067a;
assign v2303461 = hmaster2_p & v22fc96c | !hmaster2_p & v22ec71a;
assign v22fed90 = jx1_p & v230313e | !jx1_p & v23009d5;
assign v1aad4b7 = hbusreq4_p & v23fbd71 | !hbusreq4_p & v22fde04;
assign v22ef4de = hgrant3_p & v84561b | !hgrant3_p & v23f3f59;
assign v23fbac3 = hbusreq3_p & v22ee09d | !hbusreq3_p & v1e840fa;
assign v230f253 = hbusreq2_p & v23fba35 | !hbusreq2_p & v22f17eb;
assign v22f12e5 = hgrant1_p & v84564d | !hgrant1_p & !v22f991d;
assign v2305c78 = hbusreq3 & v22fb36e | !hbusreq3 & v84561b;
assign v22ecb12 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v22f56d2;
assign v22fff0a = hbusreq6 & v1aad39a | !hbusreq6 & v23f361e;
assign v23fc9d1 = hbusreq1_p & v2391d40 | !hbusreq1_p & b7b244;
assign v23fc37d = hbusreq5_p & v23fca0a | !hbusreq5_p & !v22f946f;
assign v23f56bc = hbusreq3 & v23fa215 | !hbusreq3 & b50a75;
assign fc8c27 = hbusreq5_p & v22fe1d9 | !hbusreq5_p & !v22faee9;
assign v22ef7a5 = hbusreq6 & v23f3d02 | !hbusreq6 & !v22f5198;
assign v23f9f71 = hready_p & v23f741e | !hready_p & !b11fc3;
assign v22f7375 = hmaster0_p & v22f7c44 | !hmaster0_p & v23fc3e1;
assign v150744b = hmaster0_p & af7272 | !hmaster0_p & !v23fb92b;
assign v23fc2ce = hgrant1_p & v22f7830 | !hgrant1_p & v22fb850;
assign v230dcf9 = hbusreq6 & v23f895d | !hbusreq6 & v22ff882;
assign v22feb8b = hgrant3_p & v23fbe02 | !hgrant3_p & v22fb773;
assign v23fcc1c = hmaster1_p & v22ee3ca | !hmaster1_p & v231045a;
assign v90c400 = hmaster2_p & v2305a12 | !hmaster2_p & v84561b;
assign v23fb166 = jx0_p & a452a3 | !jx0_p & v22f1cc5;
assign v23fc412 = hmaster0_p & v23f756e | !hmaster0_p & v23fc25a;
assign v23fb8ec = hmaster2_p & v23fc921 | !hmaster2_p & v22edc4f;
assign v22ee2b4 = hmaster2_p & v23fbe44 | !hmaster2_p & v2310e89;
assign v22fdbbb = hmaster0_p & v22fdd56 | !hmaster0_p & baa1eb;
assign bd951f = hgrant1_p & v22f3ed0 | !hgrant1_p & v1aae9e2;
assign v2310238 = hmaster2_p & v22fbd02 | !hmaster2_p & v22fabd2;
assign v230828c = hgrant0_p & v84561b | !hgrant0_p & v22f4700;
assign v22fe4a1 = hbusreq3_p & v230e89f | !hbusreq3_p & v84561b;
assign v22ebfcf = hgrant6_p & v22eb6c8 | !hgrant6_p & v23f36d3;
assign v23fbc9a = hbusreq3 & v23f7024 | !hbusreq3 & v84561b;
assign v23fbb58 = hlock6_p & v22f3dea | !hlock6_p & v2309305;
assign v2303886 = hmaster1_p & v23fc91d | !hmaster1_p & v84561b;
assign v890cdd = hbusreq2_p & v22ee9c4 | !hbusreq2_p & !v84561b;
assign v22fa39e = hbusreq4_p & v22fdf59 | !hbusreq4_p & v22f6053;
assign v230c653 = hbusreq4 & v23015de | !hbusreq4 & v84561b;
assign v23effa5 = hgrant5_p & v22f4bf4 | !hgrant5_p & v23fc539;
assign v22f65d5 = hlock0_p & v23fbffe | !hlock0_p & v23f4b28;
assign v1506a7a = jx0_p & v22fda63 | !jx0_p & v23096af;
assign v23f704d = hmaster2_p & v23fbf0d | !hmaster2_p & v23fbdc1;
assign v230bd05 = hgrant5_p & v2311dff | !hgrant5_p & v23fcf91;
assign a0f5d5 = hbusreq4_p & v23fbc9c | !hbusreq4_p & v23f3970;
assign v23077ec = hmaster2_p & v2313463 | !hmaster2_p & !v22fbf74;
assign v23fc1fe = hbusreq1 & v22fdf25 | !hbusreq1 & !v23fc614;
assign v22eaeab = hlock6_p & v23fceb9 | !hlock6_p & v84562b;
assign v22f004e = hlock5_p & v84564d | !hlock5_p & !v84561b;
assign v23fba42 = hmaster2_p & v23101b1 | !hmaster2_p & v239346f;
assign v22f3813 = hgrant2_p & v23f68d8 | !hgrant2_p & v84561b;
assign v22ff969 = hbusreq3_p & v22f34c1 | !hbusreq3_p & v23f8c0b;
assign v23f2a1a = stateG2_p & v2302ca3 | !stateG2_p & v2300edd;
assign v23f6c7c = hmaster0_p & v22f6629 | !hmaster0_p & v8b4671;
assign v2307e5a = hbusreq3 & v230f538 | !hbusreq3 & v84561b;
assign v23f572e = hgrant1_p & v22f9df1 | !hgrant1_p & v23fadf4;
assign v23fc69f = hbusreq6_p & v2391fc6 | !hbusreq6_p & v23fca4b;
assign v23fcb17 = hmaster2_p & v22f542d | !hmaster2_p & v22feae3;
assign v23fb593 = hlock3_p & v23ef915 | !hlock3_p & v2309733;
assign v23fcd97 = hmaster0_p & v22fda61 | !hmaster0_p & !v22ed6e1;
assign v230aa9b = hmaster1_p & v23fbf54 | !hmaster1_p & v23fd00e;
assign v23fbadd = hgrant5_p & v23f83ff | !hgrant5_p & !v84564f;
assign v23fbf24 = hbusreq2_p & v22ee660 | !hbusreq2_p & v845620;
assign v2308b14 = hbusreq3_p & v23fb578 | !hbusreq3_p & v23f7680;
assign v22f3f32 = hmaster2_p & v84561b | !hmaster2_p & v23fa0bf;
assign v22f8ec8 = hbusreq4 & v22f8cb7 | !hbusreq4 & v84561b;
assign v23f0b47 = hmaster2_p & v23101b1 | !hmaster2_p & v23fcae5;
assign v22fc964 = jx1_p & v2303982 | !jx1_p & v22ef78e;
assign v23fbb73 = hmaster2_p & v23f8928 | !hmaster2_p & v2301797;
assign v23f468c = hlock0_p & da38c1 | !hlock0_p & v84561b;
assign v230e71d = hgrant3_p & v22f8e29 | !hgrant3_p & v230d910;
assign v9e23c0 = hmaster0_p & v23f7f9d | !hmaster0_p & !v96c563;
assign v23fbd14 = hgrant1_p & v2305fe0 | !hgrant1_p & !v84561b;
assign v22f4bf5 = jx0_p & v84561b | !jx0_p & v23fc4dd;
assign v230fb43 = hbusreq3 & v23f9a81 | !hbusreq3 & v23fce7e;
assign v22fd3f7 = hgrant2_p & v22fb877 | !hgrant2_p & !v2301d10;
assign v22f5c2b = hmaster0_p & v22ed711 | !hmaster0_p & !v2302460;
assign v230d7e2 = jx2_p & v230c24b | !jx2_p & v23f5c03;
assign v23047f9 = jx1_p & v23fbc28 | !jx1_p & !v22f443a;
assign v2303982 = hmaster1_p & v23fc1db | !hmaster1_p & v23fb73e;
assign v23f619e = hlock1_p & v22ed751 | !hlock1_p & !v84561b;
assign v2308967 = hmaster2_p & v84561b | !hmaster2_p & v230a4b6;
assign v22f88c3 = hmaster2_p & v84561b | !hmaster2_p & v22f8d74;
assign v23055d9 = hmaster1_p & v23fc1be | !hmaster1_p & v230e086;
assign v22fba41 = hmaster2_p & v23f4b28 | !hmaster2_p & v23f6bc1;
assign v22f89b9 = hmaster2_p & v84561b | !hmaster2_p & v22ee8f3;
assign v22fcbac = hbusreq5_p & v230e4ef | !hbusreq5_p & v1aad518;
assign aa51ef = jx1_p & v22f04eb | !jx1_p & v230cd1c;
assign v22f5efe = hmaster0_p & v230e95c | !hmaster0_p & v2301306;
assign v230eeb5 = hbusreq3 & v23fc7e7 | !hbusreq3 & v2302131;
assign v23028fc = hmaster2_p & v23fc4f8 | !hmaster2_p & v23fcbcd;
assign v230e85f = hmaster2_p & v22eec6e | !hmaster2_p & v84561b;
assign v230b621 = hgrant1_p & v12cd9f9 | !hgrant1_p & !v23fc6ca;
assign v23058da = hgrant5_p & v84561b | !hgrant5_p & !v23fcc50;
assign v23faae7 = hbusreq3_p & v23fbadb | !hbusreq3_p & v23f86dc;
assign v12cda44 = stateA1_p & v84561b | !stateA1_p & !v23fc8a3;
assign v230b111 = hgrant3_p & v84561b | !hgrant3_p & v2303c10;
assign v230b981 = hbusreq5_p & a1fcbb | !hbusreq5_p & v84561b;
assign v23fb33a = hbusreq1_p & v23fb788 | !hbusreq1_p & v23f7796;
assign v22ee4fe = hlock0_p & v2306b74 | !hlock0_p & !v23f9ce3;
assign v2300755 = hmastlock_p & v2307460 | !hmastlock_p & v84561b;
assign v22ebf17 = hbusreq1 & v1aae087 | !hbusreq1 & v84561b;
assign v23929fd = hbusreq6_p & v2312dc5 | !hbusreq6_p & v23043b1;
assign v23038cc = hgrant4_p & v230592c | !hgrant4_p & !v84561b;
assign v22f03c8 = hbusreq6 & v23fc64c | !hbusreq6 & !v845622;
assign v2305684 = stateG10_5_p & v1e84012 | !stateG10_5_p & v22f3643;
assign v22f6d19 = hmaster2_p & v22fdc30 | !hmaster2_p & v230f63f;
assign v23fc882 = hbusreq2_p & v23fb0ba | !hbusreq2_p & !v23f86f0;
assign v22ff8ea = hbusreq0 & v1aae362 | !hbusreq0 & !v84561b;
assign v22eb265 = hmaster0_p & v23f54a0 | !hmaster0_p & !v23fbf74;
assign v23fc846 = hgrant3_p & v231330b | !hgrant3_p & v23f832b;
assign v23044cf = hmaster2_p & v23f5af5 | !hmaster2_p & v23f6411;
assign v2303253 = jx1_p & v22f8291 | !jx1_p & v84561b;
assign v2391b32 = hbusreq5_p & v84561b | !hbusreq5_p & !v230404f;
assign v22fa827 = hbusreq2_p & v22efd1a | !hbusreq2_p & v23fc199;
assign v22eb52b = hmaster0_p & be29ff | !hmaster0_p & v2300382;
assign v23f2fb7 = hbusreq3_p & v845645 | !hbusreq3_p & !v84561b;
assign v2301b99 = hbusreq4_p & v22ec502 | !hbusreq4_p & v22fd032;
assign v106aeed = hbusreq3_p & v23064ca | !hbusreq3_p & v84561b;
assign v23f55a4 = hmaster1_p & v230a407 | !hmaster1_p & v23068bb;
assign v23f2f45 = stateG2_p & v84561b | !stateG2_p & v22f197e;
assign b84511 = hbusreq3_p & v22f695c | !hbusreq3_p & v22ecab8;
assign v22eb3fd = hbusreq6 & v1e84038 | !hbusreq6 & !v23135a4;
assign v231253d = hmaster0_p & v22fba38 | !hmaster0_p & v23fc347;
assign v23fc99c = hbusreq4 & v22ee9be | !hbusreq4 & v84561b;
assign v23fb63f = hbusreq6 & v22f7e21 | !hbusreq6 & v84561b;
assign v2307bcb = hbusreq4_p & v23f46d8 | !hbusreq4_p & v12cd552;
assign v22f0545 = hmaster2_p & v23fb1a4 | !hmaster2_p & !v23fbb80;
assign v2309d59 = hmaster2_p & v13afb18 | !hmaster2_p & v22f926d;
assign v23fc3dd = hgrant5_p & v22f1905 | !hgrant5_p & !v23fb1d1;
assign v22f2624 = hbusreq1 & v23fbbf2 | !hbusreq1 & v845622;
assign v22fae9f = hmaster0_p & v22f336f | !hmaster0_p & v23f593e;
assign v22fbeea = hlock0_p & v22f13cb | !hlock0_p & v22f3789;
assign v23fc9aa = hbusreq5_p & v23f2a86 | !hbusreq5_p & v84561b;
assign v23fcf07 = hbusreq6 & v22fc0a4 | !hbusreq6 & !v84562a;
assign v22f30fe = hbusreq1 & v22f15fe | !hbusreq1 & v23f60ef;
assign v22fa73a = hbusreq3_p & v22f61f6 | !hbusreq3_p & v13aff86;
assign v23fc7d9 = hbusreq4_p & v22ff29f | !hbusreq4_p & v23fb533;
assign b00aa6 = hgrant3_p & v84561b | !hgrant3_p & v22f1244;
assign v22eb22e = hbusreq6 & v2301044 | !hbusreq6 & !v23fbeeb;
assign v230bd1c = hbusreq6_p & v23f4117 | !hbusreq6_p & v22ebc26;
assign v230faa5 = hgrant5_p & v2308b08 | !hgrant5_p & v230ff63;
assign v23fb615 = hmaster0_p & v22ede0b | !hmaster0_p & v22efc7f;
assign v22eafb2 = hbusreq1_p & v23fb591 | !hbusreq1_p & v90b913;
assign v2312628 = jx1_p & v85e5cf | !jx1_p & !v2391b34;
assign v22f397b = hbusreq6_p & v230a241 | !hbusreq6_p & v22feff6;
assign v23fc3b3 = hbusreq1_p & v23fbaf3 | !hbusreq1_p & v191aada;
assign v94508c = hbusreq6 & v2312888 | !hbusreq6 & v84561b;
assign v23fc9e4 = hlock3_p & v84561b | !hlock3_p & !v2309790;
assign v23126e2 = hgrant3_p & v84561b | !hgrant3_p & v230e37a;
assign a3cb61 = hgrant1_p & v23fb67c | !hgrant1_p & v2304672;
assign v23f507b = hmaster0_p & v23f1a86 | !hmaster0_p & bdeff3;
assign v2311be9 = hgrant1_p & v84561b | !hgrant1_p & v22fc723;
assign v23fcab7 = hbusreq3_p & v22f695c | !hbusreq3_p & v23fc365;
assign v23fcc35 = hmaster2_p & v2304b35 | !hmaster2_p & !v22ff05e;
assign v23f8345 = hbusreq3 & v230fb9e | !hbusreq3 & v845627;
assign v23f8357 = hbusreq1_p & v22f75d4 | !hbusreq1_p & v22f77e4;
assign v2313637 = jx3_p & v1aae1af | !jx3_p & v2303841;
assign v22f291f = hbusreq1_p & v22f3e93 | !hbusreq1_p & v2307205;
assign v22fdd8a = hbusreq6 & v23fb865 | !hbusreq6 & v84562a;
assign v230e606 = hbusreq0 & v23f3a55 | !hbusreq0 & v84561b;
assign v230fe6b = hmaster0_p & v22f368e | !hmaster0_p & v23fbebe;
assign v22fbd4f = hbusreq4 & v23f87e1 | !hbusreq4 & v84561b;
assign v22f9bc8 = hmaster2_p & v23fa2b5 | !hmaster2_p & v84561b;
assign v23fc638 = jx1_p & v22f8d2f | !jx1_p & v230cc95;
assign v22fa5f9 = hmaster2_p & v22ecbbd | !hmaster2_p & v230af38;
assign v2391e3e = hbusreq6 & v23f60fb | !hbusreq6 & v23f6404;
assign v1aadf44 = hmaster2_p & b9d00f | !hmaster2_p & a1fba6;
assign v23f6723 = hmaster0_p & v22f8e29 | !hmaster0_p & v230e979;
assign v22fdc60 = hburst1_p & v230371b | !hburst1_p & !v22ed56a;
assign b9d013 = hmastlock_p & v23f4b56 | !hmastlock_p & !v84561b;
assign v22ee1e6 = hbusreq0_p & v22ee2bb | !hbusreq0_p & v84561b;
assign v23f5388 = hbusreq6_p & v22fd364 | !hbusreq6_p & v23f5dfe;
assign v22ef354 = hbusreq6_p & v84561b | !hbusreq6_p & v22f1971;
assign v22ef5f1 = hgrant3_p & v23fd019 | !hgrant3_p & v23f60fb;
assign v23fb83c = hlock0_p & v23009cc | !hlock0_p & v1aadb95;
assign v23067de = hbusreq3_p & v2307e5a | !hbusreq3_p & v84561b;
assign v22f2fe1 = hlock3_p & v84561b | !hlock3_p & !v23fca7a;
assign v230c32e = jx1_p & v23fc0a7 | !jx1_p & v23055d9;
assign v22eafaa = hmaster0_p & v23096f8 | !hmaster0_p & v22ebd1b;
assign v23fc4e2 = hbusreq4_p & v23f6c83 | !hbusreq4_p & v23f74b7;
assign v22f3618 = hbusreq1_p & v22f0c1b | !hbusreq1_p & v84561b;
assign v23fb82c = hgrant0_p & v22ffb9d | !hgrant0_p & !v8ce364;
assign v22f8e0c = hbusreq3_p & v23049f8 | !hbusreq3_p & v22fe792;
assign locked = v1aacf10;
assign v2311743 = hgrant3_p & v2301b00 | !hgrant3_p & v23fc8d4;
assign v23fc273 = hmaster2_p & v230e8d3 | !hmaster2_p & v230e916;
assign v230e4ae = hgrant5_p & v230cfba | !hgrant5_p & v23fc19d;
assign v2308848 = hgrant2_p & v84564d | !hgrant2_p & v2303f9a;
assign v22f9df1 = hbusreq1_p & v23fcf46 | !hbusreq1_p & !v23fba6b;
assign b8f86b = hgrant6_p & v84561b | !hgrant6_p & v845639;
assign v23fc578 = hbusreq5_p & v23f6411 | !hbusreq5_p & v23fc503;
assign v23f7ad1 = hbusreq6 & v23fc176 | !hbusreq6 & v84561b;
assign v23f2513 = hgrant1_p & v84561b | !hgrant1_p & v2308f3d;
assign v23fcd8a = hbusreq3 & v23fc121 | !hbusreq3 & v2301319;
assign v23fce7d = hbusreq3_p & v84571e | !hbusreq3_p & !v84561b;
assign v23fcaa7 = hgrant4_p & v23fb679 | !hgrant4_p & v230cc50;
assign v23fc9c4 = hbusreq5_p & v845636 | !hbusreq5_p & v91ba6f;
assign v23f7e51 = hbusreq3 & v23fc068 | !hbusreq3 & !v84561b;
assign v22ff1cb = hbusreq4_p & v2312ebe | !hbusreq4_p & v23fcd97;
assign v230ddf3 = hmaster2_p & v84564d | !hmaster2_p & v22f4e0b;
assign v22ebe70 = hmaster1_p & v239223a | !hmaster1_p & v2303bf6;
assign v22f1154 = jx3_p & v23f47ae | !jx3_p & v23f6d75;
assign v22fc68e = jx3_p & v84561b | !jx3_p & v230dbcc;
assign v230c97c = hmaster2_p & a1fbb6 | !hmaster2_p & v22edc8d;
assign v22ef0de = hbusreq3_p & v22f2a2f | !hbusreq3_p & v23fcb7c;
assign v23fcf11 = hmaster0_p & v23fc99e | !hmaster0_p & v22f03c1;
assign v23128f3 = hbusreq6_p & v22ee8dd | !hbusreq6_p & v22f1d4f;
assign v2311d52 = hmaster2_p & v23f9414 | !hmaster2_p & v2309cdc;
assign v23f0329 = hgrant1_p & v2301511 | !hgrant1_p & b15a69;
assign v23fca35 = jx1_p & v2304764 | !jx1_p & v23fcaf8;
assign v23fc89a = hlock0_p & v22fda49 | !hlock0_p & !v845622;
assign v2392229 = hgrant5_p & v22fb8df | !hgrant5_p & !v2308356;
assign v1aae2be = hmaster2_p & v23fce57 | !hmaster2_p & v1507009;
assign v23fb54f = hgrant1_p & v84561b | !hgrant1_p & v23fbf1d;
assign v22fd124 = hbusreq1_p & bc5d21 | !hbusreq1_p & v2308bcd;
assign v2393ac5 = hbusreq5_p & v22f15fe | !hbusreq5_p & v230be24;
assign v2312d48 = stateG2_p & v84561b | !stateG2_p & v23fb8c0;
assign v23fc26a = hmaster0_p & v2306fba | !hmaster0_p & !v23fc02a;
assign v23fc3c3 = stateG10_5_p & v23fc19d | !stateG10_5_p & v845620;
assign v9ec6b5 = hgrant5_p & v22efa49 | !hgrant5_p & v23fc153;
assign v23fc3fa = hbusreq5 & v230e4ef | !hbusreq5 & v2391d40;
assign v2302d12 = hbusreq4_p & v12cd51b | !hbusreq4_p & v23fc9b2;
assign v2301655 = hbusreq2 & v22f814a | !hbusreq2 & !v84561b;
assign v23fc6a8 = hbusreq3_p & v8819d8 | !hbusreq3_p & v22f9023;
assign v22ff650 = hmaster0_p & v23f1a14 | !hmaster0_p & v22f25a1;
assign v23fc461 = hbusreq1_p & v2308d09 | !hbusreq1_p & !v22ffc69;
assign v23fb825 = hbusreq5 & v22f3643 | !hbusreq5 & v845620;
assign v2309d7a = hbusreq6_p & v22f0768 | !hbusreq6_p & v230025c;
assign v23fbf8e = hgrant3_p & v22fc6b9 | !hgrant3_p & v22f83fb;
assign v2367a45 = hbusreq1_p & v2310bf5 | !hbusreq1_p & !v84561b;
assign v230e165 = hbusreq1 & v23f63ab | !hbusreq1 & !v845636;
assign v23f0eeb = hgrant2_p & v230d5f4 | !hgrant2_p & v17a34f8;
assign v22ec9ce = hbusreq1_p & v23f2b6d | !hbusreq1_p & v2309c93;
assign v22f5088 = hlock3_p & v23f5927 | !hlock3_p & !v84561b;
assign v230e860 = hmaster2_p & v2391a57 | !hmaster2_p & !v84564d;
assign v23fc5bc = hbusreq6 & v22ebd72 | !hbusreq6 & v22f7347;
assign v22eb15f = hbusreq6_p & v2307a21 | !hbusreq6_p & v230d0ed;
assign v23f404a = hbusreq2 & v23f7efd | !hbusreq2 & v23fc1c9;
assign v2393f0d = hbusreq0_p & v22eefab | !hbusreq0_p & v23fc7ff;
assign v23f561c = hbusreq4 & v2307206 | !hbusreq4 & v845627;
assign v23f6038 = hbusreq5_p & v23fbb0f | !hbusreq5_p & v23fcce3;
assign v22f5840 = hmaster2_p & v22f0073 | !hmaster2_p & v22fda32;
assign v230a2bb = hgrant5_p & v22fa945 | !hgrant5_p & v230a941;
assign v2308f89 = hmaster0_p & v23fcbfb | !hmaster0_p & v23fad33;
assign v22f3c3d = hgrant0_p & v845622 | !hgrant0_p & v23fc1de;
assign v22ee413 = hmaster0_p & v845629 | !hmaster0_p & v23fcb28;
assign v22faac8 = stateA1_p & v23fc8a3 | !stateA1_p & v2302dd1;
assign v22f7e09 = hmaster2_p & v23fc5f4 | !hmaster2_p & v84561b;
assign v22f38db = hgrant3_p & v22f8985 | !hgrant3_p & v23f8607;
assign v22f5d45 = hmaster0_p & v23f3ce8 | !hmaster0_p & !v96c563;
assign v23f76d0 = hbusreq1_p & v22eece2 | !hbusreq1_p & !v22f5e45;
assign v230c6f1 = hlock6_p & v23034a4 | !hlock6_p & v8a6d1a;
assign ab39f4 = hbusreq4 & v22fe0a8 | !hbusreq4 & v22f28df;
assign v2311d12 = hbusreq5_p & v22f0051 | !hbusreq5_p & v84561b;
assign v22fcb7b = hmaster2_p & v22ed7a8 | !hmaster2_p & v22ffbb3;
assign v23fbff5 = hready_p & v23f1c12 | !hready_p & !v22fd0fb;
assign v231285b = hmaster2_p & v2300246 | !hmaster2_p & v84561b;
assign v845627 = hlock1_p & v84561b | !hlock1_p & !v84561b;
assign v22eb25c = hmaster2_p & v84561b | !hmaster2_p & v22f4e94;
assign v2302c6d = hlock3_p & v22ed925 | !hlock3_p & v23fc030;
assign v22f65c9 = jx1_p & v22fe1c8 | !jx1_p & v23f8186;
assign v23fcfae = hmaster2_p & v22f8235 | !hmaster2_p & !v2310271;
assign v23050c1 = hmaster2_p & v2304283 | !hmaster2_p & v23fbaaa;
assign v22ecbb2 = hbusreq3 & v23fbbec | !hbusreq3 & v22eec21;
assign v22fa027 = hready & v1aae294 | !hready & v22f197e;
assign v22fdb21 = hburst0_p & v23fc116 | !hburst0_p & !v22eff0e;
assign v2304da3 = jx2_p & v22ebf90 | !jx2_p & bb5cd7;
assign v230f75a = hbusreq1 & v22f65d5 | !hbusreq1 & v22f5583;
assign aaca7f = hmaster2_p & v22fcdf6 | !hmaster2_p & v22f9911;
assign ab4e4e = hlock5_p & v23fb598 | !hlock5_p & !v84561b;
assign v1aae0dc = hmaster1_p & v23fb0eb | !hmaster1_p & v2391735;
assign v22f4016 = hbusreq3_p & v23f80cc | !hbusreq3_p & v23fccd4;
assign v2300b80 = hgrant3_p & v230f165 | !hgrant3_p & v22febe7;
assign v230e2bb = hmaster2_p & v23fb9a9 | !hmaster2_p & v22efa93;
assign v23fbf97 = hmaster2_p & v8be441 | !hmaster2_p & !v23fa345;
assign v22eed5b = hgrant0_p & v22f3643 | !hgrant0_p & v23fb56e;
assign v23fb6a0 = jx1_p & v23fa1cd | !jx1_p & v22f6fba;
assign v22f5e63 = stateG10_5_p & v22f532c | !stateG10_5_p & v23f86f0;
assign v230464b = hbusreq1 & v23fb527 | !hbusreq1 & !v22fbe28;
assign v95fb82 = hbusreq4_p & v23fc3b8 | !hbusreq4_p & !v8fb6b6;
assign v22faefb = hlock5_p & v23f5cb3 | !hlock5_p & v23fbfb9;
assign v22f65c0 = hbusreq5_p & v230e07d | !hbusreq5_p & v23fc849;
assign v22f5974 = stateG10_5_p & v22f299f | !stateG10_5_p & v22eecf9;
assign v8bc4e1 = hmaster0_p & v22ec77a | !hmaster0_p & v22fb88d;
assign v23fb994 = hbusreq4 & v23f6470 | !hbusreq4 & v23fa2ec;
assign v2301b0c = hmaster1_p & v22fd532 | !hmaster1_p & v230cff8;
assign v23fbf1a = hbusreq5_p & v230e100 | !hbusreq5_p & v2307ab1;
assign v22f61ac = hgrant1_p & v23fb6ff | !hgrant1_p & v2302b3f;
assign v22f8fc0 = hbusreq5_p & v12cd93a | !hbusreq5_p & v84561b;
assign v99b664 = hmaster0_p & v23075dd | !hmaster0_p & !v230d674;
assign v23fcb99 = hmaster2_p & v22fa652 | !hmaster2_p & v2307d4e;
assign v191ab52 = hgrant3_p & v2310222 | !hgrant3_p & v22f4a4f;
assign b62970 = hbusreq5 & v22fafe4 | !hbusreq5 & v84561b;
assign v230cf0c = hgrant1_p & v84561b | !hgrant1_p & v2311899;
assign v23f5d34 = hbusreq1_p & v2391d40 | !hbusreq1_p & a1b75e;
assign v230ec10 = hbusreq5 & v22ed878 | !hbusreq5 & v84561b;
assign v191a90b = hburst0 & v22f80ca | !hburst0 & !v84561b;
assign v230f069 = hbusreq4_p & v23fc2da | !hbusreq4_p & v22f63e9;
assign v2309d7f = hlock3_p & v230a84b | !hlock3_p & v23fc2ae;
assign v23fbc3d = hmaster0_p & v23095df | !hmaster0_p & !v96c563;
assign v22f334e = stateG2_p & v22ec1cb | !stateG2_p & v23fb564;
assign v23f14c7 = hready_p & v23046fe | !hready_p & v23051ab;
assign v2312e30 = jx0_p & v23fcd83 | !jx0_p & v2304bcd;
assign v23fc7b4 = hbusreq3 & v23fb8e0 | !hbusreq3 & v84561b;
assign v23fc614 = hbusreq5_p & v845622 | !hbusreq5_p & v23fc839;
assign v22fbe99 = hbusreq5_p & v15071a5 | !hbusreq5_p & !v23fc463;
assign v23f471a = hbusreq1_p & v22f1faf | !hbusreq1_p & !v84561b;
assign v230c4c3 = hmaster2_p & v23fba6b | !hmaster2_p & v191a86f;
assign v23fbf8b = hgrant1_p & v23fc393 | !hgrant1_p & v230aa0d;
assign v2307701 = hmaster2_p & v23f7968 | !hmaster2_p & v22f954f;
assign v230e703 = hbusreq4_p & v23f7f51 | !hbusreq4_p & v22ee8dd;
assign v23fbcca = hbusreq3_p & v23f6588 | !hbusreq3_p & v22fc1e9;
assign v23fb9d6 = hgrant3_p & v22f2ca2 | !hgrant3_p & v230bdb9;
assign v22fa63e = hgrant6_p & v845635 | !hgrant6_p & v22ed92a;
assign v22fd559 = hmaster0_p & v22fba38 | !hmaster0_p & v23f6cdb;
assign v2302167 = hgrant5_p & v23f65bb | !hgrant5_p & v23133bb;
assign v230ee28 = stateG10_5_p & v22f61cc | !stateG10_5_p & v22edee1;
assign v22f2aff = hbusreq6 & v23fbcaa | !hbusreq6 & v22ee657;
assign v150730e = hgrant3_p & v22f690f | !hgrant3_p & v8a34ca;
assign v23fcda9 = hbusreq5_p & v22fb07c | !hbusreq5_p & v84561b;
assign v22fd663 = hmaster2_p & v895ae7 | !hmaster2_p & v84561b;
assign v23fbf6b = hmaster0_p & v22f2677 | !hmaster0_p & !v22eb933;
assign v2309561 = hmaster0_p & v22eef3f | !hmaster0_p & v2312e4e;
assign v23f34d4 = hlock0_p & v23fc8ee | !hlock0_p & !v84561b;
assign v2311196 = hmaster0_p & c1f7e4 | !hmaster0_p & !v23f89d9;
assign v22fbc0e = hbusreq4 & v22f9657 | !hbusreq4 & v84561b;
assign v23fba96 = hmaster2_p & v230eb9b | !hmaster2_p & v22fbf74;
assign a136c1 = hmaster2_p & v22f4114 | !hmaster2_p & v23f368a;
assign v23fbfaf = busreq_p & v22ee516 | !busreq_p & v845647;
assign v22fb68b = hbusreq5_p & v23f9c72 | !hbusreq5_p & v23fc5b0;
assign v2302a8c = hbusreq5 & c258f4 | !hbusreq5 & v84561b;
assign v23fa460 = hmaster0_p & v2312eaa | !hmaster0_p & !v23068cd;
assign v23fc78a = hmaster0_p & v23f592d | !hmaster0_p & v150730e;
assign v22f8f70 = jx3_p & v23f77a4 | !jx3_p & v23fcfd1;
assign v23fbcc7 = hlock0_p & v22ebee0 | !hlock0_p & a92d05;
assign v22fa7f5 = hbusreq0 & v191accc | !hbusreq0 & v23fc1de;
assign v2301585 = hgrant1_p & v230f9db | !hgrant1_p & v23fb6cf;
assign v23fc5db = hlock6_p & v239196f | !hlock6_p & !v23f14ce;
assign v23f4cc5 = hbusreq3_p & v8dd9c7 | !hbusreq3_p & aba695;
assign v22f9a51 = hmastlock_p & v2311f53 | !hmastlock_p & v84561b;
assign v23efa52 = hmastlock_p & v230d04a | !hmastlock_p & !v84561b;
assign v23fbf67 = hbusreq5 & v23fc4a5 | !hbusreq5 & v22f0add;
assign v22fd0fa = hgrant3_p & v230630c | !hgrant3_p & v23f5cfe;
assign v23fc50a = hbusreq6 & v22fea26 | !hbusreq6 & !v845625;
assign v22ecdc8 = hbusreq4_p & v2307170 | !hbusreq4_p & v23f95ba;
assign v22f3738 = hbusreq1_p & v23fb9c5 | !hbusreq1_p & v22f878c;
assign v23fc881 = hmaster2_p & v23fc765 | !hmaster2_p & v23f6c84;
assign v22ebe99 = hmaster2_p & v23fceb9 | !hmaster2_p & v22eefab;
assign v191b1e4 = hbusreq3 & v23071cd | !hbusreq3 & v84561b;
assign v23f9a37 = hgrant5_p & v230115b | !hgrant5_p & v22fe150;
assign v22f4d74 = hmaster2_p & v2300c47 | !hmaster2_p & v22f01c5;
assign v22ef0c8 = hlock3_p & v22fb511 | !hlock3_p & v2303674;
assign v22f6b4e = hbusreq4_p & v23f2856 | !hbusreq4_p & v23f37b9;
assign v22ecec6 = stateG10_5_p & v230ae19 | !stateG10_5_p & v2309c93;
assign v22f2718 = busreq_p & v23fbff3 | !busreq_p & v23fc2dd;
assign v23fcc08 = hmaster2_p & v23f3ccf | !hmaster2_p & v22ef46e;
assign v2300711 = hbusreq2 & v15071c2 | !hbusreq2 & !v23fb9be;
assign v23f2578 = hbusreq3_p & v1e83f8d | !hbusreq3_p & v23fcd66;
assign v230bc0c = hgrant0_p & v2306441 | !hgrant0_p & v22f1992;
assign v23122bc = hbusreq6_p & v23f7ef4 | !hbusreq6_p & v22f5a27;
assign v23fc048 = hmaster2_p & v9526ac | !hmaster2_p & v23fb875;
assign v22fe34f = hmaster2_p & v23fc71d | !hmaster2_p & v22f0945;
assign v22fa055 = hmaster2_p & v845647 | !hmaster2_p & !v2303393;
assign v22efa17 = hgrant1_p & v230feae | !hgrant1_p & v2307ab9;
assign v23fc9b4 = hmaster0_p & v23fb62d | !hmaster0_p & v2304048;
assign v230e3a0 = hgrant1_p & v84561b | !hgrant1_p & v22f64de;
assign v23131fd = hlock6_p & v23fca31 | !hlock6_p & v84561b;
assign v2310b4d = hbusreq6_p & v2391fc6 | !hbusreq6_p & v23fc329;
assign v22f343b = hbusreq2 & v22f7efa | !hbusreq2 & v84561b;
assign v23fccd3 = hbusreq6_p & v23f9b8f | !hbusreq6_p & !v84561b;
assign v2308b08 = hbusreq5_p & v22ed467 | !hbusreq5_p & !v22f5e63;
assign v1e840d3 = hlock0_p & b9d00f | !hlock0_p & v23fcdc0;
assign v22f7b13 = hbusreq5_p & v23fd064 | !hbusreq5_p & v230ee7d;
assign v22fb32a = hmaster2_p & v23fbd52 | !hmaster2_p & v23101b1;
assign v23fb054 = hlock2_p & v1aae56f | !hlock2_p & v84564d;
assign v23f9ce3 = hbusreq0 & v2301655 | !hbusreq0 & v84562a;
assign v230952f = hbusreq3_p & v23fc5ab | !hbusreq3_p & v23fc555;
assign v22ebffc = stateG2_p & v84561b | !stateG2_p & !v23fc8a3;
assign v23fbcb2 = hlock0_p & v22f3be4 | !hlock0_p & !v84561b;
assign v22f1117 = hbusreq3_p & v23f9758 | !hbusreq3_p & a0de1c;
assign v23f443c = jx1_p & v23f23f4 | !jx1_p & v22f1dec;
assign v230b780 = hbusreq0 & v13afe3a | !hbusreq0 & v845647;
assign v23f6dc8 = hbusreq2 & v15071c2 | !hbusreq2 & !fc8f74;
assign v23fb8cc = hbusreq3_p & v23fb60a | !hbusreq3_p & v23fcebf;
assign v22f4986 = hbusreq1_p & v191a876 | !hbusreq1_p & v191a879;
assign v230e3c5 = hbusreq3_p & v22ff538 | !hbusreq3_p & v23f660f;
assign v23fb561 = hbusreq1 & v1506ffd | !hbusreq1 & v22f1ece;
assign v23f65eb = hmaster2_p & v9d8aae | !hmaster2_p & !v23f8f21;
assign v23fc610 = hbusreq3_p & v2300f82 | !hbusreq3_p & v106ae19;
assign v23f8fd7 = hready_p & v22f3673 | !hready_p & v230de17;
assign v230d1de = hbusreq0 & v23fb978 | !hbusreq0 & v84561b;
assign v23f120d = hlock3_p & v22f2450 | !hlock3_p & v23fce8e;
assign v22ecca9 = hmaster2_p & v23f15ac | !hmaster2_p & v23f9e4f;
assign v23fbcc4 = hbusreq3 & v22fdf30 | !hbusreq3 & !v84561b;
assign v23fb074 = hbusreq3 & v22eca5d | !hbusreq3 & v84561b;
assign v2302460 = hmaster2_p & v2310e40 | !hmaster2_p & v23070c1;
assign e1d75b = hgrant3_p & v84561b | !hgrant3_p & v23fc58d;
assign v1aad31c = hbusreq3 & v23f2a5b | !hbusreq3 & v22ed5be;
assign v230e19d = hbusreq3 & v22eb8ad | !hbusreq3 & !v2301a90;
assign v2302e43 = hmaster2_p & v22ec921 | !hmaster2_p & !v84561b;
assign v23056bf = hbusreq3 & v23fbd2a | !hbusreq3 & b50a75;
assign v230e0d6 = hmaster2_p & v13afc17 | !hmaster2_p & v23f9f77;
assign v230e0c0 = hmaster0_p & v15072cc | !hmaster0_p & v2303a53;
assign v22fab80 = hgrant0_p & v845622 | !hgrant0_p & v23fc9c1;
assign v23f7f02 = hmaster2_p & v84561b | !hmaster2_p & v2304536;
assign v2309963 = stateG10_5_p & v22f4d04 | !stateG10_5_p & !v22fa5c9;
assign v1e84012 = hgrant0_p & v22f3643 | !hgrant0_p & v23fc01c;
assign v23f2fe0 = hburst0 & v22ec1cb | !hburst0 & !v84561b;
assign v22fdfde = hmaster2_p & v23f5cb3 | !hmaster2_p & !v23070c1;
assign v23f84dc = hbusreq6_p & v23fbba0 | !hbusreq6_p & v23fc7d9;
assign v22fbea4 = hbusreq0 & v22f60c6 | !hbusreq0 & !v2304ec7;
assign a1fe5e = hmaster0_p & v23f4338 | !hmaster0_p & v23fc07c;
assign bb5cd7 = jx0_p & v22ff205 | !jx0_p & v22f97f5;
assign v23fb0a1 = hbusreq6 & v22f640a | !hbusreq6 & !v84561b;
assign v191afad = hgrant5_p & v2310a41 | !hgrant5_p & !v15071d8;
assign v2309729 = hgrant1_p & v22fb1bc | !hgrant1_p & v23f134a;
assign v22eb952 = hgrant3_p & v2309d7f | !hgrant3_p & v23139c3;
assign v23faa93 = jx1_p & c17811 | !jx1_p & v84561b;
assign v2305194 = hmaster2_p & v22eec6e | !hmaster2_p & v22ee8f3;
assign v23f4961 = hbusreq4_p & v22f0db9 | !hbusreq4_p & v22ebfd3;
assign v23fb7c8 = hbusreq6_p & v230af11 | !hbusreq6_p & v23fc4d4;
assign v23fbcd8 = hbusreq6_p & v2301565 | !hbusreq6_p & v23fc598;
assign v23f9fcf = hmaster2_p & v2310e40 | !hmaster2_p & v9b93b3;
assign v22eb3e5 = hmaster2_p & v23fc596 | !hmaster2_p & v845622;
assign v22faae8 = hbusreq3_p & v23fc30d | !hbusreq3_p & v23fb77d;
assign v22f9c42 = stateG10_5_p & v23fcccd | !stateG10_5_p & v230f63f;
assign v2303ce0 = jx1_p & v85e5cf | !jx1_p & !v23f1cc0;
assign v8a0e71 = stateG10_5_p & v997ca9 | !stateG10_5_p & v17a34ff;
assign v22fdf5b = hbusreq2 & v84562b | !hbusreq2 & v84561b;
assign v22f448b = hbusreq5 & v22eb5b3 | !hbusreq5 & v84561b;
assign v23fcc43 = hlock4_p & v231182b | !hlock4_p & v23fbad7;
assign v22f2bab = hmaster2_p & v22fef4f | !hmaster2_p & v191aa68;
assign v23fcc5f = hlock3_p & v23105eb | !hlock3_p & v2303d65;
assign v23fa3b6 = hbusreq3 & v22f60da | !hbusreq3 & v84561b;
assign v23117d2 = hbusreq6_p & v22ef292 | !hbusreq6_p & v23f55c5;
assign v23fcaeb = hbusreq1 & v22f15fd | !hbusreq1 & v84561b;
assign v23f8970 = hgrant5_p & v22facbb | !hgrant5_p & v230cb7a;
assign v23fa463 = hgrant1_p & v84561b | !hgrant1_p & v230d5aa;
assign v231156b = hmaster0_p & v84561b | !hmaster0_p & v22fe792;
assign v23fa2e7 = hbusreq2_p & v22ff92f | !hbusreq2_p & !v23056b1;
assign v22f532c = hmastlock_p & v230f0a1 | !hmastlock_p & !v84561b;
assign v22fe675 = hmaster2_p & v22f79fd | !hmaster2_p & v2310e10;
assign v23f37c8 = hbusreq3_p & v22f575a | !hbusreq3_p & v22f42a5;
assign v22f57e8 = hgrant1_p & v23fc572 | !hgrant1_p & !v2306b05;
assign v2313144 = hmaster2_p & v22fef20 | !hmaster2_p & v2310108;
assign v23103f4 = jx1_p & v2301b0c | !jx1_p & v84561b;
assign v22f1259 = hbusreq4_p & v22f2cd3 | !hbusreq4_p & !v23f5c2f;
assign v22f2957 = hlock5_p & bbc337 | !hlock5_p & !v84561b;
assign v22f8d6a = hbusreq1 & v23fb952 | !hbusreq1 & v84561b;
assign v23f6843 = hbusreq3 & v22fab7c | !hbusreq3 & v84561b;
assign v22fff6e = hlock5_p & v22eec02 | !hlock5_p & !v84561b;
assign v22f25c5 = hbusreq6_p & v230824c | !hbusreq6_p & v22febde;
assign v22f05a7 = hbusreq1_p & v2312142 | !hbusreq1_p & bd9e8b;
assign v23fccec = hbusreq1 & v23fb980 | !hbusreq1 & v97808c;
assign v22f035c = hbusreq1_p & v22ee44f | !hbusreq1_p & !v23031eb;
assign v2310da0 = hlock0_p & v23fbefa | !hlock0_p & v2306885;
assign v23fb18e = hmaster2_p & v23fcf46 | !hmaster2_p & !v23f5cb3;
assign da310c = hmaster0_p & v2300d0f | !hmaster0_p & v23fbf61;
assign v2392394 = hmaster1_p & v23f42ec | !hmaster1_p & v2303d9e;
assign v231171e = hmaster0_p & v23fce0b | !hmaster0_p & !v2308fe5;
assign v23f7f0d = hbusreq1_p & v23fb788 | !hbusreq1_p & v84561b;
assign a1fe27 = hlock0_p & v22fef4f | !hlock0_p & v2300032;
assign v2346b6a = hgrant1_p & v22f3738 | !hgrant1_p & v230c233;
assign v22f12cd = hgrant2_p & v22f2f04 | !hgrant2_p & v23fc383;
assign v23f534c = hbusreq6_p & v22f7347 | !hbusreq6_p & v22f62a9;
assign v22f6187 = hbusreq1_p & v23fce72 | !hbusreq1_p & v22fb155;
assign v22eddae = hbusreq4 & v22f16ef | !hbusreq4 & v230038a;
assign v23fab20 = hlock0_p & v23fbb84 | !hlock0_p & v23fb913;
assign v23f2a86 = hlock5_p & v23f3eed | !hlock5_p & v84561b;
assign v23fc102 = hbusreq1_p & v23083d6 | !hbusreq1_p & !v84561b;
assign a1fe3e = hgrant5_p & v23fc14d | !hgrant5_p & v23fbd00;
assign v23f240a = hmaster0_p & bd74ba | !hmaster0_p & v23fa0a3;
assign v22f7f91 = hbusreq5_p & v22ef4ce | !hbusreq5_p & v23045ac;
assign v23fc253 = stateG10_5_p & v22ecf87 | !stateG10_5_p & v22ee956;
assign v23f6325 = hbusreq4_p & v23fc22c | !hbusreq4_p & v230c3ee;
assign v23fcf5b = hmaster2_p & v191a86f | !hmaster2_p & v23fbca3;
assign v22f5f09 = hbusreq1_p & v23fc17b | !hbusreq1_p & v23f7796;
assign v23f3ce8 = hbusreq6 & v22fcf52 | !hbusreq6 & v22ee657;
assign v22f6058 = hgrant0_p & a1fba6 | !hgrant0_p & v1aadb95;
assign v2308b58 = hmaster0_p & v23fb8aa | !hmaster0_p & d49f2b;
assign v2312a93 = hbusreq4 & v23fbc6a | !hbusreq4 & aa26cc;
assign v2391a62 = hbusreq5_p & v23fcf91 | !hbusreq5_p & v22f0b45;
assign v23f35c7 = hbusreq3_p & v23fc30d | !hbusreq3_p & v22efc21;
assign v22fc212 = hmaster0_p & v2308815 | !hmaster0_p & a1fbc2;
assign v2303da9 = hmaster2_p & v8912cf | !hmaster2_p & !v23fc514;
assign v23fd016 = jx0_p & v230477b | !jx0_p & v22eab03;
assign v22effdc = hmaster1_p & v23f619d | !hmaster1_p & v22f7588;
assign v2303352 = hgrant2_p & v22ede4d | !hgrant2_p & v84561b;
assign b50bc7 = hgrant5_p & v23fc4b4 | !hgrant5_p & v23f529c;
assign v23040c8 = hbusreq3 & v230fe27 | !hbusreq3 & v84561b;
assign v23fc503 = stateG10_5_p & v230d1a6 | !stateG10_5_p & v23f6411;
assign v230882d = locked_p & v23fba3a | !locked_p & v191a879;
assign v23fc383 = hbusreq2_p & v230ace0 | !hbusreq2_p & !v84561b;
assign v23038dd = hbusreq3_p & v23fb8ec | !hbusreq3_p & v22fc374;
assign v231094e = hmaster0_p & v22f2e69 | !hmaster0_p & !v23f1803;
assign v23fbfe2 = hlock1_p & v22ed4c6 | !hlock1_p & v2308235;
assign v2300a04 = hmaster2_p & v23f1db4 | !hmaster2_p & v2300b76;
assign v23f673b = hlock4_p & v1aae99f | !hlock4_p & !v23040a8;
assign v23f5d39 = hmaster1_p & v22f01b6 | !hmaster1_p & v2308d60;
assign v2303061 = hbusreq3_p & v23fb18e | !hbusreq3_p & !v23f57c1;
assign v22eb742 = hgrant5_p & v23fc1bf | !hgrant5_p & v22fb4a1;
assign v2392d4f = hgrant5_p & v23fcd22 | !hgrant5_p & v23fc612;
assign v12cc72f = hgrant0_p & v22eaafd | !hgrant0_p & v2303b4f;
assign v23fca07 = hbusreq3 & b67ed5 | !hbusreq3 & v22eb895;
assign v230539c = jx1_p & v22f036f | !jx1_p & v22f803b;
assign v23fbb8a = stateG10_5_p & v23f4fa1 | !stateG10_5_p & !v23f8383;
assign v22fda49 = hbusreq0 & v23fba6b | !hbusreq0 & v84561b;
assign v2307743 = hbusreq0_p & v230f1a7 | !hbusreq0_p & v23fb1a6;
assign v230585c = hbusreq4_p & v2307081 | !hbusreq4_p & v23efb3a;
assign v23f6769 = hbusreq3 & v230f9c2 | !hbusreq3 & v84561b;
assign v22f5576 = hmaster2_p & v84564d | !hmaster2_p & v22ed85a;
assign v23fcf79 = hbusreq5_p & v8f2065 | !hbusreq5_p & v230bbe4;
assign v230e89f = hbusreq3 & v23fa1f9 | !hbusreq3 & v84561b;
assign v23f36f1 = hbusreq5_p & v191b0a2 | !hbusreq5_p & !v84561b;
assign v2301c2a = hmaster0_p & v2313266 | !hmaster0_p & v22f4f06;
assign v23fc4f5 = hbusreq5_p & fc8e3a | !hbusreq5_p & !v84561b;
assign v22f383b = hbusreq1_p & v9a6a67 | !hbusreq1_p & !v23fb561;
assign v22f9a6b = hbusreq4_p & v23fbab6 | !hbusreq4_p & v84561b;
assign v2313264 = hburst0 & v230177d | !hburst0 & !v84561b;
assign v230935d = hbusreq1_p & v23126ae | !hbusreq1_p & v106af73;
assign v22f0050 = hbusreq3_p & v230dd35 | !hbusreq3_p & v23934f3;
assign v23fbf59 = hbusreq1 & v2312cdf | !hbusreq1 & v84561b;
assign v23fbc1a = hbusreq3_p & v230d20f | !hbusreq3_p & v84561b;
assign v23fb078 = hbusreq4_p & v23109e3 | !hbusreq4_p & v23f232d;
assign v22f17eb = hbusreq2 & v1aadb8e | !hbusreq2 & v84561b;
assign v191ab12 = hmaster2_p & v23f4b28 | !hmaster2_p & v23fca2a;
assign v23fd038 = hmaster0_p & v230d667 | !hmaster0_p & !v96c563;
assign v22f7a60 = hbusreq4_p & v22fb5f1 | !hbusreq4_p & v230c616;
assign v23024b6 = hlock0_p & v23f450b | !hlock0_p & v22ee1e6;
assign v22f7d41 = hgrant2_p & v12cd523 | !hgrant2_p & !v230e71c;
assign v22fa05b = hmaster2_p & v23f4f1e | !hmaster2_p & v230b0f5;
assign v22ff134 = hbusreq4_p & v22ed145 | !hbusreq4_p & v84561b;
assign v22f9f67 = hmaster2_p & v106a782 | !hmaster2_p & !v2307c5d;
assign v23fcaea = hmaster0_p & v231363b | !hmaster0_p & v23fd00f;
assign v22fb30f = hmaster2_p & v22f61b6 | !hmaster2_p & v23112ad;
assign v230b0f5 = hgrant1_p & v84561b | !hgrant1_p & v230104e;
assign v230910b = hbusreq5_p & v2305338 | !hbusreq5_p & v84561b;
assign v23fd00f = hbusreq6 & v2311b20 | !hbusreq6 & v23065e7;
assign v23fbcff = hbusreq5_p & a1fba6 | !hbusreq5_p & v22fc835;
assign v23fa91a = hbusreq2 & v191a876 | !hbusreq2 & v84561b;
assign v22eb75e = hbusreq3_p & v22f1b23 | !hbusreq3_p & v84561b;
assign v230ae9d = hgrant3_p & v23139ef | !hgrant3_p & v230cdf2;
assign v230e6ba = hbusreq1 & v2300071 | !hbusreq1 & v84561b;
assign v23f797b = hgrant1_p & v84561b | !hgrant1_p & v23ef89d;
assign v22f8a7e = hbusreq3_p & v23facab | !hbusreq3_p & v84561b;
assign v23fc5dd = hlock3_p & v23027f9 | !hlock3_p & v22ed8c4;
assign v23fb906 = hgrant1_p & v12cd9f9 | !hgrant1_p & !v84561b;
assign v22fcceb = hbusreq0_p & v23f7218 | !hbusreq0_p & v23fb4d1;
assign v106a84c = hgrant6_p & v84561b | !hgrant6_p & v22f25ac;
assign v22ec658 = hlock2_p & v84564d | !hlock2_p & !v84561b;
assign v23055b3 = hbusreq5_p & v23126ae | !hbusreq5_p & v22fc7c1;
assign v23f95ef = stateG10_5_p & v22fa766 | !stateG10_5_p & v22ec801;
assign v23fce11 = hgrant5_p & v23fc74c | !hgrant5_p & v84561b;
assign a1fc74 = hbusreq1_p & v23fc355 | !hbusreq1_p & !v23f14e6;
assign v10dbf64 = busreq_p & v191a86f | !busreq_p & !v191a879;
assign v2305ebc = hgrant5_p & v2306e1a | !hgrant5_p & v22fa707;
assign v23fc8f0 = stateA1_p & v22f0362 | !stateA1_p & v2300edd;
assign v23faade = hmaster0_p & v22fcdd3 | !hmaster0_p & !v23fce88;
assign v23f53a0 = hbusreq3_p & v23f522c | !hbusreq3_p & v84561b;
assign v230945e = hbusreq1_p & v9526ac | !hbusreq1_p & v23f972e;
assign v230e9d1 = hgrant3_p & v2394087 | !hgrant3_p & b09263;
assign v230bead = hbusreq3_p & v2307704 | !hbusreq3_p & v23f200c;
assign v1aae6b5 = hmaster1_p & v230fca8 | !hmaster1_p & v2312f82;
assign v22f748c = hmaster0_p & v22f87a1 | !hmaster0_p & v8fafbf;
assign v99005c = hgrant4_p & a54167 | !hgrant4_p & v23fcf45;
assign v23fcd71 = hbusreq5_p & v23fb481 | !hbusreq5_p & v2307b4c;
assign v230e880 = jx1_p & v23094a1 | !jx1_p & v84561b;
assign v23fc365 = hmaster2_p & v106a782 | !hmaster2_p & !v230eb9b;
assign v22efa5e = hmaster2_p & v22fef20 | !hmaster2_p & v230dbc9;
assign v22eeb42 = stateG10_5_p & v23fcd29 | !stateG10_5_p & v191a876;
assign v23fbcd2 = hlock4_p & be86f6 | !hlock4_p & v23f47a1;
assign v230c4bb = hbusreq5_p & v23fb0e3 | !hbusreq5_p & v23fcee9;
assign v22f0331 = hlock3_p & v23fbc1a | !hlock3_p & v22f4ebc;
assign v23f5cd3 = hbusreq3_p & v22ff9d4 | !hbusreq3_p & v23fc04f;
assign v23f1328 = hgrant4_p & v84561b | !hgrant4_p & v230a571;
assign v23004f9 = start_p & v84561b | !start_p & !v23094c6;
assign v2306e6f = hmaster0_p & v23f3bc9 | !hmaster0_p & v22fa0d4;
assign b031da = hmaster2_p & v1aad815 | !hmaster2_p & !v84561b;
assign v2309550 = hgrant1_p & v22f0755 | !hgrant1_p & v22f5e57;
assign v23f4ca0 = hgrant0_p & v84561b | !hgrant0_p & v2391b49;
assign da30fb = hmaster2_p & v23fc4f8 | !hmaster2_p & !v2312259;
assign b425f1 = hbusreq1 & v231026b | !hbusreq1 & v84561b;
assign v23fc03f = hgrant1_p & v23f5c95 | !hgrant1_p & v23fd034;
assign v2301b38 = hmaster0_p & v84561b | !hmaster0_p & !v23fbe89;
assign v230322f = hlock3_p & v22f4a1f | !hlock3_p & v22f44cc;
assign v23f8017 = hgrant5_p & v22ec5e6 | !hgrant5_p & v22f7f91;
assign v230dd28 = hmaster2_p & v23fcc72 | !hmaster2_p & v845625;
assign v23f4cf7 = hbusreq5_p & v2310a35 | !hbusreq5_p & !v84561b;
assign v23fb912 = hgrant2_p & v23fb973 | !hgrant2_p & ac37a1;
assign v23fc127 = hbusreq5_p & v23fc904 | !hbusreq5_p & v230320e;
assign v230d814 = hgrant1_p & v230d64e | !hgrant1_p & v23fcf71;
assign v2391b52 = hbusreq4_p & v23072f3 | !hbusreq4_p & v230f03c;
assign v230cf1a = hgrant0_p & v23fbb20 | !hgrant0_p & v22fb8d3;
assign v22f85c2 = hmaster0_p & v23f99a0 | !hmaster0_p & v23039c8;
assign f4076d = decide_p & v2302ffc | !decide_p & v84565b;
assign v22fb6bf = hlock5_p & v2302b44 | !hlock5_p & !v84561b;
assign v23fca0f = hmaster2_p & v230cb9a | !hmaster2_p & v22f8bd0;
assign v230358b = hready & v22fa2de | !hready & v22f60c6;
assign v2310317 = hbusreq6_p & v23f0dd4 | !hbusreq6_p & v22f25e0;
assign v22fe939 = jx1_p & v22faf49 | !jx1_p & v84561b;
assign v22fc5ad = hgrant5_p & v23f5cfd | !hgrant5_p & v23fb993;
assign v8f4f78 = hbusreq5_p & v22f6e70 | !hbusreq5_p & v84561b;
assign v23f93ee = hbusreq1 & v2307b39 | !hbusreq1 & v84561b;
assign v22fb0b7 = hbusreq5_p & v22fc091 | !hbusreq5_p & v22f65d5;
assign v23f4268 = hbusreq5_p & v2301511 | !hbusreq5_p & v230c6eb;
assign v22fc481 = hmaster1_p & v22ed1c4 | !hmaster1_p & v22ff184;
assign fc9434 = hbusreq5_p & v230cc4c | !hbusreq5_p & v84561b;
assign v22ed878 = hready & v23fc4a4 | !hready & !v84561b;
assign v106af3a = hlock3_p & v2305b34 | !hlock3_p & !v84561b;
assign v23fbfb2 = hmaster0_p & v23fbd48 | !hmaster0_p & !v23fc279;
assign v22ec960 = jx0_p & v2302608 | !jx0_p & v22f04ff;
assign v23f5ce2 = hlock0_p & v84561b | !hlock0_p & v23fc513;
assign v2312cc9 = hmaster2_p & v23f08a4 | !hmaster2_p & !v84561b;
assign v2311928 = hmaster0_p & v22eaeaf | !hmaster0_p & v22f09c4;
assign v23017a9 = hmaster1_p & e1e72e | !hmaster1_p & v150716b;
assign v2312775 = hbusreq2_p & v2307750 | !hbusreq2_p & v84561b;
assign bd9c35 = hmaster2_p & v23f77e8 | !hmaster2_p & v22f79fd;
assign v22fd364 = hmaster0_p & v23f38b7 | !hmaster0_p & !v22ecb12;
assign v22f6db5 = jx0_p & v22fc964 | !jx0_p & v23fb6b9;
assign v22ec5e6 = hbusreq5_p & v23fc4a1 | !hbusreq5_p & v230411f;
assign v2312f1b = hbusreq3_p & v230da2f | !hbusreq3_p & v22f40ef;
assign v22f264f = hgrant2_p & v22f8959 | !hgrant2_p & v22fb7bc;
assign v22f7083 = jx1_p & v85e5cf | !jx1_p & v22f2ce7;
assign v23f5ede = hgrant3_p & v230d2d8 | !hgrant3_p & v23efcf8;
assign v22fb214 = jx1_p & v230bbaf | !jx1_p & v22fbd0e;
assign v22f6529 = hmaster2_p & v22f8aec | !hmaster2_p & v22f6b4c;
assign v23f80e9 = hgrant0_p & v2310904 | !hgrant0_p & v23fcb23;
assign v23f47ca = hbusreq5_p & v23126ae | !hbusreq5_p & v22eeb42;
assign v2301f52 = hbusreq5 & v1aae087 | !hbusreq5 & v84561b;
assign v230b1a3 = hbusreq6_p & v23f3958 | !hbusreq6_p & v22ef116;
assign v23f2810 = hbusreq6 & v23f1354 | !hbusreq6 & v23f91bc;
assign v230e167 = hlock5_p & v230e651 | !hlock5_p & !v23f4e8c;
assign v23fbfd4 = hbusreq3_p & v22ed805 | !hbusreq3_p & v84561b;
assign v2311dcb = hbusreq5 & v22ed6c5 | !hbusreq5 & v84564d;
assign v23fa6f1 = hbusreq1 & v22f3643 | !hbusreq1 & v845620;
assign v22f86fc = hgrant6_p & v22f7722 | !hgrant6_p & v23f9c66;
assign v22fa768 = hbusreq6 & v22f5753 | !hbusreq6 & v84561b;
assign v23f39d9 = hmaster1_p & v230dd17 | !hmaster1_p & v1aad420;
assign v23fcf98 = stateG10_5_p & v23fd06a | !stateG10_5_p & v12cd4c6;
assign v230e7e3 = hbusreq5_p & v23fcf46 | !hbusreq5_p & v23fc7a4;
assign v22f0126 = hbusreq1_p & da38c1 | !hbusreq1_p & v230a22e;
assign v2309cdc = hbusreq1_p & v23fc361 | !hbusreq1_p & v84561b;
assign v230a24c = hmaster2_p & v22fae6e | !hmaster2_p & !v22fa870;
assign v22ffaef = hmaster2_p & v84561b | !hmaster2_p & !b8a8d7;
assign v22fd679 = hready_p & v22ed287 | !hready_p & e1e78b;
assign v22fcc32 = hbusreq1_p & v23fcd9e | !hbusreq1_p & v23fb44f;
assign v22f9ab1 = hbusreq6 & v22fcc05 | !hbusreq6 & v2301073;
assign c16bc3 = hbusreq0_p & v22ff8ea | !hbusreq0_p & !v845629;
assign v22ffa07 = jx1_p & v23fbe7d | !jx1_p & v84561b;
assign v2303b76 = hlock0_p & v2303376 | !hlock0_p & v22f931f;
assign f40cd3 = hlock2_p & b6f86d | !hlock2_p & v845620;
assign v23fc0f8 = hbusreq3_p & v2309eab | !hbusreq3_p & v23fcd8a;
assign v23f72e4 = hgrant3_p & v22feec8 | !hgrant3_p & v22eaee8;
assign v22fc0ec = hbusreq4_p & v2392898 | !hbusreq4_p & !v22fe08f;
assign v2304ec7 = locked_p & v22fe9e0 | !locked_p & v84561b;
assign v23070c0 = hmaster2_p & v230665f | !hmaster2_p & v845627;
assign v23fcb44 = hgrant5_p & v84561b | !hgrant5_p & v23030e8;
assign v2391c58 = hbusreq2 & v23fc5d5 | !hbusreq2 & v84561b;
assign v23fc457 = hlock3_p & v23f06ee | !hlock3_p & !v84561b;
assign v22f5ca6 = stateG10_5_p & v22eb5cc | !stateG10_5_p & v23fcb69;
assign v23fbab6 = hlock4_p & v86d5f2 | !hlock4_p & v84561b;
assign v22f4e94 = hgrant1_p & v84561b | !hgrant1_p & v2306c16;
assign v23fd021 = hbusreq2_p & v22ee9c4 | !hbusreq2_p & v23f4963;
assign v22ee772 = hbusreq1_p & v845620 | !hbusreq1_p & v22f79fd;
assign v23f5398 = hmaster2_p & v23fb9a9 | !hmaster2_p & v230590b;
assign v23060eb = hbusreq1 & v230913d | !hbusreq1 & !v23088b3;
assign v22ebccb = busreq_p & v22ee516 | !busreq_p & !v23fc0f5;
assign v23f84b5 = hgrant2_p & v22f2f87 | !hgrant2_p & !v84561b;
assign v23fc0ab = hmaster2_p & v22f954f | !hmaster2_p & v23f1bbf;
assign v23f707f = stateG2_p & v22f7176 | !stateG2_p & v22f2958;
assign v22eb895 = hmaster2_p & v2313247 | !hmaster2_p & v22f7808;
assign v23fbb94 = hbusreq3_p & v22efd33 | !hbusreq3_p & v84561b;
assign v22fb5a3 = hgrant5_p & v2393f08 | !hgrant5_p & v2300881;
assign v2311dc5 = hgrant3_p & v22efdf3 | !hgrant3_p & v23fc850;
assign v230c0dd = hmaster0_p & v22f654f | !hmaster0_p & v22ec77a;
assign v2300b76 = hbusreq1_p & v2301d23 | !hbusreq1_p & v22f878c;
assign v23003f5 = hbusreq4 & v23f9fa4 | !hbusreq4 & v22f5583;
assign v230936c = hmaster0_p & b00aa6 | !hmaster0_p & v2312be1;
assign v22f88aa = hbusreq2 & v2309945 | !hbusreq2 & v84561b;
assign v23027e9 = hbusreq2_p & v23f63b2 | !hbusreq2_p & !v23f8914;
assign v23fcc21 = hbusreq3_p & v230ac22 | !hbusreq3_p & !v84562e;
assign b5e222 = hbusreq5_p & v845636 | !hbusreq5_p & e1e1cb;
assign v22eeece = hmaster2_p & v84561b | !hmaster2_p & v23f87f4;
assign v22fcf35 = hmaster1_p & v23fc76e | !hmaster1_p & !v23f49cd;
assign v22ee8ee = hbusreq6_p & v23fc8f3 | !hbusreq6_p & v22f4f0f;
assign v2309b3c = hbusreq5 & v22f4e0b | !hbusreq5 & v230f5a3;
assign v22f9b67 = hmaster0_p & v22f56a5 | !hmaster0_p & !v23008f3;
assign v22fc689 = hbusreq4_p & v22fd67c | !hbusreq4_p & v22fb43e;
assign v22f2d2a = hbusreq3 & v22fe5f9 | !hbusreq3 & v23f87f4;
assign v22ff67c = hmaster2_p & v23fc4f8 | !hmaster2_p & v84561b;
assign v23fb843 = hbusreq6_p & v22ef094 | !hbusreq6_p & v84561b;
assign v23003b8 = hlock0_p & v106af4d | !hlock0_p & v2300338;
assign v230b364 = stateA1_p & v22f3294 | !stateA1_p & v23f9904;
assign v23f8a43 = hbusreq4 & v23049d7 | !hbusreq4 & v22f5fb4;
assign v23f084d = hbusreq0_p & v106ae4a | !hbusreq0_p & v230beb6;
assign v22f24f8 = hbusreq1_p & v23f8986 | !hbusreq1_p & !v84561b;
assign v2307c06 = jx1_p & v23fc9f2 | !jx1_p & v23f5109;
assign v2306d22 = hmaster2_p & v1b87673 | !hmaster2_p & v23fcba7;
assign bbc337 = hbusreq5 & v84564d | !hbusreq5 & v84561b;
assign v23fc1ef = hgrant3_p & v84561b | !hgrant3_p & v22f0fe4;
assign v23055d4 = stateA1_p & v22f80ca | !stateA1_p & v230177d;
assign v230ff8a = hgrant4_p & v1aad671 | !hgrant4_p & v23fce4d;
assign v23f651e = hmaster1_p & v23fc755 | !hmaster1_p & v23fbb0c;
assign v22fe362 = hmaster0_p & v22ebc25 | !hmaster0_p & v23fcc90;
assign v22f1d92 = hbusreq5_p & v23faaa7 | !hbusreq5_p & !v84561b;
assign v2312e4e = hmaster2_p & v191a86f | !hmaster2_p & v2392d6d;
assign v22fc2c1 = hmaster0_p & v22eef3f | !hmaster0_p & v23f1225;
assign v23fc841 = hmaster0_p & v23fbc7e | !hmaster0_p & v22fcd06;
assign v22f6d58 = hgrant5_p & v23f6130 | !hgrant5_p & v23fbc42;
assign v23f66fd = hbusreq6_p & v2301818 | !hbusreq6_p & v84561b;
assign v22f8acf = hbusreq0_p & v22fc122 | !hbusreq0_p & v23fc2ee;
assign v2305a14 = hbusreq6_p & v230f1d6 | !hbusreq6_p & v2301dad;
assign v22fba10 = hmaster0_p & v22f368e | !hmaster0_p & v22f7070;
assign v22feac9 = hmaster2_p & v230f34c | !hmaster2_p & !v84561b;
assign v230fc64 = hbusreq3_p & a9c602 | !hbusreq3_p & v23efa84;
assign v95ca80 = hgrant3_p & v22f95c3 | !hgrant3_p & v23119e3;
assign v23fcdef = hbusreq4_p & v22fb9ad | !hbusreq4_p & v23f9e84;
assign v2303a2d = jx1_p & v23fc6a6 | !jx1_p & v22fccf0;
assign v22fd693 = jx1_p & v22edbc3 | !jx1_p & v22ec2e9;
assign v23fb22d = hmaster2_p & v23fb71a | !hmaster2_p & v2367a45;
assign v22fc95b = hbusreq3_p & v2311cd1 | !hbusreq3_p & v22f4114;
assign v23fcd29 = hgrant0_p & v2312a23 | !hgrant0_p & v23f2553;
assign v23070d5 = hbusreq3_p & v22fcfed | !hbusreq3_p & v23fb84b;
assign v22fe869 = hgrant3_p & v23f4cc5 | !hgrant3_p & v1aad31a;
assign v23f6a76 = hbusreq1_p & v230e4ae | !hbusreq1_p & v2304ee5;
assign v23fbf48 = jx0_p & v230cc50 | !jx0_p & v22f8499;
assign v22ecab2 = jx0_p & v23fcb03 | !jx0_p & v23fc70f;
assign v23fba3a = stateG2_p & v2302ca3 | !stateG2_p & v22f8db2;
assign v23f710b = hgrant3_p & v84561b | !hgrant3_p & v23fa3c0;
assign v22f42a5 = hbusreq3 & v12cda11 | !hbusreq3 & v845627;
assign v2313059 = hgrant1_p & v22ecd97 | !hgrant1_p & v23f8a0e;
assign v23fb8be = hgrant1_p & v22f3ed0 | !hgrant1_p & v23fc2c8;
assign v230a3f5 = hbusreq3 & v22f779f | !hbusreq3 & v8c2b38;
assign v2391b34 = hmaster1_p & v22ed7a4 | !hmaster1_p & v23f1206;
assign v2301818 = hlock6_p & v22f856d | !hlock6_p & v22fdbdb;
assign v22fc5a9 = hbusreq6 & v230f795 | !hbusreq6 & v23fb0bb;
assign v23fcbd7 = hgrant1_p & v84561b | !hgrant1_p & v23f5156;
assign v23fba9a = hgrant1_p & v845626 | !hgrant1_p & v22f7241;
assign d7db8a = hmastlock_p & v2309099 | !hmastlock_p & v84561b;
assign v23fbeb2 = hlock3_p & v23fc261 | !hlock3_p & v23fbe7f;
assign v23f3ca5 = hlock0_p & v84561b | !hlock0_p & v23f4d54;
assign v2308a0c = hlock5_p & v230dffa | !hlock5_p & v845620;
assign ae7427 = hbusreq1_p & v2309fdb | !hbusreq1_p & v84561b;
assign v23fc976 = hbusreq0 & v2308e63 | !hbusreq0 & !v84561b;
assign v230ed3d = hgrant3_p & v230fa21 | !hgrant3_p & v23fcaff;
assign v23f869a = hgrant3_p & v84561b | !hgrant3_p & v230c404;
assign v23fc432 = hlock1_p & e1df2d | !hlock1_p & v84561b;
assign v23f07eb = hlock6_p & v84561b | !hlock6_p & v191acb4;
assign v23f8db0 = hmaster0_p & v23fccdb | !hmaster0_p & !v2302e43;
assign v22f277f = hgrant0_p & v23f2b0b | !hgrant0_p & v22f6d06;
assign v23007b3 = hbusreq0_p & v22fe421 | !hbusreq0_p & v22fc8c8;
assign v22f8e9a = hgrant1_p & v12cc2ef | !hgrant1_p & v22fb2b4;
assign v2312d33 = hmaster0_p & v23f1e38 | !hmaster0_p & v230bff5;
assign v22fec20 = hbusreq3 & v23fcd09 | !hbusreq3 & v12cdba9;
assign v22ed6e1 = hmaster2_p & v191a879 | !hmaster2_p & !v2309871;
assign v23f957b = jx1_p & v23f96d1 | !jx1_p & v23fbe03;
assign v22f8c70 = hbusreq5_p & v1aae56f | !hbusreq5_p & v13affaa;
assign v22f07ac = hlock4_p & v2311f99 | !hlock4_p & v84561b;
assign v22f568c = hbusreq6_p & v1aaddcb | !hbusreq6_p & v22f1971;
assign v23fc505 = hmaster0_p & v23fc57e | !hmaster0_p & v23fbb8f;
assign v230d346 = hgrant0_p & v2309b0f | !hgrant0_p & b9888a;
assign v22fb891 = stateG10_5_p & v22fa20a | !stateG10_5_p & a1fba6;
assign v23f15af = hgrant5_p & v23fba17 | !hgrant5_p & v23f8176;
assign f40d9e = hbusreq5_p & v23121b5 | !hbusreq5_p & v84561b;
assign v22fdf3c = hmaster0_p & v1aae22e | !hmaster0_p & v22f92a2;
assign v861565 = hmaster2_p & v23fba6b | !hmaster2_p & !v23046f7;
assign v23fbd8a = hbusreq6 & v23f1c9b | !hbusreq6 & v22f2ca2;
assign v23f47d5 = stateG10_5_p & v22f5fb8 | !stateG10_5_p & !v23f908f;
assign v23fb581 = hready & v22f5eee | !hready & v230c899;
assign v22f2254 = hmaster2_p & v22feb47 | !hmaster2_p & v22f79fd;
assign v2303822 = hmaster0_p & v22f1963 | !hmaster0_p & v22f971f;
assign v2308ced = hmaster0_p & v230d96b | !hmaster0_p & !v230ab72;
assign v23fc732 = hgrant0_p & v22f2c30 | !hgrant0_p & v23f7218;
assign v23fbd00 = hbusreq5_p & v2393c3a | !hbusreq5_p & v23f4eb4;
assign v23fc1c7 = stateG2_p & v84561b | !stateG2_p & v230b364;
assign v23fc4a3 = hgrant1_p & v23f11a3 | !hgrant1_p & v23fc117;
assign v22eaf2a = hmaster0_p & v22ed711 | !hmaster0_p & v22fdfde;
assign v23fc1c0 = hmaster0_p & v23fc23a | !hmaster0_p & v96c563;
assign v23f770f = hgrant5_p & v23fbada | !hgrant5_p & v23fb98f;
assign v23fce9d = hlock3_p & v9ce189 | !hlock3_p & !v84561b;
assign v23f5446 = hmaster0_p & v23f7e8f | !hmaster0_p & v22f10c8;
assign e1e73a = stateG10_5_p & v22feb95 | !stateG10_5_p & b5f51c;
assign v22fcd80 = hgrant3_p & v84561b | !hgrant3_p & !v230070e;
assign v230ba49 = jx1_p & v22f3a1f | !jx1_p & v22fad67;
assign v23f344d = hbusreq3 & v230ddf3 | !hbusreq3 & v23fbf1c;
assign v22f29e6 = hmaster0_p & v22f16ad | !hmaster0_p & v23110f1;
assign v23f38c4 = hmaster2_p & b16aac | !hmaster2_p & v2302225;
assign v22ff29f = hmaster0_p & v230741d | !hmaster0_p & v2305aa9;
assign v23fbe9a = stateG10_5_p & v22f3c3d | !stateG10_5_p & v845636;
assign v22fb403 = hbusreq5_p & v845636 | !hbusreq5_p & v2309b3a;
assign v23f3d02 = hlock3_p & v2312dd2 | !hlock3_p & !v84561b;
assign v22fc27d = hlock3_p & v22f1117 | !hlock3_p & a0de1c;
assign v23fba28 = hmaster0_p & v23f2810 | !hmaster0_p & v23fc1d3;
assign v230e2d8 = hbusreq1_p & v2300387 | !hbusreq1_p & v23fc3dd;
assign v22ed8b0 = hbusreq6_p & v22f6b4e | !hbusreq6_p & v22fbe9e;
assign v23fc7e2 = hmaster2_p & v22f954f | !hmaster2_p & v230e8a6;
assign v23f520c = hbusreq5_p & v23fc904 | !hbusreq5_p & !v23012e5;
assign v22f1393 = hgrant5_p & v22f05f3 | !hgrant5_p & v22eba12;
assign v22f7830 = hbusreq1_p & v23007a4 | !hbusreq1_p & !v2309c8a;
assign v23f4067 = stateG2_p & v84561b | !stateG2_p & !v23fbbf3;
assign v23fb70f = hmaster0_p & v22ffd0e | !hmaster0_p & !v22f9b75;
assign v22fba6d = hmaster2_p & v84561b | !hmaster2_p & v22f4e2e;
assign v22fdc37 = hmaster2_p & af6dff | !hmaster2_p & v23f79f6;
assign v23f4364 = hbusreq3 & v23fbcce | !hbusreq3 & v84561b;
assign v23fb954 = hgrant3_p & v22f0a24 | !hgrant3_p & v22fb49d;
assign v22ffb91 = hbusreq1 & v22f3fec | !hbusreq1 & v230466d;
assign v23fb4a5 = hbusreq4_p & v22f8f49 | !hbusreq4_p & v23fa6eb;
assign v23f9cc4 = hlock6_p & ac10e3 | !hlock6_p & v22f4b2c;
assign v22f8eb8 = hgrant3_p & v2312cf9 | !hgrant3_p & v86df86;
assign v230437d = hmaster2_p & v22f3643 | !hmaster2_p & v23105cd;
assign v23fc4ca = hmaster2_p & v84561b | !hmaster2_p & v2300815;
assign v22f3834 = hbusreq1 & fc8ab7 | !hbusreq1 & !v84561b;
assign v22facd1 = hbusreq1_p & v22f7efd | !hbusreq1_p & v23fab9b;
assign v23fc58a = hmaster2_p & v84561b | !hmaster2_p & v230658d;
assign v230b282 = hgrant1_p & v84561b | !hgrant1_p & !v23f3051;
assign v2307cdf = hmaster0_p & v1b8771f | !hmaster0_p & v22f58cd;
assign v23f66db = hlock4_p & v22ec978 | !hlock4_p & v2309bab;
assign v22f831d = hbusreq6_p & v22f9ca3 | !hbusreq6_p & bd7669;
assign v23fcf38 = hmaster2_p & v23f8928 | !hmaster2_p & v239342f;
assign v22f6719 = hbusreq3 & v23f8561 | !hbusreq3 & v84561b;
assign v230381a = hmaster0_p & v23fc33e | !hmaster0_p & v84561b;
assign v23fbd03 = hbusreq5 & v23fc4f7 | !hbusreq5 & !v230828b;
assign v23fab26 = hbusreq3_p & v22f03b1 | !hbusreq3_p & v230aa63;
assign v22f2a24 = hbusreq0_p & v845622 | !hbusreq0_p & v23fbf80;
assign v22eb097 = hbusreq1_p & v22f866f | !hbusreq1_p & !v1507464;
assign v8a3511 = hlock1_p & v84561b | !hlock1_p & v84564d;
assign v22fa49d = hmaster0_p & v23121e0 | !hmaster0_p & v23fcdf0;
assign v23fc5ad = hbusreq4 & v23f1812 | !hbusreq4 & v22ede6c;
assign v23fc00b = hbusreq6 & v23fcaef | !hbusreq6 & v230dd28;
assign v23fcd9f = hgrant5_p & v230aba5 | !hgrant5_p & v191b1f3;
assign v2303e03 = hmaster2_p & v22f8c43 | !hmaster2_p & v1aae490;
assign v23fb9d4 = hgrant6_p & v845625 | !hgrant6_p & v2307d70;
assign v2301a6d = hmaster2_p & v84561b | !hmaster2_p & !v23f34d4;
assign v23fc816 = hbusreq6_p & v23fca6f | !hbusreq6_p & v230caac;
assign v23fcce3 = hlock0_p & v84561b | !hlock0_p & v845629;
assign v23f6d93 = stateG2_p & v84561b | !stateG2_p & v23fc331;
assign v12cd93a = hbusreq5 & v23fcb5e | !hbusreq5 & v84561b;
assign v23faa23 = hbusreq1 & v2304ee5 | !hbusreq1 & v84561b;
assign v230bf51 = hmaster2_p & v23fc4d3 | !hmaster2_p & b7ab40;
assign v23fc24a = hbusreq5_p & v23fca2a | !hbusreq5_p & v22f877e;
assign v22f4fb2 = hbusreq3 & v22f5b18 | !hbusreq3 & v23007f9;
assign v23fb8f7 = jx2_p & v23fd018 | !jx2_p & v2307e41;
assign v23010b3 = hbusreq3_p & v22fc508 | !hbusreq3_p & v231051e;
assign v23fb17e = hbusreq3_p & v23fbb39 | !hbusreq3_p & !v23fa2eb;
assign fc8c3f = hgrant1_p & v231128c | !hgrant1_p & v22f214f;
assign v1aae490 = hgrant1_p & v2313965 | !hgrant1_p & v191afad;
assign a1fd0e = hbusreq6 & v23fc8a6 | !hbusreq6 & v22f0a22;
assign v22f5a6c = hbusreq5_p & v23f908f | !hbusreq5_p & !v2312343;
assign v230754a = jx2_p & bfba4f | !jx2_p & v11853ca;
assign v230c3f5 = hmaster2_p & e1e7b0 | !hmaster2_p & v84561b;
assign v23fcd2d = hbusreq5_p & v23fcc31 | !hbusreq5_p & v84564d;
assign v23f2a3d = locked_p & v84561b | !locked_p & !v23fbb74;
assign v23fbdf9 = hgrant3_p & v22f8839 | !hgrant3_p & v12cd3e7;
assign v23fc7c8 = hmaster2_p & v22f0945 | !hmaster2_p & b60876;
assign v22f533e = hgrant0_p & v23fcf46 | !hgrant0_p & v230e2f9;
assign v23fb84a = hbusreq3_p & v23fcfd3 | !hbusreq3_p & v23f8345;
assign v22f7722 = hmaster1_p & v8fac11 | !hmaster1_p & v84561b;
assign v22ff6c5 = hmaster2_p & v23f6653 | !hmaster2_p & v1506fa4;
assign v23934f0 = hgrant1_p & v9b93b3 | !hgrant1_p & v22f1a04;
assign v22eed4c = hbusreq0 & v22fc34e | !hbusreq0 & v84561b;
assign v23fb710 = hbusreq5 & v2302e32 | !hbusreq5 & v84561b;
assign v23fb786 = hbusreq5 & v22f9911 | !hbusreq5 & v84561b;
assign v22eb8b6 = hbusreq5 & v23fc7b2 | !hbusreq5 & v22ff090;
assign v22f3f06 = locked_p & v106ae4a | !locked_p & a1fba6;
assign v22f8214 = hbusreq2 & v22fdaa1 | !hbusreq2 & v84561b;
assign v22f91f1 = hgrant3_p & v84561b | !hgrant3_p & v22f595b;
assign v23fb159 = hbusreq5_p & v17a34ff | !hbusreq5_p & !bd7c53;
assign v23fb6ff = hbusreq1_p & v23fb4cb | !hbusreq1_p & !v84561b;
assign v22f03b8 = hgrant2_p & v84562a | !hgrant2_p & !v23f5f07;
assign v22f5cf0 = hmaster2_p & v22f17bb | !hmaster2_p & v230a671;
assign v2308a7d = hbusreq3_p & v22f5828 | !hbusreq3_p & !v84561b;
assign v23fb71a = hbusreq1_p & v230665f | !hbusreq1_p & !v84561b;
assign v23fcfa1 = hbusreq4_p & v230e97b | !hbusreq4_p & v2310538;
assign v22eeef8 = hmaster2_p & v84561b | !hmaster2_p & v22ed035;
assign v23fc279 = hgrant3_p & v23105b1 | !hgrant3_p & v22f2ffc;
assign v22f525a = hmaster0_p & v23fc761 | !hmaster0_p & v22ffe30;
assign v231258e = hbusreq1_p & v22fd271 | !hbusreq1_p & v230b3a5;
assign a1fd46 = hbusreq1_p & v23fc127 | !hbusreq1_p & !v23fbca3;
assign v230e932 = hmaster2_p & v23f5cb3 | !hmaster2_p & !v23fc904;
assign v23fc3aa = hbusreq3_p & v22ec354 | !hbusreq3_p & v23fb7c3;
assign v23067c1 = hbusreq5_p & v84562a | !hbusreq5_p & v230828b;
assign v230fca8 = hbusreq6_p & v23f62f2 | !hbusreq6_p & v23fbc9e;
assign v23039af = hbusreq4_p & v22ec20e | !hbusreq4_p & v84561b;
assign v2312999 = hmaster2_p & v84561b | !hmaster2_p & e1dd71;
assign v23fc99e = hbusreq6 & v23fb8f1 | !hbusreq6 & v84561b;
assign v23fcafc = hmaster0_p & v23130de | !hmaster0_p & !v84561b;
assign v23fcbb5 = hbusreq2_p & v2306d29 | !hbusreq2_p & !v191a86f;
assign v23fb9b6 = hbusreq6 & v2313077 | !hbusreq6 & !v2303db8;
assign v230e991 = hmaster1_p & v231242a | !hmaster1_p & v2308a60;
assign v230bc39 = hmaster2_p & v23fcf77 | !hmaster2_p & !v23f87f4;
assign v1aad354 = hlock6_p & fc8f90 | !hlock6_p & v845623;
assign v23067ba = stateG10_5_p & v2308356 | !stateG10_5_p & v22eb5b3;
assign v230aa99 = hlock3_p & v230e869 | !hlock3_p & v2304bc1;
assign v2304598 = hmaster0_p & v22fb335 | !hmaster0_p & v2302cf5;
assign v230c132 = hbusreq3 & e1e1d4 | !hbusreq3 & v23f7066;
assign v845653 = hgrant2_p & v84561b | !hgrant2_p & !v84561b;
assign v23fc585 = hmaster2_p & v84561b | !hmaster2_p & v22f05a7;
assign v23fc1d1 = hbusreq4_p & v22f41c4 | !hbusreq4_p & v90eab4;
assign v22fafe5 = hlock1_p & v22eea17 | !hlock1_p & v845620;
assign v22eef92 = hbusreq3_p & v23fcb3c | !hbusreq3_p & v23fcf7a;
assign v22fcc89 = hgrant3_p & v22f31b9 | !hgrant3_p & v23078ff;
assign v22fede1 = hlock0_p & v22fe59a | !hlock0_p & !v84561b;
assign v230a534 = hbusreq6_p & v23f9cc4 | !hbusreq6_p & v84561b;
assign v23f296d = hbusreq5 & v22f5037 | !hbusreq5 & v22f9927;
assign v23109fb = hgrant1_p & v230879e | !hgrant1_p & v84561b;
assign v23108a7 = hbusreq1_p & v84561b | !hbusreq1_p & v23f7796;
assign v23fb52e = stateG10_5_p & v23f8a9d | !stateG10_5_p & v22f35fa;
assign v9180fe = hmaster2_p & v84561b | !hmaster2_p & v22f35fa;
assign v23064ad = hgrant3_p & v22f5d73 | !hgrant3_p & v230c872;
assign v22f1dc9 = hgrant3_p & v84562e | !hgrant3_p & v23fc953;
assign v8c2b38 = hmaster2_p & v84561b | !hmaster2_p & fc8ab7;
assign v23f1643 = hlock3_p & v22efdae | !hlock3_p & v23fc80d;
assign v23fbb7f = hbusreq2 & v2342fc3 | !hbusreq2 & !v84561b;
assign v22eb563 = hmaster2_p & v23f972e | !hmaster2_p & v22ff732;
assign v23f82b3 = hbusreq6 & v230ab2e | !hbusreq6 & v84562f;
assign v2308d66 = hbusreq0_p & v23f7218 | !hbusreq0_p & v2303b4f;
assign v23fbc17 = hbusreq0_p & v22f56d2 | !hbusreq0_p & v230f63f;
assign v23fc528 = hgrant3_p & v84561b | !hgrant3_p & v2304477;
assign v23f1b3d = hlock0_p & v23fc6ac | !hlock0_p & v23f6f5c;
assign v22efa67 = hbusreq5_p & v230b8cd | !hbusreq5_p & v23fcf2d;
assign v22fea77 = hbusreq4_p & v22f21d0 | !hbusreq4_p & v22eddc0;
assign v23134a0 = stateG10_5_p & v23fb861 | !stateG10_5_p & !a1fba6;
assign v230892a = hbusreq6_p & v22ffcae | !hbusreq6_p & !v84561b;
assign v22f6463 = hbusreq4_p & v2308abb | !hbusreq4_p & v84561b;
assign v2308ecc = hmaster2_p & v84561b | !hmaster2_p & !v23f16fd;
assign v23f8ca4 = hgrant1_p & v22fef02 | !hgrant1_p & v23f6c41;
assign v231125d = hmaster2_p & b9d013 | !hmaster2_p & !v23026c8;
assign v23f87be = hgrant3_p & v22fe551 | !hgrant3_p & v23fc5b4;
assign af5f08 = hmaster0_p & v23fced1 | !hmaster0_p & !v23fc624;
assign v23f9d5f = hbusreq5_p & v84561b | !hbusreq5_p & !v23fb4a8;
assign v23fcdda = hlock6_p & v23f85b0 | !hlock6_p & v2309a1d;
assign v22fe22b = hmaster2_p & v8be441 | !hmaster2_p & !a39dae;
assign v23f7eaa = hbusreq1 & v22fc34e | !hbusreq1 & v84561b;
assign v22ffd22 = hbusreq0_p & v22eed66 | !hbusreq0_p & v22f94a7;
assign v23fb94a = hmaster1_p & v2310db9 | !hmaster1_p & !v23f49cd;
assign v2307061 = hmaster2_p & v23fc5a9 | !hmaster2_p & v2300aab;
assign v22f2cd3 = hlock4_p & v23008a1 | !hlock4_p & !v23f5c2f;
assign v22f62ae = hgrant1_p & v84561b | !hgrant1_p & v23fc3ee;
assign v23f87e4 = jx1_p & v1507246 | !jx1_p & v22fbc04;
assign v23f15ec = hlock5_p & v2392bc1 | !hlock5_p & v2306c80;
assign v22faef4 = hbusreq3_p & v22fcfed | !hbusreq3_p & v23fc114;
assign adc67b = hmaster2_p & v22ebedd | !hmaster2_p & !v2302693;
assign v2310fde = hbusreq2_p & v84561b | !hbusreq2_p & !v845620;
assign v1aad517 = hbusreq6_p & v230144a | !hbusreq6_p & v1aae1de;
assign v23fcf96 = hlock0_p & v84561b | !hlock0_p & v230158f;
assign v23f89fe = hgrant5_p & a1fe52 | !hgrant5_p & v22f277f;
assign v1b87690 = hbusreq5 & v23f1207 | !hbusreq5 & v845620;
assign v22f877e = stateG10_5_p & v230fa13 | !stateG10_5_p & !v23fc84b;
assign v23fbd9c = hmaster2_p & v22edaa4 | !hmaster2_p & v84561b;
assign v2300d2f = hbusreq1_p & v23f1a8d | !hbusreq1_p & v23fcb69;
assign v2304bd1 = hlock5_p & v22eb682 | !hlock5_p & v22f92b8;
assign v23fc754 = hbusreq6_p & v22f009f | !hbusreq6_p & v230385f;
assign v22f9db5 = hmaster2_p & v8912cf | !hmaster2_p & v84561b;
assign v2306d37 = hlock0_p & v106a782 | !hlock0_p & v23fc6d9;
assign v23f8e52 = hbusreq1 & v13afe3a | !hbusreq1 & !fc8ab7;
assign v22f6dfa = hbusreq3_p & v23fbe02 | !hbusreq3_p & !v22f68f1;
assign v2304fc6 = hmaster2_p & v23fcf89 | !hmaster2_p & v239342f;
assign v1506a9e = hbusreq0 & v84564d | !hbusreq0 & v23fa2ec;
assign v22f482a = hbusreq3_p & v23f5e8a | !hbusreq3_p & v2300617;
assign da3103 = hbusreq6 & v230fc36 | !hbusreq6 & v23fd015;
assign v2304cc3 = hlock0_p & b09503 | !hlock0_p & da38b9;
assign v23fc828 = hlock5_p & v84561b | !hlock5_p & v22ff8a6;
assign v22f03ce = hgrant2_p & v22f4594 | !hgrant2_p & v22f925b;
assign v1aae22e = hbusreq4 & v23f67e2 | !hbusreq4 & v23fa2ec;
assign v230f776 = busreq_p & v22f4cca | !busreq_p & v23fb4a6;
assign v22ecb28 = hbusreq3_p & v23fc23b | !hbusreq3_p & v22faf4e;
assign v231003e = hgrant3_p & v84561b | !hgrant3_p & v23fbe0e;
assign v2302520 = hbusreq5_p & v23fab2c | !hbusreq5_p & v23fc5c4;
assign v23f22f9 = stateG10_5_p & v23fcb5e | !stateG10_5_p & !v23fb1a4;
assign v1aae362 = hmastlock_p & v22f091e | !hmastlock_p & v84561b;
assign v230522a = hbusreq1_p & v23f910c | !hbusreq1_p & v23fc050;
assign v22ee247 = hlock0_p & v2391aa0 | !hlock0_p & v22f181c;
assign v23f3f73 = hmaster2_p & v22eb599 | !hmaster2_p & v22fabd2;
assign v23f06d7 = hbusreq3_p & v84562e | !hbusreq3_p & !v84561b;
assign v23f3f24 = hmaster2_p & v23fbc43 | !hmaster2_p & v22f1895;
assign v2306779 = hbusreq0_p & v2303b9a | !hbusreq0_p & !v106ae19;
assign v23f0dc7 = hbusreq6_p & v2308db0 | !hbusreq6_p & v23f3e68;
assign baf3e5 = hmaster2_p & v230aded | !hmaster2_p & v9526ac;
assign v230be96 = hmaster2_p & v22f8b01 | !hmaster2_p & v2309729;
assign v2312680 = hgrant3_p & v23fcb87 | !hgrant3_p & v22f0050;
assign v2393900 = hgrant0_p & v22ede4d | !hgrant0_p & v84561b;
assign v23fce3d = hbusreq0_p & da38c1 | !hbusreq0_p & v23058ba;
assign v23f8176 = hgrant0_p & v22ed7d1 | !hgrant0_p & v2308e3c;
assign v23fbe83 = hbusreq1_p & v84562b | !hbusreq1_p & v17a34f9;
assign v1e840fa = hmaster2_p & v84561b | !hmaster2_p & !v84564d;
assign v23fb4f0 = stateG10_5_p & v84561b | !stateG10_5_p & v23f32eb;
assign v23fbc07 = hgrant0_p & v84561b | !hgrant0_p & !v22f366a;
assign v22fb4a1 = hgrant0_p & v2306785 | !hgrant0_p & v2303535;
assign v22f28f7 = jx1_p & v230eae5 | !jx1_p & v23fc631;
assign a7e154 = jx0_p & v23047dd | !jx0_p & v22f01b7;
assign v230dde9 = hgrant5_p & v84561b | !hgrant5_p & !v23fc9b9;
assign v22f4727 = hbusreq1_p & v22f8387 | !hbusreq1_p & v231140d;
assign v23fcb80 = hmaster0_p & v23f537e | !hmaster0_p & !v2304856;
assign v22fe147 = hbusreq4_p & v23f3c84 | !hbusreq4_p & v23fc689;
assign v12cda51 = hmaster0_p & v2301be6 | !hmaster0_p & v22ed1b5;
assign v22f49ff = hgrant3_p & v23018b7 | !hgrant3_p & v23fc956;
assign v2301f5c = hbusreq3 & v23fb1a0 | !hbusreq3 & v23f7f02;
assign v23fc4eb = jx1_p & v23f651e | !jx1_p & v2306822;
assign v23028ef = jx1_p & v23fc763 | !jx1_p & v230e4c7;
assign v22f08be = hbusreq5_p & v13afa38 | !hbusreq5_p & v230f222;
assign v23fbc12 = locked_p & v2312be7 | !locked_p & !v2309c8a;
assign v23fc8a5 = hbusreq3 & v23fb0c0 | !hbusreq3 & v84561b;
assign v22fafaa = hlock2_p & v84561b | !hlock2_p & !v2391a57;
assign v15074eb = hbusreq1 & v23f8364 | !hbusreq1 & !v84561b;
assign v23f8124 = hmaster0_p & v23f350b | !hmaster0_p & abc0f5;
assign v230474b = hgrant0_p & v84561b | !hgrant0_p & v23f54ac;
assign v22eb303 = hgrant1_p & v22f3738 | !hgrant1_p & v23f9044;
assign v23057a4 = jx1_p & v23f8410 | !jx1_p & v23fb94a;
assign v22f2677 = hgrant3_p & v23fd00d | !hgrant3_p & v22f2805;
assign v23fc616 = hmaster0_p & v23fcab7 | !hmaster0_p & !v23fba96;
assign v23f9737 = hbusreq6 & v2305aa7 | !hbusreq6 & v84561b;
assign v23f3d91 = hbusreq4_p & v23fc621 | !hbusreq4_p & v22f29e6;
assign v23f7a92 = hbusreq6_p & v98151e | !hbusreq6_p & v23fc334;
assign v22fae03 = hmaster0_p & v22fe869 | !hmaster0_p & a1fdac;
assign v23f1cd5 = hbusreq2 & v23fbb74 | !hbusreq2 & v84561b;
assign v22f78ee = hbusreq5_p & v22fa70c | !hbusreq5_p & v23fc01e;
assign v2312a8d = hbusreq1_p & v906d1d | !hbusreq1_p & v22ebf17;
assign v22f389b = hgrant1_p & v84564d | !hgrant1_p & !v230ed8b;
assign v230de4d = hbusreq5 & v230358b | !hbusreq5 & v84561b;
assign v22edcce = hmaster1_p & v2310b4d | !hmaster1_p & v23fd00e;
assign v23fcc58 = hbusreq3 & v2304924 | !hbusreq3 & v84561b;
assign v22f8da3 = hbusreq1 & v22ed65e | !hbusreq1 & v84561b;
assign v23fcfb8 = hlock0_p & v23f87ea | !hlock0_p & v23f4b28;
assign v23fc8b2 = hmaster2_p & v22f9880 | !hmaster2_p & v23fb966;
assign v22fc56c = hmaster0_p & v22f7800 | !hmaster0_p & v238ab71;
assign v23f0c76 = hbusreq3 & v23fc607 | !hbusreq3 & v22f5583;
assign v2308d06 = hbusreq4_p & v23fc1f8 | !hbusreq4_p & v230ce72;
assign v2311a4a = hmaster2_p & v22f768b | !hmaster2_p & !v22f7879;
assign v23f273b = hmaster0_p & v1e840b4 | !hmaster0_p & v23f2837;
assign v23f1f6f = locked_p & v84561b | !locked_p & v23fbb74;
assign v22f39a5 = stateG10_5_p & v9f009f | !stateG10_5_p & !v22ec921;
assign v22fc5fd = hlock0_p & v2310104 | !hlock0_p & v84562b;
assign v2309ffa = hmaster0_p & v22f5b58 | !hmaster0_p & v2309270;
assign v23f74bc = hmaster2_p & v2309c93 | !hmaster2_p & v84561b;
assign v23fad13 = hbusreq4 & v23f4fa4 | !hbusreq4 & !v22ff914;
assign v2309023 = hlock5_p & v22f2f33 | !hlock5_p & v845620;
assign v23f427e = hbusreq4_p & v22f216d | !hbusreq4_p & v12cd63d;
assign v23fc28d = hmaster2_p & v84561b | !hmaster2_p & !v22f5696;
assign v23022f2 = hgrant0_p & v22f5605 | !hgrant0_p & !v23fc0ce;
assign v22fe1d9 = hbusreq5 & v2312f7e | !hbusreq5 & !v22f91c9;
assign v23104cf = hmaster0_p & v23f3bc9 | !hmaster0_p & !v23f87be;
assign v23efcfb = hgrant3_p & a7b623 | !hgrant3_p & v97f5b6;
assign v22ee946 = hmaster2_p & v23f5be9 | !hmaster2_p & v22fc8e5;
assign b208fd = hmaster0_p & v84561b | !hmaster0_p & v22ff0ce;
assign v23f1206 = hbusreq4_p & v2301e4f | !hbusreq4_p & v2309317;
assign v22f9b46 = hbusreq6 & v230fcf6 | !hbusreq6 & v84561b;
assign v22fc73a = hgrant3_p & v22fc9cb | !hgrant3_p & !v23fb1b7;
assign v23fbcfd = hlock3_p & v23070d5 | !hlock3_p & v23fb0b6;
assign v2301de9 = hbusreq3_p & v23084fa | !hbusreq3_p & v84561b;
assign b572e8 = hbusreq0 & v22fafe4 | !hbusreq0 & v84561b;
assign v22ef848 = hlock3_p & v2312cad | !hlock3_p & v84561b;
assign v23fc08f = hmaster1_p & v23f3f36 | !hmaster1_p & !v22fe147;
assign e1e358 = hgrant3_p & v23fbcaa | !hgrant3_p & v22f1e67;
assign v22fd2e8 = hmaster0_p & v22f7273 | !hmaster0_p & v22efa0f;
assign v23fbf35 = hmaster2_p & v23fbda1 | !hmaster2_p & v22f0218;
assign v23fcfcc = hgrant0_p & v84561b | !hgrant0_p & v22fa16d;
assign v2304928 = hmaster0_p & v23f67d3 | !hmaster0_p & v230dde6;
assign v23fd069 = hbusreq3_p & v23f7b86 | !hbusreq3_p & v9bbf5d;
assign v23f4d54 = hbusreq0_p & v84561b | !hbusreq0_p & v22f1389;
assign v9526ac = hmastlock_p & v22f7ca0 | !hmastlock_p & v84561b;
assign v23f4a02 = hmaster2_p & v23131e8 | !hmaster2_p & !v23027e9;
assign v230cfe2 = hburst0_p & v84561b | !hburst0_p & !v22f8fb2;
assign v23f3d47 = hbusreq1_p & v2306d29 | !hbusreq1_p & v106af73;
assign v23fbd1b = hbusreq6_p & v22eb6ca | !hbusreq6_p & v2309751;
assign v231155f = hbusreq0_p & a476c2 | !hbusreq0_p & bd5342;
assign v23f1a14 = hgrant3_p & v2302c88 | !hgrant3_p & v22f12fb;
assign v23f5dfd = hlock4_p & e1c7f2 | !hlock4_p & !v2311ed2;
assign v23fcae1 = hbusreq4_p & v23f52f2 | !hbusreq4_p & v22f580c;
assign v23f089b = hmaster2_p & v845625 | !hmaster2_p & v23fcc72;
assign v22f23e6 = jx1_p & v22fcb9d | !jx1_p & v2392867;
assign v230ea67 = jx0_p & v22ffc83 | !jx0_p & v22fe116;
assign v230edc0 = hbusreq6_p & v23fc142 | !hbusreq6_p & v23fcc8f;
assign v23fc004 = stateG10_5_p & v23fcccf | !stateG10_5_p & v191a879;
assign v22eef1f = hmaster0_p & v22fda61 | !hmaster0_p & v230b8fe;
assign v23f5ed5 = hlock0_p & v84561b | !hlock0_p & v2305628;
assign v230cef0 = hgrant5_p & v22f5836 | !hgrant5_p & v23fc36e;
assign v1aae9e1 = hbusreq6_p & v2309b67 | !hbusreq6_p & !v84561b;
assign v23fb6c2 = stateG10_5_p & v2312336 | !stateG10_5_p & v23fc4f8;
assign v13afe3a = hmastlock_p & v22fab99 | !hmastlock_p & !v84561b;
assign v22f0a76 = hbusreq4_p & v2312a98 | !hbusreq4_p & v84561b;
assign v22f9160 = hmaster2_p & b50a75 | !hmaster2_p & !v84561b;
assign v230a9d5 = hgrant5_p & v23fceb0 | !hgrant5_p & v230d346;
assign v230e43d = hbusreq3_p & v84562b | !hbusreq3_p & v22fd696;
assign v23fbbf8 = hmaster2_p & v23fc1ce | !hmaster2_p & v23f53bd;
assign v230cfed = hgrant1_p & v2301e25 | !hgrant1_p & v23026ed;
assign v23f73af = hlock4_p & v23fcc2a | !hlock4_p & !v84561b;
assign v2311f82 = hbusreq6_p & v22ff4bc | !hbusreq6_p & v22f2487;
assign v22eda43 = hready & v22f5eee | !hready & !f4067f;
assign v22ee339 = hgrant1_p & v84561b | !hgrant1_p & v2310430;
assign v22fad67 = hbusreq6_p & v23f07eb | !hbusreq6_p & !v84561b;
assign v23f3d0e = hbusreq6 & v2312dd2 | !hbusreq6 & !v22ec6e5;
assign v2311072 = hbusreq2_p & v23fbb7f | !hbusreq2_p & !v84561b;
assign v23f6646 = hbusreq4 & v22fa1a2 | !hbusreq4 & v22f0492;
assign v22f4c34 = hbusreq3_p & v23f96aa | !hbusreq3_p & v23fc53b;
assign v22ee521 = hgrant3_p & v98d402 | !hgrant3_p & v23f4bc2;
assign v23f426b = hmaster2_p & v22f5d0e | !hmaster2_p & v23fcd00;
assign v22eec2d = hmaster1_p & v23efd8a | !hmaster1_p & v23061de;
assign v1aae19c = hbusreq1_p & v23fca96 | !hbusreq1_p & v22fd9eb;
assign v23fcbf0 = hbusreq6_p & v2309c79 | !hbusreq6_p & !v84561b;
assign v23f515d = hmaster0_p & v22f7c05 | !hmaster0_p & v23f3e1b;
assign v23fc6b3 = hbusreq5_p & v106a782 | !hbusreq5_p & v22f316f;
assign v23f35de = hbusreq4_p & v22ebf32 | !hbusreq4_p & v191b1ae;
assign v23fc230 = hmaster0_p & v23fc366 | !hmaster0_p & a1ba8b;
assign v23fb062 = hbusreq6_p & v23fcfa1 | !hbusreq6_p & v23fb622;
assign v23fbdfe = busreq_p & v230c041 | !busreq_p & v22ed5e6;
assign v23126c9 = hbusreq1_p & v22f792a | !hbusreq1_p & v845620;
assign v23063b0 = hbusreq6 & v22ffa4c | !hbusreq6 & v23f869a;
assign v230b9ad = hbusreq1_p & v22f74de | !hbusreq1_p & v22f409f;
assign v23fbf12 = hbusreq3_p & v22fc8e5 | !hbusreq3_p & v2309c93;
assign v2309e42 = hmaster0_p & v230c1dd | !hmaster0_p & v22f167b;
assign v22ef45e = hgrant5_p & v22f7c09 | !hgrant5_p & v2312fc7;
assign v23fbe6c = jx1_p & v23fbb81 | !jx1_p & v22f230d;
assign v230354e = stateG10_5_p & v22f1037 | !stateG10_5_p & v23fc393;
assign v22f7f3f = hbusreq6_p & v22f8c01 | !hbusreq6_p & bd8ac4;
assign v23fca96 = hbusreq1 & v22ebdbc | !hbusreq1 & v23fa2ec;
assign v22f5317 = hgrant3_p & v84561b | !hgrant3_p & v23039c0;
assign v22fabd2 = hbusreq1_p & v23f50ec | !hbusreq1_p & v84561b;
assign v22fa654 = hlock0_p & v23f340b | !hlock0_p & v230b7c1;
assign v22ff4c3 = hbusreq5_p & v8f2065 | !hbusreq5_p & v22ecec6;
assign v22fef65 = hmaster2_p & v23fa0bf | !hmaster2_p & v2310108;
assign v23f55c5 = hbusreq4_p & v22ef292 | !hbusreq4_p & v22ec1fc;
assign v23056b1 = locked_p & v22f5fa8 | !locked_p & v106ae19;
assign v2392537 = hbusreq3_p & e1dbd6 | !hbusreq3_p & v23056bf;
assign v23089fa = hbusreq3_p & v22f6870 | !hbusreq3_p & v1aad641;
assign v2391f4b = hbusreq1_p & v230db14 | !hbusreq1_p & v2308058;
assign v23fba4d = hgrant4_p & v230716d | !hgrant4_p & v22effdc;
assign v22f68c3 = hbusreq4_p & af5f08 | !hbusreq4_p & v23f1608;
assign v23fcdd9 = hgrant5_p & v2300621 | !hgrant5_p & v23f450d;
assign v23fca95 = hgrant3_p & v22f6124 | !hgrant3_p & v230a2ae;
assign v2301a67 = hgrant3_p & v22efc9e | !hgrant3_p & v23fc7e2;
assign v22f90d2 = hmaster2_p & v1aadb8e | !hmaster2_p & v23fcf96;
assign v2312196 = hlock3_p & b9c976 | !hlock3_p & v23f8caa;
assign v23fce46 = hgrant3_p & v23fab11 | !hgrant3_p & v23fc38f;
assign v230638a = hgrant3_p & v23fc7a6 | !hgrant3_p & v23fb8d1;
assign v2309cb5 = hbusreq2_p & v23022b1 | !hbusreq2_p & v22f91c9;
assign v22f9452 = hgrant1_p & v22ecd97 | !hgrant1_p & v230e6ea;
assign v22f8d2b = hbusreq0 & v2304009 | !hbusreq0 & v23fb966;
assign v2311d6b = hbusreq3_p & v23fcf21 | !hbusreq3_p & v22ee657;
assign v23fb97a = hlock3_p & v2307a49 | !hlock3_p & v23f149d;
assign v2311c65 = hmaster1_p & v23073e4 | !hmaster1_p & v23f8368;
assign v22ff308 = hgrant1_p & v845626 | !hgrant1_p & v23fc21a;
assign v23fba6c = hgrant3_p & v230bd1b | !hgrant3_p & v22fb842;
assign v23fc203 = hgrant1_p & v22f34bd | !hgrant1_p & v230bb21;
assign v22f56ce = hgrant3_p & v12cd9b6 | !hgrant3_p & v22fea74;
assign v23fc669 = hlock2_p & v2391a57 | !hlock2_p & v84561b;
assign v23f1354 = hbusreq3_p & v22f7be4 | !hbusreq3_p & v84561b;
assign v22ef862 = start_p & v84561b | !start_p & !v863ce5;
assign v22ecaef = stateG10_5_p & v23fc382 | !stateG10_5_p & v845636;
assign v22f7319 = hbusreq3 & c0084f | !hbusreq3 & v84561b;
assign v2303b4f = hgrant2_p & v23fc11e | !hgrant2_p & v230283f;
assign v23005a9 = hmaster2_p & v22f7808 | !hmaster2_p & v22f5815;
assign v23037d2 = hbusreq5_p & v22f2c2c | !hbusreq5_p & v22fb71d;
assign v23129bb = hbusreq5 & v23fb1a4 | !hbusreq5 & !v84561b;
assign v230eb8d = hgrant0_p & v845622 | !hgrant0_p & v23fbcc7;
assign v23fc632 = hgrant0_p & v84561b | !hgrant0_p & !v22fbd4b;
assign v23fc07e = hmaster2_p & a1fba6 | !hmaster2_p & v23fb875;
assign v230ea4c = hbusreq1 & v22feb6e | !hbusreq1 & !v22ee9ac;
assign v23f617e = hbusreq0 & v23f2be7 | !hbusreq0 & v84561b;
assign v23f2b14 = hbusreq1 & v22fc2bd | !hbusreq1 & v230a671;
assign v23fc823 = hbusreq1 & v2300c3d | !hbusreq1 & !v23f9fc1;
assign v22f5e09 = hready_p & v23f98d2 | !hready_p & !v230969a;
assign v22f674b = hbusreq4 & v23f1354 | !hbusreq4 & v23f91bc;
assign v2301aa7 = hbusreq2 & v22f9911 | !hbusreq2 & v84561b;
assign v23f15fe = locked_p & b9d00f | !locked_p & a1fba6;
assign v23fc0c9 = hbusreq5_p & v23f98f8 | !hbusreq5_p & v84561b;
assign v2303cc1 = hgrant1_p & v23fc856 | !hgrant1_p & v84561b;
assign v23fb0ea = stateA1_p & v23fc116 | !stateA1_p & !v84561b;
assign v22f5109 = stateG10_5_p & v230011a | !stateG10_5_p & v22f0945;
assign v23fa8bb = hgrant2_p & v230eb9b | !hgrant2_p & !v106a782;
assign v230f904 = hgrant3_p & v84561b | !hgrant3_p & v22f743b;
assign v2309440 = hgrant3_p & v22f118e | !hgrant3_p & !v22f07d5;
assign v23fcd09 = hmaster2_p & v2308d79 | !hmaster2_p & !v2312f7e;
assign a1fcc3 = hbusreq2 & v22eda36 | !hbusreq2 & v84561b;
assign v2306d29 = locked_p & v84561b | !locked_p & !v191a86f;
assign v191abee = hmaster2_p & a3cb61 | !hmaster2_p & v23f9b8d;
assign v23f7853 = hmaster2_p & v22f3f68 | !hmaster2_p & v23fc3f1;
assign v22eecf9 = hgrant0_p & v13afebe | !hgrant0_p & v23f3310;
assign v23fbfa7 = hgrant1_p & v84561b | !hgrant1_p & v23fb1e1;
assign v86374c = hgrant3_p & v22f2ca2 | !hgrant3_p & v22f2ac8;
assign v22f4a40 = hgrant3_p & v230a71c | !hgrant3_p & v2312948;
assign v230b199 = hlock3_p & v23fcd7a | !hlock3_p & v84561b;
assign v2310406 = hbusreq6_p & v23fbe05 | !hbusreq6_p & v23f81e6;
assign v2306997 = hgrant1_p & v84561b | !hgrant1_p & !v23fb8e7;
assign v22faa7c = hgrant3_p & v230d90f | !hgrant3_p & v22f0e6b;
assign v23fcd39 = hbusreq1 & v84561b | !hbusreq1 & v845620;
assign v2300c3d = hbusreq5_p & v22f60c6 | !hbusreq5_p & v84564d;
assign v22fc0a2 = hmaster0_p & v23f90b2 | !hmaster0_p & v23fc0b3;
assign v23fc944 = hbusreq6_p & v22f251d | !hbusreq6_p & v22fc2ca;
assign v23139b9 = hbusreq4_p & v2303b86 | !hbusreq4_p & v23fb08d;
assign v2305628 = hbusreq0_p & v23f4ab8 | !hbusreq0_p & v845629;
assign v22fcef4 = hlock4_p & v22ecf16 | !hlock4_p & v845637;
assign v22ee184 = hmaster2_p & v2392ece | !hmaster2_p & v22edc4f;
assign v23f936e = hbusreq3_p & v2302fbc | !hbusreq3_p & v84561b;
assign v2307fcd = hlock3_p & v2305a26 | !hlock3_p & v9c8a7f;
assign v22eb840 = hbusreq1_p & v2308d09 | !hbusreq1_p & !v23f55ea;
assign v2312142 = hlock1_p & v23938ff | !hlock1_p & bd9e8b;
assign v2312f82 = hbusreq4_p & v22fb2dc | !hbusreq4_p & v2311928;
assign v23fb973 = hbusreq2_p & v23fc91f | !hbusreq2_p & v845620;
assign v22f28e6 = hbusreq3_p & v22f4667 | !hbusreq3_p & v84561b;
assign v23fbde1 = hbusreq6 & v23fb8e4 | !hbusreq6 & !v22f7ef7;
assign v22ef458 = hbusreq5_p & v13afad9 | !hbusreq5_p & v2304e9c;
assign v23fcec8 = hbusreq3_p & v23fc19b | !hbusreq3_p & v23fc162;
assign v22f2e0c = hmaster0_p & v13afbf0 | !hmaster0_p & v23f0db7;
assign v23f6e68 = hbusreq1_p & v230da35 | !hbusreq1_p & !b8c90d;
assign b2aff2 = hgrant5_p & v23fbd93 | !hgrant5_p & v2312acc;
assign v2303ae3 = hbusreq6 & v22edb40 | !hbusreq6 & v230b08b;
assign v23fc0d8 = hbusreq3_p & v23f558b | !hbusreq3_p & v22ecd54;
assign v23fb410 = hbusreq2_p & v106af73 | !hbusreq2_p & v191a879;
assign v2312bae = jx3_p & v23f4928 | !jx3_p & v23f818e;
assign v22f991b = hbusreq2_p & e1df2d | !hbusreq2_p & v84561b;
assign v230b375 = hgrant1_p & v230d30a | !hgrant1_p & v2304c4c;
assign v23fcc05 = hbusreq4_p & v2312faa | !hbusreq4_p & v84561b;
assign bd761f = hmaster2_p & v22fb4de | !hmaster2_p & v2313131;
assign v230aa2f = hmaster2_p & aa6574 | !hmaster2_p & !v23f763f;
assign v22ec6e5 = hmaster2_p & v23068a9 | !hmaster2_p & !v84561b;
assign v23f0776 = hgrant3_p & v22ee657 | !hgrant3_p & v1aad31c;
assign v22fb6df = hbusreq4 & v23fb856 | !hbusreq4 & v22f18f3;
assign v230c342 = hlock1_p & v23f78a4 | !hlock1_p & !v22ff457;
assign v2392d6d = hbusreq2_p & v23fc151 | !hbusreq2_p & !v191a879;
assign v22f86d2 = hmaster0_p & v84561b | !hmaster0_p & v2391e3e;
assign v22fb554 = hbusreq3_p & b9c8ff | !hbusreq3_p & v22f9c5f;
assign v23fcfe8 = hmaster1_p & v22f721f | !hmaster1_p & v230334d;
assign v23fc3bf = hgrant5_p & v191ae81 | !hgrant5_p & v22f322a;
assign v23f4015 = hmaster0_p & v2311831 | !hmaster0_p & v22f8eb8;
assign v23f7cbe = hbusreq6_p & v2306cca | !hbusreq6_p & v191acb4;
assign v22fdf59 = hlock4_p & v23066fe | !hlock4_p & v230936c;
assign v22f4ab3 = hlock5_p & da38c1 | !hlock5_p & v84561b;
assign v23fcbe3 = hbusreq1 & v2301d45 | !hbusreq1 & v230c52a;
assign v23fc744 = hbusreq1 & v230358b | !hbusreq1 & v84561b;
assign v23f8364 = locked_p & v230fdc7 | !locked_p & v84561b;
assign v23f4979 = hbusreq5_p & v23fbc5a | !hbusreq5_p & !v84561b;
assign v23fb93f = hmaster2_p & v23fbde0 | !hmaster2_p & v23f328e;
assign d7df7e = hbusreq3 & v23fca9c | !hbusreq3 & v23fc4d1;
assign v191ac87 = hbusreq6_p & v23fcbb0 | !hbusreq6_p & v84561b;
assign bdac8d = hbusreq5 & v23fbbf2 | !hbusreq5 & v845622;
assign v23fc1ce = hgrant1_p & v845626 | !hgrant1_p & v22ede16;
assign v23105aa = hbusreq3_p & v23fca08 | !hbusreq3_p & v1aad641;
assign v2305a05 = hmaster2_p & v23f572e | !hmaster2_p & v23fcf89;
assign v2305797 = hmaster0_p & v23fbb50 | !hmaster0_p & v84561b;
assign v23f069d = hgrant1_p & v94e4a6 | !hgrant1_p & v230a2b1;
assign v230154b = hlock5_p & v23fb914 | !hlock5_p & !v84561b;
assign v230eab7 = hmaster2_p & v23f7700 | !hmaster2_p & v22f0593;
assign v23f8f24 = jx3_p & v84561b | !jx3_p & v23fbe7c;
assign v23fcd34 = stateG10_5_p & v23925af | !stateG10_5_p & v230fec6;
assign v23fc324 = hbusreq3_p & v23f3d5b | !hbusreq3_p & v22fd907;
assign v22f3d67 = hmaster0_p & v23f90b2 | !hmaster0_p & !v2302cfa;
assign v23fc29d = hbusreq6 & v22ec2c4 | !hbusreq6 & v22ef062;
assign v23f9dd1 = hbusreq1_p & v23fcf49 | !hbusreq1_p & !v84561b;
assign v23fb96b = hbusreq4 & v23efac1 | !hbusreq4 & v23fc931;
assign v230159e = hmaster2_p & v23f9370 | !hmaster2_p & v2308a4b;
assign v2300b7b = hmaster0_p & v2307fcd | !hmaster0_p & v2303ae3;
assign fc8c57 = stateG10_5_p & v230828c | !stateG10_5_p & v2309c93;
assign v23fc4b7 = hbusreq4_p & v2304d08 | !hbusreq4_p & v23fb7a3;
assign v23fc449 = hlock4_p & v230a193 | !hlock4_p & v22fb147;
assign v230ce74 = hbusreq4_p & v1aadc9e | !hbusreq4_p & v23fc19e;
assign v23fcdb9 = hmastlock_p & v22eb3aa | !hmastlock_p & v84561b;
assign v22fe285 = hmaster2_p & v22feb47 | !hmaster2_p & v845620;
assign v23fc8d1 = hmaster2_p & bd74c0 | !hmaster2_p & v22f0073;
assign v23fbc7e = hgrant3_p & v22f7c9a | !hgrant3_p & v23fd069;
assign v230de17 = hmaster1_p & v22fd796 | !hmaster1_p & v230cc30;
assign v230cff9 = hready & v22f6ba1 | !hready & !v84561b;
assign v22f98e7 = hbusreq3_p & v22f8f2b | !hbusreq3_p & v22ec1f4;
assign v23f86f0 = locked_p & v230650d | !locked_p & v106ae19;
assign v2309945 = hlock2_p & v84561b | !hlock2_p & v22f60c6;
assign v22f2cf1 = hmaster2_p & v23fb98a | !hmaster2_p & !v84561b;
assign v23fbd5d = hmaster2_p & v230cb9a | !hmaster2_p & v23fbedc;
assign v23fbaef = hbusreq2 & v23fcf9b | !hbusreq2 & v84561b;
assign v23fbad7 = hmaster0_p & v2301190 | !hmaster0_p & v23fcdb6;
assign v23fb2e5 = hgrant2_p & v23f3e7f | !hgrant2_p & v23117af;
assign v22f0fcd = hbusreq4_p & bd8ac4 | !hbusreq4_p & v23fcbaf;
assign v22f752e = hmaster0_p & v2310eb0 | !hmaster0_p & v23fc587;
assign v23fc029 = hmaster0_p & v22eb711 | !hmaster0_p & v230f0de;
assign v23fb95f = hgrant3_p & v23fbef6 | !hgrant3_p & v2307553;
assign v23fcfda = hbusreq4_p & v23fcc43 | !hbusreq4_p & v23fbad7;
assign v23f593e = hbusreq6 & v23f626c | !hbusreq6 & v23fc147;
assign v22f25e6 = hgrant3_p & v22fe924 | !hgrant3_p & v23fba0f;
assign v22efef6 = hlock3_p & v22f939d | !hlock3_p & !v23fc324;
assign v2301e9a = hbusreq3_p & da38c1 | !hbusreq3_p & v230129b;
assign v2310ff6 = hbusreq3 & v23f6659 | !hbusreq3 & v84561b;
assign v22eb599 = hbusreq1_p & v23064ff | !hbusreq1_p & v22fe428;
assign v22f4e7f = hlock0_p & b572e8 | !hlock0_p & v15074df;
assign v2308d79 = busreq_p & v231066c | !busreq_p & v22fa4dd;
assign v22f53b4 = hbusreq5_p & v2309b3c | !hbusreq5_p & v2302e87;
assign v23f19b4 = hgrant0_p & v84561b | !hgrant0_p & !v88bc32;
assign v23f89f4 = hmaster1_p & v84561b | !hmaster1_p & v23fcd91;
assign v23109e3 = hlock4_p & v23fbff9 | !hlock4_p & v23f232d;
assign v23f8d53 = hbusreq6 & v22edbd5 | !hbusreq6 & v84561b;
assign v23fbd48 = hgrant3_p & v98d402 | !hgrant3_p & v22ffdc5;
assign v2302a77 = hmaster2_p & v22f11fe | !hmaster2_p & v84561b;
assign v23089ec = hbusreq1 & v230ca0f | !hbusreq1 & !v84561b;
assign v23fca15 = hbusreq5_p & v22fd8a6 | !hbusreq5_p & v22eb6ee;
assign v23fcfbf = hgrant5_p & v84561b | !hgrant5_p & v23fcbb2;
assign b09503 = hmastlock_p & v23fc32b | !hmastlock_p & v84561b;
assign v98d297 = hbusreq5 & v22efcd6 | !hbusreq5 & v23fc839;
assign v1aad8a4 = hbusreq3 & v84564d | !hbusreq3 & v22f23a1;
assign v23fbfb9 = locked_p & v230bf69 | !locked_p & v191a86f;
assign v23089cd = hmaster1_p & v23fce60 | !hmaster1_p & !v23f49cd;
assign v22fd445 = hbusreq4_p & v22f41c4 | !hbusreq4_p & v22f9f2a;
assign v22ef8af = hlock2_p & v22f53a6 | !hlock2_p & v23f0ce0;
assign v2300ba2 = hbusreq3 & ae0418 | !hbusreq3 & v84561b;
assign v2304373 = hbusreq6_p & v22fa202 | !hbusreq6_p & !v84561b;
assign v23f9127 = hlock0_p & v22fd387 | !hlock0_p & !v84561b;
assign v22f1905 = hbusreq5_p & v23fca0a | !hbusreq5_p & !v23088a4;
assign v22fe0cb = hmaster0_p & v2300d5f | !hmaster0_p & v230b38b;
assign v22ed7d3 = hbusreq2_p & v2307ff9 | !hbusreq2_p & v84561b;
assign v2300c06 = hmaster0_p & v22f0dc9 | !hmaster0_p & v22f76c6;
assign v23fc566 = hgrant3_p & v23fc75d | !hgrant3_p & v15075e0;
assign v230e916 = hbusreq5_p & v22fa76f | !hbusreq5_p & v84561b;
assign v2301aab = hbusreq0 & v23fba6b | !hbusreq0 & !v84561b;
assign v230dae4 = hmaster2_p & v191aa95 | !hmaster2_p & v84561b;
assign v23fbd80 = hlock5_p & v2311089 | !hlock5_p & v9052d9;
assign v22f166b = hgrant4_p & v845629 | !hgrant4_p & v230eaba;
assign v22f4d97 = hmaster2_p & v84561b | !hmaster2_p & !v23f301a;
assign v230bdf9 = hbusreq5_p & v1e83fd9 | !hbusreq5_p & v23f4938;
assign v22edd99 = hmaster0_p & b00aa6 | !hmaster0_p & v22ebddc;
assign v23f12d3 = hgrant3_p & v845635 | !hgrant3_p & v23fc5b6;
assign v230b8cd = hgrant0_p & v84561b | !hgrant0_p & v2391bb7;
assign v22f2db0 = hbusreq2_p & v23919a5 | !hbusreq2_p & v84561b;
assign v22ef56f = hbusreq5_p & b9d00f | !hbusreq5_p & v1e840d3;
assign v23f3922 = hbusreq4_p & v23faada | !hbusreq4_p & v22efcad;
assign v23000e2 = hbusreq1_p & v2303558 | !hbusreq1_p & !v23046f7;
assign v22ff6a2 = hmaster2_p & v23fb6e3 | !hmaster2_p & v22f1ece;
assign v2307b17 = hbusreq3_p & v2346b79 | !hbusreq3_p & v23fcd70;
assign v22ef0a0 = hmaster1_p & v23fbe8f | !hmaster1_p & !v23f49cd;
assign v23f89db = hgrant2_p & v22fa827 | !hgrant2_p & !v22eaf7a;
assign v23fc7b7 = hmaster2_p & v230b1ac | !hmaster2_p & v23fbf24;
assign v2310ada = hbusreq6 & v22ed4e1 | !hbusreq6 & v84561b;
assign v23fba79 = hgrant2_p & v2307ff5 | !hgrant2_p & v2302e32;
assign v23025aa = hbusreq0_p & v23fbb84 | !hbusreq0_p & v23fab82;
assign v23fa837 = hmaster2_p & v2312ad2 | !hmaster2_p & v2313131;
assign v22eb674 = hbusreq4_p & v23fc169 | !hbusreq4_p & v23f2199;
assign v23f56de = hgrant3_p & v23fc7a7 | !hgrant3_p & v230b68a;
assign v23f2cbe = hbusreq1 & v2301655 | !hbusreq1 & v84562a;
assign v22f2de3 = hlock3_p & v22f53e2 | !hlock3_p & v230f3e5;
assign v23fc330 = hmaster0_p & v239308e | !hmaster0_p & !v22faa86;
assign v23fb9e5 = hbusreq4_p & v84562b | !hbusreq4_p & v23fbc65;
assign v1aad323 = hbusreq3 & v22f586f | !hbusreq3 & v84561b;
assign v23fb648 = hgrant2_p & v230f253 | !hgrant2_p & v84561b;
assign v22f67ef = hbusreq1_p & v22fbc05 | !hbusreq1_p & v22f0dd6;
assign v23f9812 = hmaster1_p & v84561b | !hmaster1_p & v2311e38;
assign v23fb9ca = hbusreq3_p & v230e473 | !hbusreq3_p & v230c0e6;
assign v23fc598 = hbusreq4_p & v2307c63 | !hbusreq4_p & v23fccd7;
assign v23f5d23 = hmaster2_p & v23fc5d9 | !hmaster2_p & v22fa3e9;
assign v23fc247 = hgrant3_p & v1aad421 | !hgrant3_p & v23f53e9;
assign v22f1f6f = hlock0_p & v23f6411 | !hlock0_p & !v106ae19;
assign v230818b = hbusreq0 & v191a86f | !hbusreq0 & !v84561b;
assign v23fce81 = hbusreq1_p & v23fc9f3 | !hbusreq1_p & v1aae262;
assign v23fca3b = hmaster1_p & v84561b | !hmaster1_p & !v22fd2a3;
assign v23fc546 = hbusreq4 & v22eda3a | !hbusreq4 & v23fc6ab;
assign v22f7800 = hgrant3_p & v84561b | !hgrant3_p & v22f8af0;
assign v22f8cd9 = hbusreq3_p & b9d0a0 | !hbusreq3_p & v23fbe26;
assign v22eee99 = hmaster2_p & v23fbd52 | !hmaster2_p & v23fbaaa;
assign v230c8e9 = hbusreq1_p & v2305bb2 | !hbusreq1_p & v84561b;
assign v22f5429 = hmaster1_p & v230be9e | !hmaster1_p & v23013f8;
assign v22f3ad4 = hlock1_p & v2313463 | !hlock1_p & !v84561b;
assign v22f1b30 = hbusreq4 & v2309ca8 | !hbusreq4 & v150718d;
assign v2313a33 = hlock0_p & v23f55c0 | !hlock0_p & v2300597;
assign v22f728a = hmaster2_p & v22fc80c | !hmaster2_p & v23f79f6;
assign v22fb0c7 = hmaster2_p & v23fc6c0 | !hmaster2_p & v23080ec;
assign e1e707 = hmaster2_p & v84561b | !hmaster2_p & v23f797b;
assign v23002e0 = hbusreq1 & v23fce71 | !hbusreq1 & v84561b;
assign v22f7879 = hgrant1_p & f406c6 | !hgrant1_p & !v23fc78e;
assign v22f0139 = hbusreq1_p & v23f4154 | !hbusreq1_p & v22f3e14;
assign v22ed2f5 = hbusreq3_p & v22f61b6 | !hbusreq3_p & v23f660f;
assign v2307942 = hbusreq3_p & v230a3f5 | !hbusreq3_p & v84561b;
assign v239298e = jx0_p & v23fbb81 | !jx0_p & v23fc45d;
assign v22ed533 = hmaster2_p & v2312990 | !hmaster2_p & !v84561b;
assign v22eb06f = hbusreq1 & v23f8f21 | !hbusreq1 & !v23fbbd2;
assign v191acb4 = hbusreq4_p & v845633 | !hbusreq4_p & !v84561b;
assign v23f32eb = locked_p & v23fc3de | !locked_p & v84561b;
assign v23fc0a3 = hbusreq4 & v230b236 | !hbusreq4 & v84562f;
assign v1aae09e = hgrant1_p & v23fc5f4 | !hgrant1_p & v84561b;
assign v22f1aed = hmaster1_p & v2305a14 | !hmaster1_p & v22ed363;
assign v2308c50 = hbusreq1 & v22f31b2 | !hbusreq1 & !v23fcf77;
assign v23f8395 = hgrant2_p & v1e83fd9 | !hgrant2_p & v22f3f06;
assign v23f3508 = hmaster2_p & v23fbaaa | !hmaster2_p & v23f8e6b;
assign v96c563 = hbusreq6 & v23fc905 | !hbusreq6 & !v22fda6e;
assign v23fcfd0 = hmaster2_p & v84564d | !hmaster2_p & v22fc34e;
assign v22f5d87 = hbusreq1 & v230358b | !hbusreq1 & v2312ea7;
assign v22f70b0 = hbusreq1 & v23fa4ca | !hbusreq1 & v84561b;
assign v2303554 = jx0_p & v2392811 | !jx0_p & v230418f;
assign v22fe582 = hbusreq5_p & v23fcf46 | !hbusreq5_p & v22fa662;
assign v230fd50 = hmaster2_p & v2313131 | !hmaster2_p & v23fbdc1;
assign v230d14d = hmaster2_p & v22ed6c5 | !hmaster2_p & v1aae56f;
assign v23fab8b = hlock0_p & v23fceb9 | !hlock0_p & v23fcadd;
assign v22f7c9a = hbusreq3_p & v2309df7 | !hbusreq3_p & v23fbe21;
assign v23f28ed = hmaster0_p & v2309c9d | !hmaster0_p & v2393f05;
assign v2306f5b = hmaster2_p & v23930d2 | !hmaster2_p & !v23f63ab;
assign v23fc549 = hbusreq3 & fc88ba | !hbusreq3 & v84561b;
assign v23fce91 = stateG10_5_p & v2307e2c | !stateG10_5_p & v845636;
assign a296f8 = hmaster0_p & v898be2 | !hmaster0_p & !v96c563;
assign v2310b0b = hbusreq3 & v22ef350 | !hbusreq3 & v84561b;
assign v23106c2 = jx2_p & v23f4a0f | !jx2_p & v22f9532;
assign v23fc988 = hmaster2_p & v23fc742 | !hmaster2_p & v23f4da0;
assign v22ff63a = hbusreq4 & v230591e | !hbusreq4 & v230bece;
assign v23f4491 = hbusreq1_p & v23f25c8 | !hbusreq1_p & v22f8d8e;
assign v230226e = hmaster1_p & v22f694d | !hmaster1_p & v84561b;
assign v23fcb65 = hbusreq1_p & v2301edd | !hbusreq1_p & v84561b;
assign v230d8f3 = hmaster2_p & v84561b | !hmaster2_p & v230cfed;
assign v2303db8 = hbusreq3_p & v845636 | !hbusreq3_p & !aeff78;
assign v22f9374 = hbusreq3_p & v22efe1b | !hbusreq3_p & v230a579;
assign v230f96f = hgrant3_p & v2393332 | !hgrant3_p & v230891d;
assign v23f05ee = hmaster0_p & v191a8e5 | !hmaster0_p & v22f7347;
assign v23f963f = hbusreq3 & v22f1244 | !hbusreq3 & v22f9eb0;
assign v2303b1a = hmaster2_p & v2313463 | !hmaster2_p & !v23f908f;
assign v22f2188 = hbusreq3 & aaca7f | !hbusreq3 & v23fbf1c;
assign v932767 = hmaster2_p & v23fc4a5 | !hmaster2_p & v230c876;
assign v230ef0b = hbusreq1_p & v2301884 | !hbusreq1_p & v84561b;
assign v22f3499 = hbusreq5_p & v22eb377 | !hbusreq5_p & v90aa06;
assign v23fb43a = hmaster0_p & v22f789c | !hmaster0_p & v23f6fa8;
assign v23f68ab = hmaster2_p & v2312696 | !hmaster2_p & v23fa345;
assign bd837d = hbusreq3_p & b9d00f | !hbusreq3_p & v1aadf44;
assign v22ec801 = hbusreq5 & v22ee9be | !hbusreq5 & v84561b;
assign v22f7e59 = hbusreq1_p & v23f6e45 | !hbusreq1_p & v23fb5b4;
assign v23fc5e8 = hmaster2_p & v23fce6b | !hmaster2_p & !v84561b;
assign v23fc4ef = jx0_p & v22f0e84 | !jx0_p & v22f7ce8;
assign v230206c = hbusreq6 & v22ff0be | !hbusreq6 & v23fc84a;
assign v22f14ee = hmaster0_p & bd7ae5 | !hmaster0_p & v23f7fb6;
assign v23fc88c = hmaster2_p & v23f5af5 | !hmaster2_p & !b9d013;
assign v2300617 = hmaster2_p & v23fb0ce | !hmaster2_p & v23fbaaa;
assign v23fbe51 = hlock0_p & a1fc4e | !hlock0_p & v1507088;
assign f40d81 = hgrant2_p & e1df2d | !hgrant2_p & v84561b;
assign v23ef8ef = hgrant2_p & v22f2f87 | !hgrant2_p & !v230e78c;
assign v239223a = hgrant3_p & v84561b | !hgrant3_p & v15070ca;
assign v845639 = hbusreq6_p & v84561b | !hbusreq6_p & !v84561b;
assign v22fa23d = hlock4_p & v13afb18 | !hlock4_p & v845637;
assign v22ec5f6 = hlock5_p & v22f1b31 | !hlock5_p & bbc337;
assign v22f4266 = hgrant3_p & v84562e | !hgrant3_p & v22fdd65;
assign v22f1899 = hmaster2_p & v23f9226 | !hmaster2_p & v230590b;
assign v22fa9ce = hmaster2_p & v22f0132 | !hmaster2_p & v22fee3b;
assign v22f44cc = hbusreq3_p & v230fb0a | !hbusreq3_p & v22f61b6;
assign v23fcc1e = jx1_p & v85e5cf | !jx1_p & !v23f39d9;
assign v230d910 = hbusreq3_p & v22ff90b | !hbusreq3_p & v230080a;
assign v22f0bea = stateG2_p & v84561b | !stateG2_p & v230db9d;
assign v1aae124 = hmaster1_p & v23fc009 | !hmaster1_p & v2310037;
assign v191ac53 = hbusreq3 & v23fbcbf | !hbusreq3 & v84561b;
assign v22ff09a = hbusreq4_p & v22f20cf | !hbusreq4_p & v2301968;
assign v23f2ecd = hbusreq2_p & v23f5872 | !hbusreq2_p & v84561b;
assign v23fcdd5 = hbusreq0 & v845620 | !hbusreq0 & v23017f0;
assign v2305c1f = hgrant1_p & v84561b | !hgrant1_p & v23fc3bf;
assign v22f884c = hmaster0_p & v22f5b7c | !hmaster0_p & v2300c85;
assign v23fcadd = hbusreq0_p & v23fceb9 | !hbusreq0_p & v23fb172;
assign v22f882c = hmaster0_p & v22eb184 | !hmaster0_p & v22f3998;
assign v23fc126 = hbusreq1 & v23fa4ca | !hbusreq1 & !v84561b;
assign v23f31d3 = stateG10_5_p & v22f84ff | !stateG10_5_p & v845636;
assign v23fbe76 = hbusreq3 & v895d68 | !hbusreq3 & v22fe2ae;
assign b95000 = hmaster2_p & v84561b | !hmaster2_p & v23f908f;
assign v22ed1f3 = stateG10_5_p & v22f299f | !stateG10_5_p & v23fbb80;
assign v22ef9aa = hmaster0_p & v23081e8 | !hmaster0_p & !v23fcb43;
assign v22fab2d = jx1_p & c16602 | !jx1_p & v191acb4;
assign fc8fe6 = hmaster2_p & v230935d | !hmaster2_p & v22fe426;
assign v22fec8c = hbusreq1_p & v85d110 | !hbusreq1_p & v22eefd1;
assign v22ec240 = jx1_p & v23fcfed | !jx1_p & v22fb42c;
assign v230b086 = hmaster2_p & v2310754 | !hmaster2_p & v23fc164;
assign v230e032 = hmastlock_p & v23fc1c7 | !hmastlock_p & v84561b;
assign v2306fa2 = hbusreq2_p & v23f9a93 | !hbusreq2_p & !v22f36ff;
assign v23f17e2 = hgrant5_p & v230b750 | !hgrant5_p & v23083e6;
assign v2303c07 = hmaster2_p & v23f9789 | !hmaster2_p & v22f0945;
assign v23fb564 = hburst0_p & v84561b | !hburst0_p & v22f9cb4;
assign v22fd411 = jx3_p & v23fc3d8 | !jx3_p & v23fcb16;
assign v230e45a = hbusreq3_p & v22f2718 | !hbusreq3_p & !v84561b;
assign v22f78b4 = hbusreq6_p & v22f0d4e | !hbusreq6_p & v22f1d4f;
assign v23fc27c = hbusreq3 & v12cd692 | !hbusreq3 & !v84561b;
assign v8d360e = busreq_p & v191a86f | !busreq_p & !v23fc2dd;
assign v23fba98 = hlock5_p & v22ff613 | !hlock5_p & v845620;
assign v23f2bc0 = hbusreq3_p & v845627 | !hbusreq3_p & v22f9160;
assign v230aa0c = hmaster0_p & v22fa101 | !hmaster0_p & v22f7564;
assign v22f58cd = hbusreq4 & v22fb36e | !hbusreq4 & v84561b;
assign v230b0f9 = hmaster0_p & v23f29e9 | !hmaster0_p & v23fccb3;
assign v22f8aec = hgrant1_p & v23f6bc1 | !hgrant1_p & v23fbdac;
assign v22ff727 = hmaster1_p & v23f38b1 | !hmaster1_p & v23fc822;
assign a1fd78 = hmaster0_p & v2393c48 | !hmaster0_p & !v23fc6a7;
assign v22f6b4c = hgrant1_p & v22f0824 | !hgrant1_p & v22f7ef4;
assign v2313372 = hgrant2_p & v84561b | !hgrant2_p & v22f991b;
assign v231353a = hgrant4_p & v23934cb | !hgrant4_p & v23fce6f;
assign v23fb681 = hbusreq6_p & v23fc827 | !hbusreq6_p & v22ee524;
assign v23fc439 = hmaster2_p & v23fb6e3 | !hmaster2_p & v23f2c05;
assign v230d6fd = hgrant3_p & v84561b | !hgrant3_p & v23919c0;
assign v23fbb84 = hbusreq0 & v191accc | !hbusreq0 & v84562a;
assign v22fd169 = hmaster0_p & v22ef734 | !hmaster0_p & v23f193e;
assign v22f8105 = stateG2_p & v84561b | !stateG2_p & v23f8e0b;
assign stateG3_2 = !a1f79d;
assign v22f755a = hbusreq6 & v23fbdb9 | !hbusreq6 & v84561b;
assign v22f2450 = hbusreq3_p & v13afb18 | !hbusreq3_p & v22f4114;
assign v230095f = hmaster1_p & v23fc6be | !hmaster1_p & !v12cd586;
assign v23115e2 = hbusreq3_p & v2311967 | !hbusreq3_p & v22fcf75;
assign v22ec350 = hbusreq6 & v23f3ff9 | !hbusreq6 & v230f0de;
assign v2305782 = hmaster2_p & v84564d | !hmaster2_p & v22f1a26;
assign v23fc48a = hbusreq4_p & v1aad5ee | !hbusreq4_p & v230c440;
assign v23fcc10 = hready & v22fbf54 | !hready & v230d7b7;
assign v2302e7b = hlock4_p & v22f8c01 | !hlock4_p & !v22f9cd9;
assign v23027cd = hmaster2_p & v23fcac2 | !hmaster2_p & v22fa5fd;
assign v2305819 = hbusreq6_p & v2301450 | !hbusreq6_p & v23fb299;
assign v230cc30 = hbusreq4_p & v22f207c | !hbusreq4_p & v2311246;
assign v22ed5c5 = hgrant3_p & v2301463 | !hgrant3_p & v23fbb73;
assign v23fcbc9 = hlock3_p & v23f0a6b | !hlock3_p & v22eb338;
assign v1aad346 = hmaster1_p & v23fc1b9 | !hmaster1_p & v23fd00e;
assign v23f7898 = hgrant5_p & v84561b | !hgrant5_p & v23fcdac;
assign v23f0169 = hlock0_p & v1506a4d | !hlock0_p & v23f1ca1;
assign v22fbb0f = hbusreq4_p & v230edb2 | !hbusreq4_p & v23fbf3b;
assign v22fb10b = hgrant3_p & v13afe72 | !hgrant3_p & v2302b2c;
assign v23efcf8 = hmaster2_p & v84561b | !hmaster2_p & v23fc6c4;
assign v22f33c4 = hmaster2_p & v230a51c | !hmaster2_p & v22ee0db;
assign v2308dbf = hmaster0_p & v2306d08 | !hmaster0_p & v23037ac;
assign v230f1d6 = hbusreq4_p & v23f8d36 | !hbusreq4_p & v23fcc52;
assign v230cea0 = hgrant3_p & v230e817 | !hgrant3_p & v23fc748;
assign v22f2f44 = hbusreq5_p & v23fbb0f | !hbusreq5_p & v84561b;
assign v2303125 = hgrant0_p & v84561b | !hgrant0_p & v2307946;
assign v230894d = hbusreq1 & v22f926d | !hbusreq1 & v230c025;
assign v2300936 = hbusreq5_p & v22fc745 | !hbusreq5_p & v12cd4c6;
assign v23fc9ee = hbusreq3_p & v230c95c | !hbusreq3_p & v22f5235;
assign v22fab7c = hmaster2_p & v22f79fd | !hmaster2_p & v23f2be7;
assign v2306e28 = hbusreq3_p & d962e3 | !hbusreq3_p & v23fba9a;
assign v23fc80d = hbusreq3_p & v2307224 | !hbusreq3_p & v2300ccc;
assign v22fd372 = hbusreq1 & v23f8cd3 | !hbusreq1 & v84561b;
assign v2311089 = hbusreq5 & v22fcf71 | !hbusreq5 & v84561b;
assign v23fa4bb = hmaster2_p & v230031f | !hmaster2_p & v230de18;
assign v23fbaa8 = hbusreq3_p & v2391f3c | !hbusreq3_p & v23050c1;
assign v22ec1cb = hburst0_p & v84561b | !hburst0_p & v84563f;
assign v23fb949 = hbusreq3 & v23fcd63 | !hbusreq3 & v23f3f59;
assign v2313476 = hlock5_p & v845620 | !hlock5_p & !v84561b;
assign v2304ccc = hmaster2_p & v23fbdb0 | !hmaster2_p & v23fc48b;
assign a1fdac = hgrant3_p & v22f6ae5 | !hgrant3_p & v23f3508;
assign v22f4ee6 = hgrant3_p & v230f14b | !hgrant3_p & v23fcdc1;
assign v22ee913 = hgrant6_p & v23fce08 | !hgrant6_p & v23f1f3f;
assign v230e874 = hbusreq3 & v23fc32d | !hbusreq3 & !v23f36e9;
assign v23fc561 = hbusreq1 & v22fc5f0 | !hbusreq1 & v22f5583;
assign v23fcb3b = hgrant3_p & v22ee47d | !hgrant3_p & v23f7aea;
assign v230f0a1 = stateA1_p & v84561b | !stateA1_p & v845667;
assign v22f1943 = hbusreq2 & v23fc23d | !hbusreq2 & v84561b;
assign v230ed8b = hbusreq1_p & v22f98ad | !hbusreq1_p & v84561b;
assign v230efeb = hbusreq5_p & v9526ac | !hbusreq5_p & !v23134a0;
assign v23fcb78 = hbusreq6_p & v23fc621 | !hbusreq6_p & v23f3d91;
assign v23f0b27 = hbusreq4_p & v23fc942 | !hbusreq4_p & v84561b;
assign v23f0162 = hlock0_p & v84561b | !hlock0_p & v23fb314;
assign v2304669 = hbusreq3 & v23fcd6b | !hbusreq3 & v84561b;
assign v22feb6e = hbusreq5 & v23f8f21 | !hbusreq5 & v84561b;
assign v230a355 = hlock1_p & v23f4154 | !hlock1_p & v23f7eaa;
assign v2312f3c = hlock0_p & v22f9e5b | !hlock0_p & v22fe0ee;
assign v230e71f = hgrant2_p & v17a34ff | !hgrant2_p & !v845647;
assign a05106 = hlock4_p & v22f0974 | !hlock4_p & v230d532;
assign v22eece2 = hlock1_p & v23fb28e | !hlock1_p & v23fb574;
assign v22f4678 = hgrant0_p & v845623 | !hgrant0_p & v22fdd09;
assign v23f84b2 = hbusreq5_p & v23fc315 | !hbusreq5_p & v23f95ef;
assign v230fb76 = hmaster2_p & v22f0945 | !hmaster2_p & v23f9789;
assign v22f3eed = hmaster0_p & v22ed711 | !hmaster0_p & !v23fbe02;
assign v22f9567 = hbusreq5 & v23fb9ad | !hbusreq5 & v84561b;
assign v23fc9d3 = hgrant1_p & v23126c9 | !hgrant1_p & v84561b;
assign v1aad8c1 = hmaster2_p & v23f2513 | !hmaster2_p & v84561b;
assign v22fd030 = hgrant4_p & v23fbc19 | !hgrant4_p & v230adfa;
assign v22f20a2 = hmaster0_p & v22f853d | !hmaster0_p & v23fc75d;
assign v22f76f0 = hlock0_p & v2303d8f | !hlock0_p & v23fb4d4;
assign v22f6d45 = hgrant3_p & v230e539 | !hgrant3_p & v22eb498;
assign v23f61ba = hmaster2_p & v22f5820 | !hmaster2_p & v84561b;
assign v23fc334 = hmaster0_p & v23fcbd0 | !hmaster0_p & v230c437;
assign v22ec934 = hbusreq3_p & bd74f4 | !hbusreq3_p & v22fd196;
assign v2302c67 = hmaster2_p & v191a86f | !hmaster2_p & v23fb029;
assign stateG10_6 = !b8f86b;
assign v22f65dd = hmaster0_p & v23fcd2a | !hmaster0_p & !v23fcd24;
assign v23fc94c = hlock0_p & v23f5cb3 | !hlock0_p & v2312de4;
assign v2309099 = stateG2_p & v2302ca3 | !stateG2_p & v23fc8f0;
assign v23108aa = hgrant5_p & v2304299 | !hgrant5_p & !v22ef3d4;
assign v22fbde3 = hgrant3_p & v22ffd0e | !hgrant3_p & v23f47e3;
assign v2305d69 = hbusreq2_p & v22f1943 | !hbusreq2_p & v22f6683;
assign v22f83d7 = hmaster0_p & v23fc2b7 | !hmaster0_p & v22fda8c;
assign v230aa5d = hmaster0_p & v23fb1bb | !hmaster0_p & v23fb0a8;
assign v23133b3 = hgrant5_p & v23115bd | !hgrant5_p & v22f6090;
assign v22fced7 = hbusreq0_p & v22f6a6b | !hbusreq0_p & v23f512e;
assign v23fcef5 = hbusreq5_p & v23fbc5a | !hbusreq5_p & v84561b;
assign v2392f52 = hbusreq4 & v84561b | !hbusreq4 & v23fba11;
assign v23fcb71 = hmaster2_p & v22f7b47 | !hmaster2_p & v2309c07;
assign v2305196 = hbusreq0 & v22f9911 | !hbusreq0 & v84561b;
assign v23fbc7b = hgrant6_p & v84561b | !hgrant6_p & v23000a8;
assign v2304904 = hmaster2_p & v23fbfb9 | !hmaster2_p & v2302e32;
assign v2308e98 = hlock0_p & v22eefab | !hlock0_p & v2393f0d;
assign v230969a = jx2_p & v23fb8d7 | !jx2_p & !v22f7063;
assign v2312259 = hbusreq2_p & v22f0677 | !hbusreq2_p & !v84561b;
assign v23fbbeb = hmaster0_p & v13afeb1 | !hmaster0_p & bd7f79;
assign v23fb8a2 = hgrant1_p & v22f6b45 | !hgrant1_p & v23f3940;
assign v23f11ae = hmaster1_p & v22f03ec | !hmaster1_p & v2309d7a;
assign v23f8f1d = hbusreq3 & v23fc64c | !hbusreq3 & !v845622;
assign v23fbc9e = hbusreq4_p & v23fb0bf | !hbusreq4_p & v22eaeaf;
assign v23fc143 = hlock1_p & v23fbfe5 | !hlock1_p & v84564d;
assign v22fb260 = hmaster0_p & v23fc2b7 | !hmaster0_p & v23fc247;
assign v22f5834 = hmaster2_p & v22ed878 | !hmaster2_p & v23124cc;
assign v8ef087 = hgrant1_p & v12cd9f9 | !hgrant1_p & !v230ed8b;
assign v23f63b2 = hbusreq2 & v2312f7e | !hbusreq2 & !v23022b1;
assign v23fc512 = hbusreq5_p & v84561b | !hbusreq5_p & !v845671;
assign v2311fc9 = stateG10_5_p & v23f6bf0 | !stateG10_5_p & !v23f8274;
assign v22fc945 = hmaster2_p & v1507134 | !hmaster2_p & v23f763f;
assign v22fa36d = hmaster0_p & v231003e | !hmaster0_p & v23fcd69;
assign v12cda15 = hlock1_p & v13afb18 | !hlock1_p & v2304bc1;
assign v84564f = hgrant0_p & v84561b | !hgrant0_p & !v84561b;
assign v2305d6f = hbusreq3_p & v22f515e | !hbusreq3_p & v22ed809;
assign v22fe1e5 = hbusreq6_p & v2310538 | !hbusreq6_p & v230a0e7;
assign v23f1ad7 = hbusreq3_p & v22efdfe | !hbusreq3_p & v23fc25e;
assign v23fb5e8 = hbusreq2_p & a1fbb6 | !hbusreq2_p & a1fba6;
assign v2311cea = jx1_p & v22f800e | !jx1_p & v22fcf35;
assign v23fced9 = hbusreq1 & b50bc7 | !hbusreq1 & v84561b;
assign v23062f8 = hbusreq5_p & v23035ba | !hbusreq5_p & v23f0386;
assign v22ebe13 = hbusreq4_p & v2312e39 | !hbusreq4_p & v22fe2b6;
assign v230cc95 = hmaster1_p & v23fcdcd | !hmaster1_p & v23f78df;
assign v1aae087 = hmastlock_p & v22f334e | !hmastlock_p & v84561b;
assign v15072af = hbusreq5_p & v230f050 | !hbusreq5_p & v191b1f3;
assign v23fba32 = hlock3_p & v23fcc21 | !hlock3_p & v230f911;
assign v22ed5a5 = hmaster2_p & v22ff0d7 | !hmaster2_p & v84561b;
assign v23055c3 = hgrant3_p & v84561b | !hgrant3_p & v23f7f8d;
assign v23fc7d7 = hbusreq5_p & v23fb67c | !hbusreq5_p & v22f8dea;
assign v23fc7f0 = hbusreq1 & v23128a1 | !hbusreq1 & v84561b;
assign v22f11f6 = hgrant2_p & v12cd69f | !hgrant2_p & v23fce71;
assign v22ebbea = locked_p & bf8fe1 | !locked_p & v84561b;
assign v22edbd5 = hbusreq4 & v22edb43 | !hbusreq4 & v84561b;
assign v22f9092 = stateG10_5_p & v22f532c | !stateG10_5_p & v23056b1;
assign v22fca28 = hgrant1_p & v23fc9dd | !hgrant1_p & v23f89df;
assign v230f257 = hlock4_p & v23fc7bb | !hlock4_p & v230c3aa;
assign v23f4cd4 = stateG10_5_p & v23fa3a4 | !stateG10_5_p & v23faf8a;
assign v23051a9 = hmaster0_p & v22eb651 | !hmaster0_p & v84561b;
assign v230be8f = hbusreq3_p & v22ee6e8 | !hbusreq3_p & v23010d9;
assign v22fb450 = hgrant5_p & v23fc605 | !hgrant5_p & v23f81cf;
assign v2391735 = hbusreq4_p & v23022ab | !hbusreq4_p & v23fbc74;
assign v22eca17 = hbusreq5_p & v84564d | !hbusreq5_p & v22f0542;
assign v23fb61f = hbusreq2_p & v22ec29a | !hbusreq2_p & v22f9c73;
assign v23127b2 = hbusreq4 & v23fc197 | !hbusreq4 & v84561b;
assign v22ed34b = hbusreq4_p & v23f259c | !hbusreq4_p & !v23fcb6d;
assign v23fbb27 = jx2_p & v22ee41e | !jx2_p & v1aad441;
assign v2305ea5 = hmaster1_p & v22f52a0 | !hmaster1_p & v84561b;
assign v23f36f9 = hgrant5_p & v23fc772 | !hgrant5_p & !v84561b;
assign bdc4e2 = hgrant1_p & v23fd017 | !hgrant1_p & v22ef45e;
assign add85b = hmaster2_p & v23094a3 | !hmaster2_p & v23fbe22;
assign v23fc53e = busreq_p & v23916d6 | !busreq_p & v23003a8;
assign v23fc4d8 = hmaster1_p & v23fc5ac | !hmaster1_p & v22fdf28;
assign bd74c6 = hbusreq3_p & v23fceb9 | !hbusreq3_p & v84562b;
assign v23fc76e = hmaster0_p & v22ee657 | !hmaster0_p & !v96c563;
assign v230da35 = hlock1_p & v23f7b33 | !hlock1_p & v230cdfb;
assign v22f3a91 = hgrant4_p & v23fc0b7 | !hgrant4_p & v23fc617;
assign v8f3940 = hlock3_p & v23fc20e | !hlock3_p & v23fb8cc;
assign v2310a55 = hbusreq5_p & v23f3d14 | !hbusreq5_p & v22ee9be;
assign v230d20f = hbusreq3 & v230c65f | !hbusreq3 & v84561b;
assign v23fc776 = hmaster1_p & v230de82 | !hmaster1_p & v23fc7f4;
assign v23fbe9d = hmaster0_p & v23fb82a | !hmaster0_p & !v22f4ef7;
assign v22fbe6a = hgrant1_p & v84561b | !hgrant1_p & v22f6c1b;
assign v22f62e3 = hmaster1_p & v2302d53 | !hmaster1_p & !v23f724a;
assign v22f1841 = jx0_p & v22f6d0b | !jx0_p & v2309410;
assign v230a050 = hbusreq5_p & v2302225 | !hbusreq5_p & v23fbb6a;
assign v22f9c5f = hmaster2_p & v23fcfb8 | !hmaster2_p & v22f65d5;
assign v231232b = hlock4_p & v23f8d1a | !hlock4_p & v23fb615;
assign v22f6ed4 = hgrant3_p & v84561b | !hgrant3_p & v23fa23d;
assign v23fbdcc = stateG2_p & v84561b | !stateG2_p & !v230de5a;
assign v22f0c6d = hmaster0_p & v1b8771f | !hmaster0_p & v22efe2f;
assign v1e845ac = hbusreq5 & v22f2db0 | !hbusreq5 & v23fa2ec;
assign v22f4008 = hbusreq2 & bd9916 | !hbusreq2 & v84561b;
assign v23f6653 = hbusreq5_p & v23f6411 | !hbusreq5_p & !v106ae19;
assign v2301b2d = hgrant2_p & v845620 | !hgrant2_p & !v23fc5ba;
assign v23014fb = hbusreq5 & v23f2d8c | !hbusreq5 & v84561b;
assign v22fc477 = hbusreq4_p & v22fe01a | !hbusreq4_p & v2301e8c;
assign v22f5fa8 = stateA1_p & v84561b | !stateA1_p & !v23004f9;
assign v23940ce = stateG10_5_p & v23f9c30 | !stateG10_5_p & v84564d;
assign v22fb373 = hgrant3_p & v84562f | !hgrant3_p & v23f2dd4;
assign v22f4d04 = hgrant0_p & v2304937 | !hgrant0_p & v23fb2e5;
assign v23fb923 = hgrant3_p & v22ede34 | !hgrant3_p & v23fc2b1;
assign v22f9056 = hgrant3_p & v23f3f65 | !hgrant3_p & v23113b5;
assign v22f52c3 = hmaster2_p & v23080ec | !hmaster2_p & v22fba03;
assign v23f7891 = hmaster0_p & v23fc8d6 | !hmaster0_p & v230ba79;
assign v23fc372 = hbusreq3_p & v23117c1 | !hbusreq3_p & v23fcc3d;
assign v22fe408 = hgrant3_p & v22ffa6e | !hgrant3_p & v23fcf8a;
assign v2311094 = hbusreq3_p & v23fc664 | !hbusreq3_p & v22f61b6;
assign v23fd01f = hmaster2_p & v84561b | !hmaster2_p & !v22ff315;
assign v230c5eb = hbusreq3_p & v230681b | !hbusreq3_p & v230a735;
assign fc8f90 = hmaster0_p & v22fc8e5 | !hmaster0_p & v23fbf36;
assign v22f7098 = hmaster2_p & v84561b | !hmaster2_p & v2303679;
assign v22eeecc = hbusreq3_p & v230dacd | !hbusreq3_p & v84561b;
assign v23fcb5c = stateG10_5_p & v2312acc | !stateG10_5_p & v23f5043;
assign v22f45ac = hbusreq4_p & v23fc2f1 | !hbusreq4_p & v23fba3f;
assign v23efa84 = hmaster2_p & v191aa68 | !hmaster2_p & v2309871;
assign v22f8f2b = hmaster2_p & v2309c93 | !hmaster2_p & v2302225;
assign v1aae175 = hbusreq0 & v23fc842 | !hbusreq0 & !v84561b;
assign v23f58bb = hmaster2_p & v23f4758 | !hmaster2_p & v23f5907;
assign v23f595d = hgrant5_p & v23f5276 | !hgrant5_p & v15071a5;
assign v2303068 = hbusreq1_p & v2306d29 | !hbusreq1_p & !v191a86f;
assign v22f80b8 = hbusreq2_p & v23fcee2 | !hbusreq2_p & v9526ac;
assign v23074aa = hmaster2_p & v22f954f | !hmaster2_p & v23fb175;
assign v22f0fe5 = hgrant3_p & v230d3c2 | !hgrant3_p & v230d8f3;
assign v23f38f8 = hmaster0_p & v23f6ad0 | !hmaster0_p & v92eb35;
assign v23f8368 = hbusreq4_p & v230a3e2 | !hbusreq4_p & v23fc505;
assign v230884d = hready_p & b20f9d | !hready_p & v22fbc4e;
assign v23044e2 = stateG10_5_p & v230c649 | !stateG10_5_p & v22f0945;
assign v23060b1 = hbusreq1 & v23fc658 | !hbusreq1 & v23f5acd;
assign v22f8088 = stateA1_p & v22f79de | !stateA1_p & v23fcaaa;
assign v23f96b0 = hbusreq6 & v230fb9e | !hbusreq6 & v845627;
assign v22eefc4 = hbusreq5_p & v23fcf46 | !hbusreq5_p & v22fe260;
assign v22ecb9d = hgrant0_p & v2393723 | !hgrant0_p & v84561b;
assign v230ef7c = hbusreq5 & v23003cc | !hbusreq5 & v84561b;
assign v23078f5 = stateG10_5_p & v230848d | !stateG10_5_p & !v84561b;
assign v230d5f4 = hbusreq2_p & v23fcff0 | !hbusreq2_p & v845620;
assign v23fb793 = hbusreq1_p & v22f60c6 | !hbusreq1_p & v84564d;
assign f4066e = hbusreq6 & v84564d | !hbusreq6 & v23fc1c2;
assign v23fc23e = hgrant3_p & v23fbba8 | !hgrant3_p & v23fcaf7;
assign v1aae12f = hbusreq3 & v23025d8 | !hbusreq3 & !v230fc56;
assign v22ff92f = hlock2_p & v22f8271 | !hlock2_p & !v23056b1;
assign v2302a4d = hbusreq1_p & v22fef4f | !hbusreq1_p & v22fe62b;
assign a1fc4e = locked_p & v23fc378 | !locked_p & v22fb4e3;
assign v22f58e8 = hbusreq6_p & v2391cf3 | !hbusreq6_p & v23f9e87;
assign v2312bd0 = hready & v23114a6 | !hready & v84561b;
assign v23f83d7 = hmaster1_p & v22f7c42 | !hmaster1_p & v23f12d0;
assign v230b7f4 = hmaster2_p & v84564d | !hmaster2_p & v23fb793;
assign ae2bc6 = hmastlock_p & v2306595 | !hmastlock_p & v84561b;
assign v1aad4d7 = hbusreq1_p & v23fbadd | !hbusreq1_p & v23fb0c9;
assign v23fbc96 = hbusreq3 & v23fcd0b | !hbusreq3 & v22f3f32;
assign v23f3e38 = hmaster2_p & v23fc393 | !hmaster2_p & !v230935d;
assign v22eec11 = hbusreq6 & v949c12 | !hbusreq6 & v84561b;
assign v23fc9f2 = hmaster1_p & v84561b | !hmaster1_p & v23fa599;
assign v23f3ff7 = hbusreq3_p & v230062b | !hbusreq3_p & v22fc351;
assign v22f45d7 = hmaster2_p & v22fae6e | !hmaster2_p & !v23fbca3;
assign v2304a45 = hmaster2_p & v2306997 | !hmaster2_p & v2313131;
assign v22fedf7 = hgrant3_p & v2304f4c | !hgrant3_p & v23fade4;
assign v23fc4a1 = hlock5_p & v23f5af5 | !hlock5_p & !v2309c8a;
assign v230bbce = hgrant1_p & v22f1e91 | !hgrant1_p & v22f2319;
assign v23efac1 = hmaster2_p & v230910b | !hmaster2_p & v22f8543;
assign v2311d04 = hbusreq3 & v23f6478 | !hbusreq3 & v84561b;
assign v23f9fa4 = hmaster2_p & v22fc091 | !hmaster2_p & v22fc5f0;
assign v23f91bc = hbusreq3_p & v23fc139 | !hbusreq3_p & v84561b;
assign v22eb41e = hbusreq3_p & v191b1e4 | !hbusreq3_p & v84561b;
assign v23fcf43 = hmaster2_p & v23fbf9f | !hmaster2_p & !v84561b;
assign v23fb492 = hbusreq4_p & da310c | !hbusreq4_p & v22fed4f;
assign v23fb081 = hbusreq6 & v23efdcb | !hbusreq6 & !v106a846;
assign v22ebd88 = hbusreq3 & v22f2e41 | !hbusreq3 & v22f9add;
assign v230a9a0 = hlock0_p & v2308fe7 | !hlock0_p & !v22fa48a;
assign v22fe036 = hlock6_p & v2301da2 | !hlock6_p & v230936c;
assign v23fbf5c = hmaster0_p & v2311c0b | !hmaster0_p & v230dd15;
assign a1fd0b = hbusreq2_p & v22f60c6 | !hbusreq2_p & v84564d;
assign v22f908b = hmaster0_p & v23f76dc | !hmaster0_p & !v96c563;
assign v230f538 = hmaster2_p & v1aae56f | !hmaster2_p & v23fb9c2;
assign v230ac22 = hbusreq3 & v2305a94 | !hbusreq3 & v84561b;
assign v2306e35 = hgrant1_p & v12cd9f9 | !hgrant1_p & v2301fe9;
assign v22ec2c4 = hmaster2_p & v22ef062 | !hmaster2_p & v22ff1dd;
assign v2312888 = hmaster2_p & v23f445f | !hmaster2_p & v23f7123;
assign v22f2bb8 = hlock3_p & v23f6d50 | !hlock3_p & bd9dce;
assign v23f4ff3 = hmaster0_p & v23f9885 | !hmaster0_p & v22fda8c;
assign v230f1ae = hlock5_p & v23fbf67 | !hlock5_p & !v84561b;
assign v23fb752 = hlock1_p & v106aead | !hlock1_p & !v84561b;
assign v23f99bb = hmaster0_p & v84561b | !hmaster0_p & v23f2426;
assign v230da4a = hlock0_p & v22fda49 | !hlock0_p & !v84561b;
assign v23fc2b4 = hbusreq4 & v22f6e56 | !hbusreq4 & v23f8ca8;
assign v2309263 = stateG2_p & v84561b | !stateG2_p & v2310bf7;
assign v22ed7a5 = hbusreq3_p & v23fcaff | !hbusreq3_p & v1aae2be;
assign v94701c = hgrant1_p & v84561b | !hgrant1_p & v96bd8b;
assign v23fc03c = hmaster2_p & v84561b | !hmaster2_p & v23f0d46;
assign v2302c02 = hlock4_p & v84561b | !hlock4_p & !v2301992;
assign v22fe908 = hbusreq6 & v23fc5de | !hbusreq6 & v845645;
assign v22fc5e2 = hgrant1_p & v2311ed4 | !hgrant1_p & v230f331;
assign v23fc67f = hbusreq3_p & e1e722 | !hbusreq3_p & v2300bb5;
assign v22f2d7c = hmaster2_p & v2302e9e | !hmaster2_p & v84561b;
assign v23fbf9a = hmaster1_p & v22f1e6a | !hmaster1_p & v2311b96;
assign v22f8240 = hbusreq3 & v230cd57 | !hbusreq3 & v22f1339;
assign v22ef1a3 = hbusreq5 & v1aae29a | !hbusreq5 & v23f8364;
assign v2304bcd = jx3_p & v22f85f6 | !jx3_p & v23fbd6c;
assign v2311f44 = hbusreq6_p & v22f81a7 | !hbusreq6_p & v23f8e1c;
assign v22f4989 = hbusreq6 & v23035f1 | !hbusreq6 & v84561b;
assign v94e407 = hmaster2_p & v2301a75 | !hmaster2_p & v22ef062;
assign v23fb679 = hmaster1_p & v23fb456 | !hmaster1_p & !v22f6963;
assign v23fc463 = stateG10_5_p & v22f532c | !stateG10_5_p & v106ae19;
assign v22efe81 = hmaster2_p & v23fbfb9 | !hmaster2_p & v22eb5b3;
assign v22fb592 = hbusreq3 & v23fce3a | !hbusreq3 & !v2309d55;
assign v22f6756 = hgrant1_p & v230945e | !hgrant1_p & v22f0d2b;
assign v23fbb5f = hgrant1_p & v22f4407 | !hgrant1_p & v22eb742;
assign v230694d = hmaster0_p & v2301c51 | !hmaster0_p & !v22f383c;
assign v22faf60 = hgrant5_p & v23fc205 | !hgrant5_p & v84564f;
assign v23f8c0b = hmaster2_p & v23f1207 | !hmaster2_p & v22f98fd;
assign v22fa8e6 = hbusreq1_p & v84561b | !hbusreq1_p & v845635;
assign v22f2cb3 = hbusreq1_p & v230bd05 | !hbusreq1_p & v22f79be;
assign v845629 = hbusreq2_p & v84561b | !hbusreq2_p & !v84561b;
assign v22f082c = hbusreq6_p & v23f1e1b | !hbusreq6_p & v22f41ab;
assign v23fc709 = hmaster2_p & fc8c3f | !hmaster2_p & a6b8e0;
assign v22eb2f1 = hgrant0_p & v22f36ba | !hgrant0_p & v22fba61;
assign v2307ff5 = hbusreq2_p & v23f5cb3 | !hbusreq2_p & !v2310e40;
assign v22f1de1 = hmaster2_p & v22fa70c | !hmaster2_p & v230e4ef;
assign v23025ae = hbusreq3_p & v230a573 | !hbusreq3_p & v84562b;
assign v2306625 = hgrant3_p & v23f03d2 | !hgrant3_p & v23fbf0e;
assign v22efcc1 = hbusreq6_p & v2311b1e | !hbusreq6_p & v23fb652;
assign v231200e = hbusreq5_p & v230eb9b | !hbusreq5_p & v22fd06d;
assign v2307170 = hmaster0_p & v23fcbfb | !hmaster0_p & v23fbdd8;
assign v22f82f1 = hmaster1_p & v22f63cc | !hmaster1_p & v84561b;
assign v1507134 = hbusreq0 & v23f8f21 | !hbusreq0 & v84561b;
assign v91b2de = hmaster2_p & v22fef4f | !hmaster2_p & !v22ffc69;
assign v23fcfdb = hmaster2_p & v23101b1 | !hmaster2_p & v22f01c1;
assign v2303fd8 = hbusreq3 & v22fd8f6 | !hbusreq3 & v84561b;
assign v22f7c6f = hgrant3_p & v22f09c5 | !hgrant3_p & v230e32f;
assign v23fc1b9 = hbusreq6_p & v2391fc6 | !hbusreq6_p & v230ad18;
assign a1fcbb = hlock5_p & v191ab5f | !hlock5_p & v2310a63;
assign v230bbaf = hmaster1_p & v23fbf13 | !hmaster1_p & v23fc8e5;
assign v22f54cb = hmaster2_p & v23fa397 | !hmaster2_p & !v84561b;
assign v22f324a = hmaster2_p & v22f4986 | !hmaster2_p & !v22eaaba;
assign d97946 = hmaster0_p & v2312a90 | !hmaster0_p & v23fba11;
assign v23fc35f = hmaster2_p & v23fbf8b | !hmaster2_p & !v23fc51c;
assign v230d16b = hgrant0_p & v22f1133 | !hgrant0_p & v23f3a55;
assign v23fcdb6 = hbusreq6 & v230251b | !hbusreq6 & v84561b;
assign v230058a = hgrant1_p & v84564d | !hgrant1_p & !v23fcaf1;
assign v22fbab1 = hgrant4_p & v2308506 | !hgrant4_p & v2304c95;
assign v23f810b = hmaster0_p & v23fc81b | !hmaster0_p & v22eccfc;
assign bc87ee = hbusreq4_p & v23125a8 | !hbusreq4_p & v230e40c;
assign v23f6739 = hmaster2_p & v84561b | !hmaster2_p & v23fc7b2;
assign v22f0e00 = hbusreq1_p & v2306d29 | !hbusreq1_p & v23f4426;
assign v23fbb00 = hmaster0_p & v22f061c | !hmaster0_p & !v22ff315;
assign v23023aa = hmaster0_p & v22f50f0 | !hmaster0_p & v22f8c6b;
assign v2304965 = hmaster0_p & bd74cf | !hmaster0_p & v23f24d5;
assign v15070fa = hgrant1_p & v22ee956 | !hgrant1_p & v231140d;
assign v23fb57d = hgrant2_p & v2304074 | !hgrant2_p & v2302149;
assign v230f165 = hbusreq3_p & v22febe7 | !hbusreq3_p & v23fc02b;
assign v22fe2a8 = hbusreq3_p & v9526ac | !hbusreq3_p & v22f00c6;
assign v23124c5 = hmaster2_p & v230f9db | !hmaster2_p & !v84561b;
assign v23fbdb9 = hmaster2_p & v22ee281 | !hmaster2_p & v8f530a;
assign v2393116 = hlock2_p & b9d02f | !hlock2_p & v845620;
assign v23fc98c = hbusreq6 & v23fc320 | !hbusreq6 & v84561b;
assign v9d7c04 = hmaster0_p & v23fc442 | !hmaster0_p & v23f209f;
assign v22f606c = hmaster0_p & v22f8312 | !hmaster0_p & v23fbf94;
assign v22eea67 = hbusreq5_p & v22f4d69 | !hbusreq5_p & v23fbd94;
assign v23f4168 = hbusreq6_p & v22ff66a | !hbusreq6_p & bcc479;
assign v230d849 = hbusreq6_p & v2302f60 | !hbusreq6_p & v23fa950;
assign v22f8ad3 = hmaster2_p & v22fb0b7 | !hmaster2_p & v23fbf6c;
assign v22f316b = hbusreq5_p & v22fc5fd | !hbusreq5_p & v2300c80;
assign v191a964 = hbusreq3_p & v23fcfd3 | !hbusreq3_p & v23f56c3;
assign v22ec4d6 = hbusreq6 & v23f0178 | !hbusreq6 & !v22f05ac;
assign v23fc720 = hmaster1_p & v23fc966 | !hmaster1_p & v22edd9f;
assign v22f5d52 = hbusreq5_p & v230fab4 | !hbusreq5_p & v845620;
assign v2303199 = hmaster2_p & v22f5d52 | !hmaster2_p & v22f3b02;
assign v23f7659 = hmaster2_p & v23f86f0 | !hmaster2_p & v12cd3f4;
assign v2303102 = hmaster0_p & v23f1325 | !hmaster0_p & !v84561b;
assign v23f5055 = hgrant3_p & v230f1c8 | !hgrant3_p & v23fc2b8;
assign v2311a3e = hgrant1_p & a1fbc2 | !hgrant1_p & v2302167;
assign v191b155 = hbusreq0 & v230e9ea | !hbusreq0 & v23fbb10;
assign v22fbc47 = hmaster2_p & v23f0329 | !hmaster2_p & v2309c07;
assign v23f6215 = hmaster2_p & v23fc6c0 | !hmaster2_p & v22f7808;
assign v2305926 = stateG10_5_p & v22ef4ce | !stateG10_5_p & !v2309c8a;
assign v23f52c1 = hmaster2_p & v230d2c2 | !hmaster2_p & v23f58e5;
assign v23fba1d = hmaster1_p & v23f2849 | !hmaster1_p & v23fcbaa;
assign v22fe792 = hmaster2_p & v84561b | !hmaster2_p & !v23fb966;
assign v2300a5a = hbusreq5 & v23fc346 | !hbusreq5 & v84561b;
assign v22ff05e = hbusreq1_p & v22fcce6 | !hbusreq1_p & !v84561b;
assign v23fd014 = hgrant3_p & v23fc0a6 | !hgrant3_p & v2392ff0;
assign v22fe7ca = hmaster2_p & v22fe920 | !hmaster2_p & v23fb906;
assign v23fb5fa = stateG10_5_p & v22ed2f0 | !stateG10_5_p & v17a34ff;
assign v22efd02 = hgrant3_p & v84561b | !hgrant3_p & !v230da2f;
assign v1aad31a = hbusreq3_p & v231072a | !hbusreq3_p & v23f3c77;
assign v22fdbdb = hlock4_p & v230ccd6 | !hlock4_p & !v84563a;
assign v1506ffd = hbusreq5 & v23131e8 | !hbusreq5 & !v84561b;
assign v22efdb1 = hready & v84561b | !hready & !v23fca19;
assign v23f807d = hbusreq1_p & v106ae19 | !hbusreq1_p & b9d013;
assign v22f10c8 = hbusreq6 & v22fbc0e | !hbusreq6 & v23092cd;
assign v23fc117 = hgrant5_p & v23fc209 | !hgrant5_p & v23fb8fc;
assign v22eb338 = hbusreq3_p & v84562b | !hbusreq3_p & v22ffdd1;
assign v230ca2e = hbusreq2 & v23078cd | !hbusreq2 & v84561b;
assign v22f5216 = hbusreq4 & v23126b8 | !hbusreq4 & v84561b;
assign v23fccc5 = hbusreq6_p & v22f4507 | !hbusreq6_p & !v84561b;
assign v2307fee = hbusreq4 & v106af3a | !hbusreq4 & v22f2ca2;
assign v22ecc58 = hbusreq3_p & v23fbc40 | !hbusreq3_p & v23051cf;
assign v230c781 = hmaster2_p & v23fba93 | !hmaster2_p & v84561b;
assign v2393fc1 = hbusreq0_p & v1aae56f | !hbusreq0_p & v106ae21;
assign v22f2bc2 = hmaster0_p & v23fd051 | !hmaster0_p & v23fb7b2;
assign v23fbb9c = hbusreq6 & v22f09c4 | !hbusreq6 & v84561b;
assign v22f80ca = hburst0_p & v23fc116 | !hburst0_p & !v22fed4e;
assign v23f36a5 = hgrant0_p & v23133fa | !hgrant0_p & v23fc55f;
assign v93dace = hgrant5_p & v230439f | !hgrant5_p & v23fba08;
assign v231106e = hmaster2_p & v2308a4b | !hmaster2_p & v22f57e8;
assign v23fbba8 = hlock3_p & v22f41c0 | !hlock3_p & !v23fbf3e;
assign v2310516 = hbusreq1 & v22f8cb7 | !hbusreq1 & v84561b;
assign v23fcba1 = hmaster2_p & v8902b0 | !hmaster2_p & v230b27c;
assign v22fce73 = hbusreq1_p & v84561b | !hbusreq1_p & v22f1389;
assign v23115b1 = hbusreq6_p & v22f51b1 | !hbusreq6_p & v22ff79d;
assign v106ae87 = hmaster2_p & v22f071b | !hmaster2_p & !v23fcd0c;
assign v2308b4b = hbusreq1_p & v23fba24 | !hbusreq1_p & v23f6865;
assign v23fbba5 = hlock4_p & v23fb4af | !hlock4_p & v23f7b0a;
assign v23fc92d = hmaster0_p & v23130ea | !hmaster0_p & v13afad7;
assign v22eb711 = hbusreq4 & v230f0de | !hbusreq4 & v230aa7a;
assign v106ae3a = hbusreq4_p & v22fab90 | !hbusreq4_p & v22fdbbb;
assign v22f640a = hlock3_p & v2309282 | !hlock3_p & v84561b;
assign v22f0d4b = stateG10_5_p & v22fb71d | !stateG10_5_p & !v84561b;
assign v23fc164 = hgrant1_p & v84561b | !hgrant1_p & v230c579;
assign v230ff52 = hmaster0_p & v2312a90 | !hmaster0_p & v230f713;
assign v2310e89 = hgrant1_p & v84564d | !hgrant1_p & v2312351;
assign v22ee145 = hlock2_p & v23117af | !hlock2_p & v84564d;
assign v23fd051 = hgrant3_p & v23f56c0 | !hgrant3_p & v23fcbf3;
assign v23080ab = hbusreq5_p & v22ee956 | !hbusreq5_p & v23041c1;
assign v230bdb9 = hlock3_p & v22fb2c5 | !hlock3_p & v230105d;
assign v23f1228 = hbusreq5_p & v22f6f2b | !hbusreq5_p & !v22f654a;
assign v22f98d3 = hmaster0_p & v22f4989 | !hmaster0_p & !v230fe99;
assign v22f7ccb = hbusreq4_p & v2311027 | !hbusreq4_p & v2309c93;
assign v23f818e = jx1_p & v23fbedd | !jx1_p & v231016f;
assign v938878 = hgrant5_p & v2300c5c | !hgrant5_p & v15072af;
assign v2308331 = hmaster2_p & v22f1585 | !hmaster2_p & v2308765;
assign v230d30a = hbusreq5_p & v23f6bc1 | !hbusreq5_p & v23f4b28;
assign v23f7680 = hmaster2_p & v22f2718 | !hmaster2_p & v1aae087;
assign v23f567b = hmaster0_p & v22f1a14 | !hmaster0_p & v23f3eda;
assign v23fcfa4 = stateA1_p & v2302ca3 | !stateA1_p & v22f7078;
assign v230e635 = hmaster2_p & v22fa5fd | !hmaster2_p & v84561b;
assign v23fbfd9 = hbusreq0 & v22f03ce | !hbusreq0 & v84561b;
assign v23f74da = hbusreq6 & v23fc7e7 | !hbusreq6 & v2302131;
assign v23fc270 = hlock6_p & v230e44a | !hlock6_p & v23fcccb;
assign v2306bed = hbusreq3 & v23024ed | !hbusreq3 & !v84561b;
assign v22f9369 = stateA1_p & v2302ca3 | !stateA1_p & v23f6bf3;
assign v23fc7e8 = hmaster0_p & v22f2abb | !hmaster0_p & v2309cdc;
assign v2301be6 = hmaster2_p & v84561b | !hmaster2_p & v22eefaf;
assign v23fb21c = jx0_p & v23063de | !jx0_p & !v22f53a0;
assign v99a622 = hgrant3_p & v22f8e29 | !hgrant3_p & v23fc696;
assign v23fa1e7 = hbusreq6_p & v230e9f8 | !hbusreq6_p & v23fb935;
assign v23f7bc9 = hmaster2_p & v2302a4d | !hmaster2_p & !v22f4986;
assign v23f3978 = hbusreq2_p & v2304b4d | !hbusreq2_p & !v84561b;
assign v230124d = hbusreq4 & v12cd4c5 | !hbusreq4 & v84561b;
assign v22ee3ca = hbusreq6_p & v22ef499 | !hbusreq6_p & v23fce06;
assign v23fb215 = hlock0_p & v22fd30c | !hlock0_p & v22ff08f;
assign v23facb5 = jx2_p & v23fbfb7 | !jx2_p & v84561b;
assign v23fbfe0 = hgrant5_p & v23fc512 | !hgrant5_p & !v84561b;
assign v12cd920 = hbusreq1 & v22f9b5b | !hbusreq1 & v22f9f27;
assign v22fb653 = hmaster0_p & v23f4e63 | !hmaster0_p & v23006f8;
assign v23fcef8 = hmaster0_p & v2303fa0 | !hmaster0_p & v23f4007;
assign v22fc1be = stateG10_5_p & v22ee195 | !stateG10_5_p & v9526ac;
assign v2311ef7 = hbusreq3_p & v23f3c12 | !hbusreq3_p & v23fbe66;
assign v2304049 = hbusreq5 & v22edee1 | !hbusreq5 & v84561b;
assign v230d4d9 = hbusreq1_p & v2301d23 | !hbusreq1_p & v2309c93;
assign v22fbd0e = hmaster1_p & v23fbf13 | !hmaster1_p & v2301a76;
assign v23f65bb = hbusreq5_p & a1fbc2 | !hbusreq5_p & v22edba6;
assign v22ec330 = hbusreq3_p & v23f1e80 | !hbusreq3_p & v23fb550;
assign aacd54 = hmaster1_p & v22f9f2f | !hmaster1_p & v2310b15;
assign v22fa934 = hmaster2_p & v23fb67c | !hmaster2_p & !v230f34c;
assign v22f5c1a = hbusreq4_p & a8ec08 | !hbusreq4_p & v2302dca;
assign v23082ec = hbusreq0 & v22f925b | !hbusreq0 & v84561b;
assign v2305d6e = hbusreq3 & v22f4eeb | !hbusreq3 & v23fbd58;
assign v22f3b02 = hbusreq1_p & v22fafe5 | !hbusreq1_p & v845620;
assign v230a0ad = hmaster0_p & v22eb5a9 | !hmaster0_p & v106ae19;
assign v22f2d88 = jx2_p & v23fbc71 | !jx2_p & v2306d36;
assign v230d6b2 = hmaster0_p & v22f5b58 | !hmaster0_p & v22f0552;
assign v23fc63b = hgrant1_p & v23107b6 | !hgrant1_p & v23fc3dd;
assign v22fb442 = hmaster0_p & v2392e6c | !hmaster0_p & v23f0234;
assign v22f4d46 = hgrant0_p & v84561b | !hgrant0_p & v23fb59e;
assign v23f96d0 = hmaster2_p & v845620 | !hmaster2_p & v23fb7d1;
assign v22f0593 = hbusreq5_p & v230aa54 | !hbusreq5_p & v84561b;
assign v22f7752 = hbusreq1 & v2308d79 | !hbusreq1 & !v84561b;
assign v23f543d = hbusreq3_p & v23fba7c | !hbusreq3_p & v23f50bd;
assign v22faa21 = hlock0_p & v23094cb | !hlock0_p & !v84561b;
assign v22ef5cd = hgrant3_p & v22f52a4 | !hgrant3_p & v23f424b;
assign bee61a = hbusreq6_p & v23f1f36 | !hbusreq6_p & !v84561b;
assign v22f07fc = jx1_p & v85e5cf | !jx1_p & v23fc34a;
assign v23f240c = hbusreq4_p & v23fc787 | !hbusreq4_p & v84561b;
assign v23f4c57 = hbusreq1_p & v23064e4 | !hbusreq1_p & !v84561b;
assign v23fc6db = hbusreq3 & v22f7da7 | !hbusreq3 & v12cc30c;
assign v23f0dd4 = hmaster0_p & v2303bee | !hmaster0_p & v2312f81;
assign v23fb3a3 = hgrant3_p & v22ff969 | !hgrant3_p & v22f34c1;
assign v22f05ac = hmaster2_p & v23f75db | !hmaster2_p & v845636;
assign v23f333e = hmaster0_p & v23f67d3 | !hmaster0_p & v23fc908;
assign v2305071 = hlock1_p & v22f48a5 | !hlock1_p & v2304ec7;
assign v23fca20 = hmaster2_p & v22f4cf3 | !hmaster2_p & fc8ab7;
assign v23f7423 = hgrant3_p & v2309cdc | !hgrant3_p & v23f64db;
assign v23f9f07 = hgrant1_p & v845626 | !hgrant1_p & v23fc78b;
assign v23095df = hgrant3_p & v22ee657 | !hgrant3_p & v23051eb;
assign v23fcec2 = hbusreq5_p & v9932c2 | !hbusreq5_p & !v23fb540;
assign v23fb1b7 = hbusreq3_p & v23fb60e | !hbusreq3_p & v23f426b;
assign v2311d0c = hbusreq5_p & v23fba6b | !hbusreq5_p & v10dbf64;
assign bd8382 = hlock2_p & v230d7b7 | !hlock2_p & !v2304ec7;
assign bd7669 = hbusreq4_p & v22f9ca3 | !hbusreq4_p & v23fc1c0;
assign v22f082f = hbusreq3_p & v23fccbc | !hbusreq3_p & v23fbc96;
assign v22f227e = hmaster2_p & bdc4e2 | !hmaster2_p & v22ec89f;
assign v191b0a2 = hlock5_p & bbc337 | !hlock5_p & !v191b096;
assign v22fe8a4 = hmaster0_p & v23fbcfd | !hmaster0_p & !v2313394;
assign v23fc316 = hbusreq1_p & v22f78de | !hbusreq1_p & v2300cb6;
assign v23f8013 = hbusreq4 & v2301271 | !hbusreq4 & v22fe145;
assign v22f2ee3 = hbusreq4_p & v23fbc0c | !hbusreq4_p & v23f6723;
assign v22ed711 = hbusreq3_p & c20101 | !hbusreq3_p & v23fcc42;
assign bd3bb2 = hburst0_p & v22ed56a | !hburst0_p & !v22fdc60;
assign v23048df = hgrant2_p & v2312d11 | !hgrant2_p & v22f7f74;
assign v2305055 = hgrant5_p & v84561b | !hgrant5_p & v106a7a3;
assign v22f1f3f = hmaster2_p & v2304fe7 | !hmaster2_p & v22ffe8d;
assign ad06d5 = hbusreq6_p & v22f72ff | !hbusreq6_p & v23f6cc2;
assign v9052d9 = hbusreq5 & v230474b | !hbusreq5 & v84561b;
assign v2304962 = hgrant1_p & v84561b | !hgrant1_p & v22f23e7;
assign hgrant2 = !v12cc321;
assign v23fc9b2 = hmaster0_p & v23fce0b | !hmaster0_p & v22f2158;
assign v22ffb2b = hlock1_p & v230d109 | !hlock1_p & v99d709;
assign v23fc3b9 = jx1_p & v23091ce | !jx1_p & v2310e53;
assign v22f09ab = hgrant3_p & v22fba0e | !hgrant3_p & v23f425f;
assign v22fce06 = hbusreq0_p & v23fc14e | !hbusreq0_p & !v23fb669;
assign v23f20d3 = hmaster2_p & v230d2c2 | !hmaster2_p & v231033b;
assign v23fb64e = hgrant4_p & v2310047 | !hgrant4_p & v23050ee;
assign v2303d1d = hgrant2_p & v23fb410 | !hgrant2_p & v191a879;
assign v22ec9a7 = hbusreq5 & v13afe3a | !hbusreq5 & !v84561b;
assign v22fa7f7 = hbusreq5_p & v23faa52 | !hbusreq5_p & !v22f1553;
assign v9ae0d1 = hlock6_p & v2310a58 | !hlock6_p & v23fb0f3;
assign v23f9631 = hmaster2_p & v23f8f25 | !hmaster2_p & v23fca72;
assign v2392fa3 = hlock0_p & v84562a | !hlock0_p & v22eedf9;
assign v23fbb0f = hlock5_p & v84561b | !hlock5_p & v2391e51;
assign v22ee95f = hbusreq3 & v230cfc7 | !hbusreq3 & !v84561b;
assign v230c1e1 = hbusreq6_p & v22fb4a6 | !hbusreq6_p & v22ec1a8;
assign v22eb23c = hmaster0_p & v2308363 | !hmaster0_p & v23fc40a;
assign v22f78c3 = hbusreq3_p & v2302177 | !hbusreq3_p & !v23f946b;
assign v23fbb8f = hgrant3_p & v23fc60b | !hgrant3_p & v22efc28;
assign v123d721 = jx2_p & v22f30bb | !jx2_p & !v231029e;
assign a03e3a = hbusreq6_p & v23028be | !hbusreq6_p & v230201b;
assign v22eecbb = hbusreq3_p & v23fc083 | !hbusreq3_p & !v22ed598;
assign v22f0052 = hlock6_p & v23f8534 | !hlock6_p & !v84561b;
assign v23f68bf = hburst1 & v84561b | !hburst1 & v23fc2f3;
assign v23fc9b6 = hlock1_p & v23060eb | !hlock1_p & !v84561b;
assign v23fbf41 = hmaster0_p & v1aad69f | !hmaster0_p & v22f9ab1;
assign v23fc104 = hlock6_p & v22eaed2 | !hlock6_p & v84561b;
assign v2387c0f = jx3_p & v23fcf14 | !jx3_p & v22edccd;
assign v2302831 = hbusreq4 & v230b23c | !hbusreq4 & v84561b;
assign v22fa76f = hlock5_p & abf6b6 | !hlock5_p & bbc337;
assign v23f532f = hbusreq4 & v22f639a | !hbusreq4 & v22f475e;
assign v23fc92e = hbusreq6 & v23fa903 | !hbusreq6 & v845627;
assign v2303e9a = hgrant3_p & v23f5019 | !hgrant3_p & v23f447e;
assign v23f408c = hbusreq3 & v2306fb7 | !hbusreq3 & v84561b;
assign v22ef043 = hbusreq5 & v22ff315 | !hbusreq5 & v23fb966;
assign v1e84124 = hbusreq5_p & v22f6ba0 | !hbusreq5_p & !v22f9092;
assign v23083d6 = hbusreq1 & v22f4e0b | !hbusreq1 & v230f5a3;
assign v1506fa4 = hbusreq1_p & v23f6411 | !hbusreq1_p & !v106ae19;
assign v23fd018 = jx0_p & bd7b44 | !jx0_p & v23099b2;
assign v22f1713 = hmaster2_p & v22ffb12 | !hmaster2_p & v23fba9a;
assign v22f76c2 = hlock5_p & v23fbaf0 | !hlock5_p & !v84561b;
assign v1506a4d = hbusreq0 & v230358b | !hbusreq0 & v84561b;
assign v23fb189 = hready_p & v23f0f9a | !hready_p & v23fcb94;
assign v23fce7b = hbusreq3 & v23fc03c | !hbusreq3 & v84561b;
assign v22ee36d = hmaster0_p & v2301be6 | !hmaster0_p & v22eeb06;
assign v23f65ae = hlock0_p & v2391d40 | !hlock0_p & v22f2a24;
assign v23fba17 = hbusreq5_p & v22ede7f | !hbusreq5_p & v23f6b0f;
assign v22f30dc = hmaster0_p & v22f789c | !hmaster0_p & !v23f7632;
assign v230ccff = hmaster2_p & v23f2c05 | !hmaster2_p & !v23fa345;
assign v23028fa = hmaster0_p & v230e4da | !hmaster0_p & v23fce52;
assign v22f1f78 = hbusreq3_p & v23fc001 | !hbusreq3_p & v84561b;
assign v23f4f13 = hmaster2_p & v23fc393 | !hmaster2_p & v23f5cb3;
assign v22fd379 = hbusreq5_p & v23fc733 | !hbusreq5_p & !v23fc178;
assign v22ed83b = hbusreq3 & v230b68b | !hbusreq3 & v23fb2f8;
assign v23f9507 = hmaster2_p & v84561b | !hmaster2_p & !e1e73c;
assign v9b93b3 = hbusreq1_p & v22f56d2 | !hbusreq1_p & v230f63f;
assign v12cda32 = hbusreq5_p & v23fc947 | !hbusreq5_p & fc8c57;
assign v23fbb20 = hlock0_p & b5f51c | !hlock0_p & !v106ae19;
assign v22f01b2 = hbusreq6_p & v23f282d | !hbusreq6_p & v23fc8a9;
assign v230ec21 = stateA1_p & v23fc8d7 | !stateA1_p & !v22eced4;
assign v23fb591 = hbusreq1 & v23fcfb8 | !hbusreq1 & v22f5583;
assign v191b147 = hbusreq5_p & v22f4ab3 | !hbusreq5_p & v84561b;
assign v23091ef = hbusreq3 & v22f1de1 | !hbusreq3 & v22f8d38;
assign v23fc972 = hmaster2_p & v84561b | !hmaster2_p & v23f89f6;
assign v230562d = hbusreq4 & v23f942a | !hbusreq4 & v84561b;
assign v22f961e = hlock3_p & v230e45a | !hlock3_p & !v84561b;
assign v23fcbeb = hbusreq5_p & v23fc3f2 | !hbusreq5_p & v22f7929;
assign v22f6aa1 = hbusreq6 & v23f19ee | !hbusreq6 & v22f475e;
assign v22fa4dd = hmastlock_p & v23efe10 | !hmastlock_p & v84561b;
assign v2307578 = hlock3_p & v22f1f78 | !hlock3_p & v23fbd38;
assign v2392811 = jx1_p & v23fcb29 | !jx1_p & v23f5429;
assign v23fb5d7 = hbusreq4_p & v2312d71 | !hbusreq4_p & v22f83fd;
assign v22f4950 = jx1_p & v23f651e | !jx1_p & v22f244d;
assign v22f66cf = hgrant1_p & v22f8b43 | !hgrant1_p & v23f850a;
assign start = v2346bd3;
assign v22ec3c3 = hmaster2_p & v23fcdc9 | !hmaster2_p & !v23fcf70;
assign v2304009 = hbusreq2_p & v23f8089 | !hbusreq2_p & !v84561b;
assign v230fe8e = hgrant2_p & v23fc5f4 | !hgrant2_p & v84561b;
assign v23fc49b = hmaster2_p & v13affaa | !hmaster2_p & v23f6836;
assign v2311506 = hbusreq5_p & v22f56d2 | !hbusreq5_p & v23fb720;
assign v23fc67b = hgrant3_p & v22ff21b | !hgrant3_p & v23f3ab0;
assign v2307479 = hmaster1_p & v22f67fb | !hmaster1_p & v23f50dd;
assign v230de92 = hlock1_p & v23fc7f0 | !hlock1_p & v22fe300;
assign v23f6fed = hgrant3_p & v84561b | !hgrant3_p & e1e707;
assign v2391e8e = hbusreq4_p & v23fc063 | !hbusreq4_p & v22fb4d8;
assign v23fc888 = hmaster0_p & v23fc75d | !hmaster0_p & v231141f;
assign v23f62a8 = hmaster2_p & v2301a75 | !hmaster2_p & v22f5e91;
assign v22feb20 = hgrant1_p & v84561b | !hgrant1_p & v23f9ee2;
assign v23fce8e = hbusreq3_p & v2304bc1 | !hbusreq3_p & v22f4114;
assign a0e5e2 = hbusreq6_p & v23fca14 | !hbusreq6_p & v23fc50e;
assign v23fbcf8 = hgrant3_p & v22f368e | !hgrant3_p & v23fc676;
assign v2311dff = hbusreq5_p & v2306d29 | !hbusreq5_p & v23fcd3c;
assign v2392697 = hmaster0_p & v23fce0b | !hmaster0_p & v2309efb;
assign v23fb9dc = hbusreq2 & v23fbdb0 | !hbusreq2 & v84561b;
assign v23faa16 = hbusreq5_p & v22fc745 | !hbusreq5_p & v84562b;
assign v22eb4b3 = hmaster2_p & v845620 | !hmaster2_p & !v84561b;
assign v23f58f9 = hbusreq4 & v22f7144 | !hbusreq4 & v1aadf17;
assign v230c81f = hlock4_p & v23fcdfa | !hlock4_p & v84562b;
assign v23fbccc = hbusreq4_p & v22f1f9f | !hbusreq4_p & v84561b;
assign v22f04a6 = stateG10_5_p & v23fba61 | !stateG10_5_p & v2311810;
assign v23f7206 = hbusreq3_p & v23fbc6d | !hbusreq3_p & !v84561b;
assign v22f5521 = hmaster0_p & v230ed3d | !hmaster0_p & v230bb69;
assign v23fc5c6 = hmaster0_p & v22f063d | !hmaster0_p & v23f0d8a;
assign v23fcb56 = hbusreq3_p & v22faba5 | !hbusreq3_p & v23fcc9f;
assign v22edb96 = hbusreq6_p & v23fb7a3 | !hbusreq6_p & v23f664b;
assign bc96dd = hbusreq1_p & v23fbd53 | !hbusreq1_p & v84561b;
assign v22f71ca = hbusreq5_p & v230e311 | !hbusreq5_p & v23fd06a;
assign v23f42a6 = hmaster0_p & v22f3d79 | !hmaster0_p & a75533;
assign v23f4338 = hlock3_p & v2301e9a | !hlock3_p & v230129b;
assign v2308d5a = hmaster2_p & v22f3aa1 | !hmaster2_p & v22eec0e;
assign v23f5382 = hgrant3_p & v84561b | !hgrant3_p & v22eeff5;
assign v22ffa10 = hbusreq5_p & v23fbe0a | !hbusreq5_p & v230979f;
assign v22eb748 = hbusreq6_p & v23fc673 | !hbusreq6_p & v23fc04e;
assign v22f926d = hbusreq5_p & a8d315 | !hbusreq5_p & v84561b;
assign v22ed145 = hlock4_p & v23fb51a | !hlock4_p & v23f965d;
assign v230d5ab = hbusreq0 & v23fcf5c | !hbusreq0 & v1aadb95;
assign v23fc32e = hmaster1_p & v23fc6be | !hmaster1_p & !v23fb63e;
assign v2311606 = hbusreq1_p & v22f860b | !hbusreq1_p & v2309b39;
assign v2306fae = jx1_p & v23fbe06 | !jx1_p & v84561b;
assign v230d109 = hbusreq1 & v23003cc | !hbusreq1 & v84561b;
assign v12cc2f8 = hbusreq1_p & v23105cd | !hbusreq1_p & !v22f36ff;
assign v23021ec = hmaster0_p & v22fbde3 | !hmaster0_p & v23fbea2;
assign v22f08b7 = hgrant1_p & v2300827 | !hgrant1_p & v22f1403;
assign v22ef144 = hlock4_p & v22f7c2b | !hlock4_p & v22eaaa7;
assign v23fb5b3 = hmaster2_p & v84561b | !hmaster2_p & v845622;
assign v22f0552 = hmaster2_p & v23fcb69 | !hmaster2_p & v22ee956;
assign v23f4e8c = hbusreq5 & v230f5a3 | !hbusreq5 & v84561b;
assign b00ad2 = hbusreq2_p & v22f52c1 | !hbusreq2_p & v84561b;
assign v23f711a = hlock4_p & v84564d | !hlock4_p & !v84561b;
assign v23f4d58 = hlock5_p & v22fd8a6 | !hlock5_p & v84561b;
assign v22ee665 = hmaster0_p & v239174f | !hmaster0_p & v22fa987;
assign v12cd8ed = hbusreq4_p & v23f64dd | !hbusreq4_p & v23fbfd3;
assign v230e872 = hbusreq1 & v22ee281 | !hbusreq1 & v84561b;
assign v22eea08 = hmaster2_p & v23fbaaa | !hmaster2_p & v23fcae5;
assign v23fc4c0 = hbusreq5_p & v22fbeea | !hbusreq5_p & v23000cf;
assign v23fce86 = hbusreq0_p & v191a86f | !hbusreq0_p & !v191a879;
assign v23105eb = hbusreq3_p & v23fcae0 | !hbusreq3_p & v84561b;
assign v22ef998 = hmaster2_p & v22fe346 | !hmaster2_p & v22ffb12;
assign v23fce0d = hlock0_p & v22f2884 | !hlock0_p & v845620;
assign v23fa8d8 = hlock3_p & v2304ea9 | !hlock3_p & !v23f06d7;
assign c242c8 = jx0_p & v230e437 | !jx0_p & v23fc7a1;
assign v23fbfea = hbusreq5_p & v22fee46 | !hbusreq5_p & v12cd931;
assign v22fdc63 = hbusreq4_p & b0fc7a | !hbusreq4_p & v22efafa;
assign v22fbb54 = hgrant5_p & v23fbdb7 | !hgrant5_p & v23f3115;
assign v23fbfc3 = hmaster2_p & v23fb6e3 | !hmaster2_p & !v2312696;
assign v2301463 = hlock3_p & v23019f7 | !hlock3_p & !v23fc92f;
assign v23037ac = hgrant3_p & bd74e7 | !hgrant3_p & v22fafa5;
assign v230a180 = hbusreq2_p & b09503 | !hbusreq2_p & v84561b;
assign v230f94d = hbusreq4 & v23f9864 | !hbusreq4 & v22f3840;
assign v23fbc78 = hmaster2_p & v23f3ccf | !hmaster2_p & v23f4c57;
assign v230f9d5 = hbusreq3 & v22f60dd | !hbusreq3 & v84561b;
assign v2303bf6 = hmaster0_p & v23fb1b5 | !hmaster0_p & v239223a;
assign v2310f12 = hbusreq6_p & v23068bb | !hbusreq6_p & v22ec2c0;
assign v23fc096 = stateG10_5_p & v23052cc | !stateG10_5_p & v22efc50;
assign v23f3af2 = hmaster0_p & v23fb436 | !hmaster0_p & v23fc5ad;
assign v23f9545 = hbusreq0 & v13afe3a | !hbusreq0 & !v23fce22;
assign v22f7110 = hmaster2_p & b9d061 | !hmaster2_p & v22feae3;
assign v22fa8c6 = hgrant3_p & v84561b | !hgrant3_p & v22f9445;
assign v22fb22e = hmaster2_p & v231033b | !hmaster2_p & v2304990;
assign v22ef499 = hlock6_p & v22f37e8 | !hlock6_p & v2309840;
assign v23f460c = hmaster0_p & v22fb7ef | !hmaster0_p & a1fd9c;
assign v23051fc = hgrant3_p & v84561b | !hgrant3_p & v230322f;
assign v22fd106 = hgrant2_p & v23f4694 | !hgrant2_p & !v22f532c;
assign v22fa5f1 = hmaster0_p & v230f133 | !hmaster0_p & v2394087;
assign v23fa005 = hbusreq3 & v12ce4ac | !hbusreq3 & v22f88c3;
assign v22ff7ef = hgrant6_p & v23122b0 | !hgrant6_p & v22faa7a;
assign v23f0ce0 = hready & v22fbf54 | !hready & !v84561b;
assign v2307150 = hlock0_p & v1aae56f | !hlock0_p & v2393fc1;
assign v22eb7cc = hmaster1_p & v23f493a | !hmaster1_p & v85b90c;
assign v23f6710 = hbusreq4_p & v22f484b | !hbusreq4_p & v22f9a8b;
assign v12cd9c9 = hgrant0_p & v22f9acf | !hgrant0_p & v2302d1f;
assign v23fc799 = hgrant5_p & b9eb75 | !hgrant5_p & v2301f92;
assign v230561d = hlock2_p & v2312ea7 | !hlock2_p & v845620;
assign v23f5cd7 = hbusreq4_p & v9cf5cf | !hbusreq4_p & v23fc80c;
assign v230ee35 = hgrant5_p & v2392fbd | !hgrant5_p & !v22f5fb8;
assign v22f847c = hbusreq6_p & v23fb495 | !hbusreq6_p & v22ed55a;
assign v2307b9c = hbusreq3_p & v23fcb3c | !hbusreq3_p & v2305a05;
assign v23fc18b = hbusreq3_p & v9c8a7f | !hbusreq3_p & v22fc1e9;
assign v23045e7 = hgrant2_p & v23f1227 | !hgrant2_p & v22f0326;
assign v22f7634 = hgrant1_p & v22f1427 | !hgrant1_p & v23f8884;
assign v22fc34e = hbusreq2_p & v22ed85a | !hbusreq2_p & v84564d;
assign v2301dad = hbusreq4_p & v2310852 | !hbusreq4_p & v23fc15b;
assign v15074df = hbusreq0_p & v2304ed3 | !hbusreq0_p & v845629;
assign v2304536 = hlock0_p & v230d32d | !hlock0_p & v230d529;
assign v22ed127 = hbusreq5 & v23f3115 | !hbusreq5 & !v84561b;
assign v230a709 = hmaster2_p & v23f5f5f | !hmaster2_p & !v2309cdc;
assign v23fbb3e = hbusreq0 & v23fc926 | !hbusreq0 & v84561b;
assign v2308110 = hbusreq1_p & v22f98e3 | !hbusreq1_p & v22fe37c;
assign v22f36c5 = hmaster2_p & v22f1585 | !hmaster2_p & v22ff1dd;
assign v23fa7ba = hgrant3_p & v84561b | !hgrant3_p & v2305841;
assign v23028be = hmaster0_p & v2311524 | !hmaster0_p & b72216;
assign v23f14e6 = hbusreq1 & v22fe37c | !hbusreq1 & v23fcbeb;
assign v23fce98 = hbusreq0_p & v84561b | !hbusreq0_p & v22f1992;
assign v22ed12a = hmaster0_p & v239174f | !hmaster0_p & v22fde18;
assign v22f969f = hlock3_p & v23f022a | !hlock3_p & v22f9b0c;
assign v23fc91a = hbusreq6 & v22fc945 | !hbusreq6 & !v230aa2f;
assign v23021b9 = hmaster2_p & v22fb77d | !hmaster2_p & v22fc5f0;
assign v1aad815 = hbusreq1_p & v230fdd7 | !hbusreq1_p & v22ec745;
assign v230a70a = hmaster2_p & v23fc969 | !hmaster2_p & v845620;
assign v2308aa9 = hbusreq4_p & v23fb21a | !hbusreq4_p & v23f6114;
assign v230cb83 = hmaster1_p & v2302b5b | !hmaster1_p & !v23f49cd;
assign v1aadb45 = hbusreq6_p & v230e779 | !hbusreq6_p & v22ff6ba;
assign v23124cc = hbusreq2_p & v22edcfc | !hbusreq2_p & v84561b;
assign v22eb6ee = stateG10_5_p & v8ebd5d | !stateG10_5_p & v22f0945;
assign v22efc3c = hbusreq2 & v23fb1a4 | !hbusreq2 & !v84561b;
assign v2310eb6 = hbusreq5_p & v1506fbf | !hbusreq5_p & v84561b;
assign v191b1ba = hmaster2_p & v23f445f | !hmaster2_p & v2310108;
assign v23024ed = hmaster2_p & v84561b | !hmaster2_p & !v230c876;
assign v23014b0 = hmaster0_p & v23034c9 | !hmaster0_p & v23fc0a5;
assign v15070ca = hgrant1_p & v84561b | !hgrant1_p & v23fb0c9;
assign v23f209f = hbusreq4 & v23fcb67 | !hbusreq4 & !v845636;
assign v22fe052 = hgrant3_p & v23fc75d | !hgrant3_p & v23fbee2;
assign v23fbbcb = hbusreq3_p & ba1576 | !hbusreq3_p & v22f61d2;
assign v230a2bd = hlock2_p & v13affaa | !hlock2_p & v84564d;
assign v917514 = hbusreq3_p & v22f2bab | !hbusreq3_p & v22f5d84;
assign v230d70b = hmastlock_p & v22f63e8 | !hmastlock_p & !v22eeaaf;
assign v2392ec8 = hready_p & v23fb47d | !hready_p & v23fab81;
assign v22f7988 = jx1_p & v23047dd | !jx1_p & v22f664f;
assign v23fbf1c = hmaster2_p & v84564d | !hmaster2_p & v230f5a3;
assign v23f740f = hbusreq3_p & v22fdfdd | !hbusreq3_p & v2303811;
assign v12cd3e7 = hmaster2_p & v22fd0e6 | !hmaster2_p & v23fbab0;
assign v22fe96a = hgrant1_p & v230522a | !hgrant1_p & v23f8cd3;
assign v2306257 = hgrant0_p & v23133fa | !hgrant0_p & v23ef8ef;
assign v23f7024 = hmaster2_p & v13afe3a | !hmaster2_p & v2304009;
assign v22eb397 = hbusreq6_p & v23105ac | !hbusreq6_p & v97b313;
assign v22eddc0 = hmaster0_p & v22f09fe | !hmaster0_p & v22f092c;
assign v23035ba = hbusreq0_p & v22eb659 | !hbusreq0_p & v84561b;
assign v23fb132 = hgrant3_p & v2346b41 | !hgrant3_p & v23011c7;
assign v2311358 = hmaster0_p & v22f336f | !hmaster0_p & !v22ebb51;
assign v23fbb53 = hmaster0_p & v22fa819 | !hmaster0_p & v22fcd80;
assign v22f3dea = hmaster0_p & v23fc5d4 | !hmaster0_p & v22ff4aa;
assign v1aad671 = jx0_p & v22f324c | !jx0_p & !v23f623e;
assign v2393f41 = hbusreq1 & v23fbee9 | !hbusreq1 & v23fb8e7;
assign v2301e43 = hmaster2_p & v1aae56f | !hmaster2_p & v23f6836;
assign v2300c23 = hbusreq4_p & v2304965 | !hbusreq4_p & v23fc029;
assign v23fc2f6 = hmaster0_p & v23fc77d | !hmaster0_p & v23fb964;
assign v22f4642 = hbusreq6 & v23fc3a4 | !hbusreq6 & v2304d7a;
assign v22f5076 = hmaster0_p & v23f54f7 | !hmaster0_p & bd7497;
assign v22f4d17 = hbusreq6 & v22ecaeb | !hbusreq6 & v22f88bb;
assign v2308980 = jx1_p & v22fcf35 | !jx1_p & v230cb83;
assign fc8fd5 = hgrant3_p & v22f91a8 | !hgrant3_p & v12cc6e0;
assign v23050c3 = hbusreq4 & v22f5840 | !hbusreq4 & v22fd533;
assign b67ed5 = hmaster2_p & v2313247 | !hmaster2_p & v23fb1c1;
assign v23f87b7 = hlock0_p & v22eed4c | !hlock0_p & !v845622;
assign v12cd9b5 = hbusreq6_p & v22f3068 | !hbusreq6_p & d97946;
assign v2310c11 = hmaster2_p & v106ae1c | !hmaster2_p & v22edc8d;
assign v23fbd90 = hbusreq3 & v2312cc9 | !hbusreq3 & v23f4fcd;
assign v2304432 = hbusreq6 & v230f795 | !hbusreq6 & v84561b;
assign v23fca36 = hbusreq1 & v2300b4f | !hbusreq1 & v230c52a;
assign v22f1d8b = hbusreq1 & v22ed85a | !hbusreq1 & v84561b;
assign v22f658c = jx3_p & v84561b | !jx3_p & v2308ef6;
assign v23fb0bb = hmaster2_p & v22f0945 | !hmaster2_p & v84561b;
assign v22f426a = hbusreq5_p & b9ca3d | !hbusreq5_p & !v84561b;
assign v23fccb3 = hbusreq6 & v23f5aa7 | !hbusreq6 & v84561b;
assign v22fa68b = hmaster2_p & v22f4527 | !hmaster2_p & !v84561b;
assign v23fb992 = hgrant5_p & v23fc225 | !hgrant5_p & !v191b04d;
assign v22fe552 = hgrant5_p & v230d25c | !hgrant5_p & !v84561b;
assign v23fbc6a = hgrant3_p & a4c16b | !hgrant3_p & v23f30b2;
assign v22f1963 = hmaster2_p & v22f0c59 | !hmaster2_p & v845627;
assign v22fb3c8 = hmaster1_p & v23fbf13 | !hmaster1_p & v2392023;
assign v2311bc4 = hbusreq3 & v23f4fbf | !hbusreq3 & v23fc988;
assign v230a9eb = hbusreq2_p & v23f6411 | !hbusreq2_p & !b9d013;
assign v22fc564 = hbusreq1_p & v23fc3f2 | !hbusreq1_p & v23fcbeb;
assign v23fc686 = hlock0_p & v84561b | !hlock0_p & v23fc73e;
assign v23ef987 = hmaster0_p & v23fa7ba | !hmaster0_p & v22fb151;
assign v23f3fb6 = hbusreq3_p & v2307d7f | !hbusreq3_p & !v84561b;
assign v231256a = hmaster2_p & v22f1244 | !hmaster2_p & v23fc04a;
assign v23fbd34 = hbusreq3_p & v22ffea6 | !hbusreq3_p & v23f660f;
assign v23fca63 = hbusreq6 & v23f90bc | !hbusreq6 & v845645;
assign v230a15d = hbusreq4_p & v22fa23d | !hbusreq4_p & v845637;
assign v22ed5fd = hbusreq3 & v191abee | !hbusreq3 & bfb87c;
assign v85bd38 = hbusreq5 & v2311255 | !hbusreq5 & v84561b;
assign v23fcb28 = hmaster2_p & v845629 | !hmaster2_p & !v84561b;
assign v230ae4f = hbusreq3_p & v8819d8 | !hbusreq3_p & v230159e;
assign v23facd7 = hbusreq3_p & v23fa005 | !hbusreq3_p & v23fbe76;
assign v23f0b74 = hbusreq4_p & v9d0518 | !hbusreq4_p & v23f60ba;
assign v22fd1a7 = hmaster2_p & v23fbe39 | !hmaster2_p & !v22f1ae5;
assign v230e509 = hbusreq5 & v23128a1 | !hbusreq5 & v84561b;
assign v23fc842 = hgrant2_p & v23fbbc7 | !hgrant2_p & v84564d;
assign v23f75e9 = hgrant5_p & v23fcbab | !hgrant5_p & v13afa38;
assign v22f0810 = hlock2_p & v22f037a | !hlock2_p & !v84561b;
assign v23f9033 = hgrant3_p & v84561b | !hgrant3_p & v23fbe0b;
assign b9c9ef = hlock0_p & v23f60ef | !hlock0_p & v23f039f;
assign v1aadad9 = hmaster2_p & v22f17ca | !hmaster2_p & v2304990;
assign v23f1cc0 = hmaster1_p & v22fbdcf | !hmaster1_p & v23108cb;
assign v230f14b = hlock3_p & v2309e57 | !hlock3_p & v2304bc1;
assign v230630c = hlock3_p & bd74c6 | !hlock3_p & v84562b;
assign v106ae43 = hready & v22f9527 | !hready & !v84561b;
assign v22f88f9 = hbusreq6_p & v22ed674 | !hbusreq6_p & v1506ec2;
assign v23fcca7 = hbusreq6_p & v95fb82 | !hbusreq6_p & v22f1259;
assign v23fb5a1 = hgrant1_p & v23fa2ec | !hgrant1_p & v23fcd4a;
assign v230859e = hmaster2_p & v22f5242 | !hmaster2_p & b50a75;
assign v23089a5 = hmaster2_p & v22f8c70 | !hmaster2_p & v22fe71e;
assign v230330a = hbusreq5 & v84561b | !hbusreq5 & fc8ab7;
assign v23f21c1 = hmaster2_p & v23fce6b | !hmaster2_p & v84561b;
assign v23fbcaa = hbusreq3 & v22eb4b3 | !hbusreq3 & v23fba11;
assign v22f0acc = hmaster0_p & v23027b1 | !hmaster0_p & v23fbb28;
assign v23fbd92 = hbusreq4_p & abf9f6 | !hbusreq4_p & v23fcb80;
assign v23fcbfb = hgrant3_p & v23fc3e8 | !hgrant3_p & adc67b;
assign v23fc60e = hmaster1_p & v23f437d | !hmaster1_p & v23fba0a;
assign v22f7289 = jx3_p & v23075bd | !jx3_p & v23f3ac8;
assign v23057e6 = hgrant5_p & v23fcc1f | !hgrant5_p & v23fbfe4;
assign v22efcbf = jx1_p & v2307fb2 | !jx1_p & v23f7ba2;
assign v23fb8c9 = hmaster0_p & baa026 | !hmaster0_p & v22f52a4;
assign v23f266b = hbusreq3_p & v2310bdf | !hbusreq3_p & v23fac5a;
assign v23920d8 = hgrant0_p & v23f0135 | !hgrant0_p & v84561b;
assign v23021af = hbusreq3_p & v23f7698 | !hbusreq3_p & !v84561b;
assign v95aaca = hbusreq4 & v22f6741 | !hbusreq4 & v84561b;
assign v23f1d8b = hgrant0_p & v23fa75a | !hgrant0_p & v23048df;
assign v230a5f5 = hbusreq4_p & v23fcabe | !hbusreq4_p & v22f0ad8;
assign v22fb8df = hbusreq5_p & v23fc904 | !hbusreq5_p & !v23067ba;
assign v22eb659 = hbusreq0 & v22f3643 | !hbusreq0 & v84561b;
assign v22fd7dd = hready & v22fa2de | !hready & v230d7b7;
assign v23f46ba = stateG10_5_p & v23fd03b | !stateG10_5_p & v23f5af5;
assign v22edc14 = hmaster0_p & v23107f5 | !hmaster0_p & v22f4b91;
assign v22fb49d = hmaster2_p & v23fc362 | !hmaster2_p & v23fb175;
assign v22f411f = hgrant1_p & v84561b | !hgrant1_p & v230a2bb;
assign v22f0b42 = hgrant1_p & v84561b | !hgrant1_p & !v22f135c;
assign v23f66a4 = hbusreq5_p & v84564d | !hbusreq5_p & v2302e87;
assign v22f9248 = hbusreq5_p & v22fb3c1 | !hbusreq5_p & v23f40ba;
assign v22f654e = hbusreq0 & v22f3959 | !hbusreq0 & !v84561b;
assign stateG10_1 = !v17cf286;
assign v230c6eb = stateG10_5_p & v22f69cc | !stateG10_5_p & v2301511;
assign v23fa23d = hbusreq3_p & v230e41f | !hbusreq3_p & v84561b;
assign v230dec9 = hmaster0_p & v23f76a5 | !hmaster0_p & !v230df28;
assign v230bb08 = hlock3_p & v23f8529 | !hlock3_p & v23094b2;
assign v22fc690 = hmaster1_p & v22fe315 | !hmaster1_p & v2308bfc;
assign v23fd067 = hbusreq5 & v2308e63 | !hbusreq5 & !v84561b;
assign v2307ffd = hmaster1_p & v22fa4a3 | !hmaster1_p & v23fd00e;
assign v230e80e = hmaster0_p & v23139e3 | !hmaster0_p & v23f6949;
assign v23fcecb = hbusreq3 & v23f4a02 | !hbusreq3 & !v84561b;
assign v84562e = hbusreq3 & v84561b | !hbusreq3 & !v84561b;
assign v22fd86e = hbusreq2 & v23fbfd0 | !hbusreq2 & v84561b;
assign v230fe27 = hmaster2_p & v191a86f | !hmaster2_p & v231228e;
assign v2310d1e = jx1_p & v23fc678 | !jx1_p & v23f9812;
assign v230c5ea = hbusreq1_p & v2306494 | !hbusreq1_p & v23f6ac5;
assign v23fb787 = hmaster0_p & v22ede34 | !hmaster0_p & v22fe392;
assign v23f4937 = hmaster0_p & v22ef4f0 | !hmaster0_p & !v2301a6d;
assign v22f8012 = hlock3_p & v23028f6 | !hlock3_p & v23fc99a;
assign v845622 = hbusreq0 & v84561b | !hbusreq0 & !v84561b;
assign v23fb314 = hbusreq0_p & v84561b | !hbusreq0_p & v23fa8bb;
assign v23fc265 = hbusreq0 & v23f8364 | !hbusreq0 & !v84561b;
assign v23fce29 = hbusreq6_p & v230a15d | !hbusreq6_p & v2302943;
assign v22f7e7a = hmaster2_p & v84562a | !hmaster2_p & v22f4527;
assign v2303507 = hmaster0_p & v22f2564 | !hmaster0_p & v23fbb5b;
assign v230ffae = hbusreq1_p & v23fb555 | !hbusreq1_p & !v84561b;
assign v230ff7d = hgrant1_p & v22eafb2 | !hgrant1_p & v230db14;
assign v22f4e64 = hmaster2_p & v23f80c1 | !hmaster2_p & v84561b;
assign v23f70c6 = hbusreq3 & v23f9c7f | !hbusreq3 & v23f9666;
assign v230ff63 = hbusreq5_p & v15071a5 | !hbusreq5_p & !v23fbde8;
assign v23f36e9 = hmaster2_p & v2309d55 | !hmaster2_p & v22fc13d;
assign v22edc85 = hbusreq6 & v23fbe8e | !hbusreq6 & v22ed5a5;
assign v230ba85 = hbusreq3 & v22ff3d1 | !hbusreq3 & v23fbc78;
assign v22ef810 = hlock1_p & v22fc42e | !hlock1_p & v84564d;
assign v23f1e38 = hbusreq6 & v22f8ad3 | !hbusreq6 & v22f5583;
assign v2306798 = hready_p & v22fa63e | !hready_p & v23fc0eb;
assign v22f176d = hmaster2_p & v22f61b6 | !hmaster2_p & v22ec894;
assign v23fac2d = hgrant3_p & v2346b41 | !hgrant3_p & v22fcad1;
assign f4067f = hmastlock_p & v23fc8a3 | !hmastlock_p & !v84561b;
assign v23fa0bf = hlock1_p & v191ad59 | !hlock1_p & !v84561b;
assign v23fcfa6 = hlock1_p & v23068a9 | !hlock1_p & v84561b;
assign v2310e81 = hgrant1_p & v23f646e | !hgrant1_p & v2303516;
assign v22f0d8d = hlock2_p & v22f1389 | !hlock2_p & v1aae087;
assign v23f710d = hbusreq4_p & v22fe362 | !hbusreq4_p & v84561b;
assign v22f4638 = hbusreq1_p & v230bd05 | !hbusreq1_p & v23fbbbd;
assign v22f366a = hgrant2_p & v2305fe0 | !hgrant2_p & !v84561b;
assign v23fc974 = hbusreq0 & v22f1389 | !hbusreq0 & v84561b;
assign v22f91f3 = stateG2_p & v23023b3 | !stateG2_p & !v22f349a;
assign v22f991d = hbusreq1_p & v23f8c22 | !hbusreq1_p & v84561b;
assign v22ec96a = hbusreq3_p & v22ecbb2 | !hbusreq3_p & v84561b;
assign v22f4700 = hlock0_p & v84561b | !hlock0_p & v230037d;
assign v230339f = hmaster0_p & v2312f45 | !hmaster0_p & v23fb5ee;
assign a5d081 = hbusreq1_p & v23f0bd2 | !hbusreq1_p & v23fc98a;
assign v23fc8d8 = hmaster2_p & v2312696 | !hmaster2_p & a39dae;
assign v22ee703 = hgrant1_p & v845626 | !hgrant1_p & b0df38;
assign v230c2ff = hmaster2_p & v23fa2ec | !hmaster2_p & v2305a12;
assign v2311027 = hlock4_p & v23fc390 | !hlock4_p & v2309c93;
assign v22ebedc = stateG10_5_p & v22f7f74 | !stateG10_5_p & v191a876;
assign v22f9d85 = hbusreq2 & v8b7fb1 | !hbusreq2 & v84562b;
assign v22f336f = hbusreq3_p & v230ba85 | !hbusreq3_p & v23fcc95;
assign v23fbddb = hgrant5_p & v23f7372 | !hgrant5_p & v230e07e;
assign v2312ac8 = hbusreq4 & v22f36c5 | !hbusreq4 & v23f44d0;
assign v2312c77 = hgrant1_p & v84561b | !hgrant1_p & v2306f84;
assign v23f5caf = hbusreq5_p & v23fb960 | !hbusreq5_p & v22f6372;
assign v2310782 = hmaster2_p & v23fab18 | !hmaster2_p & v84561b;
assign v23f85d7 = hbusreq1 & v13afe3a | !hbusreq1 & !v23fce22;
assign v2387c09 = hgrant1_p & v22f80b4 | !hgrant1_p & v22f0d2b;
assign v2309b3e = hbusreq1 & v2312912 | !hbusreq1 & v2391eaa;
assign v23f688e = hlock1_p & b5f51c | !hlock1_p & !v106ae19;
assign v22f0e5e = hbusreq5_p & v13afa38 | !hbusreq5_p & v22f7cab;
assign v23126fc = hgrant1_p & v84561b | !hgrant1_p & v23086c5;
assign v22fcf5b = hbusreq1_p & v23fb99b | !hbusreq1_p & v845620;
assign v23fc29b = hbusreq6_p & v23fcf62 | !hbusreq6_p & !v23f95bd;
assign v230abf3 = hlock0_p & v22f6a6b | !hlock0_p & v22fced7;
assign v2306bf9 = hgrant5_p & v84561b | !hgrant5_p & v22f0360;
assign v22fb29c = hmaster2_p & v22f0acd | !hmaster2_p & v2303a76;
assign v22f5cd9 = hbusreq6_p & v22ee142 | !hbusreq6_p & v23066bc;
assign v22fb631 = jx1_p & v23f8294 | !jx1_p & v22f70bf;
assign v230b750 = hbusreq5_p & v22f3643 | !hbusreq5_p & v2305684;
assign v23fcafe = hgrant0_p & v23133fa | !hgrant0_p & v22f7e80;
assign v23fc403 = jx0_p & v23fb522 | !jx0_p & v8eb4b5;
assign v23fb965 = hmaster0_p & v22f3b15 | !hmaster0_p & !v22f2005;
assign v22f6090 = hbusreq5_p & v84561b | !hbusreq5_p & v22f4d68;
assign v2312679 = hgrant3_p & v230b3ec | !hgrant3_p & v23f07f9;
assign v23f8fd0 = hmaster0_p & v22eec11 | !hmaster0_p & v22f9340;
assign v2301bdb = hmaster2_p & v84561b | !hmaster2_p & v2313118;
assign v22fa819 = hgrant3_p & v84561b | !hgrant3_p & !v22f57d4;
assign v23f8638 = hbusreq0 & v23131e8 | !hbusreq0 & v2306220;
assign v22fd799 = hmaster2_p & v23f55ea | !hmaster2_p & !v23fb029;
assign v22f2822 = hbusreq1 & v23f1207 | !hbusreq1 & b6f86d;
assign v23fc017 = hlock0_p & v191b0e4 | !hlock0_p & v2306885;
assign v2305ee5 = hbusreq3 & v23045f5 | !hbusreq3 & v84561b;
assign v2394087 = hbusreq3_p & v22ff21b | !hbusreq3_p & v23fc20d;
assign v23fb861 = hmastlock_p & v845667 | !hmastlock_p & !v84561b;
assign v230af72 = hbusreq5 & v2302e32 | !hbusreq5 & !v84561b;
assign a1ff0e = hbusreq3_p & v2382e8c | !hbusreq3_p & !v106ae19;
assign v23fb952 = hgrant5_p & v230b750 | !hgrant5_p & v1e84012;
assign v23fcae5 = hgrant1_p & v22ee956 | !hgrant1_p & v22fa155;
assign v22fcfee = jx2_p & v23f1328 | !jx2_p & v23f712d;
assign v22fc398 = hmaster0_p & v2302177 | !hmaster0_p & v13afb18;
assign v23f52f2 = hmaster0_p & v22ec354 | !hmaster0_p & v22f7ec9;
assign v23916fa = stateG10_5_p & v23f4eb4 | !stateG10_5_p & !v2310283;
assign v230d664 = hbusreq3_p & v230e932 | !hbusreq3_p & v23130d6;
assign v22ed4c6 = hbusreq1 & v22f5a08 | !hbusreq1 & v84561b;
assign v23f836b = hbusreq4 & b9c9cc | !hbusreq4 & v84561b;
assign v1507246 = hmaster1_p & v2305992 | !hmaster1_p & v23fc03d;
assign v23fcba3 = hgrant1_p & v84561b | !hgrant1_p & v2392d14;
assign v23fc7df = hlock2_p & v23f5af5 | !hlock2_p & !v2309c8a;
assign v23f1a4c = hmaster0_p & v23f1a14 | !hmaster0_p & v23094f0;
assign v23065e7 = hgrant3_p & b00ac7 | !hgrant3_p & v2393b99;
assign v22fdc80 = hmaster2_p & v22f7b47 | !hmaster2_p & v84561b;
assign v230adb7 = hmaster2_p & v23fbfd0 | !hmaster2_p & v23fc023;
assign v230c58d = hbusreq2_p & v23f95e1 | !hbusreq2_p & !v84561b;
assign v23fc277 = hbusreq3_p & v23fced1 | !hbusreq3_p & v22f2ed0;
assign v2302f63 = hlock3_p & bd837d | !hlock3_p & v2303cd6;
assign v2393495 = hbusreq4 & v1aadad9 | !hbusreq4 & v2310d04;
assign v23f67bd = hgrant0_p & v23fc246 | !hgrant0_p & !v23064ae;
assign v22fcea3 = hmaster0_p & v23f58bb | !hmaster0_p & a9c602;
assign v23fb41a = hbusreq3_p & v22ecf6c | !hbusreq3_p & !v84561b;
assign v22f768b = hgrant1_p & v22f86f3 | !hgrant1_p & !v22ec686;
assign v22f50f0 = hbusreq6 & v23f2843 | !hbusreq6 & a7dd55;
assign v23fbf17 = hgrant3_p & v23029bb | !hgrant3_p & v23fc6a8;
assign v23f65b4 = locked_p & v22fb157 | !locked_p & v191a86f;
assign v22f6f2b = hlock5_p & v23efc03 | !hlock5_p & v23f12fa;
assign v23fc25e = hbusreq3 & b9c9cc | !hbusreq3 & v84561b;
assign v2391f3b = hburst0 & v84561b | !hburst0 & !v22ec1cb;
assign v23fb0f0 = hbusreq3_p & v23fce88 | !hbusreq3_p & v23025e4;
assign v12cd4be = hmaster2_p & v230c727 | !hmaster2_p & v231007b;
assign v22ff982 = hlock3_p & v2306728 | !hlock3_p & !v84561b;
assign v23faece = hgrant5_p & v23fcd81 | !hgrant5_p & v230b52c;
assign v23fbb11 = hlock2_p & v22eda43 | !hlock2_p & v23fb581;
assign v23fb90b = hmaster0_p & v23fb8f3 | !hmaster0_p & v84561b;
assign v23fb505 = hgrant5_p & v84561b | !hgrant5_p & v22fa771;
assign v22f71ee = hbusreq3_p & v23fbb9d | !hbusreq3_p & v84561b;
assign v2303f37 = hbusreq1_p & v2392c41 | !hbusreq1_p & v23f99cf;
assign v22f128d = hbusreq3 & v23fcf88 | !hbusreq3 & v23002bf;
assign v22f56a5 = hlock3_p & v23fc8ba | !hlock3_p & v23f8d79;
assign v23fca75 = hbusreq5_p & v22eb32b | !hbusreq5_p & !v84561b;
assign v2304452 = hbusreq4 & v23fbcce | !hbusreq4 & v84561b;
assign v23119e0 = hburst1_p & v22f4e3c | !hburst1_p & v84561b;
assign v2312f45 = hgrant3_p & v23fc0d8 | !hgrant3_p & v23fbaa8;
assign v22f28d6 = hlock1_p & v23027c2 | !hlock1_p & v2305568;
assign v23030fc = hbusreq1_p & v23126de | !hbusreq1_p & v84561b;
assign v22fe0c1 = hlock5_p & v84561b | !hlock5_p & v23fba09;
assign v230b93b = hlock6_p & v23fbba0 | !hlock6_p & !v23fcae1;
assign bd77c5 = hbusreq6_p & b535c6 | !hbusreq6_p & b00a55;
assign v22f0323 = hbusreq5_p & v22f3643 | !hbusreq5_p & v23fbfcf;
assign v23f7f9d = hbusreq6 & v23008e6 | !hbusreq6 & !v84562e;
assign v23105cd = hready & v22f587e | !hready & v84561b;
assign v23fb6cf = hbusreq1_p & v22fc61a | !hbusreq1_p & v22fdc74;
assign v23f6ec6 = hmaster1_p & v15071f7 | !hmaster1_p & !v23f49cd;
assign v23fcf5d = hbusreq3 & v22f3643 | !hbusreq3 & v84561b;
assign v23fc917 = jx3_p & v23fbd51 | !jx3_p & v23faa11;
assign v239313a = hbusreq3_p & v2391e0c | !hbusreq3_p & v230a226;
assign v23f7997 = hbusreq6 & v2311568 | !hbusreq6 & v22fb3f4;
assign v23130f6 = hbusreq6_p & v2308164 | !hbusreq6_p & v23fcc68;
assign v2300b33 = jx1_p & v2309bda | !jx1_p & v23f83af;
assign v23fc956 = hbusreq3_p & v230ed85 | !hbusreq3_p & v230216e;
assign v23fbdd8 = hgrant3_p & v22f7dbc | !hgrant3_p & v23126b1;
assign v22f6397 = hbusreq5 & v1aad5ad | !hbusreq5 & v2312775;
assign v23fb81f = hbusreq3 & v23fb1fc | !hbusreq3 & v22fab50;
assign v23fc249 = stateA1_p & v2305aa1 | !stateA1_p & !v845649;
assign v23f957f = hbusreq6_p & v22f583d | !hbusreq6_p & v23083ee;
assign bd7535 = hmaster1_p & v23fc944 | !hmaster1_p & v2305c43;
assign v22fe940 = hgrant1_p & v23fb6ff | !hgrant1_p & v22f1393;
assign v22edbe0 = hlock5_p & v8ebd5d | !hlock5_p & v15070f7;
assign v22f0646 = hmaster2_p & v22eda43 | !hmaster2_p & v84561b;
assign v22efce1 = hmaster1_p & v22fc212 | !hmaster1_p & v230056c;
assign v22fa16d = hbusreq0_p & bd7b37 | !hbusreq0_p & v84561b;
assign v23fba04 = hbusreq4 & v23fb938 | !hbusreq4 & v2310ffa;
assign v23122cd = hmaster2_p & v2304c77 | !hmaster2_p & v22fab30;
assign v22feb98 = hbusreq1 & v22fef02 | !hbusreq1 & v84561b;
assign v2300d67 = hbusreq3 & v22ecca9 | !hbusreq3 & v23f182c;
assign v23fb667 = hbusreq3 & v23fc497 | !hbusreq3 & v84561b;
assign v2305741 = hmaster0_p & v23f6b2f | !hmaster0_p & !v84561b;
assign v23fc1d3 = hbusreq6 & v22ed494 | !hbusreq6 & v23f91bc;
assign v230e882 = hbusreq3_p & v230eeb5 | !hbusreq3_p & v2308c3d;
assign v23f69e4 = hmaster0_p & v23fbcf8 | !hmaster0_p & v23fccb7;
assign v230e539 = hbusreq3_p & v22f7dbc | !hbusreq3_p & !v23f39e6;
assign v2309856 = hmaster0_p & v22f5b58 | !hmaster0_p & v230b38b;
assign v230e821 = hbusreq1_p & v23f616b | !hbusreq1_p & !v2307a62;
assign v1507464 = hbusreq1 & v23930d2 | !hbusreq1 & v150745f;
assign v23f2426 = hmaster2_p & v84561b | !hmaster2_p & !v2303ebe;
assign v230bd77 = hgrant3_p & v230d8af | !hgrant3_p & v23fcbc3;
assign v191ab5f = hbusreq5 & v23fce71 | !hbusreq5 & v84561b;
assign v22f8fe0 = hbusreq0_p & a1fbc2 | !hbusreq0_p & v22eb377;
assign v22f5f7e = hbusreq1 & v23fbdb0 | !hbusreq1 & v84561b;
assign v23fcd3c = stateG10_5_p & v23fcf91 | !stateG10_5_p & v2306d29;
assign v230200a = hmaster2_p & v23126ae | !hmaster2_p & v22f56d2;
assign v23fbd52 = hgrant1_p & a1fba6 | !hgrant1_p & v22f0295;
assign v230b4ad = hmaster2_p & v23fc393 | !hmaster2_p & !v23065ad;
assign v22fa101 = hmaster2_p & v84561b | !hmaster2_p & v23017ee;
assign v230dc17 = hmaster2_p & v23108b7 | !hmaster2_p & !v22f5583;
assign v23018b7 = hbusreq3_p & v191ab12 | !hbusreq3_p & v2392f80;
assign v22fa064 = hgrant1_p & v22f24f8 | !hgrant1_p & v2312351;
assign v23fca52 = hbusreq1_p & v2302225 | !hbusreq1_p & v230a050;
assign v22fd8f6 = hmaster2_p & v2312f7e | !hmaster2_p & v23fc017;
assign b7ab40 = hgrant1_p & v845635 | !hgrant1_p & v230b3a5;
assign v22efadc = hmaster0_p & v9122cc | !hmaster0_p & v22f8cb9;
assign v23fc060 = hbusreq6 & v23022d0 | !hbusreq6 & v84561b;
assign v23120a5 = hbusreq1_p & v22f7aff | !hbusreq1_p & !v230ca0f;
assign v2303ae8 = hmaster2_p & v22fb1bc | !hmaster2_p & v23fcd14;
assign v15075e0 = hbusreq3_p & v22f891a | !hbusreq3_p & v22f859d;
assign v22f8e5d = hbusreq5 & v84561b | !hbusreq5 & !v23fb4bd;
assign v23fd00d = hlock3_p & v231363c | !hlock3_p & !v22f07d3;
assign v23fb4a8 = stateG10_5_p & v23f67bd | !stateG10_5_p & !v23064ae;
assign v22eec8b = hbusreq1_p & v23fd01b | !hbusreq1_p & !v106ae19;
assign v23fc11a = hgrant3_p & v22f6d82 | !hgrant3_p & v89e88b;
assign v23fbca0 = hbusreq3 & v23f1816 | !hbusreq3 & v2311fb5;
assign v23fb61d = hbusreq3_p & v22f07d5 | !hbusreq3_p & v23f7d2e;
assign v22ee50f = hbusreq1 & v22f2718 | !hbusreq1 & v84561b;
assign v22f90a5 = hmaster2_p & v84561b | !hmaster2_p & v22f274e;
assign v23fc318 = hlock3_p & v22f082f | !hlock3_p & v2302b3e;
assign v230da69 = hmaster2_p & v23fc51c | !hmaster2_p & v230e8a6;
assign v22fa20a = hgrant0_p & a1fba6 | !hgrant0_p & v22f1874;
assign v23fc034 = hgrant3_p & v84561b | !hgrant3_p & v23fcedb;
assign v23116cd = hbusreq4_p & v23fc5bf | !hbusreq4_p & f4064b;
assign v23f83f3 = hbusreq1_p & v22f7241 | !hbusreq1_p & v23fba3e;
assign v2302de2 = hmaster1_p & v23f38b1 | !hmaster1_p & v23016dc;
assign v23fa2ec = hbusreq2_p & v15072de | !hbusreq2_p & v84561b;
assign v231057b = hgrant1_p & v23fc3d4 | !hgrant1_p & v22f0d2b;
assign v2305d92 = hmaster2_p & v22f26fc | !hmaster2_p & v23f3b1e;
assign v22fc53d = hbusreq3_p & a8e3ee | !hbusreq3_p & !v84561b;
assign v23fb914 = hbusreq5 & v230913d | !hbusreq5 & !v22f8ac3;
assign v23fb92b = hmaster2_p & v23f5cb3 | !hmaster2_p & !v22fe426;
assign v2310ffa = hgrant3_p & v2301652 | !hgrant3_p & v23015c2;
assign v23f5ce0 = hlock5_p & v84561b | !hlock5_p & v2312d20;
assign v23fcdac = hgrant0_p & v84561b | !hgrant0_p & v191b155;
assign v22fee9e = hgrant3_p & v2306bfb | !hgrant3_p & c0e31a;
assign v230a742 = hbusreq6_p & v23f839a | !hbusreq6_p & v84561b;
assign v23043ec = hbusreq1_p & v23f763f | !hbusreq1_p & v230e23c;
assign v230627c = hbusreq3_p & v22f854f | !hbusreq3_p & v861565;
assign v2393321 = hmaster2_p & v2307a5e | !hmaster2_p & v22ecbbd;
assign v23fba35 = hbusreq2 & v84561b | !hbusreq2 & b5e598;
assign v22f0fd7 = hbusreq0_p & v23fb47c | !hbusreq0_p & v84561b;
assign v22f0e99 = hmaster2_p & v23f646e | !hmaster2_p & v106af73;
assign v23041ed = jx1_p & v2310c61 | !jx1_p & v2309bcf;
assign v2302937 = locked_p & v12cd9cd | !locked_p & v84561b;
assign v23f9c04 = hmaster0_p & v23127b2 | !hmaster0_p & v23fc99c;
assign v230b1ab = hbusreq4_p & v23f673b | !hbusreq4_p & v84561b;
assign v23f18fc = hmaster0_p & v22f5b58 | !hmaster0_p & v22f6ae5;
assign b9d02f = hready & v23fb95d | !hready & !v23f2508;
assign v22fc893 = hbusreq3_p & v23fcc67 | !hbusreq3_p & v845620;
assign v22fdb97 = hmaster1_p & v22f54a0 | !hmaster1_p & v23f8328;
assign v23fca48 = hbusreq0 & v22ee0c4 | !hbusreq0 & !v84561b;
assign v230f403 = hmaster0_p & v23f5af8 | !hmaster0_p & v22f9e08;
assign v22eb8e1 = hbusreq6_p & v23fc53d | !hbusreq6_p & v84561b;
assign v23044d2 = hmaster2_p & v23fc393 | !hmaster2_p & !v23126ae;
assign v23fcf88 = hmaster2_p & v22f65d5 | !hmaster2_p & v84561b;
assign v2311a34 = hmaster2_p & v22fd008 | !hmaster2_p & v23126f2;
assign v23fcd0e = hbusreq1 & v22eb5b3 | !hbusreq1 & !v84561b;
assign v230bd1b = hmaster2_p & v2301511 | !hmaster2_p & v84561b;
assign v23f22a1 = hbusreq5 & v845620 | !hbusreq5 & !v84561b;
assign v22f7929 = hlock0_p & v23fc265 | !hlock0_p & v84561b;
assign v2305338 = hbusreq5 & v23fbfd0 | !hbusreq5 & v84561b;
assign v23f83af = hmaster1_p & v23fc550 | !hmaster1_p & v22ff0ef;
assign v23f5a68 = hlock6_p & v2309e7a | !hlock6_p & v230f5a4;
assign v23f1193 = hbusreq3_p & v23fc23b | !hbusreq3_p & v84561b;
assign v22fb5f1 = hmaster0_p & v23fb923 | !hmaster0_p & v1507557;
assign v22ef116 = hbusreq4_p & v2300b7b | !hbusreq4_p & v22ffcec;
assign v23f3724 = hgrant5_p & v84561b | !hgrant5_p & v23f4ca0;
assign v2310cbb = hbusreq4_p & v23f88d9 | !hbusreq4_p & v22fc3c7;
assign v2393b93 = hbusreq0 & v23fc7b2 | !hbusreq0 & v22ff090;
assign v230b879 = hbusreq3_p & v86c778 | !hbusreq3_p & v23fc6db;
assign v23f8534 = hmaster0_p & v2308dcf | !hmaster0_p & v23f302c;
assign v22ff0ce = hbusreq6 & v22f4d97 | !hbusreq6 & v23fb4cf;
assign v23fc39f = hmaster0_p & v22f97c3 | !hmaster0_p & v22f3b8c;
assign v22fc374 = hmaster2_p & v2308a4b | !hmaster2_p & v23fc06c;
assign v22ff400 = hmaster0_p & v2302f63 | !hmaster0_p & v22f0e4e;
assign v230f47e = hmaster2_p & v84561b | !hmaster2_p & v22ed000;
assign v23f4fa9 = hbusreq6_p & v2312e39 | !hbusreq6_p & v23f9dba;
assign v22f4f06 = hgrant3_p & v22f46ff | !hgrant3_p & v23fc039;
assign v23f6926 = hbusreq0_p & c16191 | !hbusreq0_p & !v2312259;
assign v23000a8 = hgrant4_p & v84561b | !hgrant4_p & v23fc9a4;
assign v23fa94e = hmaster2_p & v2306d29 | !hmaster2_p & v9b93b3;
assign v22fca43 = jx1_p & v2311790 | !jx1_p & v22fbc04;
assign v22ed467 = hlock5_p & v22f1b4e | !hlock5_p & !v23056b1;
assign v23fcc7c = hmaster0_p & v231354e | !hmaster0_p & !v23f7be0;
assign v23f9a46 = hbusreq3 & a8a256 | !hbusreq3 & v84564d;
assign v23fbef6 = hlock3_p & v230cb0f | !hlock3_p & v230ed08;
assign v2309410 = hmaster1_p & v23055c3 | !hmaster1_p & v23103e6;
assign v22f0824 = hbusreq0_p & v23fc681 | !hbusreq0_p & v84561b;
assign v1aae2c1 = hbusreq6_p & v23fb599 | !hbusreq6_p & v22f62a9;
assign v22ede4d = locked_p & v22ef2c3 | !locked_p & v84561b;
assign v23f41af = jx0_p & v23f6aab | !jx0_p & c098a9;
assign v230a193 = hmaster0_p & v239160b | !hmaster0_p & !v230065b;
assign v230f7ff = hmaster2_p & v22fbd02 | !hmaster2_p & v23f445f;
assign v2308b7c = hbusreq5 & v23131e8 | !hbusreq5 & v2306220;
assign v23fbcd4 = hmaster2_p & v22fd0e6 | !hmaster2_p & v230ce60;
assign v230e8ea = hmaster0_p & v23fcb9f | !hmaster0_p & v231256b;
assign v22fa999 = hbusreq1_p & v2309fb1 | !hbusreq1_p & v230e165;
assign v23fcdc9 = hbusreq1_p & v22f343b | !hbusreq1_p & v2302071;
assign v23f33c7 = hmaster0_p & v230eeb6 | !hmaster0_p & v23f96d0;
assign v23f7700 = hbusreq5_p & v231086d | !hbusreq5_p & v84561b;
assign v22f2730 = hbusreq5_p & v106a782 | !hbusreq5_p & v23fba9b;
assign v22f8ee3 = hmaster2_p & v2304074 | !hmaster2_p & v22ee956;
assign v230b9fc = hbusreq6_p & v23fce89 | !hbusreq6_p & v230a87b;
assign v230fdd7 = hlock1_p & v191ac91 | !hlock1_p & v23060b1;
assign v239157f = hmaster0_p & v23fbed7 | !hmaster0_p & v22ef5f1;
assign v23f0872 = hmaster2_p & v23fba9a | !hmaster2_p & v23fb624;
assign v22fb44a = hbusreq4 & v23fcc5f | !hbusreq4 & v84561b;
assign b9d0ca = hbusreq3_p & v2308ecc | !hbusreq3_p & v23fbfb5;
assign v23002bf = hmaster2_p & v22f5583 | !hmaster2_p & v84561b;
assign v230cd34 = hgrant3_p & v230d45f | !hgrant3_p & v22f6529;
assign v2308237 = hbusreq3_p & v22f90d2 | !hbusreq3_p & !v84561b;
assign v23f988f = hbusreq5 & v230bc8b | !hbusreq5 & v23fcb5e;
assign v2301ac0 = hgrant3_p & v23047e5 | !hgrant3_p & v23fce5f;
assign v230e312 = hready_p & v230933a | !hready_p & v23fbf83;
assign v22feff6 = hbusreq4_p & v23f8ba7 | !hbusreq4_p & v22edbd4;
assign v22fe415 = hbusreq3_p & v23051f6 | !hbusreq3_p & v23122cd;
assign v23f4526 = hmaster2_p & v23f9789 | !hmaster2_p & v84561b;
assign v2312925 = hbusreq3_p & v22f0538 | !hbusreq3_p & v2393321;
assign v2300597 = hbusreq0_p & v23fc2fd | !hbusreq0_p & v84561b;
assign v2310319 = hgrant3_p & v230b8fb | !hgrant3_p & v23fb5ec;
assign v230f5e2 = hlock0_p & v2307582 | !hlock0_p & v23fb4b6;
assign v2303220 = jx2_p & v23fc517 | !jx2_p & v22eb993;
assign v2304f4c = hmaster2_p & v23f6411 | !hmaster2_p & v22ffbb3;
assign v23fcf9b = hready & v23fc90f | !hready & !v84561b;
assign f405d5 = hbusreq1_p & v230d109 | !hbusreq1_p & v2310516;
assign v2305a91 = hmaster0_p & v23fccc1 | !hmaster0_p & v23fc521;
assign v2300562 = hgrant3_p & v84561b | !hgrant3_p & !v22fd621;
assign v22ed59e = hbusreq1_p & v12cd54c | !hbusreq1_p & !v84561b;
assign v22f0470 = hbusreq0_p & v23fba79 | !hbusreq0_p & v22ee750;
assign v21b0f6a = hbusreq5 & v2301655 | !hbusreq5 & v84562a;
assign v2312e57 = stateG10_5_p & v23920d8 | !stateG10_5_p & v845620;
assign v22fec81 = hbusreq1_p & v23f16fd | !hbusreq1_p & v23fc30e;
assign v22f6219 = hbusreq3_p & v22fa3df | !hbusreq3_p & v230a226;
assign v2393aca = hgrant5_p & v2304db3 | !hgrant5_p & v22f9248;
assign v22eb8ae = hbusreq3_p & v23f3346 | !hbusreq3_p & v23122cf;
assign v22fb842 = hmaster2_p & v23f0329 | !hmaster2_p & v84561b;
assign v23091ce = hmaster1_p & v22f95ec | !hmaster1_p & v230e97b;
assign v84564d = locked_p & v84561b | !locked_p & !v84561b;
assign v22f161f = jx3_p & v2300687 | !jx3_p & v22fe939;
assign v23fca9d = hbusreq6 & v23fcfbe | !hbusreq6 & v84561b;
assign v23f3a07 = hlock5_p & v1aad4fc | !hlock5_p & !v84561b;
assign v230d379 = hbusreq5 & v23f36a5 | !hbusreq5 & v84561b;
assign v23f3e77 = hmaster0_p & v23fbaed | !hmaster0_p & v23f3de0;
assign c26df3 = hmaster1_p & v22f32df | !hmaster1_p & v231138f;
assign v22f16ad = hgrant3_p & v2393527 | !hgrant3_p & v23faae7;
assign v23fc3af = hbusreq6 & v22f8ebe | !hbusreq6 & v84561b;
assign v1e8408b = stateG2_p & v84561b | !stateG2_p & !v845649;
assign v22f82cd = hmaster2_p & v22f4aa2 | !hmaster2_p & v22efb77;
assign v85c335 = hbusreq3 & v22eb4b3 | !hbusreq3 & v84561b;
assign v23f53bd = hgrant1_p & v845626 | !hgrant1_p & v23fc3f5;
assign v22eb933 = hgrant3_p & v22f1ee0 | !hgrant3_p & v231125d;
assign v23127fb = hbusreq5 & v2302048 | !hbusreq5 & v84561b;
assign v230a58f = hbusreq4_p & v22f14ee | !hbusreq4_p & !v84563a;
assign v23f4b99 = hmaster2_p & v845647 | !hmaster2_p & !v2307758;
assign v22eff51 = hmaster2_p & b9d00f | !hmaster2_p & v22f4f42;
assign v23fc065 = hbusreq6_p & v23fc79a | !hbusreq6_p & v23f4b9c;
assign v22f2b42 = hlock4_p & v2306e3c | !hlock4_p & v23f28ed;
assign v23f8529 = hbusreq3_p & v22f2bab | !hbusreq3_p & v23f7bc9;
assign v22f2ac8 = hlock3_p & v22fb081 | !hlock3_p & v23fb958;
assign v23fb810 = hbusreq6 & v22fea98 | !hbusreq6 & v84561b;
assign v2302e32 = hbusreq2_p & v191a86f | !hbusreq2_p & !v191a876;
assign v22fccd1 = hmaster2_p & v13afc17 | !hmaster2_p & v22fee3b;
assign v22ecff3 = hmaster2_p & v84561b | !hmaster2_p & v230835d;
assign v23f8186 = hmaster1_p & v22fe1c8 | !hmaster1_p & v23f846c;
assign v239228f = hmaster2_p & v22f7466 | !hmaster2_p & e1e250;
assign v22f18b1 = hgrant0_p & v845623 | !hgrant0_p & v23f5ed5;
assign v22ebe7f = hbusreq5 & v106ae21 | !hbusreq5 & v84564d;
assign v22edfb7 = hbusreq5 & v22fc2bd | !hbusreq5 & b16aac;
assign v2313429 = hmaster1_p & v23122bc | !hmaster1_p & v2304c8b;
assign v23fb2f8 = hmaster2_p & v22fa70c | !hmaster2_p & v23f4722;
assign v2300686 = hbusreq4 & v22fb22e | !hbusreq4 & v2310d04;
assign v23fa3e0 = hlock6_p & b355fd | !hlock6_p & !v84561b;
assign v106a7d8 = jx1_p & v23fc720 | !jx1_p & v23f0db6;
assign v22f52a4 = hmaster2_p & v106a782 | !hmaster2_p & !v230fec6;
assign v106af73 = locked_p & v84561b | !locked_p & v191a879;
assign v2301f63 = hgrant3_p & v2393527 | !hgrant3_p & v23fbadb;
assign v2312441 = hgrant0_p & v23f6721 | !hgrant0_p & !v84561b;
assign v23fccca = stateG10_5_p & v23f7094 | !stateG10_5_p & v845636;
assign v23fc942 = hlock4_p & v22fff51 | !hlock4_p & v84561b;
assign v23043b1 = hbusreq4_p & v23f8f18 | !hbusreq4_p & v22f7303;
assign v22f3262 = hbusreq3_p & v230a4f1 | !hbusreq3_p & a136c1;
assign v230c6c7 = hgrant3_p & v84561b | !hgrant3_p & v23fb6bb;
assign v23f5a4e = hlock6_p & v239158e | !hlock6_p & v84561b;
assign v230e869 = hbusreq3_p & v2311cd1 | !hbusreq3_p & v2304bc1;
assign v23fb9e7 = hgrant3_p & v22f988a | !hgrant3_p & v22f679a;
assign v23fc783 = hbusreq3_p & v23f79a7 | !hbusreq3_p & v23fcd49;
assign v23fb975 = hmaster0_p & v23139e3 | !hmaster0_p & !v23fbbf9;
assign v22f3cf2 = hbusreq3_p & v230a573 | !hbusreq3_p & v22fd696;
assign v22ec890 = hgrant3_p & v23035ba | !hgrant3_p & v23fbd70;
assign v23046f7 = locked_p & v23fb136 | !locked_p & v191a879;
assign v23fccd6 = hmaster2_p & v23128a1 | !hmaster2_p & v23fc023;
assign v23f1688 = hmaster0_p & v22fba38 | !hmaster0_p & !v239387a;
assign v22eb9e7 = stateG10_5_p & v23fb98f | !stateG10_5_p & v230a9eb;
assign v22ff8a6 = hbusreq5 & v84561b | !hbusreq5 & !v23068a9;
assign v22ec552 = hbusreq4 & v22f367c | !hbusreq4 & v22f8ba5;
assign v22fe19a = hmaster2_p & v9d8aae | !hmaster2_p & v23fbbd2;
assign v22f95e4 = hbusreq6_p & b61053 | !hbusreq6_p & v22ebc8f;
assign v23fc9db = hbusreq2_p & v22eab01 | !hbusreq2_p & !v84561b;
assign v23f909e = hbusreq1 & v23fc530 | !hbusreq1 & !v84562a;
assign v2312268 = hbusreq6 & v23fb9ad | !hbusreq6 & v84561b;
assign v22fb638 = hready_p & v22ff7ef | !hready_p & v23f8b2b;
assign v23008a6 = hgrant3_p & v23fc1b3 | !hgrant3_p & v23fc03c;
assign v23064bf = hbusreq4_p & v23fc2f6 | !hbusreq4_p & v23fc029;
assign v23060c7 = hbusreq5_p & v23fbd80 | !hbusreq5_p & v84561b;
assign v22ff457 = hbusreq5_p & v106ae19 | !hbusreq5_p & b9d013;
assign v230e851 = hbusreq5_p & v23fbd26 | !hbusreq5_p & !v23fce66;
assign v230e760 = hmaster2_p & v231009b | !hmaster2_p & !v23fb9ad;
assign v230c6c0 = hmaster2_p & v23fcf46 | !hmaster2_p & v2310e40;
assign v22ee657 = hbusreq3 & v845645 | !hbusreq3 & v84561b;
assign v9ed019 = hgrant3_p & v84561b | !hgrant3_p & !v23fc880;
assign e1dd6a = hgrant0_p & v23fbe51 | !hgrant0_p & !v22f753d;
assign v2307788 = hgrant5_p & v22f05f3 | !hgrant5_p & v23fcedd;
assign v2309e7a = hbusreq4_p & v23090a6 | !hbusreq4_p & v23fc826;
assign v23041e2 = hbusreq1_p & v22ecc15 | !hbusreq1_p & v2392d6d;
assign v22f668b = hmaster0_p & v22ef1f3 | !hmaster0_p & bd1c32;
assign v23fbd5b = hmaster0_p & v2303c5a | !hmaster0_p & v2304048;
assign v22f31b2 = hbusreq5_p & v23fb786 | !hbusreq5_p & v84561b;
assign v230e9be = hlock6_p & a1fc9e | !hlock6_p & v22ec77a;
assign v2310a7e = hlock0_p & v23fceb9 | !hlock0_p & v84562b;
assign v23011c7 = hmaster2_p & v23fb4be | !hmaster2_p & !v84561b;
assign v23f5d7f = hbusreq2_p & v230b78b | !hbusreq2_p & v23fbcef;
assign v23101f4 = hbusreq6 & v23fd014 | !hbusreq6 & be7d90;
assign v23105ac = hlock6_p & v22fc2c1 | !hlock6_p & v2309561;
assign v230a942 = hbusreq4 & v23fb862 | !hbusreq4 & v84561b;
assign v22f1ab6 = hgrant3_p & v230b38b | !hgrant3_p & v23106e3;
assign v230f537 = hgrant1_p & v22ecd97 | !hgrant1_p & v23fbe09;
assign v22f3cc0 = hgrant3_p & v230f883 | !hgrant3_p & v23f3ff7;
assign v2305630 = jx3_p & v9b1253 | !jx3_p & v2310d1e;
assign v23f3c20 = hburst0 & v22fdb21 | !hburst0 & !v23fc8d7;
assign v23faaef = hbusreq1 & v1aae29a | !hbusreq1 & v23f8364;
assign v23fcbe1 = hlock0_p & v23fb66a | !hlock0_p & v23fc370;
assign v22f8986 = stateG10_5_p & v22ee195 | !stateG10_5_p & v2304074;
assign v23133bb = hgrant0_p & a1fbc2 | !hgrant0_p & v22f2271;
assign v2304781 = hgrant1_p & v23f908f | !hgrant1_p & v23051fd;
assign v191b1f3 = hgrant0_p & v22efc2a | !hgrant0_p & !v22fdbf7;
assign v2312392 = hbusreq5 & v84561b | !hbusreq5 & !v12cc72f;
assign v23fbe11 = hgrant6_p & v84562d | !hgrant6_p & v23fc59e;
assign v230dce6 = hgrant3_p & v84561b | !hgrant3_p & v99ce01;
assign v22f5611 = hbusreq5 & v1aae56f | !hbusreq5 & v84561b;
assign v23fbfe5 = hbusreq1 & v22f1389 | !hbusreq1 & v84561b;
assign v231262c = hgrant5_p & v84561b | !hgrant5_p & !v23060a6;
assign v23f613e = hbusreq4_p & b0fc7a | !hbusreq4_p & v22eff53;
assign v22fd522 = hbusreq3_p & v22fd6c8 | !hbusreq3_p & v23f692f;
assign v22f349c = hgrant5_p & v22f43cf | !hgrant5_p & v84561b;
assign v22f5afa = hmaster2_p & v23fba25 | !hmaster2_p & v9442ad;
assign v23fc7ff = hbusreq2_p & v23fc7e5 | !hbusreq2_p & !v84561b;
assign v23fc642 = hgrant4_p & v23f1a83 | !hgrant4_p & v23f41af;
assign v2303b17 = hbusreq5 & v23f301a | !hbusreq5 & v22fede1;
assign v22ef648 = hmaster2_p & v23fa0aa | !hmaster2_p & v231057b;
assign v2303fa1 = hbusreq6_p & v22fd0b6 | !hbusreq6_p & v22fc7e5;
assign v23fc890 = hmaster2_p & v23fcfbe | !hmaster2_p & v845620;
assign v23fbfa5 = jx0_p & v2308980 | !jx0_p & v23fc647;
assign v22ff78b = hbusreq4_p & v230f403 | !hbusreq4_p & v84561b;
assign v23fc6f0 = hlock6_p & v2305dde | !hlock6_p & v23fcaec;
assign v23fcfcd = hbusreq2 & v2312f7e | !hbusreq2 & v84561b;
assign v2306441 = hlock0_p & v23fc974 | !hlock0_p & v230fa92;
assign v23fcdcd = hbusreq6_p & v23fc78a | !hbusreq6_p & v23fcf22;
assign v12cd68e = hgrant1_p & v23f78a4 | !hgrant1_p & a1fcc9;
assign v22ec39f = hmaster0_p & v22f6629 | !hmaster0_p & !v23f9fcf;
assign v22f8013 = hbusreq4_p & v230e352 | !hbusreq4_p & v2307b64;
assign v2312397 = jx1_p & v23047dd | !jx1_p & v23031bc;
assign v22ee124 = hbusreq6 & v23049d7 | !hbusreq6 & v22f5fb4;
assign v22ede16 = hgrant5_p & v22f0380 | !hgrant5_p & v22fab80;
assign v22edadc = hmaster2_p & v230f537 | !hmaster2_p & v22f9452;
assign v22faa7a = jx2_p & v23fc642 | !jx2_p & v22fd3c7;
assign v22ec753 = hbusreq1_p & v23fb752 | !hbusreq1_p & !v84561b;
assign v230ada5 = hbusreq6 & v2305a09 | !hbusreq6 & v23fba11;
assign v2309599 = hmaster0_p & v23fccdb | !hmaster0_p & v90c400;
assign v23fb97f = hlock0_p & v23fceb9 | !hlock0_p & v23fbab2;
assign v22fff04 = hbusreq5_p & v17a34ff | !hbusreq5_p & v23fb5fa;
assign baa1eb = hgrant3_p & v84562e | !hgrant3_p & v23f69a3;
assign v23f847c = hbusreq5 & v22f925b | !hbusreq5 & v84564d;
assign v2312b57 = hbusreq6_p & v2310b15 | !hbusreq6_p & v22ff1cb;
assign v23fc949 = hbusreq0_p & v23fbd5f | !hbusreq0_p & v84561b;
assign v22f0ad8 = hmaster0_p & v23127b2 | !hmaster0_p & v23f836b;
assign v23fc52e = hmaster0_p & v230f18c | !hmaster0_p & v22f8cb9;
assign v22edb60 = hmaster2_p & v22ed85a | !hmaster2_p & v23fc48b;
assign v23f8825 = hgrant5_p & v23fbfea | !hgrant5_p & v22f6fb8;
assign v22faa19 = hmaster0_p & v2306593 | !hmaster0_p & v230b38b;
assign v23105b6 = hbusreq5_p & v23f3f46 | !hbusreq5_p & !v23fc706;
assign v23fbe61 = hgrant2_p & v84561b | !hgrant2_p & v23f68d8;
assign v23fb555 = hlock1_p & b0d6e5 | !hlock1_p & !v84561b;
assign v23fc3e7 = hmaster0_p & v1aad69f | !hmaster0_p & v22fad0f;
assign v22f38ab = hgrant3_p & v22eaee1 | !hgrant3_p & v22ecbc1;
assign v23017c7 = hbusreq3 & v22f9ddc | !hbusreq3 & v23f6215;
assign v22fc2ca = hbusreq4_p & v23fc575 | !hbusreq4_p & !v230a0ad;
assign v23fb9f0 = hgrant3_p & v84561b | !hgrant3_p & v22f0b50;
assign v230b930 = hmaster2_p & v2308d79 | !hmaster2_p & v845647;
assign v230a435 = hmaster2_p & v23f6f88 | !hmaster2_p & v23fc7ba;
assign v23fa9b8 = hbusreq3_p & v23efe71 | !hbusreq3_p & e1e70f;
assign v22f5f72 = hgrant4_p & v22fd6ad | !hgrant4_p & v23fc7fe;
assign v23f9a06 = hbusreq5_p & a1fba6 | !hbusreq5_p & v23fbbcf;
assign v22f2903 = locked_p & v22fef4f | !locked_p & v23fc393;
assign v230eaba = hgrant3_p & v845629 | !hgrant3_p & v2302d9a;
assign v23fbcde = hbusreq6 & v23fba78 | !hbusreq6 & v84561b;
assign v230bd96 = hbusreq5_p & v22ef983 | !hbusreq5_p & !v22fa440;
assign v22eccee = hbusreq0 & v8912cf | !hbusreq0 & !v84561b;
assign v2305a37 = hbusreq3_p & v22ed1a8 | !hbusreq3_p & v84561b;
assign v23fc346 = hbusreq2_p & v84561b | !hbusreq2_p & v1aae087;
assign v23101b1 = hgrant1_p & a1fbc2 | !hgrant1_p & v23001a4;
assign v230f073 = hmaster1_p & v23fbbc0 | !hmaster1_p & v22f25fa;
assign v22f346d = hmaster2_p & v191a86f | !hmaster2_p & v22f7d4e;
assign v22f8556 = hmaster0_p & v23f4e63 | !hmaster0_p & v23f6a00;
assign c25c58 = hbusreq5_p & v84564d | !hbusreq5_p & v23fbb3c;
assign bd7497 = hbusreq6 & v23f93e7 | !hbusreq6 & v2310d04;
assign v2300b96 = hlock5_p & v84561b | !hlock5_p & !v22fa4b4;
assign v23fcc64 = hmaster1_p & v1e84b3e | !hmaster1_p & v231251d;
assign v2312187 = hbusreq0_p & v1aae175 | !hbusreq0_p & v23fc2ee;
assign v23fc3f2 = hlock0_p & v23fc265 | !hlock0_p & v845622;
assign v23fd034 = hgrant5_p & v23f1861 | !hgrant5_p & !v230e8d0;
assign b11fc3 = hgrant6_p & v2308be0 | !hgrant6_p & v22f118f;
assign v23fc965 = hbusreq4_p & v23fba28 | !hbusreq4_p & v23fb828;
assign v23fa66e = hmaster0_p & v22f21f6 | !hmaster0_p & v23fc9ee;
assign v22fe0ef = hmaster2_p & v13afe3a | !hmaster2_p & e1e73c;
assign v23070de = hgrant3_p & v84561b | !hgrant3_p & v231256a;
assign v23fc4d1 = hmaster2_p & v84561b | !hmaster2_p & !v2391d17;
assign v22f0132 = hbusreq1_p & v22f5f7e | !hbusreq1_p & v84561b;
assign v23fc437 = hbusreq6 & v23f46b3 | !hbusreq6 & v84561b;
assign v23f91e7 = hmaster2_p & v23fcaf0 | !hmaster2_p & v22f2f44;
assign v22ec6d9 = hgrant2_p & v22ed7d3 | !hgrant2_p & v84561b;
assign v23faaa7 = hlock5_p & v22fb890 | !hlock5_p & !v84561b;
assign v239350a = hbusreq3_p & v22fffe4 | !hbusreq3_p & v23041ee;
assign v22ff745 = hmaster2_p & v230ff7d | !hmaster2_p & v23fc63b;
assign v23fb8da = hgrant5_p & v2308fc5 | !hgrant5_p & !v23041b6;
assign v239299c = hbusreq4_p & v22f8894 | !hbusreq4_p & v2302244;
assign v22f6246 = hgrant5_p & v2309ab5 | !hgrant5_p & v22f299f;
assign v23fbd2f = hbusreq2_p & v84562a | !hbusreq2_p & !v22ee59c;
assign v22f33d3 = hbusreq5_p & v230d16b | !hbusreq5_p & v22f2e64;
assign v22fa48a = hbusreq0 & v23f022d | !hbusreq0 & v22eedf9;
assign v23fc6bd = hmaster2_p & v2306e35 | !hmaster2_p & v2305148;
assign v2303a58 = hmaster0_p & v23f85a9 | !hmaster0_p & v106a888;
assign v22edf31 = hlock3_p & v22fab7c | !hlock3_p & !v84561b;
assign v22f94a7 = hgrant2_p & v22eb377 | !hgrant2_p & a1fba6;
assign v23fc98e = hbusreq1_p & v22f9927 | !hbusreq1_p & v2311374;
assign v23fbc1d = hbusreq1 & v23fcf83 | !hbusreq1 & v84561b;
assign v230c521 = hmaster2_p & v23fbbe7 | !hmaster2_p & !b9d013;
assign v22ed7d1 = hlock0_p & v230a9eb | !hlock0_p & !v12cd3f4;
assign v2308a4b = hgrant1_p & v22f0af2 | !hgrant1_p & !v191aada;
assign v23fc1df = hgrant1_p & v84561b | !hgrant1_p & v22fac26;
assign v23fbf6d = hgrant3_p & v22f8e29 | !hgrant3_p & v22fadf8;
assign a3aa64 = hlock3_p & v2308237 | !hlock3_p & !v84561b;
assign v23fbfb7 = jx0_p & v230e2bd | !jx0_p & v84561b;
assign v2307582 = hgrant2_p & v23fc9c6 | !hgrant2_p & !v22ec29a;
assign v23fb7a3 = hmaster0_p & v22f9cee | !hmaster0_p & v2391a45;
assign v22f2ffc = hmaster2_p & v23fc51c | !hmaster2_p & v23934f0;
assign v22f6403 = hbusreq6_p & v22f5fe4 | !hbusreq6_p & v22f0445;
assign v23f4dc4 = hmaster0_p & v22fc73a | !hmaster0_p & v23019b7;
assign v1aae9b5 = hbusreq5_p & v23f200b | !hbusreq5_p & v22f878c;
assign v22f05b9 = hmaster2_p & v2392f6b | !hmaster2_p & v2393508;
assign v23f4ae1 = hbusreq0 & v23023c9 | !hbusreq0 & v23017f0;
assign v22fb757 = hbusreq6 & v2306944 | !hbusreq6 & v2309726;
assign v23059c5 = jx0_p & v23f2298 | !jx0_p & v23fca45;
assign v22fcd7c = hbusreq1_p & v2303dcb | !hbusreq1_p & v23f89df;
assign v23f88a1 = hbusreq6_p & v22f6e51 | !hbusreq6_p & v23fa599;
assign v23fcd2a = hlock3_p & v23fc152 | !hlock3_p & v23f8d9f;
assign v22ff106 = hlock0_p & v23110b9 | !hlock0_p & !v84561b;
assign v23fc77b = hbusreq3_p & e1e7a3 | !hbusreq3_p & v231106e;
assign v23fb6a4 = hbusreq1_p & v22ed85a | !hbusreq1_p & v84564d;
assign v22fc42e = hbusreq1 & v23113a4 | !hbusreq1 & v84561b;
assign v22f79fd = hready & v23f8134 | !hready & !v84561b;
assign v22fac2f = hbusreq1_p & v23fba24 | !hbusreq1_p & v22ed741;
assign v2302779 = hlock0_p & v23fcd76 | !hlock0_p & v22f3e94;
assign v22f16d5 = hbusreq1 & v23fc26f | !hbusreq1 & v84561b;
assign v22f0eec = stateG2_p & v2302ca3 | !stateG2_p & !v23fcb5d;
assign v2305fe0 = locked_p & v845647 | !locked_p & !v84561b;
assign v150748b = hgrant5_p & da30f9 | !hgrant5_p & v22f90bf;
assign v1507045 = hmaster2_p & v23f2e42 | !hmaster2_p & v22ffe8d;
assign v22f372e = hmaster2_p & v84564d | !hmaster2_p & !v22ebbea;
assign v23fc83e = hmaster0_p & v230e02e | !hmaster0_p & v230c73d;
assign v23fc223 = hgrant3_p & v23fba11 | !hgrant3_p & v22f8f8c;
assign v23fa3c0 = hmaster2_p & v84561b | !hmaster2_p & v22f4998;
assign v230eaa1 = hmaster2_p & v2306220 | !hmaster2_p & !v22fdc17;
assign v23fc90f = hmastlock_p & v2306d5c | !hmastlock_p & v84561b;
assign v23006de = hbusreq1 & v23fbacf | !hbusreq1 & v22ec299;
assign v23f7148 = hbusreq5 & v85d110 | !hbusreq5 & v84561b;
assign v22fdafe = hmaster2_p & a07f9b | !hmaster2_p & a1fbc2;
assign v23f8efa = hmaster2_p & v10dbf64 | !hmaster2_p & v23fbfb9;
assign v22f0f36 = hgrant3_p & v23f2c65 | !hgrant3_p & v23fc02d;
assign v230d3a4 = hbusreq3 & v23fba9a | !hbusreq3 & v22fab50;
assign v22ee93b = hbusreq6_p & v23fc17f | !hbusreq6_p & v22f5c4c;
assign v23f9c7f = hmaster2_p & v84561b | !hmaster2_p & !v23fc93b;
assign v2310e5d = hbusreq3 & v230f863 | !hbusreq3 & !v84561b;
assign a1fde3 = hbusreq0_p & v22ebe16 | !hbusreq0_p & v84561b;
assign v23fc97f = hbusreq6_p & v2310c98 | !hbusreq6_p & v23f3c98;
assign v2305483 = hbusreq4 & v23fbd5d | !hbusreq4 & v2300f25;
assign v1507446 = hgrant3_p & v230d8af | !hgrant3_p & v23fba42;
assign v230b2a4 = hgrant3_p & v230a7a5 | !hgrant3_p & v2303199;
assign v2309df7 = hmaster2_p & v23f87f4 | !hmaster2_p & v22ef403;
assign v23fc550 = hbusreq6_p & v22fb260 | !hbusreq6_p & v230b7c8;
assign v22f91ef = hmaster2_p & v23fbfb9 | !hmaster2_p & v23fcc36;
assign v22f97fe = hmaster2_p & v22fab30 | !hmaster2_p & v230e3a0;
assign v22f9f47 = hbusreq4 & v230f795 | !hbusreq4 & v23f4526;
assign v239253c = hbusreq5_p & v23f646e | !hbusreq5_p & v23fc7a4;
assign v2304ee5 = hgrant5_p & v23f730d | !hgrant5_p & v22edee1;
assign v23fc6a7 = hgrant3_p & v17a34ff | !hgrant3_p & v22f1491;
assign v23fc341 = hgrant5_p & v84561b | !hgrant5_p & v230415a;
assign v2309295 = hmastlock_p & bd757c | !hmastlock_p & v84561b;
assign v2306b1d = jx1_p & v23fc781 | !jx1_p & !v23fbb1b;
assign v23f529c = hgrant0_p & v22f1133 | !hgrant0_p & v22f264f;
assign v23f7372 = hbusreq5_p & e1dcf6 | !hbusreq5_p & v23fafc1;
assign v23fcdb8 = hbusreq4_p & v2309294 | !hbusreq4_p & v230b0f9;
assign v23f480d = hgrant5_p & v22ff9d9 | !hgrant5_p & v23fcccd;
assign v9442ad = hbusreq1_p & a1fbcb | !hbusreq1_p & !v84561b;
assign jx0 = v106a8b9;
assign v23fb848 = hbusreq5_p & v13afa38 | !hbusreq5_p & v23fb1d4;
assign v23f16dc = hlock3_p & v1aad8a8 | !hlock3_p & v22fc37d;
assign v230bc37 = hbusreq6_p & v22fc231 | !hbusreq6_p & v231210f;
assign v2313564 = hgrant1_p & v23093a7 | !hgrant1_p & v2392095;
assign v230a919 = hbusreq3 & v22f881b | !hbusreq3 & v2307632;
assign v2307646 = stateG10_5_p & v2313618 | !stateG10_5_p & !v23fc904;
assign v230efa2 = hmaster1_p & v22f9f01 | !hmaster1_p & v23929fd;
assign v23fc530 = hlock0_p & v230446f | !hlock0_p & v87cfb8;
assign v230bece = hgrant3_p & v2303ae8 | !hgrant3_p & v23005a9;
assign v23fcd16 = hbusreq5 & v23efe0a | !hbusreq5 & v84561b;
assign v22f249f = hgrant1_p & a1fd46 | !hgrant1_p & v230d5be;
assign v23fb7d1 = hlock0_p & v9e3170 | !hlock0_p & v845620;
assign v230a951 = hbusreq1 & v230e8d3 | !hbusreq1 & v23f87f4;
assign v230e857 = hmaster2_p & v9526ac | !hmaster2_p & v22ee956;
assign v22fbe9e = hbusreq4_p & v23f2856 | !hbusreq4_p & v230f857;
assign v230f050 = hgrant0_p & v23fc914 | !hgrant0_p & !v22ee34a;
assign v22f3092 = hbusreq3 & v22fd663 | !hbusreq3 & v84561b;
assign v23f89fc = hbusreq4 & v23fc180 | !hbusreq4 & !v1aad988;
assign v22f8da5 = hgrant5_p & v2303388 | !hgrant5_p & v23fbc07;
assign v23fc6d9 = hbusreq0_p & v106a782 | !hbusreq0_p & v22ed346;
assign v230adfa = jx0_p & v22f7b24 | !jx0_p & v22f5898;
assign v23fc01f = hmaster0_p & v230f133 | !hmaster0_p & v23f5066;
assign v23f133b = hgrant5_p & v22fc3c4 | !hgrant5_p & v230eb8d;
assign v22ebd0b = hbusreq6_p & v1aad9cb | !hbusreq6_p & v23f682c;
assign v960676 = hmaster2_p & v22f0218 | !hmaster2_p & v23fc957;
assign v23fc15f = hbusreq6 & v22f28c4 | !hbusreq6 & v84561b;
assign v23fc1ab = hgrant3_p & v84561b | !hgrant3_p & v22f3b00;
assign v22f94ba = stateG10_5_p & v23f1d8b | !stateG10_5_p & v23fcd29;
assign v230248b = hbusreq2 & v23fc514 | !hbusreq2 & !v23022b1;
assign v23fc5a3 = hbusreq5_p & v23052cc | !hbusreq5_p & v23fc096;
assign v2304cd0 = hbusreq4 & v23fbe1c | !hbusreq4 & v23f87f4;
assign v2309456 = hgrant1_p & v23fccbe | !hgrant1_p & v23fb6a7;
assign v23f9f68 = stateG10_5_p & v230c428 | !stateG10_5_p & v23fb562;
assign v2311826 = hbusreq3_p & v22ffe44 | !hbusreq3_p & v2304b1d;
assign v23f2fd2 = hbusreq3_p & v22f1754 | !hbusreq3_p & v239288d;
assign v22f721f = hbusreq6_p & v23f3e44 | !hbusreq6_p & v2311eaa;
assign v22f8629 = hgrant5_p & v84561b | !hgrant5_p & !v22fb95e;
assign v22f3feb = hbusreq3_p & v22ffea6 | !hbusreq3_p & v22f61b6;
assign v23fc7b9 = hbusreq4 & v2313077 | !hbusreq4 & !v2303db8;
assign v23fc1be = hbusreq6_p & v22fc0a2 | !hbusreq6_p & v2307572;
assign v22eb72a = stateG10_5_p & v23f3adc | !stateG10_5_p & v2300a5a;
assign v23fb1d1 = hgrant0_p & v22ec303 | !hgrant0_p & !v2313a33;
assign v23fb5c0 = jx0_p & v23fd013 | !jx0_p & !v23f623e;
assign v2308f3d = hgrant5_p & v84561b | !hgrant5_p & v23f7499;
assign v22f8ebe = hbusreq4 & v2311743 | !hbusreq4 & v22ec1ef;
assign v23f022a = hbusreq3_p & v230709c | !hbusreq3_p & v84561b;
assign v22f7793 = hmaster2_p & v84561b | !hmaster2_p & v22fef02;
assign b00ac4 = hmaster2_p & a1fba6 | !hmaster2_p & a1fbc2;
assign e1ddd0 = hgrant2_p & v22f8209 | !hgrant2_p & v84564d;
assign v23fb966 = hbusreq2_p & v22f9d85 | !hbusreq2_p & !v84561b;
assign v22f012b = stateG10_5_p & v15071a5 | !stateG10_5_p & !v106ae19;
assign v22f7c05 = hlock3_p & v23f1279 | !hlock3_p & v23fc6b6;
assign v23f6045 = hbusreq1_p & b7427f | !hbusreq1_p & v84561b;
assign v22f2481 = hbusreq0_p & v2304ed3 | !hbusreq0_p & v84561b;
assign v22f4667 = hbusreq3 & v23fc16b | !hbusreq3 & v84561b;
assign v23f0734 = hbusreq1 & v230882d | !hbusreq1 & v23f8364;
assign v23f8e0b = stateA1_p & v84561b | !stateA1_p & v23f2216;
assign v22f1fdb = hgrant3_p & v84561b | !hgrant3_p & v2303f50;
assign v2312ea4 = hbusreq6_p & v230dcd9 | !hbusreq6_p & v2307bcb;
assign v230fcad = hbusreq1 & v23fc3f5 | !hbusreq1 & v22f7241;
assign d79b38 = hmaster2_p & v230f347 | !hmaster2_p & v23fc38f;
assign v22f1dc4 = hmaster2_p & v2306220 | !hmaster2_p & !v2392974;
assign v8a34ca = hmaster2_p & v22ec89f | !hmaster2_p & v84561b;
assign v22fe116 = jx1_p & v2301bda | !jx1_p & v23fc08f;
assign v23faaa0 = hmaster2_p & v230bdd0 | !hmaster2_p & v845627;
assign v2312990 = hbusreq1_p & v22edaa4 | !hbusreq1_p & v84561b;
assign v22f9497 = hbusreq2 & v84561b | !hbusreq2 & !v845620;
assign v23fc0e4 = hbusreq3 & v22ec354 | !hbusreq3 & !v84561b;
assign v230f222 = hgrant0_p & v22f021c | !hgrant0_p & v230f5e2;
assign v23fbe85 = jx3_p & v23080be | !jx3_p & v23fa031;
assign v230d4c3 = hbusreq1_p & v2392fd0 | !hbusreq1_p & v23fcd3a;
assign v22f068b = hgrant1_p & v84561b | !hgrant1_p & v231262c;
assign v23fcfab = hbusreq6 & v84564d | !hbusreq6 & v2302131;
assign v23f8294 = hmaster1_p & v230446b | !hmaster1_p & v23fc7d9;
assign v23f982d = hbusreq6 & v23f68ab | !hbusreq6 & !v230ccff;
assign v22f891a = hmaster2_p & v2312dc1 | !hmaster2_p & v22f62ae;
assign v99d709 = hbusreq1 & v2300de3 | !hbusreq1 & v84561b;
assign v22fe4be = hbusreq1_p & v23f595d | !hbusreq1_p & !b9d013;
assign v23f111b = hmaster2_p & v22fe5b1 | !hmaster2_p & v22f9927;
assign v230e41f = hbusreq3 & v23f6089 | !hbusreq3 & v84561b;
assign v230267d = hbusreq4_p & v22f4089 | !hbusreq4_p & v23040a5;
assign v22fcabc = hbusreq3_p & v230c3f5 | !hbusreq3_p & v231285b;
assign v230f010 = hbusreq5_p & v22faba3 | !hbusreq5_p & v84561b;
assign v22f091e = stateG2_p & v84561b | !stateG2_p & v22f80ca;
assign v2303ebe = hbusreq5_p & v23f384c | !hbusreq5_p & v23fb966;
assign v23fb85c = hbusreq1 & v22f8c70 | !hbusreq1 & v84564d;
assign v2300834 = hmaster0_p & v23fc357 | !hmaster0_p & v86e576;
assign v22fbdda = hmaster2_p & v13afe3a | !hmaster2_p & v1aad847;
assign v22ed400 = hgrant3_p & v2393332 | !hgrant3_p & v23f179d;
assign bad6eb = hbusreq4 & v23fc69b | !hbusreq4 & v23fba11;
assign v22f3673 = hgrant6_p & v22ee274 | !hgrant6_p & bebe64;
assign v22eddd9 = hmaster2_p & v22f23a1 | !hmaster2_p & !v230104a;
assign v23fbe99 = hmaster0_p & v23928ae | !hmaster0_p & !v230a934;
assign v22fd15a = hbusreq4_p & v23fc3ac | !hbusreq4_p & v23f632e;
assign v23f3d38 = hlock3_p & v2312060 | !hlock3_p & baa026;
assign v23f79d2 = hlock1_p & v1aadb8e | !hlock1_p & !v84561b;
assign v230e75b = hmaster2_p & v22fd25c | !hmaster2_p & !v22eb1f5;
assign v23fcfb6 = hbusreq3_p & v23fcb3c | !hbusreq3_p & v22fd196;
assign v2308364 = hbusreq3_p & v23f7024 | !hbusreq3_p & v22fbdda;
assign v23f1cf2 = hbusreq6_p & v23f613e | !hbusreq6_p & v22fdc63;
assign v23fcd4a = hgrant5_p & v23fa155 | !hgrant5_p & v23fc619;
assign v22ec882 = hmaster2_p & v2309c8a | !hmaster2_p & v23056b1;
assign v230d1ff = hgrant4_p & v22eb8fb | !hgrant4_p & v22f85f2;
assign v2392f80 = hmaster2_p & v23f4b28 | !hmaster2_p & !v23fc84b;
assign v230f5a4 = hbusreq4_p & v22fb442 | !hbusreq4_p & v23f34b8;
assign v23f3c12 = hmaster2_p & v22f15fe | !hmaster2_p & !v84561b;
assign v23fb104 = hbusreq2 & v230a2bd | !hbusreq2 & v84561b;
assign v22f4527 = hbusreq2 & v23fca06 | !hbusreq2 & !v84561b;
assign v22f322a = hgrant0_p & v84561b | !hgrant0_p & !v23f316e;
assign v2306b2e = hbusreq0 & v191a86f | !hbusreq0 & v84561b;
assign v22f7022 = hmaster2_p & v191aa68 | !hmaster2_p & v23fb029;
assign v22f7be4 = hbusreq3 & v191aed3 | !hbusreq3 & v84561b;
assign v23fc087 = hbusreq6_p & v230b93b | !hbusreq6_p & !v22fcabb;
assign v22f8824 = hbusreq4_p & v22eebd6 | !hbusreq4_p & v23fc39f;
assign v23f0fd1 = hready & v22f5280 | !hready & v9526ac;
assign v23f95ba = hmaster0_p & v23fcbfb | !hmaster0_p & a1fcb8;
assign v23f40d6 = hgrant1_p & v84561b | !hgrant1_p & v2391728;
assign v230db4d = hbusreq5 & v230b089 | !hbusreq5 & v84561b;
assign v22eb015 = jx1_p & v22f4619 | !jx1_p & v230e896;
assign c16218 = hmaster2_p & f40d66 | !hmaster2_p & v23f717f;
assign v23fb0cd = hbusreq5_p & v84561b | !hbusreq5_p & v23fb80a;
assign v2307852 = hgrant1_p & v23fbf10 | !hgrant1_p & !v2308b4b;
assign v23fbcfb = hgrant1_p & v1e83fd9 | !hgrant1_p & v2391dfa;
assign v2310657 = hbusreq0 & v2391b49 | !hbusreq0 & v84561b;
assign v22f5405 = hmaster2_p & v23fc4f8 | !hmaster2_p & v23fa2ec;
assign v23045ae = hmaster2_p & v23f58e5 | !hmaster2_p & v23fc5ff;
assign v23fcb5e = hgrant0_p & v84564d | !hgrant0_p & v2308848;
assign v22ecb49 = hmaster2_p & v23f0169 | !hmaster2_p & v84561b;
assign v22fa0d4 = hgrant3_p & v22ef31d | !hgrant3_p & v23fc019;
assign v230c404 = hmaster2_p & v22f61b6 | !hmaster2_p & v22f7ab4;
assign v23f5fb9 = hbusreq6_p & v2393031 | !hbusreq6_p & v2311b32;
assign v22f7378 = hgrant5_p & v84561b | !hgrant5_p & v23fb0e3;
assign v22ecdfe = hbusreq1_p & v22feee5 | !hbusreq1_p & v845620;
assign v23f8679 = hgrant1_p & v23fbd0e | !hgrant1_p & v2303707;
assign v9f009f = hgrant2_p & v84561b | !hgrant2_p & v23fa2ec;
assign v23fcfd2 = hgrant3_p & v84561b | !hgrant3_p & v22ee6e8;
assign v2309cfe = hbusreq2 & v23105cd | !hbusreq2 & !v230e6ee;
assign b3865a = hlock1_p & v23f6411 | !hlock1_p & !v106ae19;
assign v22f7195 = hmaster2_p & v22f7da7 | !hmaster2_p & v22f7b47;
assign v23fc746 = hmaster2_p & v22fd696 | !hmaster2_p & v23fbe83;
assign v22f7dd1 = stateG10_5_p & v22f2195 | !stateG10_5_p & v22ff732;
assign v23fc205 = hbusreq5_p & v84561b | !hbusreq5_p & v23fc577;
assign v230db5e = hmaster2_p & v22eec6e | !hmaster2_p & v1e84174;
assign v22f5b75 = hmaster2_p & v22f61b6 | !hmaster2_p & v23fca70;
assign v22fa0ec = hbusreq3_p & c20101 | !hbusreq3_p & v23044d2;
assign v23049cc = hmaster1_p & v9aa6cf | !hmaster1_p & v1aae9e1;
assign v230b6e3 = hmaster2_p & v106a782 | !hmaster2_p & !v2304781;
assign v23f31a9 = hbusreq3 & v23fb2e9 | !hbusreq3 & v84561b;
assign v2306932 = hbusreq0_p & v22f18ad | !hbusreq0_p & v84561b;
assign v22f7c42 = hbusreq6_p & v22eb52b | !hbusreq6_p & v230842d;
assign v23fc1e3 = hlock0_p & v23fc93e | !hlock0_p & v22f06fc;
assign v22f70f4 = hlock2_p & v2304ec7 | !hlock2_p & v84561b;
assign v22eddb2 = hbusreq0 & v23fd021 | !hbusreq0 & v23fb966;
assign v23f280c = hgrant2_p & v22f3396 | !hgrant2_p & !v2301d10;
assign v23f5622 = hgrant5_p & v22ee7e0 | !hgrant5_p & !v23fc133;
assign v22f2b78 = hgrant1_p & v23fc4f8 | !hgrant1_p & v230522c;
assign v23fcb83 = hbusreq1_p & v23001c7 | !hbusreq1_p & v84561b;
assign v23f99a0 = hbusreq6 & v22f0567 | !hbusreq6 & v2310d04;
assign v23fc5b4 = hmaster2_p & v106ae19 | !hmaster2_p & !v979b7c;
assign v2305e51 = hbusreq1_p & v22fed24 | !hbusreq1_p & v23facdf;
assign v22ef867 = stateA1_p & v2302ca3 | !stateA1_p & !v84561b;
assign v23087bc = hbusreq6 & v22ff94b | !hbusreq6 & !v845636;
assign v106a846 = hmaster2_p & v23f4722 | !hmaster2_p & !v23f763f;
assign v2312282 = hmaster1_p & v230b3a5 | !hmaster1_p & v22fb112;
assign v230f75b = hbusreq6 & b00aa6 | !hbusreq6 & v22f1962;
assign v22fdd09 = hlock0_p & v84561b | !hlock0_p & v22efd62;
assign e1df52 = hbusreq6_p & v22fe098 | !hbusreq6_p & v23fb9c7;
assign v22ebb79 = hbusreq1_p & v23f7db8 | !hbusreq1_p & v84561b;
assign be7d90 = hbusreq4 & v23fd014 | !hbusreq4 & v2307d08;
assign a1fbe9 = hgrant3_p & v23fce1e | !hgrant3_p & d79b38;
assign v231160c = hmaster1_p & v22ebb15 | !hmaster1_p & v239268e;
assign v23fc2d2 = busreq_p & v1b87673 | !busreq_p & !v23fcdb9;
assign v22f9d95 = hmaster2_p & v84561b | !hmaster2_p & v22f0870;
assign v22eca5d = hmaster2_p & v230358b | !hmaster2_p & v23003cc;
assign v23f1495 = hbusreq4 & v230420d | !hbusreq4 & v84562f;
assign v22f3196 = hbusreq3 & v2308d79 | !hbusreq3 & !v84561b;
assign v106ae21 = locked_p & v84561b | !locked_p & !v13afe8f;
assign v23f7d51 = hlock2_p & v23f1f6f | !hlock2_p & v23fbb74;
assign v22fe816 = hmaster0_p & v2302f63 | !hmaster0_p & v2392067;
assign v230466c = hmaster0_p & v22f4c34 | !hmaster0_p & v22fb1bc;
assign v231251d = hbusreq4_p & v23fbba5 | !hbusreq4_p & v23f7b0a;
assign v23109c8 = hbusreq4_p & v22ef3aa | !hbusreq4_p & v23015c7;
assign v2308fe5 = hbusreq3_p & v22f03a2 | !hbusreq3_p & !v84561b;
assign v22fcf46 = hbusreq4 & v23f97bb | !hbusreq4 & v84561b;
assign v23f66cf = jx1_p & v22feca2 | !jx1_p & v22f2a85;
assign v23fca2a = hbusreq0_p & v23fcf05 | !hbusreq0_p & v84561b;
assign v230fe65 = hmaster0_p & v23fc1ef | !hmaster0_p & v22ebc57;
assign v23111c2 = hbusreq5_p & v2301e25 | !hbusreq5_p & v22fb88e;
assign v2310116 = hbusreq2_p & v23fc7df | !hbusreq2_p & !v2309c8a;
assign v2311810 = hlock0_p & v84561b | !hlock0_p & a1fba6;
assign v22f6c01 = hlock6_p & v22f0a76 | !hlock6_p & v2391c55;
assign v2312cad = hbusreq3_p & v230d1c3 | !hbusreq3_p & v84561b;
assign v22f11cc = hbusreq4_p & v23fc30a | !hbusreq4_p & v9d7c04;
assign v2304474 = hbusreq6 & v23fbb9b | !hbusreq6 & v84561b;
assign v22ff08f = hbusreq0_p & v22fd30c | !hbusreq0_p & v23056e9;
assign v2313077 = hbusreq3_p & c043dc | !hbusreq3_p & v2310051;
assign v2305cc1 = hgrant3_p & v23fb85a | !hgrant3_p & v1aadf33;
assign v230ace0 = hbusreq2 & v22fafd7 | !hbusreq2 & !v84561b;
assign v23fadf4 = hbusreq1_p & v23f75e9 | !hbusreq1_p & v22f4ef1;
assign v230153d = hbusreq0 & v23fbfd0 | !hbusreq0 & v22f0add;
assign v22f0a22 = hbusreq3_p & v23f3297 | !hbusreq3_p & v23fc016;
assign v23fbeb4 = hburst1 & v23fa931 | !hburst1 & v23f5bdc;
assign v23f384c = hlock5_p & v22ef043 | !hlock5_p & v23fcd1e;
assign v22ef403 = hbusreq5_p & v230b1db | !hbusreq5_p & v84561b;
assign v22feecb = hgrant0_p & v2310a5e | !hgrant0_p & v84561b;
assign v23f5c60 = hmaster2_p & v23f5f5f | !hmaster2_p & !v23f3997;
assign v9b33d9 = hmaster0_p & v2304474 | !hmaster0_p & v230fa04;
assign v23f5d1a = hmaster0_p & v22f2f3e | !hmaster0_p & !v22fdfde;
assign v22f2f87 = hbusreq2_p & v22ec658 | !hbusreq2_p & !v84561b;
assign bd772c = hbusreq4_p & v23fc00a | !hbusreq4_p & v23f5f4d;
assign v2310d04 = hbusreq1_p & v23fa623 | !hbusreq1_p & v84561b;
assign v2313041 = hbusreq3_p & v230426b | !hbusreq3_p & v22ff745;
assign v22f2f19 = hbusreq5_p & v84564d | !hbusreq5_p & v230e9a6;
assign v23fbacf = hgrant5_p & v84561b | !hgrant5_p & v230b611;
assign v2307a49 = hbusreq3_p & v22f2d2a | !hbusreq3_p & v23f149d;
assign v1aae262 = hbusreq1 & v2310a55 | !hbusreq1 & v84561b;
assign v2391f9b = hlock4_p & v23065db | !hlock4_p & !v84561b;
assign v22f0de4 = hmaster0_p & v22fcc78 | !hmaster0_p & v23f99bc;
assign v230886c = hmaster2_p & v22eb599 | !hmaster2_p & v23fa0bf;
assign v23f8d79 = hbusreq3_p & v23fc19b | !hbusreq3_p & v230dc43;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hbusreq2_p = 0;
  hlock2_p = 0;
  hbusreq3_p = 0;
  hlock3_p = 0;
  hbusreq4_p = 0;
  hlock4_p = 0;
  hbusreq5_p = 0;
  hlock5_p = 0;
  hbusreq6_p = 0;
  hlock6_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmaster1_p = 0;
  hmaster2_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  hgrant2_p = 0;
  hgrant3_p = 0;
  hgrant4_p = 0;
  hgrant5_p = 0;
  hgrant6_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  stateG10_2_p = 0;
  stateG10_3_p = 0;
  stateG10_4_p = 0;
  stateG10_5_p = 0;
  stateG10_6_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
  jx3_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hbusreq2_p = hbusreq2;
  hlock2_p = hlock2;
  hbusreq3_p = hbusreq3;
  hlock3_p = hlock3;
  hbusreq4_p = hbusreq4;
  hlock4_p = hlock4;
  hbusreq5_p = hbusreq5;
  hlock5_p = hlock5;
  hbusreq6_p = hbusreq6;
  hlock6_p = hlock6;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmaster1_p = hmaster1;
  hmaster2_p = hmaster2;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  hgrant2_p = hgrant2;
  hgrant3_p = hgrant3;
  hgrant4_p = hgrant4;
  hgrant5_p = hgrant5;
  hgrant6_p = hgrant6;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  stateG10_2_p = stateG10_2;
  stateG10_3_p = stateG10_3;
  stateG10_4_p = stateG10_4;
  stateG10_5_p = stateG10_5;
  stateG10_6_p = stateG10_6;
  jx0_p = jx0;
  jx1_p = jx1;
  jx2_p = jx2;
  jx3_p = jx3;
    end
endmodule

