module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, StoB_REQ4_n, StoB_REQ5_n, StoB_REQ6_n, StoB_REQ7_n, StoB_REQ8_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoS_ACK4_n, BtoS_ACK5_n, BtoS_ACK6_n, BtoS_ACK7_n, BtoS_ACK8_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, SLC2_n, SLC3_n, jx0_n, jx1_n, jx2_n, jx3_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844fbb;
  wire v8e58fd;
  wire v85e3a6;
  wire v844fa1;
  wire v8b555e;
  wire v8991aa;
  wire v8451c3;
  wire v8b5773;
  wire v8e55e7;
  wire v8573c8;
  wire v85d2c4;
  wire v8cce0d;
  wire v8e58ae;
  wire v889f0f;
  wire v8585f1;
  wire v8565ea;
  wire v85667b;
  wire v85dc42;
  wire v85702d;
  wire v86290d;
  wire v8a87cd;
  wire v844f9f;
  wire v8e519b;
  wire v8e19f0;
  wire v8b56ce;
  wire v844f9d;
  wire v8b5875;
  wire v8e3883;
  wire v8e4a1f;
  wire v85aea7;
  wire v889f88;
  wire v8e58d2;
  wire v883cf8;
  wire v85e653;
  wire v8b5768;
  wire v844f9b;
  wire v8e4637;
  wire v8e4831;
  wire v85ffcd;
  wire v885341;
  wire v8e1d42;
  wire v8e570f;
  wire v856765;
  wire v8e17d6;
  wire v85e4bb;
  wire v85da27;
  wire v85b9de;
  wire v8e1933;
  wire v8e2121;
  wire v8e3f65;
  wire v85697c;
  wire v8e3b37;
  wire v85f42f;
  wire v8e4f80;
  wire v85b2a9;
  wire v8e1d5c;
  wire v856656;
  wire v856ce2;
  wire v8e5a35;
  wire v87aaa9;
  wire v844fb7;
  wire v85ea8d;
  wire v8b56bd;
  wire v8e5a72;
  wire v85dffb;
  wire v8e4e35;
  wire v8af0ec;
  wire v8dc5fb;
  wire v8e45f5;
  wire v85e9b9;
  wire v8af41c;
  wire v85dff8;
  wire v8e58cc;
  wire v8e3e4b;
  wire v8e5a59;
  wire v8af160;
  wire v85cd1c;
  wire v856e07;
  wire v8af15c;
  wire v8e4943;
  wire v856eb7;
  wire v8e198d;
  wire v85a4ae;
  wire v8e1ffd;
  wire v8e5896;
  wire v85d69a;
  wire v8564fa;
  wire v8e59c9;
  wire v8e3cda;
  wire v85f343;
  wire v85767f;
  wire v8b582b;
  wire v8af369;
  wire v845037;
  wire v8564f5;
  wire v856b4b;
  wire v85dcb5;
  wire v8e50c2;
  wire v85660f;
  wire v85b898;
  wire v8e5a75;
  wire v8650c5;
  wire v8e4fff;
  wire v85a1ee;
  wire v8451cf;
  wire v8b55c2;
  wire v8e1f2b;
  wire v8af3f2;
  wire v8572c2;
  wire v8b5841;
  wire v85e23a;
  wire v856eba;
  wire v8e59c0;
  wire v8dc552;
  wire v8b5544;
  wire v85e5cf;
  wire v88d6ad;
  wire v8b54e6;
  wire v8e1a9b;
  wire v8e4b9b;
  wire v86695b;
  wire v889f78;
  wire v8e3d4a;
  wire v8e1bda;
  wire v8e4497;
  wire v8565a2;
  wire v8e1852;
  wire v8b5814;
  wire v865770;
  wire v85aa14;
  wire v85ab00;
  wire v8e5000;
  wire v86e8c2;
  wire v8a5c02;
  wire v85b2d3;
  wire v85d8f4;
  wire v84507b;
  wire v85cdc5;
  wire v8b54d3;
  wire v8e4d0b;
  wire v8b54d6;
  wire v8566f3;
  wire v8b565c;
  wire v856919;
  wire v8b5763;
  wire v8b56a4;
  wire v8e4fc9;
  wire v8e5b48;
  wire v8e1755;
  wire v8e482a;
  wire v88e4cb;
  wire v88c352;
  wire v8b5684;
  wire v8e1964;
  wire v85d42c;
  wire v85ca37;
  wire v8e57de;
  wire v856fdd;
  wire v8e198b;
  wire v8e1e8f;
  wire v8b5804;
  wire v867a97;
  wire v8893ab;
  wire v8e58e9;
  wire v845281;
  wire v85dcb6;
  wire v8893b1;
  wire v844fc9;
  wire v844fcb;
  wire v8b57bd;
  wire v89a257;
  wire v8e59f5;
  wire v8b5850;
  wire v85c6d3;
  wire v8967e3;
  wire v85dee1;
  wire v8e4b4d;
  wire v85dbda;
  wire v8e16f6;
  wire v8af325;
  wire v8a5bf8;
  wire v8e3ca1;
  wire v85a6a9;
  wire v86baf9;
  wire v883566;
  wire v85e383;
  wire v85bd67;
  wire v85f5e7;
  wire v856803;
  wire v8dc58d;
  wire v8e3a26;
  wire v8e4764;
  wire v881aaf;
  wire v8e4fad;
  wire v8b584a;
  wire v85dbef;
  wire v85e4ac;
  wire v8e1764;
  wire v8e4cae;
  wire v8e20d0;
  wire v8cc8b1;
  wire v856ff6;
  wire v8e5350;
  wire v856dc8;
  wire v8e508f;
  wire v8b5630;
  wire v89929e;
  wire v856a38;
  wire v856ea9;
  wire v8e4189;
  wire v85fa19;
  wire v8893a8;
  wire v8e4416;
  wire v8e4800;
  wire v85f50b;
  wire v8a5c2b;
  wire v8e3916;
  wire v8e4a14;
  wire v8e599e;
  wire v89928e;
  wire v86513d;
  wire v8e58d4;
  wire v8e5a07;
  wire v8e5372;
  wire v85710e;
  wire v85adf5;
  wire v8e48b6;
  wire v85aeb5;
  wire v865836;
  wire v8b5615;
  wire v8e4e25;
  wire v8e4036;
  wire v8e4432;
  wire v8e4022;
  wire v8b55a7;
  wire v8e3dde;
  wire v8845c4;
  wire v8e52a2;
  wire v8e4ca0;
  wire v8e1106;
  wire v8b3618;
  wire v8e4aa2;
  wire v8e4959;
  wire v865764;
  wire v8e54de;
  wire v8b562d;
  wire v8b5809;
  wire v856725;
  wire v8e21b3;
  wire v860886;
  wire v8e4579;
  wire v8e59e6;
  wire v8e52f2;
  wire v8e4574;
  wire v85acf3;
  wire v844fa0;
  wire v85dbdd;
  wire v85ad39;
  wire v8e4337;
  wire v844f99;
  wire v8dc594;
  wire v844f97;
  wire v8b57d0;
  wire v8e5033;
  wire v8e3911;
  wire v845146;
  wire v8b5577;
  wire v845222;
  wire v8a5c84;
  wire v8b56ee;
  wire v8e4523;
  wire v8cce3b;
  wire v88bcd0;
  wire v86f9a1;
  wire v8a54f3;
  wire v8e3c81;
  wire v8b5757;
  wire v88d5d7;
  wire v88c2b9;
  wire v85ba51;
  wire v8e5298;
  wire v856801;
  wire v8e4191;
  wire v85d3e1;
  wire v8e18e6;
  wire v8e1a97;
  wire v8e594f;
  wire v8573b2;
  wire v85e7be;
  wire v86f856;
  wire v8e1084;
  wire v85df5a;
  wire v8e51d9;
  wire v85f218;
  wire v8b5789;
  wire v8ca6f1;
  wire v8e45a8;
  wire v8e228f;
  wire v8e1090;
  wire v8b55d5;
  wire v8e3a68;
  wire v8cc8cf;
  wire v8e392a;
  wire v8e3e8e;
  wire v8b57ac;
  wire v86f694;
  wire v883d05;
  wire v8e5a3c;
  wire v8af186;
  wire v8e5962;
  wire v8b56eb;
  wire v8e1f02;
  wire v8b5701;
  wire v8e1d78;
  wire v85e858;
  wire v8b5527;
  wire v8af36d;
  wire v8b5565;
  wire v888cd4;
  wire v8e4916;
  wire v8b5699;
  wire v8b42e6;
  wire v8a5c45;
  wire v8e5bd2;
  wire v85f2f8;
  wire v8e5965;
  wire v8e213d;
  wire v8e5a51;
  wire v856b48;
  wire v8e3d7b;
  wire v85ccf0;
  wire v85f59b;
  wire v85e259;
  wire v8e52b0;
  wire v85c971;
  wire v8be123;
  wire v8e42c6;
  wire v8e1be3;
  wire v8b55ff;
  wire v86584f;
  wire v8e1a00;
  wire v8b575f;
  wire v8b5812;
  wire v8dc6a0;
  wire v8e5982;
  wire v8e1d73;
  wire v870e66;
  wire v8e53a5;
  wire v858482;
  wire v85a894;
  wire v8af3c9;
  wire v8b56ae;
  wire v881b59;
  wire v8e1f36;
  wire v8564bf;
  wire v8b5790;
  wire v8e1800;
  wire v8e499d;
  wire v85c9c5;
  wire v8b5517;
  wire v8e464c;
  wire v8e3cf8;
  wire v8e39ff;
  wire v8e3c27;
  wire v8e4662;
  wire v85d7bb;
  wire v867a93;
  wire v85d2e2;
  wire v8a6915;
  wire v8e4e0b;
  wire v8e5426;
  wire v88c32b;
  wire v8b56fa;
  wire v8847b9;
  wire v8b5698;
  wire v8e5952;
  wire v8b579f;
  wire v8b570f;
  wire v85e4fc;
  wire v8b54c7;
  wire v8e157d;
  wire v889270;
  wire v85f3fb;
  wire v85ba2f;
  wire v85dfad;
  wire v856eb5;
  wire v85ea99;
  wire v8e1678;
  wire v8e5611;
  wire v8569a8;
  wire v85d7b1;
  wire v8e3c39;
  wire v8cc8e8;
  wire v8860f1;
  wire v84514a;
  wire v8b56e5;
  wire v8b5799;
  wire v8e1de6;
  wire v85cda6;
  wire v85672e;
  wire v8e23b9;
  wire v8dc607;
  wire v8b54c0;
  wire v856763;
  wire v8564e9;
  wire v8e1fe7;
  wire v8e4fa6;
  wire v8b55ca;
  wire v8e3ee9;
  wire v85f3dd;
  wire v8e4e9e;
  wire v8e5a2b;
  wire v8b573a;
  wire v8b582a;
  wire v88c2c4;
  wire v8e58ac;
  wire v870b4c;
  wire v8e3f8b;
  wire v8b55e6;
  wire v865810;
  wire v89924f;
  wire v8e2395;
  wire v85dee3;
  wire v8e5b68;
  wire v85d3c7;
  wire v866552;
  wire v8e5aa4;
  wire v85c771;
  wire v86e720;
  wire v8af0f7;
  wire v8b5784;
  wire v8566db;
  wire v8565bb;
  wire v8e3b88;
  wire v8e238b;
  wire v8af1a0;
  wire v862911;
  wire v8b54ec;
  wire v85f194;
  wire v8e165a;
  wire v8af389;
  wire v85e93d;
  wire v8e4b64;
  wire v8e38b0;
  wire v8b5771;
  wire v85d7a7;
  wire v880b7a;
  wire v8e45a4;
  wire v85eb04;
  wire v8e59c6;
  wire v8e46e5;
  wire v8b5817;
  wire v8e4dcf;
  wire v8e51cd;
  wire v8e4261;
  wire v8e4f28;
  wire v8575ef;
  wire v8b564d;
  wire v8be114;
  wire v85ae38;
  wire v8572f8;
  wire v8984b0;
  wire v845249;
  wire v85b5fb;
  wire v8b5693;
  wire v8e19a8;
  wire v8e559d;
  wire v8cce31;
  wire v8451d7;
  wire v85ceaf;
  wire v8e5171;
  wire v863e80;
  wire v8451d8;
  wire v8587ce;
  wire v8af292;
  wire v856bd5;
  wire v8e44d0;
  wire v8e438d;
  wire v8b5506;
  wire v88934b;
  wire v8b5530;
  wire v8e3d91;
  wire v85cb8e;
  wire v85b60a;
  wire v85e905;
  wire v8b584f;
  wire v8b559d;
  wire v8b5662;
  wire v8e53e7;
  wire v8e41d9;
  wire v856264;
  wire v8e59d1;
  wire v89921c;
  wire v85dee5;
  wire v85d3cb;
  wire v8e2355;
  wire v8e4c11;
  wire v8626fe;
  wire v8b5651;
  wire v8e589d;
  wire v8af37f;
  wire v8e1982;
  wire v85a07c;
  wire v85d6a8;
  wire v88c339;
  wire v8dc5be;
  wire v85f49e;
  wire v8b5668;
  wire v8cce41;
  wire v85e355;
  wire v8e3ed3;
  wire v84520f;
  wire v8600af;
  wire v85c593;
  wire v8be143;
  wire v8cce46;
  wire v85a277;
  wire v8b54f0;
  wire v8b5563;
  wire v85e281;
  wire v8565b3;
  wire v8e438a;
  wire v85bd37;
  wire v85f2f0;
  wire v8b5667;
  wire v8e5a98;
  wire v85d35a;
  wire v8892d3;
  wire v8e4187;
  wire v8b57b7;
  wire v8e4096;
  wire v865261;
  wire v844fb1;
  wire v85b642;
  wire v8e4086;
  wire v8e2158;
  wire v8af46c;
  wire v85daf5;
  wire v856f73;
  wire v8e4988;
  wire v85d3e9;
  wire v8e585b;
  wire v8b5526;
  wire v8e1c26;
  wire v86cb45;
  wire v866ae1;
  wire v8e20a6;
  wire v8b55d8;
  wire v85d701;
  wire v8e1d85;
  wire v8e15cb;
  wire v8b57a9;
  wire v85740b;
  wire v85ca46;
  wire v8b571f;
  wire v88934d;
  wire v8e4cf4;
  wire v860053;
  wire v8e572f;
  wire v8e19fe;
  wire v8be0ec;
  wire v8e5aa3;
  wire v8b588b;
  wire v8e2136;
  wire v8a5b4f;
  wire v8dc580;
  wire v8e5a1c;
  wire v8e1b44;
  wire v8e2267;
  wire v8af47a;
  wire v8e4f71;
  wire v8dc58b;
  wire v865820;
  wire v8e46de;
  wire v8e1c52;
  wire v8b54f4;
  wire v85f334;
  wire v85653c;
  wire v85a008;
  wire v899197;
  wire v856878;
  wire v884771;
  wire v8a5cca;
  wire v88c371;
  wire v8e594d;
  wire v85699e;
  wire v8b5525;
  wire v8af243;
  wire v8e5754;
  wire v8e54a9;
  wire v85eac4;
  wire v85da38;
  wire v8af402;
  wire v856a03;
  wire v856452;
  wire v8b5543;
  wire v8e1ead;
  wire v85ca40;
  wire v8e4212;
  wire v85ddb7;
  wire v8e5708;
  wire v8bf293;
  wire v8e44eb;
  wire v8e4059;
  wire v8a5bd1;
  wire v8e5486;
  wire v85d757;
  wire v8e58f8;
  wire v8e5b65;
  wire v85d794;
  wire v85d433;
  wire v8e5a33;
  wire v87c63a;
  wire v856575;
  wire v8b55c1;
  wire v85b739;
  wire v85b3c3;
  wire v8af176;
  wire v85e103;
  wire v8e3d1a;
  wire v8e472c;
  wire v8a554f;
  wire v8e162b;
  wire v8e3ea1;
  wire v8b57d9;
  wire v8e5ba4;
  wire v8e4b2a;
  wire v88c355;
  wire v86d6bd;
  wire v85b66d;
  wire v8e1857;
  wire v88bbf7;
  wire v8e1cfb;
  wire v8e4db6;
  wire v889f0e;
  wire v880b8e;
  wire v873e9c;
  wire v8b583b;
  wire v8e4b5f;
  wire v8b54da;
  wire v85eb45;
  wire v8e570a;
  wire v85b5db;
  wire v8b3615;
  wire v8e5914;
  wire v85658e;
  wire v85abee;
  wire v8e1542;
  wire v85fa6e;
  wire v85df70;
  wire v8b585d;
  wire v85b4ff;
  wire v85d52e;
  wire v856799;
  wire v8b56cf;
  wire v8e19b0;
  wire v8b55a3;
  wire v85e4d3;
  wire v8e4b2c;
  wire v8e41fc;
  wire v856f27;
  wire v881b42;
  wire v856b71;
  wire v8cc95b;
  wire v8e5a08;
  wire v85f12d;
  wire v8e589c;
  wire v85aeed;
  wire v856354;
  wire v8e21c5;
  wire v8e4918;
  wire v8e2288;
  wire v8e569c;
  wire v856f79;
  wire v8e4345;
  wire v8b55ef;
  wire v85ba36;
  wire v8b5500;
  wire v8e243e;
  wire v899219;
  wire v8e44b5;
  wire v8e595c;
  wire v8e58d9;
  wire v865f86;
  wire v85f133;
  wire v885f57;
  wire v85cb89;
  wire v8e17c4;
  wire v8e474f;
  wire v8b56a9;
  wire v85f7ea;
  wire v85eaf9;
  wire v85df5b;
  wire v85c7da;
  wire v8e56ca;
  wire v85dd8c;
  wire v8b54d5;
  wire v8e58b1;
  wire v8e4f0c;
  wire v8e3db6;
  wire v856353;
  wire v845027;
  wire v8b564c;
  wire v88e277;
  wire v8e3ff5;
  wire v8563f1;
  wire v85df15;
  wire v8e5a2f;
  wire v8e45e3;
  wire v856406;
  wire v86bc13;
  wire v8a8822;
  wire v85da8e;
  wire v85d886;
  wire v8618f2;
  wire v8e5be4;
  wire v8b5601;
  wire v85cc2a;
  wire v85e619;
  wire v8e4cb9;
  wire v85e9c5;
  wire v8e599d;
  wire v85dce5;
  wire v856c55;
  wire v8565cc;
  wire v8cce04;
  wire v85ba35;
  wire v85cc48;
  wire v8892a6;
  wire v8e4ad3;
  wire v85aaed;
  wire v85f59c;
  wire v8b56ca;
  wire v866529;
  wire v8e5833;
  wire v8e40ce;
  wire v85a25b;
  wire v8e4021;
  wire v8b55cf;
  wire v85643a;
  wire v8af0dd;
  wire v85654c;
  wire v8e59fd;
  wire v8e522a;
  wire v8e44a2;
  wire v8e5194;
  wire v8af3db;
  wire v8b55f0;
  wire v8b54f9;
  wire v881ad8;
  wire v8845b3;
  wire v8b5736;
  wire v85da9f;
  wire v85dfb4;
  wire v8e4668;
  wire v8b56ab;
  wire v8e59cc;
  wire v85ff96;
  wire v8b5691;
  wire v8e58c1;
  wire v8a555c;
  wire v8e1f0e;
  wire v8563cb;
  wire v8cc9b5;
  wire v844fbf;
  wire v844fa5;
  wire v8b55a4;
  wire v8b5732;
  wire v8e5a21;
  wire v8601d6;
  wire v8e19ae;
  wire v8e3a67;
  wire v8e1c59;
  wire v8a552d;
  wire v8b5848;
  wire v8e455f;
  wire v857107;
  wire v8e3af2;
  wire v8b589f;
  wire v8e3a16;
  wire v8e5208;
  wire v8b5579;
  wire v8585db;
  wire v8e1695;
  wire v8b585b;
  wire v856913;
  wire v8e598b;
  wire v85cc2b;
  wire v88bc2b;
  wire v85b670;
  wire v864a5d;
  wire v8e17e8;
  wire v8e1841;
  wire v8a54eb;
  wire v8e5917;
  wire v8e589b;
  wire v8b57c1;
  wire v8e3a36;
  wire v8b58a7;
  wire v8e4131;
  wire v8af277;
  wire v8e5920;
  wire v8e5c6a;
  wire v8b571d;
  wire v8b5551;
  wire v857271;
  wire v857943;
  wire v8992a4;
  wire v8e409a;
  wire v8563df;
  wire v8af190;
  wire v8b56e1;
  wire v8e5949;
  wire v8e3b2b;
  wire v8e59d8;
  wire v8e5a60;
  wire v8e5413;
  wire v8e4153;
  wire v85d73d;
  wire v8b5887;
  wire v860551;
  wire v8b553b;
  wire v889f6d;
  wire v85cb94;
  wire v8e43f1;
  wire v845379;
  wire v8b5837;
  wire v8e4411;
  wire v8b550b;
  wire v8e10b7;
  wire v8e1aee;
  wire v8e118d;
  wire v8e1bf6;
  wire v8e1acc;
  wire v8569c7;
  wire v85659e;
  wire v8e55a6;
  wire v8e425a;
  wire v8566be;
  wire v85f3b1;
  wire v85af2b;
  wire v8e5900;
  wire v856960;
  wire v8e1c5f;
  wire v8b54d8;
  wire v8b57bb;
  wire v8e46a3;
  wire v85b5c5;
  wire v86c57a;
  wire v8450c0;
  wire v85c3e3;
  wire v8b5808;
  wire v8e3c23;
  wire v8e1fa5;
  wire v8e4996;
  wire v85f79e;
  wire v8e4394;
  wire v8e3d36;
  wire v8b5760;
  wire v8e59af;
  wire v8450b6;
  wire v8e1730;
  wire v8b587a;
  wire v8b57f3;
  wire v8cc8fa;
  wire v8e4f0b;
  wire v8e4236;
  wire v85b9a7;
  wire v856902;
  wire v8e4472;
  wire v8e3dd3;
  wire v85ce79;
  wire v8b5884;
  wire v8e4f2e;
  wire v8e588f;
  wire v8dc6bf;
  wire v8e5b16;
  wire v8e1862;
  wire v86006a;
  wire v8e5a54;
  wire v845235;
  wire v85ca8a;
  wire v8bf910;
  wire v85c632;
  wire v856594;
  wire v8e5989;
  wire v8e4636;
  wire v8e4602;
  wire v864f49;
  wire v889f82;
  wire v845074;
  wire v85cdc8;
  wire v8af44d;
  wire v8e47dd;
  wire v8e4b24;
  wire v8e5924;
  wire v8e1a90;
  wire v8e44a1;
  wire v8af34f;
  wire v8e1b23;
  wire v856ec1;
  wire v8e3c8e;
  wire v8af3c1;
  wire v8e5510;
  wire v8e5c10;
  wire v85c6f5;
  wire v8e3a2f;
  wire v8e40a9;
  wire v84507a;
  wire v8e58d6;
  wire v8b5687;
  wire v85c6ec;
  wire v8e5a7f;
  wire v85a8af;
  wire v8e400a;
  wire v899202;
  wire v85e000;
  wire v8e4c04;
  wire v86e4e7;
  wire v8e16ea;
  wire v85f287;
  wire v8e52f8;
  wire v8e466e;
  wire v8e5a10;
  wire v8e1701;
  wire v8e56eb;
  wire v8dc5ec;
  wire v8af327;
  wire v85f53b;
  wire v88c36f;
  wire v856b75;
  wire v8e5891;
  wire v883ca3;
  wire v8b556f;
  wire v8e3d0c;
  wire v8567bb;
  wire v8e1e6a;
  wire v88475f;
  wire v8568a1;
  wire v8e3dc6;
  wire v8e1eb9;
  wire v8e5996;
  wire v8e49ee;
  wire v8b5663;
  wire v8b577d;
  wire v8e45c6;
  wire v8e422f;
  wire v8e1d94;
  wire v8e3af1;
  wire v8e3bf3;
  wire v85ea86;
  wire v845189;
  wire v8e4397;
  wire v8af2e0;
  wire v8e5bb2;
  wire v85f6bc;
  wire v8e5bed;
  wire v85641f;
  wire v8b54db;
  wire v85df78;
  wire v8e4d75;
  wire v8e42fd;
  wire v8e5908;
  wire v86653e;
  wire v85e7d3;
  wire v8e4caf;
  wire v8e49c8;
  wire v85df40;
  wire v85aab4;
  wire v8967e2;
  wire v8b565d;
  wire v845150;
  wire v88c39f;
  wire v8e56dc;
  wire v8572f7;
  wire v8a747c;
  wire v8e54e0;
  wire v8a5bca;
  wire v8e3972;
  wire v8e42df;
  wire v8b5895;
  wire v8a5cb5;
  wire v8562ad;
  wire v84530d;
  wire v8a87ae;
  wire v8be15d;
  wire v8b5750;
  wire v85dda8;
  wire v8e588e;
  wire v8e1a1d;
  wire v8e4185;
  wire v8e1ea1;
  wire v8e1598;
  wire v8e1969;
  wire v870cce;
  wire v8b57d1;
  wire v8e2248;
  wire v8e58c2;
  wire v8e5a66;
  wire v86582c;
  wire v8e4d5c;
  wire v85ad92;
  wire v8e5155;
  wire v857553;
  wire v85d2bd;
  wire v85df2b;
  wire v8b56b7;
  wire v8e1975;
  wire v858462;
  wire v85b29f;
  wire v8e59d0;
  wire v8b5641;
  wire v8dc67d;
  wire v89925a;
  wire v8e4003;
  wire v8e3de2;
  wire v8b558d;
  wire v867a58;
  wire v880dfd;
  wire v85e1b8;
  wire v85adaf;
  wire v8e5c47;
  wire v8e1bc6;
  wire v8e408d;
  wire v867b8d;
  wire v857615;
  wire v8451c4;
  wire v8e1d33;
  wire v8e5bd5;
  wire v863b40;
  wire v889f58;
  wire v85d917;
  wire v889f6b;
  wire v85705c;
  wire v85f62f;
  wire v85dac7;
  wire v8dc68b;
  wire v8e4786;
  wire v8e1add;
  wire v85c416;
  wire v85fb40;
  wire v8e3c73;
  wire v8e587f;
  wire v8b57ff;
  wire v856b08;
  wire v8a87d6;
  wire v85ad35;
  wire v8e1e8c;
  wire v8e3a0e;
  wire v8e5a80;
  wire v8e4cb1;
  wire v8caede;
  wire v85e340;
  wire v8e20ff;
  wire v85f689;
  wire v867a75;
  wire v85fc5a;
  wire v8571d0;
  wire v8af3cb;
  wire v8e18bd;
  wire v8e58c9;
  wire v89b438;
  wire v8e2035;
  wire v8e4254;
  wire v85ccc3;
  wire v856edd;
  wire v85714b;
  wire v85d5a0;
  wire v8e466b;
  wire v8e3e3a;
  wire v885fa8;
  wire v885455;
  wire v8e5428;
  wire v8af0d0;
  wire v8cc8c9;
  wire v8a5bb4;
  wire v8e5344;
  wire v8e199b;
  wire v8e4603;
  wire v8e14dc;
  wire v8e5959;
  wire v8e503a;
  wire v87f6a7;
  wire v885d2d;
  wire v85680b;
  wire v8e59b1;
  wire v8e4ca6;
  wire v8b55cb;
  wire v8e49b1;
  wire v8567fa;
  wire v8cc8fb;
  wire v8be11a;
  wire v8b585f;
  wire v8e59be;
  wire v868a25;
  wire v865862;
  wire v8b5840;
  wire v8574d0;
  wire v8e592f;
  wire v88173a;
  wire v85f2cd;
  wire v86f85b;
  wire v85c6e4;
  wire v8e45fa;
  wire v85a863;
  wire v8e57b4;
  wire v85ea88;
  wire v85cb96;
  wire v8b55a2;
  wire v8e1fdc;
  wire v8e5a64;
  wire v85e994;
  wire v8e38a9;
  wire v8a5b8c;
  wire v8b5826;
  wire v8e5810;
  wire v8e54fe;
  wire v856fa4;
  wire v8e58ad;
  wire v88c2da;
  wire v864623;
  wire v8852fd;
  wire v857374;
  wire v8e416f;
  wire v8db8b5;
  wire v8b576f;
  wire v8b5516;
  wire v8b56fd;
  wire v8e1f00;
  wire v85c986;
  wire v866812;
  wire v8e576d;
  wire v85e111;
  wire v8b577b;
  wire v8e22de;
  wire v85d441;
  wire v8b553e;
  wire v8b55ab;
  wire v8a5b53;
  wire v856959;
  wire v85bdb6;
  wire v876a22;
  wire v856f22;
  wire v8ccdf7;
  wire v8e451f;
  wire v8b572b;
  wire v8e1b43;
  wire v8e5a27;
  wire v8b572d;
  wire v8e59f7;
  wire v88924e;
  wire v8e3b31;
  wire v8e4e75;
  wire v8e179a;
  wire v85f646;
  wire v85dd9f;
  wire v8e4b93;
  wire v8e17b2;
  wire v8e111b;
  wire v85e566;
  wire v85fc19;
  wire v85dbbe;
  wire v8e570e;
  wire v85f223;
  wire v8e45d6;
  wire v86066c;
  wire v8e3c11;
  wire v8e1f7b;
  wire v85dd22;
  wire v8b54f5;
  wire v856c71;
  wire v8e2451;
  wire v85e7ea;
  wire v8e1902;
  wire v8e209c;
  wire v8e1f7f;
  wire v899283;
  wire v85ab77;
  wire v8e520c;
  wire v8b56af;
  wire v8e2303;
  wire v85d43b;
  wire v86e0c8;
  wire v8e44d3;
  wire v85b99e;
  wire v8af107;
  wire v8e4a48;
  wire v85bbcc;
  wire v8e438f;
  wire v8b554e;
  wire v8e2222;
  wire v85d9cc;
  wire v85f386;
  wire v8e5a3f;
  wire v856bb4;
  wire v8e3b5f;
  wire v8e593d;
  wire v88460a;
  wire v8e39cc;
  wire v85b9a9;
  wire v85ada7;
  wire v85e282;
  wire v85b238;
  wire v8e58e0;
  wire v8b5720;
  wire v899fb0;
  wire v85736b;
  wire v845373;
  wire v8e4224;
  wire v8e4294;
  wire v8e55c9;
  wire v8564b7;
  wire v8e38f1;
  wire v867a71;
  wire v85dd8e;
  wire v85bbb6;
  wire v8e407e;
  wire v85dbb6;
  wire v85d475;
  wire v86ae81;
  wire v8e4885;
  wire v86d1ff;
  wire v8984a8;
  wire v85dbe7;
  wire v8cf114;
  wire v8e592e;
  wire v8b573f;
  wire v8b580b;
  wire v85c4c3;
  wire v8e1f2f;
  wire v8e3d40;
  wire v8b5707;
  wire v8e5a4b;
  wire v8b57c9;
  wire v8e55a8;
  wire v8e59bd;
  wire v8e4d0c;
  wire v8b54ea;
  wire v8e190d;
  wire v8e2181;
  wire v8e3c9e;
  wire v8b56ef;
  wire v85c433;
  wire v8e4bdc;
  wire v856895;
  wire v8af2e6;
  wire v8e56d9;
  wire v8e1bc1;
  wire v85fedf;
  wire v8a5561;
  wire v8e5a09;
  wire v8e5c0a;
  wire v85e946;
  wire v8e59e5;
  wire v8e4a96;
  wire v8e58ce;
  wire v85aa21;
  wire v8b588c;
  wire v86e347;
  wire v8e4d7d;
  wire v8e5c1b;
  wire v8e530b;
  wire v8b55f4;
  wire v8e5723;
  wire v8e4670;
  wire v8e46fa;
  wire v85f401;
  wire v8e22b0;
  wire v8567f9;
  wire v85f411;
  wire v8cc8e9;
  wire v85db32;
  wire v85bd7c;
  wire v8e1ebe;
  wire v8b573e;
  wire v8e46da;
  wire v8568f6;
  wire v87ee2b;
  wire v856813;
  wire v8e516c;
  wire v8b5669;
  wire v856951;
  wire v86c2ed;
  wire v85da55;
  wire v8e5ace;
  wire v8672b3;
  wire v845187;
  wire v8e5778;
  wire v8e59f0;
  wire v8e5a73;
  wire v8e5906;
  wire v86582f;
  wire v8e3a6a;
  wire v8e1d76;
  wire v85cdaa;
  wire v8b56b2;
  wire v8e5a2d;
  wire v8e473e;
  wire v8e5646;
  wire v8b5820;
  wire v8e42a4;
  wire v85da20;
  wire v856867;
  wire v8b5505;
  wire v8563e3;
  wire v880b9c;
  wire v8b57a8;
  wire v8e148a;
  wire v8563a2;
  wire v8e10aa;
  wire v8e4c73;
  wire v85b380;
  wire v8b55cc;
  wire v85fabb;
  wire v8e45b5;
  wire v85aba0;
  wire v845160;
  wire v85a600;
  wire v899fe9;
  wire v85c6f0;
  wire v856b36;
  wire v8e56a0;
  wire v8e58f5;
  wire v85665c;
  wire v8e57c2;
  wire v8db551;
  wire v85ae84;
  wire v8e40eb;
  wire v85b5f3;
  wire v8af209;
  wire v856819;
  wire v8a5c04;
  wire v8a5564;
  wire v844fb3;
  wire v8573cd;
  wire v8984a5;
  wire v8e23b1;
  wire v8e5998;
  wire v8a3c77;
  wire v86dabf;
  wire v866544;
  wire v8b5844;
  wire v8af14f;
  wire v85dddb;
  wire v85e8a6;
  wire v8b57fc;
  wire v8e59d4;
  wire v8b54d7;
  wire v8e599c;
  wire v8452da;
  wire v8e572e;
  wire v8e42f6;
  wire v8e2429;
  wire v85f2b2;
  wire v859ffa;
  wire v85fc37;
  wire v85ae77;
  wire v8e18ff;
  wire v8dc668;
  wire v8e1f59;
  wire v8e56e1;
  wire v882912;
  wire v84530b;
  wire v8451a1;
  wire v8e59ee;
  wire v8e4d7b;
  wire v8dc599;
  wire v8e59df;
  wire v8e10a4;
  wire v8e388e;
  wire v8b57df;
  wire v8e41ec;
  wire v865856;
  wire v8cce1f;
  wire v86c65e;
  wire v8b55b0;
  wire v85a51c;
  wire v8b565b;
  wire v8e597a;
  wire v856809;
  wire v8e4c7f;
  wire v8b5794;
  wire v85f35f;
  wire v8e2040;
  wire v8a5b25;
  wire v8b56f5;
  wire v8af40e;
  wire v8af18f;
  wire v8b56b6;
  wire v8b5685;
  wire v86a790;
  wire v8574d6;
  wire v8571db;
  wire v8e2025;
  wire v89920d;
  wire v8e5b0f;
  wire v85b09e;
  wire v85c435;
  wire v8984d7;
  wire v8b566c;
  wire v8e14bc;
  wire v881baf;
  wire v8e5b58;
  wire v8af11e;
  wire v8e5a7e;
  wire v8b56de;
  wire v8e58cb;
  wire v85e006;
  wire v85c120;
  wire v8e4a6c;
  wire v8e212d;
  wire v856b41;
  wire v8e23df;
  wire v8e592b;
  wire v86cbc7;
  wire v8b5682;
  wire v8cce2b;
  wire v8e5223;
  wire v8991c0;
  wire v8a5c49;
  wire v8e5a02;
  wire v8e4e2c;
  wire v8e59a9;
  wire v85727c;
  wire v8b568e;
  wire v8e47f2;
  wire v8e5816;
  wire v85ccfd;
  wire v85e1a0;
  wire v856fe8;
  wire v856a2e;
  wire v8e5707;
  wire v8e1d1f;
  wire v85b724;
  wire v8803e2;
  wire v856ad9;
  wire v8984af;
  wire v8892a1;
  wire v85cde3;
  wire v8563a9;
  wire v85ad8b;
  wire v85e664;
  wire v85e1a3;
  wire v8e5a94;
  wire v85f81e;
  wire v8e591a;
  wire v85e947;
  wire v8574ed;
  wire v8562b6;
  wire v8e5942;
  wire v8b588a;
  wire v85e0ba;
  wire v8b565e;
  wire v8b553d;
  wire v8e4c64;
  wire v856901;
  wire v8b56ad;
  wire v8e55ec;
  wire v8e5a8f;
  wire v8e5032;
  wire v8dc5ad;
  wire v8e1b02;
  wire v8b577f;
  wire v8b5899;
  wire v85d792;
  wire v8dc5d5;
  wire v8e58f9;
  wire v8e57d3;
  wire v8b5518;
  wire v856395;
  wire v8b582f;
  wire v8e15ab;
  wire v8e5a1f;
  wire v8e3f7f;
  wire v8451f9;
  wire v85dc95;
  wire v85768f;
  wire v8e453e;
  wire v8e4f3b;
  wire v85af76;
  wire v8e1650;
  wire v8b5724;
  wire v8cce49;
  wire v8e4d72;
  wire v8e3bdc;
  wire v8b555f;
  wire v8af461;
  wire v8b5813;
  wire v8573cf;
  wire v8e1f0d;
  wire v85aef4;
  wire v8e4792;
  wire v8af47b;
  wire v8e5022;
  wire v85f340;
  wire v8e58fa;
  wire v85d428;
  wire v856473;
  wire v889350;
  wire v8b569c;
  wire v8e4267;
  wire v8e3c83;
  wire v8e5a23;
  wire v865772;
  wire v8e1956;
  wire v85d9d8;
  wire v8b580f;
  wire v8b5683;
  wire v8b58ab;
  wire v881bc6;
  wire v8b35f0;
  wire v844fe7;
  wire v8b585a;
  wire v8b5756;
  wire v8b5801;
  wire v8892a8;
  wire v85da46;
  wire v8dc673;
  wire v85c9fb;
  wire v8af4c2;
  wire v8dc554;
  wire v889290;
  wire v85a10a;
  wire v8e4e02;
  wire v845047;
  wire v85c754;
  wire v85fa42;
  wire v8b57fa;
  wire v85696e;
  wire v8af26f;
  wire v863db8;
  wire v8e1a88;
  wire v8b55db;
  wire v8e4be4;
  wire v8e4f00;
  wire v8e158b;
  wire v85695e;
  wire v865b8f;
  wire v8562d4;
  wire v85d7a6;
  wire v8e4941;
  wire v85dbf1;
  wire v889fea;
  wire v8e3f84;
  wire v8a5bcf;
  wire v85c469;
  wire v8e4188;
  wire v8e4913;
  wire v865d5b;
  wire v856255;
  wire v8e4b00;
  wire v85dd64;
  wire v857625;
  wire v8b57b2;
  wire v8e5244;
  wire v85fa63;
  wire v8e1a57;
  wire v85e836;
  wire v8e59ca;
  wire v8e593b;
  wire v8b57ce;
  wire v8a5bbf;
  wire v85e1dd;
  wire v85e332;
  wire v85ccb4;
  wire v85f8f2;
  wire v8a5c15;
  wire v8b554b;
  wire v88c2d2;
  wire v86b9f0;
  wire v8b55d4;
  wire v8e58c4;
  wire v8b5764;
  wire v8e1756;
  wire v8e49d3;
  wire v8e5799;
  wire v8e51ad;
  wire v8b58b3;
  wire v86299d;
  wire v8db83f;
  wire v85744d;
  wire v8b56a6;
  wire v8e48d8;
  wire v8b56e8;
  wire v856558;
  wire v85733c;
  wire v8b5796;
  wire v8b554a;
  wire v8b569f;
  wire v8e3fa0;
  wire v8e3a10;
  wire v8af185;
  wire v8b56a2;
  wire v8e1ed4;
  wire v8b5891;
  wire v8e20fa;
  wire v8e222b;
  wire v85ad10;
  wire v85d42f;
  wire v8e19b1;
  wire v8b55e1;
  wire v85b07e;
  wire v8b560e;
  wire v8b55c5;
  wire v8842d0;
  wire v8e5943;
  wire v8e2059;
  wire v8e58bd;
  wire v8ce3d5;
  wire v8e4db2;
  wire v8e1f19;
  wire v85f123;
  wire v8e4f56;
  wire v8991c9;
  wire v85670f;
  wire v8b56d2;
  wire v85dbad;
  wire v8e424e;
  wire v8e14e0;
  wire v8b5681;
  wire v8e5607;
  wire v85e5db;
  wire v8b5728;
  wire v8e16f2;
  wire v8e4638;
  wire v8b57b5;
  wire v85b6c8;
  wire v85afc8;
  wire v8b54d4;
  wire v89954f;
  wire v85db5c;
  wire v8672d0;
  wire v8b5893;
  wire v8e22c7;
  wire v8e4e4e;
  wire v8e58d8;
  wire v8e2431;
  wire v8e4391;
  wire v8e59b7;
  wire v8e479e;
  wire v84513a;
  wire v882429;
  wire v8b560a;
  wire v8e3977;
  wire v85e08e;
  wire v85d309;
  wire v8e1651;
  wire v856669;
  wire v8b556b;
  wire v8b5831;
  wire v86654a;
  wire v8e4c9d;
  wire v8572ac;
  wire v8e509c;
  wire v856a23;
  wire v8e3eb2;
  wire v8bf0c7;
  wire v8a87b4;
  wire v8af226;
  wire v8b550c;
  wire v8573f7;
  wire v8e5971;
  wire v86c74d;
  wire v85d7bd;
  wire v8e3e82;
  wire v8b5554;
  wire v8cce20;
  wire v8e4051;
  wire v8e552e;
  wire v85cbea;
  wire v85b5f6;
  wire v8b57f5;
  wire v8a9208;
  wire v85677f;
  wire v8e5b11;
  wire v8b576c;
  wire v8b5889;
  wire v845183;
  wire v8e58aa;
  wire v882bc3;
  wire v85aa18;
  wire v8e4a68;
  wire v8e14ab;
  wire v8e48d7;
  wire v856edf;
  wire v8b5672;
  wire v8e3db0;
  wire v8e1579;
  wire v8b35e8;
  wire v856556;
  wire v8e193b;
  wire v8b587e;
  wire v8b5626;
  wire v8e4c46;
  wire v8e4ece;
  wire v8b5721;
  wire v8e5979;
  wire v8b55a1;
  wire v8e1813;
  wire v85e942;
  wire v889f73;
  wire v8b5851;
  wire v8bf339;
  wire v8e502c;
  wire v884d71;
  wire v8e19c2;
  wire v8b5829;
  wire v85c5cf;
  wire v85c941;
  wire v8a6914;
  wire v84523d;
  wire v865827;
  wire v8e1810;
  wire v8e56ef;
  wire v86ce9d;
  wire v8e5367;
  wire v8b589b;
  wire v8e3b66;
  wire v8e5054;
  wire v8b5508;
  wire v8e4589;
  wire v85a0da;
  wire v85faba;
  wire v8e4bb0;
  wire v857549;
  wire v8b57e3;
  wire v8b54d9;
  wire v85acdb;
  wire v8e59db;
  wire v8dc59e;
  wire v8b5807;
  wire v8665a9;
  wire v8e3dec;
  wire v8e5173;
  wire v88424e;
  wire v8e583f;
  wire v8af268;
  wire v8b5836;
  wire v85649c;
  wire v85679b;
  wire v8e58d7;
  wire v8e4163;
  wire v856b4f;
  wire v8b5610;
  wire v8b57fb;
  wire v8e460d;
  wire v8b5827;
  wire v85f8fd;
  wire v8e59fb;
  wire v85e0a1;
  wire v85b400;
  wire v86d72e;
  wire v8b55b8;
  wire v8e3b75;
  wire v84523b;
  wire v880bdf;
  wire v8e5a7a;
  wire v8b57a5;
  wire v8b57be;
  wire v85b2e6;
  wire v85c8b5;
  wire v8e3ac5;
  wire v8e3c3e;
  wire v8e41df;
  wire v85b2d5;
  wire v8e41c1;
  wire v8b55ea;
  wire v8e59b9;
  wire v8e47e7;
  wire v845069;
  wire v8e1961;
  wire v8af355;
  wire v8b5795;
  wire v8b57fe;
  wire v8e4217;
  wire v85b2ae;
  wire v8e5678;
  wire v85b073;
  wire v856474;
  wire v8e1a8c;
  wire v85f57e;
  wire v8e1f55;
  wire v8e4a85;
  wire v85fa3e;
  wire v85f2ba;
  wire v8e5928;
  wire v8e4b68;
  wire v8e53c7;
  wire v8b56c3;
  wire v8b570c;
  wire v882156;
  wire v8e58a0;
  wire v85dcd6;
  wire v8b55e3;
  wire v845033;
  wire v85a880;
  wire v8b5805;
  wire v845136;
  wire v8b561b;
  wire v8e5a63;
  wire v8e3dad;
  wire v8af1e3;
  wire v8b552a;
  wire v885308;
  wire v8e1f43;
  wire v8e192f;
  wire v8b5533;
  wire v8b562a;
  wire v85e652;
  wire v8b54c1;
  wire v8e160f;
  wire v8e415b;
  wire v8570f0;
  wire v8569c1;
  wire v8b57b3;
  wire v85d3cc;
  wire v8cc909;
  wire v85d7e9;
  wire v8e58ef;
  wire v8b56e4;
  wire v84515d;
  wire v85660c;
  wire v8e4b4e;
  wire v8e58cf;
  wire v8e4e81;
  wire v8b5658;
  wire v8e1931;
  wire v85d2e8;
  wire v8e1ae8;
  wire v845109;
  wire v84518e;
  wire v8e4f99;
  wire v85dd7f;
  wire v86290f;
  wire v8b5743;
  wire v8e519d;
  wire v8b57f2;
  wire v8e47ef;
  wire v8e3b0a;
  wire v8e1934;
  wire v8b54c4;
  wire v8e4832;
  wire v8e199a;
  wire v8e59e7;
  wire v85e7f0;
  wire v85c73b;
  wire v8b578f;
  wire v880b12;
  wire v8e2440;
  wire v8e5569;
  wire v8dc555;
  wire v8e1667;
  wire v8451b6;
  wire v8e55cf;
  wire v8e535e;
  wire v8812e9;
  wire v8e432e;
  wire v85626a;
  wire v8e15a0;
  wire v85aa15;
  wire v86824f;
  wire v8e527e;
  wire v8e51f4;
  wire v85f1cb;
  wire v856883;
  wire v8b5758;
  wire v8b56ec;
  wire v8b562e;
  wire v85d72c;
  wire v86654f;
  wire v8e5a3b;
  wire v85daa5;
  wire v8e38c7;
  wire v8e5960;
  wire v8e59e4;
  wire v8b587d;
  wire v8e46b8;
  wire v8e58f1;
  wire v8e1199;
  wire v856bc8;
  wire v8a5c52;
  wire v8e4eba;
  wire v8a881f;
  wire v8be142;
  wire v8b56fe;
  wire v8e469f;
  wire v8e16ce;
  wire v8cce79;
  wire v8e5a68;
  wire v8e58d3;
  wire v85df0b;
  wire v8564db;
  wire v8b56be;
  wire v8af21d;
  wire v8e3e66;
  wire v8b56e0;
  wire v85bbe5;
  wire v85d8ae;
  wire v85fa37;
  wire v8e4e15;
  wire v8e51d0;
  wire v8a5c58;
  wire v8e2079;
  wire v899224;
  wire v85e1f5;
  wire v8e5a61;
  wire v8be0f9;
  wire v8b5569;
  wire v85d3d0;
  wire v8ca185;
  wire v85dd3e;
  wire v8566f1;
  wire v8e3e49;
  wire v84507d;
  wire v8b54e9;
  wire v8e5a71;
  wire v8e5b2c;
  wire v88c2f2;
  wire v85c83d;
  wire v8e5a15;
  wire v8e240d;
  wire v85b6c9;
  wire v8b5775;
  wire v8b57f9;
  wire v85ce6f;
  wire v8e4d04;
  wire v85d3f6;
  wire v863508;
  wire v8e4c29;
  wire v8572b6;
  wire v8e59d6;
  wire v8563a6;
  wire v8e5252;
  wire v8e21a2;
  wire v8e3a7c;
  wire v8af3b8;
  wire v84510d;
  wire v85a4f0;
  wire v845101;
  wire v8e56ac;
  wire v8e4baa;
  wire v8e3926;
  wire v8e2144;
  wire v85760e;
  wire v85dfaa;
  wire v8e5b8b;
  wire v8b551c;
  wire v85724c;
  wire v8e1d49;
  wire v8e3fca;
  wire v85f567;
  wire v85d543;
  wire v8566fa;
  wire v8e42ab;
  wire v8e20ba;
  wire v85d750;
  wire v8b56d1;
  wire v8e21da;
  wire v8dc6c6;
  wire v844fbd;
  wire v8562d0;
  wire v844fa3;
  wire v85dfb7;
  wire v8cc8c3;
  wire v85f9b8;
  wire v8b5798;
  wire v860006;
  wire v860057;
  wire v8e17ae;
  wire v8e598e;
  wire v8e1cd8;
  wire v86514d;
  wire v8e4fe9;
  wire v85da5d;
  wire v8e5967;
  wire v85d8ba;
  wire v85e2b5;
  wire v856ef1;
  wire v85f5a7;
  wire v87f854;
  wire v85b036;
  wire v8b5863;
  wire v85dd7c;
  wire v8b5696;
  wire v8b5621;
  wire v85dcf5;
  wire v8be101;
  wire v8565ce;
  wire v8b5857;
  wire v8e4617;
  wire v85e0e3;
  wire v85f816;
  wire v85f4e0;
  wire v8e596c;
  wire v85dba0;
  wire v8e5606;
  wire v85631f;
  wire v8e51f8;
  wire v8e2177;
  wire v8e58b3;
  wire v8b5892;
  wire v8e1985;
  wire v8e4ac8;
  wire v8b568f;
  wire v8e2416;
  wire v889f3b;
  wire v86658f;
  wire v883cc4;
  wire v85da2e;
  wire v8e3a74;
  wire v8e5a0b;
  wire v845245;
  wire v8b568d;
  wire v845230;
  wire v8e1c12;
  wire v8e4255;
  wire v85c1d4;
  wire v86531f;
  wire v8b57c8;
  wire v8dc5e7;
  wire v8e593f;
  wire v861611;
  wire v86c2d3;
  wire v8dc55f;
  wire v8e58dd;
  wire v85769d;
  wire v85db04;
  wire v8e4d94;
  wire v8b5830;
  wire v8e5a76;
  wire v8e3bba;
  wire v857542;
  wire v857309;
  wire v8e47f9;
  wire v8563b7;
  wire v8b58aa;
  wire v8b54e1;
  wire v8e53ec;
  wire v8b5678;
  wire v8a923a;
  wire v867c19;
  wire v8b55a5;
  wire v85d6fe;
  wire v8e5a82;
  wire v8e5a5a;
  wire v8e579b;
  wire v8e5958;
  wire v880b6e;
  wire v8af12b;
  wire v85d6ea;
  wire v8b5645;
  wire v8e3992;
  wire v8b5659;
  wire v8e59ae;
  wire v845064;
  wire v85664e;
  wire v8af2f2;
  wire v8b574d;
  wire v8e4071;
  wire v85e1fe;
  wire v8af4b7;
  wire v8b569b;
  wire v84501d;
  wire v8e3d66;
  wire v8e5a19;
  wire v85d3b1;
  wire v8e44ed;
  wire v8af480;
  wire v8e591c;
  wire v84521e;
  wire v8b5613;
  wire v8cce8a;
  wire v844faf;
  wire v8b55bd;
  wire v85afc0;
  wire v8b5607;
  wire v844f95;
  wire v85de51;
  wire v883b69;
  wire v8565a3;
  wire v8e3899;
  wire v8b5501;
  wire v8e1c72;
  wire v8b5666;
  wire v85f52f;
  wire v8e17fe;
  wire v8e1d09;
  wire v8b55ac;
  wire v8e1f1b;
  wire v8e3cfe;
  wire v8e436f;
  wire v8e48fc;
  wire v8e240e;
  wire v85ae46;
  wire v85c73d;
  wire v85e3d2;
  wire v85deeb;
  wire v8e598d;
  wire v8a54e5;
  wire v8b5879;
  wire v8e2381;
  wire v8b5786;
  wire v8e40df;
  wire v8b5765;
  wire v8af23a;
  wire v8b55bf;
  wire v8e162c;
  wire v8b57d5;
  wire v85d805;
  wire v8664e6;
  wire v860007;
  wire v8e4040;
  wire v85e66e;
  wire v8e5861;
  wire v8e549e;
  wire v856f8d;
  wire v8b5860;
  wire v85e1e9;
  wire v866503;
  wire v8be0f6;
  wire v8e594c;
  wire v8af46d;
  wire v8b5778;
  wire v86e38c;
  wire v88c32e;
  wire v84535e;
  wire v8e5956;
  wire v8e4c6e;
  wire v8e41ae;
  wire v8b5727;
  wire v8b5609;
  wire v88486d;
  wire v865d55;
  wire v85fac2;
  wire v85f48a;
  wire v8e4be1;
  wire v8b55a6;
  wire v85ccc2;
  wire v86d019;
  wire v8b56f8;
  wire v8b5792;
  wire v8e4142;
  wire v8e59d5;
  wire v85b49f;
  wire v8e1ccb;
  wire v8e58e4;
  wire v8e1b90;
  wire v85a23c;
  wire v856fc9;
  wire v88c2be;
  wire v8e5060;
  wire v8e21d3;
  wire v8af37d;
  wire v85722b;
  wire v85c47d;
  wire v8e5242;
  wire v8e41db;
  wire v8a5bcc;
  wire v85dcee;
  wire v8e41d0;
  wire v8e176c;
  wire v85b514;
  wire v8564ef;
  wire v8e5b7d;
  wire v85f34e;
  wire v85ad1a;
  wire v8e4ba8;
  wire v85d8ad;
  wire v8e1eab;
  wire v860902;
  wire v8e4cfe;
  wire v85b2bc;
  wire v8b5586;
  wire v8e22d4;
  wire v8e59de;
  wire v8e531e;
  wire v85e8bf;
  wire v8565fe;
  wire v884319;
  wire v85deb3;
  wire v8e1abd;
  wire v8e1765;
  wire v8831e7;
  wire v85db08;
  wire v8e5a43;
  wire v8b588e;
  wire v8b572e;
  wire v8e3bee;
  wire v862719;
  wire v8e539f;
  wire v85dcb9;
  wire v8b54fa;
  wire v8bf8d8;
  wire v8b562f;
  wire v8b58ad;
  wire v8b572a;
  wire v8af29a;
  wire v8b57e2;
  wire v85db26;
  wire v8e5753;
  wire v8e415a;
  wire v8e4877;
  wire v8e1770;
  wire v85bbb8;
  wire v85c7af;
  wire v85a9b1;
  wire v8b5555;
  wire v8b55d2;
  wire v8af102;
  wire v8af40a;
  wire v85b5f8;
  wire v8b58ba;
  wire v8e4dbe;
  wire v8b578a;
  wire v8e1be0;
  wire v8e5881;
  wire v8e3fce;
  wire v8b5665;
  wire v8e1778;
  wire v8b54ed;
  wire v85668b;
  wire v8e3b74;
  wire v85666e;
  wire v85b906;
  wire v857423;
  wire v8be173;
  wire v8e57a1;
  wire v866511;
  wire v8b5776;
  wire v8e1eb3;
  wire v8a8877;
  wire v8b5880;
  wire v8e4e6e;
  wire v859fe9;
  wire v8e436b;
  wire v8b58bb;
  wire v8b552b;
  wire v8b54e8;
  wire v88c324;
  wire v8e5a48;
  wire v85b04f;
  wire v8b56d7;
  wire v8e4fe5;
  wire v8e3bda;
  wire v8e57c9;
  wire v8b586b;
  wire v85d79a;
  wire v8e4805;
  wire v8e54cf;
  wire v8b55ed;
  wire v8af457;
  wire v856653;
  wire v85f27b;
  wire v8b55e9;
  wire v8b5585;
  wire v85d6b7;
  wire v8dc5b0;
  wire v8e4468;
  wire v88c326;
  wire v85de64;
  wire v8b5806;
  wire v8b563d;
  wire v8e5939;
  wire v8e1b05;
  wire v8af4aa;
  wire v8b5548;
  wire v85737f;
  wire v8b5542;
  wire v8e4aec;
  wire v8b5762;
  wire v88bcc8;
  wire v8e58e6;
  wire v86c874;
  wire v8cf0f4;
  wire v8e3cb6;
  wire v857540;
  wire v85a24b;
  wire v8be150;
  wire v85673d;
  wire v8e5883;
  wire v8e5957;
  wire v8e59aa;
  wire v8450f2;
  wire v8b57d3;
  wire v8e5973;
  wire v8584f3;
  wire v86ea54;
  wire v8a5bc5;
  wire v8b55a9;
  wire v8e1da5;
  wire v88c2e1;
  wire v8e4172;
  wire v8e4f40;
  wire v86349c;
  wire v8e42dc;
  wire v8b57d8;
  wire v85dc0d;
  wire v8e5bbe;
  wire v8b57de;
  wire v8af147;
  wire v8e242d;
  wire v85a622;
  wire v8b5624;
  wire v8af31b;
  wire v85f647;
  wire v8b56a0;
  wire v8562ab;
  wire v8a554b;
  wire v8e4976;
  wire v85e152;
  wire v8e3979;
  wire v85db39;
  wire v8e1664;
  wire v89b6ce;
  wire v86e551;
  wire v856d2f;
  wire v8b5627;
  wire v85aad0;
  wire v8e222f;
  wire v8563e4;
  wire v8e520d;
  wire v88bc46;
  wire v8e5a5f;
  wire v8e5913;
  wire v8e548f;
  wire v8e1a78;
  wire v8a691b;
  wire v8e44c7;
  wire v85d914;
  wire v8562f2;
  wire v8b578b;
  wire v85cd17;
  wire v8af4a4;
  wire v861da7;
  wire v8892d9;
  wire v88928c;
  wire v8e38b1;
  wire v856345;
  wire v856eb9;
  wire v8e4f36;
  wire v856a21;
  wire v8e56cb;
  wire v8e159f;
  wire v8b5816;
  wire v8e22f8;
  wire v85a648;
  wire v8dc5b6;
  wire v8b57ab;
  wire v8e5049;
  wire v8a880e;
  wire v8bf437;
  wire v8e2154;
  wire v857144;
  wire v856275;
  wire v85e0c2;
  wire v8b5846;
  wire v8568a8;
  wire v88c2c2;
  wire v8565e5;
  wire v8b56db;
  wire v8606a9;
  wire v8e44f7;
  wire v865121;
  wire v8e5c69;
  wire v85e60f;
  wire v86bbca;
  wire v85b512;
  wire v8af4c4;
  wire v8e2098;
  wire v8e3c65;
  wire v8b564f;
  wire v85a4be;
  wire v8e55ba;
  wire v85ffb3;
  wire v85ddb8;
  wire v8b567f;
  wire v8e1823;
  wire v8b555a;
  wire v8e5968;
  wire v8e1d21;
  wire v86d0c6;
  wire v8e3af6;
  wire v8e4dae;
  wire v8caee0;
  wire v85fc4e;
  wire v864971;
  wire v85e8b5;
  wire v8a5b1b;
  wire v8b587b;
  wire v8e55ef;
  wire v8af1a3;
  wire v8991fe;
  wire v8e511b;
  wire v856f89;
  wire v85c895;
  wire v85735b;
  wire v8e23ce;
  wire v8892c0;
  wire v8e587b;
  wire v8e5588;
  wire v8e43dc;
  wire v85696d;
  wire v8af2be;
  wire v8b55a0;
  wire v8af19b;
  wire v889f94;
  wire v85c93d;
  wire v8e5a6a;
  wire v8e40af;
  wire v856cac;
  wire v85f4fb;
  wire v8a87fd;
  wire v856358;
  wire v8b583c;
  wire v8e3e1e;
  wire v8e57a4;
  wire v85db1a;
  wire v8b575b;
  wire v889f8a;
  wire v8e57a6;
  wire v8e59ec;
  wire v8e181b;
  wire v8e58b7;
  wire v8892cb;
  wire v8e4b6f;
  wire v8e56dd;
  wire v8b56ff;
  wire v8e14ca;
  wire v8e41a5;
  wire v856314;
  wire v8e5985;
  wire v8dc571;
  wire v85fbec;
  wire v8e3aa7;
  wire v85c436;
  wire v85f2a6;
  wire v85f839;
  wire v8b58b1;
  wire v856c6c;
  wire v8e39eb;
  wire v8e197c;
  wire v85f8da;
  wire v85cdde;
  wire v861ca6;
  wire v8a887e;
  wire v8e501a;
  wire v856312;
  wire v85b863;
  wire v85b69f;
  wire v8e3b8b;
  wire v8e4f5f;
  wire v8572d0;
  wire v857499;
  wire v8e2265;
  wire v8b5722;
  wire v8e5a2c;
  wire v8e15b2;
  wire v8e57ab;
  wire v856386;
  wire v8b558a;
  wire v8e40f6;
  wire v85b6b7;
  wire v85e548;
  wire v85da91;
  wire v85a0d2;
  wire v881da6;
  wire v8af188;
  wire v8e57d8;
  wire v8e58ed;
  wire v8b5704;
  wire v8e3eb5;
  wire v8e109f;
  wire v8b566b;
  wire v8e59a8;
  wire v85a893;
  wire v85dcb8;
  wire v8af432;
  wire v8e4103;
  wire v8e503e;
  wire v8e16e1;
  wire v85f5cc;
  wire v8dc6c4;
  wire v8e550e;
  wire v867aa7;
  wire v8e59f6;
  wire v8af418;
  wire v85725c;
  wire v8e4632;
  wire v8b5823;
  wire v85e0b0;
  wire v85e237;
  wire v85a4fc;
  wire v8b557e;
  wire v8e3c2f;
  wire v889264;
  wire v8e3a9d;
  wire v85f230;
  wire v8567ae;
  wire v8569ee;
  wire v8e4235;
  wire v8452fa;
  wire v85f448;
  wire v85d59f;
  wire v84521c;
  wire v88e287;
  wire v8bf8d3;
  wire v85d5b1;
  wire v8e46ed;
  wire v8b57cc;
  wire v865897;
  wire v8b54fc;
  wire v85b0a3;
  wire v85e61d;
  wire v85d860;
  wire v8e47d6;
  wire v8b5674;
  wire v8dc57c;
  wire v8e54a4;
  wire v85e887;
  wire v85ccec;
  wire v889ec1;
  wire v85a0f8;
  wire v8e43ad;
  wire v8e59c7;
  wire v8e5692;
  wire v8e4270;
  wire v856367;
  wire v8575eb;
  wire v8b5733;
  wire v881a3e;
  wire v8e10ed;
  wire v8e1a2e;
  wire v85e694;
  wire v8e1f76;
  wire v85d971;
  wire v8b56ba;
  wire v8e201e;
  wire v8b553c;
  wire v8b56d3;
  wire v8e44c8;
  wire v8b5595;
  wire v8dc5cb;
  wire v8e207d;
  wire v85a51b;
  wire v8564de;
  wire v845351;
  wire v8e2045;
  wire v8e438b;
  wire v8af383;
  wire v8b5862;
  wire v8892b3;
  wire v88926c;
  wire v8e40a5;
  wire v85d9d4;
  wire v856443;
  wire v8e4761;
  wire v8b5689;
  wire v856f08;
  wire v8b5656;
  wire v8e57e7;
  wire v8af493;
  wire v845039;
  wire v8635e4;
  wire v8af0dc;
  wire v8e23c6;
  wire v85d53f;
  wire v88924d;
  wire v85afea;
  wire v8e1b8d;
  wire v8e46b2;
  wire v8e5650;
  wire v8e5075;
  wire v8e4d85;
  wire v8b581e;
  wire v8b577c;
  wire v8e5a31;
  wire v85e9ee;
  wire v8e1480;
  wire v8e4d8f;
  wire v8e1c87;
  wire v8e460c;
  wire v8e4229;
  wire v87c63e;
  wire v880b52;
  wire v8e5a55;
  wire v8e4cc0;
  wire v8e4588;
  wire v8e1d32;
  wire v860064;
  wire v8e51cf;
  wire v859fe5;
  wire v85afbc;
  wire v8e57ee;
  wire v8e2091;
  wire v85ace0;
  wire v8cafe0;
  wire v8e5936;
  wire v8e493e;
  wire v8e45c9;
  wire v8e3ffc;
  wire v8e1dbf;
  wire v85cc98;
  wire v8dc575;
  wire v8564c4;
  wire v857056;
  wire v8b584e;
  wire v8e492c;
  wire v85db90;
  wire v85f422;
  wire v8e1f2a;
  wire v8e1df8;
  wire v85dbf8;
  wire v856eeb;
  wire v85684d;
  wire v85e0b5;
  wire v8e5a00;
  wire v8b553f;
  wire v8a5bfd;
  wire v8b54de;
  wire v8b5640;
  wire v8b55fc;
  wire v8e5a01;
  wire v85db0d;
  wire v8e4d0d;
  wire v8b589d;
  wire v8dc65c;
  wire v8650b9;
  wire v8b5883;
  wire v8e1c1c;
  wire v8b55dd;
  wire v8e428a;
  wire v8e4a30;
  wire v8e1f8f;
  wire v8af330;
  wire v8a5cb3;
  wire v85a88e;
  wire v8e59d3;
  wire v8cc8f2;
  wire v8e1f47;
  wire v8e55d6;
  wire v8e53be;
  wire v8a5c2d;
  wire v85b5bc;
  wire v8b5859;
  wire v85f953;
  wire v85a0ae;
  wire v8af231;
  wire v8e10fb;
  wire v8e20a4;
  wire v8b55c7;
  wire v8e541f;
  wire v88c2f6;
  wire v8dc5de;
  wire v85761b;
  wire v8cce37;
  wire v8b5838;
  wire v85db8a;
  wire v8e5a3e;
  wire v880bc4;
  wire v8b5557;
  wire v8af18b;
  wire v8b57ea;
  wire v8b5719;
  wire v8cc8ad;
  wire v8e20e3;
  wire v8563be;
  wire v85d34c;
  wire v8e595b;
  wire v8b579c;
  wire v85f427;
  wire v8dc606;
  wire v8e229e;
  wire v8e1718;
  wire v856fbd;
  wire v8b54dc;
  wire v85cccf;
  wire v858f70;
  wire v8e39e6;
  wire v85f814;
  wire v8e4a57;
  wire v85dbf7;
  wire v8b54c2;
  wire v8e3cd1;
  wire v8b5679;
  wire v8be0ea;
  wire v8e5a5c;
  wire v861ed7;
  wire v8e2229;
  wire v8e5a11;
  wire v8e58ec;
  wire v8b54eb;
  wire v8b572c;
  wire v8e5880;
  wire v8e5698;
  wire v845360;
  wire v889ec2;
  wire v8b5800;
  wire v856598;
  wire v85a05d;
  wire v8e3d83;
  wire v85d98f;
  wire v8e59f9;
  wire v8b5643;
  wire v8b56fb;
  wire v8b5897;
  wire v856b0d;
  wire v85d6ab;
  wire v85cb88;
  wire v856479;
  wire v85cc56;
  wire v85a0bf;
  wire v85acfd;
  wire v859ffb;
  wire v85d376;
  wire v8dc5ab;
  wire v85e951;
  wire v8e47f8;
  wire v8e5498;
  wire v8e229f;
  wire v85db87;
  wire v8b5712;
  wire v845386;
  wire v88927c;
  wire v8cc95a;
  wire v8e59c5;
  wire v8e1aa8;
  wire v85726b;
  wire v856be5;
  wire v8b56bb;
  wire v8b5670;
  wire v88c3ad;
  wire v8e463e;
  wire v8a5b9b;
  wire v8e38c8;
  wire v8e3ab5;
  wire v8b582d;
  wire v8b566d;
  wire v85f170;
  wire v8e2147;
  wire v889244;
  wire v856261;
  wire v858981;
  wire v8e1c7f;
  wire v8e4f78;
  wire v8e431c;
  wire v8b55ec;
  wire v85ccc6;
  wire v8e5950;
  wire v8e17a8;
  wire v8b576a;
  wire v85c77b;
  wire v8e3fe8;
  wire v85bd3d;
  wire v856404;
  wire v8e39e1;
  wire v8e4514;
  wire v8e4c47;
  wire v85e091;
  wire v8b56e6;
  wire v85de53;
  wire v85dfab;
  wire v8dc5ff;
  wire v85c7c5;
  wire v8e5946;
  wire v8e3df4;
  wire v865833;
  wire v85de34;
  wire v85e18a;
  wire v85b6b5;
  wire v85f2c8;
  wire v86007f;
  wire v865131;
  wire v8e1654;
  wire v8e396e;
  wire v8e1cd3;
  wire v85e8fd;
  wire v8e58b4;
  wire v8e595d;
  wire v85f594;
  wire v8e1f73;
  wire v8af34b;
  wire v85b938;
  wire v8e5a84;
  wire v8cdce6;
  wire v8e2000;
  wire v8452cd;
  wire v8e197f;
  wire v863b23;
  wire v85e565;
  wire v85d434;
  wire v8e1a5a;
  wire v856a1f;
  wire v85ad82;
  wire v8e18dd;
  wire v8e3f79;
  wire v85d671;
  wire v8b5856;
  wire v8e1d99;
  wire v8e5977;
  wire v889fde;
  wire v8e462b;
  wire v856663;
  wire v8b586a;
  wire v8e22fd;
  wire v8e50df;
  wire v85d314;
  wire v85a153;
  wire v8e239b;
  wire v85fc09;
  wire v8b5872;
  wire v8e53c6;
  wire v8e4cfc;
  wire v8b57e0;
  wire v8e15a4;
  wire v8b5549;
  wire v85c80b;
  wire v8cce52;
  wire v8e1e0e;
  wire v85cbd3;
  wire v8e4a06;
  wire v88c31b;
  wire v8b55f8;
  wire v8be124;
  wire v8e5aa0;
  wire v8b57e9;
  wire v8e3d20;
  wire v8e17e6;
  wire v8cce02;
  wire v8892b6;
  wire v889ec0;
  wire v8e51e4;
  wire v8e4ffe;
  wire v8e1f66;
  wire v856ecb;
  wire v8e5366;
  wire v85c639;
  wire v8e50a2;
  wire v8e597e;
  wire v8e1abc;
  wire v8e1a74;
  wire v8b54c5;
  wire v8e3b4c;
  wire v8e1692;
  wire v8b5852;
  wire v85d90a;
  wire v8e42fe;
  wire v8b56d6;
  wire v8e477d;
  wire v8b5793;
  wire v8e5a22;
  wire v8b56c8;
  wire v856fe9;
  wire v8e469a;
  wire v8e214e;
  wire v85b1c3;
  wire v857010;
  wire v8e436c;
  wire v85abc1;
  wire v85c96a;
  wire v8e4050;
  wire v8e4184;
  wire v86bf1f;
  wire v8e1c07;
  wire v8e4d32;
  wire v85655b;
  wire v8e188a;
  wire v8e38c3;
  wire v8e57f0;
  wire v8e5887;
  wire v8e3de0;
  wire v8e5a5e;
  wire v85ea90;
  wire v8e3ec6;
  wire v8e4f37;
  wire v85aa47;
  wire v8b57ef;
  wire v8567a3;
  wire v856481;
  wire v8e1b83;
  wire v85e80e;
  wire v8b5754;
  wire v857578;
  wire v8b586f;
  wire v8e566a;
  wire v8b563f;
  wire v8e51c8;
  wire v8e3d2a;
  wire v85ac27;
  wire v884bb3;
  wire v85e27e;
  wire v85af8a;
  wire v86583e;
  wire v8566fb;
  wire v85de73;
  wire v8b5648;
  wire v8e3a58;
  wire v8e45ab;
  wire v8e1ec6;
  wire v8e591f;
  wire v8563b6;
  wire v8b54c6;
  wire v85a3a4;
  wire v8e1c27;
  wire v8e1995;
  wire v8e10c3;
  wire v856c3d;
  wire v8e589a;
  wire v85b4e6;
  wire v8e3c75;
  wire v856705;
  wire v8b5567;
  wire v85e362;
  wire v8e4118;
  wire v8e5085;
  wire v856390;
  wire v8b5571;
  wire v8e4b9f;
  wire v85fb1e;
  wire v8b5832;
  wire v8b571e;
  wire v8e21c8;
  wire v8e4d59;
  wire v85e68a;
  wire v899550;
  wire v856cd5;
  wire v8b5644;
  wire v85ffdf;
  wire v8e20a2;
  wire v8e5a69;
  wire v8b54d1;
  wire v8e5600;
  wire v8e5c2a;
  wire v8e1f7e;
  wire v8b5896;
  wire v867a85;
  wire v8450f8;
  wire v8e1504;
  wire v8cc8ae;
  wire v8e5a62;
  wire v85d8e2;
  wire v85e99d;
  wire v8b55f2;
  wire v8e3e83;
  wire v85b57e;
  wire v8e568f;
  wire v856688;
  wire v85b540;
  wire v8e5b0d;
  wire v86e828;
  wire v8b572f;
  wire v8e1eb4;
  wire v84518f;
  wire v8e22c3;
  wire v8452dc;
  wire v8b35f5;
  wire v85da56;
  wire v8dc551;
  wire v85fa41;
  wire v85c73e;
  wire v856a93;
  wire v8672c1;
  wire v8e46d9;
  wire v8b5605;
  wire v8e3ff2;
  wire v8563c0;
  wire v8e1abe;
  wire v856be2;
  wire v857037;
  wire v8b5686;
  wire v8e1d00;
  wire v8e3b87;
  wire v856cb3;
  wire v8e22bd;
  wire v8e1f74;
  wire v8b55e8;
  wire v8e1bf5;
  wire v8e5769;
  wire v8b5559;
  wire v8b55b1;
  wire v8e43fa;
  wire v8e420f;
  wire v8b5847;
  wire v8e212b;
  wire v8e5a6f;
  wire v85d533;
  wire v85767e;
  wire v88934e;
  wire v8e44d9;
  wire v8e1c96;
  wire v85b06b;
  wire v85c4b8;
  wire v8e3bef;
  wire v861740;
  wire v8cce14;
  wire v845268;
  wire v85df25;
  wire v8a6d22;
  wire v8e4791;
  wire v85d382;
  wire v8e5907;
  wire v8e18fe;
  wire v8e1590;
  wire v8e44dd;
  wire v8b57da;
  wire v856b8f;
  wire v8e544a;
  wire v89920a;
  wire v856466;
  wire v8e417e;
  wire v85f697;
  wire v8b58ae;
  wire v85650e;
  wire v8e2282;
  wire v845380;
  wire v8dc593;
  wire v8e4c41;
  wire v8e3ea2;
  wire v8e4ebc;
  wire v85724d;
  wire v8819a3;
  wire v8b35f2;
  wire v8691fd;
  wire v8e1b00;
  wire v8b570e;
  wire v85e3a8;
  wire v85c47a;
  wire v863949;
  wire v856bc1;
  wire v8b586c;
  wire v87356b;
  wire v8e44a9;
  wire v8b57ae;
  wire v8e1e6c;
  wire v8892bc;
  wire v8e38a7;
  wire v8e58d5;
  wire v8b567b;
  wire v85de0b;
  wire v8b556d;
  wire v85b54e;
  wire v8e1638;
  wire v85ba99;
  wire v8e1cc4;
  wire v88c38a;
  wire v8b55c3;
  wire v8571d6;
  wire v85d9f0;
  wire v8e3b2f;
  wire v85e272;
  wire v8e114b;
  wire v8e58b8;
  wire v8e5a56;
  wire v8e2475;
  wire v8e1d80;
  wire v8cce39;
  wire v85cbe8;
  wire v8e5a13;
  wire v856364;
  wire v856b8e;
  wire v8b5858;
  wire v8af3e3;
  wire v8e4b49;
  wire v8992c3;
  wire v8e5a9d;
  wire v8e21d0;
  wire v8e4e45;
  wire v856ca7;
  wire v856e1f;
  wire v85deb5;
  wire v8e3df8;
  wire v85ad62;
  wire v8e58a6;
  wire v8b58b7;
  wire v85da0f;
  wire v8e4007;
  wire v8b5589;
  wire v8e55ca;
  wire v85e45f;
  wire v8e5494;
  wire v899247;
  wire v8e5a39;
  wire v85ca01;
  wire v8dc612;
  wire v8e388a;
  wire v85a98f;
  wire v85ccc4;
  wire v85ca3a;
  wire v8e4a22;
  wire v8e23ae;
  wire v856b6d;
  wire v85b5d9;
  wire v85d539;
  wire v8e22ae;
  wire v8e41c2;
  wire v85ffb2;
  wire v85638e;
  wire v856eca;
  wire v8e14db;
  wire v85f64e;
  wire v85659c;
  wire v86b6cf;
  wire v8e55a3;
  wire v8b5625;
  wire v8b5839;
  wire v8dc5d8;
  wire v8e1893;
  wire v8e41a7;
  wire v8e565f;
  wire v8b584c;
  wire v8e10c0;
  wire v8b57c6;
  wire v8b55fa;
  wire v8ccdf5;
  wire v8dc60e;
  wire v8562b8;
  wire v8e1811;
  wire v8e10f9;
  wire v8e59b4;
  wire v8e57dd;
  wire v8e5a2a;
  wire v85c7b4;
  wire v8b5515;
  wire v8b55e7;
  wire v8b55d1;
  wire v8e4f8b;
  wire v8e20f6;
  wire v8af419;
  wire v8b55c0;
  wire v8e4e95;
  wire v8e484a;
  wire v85bbe2;
  wire v8b588f;
  wire v85ddc7;
  wire v8e5266;
  wire v85d340;
  wire v85a34c;
  wire v8574cc;
  wire v8e5212;
  wire v8e5897;
  wire v8e5468;
  wire v85b979;
  wire v8892c1;
  wire v85d933;
  wire v8e5aa8;
  wire v856bd4;
  wire v8b5611;
  wire v8e152b;
  wire v8e200b;
  wire v8e42b2;
  wire v85fa64;
  wire v85a1f0;
  wire v8af2da;
  wire v8e5a78;
  wire v8e3b4b;
  wire v8e38ea;
  wire v8b56b3;
  wire v8dc56c;
  wire v8b56c2;
  wire v8833ba;
  wire v867398;
  wire v8e53de;
  wire v8b557d;
  wire v8e23a9;
  wire v8af213;
  wire v880b59;
  wire v86650a;
  wire v8e3d3c;
  wire v8e1c84;
  wire v85e274;
  wire v8b55bc;
  wire v85688c;
  wire v862c12;
  wire v8e5ad2;
  wire v8564ad;
  wire v8e3dac;
  wire v8e2373;
  wire v8e42b6;
  wire v85b3a4;
  wire v85adad;
  wire v8e1bb4;
  wire v8b567a;
  wire v8e1aea;
  wire v8b576e;
  wire v8dc639;
  wire v8be167;
  wire v8e4a8a;
  wire v85d45f;
  wire v883ca1;
  wire v85fbed;
  wire v8e1484;
  wire v877314;
  wire v8b5745;
  wire v8e5098;
  wire v885465;
  wire v8e58a7;
  wire v85d7c8;
  wire v8e57d0;
  wire v8665a0;
  wire v8567d9;
  wire v8a5552;
  wire v8e4a83;
  wire v889f95;
  wire v8b5596;
  wire v8e3e0e;
  wire v85dbd4;
  wire v8e1618;
  wire v8e4eef;
  wire v87d771;
  wire v8b5761;
  wire v8e572b;
  wire v8846fb;
  wire v8672c7;
  wire v856ba0;
  wire v8b5649;
  wire v8e19b2;
  wire v8e4872;
  wire v8e5a9f;
  wire v88c2fb;
  wire v8e49eb;
  wire v8b5558;
  wire v8b5822;
  wire v8e21d1;
  wire v85ce72;
  wire v8e1e94;
  wire v880bc3;
  wire v85e81e;
  wire v8e2239;
  wire v86ed0b;
  wire v8e3f4c;
  wire v8e205f;
  wire v85d598;
  wire v8e4e0e;
  wire v8e543c;
  wire v899261;
  wire v8b569a;
  wire v8b561f;
  wire v85663a;
  wire v8e5a6e;
  wire v856dbe;
  wire v8cce0a;
  wire v8e5909;
  wire v8e5364;
  wire v85a990;
  wire v8e1e59;
  wire v8e1c8a;
  wire v8b55f7;
  wire v8e1d7d;
  wire v8e4d9f;
  wire v8e4461;
  wire v8b5622;
  wire v87c649;
  wire v844fb5;
  wire v8e38d9;
  wire v85ad2e;
  wire v865125;
  wire v85cd1f;
  wire v8b56a3;
  wire v85ba14;
  wire v889f3d;
  wire v85fc4d;
  wire v8b56f7;
  wire v8e3f6f;
  wire v8e3ae7;
  wire v85630a;
  wire v8b552d;
  wire v8e4b0e;
  wire v8e1f85;
  wire v8e5889;
  wire v8b58b2;
  wire v8b5546;
  wire v856c90;
  wire v8b5614;
  wire v85fb12;
  wire v8658a0;
  wire v889f9b;
  wire v8569df;
  wire v8b54cb;
  wire v8e1c89;
  wire v8b57a6;
  wire v8e58b0;
  wire v856afe;
  wire v8b5522;
  wire v8e4ed1;
  wire v8e4eb5;
  wire v889f96;
  wire v85c8f2;
  wire v8e501b;
  wire v8b5600;
  wire v86972a;
  wire v85aea9;
  wire v8e4a95;
  wire v8dc617;
  wire v8e2436;
  wire v8e17b8;
  wire v85758c;
  wire v85b421;
  wire v8e5048;
  wire v8e564d;
  wire v8e2470;
  wire v85cea0;
  wire v845026;
  wire v8b5503;
  wire v8e238d;
  wire v8568c2;
  wire v856c62;
  wire v8e5259;
  wire v889e03;
  wire v85b3fb;
  wire v845060;
  wire v889fca;
  wire v8b5677;
  wire v8e3917;
  wire v8e484f;
  wire v8565ab;
  wire v8e5895;
  wire v85df05;
  wire v85708d;
  wire v85e4af;
  wire v8b55c6;
  wire v8e39c1;
  wire v85bdac;
  wire v85dd89;
  wire v8e233b;
  wire v8e488c;
  wire v8be147;
  wire v8b56cd;
  wire v85f4ff;
  wire v8e1d5f;
  wire v8569ce;
  wire v85630d;
  wire v85ba1d;
  wire v898498;
  wire v85dd75;
  wire v85c718;
  wire v8e441a;
  wire v857558;
  wire v8e2060;
  wire v8b5779;
  wire v8566b6;
  wire v8e4605;
  wire v8e164c;
  wire v8b55e4;
  wire v8e590b;
  wire v8e19e8;
  wire v8b56ed;
  wire v8e1ee5;
  wire v845079;
  wire v8b56f1;
  wire v85e82e;
  wire v8b583e;
  wire v8e1e0a;
  wire v8e47b7;
  wire v858ae4;
  wire v8e5b6b;
  wire v8e4cc7;
  wire v85b390;
  wire v85a6d2;
  wire v8b57ec;
  wire v8a5c22;
  wire v8e50d1;
  wire v8e58a1;
  wire v8e3bbb;
  wire v866593;
  wire v85d812;
  wire v8b5538;
  wire v856c2e;
  wire v8cb249;
  wire v8e3f1b;
  wire v8b57a0;
  wire v8e3bf7;
  wire v85da6c;
  wire v8e1cd2;
  wire v8af271;
  wire v8e58b6;
  wire v85e895;
  wire v8e5b6d;
  wire v8e1088;
  wire v8e16d2;
  wire v8e1ad8;
  wire v85bdbc;
  wire v8e58cd;
  wire v86d36d;
  wire v85a0f3;
  wire v8e5a18;
  wire v85e33b;
  wire v8e444a;
  wire v8451d1;
  wire v856ae7;
  wire v8e597b;
  wire v8b558c;
  wire v8b55d7;
  wire v8e5625;
  wire v8e583d;
  wire v8e420a;
  wire v85f1ac;
  wire v889f6e;
  wire v85e8f4;
  wire v85e8f2;
  wire v8e5b23;
  wire v8b5578;
  wire v85bbd9;
  wire v856b8b;
  wire v8e202c;
  wire v86cf33;
  wire v8840fd;
  wire v84520b;
  wire v8e17f5;
  wire v8e3c25;
  wire v8e4c34;
  wire v8e597f;
  wire v8e3bb9;
  wire v8e5b63;
  wire v85bd68;
  wire v85abc2;
  wire v8b5675;
  wire v8b551a;
  wire v85ba2c;
  wire v8b42e8;
  wire v8b57b8;
  wire v8e5903;
  wire v8af0de;
  wire v8b5731;
  wire v85ba47;
  wire v860037;
  wire v8e5930;
  wire v85f43b;
  wire v85f33d;
  wire v8b56a8;
  wire v85f244;
  wire v85df7f;
  wire v8a87f0;
  wire v8e19fd;
  wire v8e3dcc;
  wire v85da39;
  wire v883e72;
  wire v856c6d;
  wire v8e48a0;
  wire v8e58e8;
  wire v8a6968;
  wire v8e53b1;
  wire v865802;
  wire v8e19c3;
  wire v856c3c;
  wire v8e590d;
  wire v8b5697;
  wire v86b0d6;
  wire v88bc4c;
  wire v85b6e3;
  wire v85e618;
  wire v8e413b;
  wire v8b5873;
  wire v8e19c4;
  wire v8b56a5;
  wire v8e2399;
  wire v85e50d;
  wire v859fe4;
  wire v8a691d;
  wire v8e21cf;
  wire v8b57ad;
  wire v85e545;
  wire v8e4ea5;
  wire v8e4e56;
  wire v85b9a0;
  wire v8b54f2;
  wire v85ccdf;
  wire v8e19c7;
  wire v857139;
  wire v85e1bb;
  wire v85ce5c;
  wire v8ce34d;
  wire v889f4f;
  wire v8b5749;
  wire v8e4e99;
  wire v8a5b9d;
  wire v8e5069;
  wire v8e465f;
  wire v8e2213;
  wire v856fdc;
  wire v85dc21;
  wire v8e4bc9;
  wire v85a5e3;
  wire v8e15fd;
  wire v8e4599;
  wire v85ad0c;
  wire v8e1bf9;
  wire v85f6b4;
  wire v8e4d29;
  wire v85f2aa;
  wire v8e1e31;
  wire v856fba;
  wire v8e3ad8;
  wire v889f5a;
  wire v8af41e;
  wire v8b574f;
  wire v85eae6;
  wire v8e4f16;
  wire v85d57d;
  wire v8b550e;
  wire v8e58a8;
  wire v85d507;
  wire v8e20ac;
  wire v85dc22;
  wire v8e53d3;
  wire v8e5433;
  wire v8e45f1;
  wire v8e14ea;
  wire v8b5842;
  wire v8e38cd;
  wire v8b54f7;
  wire v85d2dd;
  wire v85a5eb;
  wire v8b5545;
  wire v8e39bb;
  wire v8680cc;
  wire v88bcc9;
  wire v8e48f1;
  wire v865dba;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg StoB_REQ4_p;
  input StoB_REQ4_n;
  reg StoB_REQ5_p;
  input StoB_REQ5_n;
  reg StoB_REQ6_p;
  input StoB_REQ6_n;
  reg StoB_REQ7_p;
  input StoB_REQ7_n;
  reg StoB_REQ8_p;
  input StoB_REQ8_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoS_ACK4_p;
  output BtoS_ACK4_n;
  reg BtoS_ACK5_p;
  output BtoS_ACK5_n;
  reg BtoS_ACK6_p;
  output BtoS_ACK6_n;
  reg BtoS_ACK7_p;
  output BtoS_ACK7_n;
  reg BtoS_ACK8_p;
  output BtoS_ACK8_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg SLC2_p;
  output SLC2_n;
  reg SLC3_p;
  output SLC3_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  reg jx3_p;
  output jx3_n;
  wire ENQ_n;
  wire SLC3_n;

assign v857943 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & v85cd1c;
assign v8db8b5 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v85ea8d;
assign v8be15d = jx0_p & v8af44d | !jx0_p & !v84507a;
assign v8e59b4 = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v8e10f9;
assign v8e2025 = jx2_p & v8574d6 | !jx2_p & v8571db;
assign v8e22fd = jx0_p & v8e4fad | !jx0_p & !v8b586a;
assign v8e54a4 = BtoS_ACK0_p & v8e550e | !BtoS_ACK0_p & v8dc57c;
assign v85c3e3 = BtoS_ACK0_p & v8e4637 | !BtoS_ACK0_p & v8450c0;
assign v8e5a07 = ENQ_p & v8e3a26 | !ENQ_p & v8e58d4;
assign v8585db = BtoS_ACK8_p & v86290d | !BtoS_ACK8_p & v844f91;
assign v8b5656 = BtoS_ACK6_p & v865897 | !BtoS_ACK6_p & v856f08;
assign v8e176c = jx2_p & v844f91 | !jx2_p & v8e41d0;
assign v8e5754 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8af243;
assign v8cf114 = BtoS_ACK0_p & v8e5a10 | !BtoS_ACK0_p & v85dbe7;
assign v8b5571 = StoB_REQ7_p & v86007f | !StoB_REQ7_p & v856390;
assign v86e828 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e5b0d;
assign v8b5546 = BtoS_ACK6_p & v8e3ae7 | !BtoS_ACK6_p & v8b58b2;
assign v8b5847 = BtoS_ACK6_p & v8e4f37 | !BtoS_ACK6_p & v8e420f;
assign v85767f = jx1_p & v85f42f | !jx1_p & v85e653;
assign v88c39f = jx1_p & v8b56ee | !jx1_p & v845150;
assign v8e3ad8 = BtoS_ACK8_p & v8e15fd | !BtoS_ACK8_p & v856fba;
assign v85a153 = jx0_p & v85d314 | !jx0_p & !v844f91;
assign v85aea9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86972a;
assign v85ad0c = BtoS_ACK7_p & v8e420a | !BtoS_ACK7_p & v8e4599;
assign v8e5971 = StoB_REQ1_p & v8e3d7b | !StoB_REQ1_p & v8573f7;
assign v8b571f = stateG12_p & v8b57a9 | !stateG12_p & v844f91;
assign v8e40a5 = StoB_REQ0_p & v8892b3 | !StoB_REQ0_p & v88926c;
assign v8e4a96 = StoB_REQ7_p & v8e2181 | !StoB_REQ7_p & v8e59e5;
assign v8e5959 = BtoS_ACK6_p & v8e58c2 | !BtoS_ACK6_p & v8e14dc;
assign BtoS_ACK8_n = v8bf910;
assign v8e5aa4 = jx0_p & v8b5698 | !jx0_p & v866552;
assign v8e5a2f = BtoS_ACK0_p & v86290d | !BtoS_ACK0_p & !v88d5d7;
assign v85dee5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e5033;
assign v8b5589 = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v8e4007;
assign v8e4dbe = jx1_p & v8b58ba | !jx1_p & v844f91;
assign v86583e = jx2_p & v85af8a | !jx2_p & v8e188a;
assign v85e905 = jx1_p & v86290d | !jx1_p & v85f2f8;
assign v8b54fc = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v857499;
assign v8b57f9 = StoB_REQ8_p & v8e5a61 | !StoB_REQ8_p & v8b5775;
assign v85dfb4 = StoB_REQ8_p & v8a8822 | !StoB_REQ8_p & v85da9f;
assign v85a990 = RtoB_ACK1_p & v8e543c | !RtoB_ACK1_p & !v8e5364;
assign v85ce5c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e1bb;
assign v8e5928 = BtoS_ACK1_p & v8e3d7b | !BtoS_ACK1_p & v85f2ba;
assign v867b8d = jx0_p & v8e4003 | !jx0_p & !v8e408d;
assign v8e3f65 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e2121;
assign v8e5a1f = jx1_p & v8e15ab | !jx1_p & v844f91;
assign v8e415b = BtoS_ACK2_p & v8b550c | !BtoS_ACK2_p & v8e160f;
assign v8e2355 = jx1_p & v8dc6a0 | !jx1_p & v85d3cb;
assign v85c436 = BtoS_ACK8_p & v856cac | !BtoS_ACK8_p & v8e3aa7;
assign v8a747c = jx1_p & v8572f7 | !jx1_p & !v88d5d7;
assign v88934e = EMPTY_p & v85767e | !EMPTY_p & v8b55f2;
assign v8e1da5 = BtoS_ACK0_p & v85de64 | !BtoS_ACK0_p & v8b55a9;
assign v8e3b87 = StoB_REQ2_p & v8b572f | !StoB_REQ2_p & v8e1d00;
assign v88c2f6 = BtoR_REQ0_p & v8e541f | !BtoR_REQ0_p & v8b55c7;
assign v8a5564 = jx3_p & v8e5c10 | !jx3_p & v8a5c04;
assign v8e5a66 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8e519b;
assign v8e4589 = StoB_REQ7_p & v8e5982 | !StoB_REQ7_p & v8e22c7;
assign v8af3db = ENQ_p & v8af46c | !ENQ_p & v8e5194;
assign v8e229f = jx2_p & v8e5498 | !jx2_p & v844f91;
assign v8b5820 = jx2_p & v8e5646 | !jx2_p & v86290d;
assign v85b2d5 = StoB_REQ7_p & v8e5a7a | !StoB_REQ7_p & v8e41df;
assign v8e44f7 = BtoS_ACK7_p & v85737f | !BtoS_ACK7_p & v8606a9;
assign v8e3899 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v844fb3 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v8450b6 = jx2_p & v85cb8e | !jx2_p & v844f91;
assign v8b55d2 = BtoS_ACK7_p & v85db26 | !BtoS_ACK7_p & v8b5555;
assign v8af160 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9b;
assign v8e3c27 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e39ff;
assign v88486d = BtoS_ACK7_p & v8e594c | !BtoS_ACK7_p & !v8b5609;
assign v85f8f2 = BtoS_ACK7_p & v856255 | !BtoS_ACK7_p & v85ccb4;
assign v85fac2 = BtoS_ACK8_p & v8e162c | !BtoS_ACK8_p & v865d55;
assign v8a54e5 = StoB_REQ6_p & v8e598d | !StoB_REQ6_p & v844f95;
assign v85d8ba = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v844f91;
assign v8b5754 = BtoS_ACK3_p & v8e16ea | !BtoS_ACK3_p & v8e3d20;
assign v8e5861 = StoB_REQ0_p & v8a54f3 | !StoB_REQ0_p & v844f91;
assign v8b56b2 = BtoS_ACK8_p & v8cc8e9 | !BtoS_ACK8_p & v85cdaa;
assign v85d98f = jx0_p & v8e3d83 | !jx0_p & !v844f91;
assign v8b56a5 = jx2_p & v8e19c4 | !jx2_p & !v8e238d;
assign v8af271 = BtoS_ACK0_p & v86972a | !BtoS_ACK0_p & v8e1cd2;
assign v8b5704 = BtoS_ACK7_p & v8e15b2 | !BtoS_ACK7_p & v8e58ed;
assign v88475f = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v8e40a9;
assign v8e4b64 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85e93d;
assign v8e5367 = StoB_REQ6_p & v8a6914 | !StoB_REQ6_p & !v86ce9d;
assign v8562d4 = BtoR_REQ0_p & v865b8f | !BtoR_REQ0_p & v85f2b2;
assign v85f3dd = jx2_p & v8569a8 | !jx2_p & !v8e3ee9;
assign v8e1c59 = ENQ_p & v844fbf | !ENQ_p & !v865764;
assign v856819 = RtoB_ACK0_p & v8567f9 | !RtoB_ACK0_p & v8af209;
assign v8e3bf3 = StoB_REQ0_p & v8e5033 | !StoB_REQ0_p & v856594;
assign v8e1abe = StoB_REQ2_p & v85b540 | !StoB_REQ2_p & v8563c0;
assign v8e40df = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5786;
assign v8af4a4 = BtoS_ACK7_p & v85737f | !BtoS_ACK7_p & v85cd17;
assign v85d757 = BtoS_ACK0_p & v8e5a1c | !BtoS_ACK0_p & v8e5486;
assign v856ff6 = ENQ_p & v8e3a26 | !ENQ_p & v8cc8b1;
assign v8b54ed = EMPTY_p & v8e5881 | !EMPTY_p & v8b5665;
assign v85d539 = jx2_p & v856b6d | !jx2_p & v85b5d9;
assign v8e5244 = BtoS_ACK3_p & v85dbdd | !BtoS_ACK3_p & v8b57b2;
assign v85daa5 = jx0_p & v8b5758 | !jx0_p & v8e5a3b;
assign v8e17e6 = StoB_REQ2_p & v867a58 | !StoB_REQ2_p & v8e3d20;
assign v8b42e8 = BtoS_ACK0_p & v86972a | !BtoS_ACK0_p & v85ba2c;
assign v8e5b63 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8e3bb9;
assign v85da56 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8b586a;
assign v8e4189 = BtoS_ACK7_p & v8e4764 | !BtoS_ACK7_p & v856ea9;
assign v8e58ad = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8b5687;
assign v8e4c47 = jx0_p & v844f9f | !jx0_p & !v844f9d;
assign v85dbbe = BtoS_ACK0_p & v8568a1 | !BtoS_ACK0_p & v85fc19;
assign v8a5b8c = BtoS_ACK6_p & v8b5840 | !BtoS_ACK6_p & v8e38a9;
assign v8a5bca = BtoS_ACK6_p & v8e42fd | !BtoS_ACK6_p & v8e54e0;
assign v8e58b1 = BtoS_ACK6_p & v8b583b | !BtoS_ACK6_p & v8b54d5;
assign v8e1b83 = StoB_REQ1_p & v8e214e | !StoB_REQ1_p & v856481;
assign v8dc607 = BtoS_ACK0_p & v8e4831 | !BtoS_ACK0_p & v8e23b9;
assign v8e19c2 = jx1_p & v8e509c | !jx1_p & v8e4051;
assign v8e590d = BtoS_ACK6_p & v860037 | !BtoS_ACK6_p & v856c3c;
assign v8cf0f4 = jx0_p & v844f91 | !jx0_p & v8e4831;
assign v8b5596 = StoB_REQ0_p & v8e42b6 | !StoB_REQ0_p & v889f95;
assign v8b587b = jx1_p & v8a5b1b | !jx1_p & v85a8af;
assign v8e1de6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5799;
assign v8e3aa7 = StoB_REQ8_p & v85e8b5 | !StoB_REQ8_p & v85fbec;
assign v881b42 = EMPTY_p & v8e5ba4 | !EMPTY_p & v856f27;
assign v8cc8c9 = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & v8af44d;
assign v8e5a5e = jx2_p & v8e3de0 | !jx2_p & v85dfab;
assign v8e1e0e = jx1_p & v8b56ee | !jx1_p & v8cce52;
assign v8691fd = BtoS_ACK0_p & v85d90a | !BtoS_ACK0_p & v8b35f2;
assign v8b58ba = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af29a;
assign v8be101 = jx2_p & v85dcf5 | !jx2_p & !v85b036;
assign v8e5b0f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v89920d;
assign v8565b3 = BtoS_ACK6_p & v85e281 | !BtoS_ACK6_p & v85d6a8;
assign v8b562d = stateG12_p & v8e54de | !stateG12_p & !v865764;
assign v8e57de = EMPTY_p & v85ca37 | !EMPTY_p & v8e4497;
assign v856cb3 = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & !v8e3b87;
assign v8e4523 = jx1_p & v8b56ee | !jx1_p & v85ad39;
assign v8b5895 = jx1_p & v8e45c6 | !jx1_p & v85ea86;
assign v8e1bf5 = StoB_REQ0_p & v8e22c3 | !StoB_REQ0_p & v8b55e8;
assign v8563b7 = jx1_p & v85d8ba | !jx1_p & !v8e47f9;
assign v8563f1 = jx1_p & v8e5aa3 | !jx1_p & v844f91;
assign v8e39e6 = jx1_p & v85db8a | !jx1_p & !v8af0dc;
assign v889264 = StoB_REQ6_p & v85e237 | !StoB_REQ6_p & v8e3c2f;
assign v85a4f0 = DEQ_p & v84510d | !DEQ_p & v86290f;
assign v85dfb7 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844fa3;
assign v8af34b = BtoS_ACK8_p & v8dc5ff | !BtoS_ACK8_p & !v8e1f73;
assign v8cce79 = jx0_p & v8e4637 | !jx0_p & !v8b5893;
assign v8b5806 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85de64;
assign v8e4605 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e1e8c;
assign v8e54fe = jx1_p & v8e5810 | !jx1_p & !v8e1701;
assign v8e4051 = StoB_REQ6_p & v85d7bd | !StoB_REQ6_p & v8cce20;
assign v8569c7 = jx2_p & v8b550b | !jx2_p & v8e1acc;
assign v8b56e0 = StoB_REQ8_p & v8e432e | !StoB_REQ8_p & v8e3e66;
assign v84530d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8562ad;
assign v889f6e = jx1_p & v85f1ac | !jx1_p & !v844f91;
assign v85b3fb = BtoS_ACK1_p & v8b5600 | !BtoS_ACK1_p & v889e03;
assign v8b572e = StoB_REQ8_p & v8e1abd | !StoB_REQ8_p & !v8b588e;
assign v8e593f = EMPTY_p & v8e1985 | !EMPTY_p & v8dc5e7;
assign v8e5c0a = StoB_REQ0_p & v8e39cc | !StoB_REQ0_p & v8e5a09;
assign v8b5683 = BtoS_ACK0_p & v89920d | !BtoS_ACK0_p & v8b580f;
assign v880bc4 = jx2_p & v8e5a3e | !jx2_p & v856386;
assign v8b5838 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8892b3;
assign v8b5839 = StoB_REQ0_p & v8e4a22 | !StoB_REQ0_p & v8b5625;
assign v8b564d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8575ef;
assign v8e57a1 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844fb7;
assign v85cc48 = BtoS_ACK6_p & v8e4cb9 | !BtoS_ACK6_p & v85ba35;
assign v85d433 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85d794;
assign v8b5768 = jx1_p & v8a87cd | !jx1_p & v85e653;
assign v8e16e1 = EMPTY_p & v85a893 | !EMPTY_p & v8e503e;
assign v8be11a = jx2_p & v8e4ca6 | !jx2_p & v8cc8fb;
assign v8e568f = BtoR_REQ1_p & v8b54c6 | !BtoR_REQ1_p & v85b57e;
assign v884bb3 = StoB_REQ6_p & v8e4050 | !StoB_REQ6_p & v85ac27;
assign v856ef1 = jx1_p & v85d8ba | !jx1_p & !v85e2b5;
assign v856c6d = BtoS_ACK0_p & v8b585f | !BtoS_ACK0_p & v883e72;
assign v8b54cb = DEQ_p & v889f9b | !DEQ_p & v8569df;
assign v85e152 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e4976;
assign v85e4fc = jx0_p & v8b5698 | !jx0_p & v8b570f;
assign v85fa37 = jx1_p & v856a23 | !jx1_p & !v844f91;
assign v8845b3 = jx2_p & v8b5601 | !jx2_p & v881ad8;
assign v8451cf = BtoS_ACK1_p & v8e4a1f | !BtoS_ACK1_p & v85a1ee;
assign v8b5666 = BtoS_ACK6_p & v8565a3 | !BtoS_ACK6_p & v8e1c72;
assign v85a4ae = StoB_REQ6_p & v8e198d | !StoB_REQ6_p & v844f91;
assign v856ecb = StoB_REQ6_p & v8e462b | !StoB_REQ6_p & v8e1f66;
assign v856b4f = jx0_p & v8b587e | !jx0_p & v8e4163;
assign v8e58b7 = BtoS_ACK7_p & v8a87fd | !BtoS_ACK7_p & v8e181b;
assign v8e591f = ENQ_p & v8af34b | !ENQ_p & v8e1ec6;
assign v8a5cb5 = jx2_p & v8e42df | !jx2_p & !v8b5895;
assign v8b553f = jx0_p & v8e4d94 | !jx0_p & !v8e5a00;
assign v8e462b = BtoS_ACK0_p & v8e4c47 | !BtoS_ACK0_p & v889fde;
assign v8e58a7 = BtoS_ACK6_p & v85f64e | !BtoS_ACK6_p & v885465;
assign v8b559d = BtoS_ACK6_p & v8b584f | !BtoS_ACK6_p & v85b60a;
assign v8e4a1f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e3883;
assign v8e42fe = StoB_REQ0_p & v8e4c47 | !StoB_REQ0_p & v85d90a;
assign v8e38a9 = jx2_p & v85a863 | !jx2_p & v85e994;
assign v85f42f = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v844fa1;
assign v8e4f36 = jx2_p & v856eb9 | !jx2_p & v8b552b;
assign v8803e2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85727c;
assign v85ad1a = BtoS_ACK7_p & v8e176c | !BtoS_ACK7_p & v85f34e;
assign v8e3bb9 = StoB_REQ3_p & v8e5000 | !StoB_REQ3_p & !v844f91;
assign v8b566b = ENQ_p & v8572d0 | !ENQ_p & v8e109f;
assign v889f8a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b575b;
assign v85b390 = StoB_REQ6_p & v858ae4 | !StoB_REQ6_p & v8e4cc7;
assign v8e1c7f = EMPTY_p & v858981 | !EMPTY_p & v889244;
assign v8e38c8 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e463e;
assign v8e1a78 = StoB_REQ6_p & v85a8af | !StoB_REQ6_p & v8e548f;
assign v85737f = jx2_p & v8b5548 | !jx2_p & v844f91;
assign v8e3fa0 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8b569f;
assign v87f854 = StoB_REQ7_p & v8e5982 | !StoB_REQ7_p & v844f91;
assign v8e15b2 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e5a2c;
assign v85d7a7 = jx1_p & v85acf3 | !jx1_p & v8b5771;
assign v8b5586 = StoB_REQ0_p & v85b2bc | !StoB_REQ0_p & v844f91;
assign v85afc8 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v85b6c8;
assign v883ca3 = jx0_p & v844f9b | !jx0_p & !v844f91;
assign v8e3e0e = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8b5596;
assign v856b0d = BtoS_ACK7_p & v8e4235 | !BtoS_ACK7_p & v8b5897;
assign v85f953 = BtoS_ACK6_p & v8e5650 | !BtoS_ACK6_p & v8b5859;
assign v8b5554 = jx0_p & v8a87b4 | !jx0_p & v8e3e82;
assign v85b3a4 = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8e42b6;
assign v8b586a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f99;
assign v8b565e = BtoS_ACK8_p & v85e947 | !BtoS_ACK8_p & v85e0ba;
assign BtoS_ACK7_n = !v8cce8a;
assign v8dc593 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e3d20;
assign v8e58bd = ENQ_p & v8e2059 | !ENQ_p & !v844f91;
assign v845235 = RtoB_ACK0_p & v8e59af | !RtoB_ACK0_p & v8e5a54;
assign v85adad = jx1_p & v85dee1 | !jx1_p & !v85b3a4;
assign v89b6ce = BtoS_ACK0_p & v8e1664 | !BtoS_ACK0_p & v8e5a48;
assign v85e836 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e1a57;
assign v856bb4 = jx0_p & v8e5a3f | !jx0_p & !v85f2cd;
assign v8af1a3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e3979;
assign v8dc5e7 = DEQ_p & v8b57c8 | !DEQ_p & v860057;
assign v8bf437 = BtoS_ACK8_p & v85d914 | !BtoS_ACK8_p & v8a880e;
assign v85d805 = jx2_p & v8b57d5 | !jx2_p & v8b55bf;
assign v85cb96 = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & !v85ea88;
assign v885341 = StoB_REQ6_p & v85ffcd | !StoB_REQ6_p & v844f91;
assign v865772 = jx1_p & v8e5a23 | !jx1_p & v8e59df;
assign v85a1ee = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4fff;
assign BtoS_ACK0_n = !v8be173;
assign v8af226 = StoB_REQ1_p & v8a87b4 | !StoB_REQ1_p & v844f9f;
assign v8b5778 = BtoS_ACK0_p & v8af46d | !BtoS_ACK0_p & !v844f95;
assign v8b5831 = RtoB_ACK0_p & v8b556b | !RtoB_ACK0_p & !v844f91;
assign v8e4fad = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v881aaf;
assign v8e20a2 = StoB_REQ1_p & v8e214e | !StoB_REQ1_p & v85ffdf;
assign v8b57d5 = jx1_p & v844f91 | !jx1_p & v8b5786;
assign v85b9a9 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8e1e8c;
assign v8cce37 = jx2_p & v85761b | !jx2_p & v844f91;
assign v8e54de = ENQ_p & v844f91 | !ENQ_p & !v865764;
assign v8e1e31 = BtoS_ACK7_p & v8b54f2 | !BtoS_ACK7_p & v85f2aa;
assign v856594 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v85c632;
assign v8e5022 = jx0_p & v844f91 | !jx0_p & !v8af47b;
assign v85ad2e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8e38d9;
assign v85a23c = jx1_p & v8565a3 | !jx1_p & v8e40df;
assign v8e42c6 = StoB_REQ0_p & v85f2f8 | !StoB_REQ0_p & v8be123;
assign v8e3bdc = StoB_REQ8_p & v85dc95 | !StoB_REQ8_p & v8e4d72;
assign v8b57ec = jx1_p & v8b56f1 | !jx1_p & !v85a6d2;
assign v856a93 = jx1_p & v85fa41 | !jx1_p & !v85c73e;
assign v8e1841 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e17e8;
assign v8b56de = jx1_p & v8e59d4 | !jx1_p & v8e5a7e;
assign v85630a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v85ea88;
assign v85f27b = stateG12_p & v8b55ed | !stateG12_p & v844f91;
assign v8e408d = BtoS_ACK1_p & v8e52f8 | !BtoS_ACK1_p & v8e1bc6;
assign v856663 = jx1_p & v8e4514 | !jx1_p & v8e462b;
assign v8ca6f1 = BtoS_ACK6_p & v8cce3b | !BtoS_ACK6_p & v8b5789;
assign v8e1651 = BtoS_ACK8_p & v8e58d8 | !BtoS_ACK8_p & !v85d309;
assign v85df0b = StoB_REQ7_p & v8e1fe7 | !StoB_REQ7_p & v8e58d3;
assign v8b553b = jx1_p & v860551 | !jx1_p & v85dee5;
assign v8e50c2 = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v85dcb5;
assign v8e4f28 = StoB_REQ0_p & v8e38b0 | !StoB_REQ0_p & v8e4261;
assign v8572b6 = BtoS_ACK6_p & v8e4c29 | !BtoS_ACK6_p & v8a5c58;
assign v8e3f6f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b56f7;
assign v85db39 = jx0_p & v88c324 | !jx0_p & v8b56ce;
assign v8e4ac8 = StoB_REQ7_p & v85ffcd | !StoB_REQ7_p & v844f91;
assign v8e1f7f = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85ea88;
assign v8b5506 = BtoS_ACK8_p & v8e165a | !BtoS_ACK8_p & !v8e438d;
assign v8b5761 = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v87d771;
assign v8846fb = StoB_REQ8_p & v8dc639 | !StoB_REQ8_p & v8e572b;
assign v85dbf8 = BtoS_ACK6_p & v8e4235 | !BtoS_ACK6_p & v8e1df8;
assign v8e1ae8 = jx2_p & v8b56e4 | !jx2_p & v85d2e8;
assign v8e4472 = BtoS_ACK6_p & v856902 | !BtoS_ACK6_p & v8450b6;
assign v85e259 = StoB_REQ0_p & v85f2f8 | !StoB_REQ0_p & v85f59b;
assign v85da0f = jx1_p & v85e383 | !jx1_p & v8b58b7;
assign v85fabb = jx2_p & v8b55cc | !jx2_p & v86290d;
assign v8e56d9 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v85e340;
assign v8e5a4b = BtoS_ACK0_p & v8e5a10 | !BtoS_ACK0_p & v8b5707;
assign v8e16f6 = jx1_p & v85dbda | !jx1_p & v844f91;
assign v8b57a9 = ENQ_p & v8af46c | !ENQ_p & v844f91;
assign v881b59 = jx1_p & v85acf3 | !jx1_p & v85f2f8;
assign v85df78 = jx2_p & v85641f | !jx2_p & !v8b54db;
assign v8573cd = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844fb3;
assign v857553 = jx0_p & v8af44d | !jx0_p & v8e5155;
assign v8dc575 = EMPTY_p & v8635e4 | !EMPTY_p & v85cc98;
assign v85630d = jx2_p & v8569ce | !jx2_p & !v85cea0;
assign v85c6e4 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v86f85b;
assign v865810 = jx1_p & v8e5962 | !jx1_p & v88c2c4;
assign v8e5942 = jx2_p & v844f91 | !jx2_p & v8562b6;
assign v8b57ad = jx2_p & v844f91 | !jx2_p & !v8e21cf;
assign v8e58c4 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b55d4;
assign v8af389 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9d;
assign v8cc8fb = jx1_p & v8e422f | !jx1_p & v8567fa;
assign v8e45c6 = StoB_REQ6_p & v8e3dc6 | !StoB_REQ6_p & v8b577d;
assign v85b4ff = BtoS_ACK0_p & v8e4f71 | !BtoS_ACK0_p & v8b585d;
assign v85740b = DEQ_p & v8e15cb | !DEQ_p & v8b57a9;
assign v85f64e = jx2_p & v8e14db | !jx2_p & v8e4e45;
assign v8e4e45 = jx1_p & v85dbda | !jx1_p & !v8b57d0;
assign v8dc6c4 = RtoB_ACK1_p & v8af432 | !RtoB_ACK1_p & v85f5cc;
assign v85f79e = BtoS_ACK7_p & v889f6d | !BtoS_ACK7_p & !v8e4996;
assign v8b558c = BtoS_ACK8_p & v8e3f1b | !BtoS_ACK8_p & v8e597b;
assign v8e4b0e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b552d;
assign v8e1b23 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8af34f;
assign v85b4e6 = StoB_REQ2_p & v8e4224 | !StoB_REQ2_p & v8e589a;
assign v8600af = jx2_p & v84520f | !jx2_p & !v85ffcd;
assign v8e559d = BtoS_ACK0_p & v8e4831 | !BtoS_ACK0_p & v8e19a8;
assign v8e51f8 = BtoS_ACK6_p & v8be101 | !BtoS_ACK6_p & v85631f;
assign v8e4040 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v860007;
assign v8e4941 = RtoB_ACK0_p & v8e1f0d | !RtoB_ACK0_p & v85d7a6;
assign v85ad10 = BtoS_ACK1_p & v844fa0 | !BtoS_ACK1_p & v8e222b;
assign v85eac4 = StoB_REQ6_p & v8b5525 | !StoB_REQ6_p & !v8e54a9;
assign v85cbe8 = BtoS_ACK8_p & v8dc5ff | !BtoS_ACK8_p & v8e15a4;
assign v8e5a61 = BtoS_ACK7_p & v8a5c58 | !BtoS_ACK7_p & v85e1f5;
assign v85684d = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v880dfd;
assign v8caee0 = jx1_p & v844f91 | !jx1_p & v8e4dae;
assign v8b54d5 = jx2_p & v8e17c4 | !jx2_p & v85dd8c;
assign v8e4668 = BtoS_ACK8_p & v8e5833 | !BtoS_ACK8_p & v85dfb4;
assign v8b55f4 = jx1_p & v8e4a96 | !jx1_p & v8e530b;
assign v8e5a54 = BtoR_REQ1_p & v8dc6bf | !BtoR_REQ1_p & v86006a;
assign v8af18b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5557;
assign v8e58e0 = jx1_p & v85b238 | !jx1_p & !v85aeed;
assign v8b5557 = jx0_p & v844f91 | !jx0_p & v8e47d6;
assign v8e5a43 = BtoS_ACK6_p & v856fc9 | !BtoS_ACK6_p & v85db08;
assign v845033 = BtoS_ACK6_p & v8e4a85 | !BtoS_ACK6_p & v8b55e3;
assign v8e38f1 = BtoS_ACK0_p & v85a8af | !BtoS_ACK0_p & v8564b7;
assign v85abc1 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8e436c;
assign v8e1f7b = StoB_REQ0_p & v8e57b4 | !StoB_REQ0_p & v8e3c11;
assign v85c1d4 = StoB_REQ8_p & v8b5621 | !StoB_REQ8_p & v8e4255;
assign v8e21c5 = jx2_p & v844f91 | !jx2_p & v856354;
assign v8e158b = stateG7_1_p & v8e1a88 | !stateG7_1_p & v8e4f00;
assign v8e4a22 = jx0_p & v8b5856 | !jx0_p & v844f91;
assign v8e3977 = BtoS_ACK6_p & v8e2431 | !BtoS_ACK6_p & v8b560a;
assign v8565ea = DEQ_p & v8585f1 | !DEQ_p & v8cce0d;
assign v85e091 = jx1_p & v8e4514 | !jx1_p & v8e4c47;
assign v85ffdf = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8b5644;
assign v8e5903 = jx1_p & v85b238 | !jx1_p & !v844f91;
assign v85d441 = BtoS_ACK1_p & v8e52f8 | !BtoS_ACK1_p & v8e22de;
assign v8e209c = BtoS_ACK0_p & v8b55cb | !BtoS_ACK0_p & !v8e1902;
assign v8e198b = BtoR_REQ0_p & v8e57de | !BtoR_REQ0_p & v856fdd;
assign v85c47a = jx2_p & v85e3a8 | !jx2_p & v856b8f;
assign v85ba1d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8e49c8;
assign v85c416 = StoB_REQ2_p & v8af160 | !StoB_REQ2_p & !v844f91;
assign v85e2b5 = StoB_REQ7_p & v8e3eb2 | !StoB_REQ7_p & v844f91;
assign v85a0ae = BtoS_ACK7_p & v8e1b8d | !BtoS_ACK7_p & v85f953;
assign v8e40a9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v8e5a59 = jx1_p & v85f42f | !jx1_p & v8e3e4b;
assign v856765 = jx1_p & v8a87cd | !jx1_p & v844f91;
assign v8e4632 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85725c;
assign v8e10a4 = jx1_p & v8e59ee | !jx1_p & v8e59df;
assign v85c80b = jx2_p & v8b5549 | !jx2_p & v85dfab;
assign v8e587f = StoB_REQ0_p & v8e56dc | !StoB_REQ0_p & v8e3c73;
assign v8b567b = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e58d5;
assign v8a6d22 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85df25;
assign v856a03 = jx2_p & v8af402 | !jx2_p & v8b54f4;
assign v85df7f = StoB_REQ0_p & v8e39cc | !StoB_REQ0_p & v85f244;
assign v8a923a = BtoS_ACK6_p & v8be101 | !BtoS_ACK6_p & v8b5678;
assign v8626fe = jx0_p & v844f91 | !jx0_p & !v8dc552;
assign v8e1fa5 = jx2_p & v85b5c5 | !jx2_p & v8e3c23;
assign v8e1df8 = jx2_p & v8e1f2a | !jx2_p & v844f91;
assign v8b5517 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v85c9c5;
assign v8e472c = jx2_p & v8e5b65 | !jx2_p & v8e3d1a;
assign v8566db = jx2_p & v8b5784 | !jx2_p & !v85e5cf;
assign v8b57cc = jx1_p & v85d5b1 | !jx1_p & !v8e46ed;
assign v8860f1 = jx0_p & v8e3c39 | !jx0_p & v8cc8e8;
assign v856ea9 = BtoS_ACK6_p & v8af325 | !BtoS_ACK6_p & v856a38;
assign v8e5a7a = BtoS_ACK0_p & v8af190 | !BtoS_ACK0_p & v8564e9;
assign v8e4f0b = StoB_REQ8_p & v8cc8fa | !StoB_REQ8_p & v844f91;
assign v85dd89 = StoB_REQ0_p & v8e4eb5 | !StoB_REQ0_p & v889f3d;
assign v8b56ce = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e19f0;
assign v8b54c6 = EMPTY_p & v8e3b4c | !EMPTY_p & v8563b6;
assign v8af3cb = BtoS_ACK0_p & v8b5663 | !BtoS_ACK0_p & v8571d0;
assign v8e588f = DEQ_p & v8e4f2e | !DEQ_p & v8601d6;
assign v8b5883 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v8650b9;
assign v85cdaa = StoB_REQ8_p & v8b573e | !StoB_REQ8_p & v8e1d76;
assign v85e45f = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & !v8e55ca;
assign v8b5856 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85d671;
assign v8b586f = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v857578;
assign v8567ae = jx2_p & v85f230 | !jx2_p & v8e57ab;
assign v85a0f8 = BtoS_ACK1_p & v8e16ea | !BtoS_ACK1_p & v889ec1;
assign v8564bf = BtoS_ACK6_p & v8b56ae | !BtoS_ACK6_p & v8e1f36;
assign v861da7 = StoB_REQ6_p & v88c326 | !StoB_REQ6_p & v859fe9;
assign v882912 = jx0_p & v8b55cb | !jx0_p & v844f91;
assign v8b5829 = jx1_p & v8e5b11 | !jx1_p & !v8b5889;
assign v8dc5ad = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8e5032;
assign v8e52f2 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v8e59e6;
assign v8e1778 = EMPTY_p & v85b5f8 | !EMPTY_p & v8b5665;
assign v85a34c = ENQ_p & v85e45f | !ENQ_p & v85d340;
assign v8e1902 = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & v85e7ea;
assign v85ccfd = BtoS_ACK0_p & v8e3d0c | !BtoS_ACK0_p & v8e5816;
assign v8e595b = BtoS_ACK7_p & v8e4235 | !BtoS_ACK7_p & v85d34c;
assign v845069 = StoB_REQ8_p & v884d71 | !StoB_REQ8_p & v8e47e7;
assign v86f694 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v8b57ac;
assign v8b5860 = jx2_p & v85e66e | !jx2_p & v856f8d;
assign v8b5795 = StoB_REQ7_p & v8e3eb2 | !StoB_REQ7_p & v8af355;
assign v85659c = BtoS_ACK2_p & v8bf0c7 | !BtoS_ACK2_p & v8b55f8;
assign v85cda6 = BtoS_ACK0_p & v8e4831 | !BtoS_ACK0_p & v8e1de6;
assign v85db0d = BtoS_ACK1_p & v8e4632 | !BtoS_ACK1_p & v8e5a01;
assign v8451c3 = BtoS_ACK7_p & v844fa1 | !BtoS_ACK7_p & !v8991aa;
assign v8e5968 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9d;
assign v8e5a80 = jx0_p & v8a87d6 | !jx0_p & v8e3a0e;
assign v8e4c73 = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v8e10aa;
assign v85f4ff = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b56cd;
assign v8e22c7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5893;
assign v85b9a0 = jx1_p & v8e4e56 | !jx1_p & v844f91;
assign v8e3cb6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cf0f4;
assign v8e466e = StoB_REQ1_p & v86e4e7 | !StoB_REQ1_p & v8e52f8;
assign v8e3ff5 = BtoR_REQ0_p & v8b564c | !BtoR_REQ0_p & v88e277;
assign v8e4dae = BtoS_ACK0_p & v85a8af | !BtoS_ACK0_p & v8e3af6;
assign v8e58ed = BtoS_ACK6_p & v856386 | !BtoS_ACK6_p & v8e57d8;
assign v8e54cf = stateG12_p & v8e4805 | !stateG12_p & v85d79a;
assign v8e1084 = jx0_p & v85e7be | !jx0_p & v86f856;
assign v85b938 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v8e16ea;
assign v8e5a5f = ENQ_p & v8e4e6e | !ENQ_p & v88bc46;
assign v8e2395 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v856b48;
assign v85e4ac = jx1_p & v85dbef | !jx1_p & v844f91;
assign v8e2267 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e1b44;
assign v8ca185 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8a6914;
assign v8984b0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8572f8;
assign v8e2213 = StoB_REQ8_p & v8e4ea5 | !StoB_REQ8_p & v8e465f;
assign v8af44d = BtoS_ACK1_p & v85c632 | !BtoS_ACK1_p & !v85cdc8;
assign v85d598 = EMPTY_p & v8e205f | !EMPTY_p & v85e81e;
assign v8af209 = BtoR_REQ1_p & v85ae84 | !BtoR_REQ1_p & v85b5f3;
assign v8e39cc = jx0_p & v86baf9 | !jx0_p & !v844f91;
assign v8b54e8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e1ead;
assign v8cce39 = stateG7_1_p & v8e5a56 | !stateG7_1_p & v8e1d80;
assign v85df5a = BtoS_ACK0_p & v8dc594 | !BtoS_ACK0_p & v8e1084;
assign v8cce46 = StoB_REQ8_p & v8b5662 | !StoB_REQ8_p & v8be143;
assign v86290d = jx0_p & v844f91 | !jx0_p & !v844f91;
assign v85a88e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a5cb3;
assign v8e5b65 = jx1_p & v86cb45 | !jx1_p & v8e58f8;
assign v860902 = EMPTY_p & v85f48a | !EMPTY_p & v8e1eab;
assign v856404 = RtoB_ACK0_p & v8b55ec | !RtoB_ACK0_p & !v85bd3d;
assign v8b5525 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85699e;
assign v8568f6 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8e46da;
assign v8e451f = jx0_p & v8e4003 | !jx0_p & !v8ccdf7;
assign v85dc42 = RtoB_ACK0_p & v889f0f | !RtoB_ACK0_p & v85667b;
assign v8e5000 = StoB_REQ5_p & v844fb7 | !StoB_REQ5_p & v844f91;
assign v8e38c7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85daa5;
assign v86e38c = StoB_REQ6_p & v8af46d | !StoB_REQ6_p & v8b5778;
assign v85afc0 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b55bd;
assign v85b1c3 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e214e;
assign v85e282 = StoB_REQ0_p & v8e39cc | !StoB_REQ0_p & v85ada7;
assign v8e17b2 = StoB_REQ1_p & v86f9a1 | !StoB_REQ1_p & v85ea88;
assign v8572f8 = jx0_p & v8e4943 | !jx0_p & !v85ae38;
assign v85699e = jx0_p & v844f91 | !jx0_p & !v844f97;
assign v8a691d = BtoS_ACK0_p & v883ca3 | !BtoS_ACK0_p & v859fe4;
assign v8b35f2 = StoB_REQ0_p & v8e4791 | !StoB_REQ0_p & v8819a3;
assign v88924d = StoB_REQ6_p & v867aa7 | !StoB_REQ6_p & v8e5a2c;
assign v8e2429 = stateG12_p & v8e42f6 | !stateG12_p & v8e572e;
assign v8b54f2 = jx2_p & v85b9a0 | !jx2_p & !v8e238d;
assign v8e5996 = StoB_REQ1_p & v8b556f | !StoB_REQ1_p & v8e1eb9;
assign v8e1a57 = BtoS_ACK2_p & v8a5bcf | !BtoS_ACK2_p & v85fa63;
assign v8e45f5 = BtoS_ACK1_p & v8e4a1f | !BtoS_ACK1_p & v8dc5fb;
assign v856eb7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4943;
assign v85f839 = EMPTY_p & v85f2a6 | !EMPTY_p & v8e14ca;
assign v8be0f9 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8a6914;
assign v8e3d1a = jx1_p & v8b55c1 | !jx1_p & v85e103;
assign v85e618 = EMPTY_p & v85b6e3 | !EMPTY_p & v8e5625;
assign v8b586c = StoB_REQ8_p & v856466 | !StoB_REQ8_p & v856bc1;
assign v8b57ef = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v85aa47;
assign v85b036 = jx1_p & v85f5a7 | !jx1_p & v87f854;
assign v8b55bf = jx1_p & v8af23a | !jx1_p & v8e1d94;
assign v85b69f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85b863;
assign v8e1e8c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85ad35;
assign v8b55db = BtoS_ACK8_p & v8af4c2 | !BtoS_ACK8_p & v8b5801;
assign v85e383 = BtoS_ACK0_p & v85dbda | !BtoS_ACK0_p & v883566;
assign v8e4eb5 = jx0_p & v889f3d | !jx0_p & v844f91;
assign v85f230 = jx1_p & v8e59f6 | !jx1_p & !v8e3a9d;
assign v85db32 = jx1_p & v86290d | !jx1_p & v8e5bed;
assign v8b56e6 = jx0_p & v844f9b | !jx0_p & !v844f99;
assign v8e4b5f = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v85ddb7;
assign v856466 = BtoS_ACK7_p & v8e1a5a | !BtoS_ACK7_p & v89920a;
assign v8e460d = StoB_REQ6_p & v85649c | !StoB_REQ6_p & v8b57fb;
assign v8e55a8 = StoB_REQ7_p & v8e38f1 | !StoB_REQ7_p & v8b57c9;
assign v85e548 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85b6b7;
assign v8e4988 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v856f73;
assign v85724d = BtoS_ACK1_p & v8e1692 | !BtoS_ACK1_p & v8e4ebc;
assign v8450c0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86c57a;
assign v8e4b4e = StoB_REQ6_p & v85660c | !StoB_REQ6_p & v8e58a0;
assign v844fe7 = jx2_p & v8b35f0 | !jx2_p & v8e58fa;
assign v8e157d = BtoS_ACK0_p & v85f59b | !BtoS_ACK0_p & v8b54c7;
assign v8e527e = BtoS_ACK1_p & v8b5875 | !BtoS_ACK1_p & v86824f;
assign v8af15c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v856e07;
assign v865833 = jx2_p & v8e3df4 | !jx2_p & v85dfab;
assign v8e4185 = jx0_p & v899202 | !jx0_p & !v8dc5ec;
assign v85b54e = jx0_p & v8b556d | !jx0_p & !v85724d;
assign v85ba35 = jx2_p & v8cce04 | !jx2_p & v8e45e3;
assign v8e4c9d = jx0_p & v8b5893 | !jx0_p & !v844f91;
assign v845039 = BtoS_ACK8_p & v8567ae | !BtoS_ACK8_p & v8af493;
assign v85f5cc = RtoB_ACK0_p & v8af432 | !RtoB_ACK0_p & v8e16e1;
assign v8b55e3 = jx2_p & v8b570c | !jx2_p & v85dcd6;
assign v8e5a3f = BtoS_ACK1_p & v85e000 | !BtoS_ACK1_p & v85f386;
assign v85e565 = jx2_p & v863b23 | !jx2_p & v85dfab;
assign v8e4b68 = jx0_p & v8b587e | !jx0_p & v8e5928;
assign v8b5648 = StoB_REQ8_p & v8e5887 | !StoB_REQ8_p & v85de73;
assign v8e3c2f = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8b557e;
assign v8b5600 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8bf0c7;
assign v8b5577 = jx2_p & v8e4337 | !jx2_p & v845146;
assign v8b55f0 = EMPTY_p & v8af3db | !EMPTY_p & v8e522a;
assign v8e41df = StoB_REQ6_p & v85b2e6 | !StoB_REQ6_p & v8e3c3e;
assign v865802 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e53b1;
assign v85f43b = jx1_p & v8b58b2 | !jx1_p & v8e5930;
assign v8a54f3 = jx0_p & v88bcd0 | !jx0_p & !v86f9a1;
assign v85ba47 = BtoS_ACK7_p & v8e3bf7 | !BtoS_ACK7_p & v8b5731;
assign v8e114b = BtoS_ACK8_p & v8e5a22 | !BtoS_ACK8_p & v85e272;
assign v85b57e = BtoR_REQ0_p & v8e3e83 | !BtoR_REQ0_p & v8b54c6;
assign v85d7bd = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86c74d;
assign v8af0dd = BtoS_ACK8_p & v8e5833 | !BtoS_ACK8_p & v85643a;
assign v8e4e99 = jx1_p & v8b5749 | !jx1_p & v844f91;
assign v8e5887 = BtoS_ACK7_p & v8e1a5a | !BtoS_ACK7_p & v8e57f0;
assign v8b5549 = jx1_p & v8a87cd | !jx1_p & v8452cd;
assign v85e18a = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85de34;
assign v8af46d = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v844f91;
assign v85d8ad = ENQ_p & v8b5607 | !ENQ_p & v8e4ba8;
assign v8e1eab = DEQ_p & v8e41db | !DEQ_p & v85d8ad;
assign v856803 = BtoS_ACK6_p & v8af325 | !BtoS_ACK6_p & v85f5e7;
assign v85dd7f = BtoS_ACK8_p & v8e1a8c | !BtoS_ACK8_p & !v8e4f99;
assign v8e212d = jx2_p & v8b56de | !jx2_p & v8e4a6c;
assign v85710e = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v881aaf;
assign v85e0c2 = ENQ_p & v8e4e6e | !ENQ_p & v85737f;
assign v8b56c3 = BtoS_ACK0_p & v85aa18 | !BtoS_ACK0_p & v8e53c7;
assign v84507b = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v85d8f4;
assign v8566fb = BtoS_ACK6_p & v8e4f37 | !BtoS_ACK6_p & v86583e;
assign v88c2d2 = StoB_REQ5_n & v844f91 | !StoB_REQ5_n & !v85ea8d;
assign v8b585a = BtoS_ACK6_p & v8e1956 | !BtoS_ACK6_p & v844fe7;
assign v8be0f6 = jx1_p & v8a54e5 | !jx1_p & !v8b5786;
assign v85f50b = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8e4800;
assign v8e2399 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8af160;
assign v88bcc8 = BtoS_ACK7_p & v85737f | !BtoS_ACK7_p & v8b5762;
assign v8e59b7 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & !v8e4391;
assign v8e53be = StoB_REQ6_p & v8dc65c | !StoB_REQ6_p & v8e55d6;
assign v8cb249 = jx1_p & v8e59be | !jx1_p & !v85fc4d;
assign v8b5857 = BtoS_ACK1_p & v8b5875 | !BtoS_ACK1_p & v8565ce;
assign v8e4d59 = BtoS_ACK8_p & v8e5a22 | !BtoS_ACK8_p & !v8e21c8;
assign v8dc67d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v899202;
assign v8b57f3 = BtoS_ACK6_p & v8b587a | !BtoS_ACK6_p & v8450b6;
assign v8571d0 = StoB_REQ0_p & v8e56dc | !StoB_REQ0_p & v85fc5a;
assign v85e887 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e54a4;
assign v8e53de = BtoR_REQ0_p & v867398 | !BtoR_REQ0_p & v8b5611;
assign v8984a8 = jx0_p & v85dd8e | !jx0_p & !v86d1ff;
assign v8af176 = BtoS_ACK0_p & v8af243 | !BtoS_ACK0_p & v85b739;
assign v88c2c2 = BtoR_REQ1_p & v856275 | !BtoR_REQ1_p & v8568a8;
assign v84520f = jx1_p & v8e59d1 | !jx1_p & v88c2c4;
assign v8e4b49 = RtoB_ACK1_p & v8e568f | !RtoB_ACK1_p & v8af3e3;
assign v8e4662 = BtoS_ACK0_p & v8e3cf8 | !BtoS_ACK0_p & v8e3c27;
assign v8a5bb4 = BtoS_ACK0_p & v8af0d0 | !BtoS_ACK0_p & v8cc8c9;
assign v85bdbc = jx2_p & v8e1ad8 | !jx2_p & !v8cb249;
assign v8e222b = BtoS_ACK2_p & v844fa0 | !BtoS_ACK2_p & v8e20fa;
assign v85dee1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v86290d;
assign v8a5bfd = BtoS_ACK0_p & v8af418 | !BtoS_ACK0_p & v8b553f;
assign v8e190d = StoB_REQ0_p & v8e39cc | !StoB_REQ0_p & v8b54ea;
assign v85f170 = stateG12_p & v8b566d | !stateG12_p & !v8e38c8;
assign v85e947 = jx2_p & v844f91 | !jx2_p & v8e591a;
assign v8e2373 = BtoR_REQ1_p & v8564ad | !BtoR_REQ1_p & v8e3dac;
assign v8e1695 = ENQ_p & v8585db | !ENQ_p & v844f91;
assign v873e9c = jx1_p & v85d3e9 | !jx1_p & v8e2267;
assign v85d45f = BtoS_ACK1_p & v8a87b4 | !BtoS_ACK1_p & v8e4a8a;
assign v8e5625 = DEQ_p & v8b55d7 | !DEQ_p & v8569df;
assign v8b55ed = ENQ_p & v8e4e6e | !ENQ_p & v844f91;
assign v8562b8 = BtoS_ACK0_p & v8b57d0 | !BtoS_ACK0_p & v8e239b;
assign v8e1c5f = BtoS_ACK1_p & v8a5b4f | !BtoS_ACK1_p & v8e44b5;
assign v8e3b4c = ENQ_p & v8af34b | !ENQ_p & v8b54c5;
assign v8af147 = BtoS_ACK0_p & v85a8af | !BtoS_ACK0_p & v8b57de;
assign v85c47d = StoB_REQ8_p & v8e1b90 | !StoB_REQ8_p & !v85722b;
assign v8e1ffd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85a4ae;
assign v85b5d9 = jx1_p & v85dbef | !jx1_p & !v8e239b;
assign v8b579f = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8e5952;
assign v8b54d1 = jx0_p & v8e5a69 | !jx0_p & !v8b563f;
assign v862c12 = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & v85688c;
assign v8e1bb4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8e239b;
assign v85da38 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85eac4;
assign v8e53c7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4b68;
assign v8e5a2a = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8e4a06;
assign v85faba = jx2_p & v8e5054 | !jx2_p & v85a0da;
assign v8e3c23 = jx1_p & v85c3e3 | !jx1_p & !v8b5808;
assign v8992c3 = jx3_p & v8e39e1 | !jx3_p & !v8e4b49;
assign v85d6ea = StoB_REQ7_p & v85dee5 | !StoB_REQ7_p & v844f91;
assign v8e4e2c = jx0_p & v85a51c | !jx0_p & v8e5a02;
assign v8e58ce = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8e2035;
assign v85c632 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e519b;
assign v8e5611 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e1678;
assign v84520b = jx0_p & v844f9b | !jx0_p & !v8840fd;
assign v8e593d = BtoS_ACK0_p & v85f6bc | !BtoS_ACK0_p & v8e3b5f;
assign v85c718 = jx0_p & v85b3fb | !jx0_p & v85dd75;
assign v8b56d1 = RtoB_ACK0_p & v85d8ae | !RtoB_ACK0_p & v85d750;
assign v845136 = jx1_p & v8e5678 | !jx1_p & !v8b5889;
assign v8b55a1 = BtoS_ACK0_p & v85aa18 | !BtoS_ACK0_p & v8e5979;
assign v8b576c = StoB_REQ7_p & v85b5f6 | !StoB_REQ7_p & v8e5b11;
assign v8b584f = jx2_p & v85e905 | !jx2_p & !v844f91;
assign v85f59b = jx0_p & v8e5a51 | !jx0_p & v85ccf0;
assign v8be0ea = jx1_p & v8b5679 | !jx1_p & !v8e400a;
assign v8e407e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v85bbb6;
assign v8e58b6 = jx1_p & v844f91 | !jx1_p & v8af271;
assign v85c6f5 = jx0_p & v856594 | !jx0_p & !v844f91;
assign v8b583c = jx2_p & v856358 | !jx2_p & v8b552b;
assign v8b5798 = ENQ_p & v8562d0 | !ENQ_p & !v85f9b8;
assign v8b587e = BtoS_ACK1_p & v8a87b4 | !BtoS_ACK1_p & v8e193b;
assign v8b55cc = jx1_p & v85b380 | !jx1_p & v86290d;
assign v8e1d78 = BtoS_ACK7_p & v8e5a3c | !BtoS_ACK7_p & v8b5701;
assign v856dc8 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8e5350;
assign v8e579b = EMPTY_p & v8e5a82 | !EMPTY_p & v8dc55f;
assign v8e4a14 = jx1_p & v8e3916 | !jx1_p & v844f91;
assign v8e205f = ENQ_p & v8e3f4c | !ENQ_p & !v86290d;
assign v8b570e = StoB_REQ7_p & v85d382 | !StoB_REQ7_p & v8e1b00;
assign v8e5816 = StoB_REQ0_p & v8e47f2 | !StoB_REQ0_p & v8e4e75;
assign v8e4599 = BtoS_ACK6_p & v8e3bf7 | !BtoS_ACK6_p & v85e8f4;
assign v85bbd9 = ENQ_p & v85ba14 | !ENQ_p & v8b5578;
assign v8e5aa0 = StoB_REQ1_p & v85d671 | !StoB_REQ1_p & v8be124;
assign v8e45fa = BtoS_ACK0_p & v85f6bc | !BtoS_ACK0_p & v85c6e4;
assign v85e68a = ENQ_p & v8e4d59 | !ENQ_p & v8b54c5;
assign v85dfad = jx0_p & v8b5698 | !jx0_p & v85ba2f;
assign v8b56fe = StoB_REQ6_p & v8e1199 | !StoB_REQ6_p & v8be142;
assign v8e4792 = jx2_p & v85aef4 | !jx2_p & v8e591a;
assign v8e148a = jx0_p & v844f91 | !jx0_p & !v8af44d;
assign v8b55c3 = jx1_p & v8e4514 | !jx1_p & v88c38a;
assign v8b56ad = BtoR_REQ1_p & v85f81e | !BtoR_REQ1_p & v856901;
assign v8b57a0 = jx1_p & v8e59be | !jx1_p & !v844f91;
assign v8e43f1 = BtoS_ACK1_p & v8a5b4f | !BtoS_ACK1_p & v85eb45;
assign v8e3dac = EMPTY_p & v8e5ad2 | !EMPTY_p & v856bd4;
assign v8e492c = BtoR_REQ1_p & v8dc575 | !BtoR_REQ1_p & v8b584e;
assign v856b41 = BtoS_ACK6_p & v8af11e | !BtoS_ACK6_p & v8e212d;
assign v85f2ba = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & v85fa3e;
assign v8e1bda = ENQ_p & v85e3a6 | !ENQ_p & v8e3d4a;
assign v88c2c4 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85e259;
assign v8e53ec = jx1_p & v8b58aa | !jx1_p & !v8b54e1;
assign v8cc8c3 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v85dfb7;
assign v8e14e0 = BtoS_ACK6_p & v8cce3b | !BtoS_ACK6_p & v8e424e;
assign v8e2303 = StoB_REQ6_p & v8e520c | !StoB_REQ6_p & v8b56af;
assign v8b56af = BtoS_ACK0_p & v856594 | !BtoS_ACK0_p & !v8cc8c9;
assign v85a277 = BtoS_ACK8_p & v8e3ed3 | !BtoS_ACK8_p & v8cce46;
assign v8b557d = BtoR_REQ1_p & v8b5611 | !BtoR_REQ1_p & v8e53de;
assign v85e652 = BtoS_ACK0_p & v8e3eb2 | !BtoS_ACK0_p & v8b562a;
assign v85b073 = StoB_REQ7_p & v8e4217 | !StoB_REQ7_p & v8e5678;
assign v8b5563 = EMPTY_p & v8b5668 | !EMPTY_p & v8b54f0;
assign v8b5558 = EMPTY_p & v8e49eb | !EMPTY_p & v8e5aa8;
assign v8b56eb = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v85e5cf;
assign v85b6e3 = ENQ_p & v85ba14 | !ENQ_p & v88bc4c;
assign v8e5810 = StoB_REQ6_p & v8e3a2f | !StoB_REQ6_p & v8e5989;
assign v8e5b7d = jx2_p & v844f91 | !jx2_p & v8564ef;
assign v8e4394 = StoB_REQ8_p & v85f79e | !StoB_REQ8_p & !v844f91;
assign v85d2c4 = stateG12_p & v8573c8 | !stateG12_p & v8e55e7;
assign v8b588c = BtoS_ACK0_p & v85aa21 | !BtoS_ACK0_p & v8e3e3a;
assign v85cbea = jx1_p & v856a23 | !jx1_p & !v8e552e;
assign v8e59f7 = jx1_p & v8e416f | !jx1_p & v8b572d;
assign v8e1d99 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v867a58;
assign v8b56d3 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8b553c;
assign v8e2451 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86f9a1;
assign v8e3bee = BtoS_ACK8_p & v8b55a6 | !BtoS_ACK8_p & v8b572e;
assign v8e5956 = jx2_p & v84535e | !jx2_p & v8b55bf;
assign v8af355 = StoB_REQ6_p & v85d7bd | !StoB_REQ6_p & v8e4a68;
assign v8b556b = EMPTY_p & v8e1651 | !EMPTY_p & v856669;
assign v8e5607 = BtoS_ACK8_p & v8b5577 | !BtoS_ACK8_p & !v8b5681;
assign v85a5e3 = jx1_p & v8e4bc9 | !jx1_p & v844f91;
assign v8e4f99 = StoB_REQ8_p & v85a880 | !StoB_REQ8_p & v84518e;
assign v8e58dd = EMPTY_p & v8e1985 | !EMPTY_p & v8dc55f;
assign v8b5662 = BtoS_ACK7_p & v85b60a | !BtoS_ACK7_p & v8b559d;
assign v85e8f4 = jx2_p & v844f91 | !jx2_p & !v889f6e;
assign v85ffcd = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4831;
assign v8e3ffc = BtoS_ACK8_p & v85d53f | !BtoS_ACK8_p & v8e45c9;
assign v8e4c7f = jx0_p & v85a51c | !jx0_p & v856809;
assign v8e51e4 = jx0_p & v8b57e9 | !jx0_p & !v889ec0;
assign v8af4c2 = jx2_p & v85c9fb | !jx2_p & v8e591a;
assign v8e58ac = jx1_p & v8af186 | !jx1_p & v88c2c4;
assign v8e59aa = jx1_p & v8e5957 | !jx1_p & v85a8af;
assign v85e1f5 = BtoS_ACK6_p & v899224 | !BtoS_ACK6_p & v8a5c58;
assign v85b5f6 = StoB_REQ0_p & v8dc594 | !StoB_REQ0_p & v865820;
assign v8e5588 = jx1_p & v8e587b | !jx1_p & v8e4dae;
assign v8e16f2 = EMPTY_p & v8e58bd | !EMPTY_p & !v8b5728;
assign v856b75 = StoB_REQ7_p & v85a8af | !StoB_REQ7_p & v88c36f;
assign v8e52b0 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v844f91;
assign v85b421 = jx1_p & v8e501b | !jx1_p & v85758c;
assign v85c433 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8e3a0e;
assign v8b58ae = StoB_REQ2_p & v8e3bef | !StoB_REQ2_p & v85f697;
assign v85e1fe = StoB_REQ8_p & v8b5621 | !StoB_REQ8_p & v8e4071;
assign v845386 = StoB_REQ8_p & v856b0d | !StoB_REQ8_p & v8b5712;
assign v8e4191 = jx2_p & v8e4337 | !jx2_p & v856801;
assign v8b5693 = jx0_p & v8e4943 | !jx0_p & v85b5fb;
assign v8e57dd = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v8e59b4;
assign v8e436b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v859fe9;
assign v8e1bf6 = BtoS_ACK0_p & v8e5033 | !BtoS_ACK0_p & v8b56e1;
assign v8a87cd = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v844f91;
assign v8672d0 = jx3_p & v8b5891 | !jx3_p & v85db5c;
assign v8e59e4 = StoB_REQ6_p & v8e5960 | !StoB_REQ6_p & v880b12;
assign v87c63e = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8e4229;
assign v85f5a7 = StoB_REQ7_p & v8b5812 | !StoB_REQ7_p & v844f91;
assign v8af4aa = jx2_p & v8e1b05 | !jx2_p & v8b58bb;
assign v845027 = ENQ_p & v8af46c | !ENQ_p & v856353;
assign v8991c9 = jx0_p & v86baf9 | !jx0_p & !v8e4d0c;
assign v8e569c = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v8e5000;
assign v8e3eb5 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8b5704;
assign v8672b3 = jx0_p & v844f91 | !jx0_p & !v8e5155;
assign v8e162b = BtoS_ACK7_p & v8e594d | !BtoS_ACK7_p & v8a554f;
assign v8e1bf9 = jx1_p & v85ccdf | !jx1_p & v8b5538;
assign v882bc3 = jx2_p & v85cbea | !jx2_p & v8e58aa;
assign v86d019 = StoB_REQ0_p & v85ccc2 | !StoB_REQ0_p & v844f91;
assign v85c7da = BtoS_ACK0_p & v85699e | !BtoS_ACK0_p & v85b739;
assign v8e1be0 = BtoS_ACK8_p & v8b578a | !BtoS_ACK8_p & v8af102;
assign v8e240e = stateG12_p & v8e3cfe | !stateG12_p & v844f91;
assign v8e4b93 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v85dd9f;
assign v85d3d0 = jx2_p & v8b5569 | !jx2_p & v86290f;
assign v8b55ea = jx2_p & v85f8fd | !jx2_p & v8e41c1;
assign v8e1598 = StoB_REQ7_p & v85a8af | !StoB_REQ7_p & v8e1ea1;
assign v8e4fff = BtoS_ACK2_p & v8e3883 | !BtoS_ACK2_p & v8650c5;
assign v856cd5 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v899550;
assign v899219 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e243e;
assign v8dc58b = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v8e1cc4 = StoB_REQ6_p & v85d382 | !StoB_REQ6_p & v85ba99;
assign v8cce0a = BtoR_REQ0_p & v856dbe | !BtoR_REQ0_p & !v8e2239;
assign v85cb8e = jx1_p & v8e4574 | !jx1_p & v844f91;
assign v8e41ae = jx1_p & v8e1c72 | !jx1_p & v8e4c6e;
assign v86824f = BtoS_ACK2_p & v8b5875 | !BtoS_ACK2_p & !v85aa15;
assign v8af37d = BtoS_ACK6_p & v856fc9 | !BtoS_ACK6_p & v8e21d3;
assign v84507d = jx2_p & v85dd3e | !jx2_p & v8e3e49;
assign v85ccb4 = BtoS_ACK6_p & v85dd64 | !BtoS_ACK6_p & v85e332;
assign v85d3f6 = jx1_p & v8e4d04 | !jx1_p & !v844f91;
assign v85dc21 = ENQ_p & v85ba14 | !ENQ_p & v856fdc;
assign v86650a = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v880b59;
assign v8e238b = StoB_REQ8_p & v8b5790 | !StoB_REQ8_p & v8e3b88;
assign v8e22c3 = jx0_p & v86e828 | !jx0_p & !v84518f;
assign v8b5658 = StoB_REQ6_p & v8e4e81 | !StoB_REQ6_p & v84513a;
assign v86ae81 = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v85d475;
assign v85727c = BtoS_ACK0_p & v8e4d7b | !BtoS_ACK0_p & v8e59a9;
assign v8572d0 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e4f5f;
assign v8e58d6 = jx0_p & v856594 | !jx0_p & v84507a;
assign v8b55ff = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e1be3;
assign v8e5b23 = BtoS_ACK7_p & v8e420a | !BtoS_ACK7_p & v85e8f2;
assign v85d2bd = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v857553;
assign v885465 = jx2_p & v8e5098 | !jx2_p & v8b567a;
assign v86c2d3 = ENQ_p & v8562d0 | !ENQ_p & !v861611;
assign v8e550e = jx0_p & v8b5722 | !jx0_p & v844f91;
assign v856b8b = DEQ_p & v8b55d7 | !DEQ_p & v85bbd9;
assign v8e1ad8 = jx1_p & v85c8f2 | !jx1_p & v85aea9;
assign v8e3bf7 = jx2_p & v8b5503 | !jx2_p & !v8b57a0;
assign v8565ce = BtoS_ACK2_p & v8b5875 | !BtoS_ACK2_p & !v8b56bd;
assign v8e58e8 = StoB_REQ7_p & v8a87f0 | !StoB_REQ7_p & v8e48a0;
assign v85f594 = BtoS_ACK6_p & v865833 | !BtoS_ACK6_p & v8e595d;
assign v85677f = StoB_REQ0_p & v8dc594 | !StoB_REQ0_p & v8a9208;
assign v8cce04 = jx1_p & v8565cc | !jx1_p & v844f91;
assign v8e4cf4 = EMPTY_p & v8b57a9 | !EMPTY_p & v88934d;
assign v8e1cd2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85da6c;
assign v85e80e = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e1b83;
assign v8e4d9f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e1e59;
assign v8b5686 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v857037;
assign v8e2229 = BtoS_ACK7_p & v858f70 | !BtoS_ACK7_p & v861ed7;
assign v8e19e8 = jx0_p & v88bcd0 | !jx0_p & !v85630a;
assign v88c3ad = jx3_p & v8dc6c4 | !jx3_p & v8b5670;
assign v8b57d8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e42dc;
assign v85a8af = jx0_p & v844f91 | !jx0_p & !v844f9d;
assign v85c593 = BtoS_ACK6_p & v8600af | !BtoS_ACK6_p & v85d6a8;
assign v85ddc7 = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v8b588f;
assign v8e59d3 = BtoS_ACK1_p & v8e4632 | !BtoS_ACK1_p & v85a88e;
assign v8b56f1 = StoB_REQ7_p & v8572f7 | !StoB_REQ7_p & v845079;
assign v85e4af = jx1_p & v8e564d | !jx1_p & !v85fc4d;
assign v8cdce6 = jx0_p & v844f9f | !jx0_p & !v8e5a84;
assign v8b5615 = jx2_p & v8e4b4d | !jx2_p & !v865836;
assign v8a87ae = StoB_REQ0_p & v85c6f5 | !StoB_REQ0_p & v8e58d6;
assign v85e0b5 = BtoS_ACK2_p & v8e16ea | !BtoS_ACK2_p & v85684d;
assign v8e587b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8892c0;
assign v8e55ec = jx2_p & v8cce2b | !jx2_p & v8e41ec;
assign v8984a5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8573cd;
assign v85fc4e = jx2_p & v8caee0 | !jx2_p & v844f91;
assign v8e1d73 = StoB_REQ7_p & v8e5982 | !StoB_REQ7_p & v85ffcd;
assign v8b573f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e592e;
assign v8e594d = jx2_p & v88c371 | !jx2_p & v8b54f4;
assign v8e55d6 = BtoS_ACK0_p & v85e0b0 | !BtoS_ACK0_p & v8e1f47;
assign v857271 = jx1_p & v85acf3 | !jx1_p & v8b5551;
assign v8e1d00 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8e3d20;
assign v8e541f = EMPTY_p & v8e20a4 | !EMPTY_p & v85cc98;
assign v8e1e0a = StoB_REQ0_p & v8e39c1 | !StoB_REQ0_p & v8b583e;
assign v85da55 = jx1_p & v86c2ed | !jx1_p & v8e1598;
assign v8e58a1 = BtoS_ACK7_p & v8b55c6 | !BtoS_ACK7_p & v8e50d1;
assign v8e5917 = jx0_p & v8e4637 | !jx0_p & v844f99;
assign v8a552d = DEQ_p & v8e5a21 | !DEQ_p & v8e1c59;
assign v8991fe = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af1a3;
assign v85d543 = BtoS_ACK8_p & v863508 | !BtoS_ACK8_p & v85f567;
assign v8e51f4 = jx0_p & v8e15a0 | !jx0_p & v8e527e;
assign v8e44d3 = jx2_p & v8e59f7 | !jx2_p & v86e0c8;
assign v85fa6e = StoB_REQ1_p & v856eba | !StoB_REQ1_p & v844f91;
assign v8e3ee9 = jx1_p & v856763 | !jx1_p & !v8b55ca;
assign v8b552d = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & v85630a;
assign v8e4254 = BtoS_ACK0_p & v89b438 | !BtoS_ACK0_p & v8e2035;
assign v857374 = jx2_p & v88c2da | !jx2_p & v8852fd;
assign v8e1d5c = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v85b2a9;
assign v85a0da = jx1_p & v8b5508 | !jx1_p & !v8e4589;
assign v8e23a9 = BtoS_ACK0_p & v86290d | !BtoS_ACK0_p & !v8e239b;
assign v8b572b = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8e451f;
assign v8e1bc6 = StoB_REQ1_p & v8b558d | !StoB_REQ1_p & v8e5c47;
assign v8e5920 = BtoS_ACK1_p & v8a5b4f | !BtoS_ACK1_p & v8bf293;
assign v8e4086 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v85b642;
assign v8b56a9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8e474f;
assign v8e463e = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v86290d;
assign v85f2b2 = ENQ_p & v8a3c77 | !ENQ_p & v844f91;
assign v85e653 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v883cf8;
assign v8b5727 = jx2_p & v8e41ae | !jx2_p & v856f8d;
assign v8e1a97 = BtoS_ACK8_p & v8b5577 | !BtoS_ACK8_p & !v8e18e6;
assign v85d73d = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v8e4153;
assign v8b5670 = RtoB_ACK1_p & v8e492c | !RtoB_ACK1_p & v8b56bb;
assign v8b58ab = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b5683;
assign v8e5a23 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5b0f;
assign v889270 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8e3d7b;
assign v8e2436 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dc617;
assign v889f3b = BtoS_ACK3_p & v8b5875 | !BtoS_ACK3_p & !v8b56bd;
assign v8e2470 = StoB_REQ7_p & v883ca3 | !StoB_REQ7_p & v8e564d;
assign v8e4f8b = jx0_p & v8b55d1 | !jx0_p & v844f91;
assign v8e5880 = DEQ_p & v8b54eb | !DEQ_p & v8b572c;
assign v8e4f3b = jx1_p & v8e59d4 | !jx1_p & v8e453e;
assign v8b589f = FULL_p & v8601d6 | !FULL_p & v8e1c59;
assign v8be173 = jx3_p & v85deeb | !jx3_p & v857423;
assign v85dba0 = StoB_REQ7_p & v8e5a7a | !StoB_REQ7_p & v844f91;
assign v8e50a2 = jx2_p & v85c639 | !jx2_p & v8e53c6;
assign v844fcb = DEQ_p & v844f91 | !DEQ_p & !v844f91;
assign v84523d = jx0_p & v8b5893 | !jx0_p & v844f91;
assign v8b5841 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8572c2;
assign v8e5364 = RtoB_ACK0_p & v899261 | !RtoB_ACK0_p & !v8e5909;
assign v8e3c75 = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & !v85b4e6;
assign v8e431c = BtoR_REQ1_p & v856261 | !BtoR_REQ1_p & !v8e4f78;
assign v889244 = DEQ_p & v85f170 | !DEQ_p & v8e2147;
assign v8e1f76 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85e694;
assign v8e1810 = jx0_p & v8e59b7 | !jx0_p & !v8b5893;
assign v8b562f = jx2_p & v8bf8d8 | !jx2_p & v8e41d0;
assign v8be123 = jx0_p & v8e5a51 | !jx0_p & v85c971;
assign v85b898 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v85660f;
assign v8af2e6 = BtoS_ACK0_p & v8568a1 | !BtoS_ACK0_p & v856895;
assign v85d309 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v85e08e;
assign v85b5db = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8e570a;
assign v8e4e15 = jx2_p & v85fa37 | !jx2_p & v86290f;
assign v8e45b5 = BtoS_ACK6_p & v8b57a8 | !BtoS_ACK6_p & v85fabb;
assign v85fc09 = StoB_REQ0_p & v85a153 | !StoB_REQ0_p & v8e239b;
assign v8e4e4e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8e22c7;
assign v85ffb2 = jx1_p & v844f91 | !jx1_p & !v85ca01;
assign v8e4b00 = StoB_REQ7_p & v86290d | !StoB_REQ7_p & v856255;
assign v8892b3 = jx0_p & v844f91 | !jx0_p & v8b5722;
assign v8b5745 = StoB_REQ7_p & v85b3a4 | !StoB_REQ7_p & v877314;
assign v8e5085 = BtoS_ACK0_p & v85d90a | !BtoS_ACK0_p & v8e4118;
assign v88c32b = StoB_REQ2_p & v8e4f80 | !StoB_REQ2_p & v8e5426;
assign v8e3c83 = jx2_p & v8e4267 | !jx2_p & v8e591a;
assign v8e23b9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85672e;
assign v8e44c8 = BtoS_ACK0_p & v8b557e | !BtoS_ACK0_p & v8b56d3;
assign v858981 = ENQ_p & v8b55a4 | !ENQ_p & !v8e38c8;
assign v8b574d = BtoS_ACK6_p & v8e2416 | !BtoS_ACK6_p & v8af12b;
assign v86582c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e5a66;
assign v8e19b0 = BtoS_ACK6_p & v8b583b | !BtoS_ACK6_p & v8b56cf;
assign v889ec2 = stateG7_1_p & v8e5698 | !stateG7_1_p & v845360;
assign v8b54c2 = BtoS_ACK0_p & v8892b3 | !BtoS_ACK0_p & v85dbf7;
assign v856ce2 = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v856656;
assign v85758c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e17b8;
assign v8b56ef = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8e3c9e;
assign v8b56e4 = jx1_p & v8b560a | !jx1_p & !v8e58ef;
assign v8e5a10 = jx0_p & v8e4c04 | !jx0_p & !v8e466e;
assign v8e2098 = jx2_p & v8af4c4 | !jx2_p & v8e4fe5;
assign v8e5b58 = jx1_p & v881baf | !jx1_p & v8e59df;
assign v899fe9 = DEQ_p & v85a600 | !DEQ_p & v86290d;
assign v8b5750 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8be15d;
assign v8e4636 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e5989;
assign v8e4832 = BtoS_ACK1_p & v8a87b4 | !BtoS_ACK1_p & v8b54c4;
assign v884d71 = BtoS_ACK7_p & v8b5672 | !BtoS_ACK7_p & !v8e502c;
assign v8e1f19 = jx0_p & v85ad10 | !jx0_p & v8e4db2;
assign v85ea99 = BtoS_ACK0_p & v8be123 | !BtoS_ACK0_p & v856eb5;
assign v8b55a4 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v844fa5;
assign v8b5625 = jx0_p & v8e55a3 | !jx0_p & v844f91;
assign v8e23b1 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8984a5;
assign v8e23ae = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8e4a22;
assign v85db8a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5838;
assign v8b5837 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v845379;
assign v8e49c8 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e4caf;
assign v8e20d0 = BtoS_ACK7_p & v8e4764 | !BtoS_ACK7_p & v8e4cae;
assign v8e56ca = StoB_REQ7_p & v85df5b | !StoB_REQ7_p & v85c7da;
assign v85f81e = EMPTY_p & v8b5682 | !EMPTY_p & v8e5a94;
assign v8e5692 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v880dfd;
assign v8e40eb = EMPTY_p & v85a600 | !EMPTY_p & v899fe9;
assign v85dd22 = BtoS_ACK0_p & v8b5663 | !BtoS_ACK0_p & v8e1f7b;
assign v8e4638 = BtoR_REQ0_p & v8b57bd | !BtoR_REQ0_p & v8e16f2;
assign v8e592e = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e5bd5;
assign v8b56ca = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85da8e;
assign v876a22 = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v85bdb6;
assign v8b578a = jx2_p & v8e4dbe | !jx2_p & v8e41d0;
assign v86bc13 = BtoS_ACK6_p & v85a008 | !BtoS_ACK6_p & v856406;
assign v8e1088 = BtoS_ACK6_p & v8e3bf7 | !BtoS_ACK6_p & v8e5b6d;
assign v8b5503 = jx1_p & v844f91 | !jx1_p & v85aea9;
assign v845047 = BtoS_ACK6_p & v85a10a | !BtoS_ACK6_p & v8e4e02;
assign v8b55bc = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v85e274;
assign v8e58c9 = StoB_REQ7_p & v8b57ff | !StoB_REQ7_p & v8e18bd;
assign v8e42df = jx1_p & v85c6ec | !jx1_p & !v88c36f;
assign v8e5891 = jx1_p & v8e5a7f | !jx1_p & v856b75;
assign v8b5765 = jx1_p & v8b5879 | !jx1_p & v8e40df;
assign v8e50d1 = BtoS_ACK6_p & v85630d | !BtoS_ACK6_p & v8a5c22;
assign v85aab4 = BtoS_ACK1_p & v8e5bb2 | !BtoS_ACK1_p & v85df40;
assign v86972a = jx0_p & v8b5600 | !jx0_p & v8e5bb2;
assign v884771 = BtoS_ACK6_p & v85a008 | !BtoS_ACK6_p & v856878;
assign v857056 = DEQ_p & v8e1dbf | !DEQ_p & v8564c4;
assign v863b40 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e5bd5;
assign v8e591a = jx1_p & v8e388e | !jx1_p & v844f91;
assign v8b551a = jx0_p & v8b5675 | !jx0_p & v85f2cd;
assign v845109 = BtoS_ACK6_p & v885308 | !BtoS_ACK6_p & v8e1ae8;
assign v88d6ad = StoB_REQ6_p & v85e5cf | !StoB_REQ6_p & v844f91;
assign v8893b1 = jx3_p & v85702d | !jx3_p & v85dcb6;
assign v8e58d9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8e595c;
assign v8b5896 = StoB_REQ7_p & v8e4050 | !StoB_REQ7_p & v8e1f7e;
assign v8b57c9 = StoB_REQ6_p & v8cf114 | !StoB_REQ6_p & v8e5a4b;
assign v85d701 = BtoS_ACK8_p & v8e4988 | !BtoS_ACK8_p & v8b55d8;
assign v88c36f = StoB_REQ6_p & v8e1701 | !StoB_REQ6_p & v85f53b;
assign BtoS_ACK4_n = !v8a887e;
assign v8e3a9d = StoB_REQ7_p & v8af418 | !StoB_REQ7_p & v889264;
assign v8e43dc = jx2_p & v8e5588 | !jx2_p & v844f91;
assign v85dd8e = BtoS_ACK1_p & v85e000 | !BtoS_ACK1_p & v867a71;
assign v8e55ca = BtoS_ACK7_p & v85deb5 | !BtoS_ACK7_p & !v8b5589;
assign v8e2147 = stateG12_p & v8b566d | !stateG12_p & !v8e3ab5;
assign BtoR_REQ1_n = !v883d05;
assign v8e3df4 = jx1_p & v85dee1 | !jx1_p & v8e4c47;
assign v8e57e7 = BtoS_ACK7_p & v85f448 | !BtoS_ACK7_p & v8b5656;
assign v85f194 = EMPTY_p & v8b582a | !EMPTY_p & v8b54ec;
assign v8e22d4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b5586;
assign v856314 = jx1_p & v889f8a | !jx1_p & v8e4dae;
assign v8e3f4c = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v86ed0b;
assign v8b5665 = DEQ_p & v8e5881 | !DEQ_p & v8e3fce;
assign v8e59d8 = jx2_p & v857271 | !jx2_p & v8e3b2b;
assign v8564ad = EMPTY_p & v8e5ad2 | !EMPTY_p & v8833ba;
assign v8563df = BtoS_ACK0_p & v8e5917 | !BtoS_ACK0_p & v8e409a;
assign v8e1aea = jx2_p & v85adad | !jx2_p & v8b567a;
assign v85de53 = StoB_REQ0_p & v8e5033 | !StoB_REQ0_p & v8b57d0;
assign BtoS_ACK2_n = !v889fea;
assign v85b04f = BtoS_ACK0_p & v8b56ce | !BtoS_ACK0_p & v8e5a48;
assign v856f79 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8e569c;
assign v881a3e = jx0_p & v844f9f | !jx0_p & !v8b5733;
assign v8b570f = BtoS_ACK1_p & v8e3d7b | !BtoS_ACK1_p & v8b579f;
assign v8e21cf = jx1_p & v8a691d | !jx1_p & !v844f91;
assign v8a5c84 = jx2_p & v845222 | !jx2_p & !v845146;
assign v857540 = StoB_REQ0_p & v8e4468 | !StoB_REQ0_p & v85de64;
assign v8e2431 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e22c7;
assign v8e42fd = jx2_p & v8e4d75 | !jx2_p & v8b54db;
assign v85b5f8 = ENQ_p & v8b5607 | !ENQ_p & v8af40a;
assign v8e58d8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e4e4e;
assign v85e8fd = BtoS_ACK0_p & v86290d | !BtoS_ACK0_p & v8e1cd3;
assign v85a894 = jx2_p & v858482 | !jx2_p & v844f91;
assign v845249 = BtoS_ACK0_p & v8b575f | !BtoS_ACK0_p & v8984b0;
assign v8e2177 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8e51f8;
assign v8b55a9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a5bc5;
assign v8e3bba = BtoS_ACK1_p & v8b5875 | !BtoS_ACK1_p & v8e5a76;
assign v8e44eb = StoB_REQ1_p & v8bf293 | !StoB_REQ1_p & v844f91;
assign v8e201e = BtoS_ACK1_p & v8e56eb | !BtoS_ACK1_p & v8b56ba;
assign v85d792 = BtoS_ACK1_p & v8e52b0 | !BtoS_ACK1_p & v8b5899;
assign v8b5538 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85aea9;
assign v85fa41 = BtoS_ACK0_p & v8b56e6 | !BtoS_ACK0_p & v8dc551;
assign v8b56bb = RtoB_ACK0_p & v8dc5de | !RtoB_ACK0_p & v856be5;
assign v85d428 = jx2_p & v844f91 | !jx2_p & v8e58fa;
assign v8450f8 = jx2_p & v867a85 | !jx2_p & v8e188a;
assign v8e20e3 = jx1_p & v8cc8ad | !jx1_p & !v8e400a;
assign v8e1d09 = BtoS_ACK8_p & v883b69 | !BtoS_ACK8_p & v8e17fe;
assign v860006 = stateG12_p & v8b5798 | !stateG12_p & !v85f9b8;
assign v8b553e = jx0_p & v8e4003 | !jx0_p & !v85d441;
assign v8b5786 = StoB_REQ0_p & v8e2381 | !StoB_REQ0_p & v844f91;
assign v8b558d = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8e3de2;
assign v85aa47 = StoB_REQ3_p & v856fe9 | !StoB_REQ3_p & v844f9f;
assign v8e2222 = jx2_p & v8e4ca6 | !jx2_p & v8e4397;
assign v8b5613 = RtoB_ACK1_p & v85769d | !RtoB_ACK1_p & v84521e;
assign v856556 = StoB_REQ2_p & v8b35e8 | !StoB_REQ2_p & v8e5426;
assign v8a5c45 = StoB_REQ6_p & v8b42e6 | !StoB_REQ6_p & v85ffcd;
assign v8e1add = jx1_p & v8e1975 | !jx1_p & v8e4786;
assign v8e213d = StoB_REQ2_p & v8e4f80 | !StoB_REQ2_p & v8e5965;
assign v8b5526 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v8e585b;
assign v8b57bb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b54d8;
assign v8606a9 = BtoS_ACK6_p & v85737f | !BtoS_ACK6_p & v8b56db;
assign v8b5678 = jx2_p & v8563b7 | !jx2_p & !v8e53ec;
assign v880dfd = StoB_REQ5_p & v867a58 | !StoB_REQ5_p & v844f91;
assign v8e1c12 = BtoS_ACK6_p & v8e2416 | !BtoS_ACK6_p & v845230;
assign v867aa7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e550e;
assign v8e5b48 = StoB_REQ6_p & v8e4fc9 | !StoB_REQ6_p & v844f91;
assign v86654a = RtoB_ACK1_p & v8b556b | !RtoB_ACK1_p & v8b5831;
assign v8e3cd1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b54c2;
assign v85f4fb = jx1_p & v85c93d | !jx1_p & v85a8af;
assign v8b54e9 = jx0_p & v844f91 | !jx0_p & v8e59b7;
assign v8e58a8 = StoB_REQ8_p & v8e4ea5 | !StoB_REQ8_p & v8b550e;
assign v8b55a5 = StoB_REQ8_p & v8b5621 | !StoB_REQ8_p & v867c19;
assign v85d7b1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85cd1c;
assign v856a38 = jx2_p & v8e4b4d | !jx2_p & !v89929e;
assign v8dc5be = BtoS_ACK7_p & v856264 | !BtoS_ACK7_p & v88c339;
assign v8e5bed = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v85f6bc;
assign v856395 = jx0_p & v844f91 | !jx0_p & v8e4d0c;
assign v8b5518 = jx1_p & v844f91 | !jx1_p & v8e57d3;
assign v85e1dd = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v8a5bbf;
assign v8e5914 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b3615;
assign v8e4913 = jx0_p & v8e4188 | !jx0_p & !v844f91;
assign v8e21d0 = jx1_p & v85dee1 | !jx1_p & !v8e5a9d;
assign v8b5899 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8b577f;
assign v8e2181 = BtoS_ACK0_p & v8e3d0c | !BtoS_ACK0_p & v8e190d;
assign v86654f = StoB_REQ1_p & v8e59e7 | !StoB_REQ1_p & v85d72c;
assign v845183 = StoB_REQ7_p & v8e5982 | !StoB_REQ7_p & v8b5889;
assign v8e179a = StoB_REQ0_p & v8e57b4 | !StoB_REQ0_p & v8e4e75;
assign v85e1a3 = ENQ_p & v8a3c77 | !ENQ_p & v85e664;
assign v85d7a6 = BtoR_REQ1_p & v8e158b | !BtoR_REQ1_p & v8562d4;
assign v8e5428 = jx0_p & v8af44d | !jx0_p & !v856594;
assign v8e59ae = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8b5659;
assign v8e14ab = jx1_p & v8a87cd | !jx1_p & v8e4a68;
assign v85d507 = BtoS_ACK8_p & v8e15fd | !BtoS_ACK8_p & v8e58a8;
assign v8e58b8 = ENQ_p & v8af34b | !ENQ_p & v8e114b;
assign v85b9de = jx1_p & v8a87cd | !jx1_p & v883cf8;
assign v85e274 = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v8e1c84;
assign v8af23a = StoB_REQ0_p & v8dc594 | !StoB_REQ0_p & v844f91;
assign v8e3f1b = jx2_p & v856c2e | !jx2_p & !v8cb249;
assign v865dba = jx3_p & v8e4ed1 | !jx3_p & v8e48f1;
assign v85dd75 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v898498;
assign v85702d = RtoB_ACK1_p & v889f0f | !RtoB_ACK1_p & v85dc42;
assign v844fa5 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v844f91;
assign v8e10aa = BtoS_ACK0_p & v8b5669 | !BtoS_ACK0_p & v8563a2;
assign v8564e9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8b5757;
assign v8b55c0 = StoB_REQ6_p & v8e23ae | !StoB_REQ6_p & v8af419;
assign v85d8e2 = BtoS_ACK8_p & v8e5a22 | !BtoS_ACK8_p & v8e5a62;
assign v856452 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8e519b;
assign v8e57d0 = StoB_REQ8_p & v8dc639 | !StoB_REQ8_p & v85d7c8;
assign v8e1d21 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8e5968;
assign v857107 = BtoR_REQ0_p & v8e3a67 | !BtoR_REQ0_p & v8b5848;
assign v8e4d29 = jx2_p & v8e4e99 | !jx2_p & !v889f6e;
assign v856ae7 = BtoS_ACK7_p & v85bdbc | !BtoS_ACK7_p & v8451d1;
assign v8b54ea = jx0_p & v8e3b31 | !jx0_p & v8e4d0c;
assign v8af325 = jx2_p & v8e4b4d | !jx2_p & !v8e16f6;
assign v8e197c = BtoR_REQ0_p & v8e39eb | !BtoR_REQ0_p & v8b55ed;
assign v8812e9 = BtoS_ACK6_p & v8e4a85 | !BtoS_ACK6_p & v8e535e;
assign v8e4a85 = jx2_p & v8e3db0 | !jx2_p & v85f57e;
assign v85e545 = BtoS_ACK6_p & v8568c2 | !BtoS_ACK6_p & v8b57ad;
assign v8e477d = StoB_REQ7_p & v8e4c47 | !StoB_REQ7_p & v8b56d6;
assign v8e4103 = stateG12_p & v85a893 | !stateG12_p & v844f91;
assign v8b54c0 = StoB_REQ6_p & v85cda6 | !StoB_REQ6_p & v8dc607;
assign v8af0d0 = StoB_REQ0_p & v885455 | !StoB_REQ0_p & v8e5428;
assign v8b585d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85df70;
assign v8b5605 = BtoS_ACK7_p & v8e1a5a | !BtoS_ACK7_p & v8e46d9;
assign v8e45c9 = StoB_REQ8_p & v8e4235 | !StoB_REQ8_p & v8e493e;
assign v8e59be = StoB_REQ0_p & v883ca3 | !StoB_REQ0_p & v8b585f;
assign v85d933 = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & v8892c1;
assign v8e3c65 = BtoS_ACK6_p & v8e4f36 | !BtoS_ACK6_p & v8e2098;
assign v85c8f2 = StoB_REQ6_p & v889f96 | !StoB_REQ6_p & v85fc4d;
assign v8450f2 = jx2_p & v8e59aa | !jx2_p & v8b552b;
assign v8e42f6 = ENQ_p & v8a3c77 | !ENQ_p & v8e572e;
assign v86ea54 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & v8584f3;
assign v8e416f = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v8e5924;
assign v8af41e = FULL_p & v8569df | !FULL_p & v85bbd9;
assign v85adf5 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v85710e;
assign v8e3b31 = BtoS_ACK1_p & v8b556f | !BtoS_ACK1_p & v88924e;
assign v85c4b8 = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & v8b5800;
assign v8e40f6 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8b558a;
assign v8e1650 = jx1_p & v8e15ab | !jx1_p & v85af76;
assign v8e3b37 = jx2_p & v85697c | !jx2_p & v844f91;
assign v8af2f2 = ENQ_p & v8562d0 | !ENQ_p & !v85664e;
assign v8b55cf = BtoS_ACK7_p & v8618f2 | !BtoS_ACK7_p & v8e4021;
assign v8a5cca = BtoS_ACK7_p & v85a008 | !BtoS_ACK7_p & v884771;
assign v85c469 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a5bcf;
assign v8e5778 = BtoS_ACK0_p & v8e46da | !BtoS_ACK0_p & v845187;
assign v85f1ac = BtoS_ACK0_p & v883ca3 | !BtoS_ACK0_p & v8e57b4;
assign v8650b9 = StoB_REQ3_p & v8e5000 | !StoB_REQ3_p & !v844f9f;
assign v85f3fb = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v889270;
assign v88c371 = jx1_p & v8be0ec | !jx1_p & v8e1b44;
assign v8b56b3 = StoB_REQ8_p & v8892c1 | !StoB_REQ8_p & v8e38ea;
assign v85760e = BtoS_ACK8_p & v863508 | !BtoS_ACK8_p & v8e2144;
assign v86299d = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v8b58b3;
assign v857423 = RtoB_ACK1_p & v8e4cfe | !RtoB_ACK1_p & v85b906;
assign v85dbb6 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v85e1b8;
assign v8e3dd3 = BtoS_ACK7_p & v8450b6 | !BtoS_ACK7_p & v8e4472;
assign v8b54f5 = StoB_REQ6_p & v85dbbe | !StoB_REQ6_p & v85dd22;
assign v85e619 = jx1_p & v88c355 | !jx1_p & !v85cc2a;
assign v8dc5de = BtoR_REQ1_p & v8b55c7 | !BtoR_REQ1_p & v88c2f6;
assign v8e493e = BtoS_ACK7_p & v8e1b8d | !BtoS_ACK7_p & v8e5936;
assign v8e3c3e = BtoS_ACK0_p & v8e3ac5 | !BtoS_ACK0_p & v8e479e;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v8e57c9 = BtoS_ACK7_p & v8e436b | !BtoS_ACK7_p & v8e3bda;
assign v85bbb8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e1770;
assign v85bd3d = BtoR_REQ1_p & v856261 | !BtoR_REQ1_p & !v8e3fe8;
assign v85b514 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8af46d;
assign v856364 = EMPTY_p & v8e5a13 | !EMPTY_p & v8e591f;
assign v8e4588 = BtoS_ACK2_p & v85725c | !BtoS_ACK2_p & v8e4cc0;
assign v8567fa = StoB_REQ7_p & v8e49b1 | !StoB_REQ7_p & v85ea86;
assign v89924f = jx2_p & v865810 | !jx2_p & !v85ffcd;
assign v85d533 = BtoS_ACK8_p & v8e5a22 | !BtoS_ACK8_p & v8e5a6f;
assign v8b5789 = jx2_p & v8e4337 | !jx2_p & v85f218;
assign v8e3883 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b5875;
assign v859fe5 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8e51cf;
assign v8e4096 = RtoB_ACK1_p & v85f194 | !RtoB_ACK1_p & v8b57b7;
assign v860053 = RtoB_ACK0_p & v85ca46 | !RtoB_ACK0_p & v8e4cf4;
assign v85d914 = jx2_p & v8e44c7 | !jx2_p & v8b58bb;
assign v8dc57c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5674;
assign v8e4f5f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e3b8b;
assign v84513a = BtoS_ACK0_p & v8b5893 | !BtoS_ACK0_p & v8e479e;
assign v8e4db2 = BtoS_ACK1_p & v85dbdd | !BtoS_ACK1_p & v8ce3d5;
assign v8dc599 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4d7b;
assign v8b54f9 = stateG7_1_p & v8e44a2 | !stateG7_1_p & v8b55f0;
assign v8e1f0e = RtoB_ACK0_p & v8e3ff5 | !RtoB_ACK0_p & v8a555c;
assign v8e1f74 = BtoS_ACK1_p & v8e1692 | !BtoS_ACK1_p & v8e22bd;
assign v8af457 = DEQ_p & v8e54cf | !DEQ_p & v8b55ed;
assign v85cdde = RtoB_ACK0_p & v8e1823 | !RtoB_ACK0_p & v85f8da;
assign v85e3d2 = RtoB_ACK0_p & v8e48fc | !RtoB_ACK0_p & v85c73d;
assign v8e5298 = BtoS_ACK0_p & v88d5d7 | !BtoS_ACK0_p & v85ba51;
assign v8e438f = DEQ_p & v85bbcc | !DEQ_p & v86290d;
assign v8e5366 = StoB_REQ7_p & v8e462b | !StoB_REQ7_p & v856ecb;
assign v8a5bc5 = jx0_p & v88c324 | !jx0_p & v86ea54;
assign v8e4bb0 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8b35e8;
assign v85c7b4 = StoB_REQ2_p & v8e3f79 | !StoB_REQ2_p & v8e5a2a;
assign v8e4188 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85c469;
assign v8b5505 = jx1_p & v8e5a2d | !jx1_p & v86290d;
assign v8e5a76 = BtoS_ACK2_p & v8b5875 | !BtoS_ACK2_p & !v8b5830;
assign v8dc552 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & v8e59c0;
assign v85ea86 = StoB_REQ6_p & v8e3af1 | !StoB_REQ6_p & v8e3bf3;
assign v8e4bc9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e4e56;
assign v8e59fd = FULL_p & v8b57a9 | !FULL_p & v8cc95b;
assign v85df15 = jx2_p & v8563f1 | !jx2_p & v85653c;
assign v85a05d = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856598;
assign v85667b = EMPTY_p & v8cce0d | !EMPTY_p & v8565ea;
assign v856c55 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85dce5;
assign v8e41d0 = jx1_p & v844f91 | !jx1_p & v8af46d;
assign v85d3b1 = EMPTY_p & v8b569b | !EMPTY_p & v8e3d66;
assign v8e4cb9 = jx2_p & v8b5601 | !jx2_p & v85e619;
assign v8e20ba = stateG7_1_p & v8566fa | !stateG7_1_p & v8e42ab;
assign v85c83d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88c2f2;
assign v85d72c = BtoS_ACK2_p & v8b550c | !BtoS_ACK2_p & !v8b562e;
assign v86e0c8 = jx1_p & v856c71 | !jx1_p & v85d43b;
assign v8e152b = jx0_p & v8e5a69 | !jx0_p & v844f91;
assign v8e5881 = ENQ_p & v8b5607 | !ENQ_p & v8e1be0;
assign v8e5998 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e23b1;
assign v845079 = StoB_REQ6_p & v8e590b | !StoB_REQ6_p & v8e1ee5;
assign v89920d = jx0_p & v844f91 | !jx0_p & v8b55cb;
assign v8b5707 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8e3d40;
assign v85d79a = BtoS_ACK8_p & v8b58bb | !BtoS_ACK8_p & v8b586b;
assign v8e4345 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856f79;
assign v8e5155 = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & !v85ad92;
assign v85d2e2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e42c6;
assign v8e59af = EMPTY_p & v8b5760 | !EMPTY_p & v85af2b;
assign v8b55ec = BtoR_REQ1_p & v8e1c7f | !BtoR_REQ1_p & !v856261;
assign v8e4cc0 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e5a55;
assign v8a5c2b = jx0_p & v85f50b | !jx0_p & v844f91;
assign v8a5bd1 = jx0_p & v8e4212 | !jx0_p & v8e4059;
assign v8b56e8 = BtoS_ACK8_p & v8e4b00 | !BtoS_ACK8_p & v8e48d8;
assign v85df40 = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & v8e49c8;
assign v8e18ff = DEQ_p & v85ae77 | !DEQ_p & v85f2b2;
assign v85df5b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85b739;
assign v8e1abd = BtoS_ACK7_p & v85d805 | !BtoS_ACK7_p & v85deb3;
assign v8b35f0 = jx1_p & v881bc6 | !jx1_p & v844f91;
assign v888cd4 = RtoB_ACK0_p & v8b5565 | !RtoB_ACK0_p & !v844f91;
assign v85fc4d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v889f3d;
assign v8e5a31 = BtoS_ACK0_p & v8af418 | !BtoS_ACK0_p & v8b577c;
assign v85f340 = BtoS_ACK0_p & v8e388e | !BtoS_ACK0_p & v8e5022;
assign v860886 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8e21b3;
assign v856883 = StoB_REQ1_p & v8b54c4 | !StoB_REQ1_p & v85626a;
assign v8563cb = RtoB_ACK1_p & v8e589c | !RtoB_ACK1_p & v8e1f0e;
assign v8e5212 = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8574cc;
assign v85dfaa = EMPTY_p & v85760e | !EMPTY_p & v85a4f0;
assign v8e588e = StoB_REQ6_p & v84530d | !StoB_REQ6_p & !v85dda8;
assign v85a1f0 = StoB_REQ7_p & v8e5212 | !StoB_REQ7_p & v85fa64;
assign v85deeb = RtoB_ACK1_p & v8e48fc | !RtoB_ACK1_p & v85e3d2;
assign v85e3a8 = jx1_p & v8e4514 | !jx1_p & v8b570e;
assign v8b57fa = BtoS_ACK8_p & v8af4c2 | !BtoS_ACK8_p & v85fa42;
assign v880bc3 = jx3_p & v844f91 | !jx3_p & !v8e1e94;
assign v8e111b = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & !v8e17b2;
assign v8574d0 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8e4caf;
assign v8e20f6 = StoB_REQ0_p & v8e4a22 | !StoB_REQ0_p & v8e4f8b;
assign v8e46b2 = jx1_p & v8e59f6 | !jx1_p & !v8af0dc;
assign v8e5939 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b563d;
assign v8564ef = jx1_p & v844f91 | !jx1_p & v85b514;
assign v8b5809 = DEQ_p & v8b562d | !DEQ_p & v844f91;
assign v85af8a = jx1_p & v8e4514 | !jx1_p & v85e27e;
assign v856b71 = BtoS_ACK8_p & v85a008 | !BtoS_ACK8_p & v889f0e;
assign v8b56b7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v85df2b;
assign v8af3c1 = EMPTY_p & v856ec1 | !EMPTY_p & v8e3c8e;
assign v85dc0d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b57d8;
assign v85769d = BtoR_REQ1_p & v8e593f | !BtoR_REQ1_p & v8e58dd;
assign v8e5a3e = jx1_p & v85db8a | !jx1_p & !v8e46ed;
assign v85ba2c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b551a;
assign v8e4791 = jx0_p & v8cce14 | !jx0_p & !v8a6d22;
assign v8e566a = StoB_REQ1_p & v8e436c | !StoB_REQ1_p & v8b586f;
assign v856edd = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8e1e8c;
assign v85ac27 = BtoS_ACK0_p & v85d90a | !BtoS_ACK0_p & v8e3d2a;
assign v8e1a5a = jx2_p & v85d434 | !jx2_p & v85dfab;
assign v8e4fe9 = EMPTY_p & v860057 | !EMPTY_p & v86514d;
assign v85deb5 = jx2_p & v856e1f | !jx2_p & !v8e4e45;
assign v8e58fa = jx1_p & v85f340 | !jx1_p & v844f91;
assign v8b583e = jx0_p & v85e82e | !jx0_p & v889f3d;
assign v85e858 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v8e1d78;
assign v856b4b = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8564f5;
assign v85d52e = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v85b739;
assign v8847b9 = StoB_REQ1_p & v8e4f80 | !StoB_REQ1_p & v8b56fa;
assign v8e4007 = jx2_p & v8e58a6 | !jx2_p & v85da0f;
assign v8571db = jx1_p & v8b57df | !jx1_p & v86dabf;
assign v8b5585 = EMPTY_p & v8b55ed | !EMPTY_p & v8b55e9;
assign v8e38d9 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844fb5;
assign v8e1b8d = jx2_p & v85afea | !jx2_p & v8e15b2;
assign v8e23df = BtoS_ACK7_p & v8e2025 | !BtoS_ACK7_p & v856b41;
assign v85e281 = jx2_p & v84520f | !jx2_p & !v8e2355;
assign v8e4ebc = StoB_REQ1_p & v85df25 | !StoB_REQ1_p & v8e3ea2;
assign v8b55fc = BtoS_ACK2_p & v85725c | !BtoS_ACK2_p & v8b5640;
assign v85dbf1 = RtoB_ACK1_p & v8b56ad | !RtoB_ACK1_p & v8e4941;
assign v85dcb6 = RtoB_ACK1_p & v85ab00 | !RtoB_ACK1_p & v845281;
assign v8892bc = EMPTY_p & v8e44a9 | !EMPTY_p & v8e1e6c;
assign v8e4831 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4637;
assign v86514d = DEQ_p & v8e1cd8 | !DEQ_p & v860057;
assign v8b5794 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4c7f;
assign v85a648 = jx1_p & v8e4fe5 | !jx1_p & v8e22f8;
assign v8e17fe = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v85f52f;
assign v8e3b0a = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8e47ef;
assign v8dc571 = BtoS_ACK6_p & v8b583c | !BtoS_ACK6_p & v8e5985;
assign v8e1d94 = StoB_REQ0_p & v8e5033 | !StoB_REQ0_p & v844f91;
assign v85670f = BtoS_ACK0_p & v8dc594 | !BtoS_ACK0_p & v8991c9;
assign v8e5c1b = StoB_REQ6_p & v8b588c | !StoB_REQ6_p & v8e4d7d;
assign v8e14bc = StoB_REQ6_p & v8e5b0f | !StoB_REQ6_p & v8b566c;
assign v8e4cfe = BtoR_REQ1_p & v85dcee | !BtoR_REQ1_p & v860902;
assign v8e3b2f = BtoS_ACK7_p & v8e5a5e | !BtoS_ACK7_p & v85d9f0;
assign v88c32e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v86e38c;
assign v8e482a = jx1_p & v85f42f | !jx1_p & v8e1755;
assign v85d6a8 = jx2_p & v85a07c | !jx2_p & !v844f91;
assign v85c7af = jx1_p & v85bbb8 | !jx1_p & v844f91;
assign v85daf5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f97;
assign v8b5832 = BtoS_ACK6_p & v8e10c3 | !BtoS_ACK6_p & v85fb1e;
assign v8b54e1 = StoB_REQ7_p & v8e1fe7 | !StoB_REQ7_p & !v844f91;
assign v8574d6 = jx1_p & v8451a1 | !jx1_p & v8dc599;
assign v8e4036 = BtoS_ACK7_p & v8e4764 | !BtoS_ACK7_p & v8e4e25;
assign v85a6d2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85b390;
assign v85725c = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8e16ea;
assign v8563c0 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v8e3ff2;
assign v88bc46 = BtoS_ACK8_p & v8af4aa | !BtoS_ACK8_p & v8e520d;
assign v8e4d8f = BtoS_ACK2_p & v85725c | !BtoS_ACK2_p & v8e1480;
assign v8e3b5f = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v856bb4;
assign v844faf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v86c57a = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & !v856e07;
assign v8b589b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5367;
assign v85dff8 = BtoS_ACK0_p & v889f88 | !BtoS_ACK0_p & v8af41c;
assign v8e4f16 = jx2_p & v8e1bf9 | !jx2_p & !v8e4c34;
assign v8a87fd = jx2_p & v85f4fb | !jx2_p & v844f91;
assign v8e3af2 = stateG12_p & v8e1c59 | !stateG12_p & !v865764;
assign v8e2282 = StoB_REQ1_p & v861740 | !StoB_REQ1_p & v85650e;
assign v8e5060 = jx1_p & v8e1c72 | !jx1_p & v88c2be;
assign v8e57b4 = jx0_p & v85e7be | !jx0_p & !v844f91;
assign v8585f1 = stateG12_p & v8cce0d | !stateG12_p & v844f91;
assign v85d340 = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & v8e5266;
assign v85658e = BtoS_ACK0_p & v8e5a1c | !BtoS_ACK0_p & v8e5914;
assign v8e3917 = jx1_p & v844f91 | !jx1_p & v8b5677;
assign v8e3b75 = BtoS_ACK0_p & v8a9208 | !BtoS_ACK0_p & v8b55b8;
assign v8a554f = BtoS_ACK6_p & v856a03 | !BtoS_ACK6_p & v8e472c;
assign v8b577d = StoB_REQ0_p & v883ca3 | !StoB_REQ0_p & v8b5663;
assign v85dbf7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4a57;
assign v8e4e75 = jx0_p & v8e3b31 | !jx0_p & !v86f856;
assign v856353 = BtoS_ACK8_p & v85b66d | !BtoS_ACK8_p & v8e3db6;
assign v8e3b8b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v85b69f;
assign v8e1dbf = ENQ_p & v8572d0 | !ENQ_p & v8e3ffc;
assign v85e4bb = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8e17d6;
assign v85dce5 = BtoS_ACK0_p & v85699e | !BtoS_ACK0_p & v8e599d;
assign v85dd7c = jx1_p & v8b56ee | !jx1_p & !v844f91;
assign v863508 = jx2_p & v85d3f6 | !jx2_p & v86290f;
assign v8e1667 = StoB_REQ0_p & v8991c9 | !StoB_REQ0_p & v8dc555;
assign v8e598b = EMPTY_p & v8601d6 | !EMPTY_p & v856913;
assign v8e4a48 = StoB_REQ8_p & v8b5826 | !StoB_REQ8_p & v8af107;
assign v8af2e0 = jx2_p & v8e5891 | !jx2_p & v8e4397;
assign v845150 = BtoS_ACK0_p & v85f6bc | !BtoS_ACK0_p & v8b565d;
assign v8e39ff = jx0_p & v8dc552 | !jx0_p & v8e4831;
assign v86066c = BtoS_ACK1_p & v85c632 | !BtoS_ACK1_p & !v867a75;
assign v85e8b5 = BtoS_ACK7_p & v85737f | !BtoS_ACK7_p & v864971;
assign v8e5054 = jx1_p & v8b589b | !jx1_p & !v8e3b66;
assign v8e5032 = StoB_REQ2_p & v8e5a8f | !StoB_REQ2_p & v844f91;
assign v8e1f2a = jx1_p & v844f91 | !jx1_p & !v85f422;
assign v8af107 = BtoS_ACK7_p & v856fa4 | !BtoS_ACK7_p & !v85b99e;
assign v85ffb3 = ENQ_p & v8e4e6e | !ENQ_p & v8e55ba;
assign v8e5958 = BtoR_REQ0_p & v8e5a5a | !BtoR_REQ0_p & v8e579b;
assign v856eb5 = StoB_REQ0_p & v85f2f8 | !StoB_REQ0_p & v85dfad;
assign v8e47e7 = BtoS_ACK7_p & v85c5cf | !BtoS_ACK7_p & !v8e59b9;
assign v8e10b7 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & v856eba;
assign v864623 = StoB_REQ7_p & v8e49b1 | !StoB_REQ7_p & v8e3bf3;
assign v85e694 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v8e1d33;
assign v8e5982 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v844f97;
assign v8572c2 = StoB_REQ6_p & v8af3f2 | !StoB_REQ6_p & v844f91;
assign v8af268 = jx0_p & v8b5807 | !jx0_p & v8e583f;
assign v8b5801 = StoB_REQ8_p & v889350 | !StoB_REQ8_p & v8b5756;
assign v867a93 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85d7bb;
assign v8b5830 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8b56bd;
assign BtoR_REQ0_n = !v8672d0;
assign v865856 = jx2_p & v8e10a4 | !jx2_p & v8e41ec;
assign v8a691b = StoB_REQ7_p & v85a8af | !StoB_REQ7_p & v8e1a78;
assign v8e596c = StoB_REQ7_p & v8b56e5 | !StoB_REQ7_p & v844f91;
assign v85aef4 = jx1_p & v8e59ee | !jx1_p & v844f91;
assign v8e530b = StoB_REQ7_p & v8e58ce | !StoB_REQ7_p & !v8e5c1b;
assign v8452cd = StoB_REQ6_p & v8e4c47 | !StoB_REQ6_p & v8e2000;
assign v865f86 = jx0_p & v8b5500 | !jx0_p & v8e58d9;
assign v8e1765 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e22d4;
assign v8e4021 = BtoS_ACK6_p & v8e40ce | !BtoS_ACK6_p & v85a25b;
assign v8e5498 = jx1_p & v8b5679 | !jx1_p & !v8e47f8;
assign v8b571d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e5c6a;
assign v899202 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v844f91;
assign v8e5833 = jx2_p & v866529 | !jx2_p & v85653c;
assign v85e006 = BtoS_ACK0_p & v8e58cb | !BtoS_ACK0_p & v85dddb;
assign v8e1800 = jx1_p & v8a5c45 | !jx1_p & !v8e1be3;
assign v8e5909 = BtoR_REQ1_p & v8e2239 | !BtoR_REQ1_p & !v8cce0a;
assign v8b5762 = BtoS_ACK6_p & v85737f | !BtoS_ACK6_p & v8e4aec;
assign v85ae77 = stateG12_p & v85f2b2 | !stateG12_p & v844f91;
assign v845281 = RtoB_ACK0_p & v8e198b | !RtoB_ACK0_p & v8e58e9;
assign v8e3d20 = StoB_REQ3_p & v867a58 | !StoB_REQ3_p & v880dfd;
assign v86e720 = BtoS_ACK0_p & v85f59b | !BtoS_ACK0_p & v85c771;
assign v863b23 = jx1_p & v8e4514 | !jx1_p & v8e197f;
assign v8e511b = jx1_p & v8991fe | !jx1_p & v85a8af;
assign v8e2079 = jx1_p & v86290d | !jx1_p & !v8e4a68;
assign v8e59c9 = StoB_REQ8_p & v85da27 | !StoB_REQ8_p & v8564fa;
assign v8e53e7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b5517;
assign v856473 = BtoS_ACK6_p & v8b55b0 | !BtoS_ACK6_p & v85d428;
assign v85dbdd = StoB_REQ5_n & v844f91 | !StoB_REQ5_n & v844f9d;
assign v88927c = BtoS_ACK8_p & v8b54dc | !BtoS_ACK8_p & v845386;
assign v85af76 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85e8a6;
assign v844f9f = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & !v844f91;
assign v8e19c7 = jx1_p & v85ccdf | !jx1_p & v8e1d5f;
assign v89928e = BtoS_ACK6_p & v8af325 | !BtoS_ACK6_p & v8e599e;
assign v865125 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85ad2e;
assign v85e1bb = jx0_p & v844f91 | !jx0_p & v8b552d;
assign v8e3e66 = BtoS_ACK7_p & v8b561b | !BtoS_ACK7_p & !v8af21d;
assign v85e895 = jx1_p & v8e5a64 | !jx1_p & !v844f91;
assign v8b5533 = BtoS_ACK1_p & v8b5875 | !BtoS_ACK1_p & v8e192f;
assign v856b8f = jx1_p & v8e44dd | !jx1_p & v8b57da;
assign v8b5682 = ENQ_p & v8a3c77 | !ENQ_p & v86cbc7;
assign v8e3c81 = BtoS_ACK0_p & v8dc594 | !BtoS_ACK0_p & v8a54f3;
assign v8b5522 = RtoB_ACK0_p & v8e1c89 | !RtoB_ACK0_p & v856afe;
assign v85a880 = BtoS_ACK7_p & v8e1f55 | !BtoS_ACK7_p & !v845033;
assign v85ca01 = StoB_REQ6_p & v8e5a9d | !StoB_REQ6_p & v8e5a39;
assign v889f73 = BtoS_ACK0_p & v8e5917 | !BtoS_ACK0_p & v85e942;
assign v8b567a = jx1_p & v85aeb5 | !jx1_p & !v8e1bb4;
assign v8e2091 = StoB_REQ7_p & v8e5a31 | !StoB_REQ7_p & v8e57ee;
assign v85e50d = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8e2399;
assign v8e1199 = BtoS_ACK0_p & v8e4f71 | !BtoS_ACK0_p & v8e58f1;
assign v84518f = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8e1eb4;
assign v845379 = jx0_p & v8af277 | !jx0_p & v8e43f1;
assign v85e8f2 = BtoS_ACK6_p & v8e420a | !BtoS_ACK6_p & v85e8f4;
assign v8af188 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v881da6;
assign v8e3c25 = StoB_REQ7_p & v8e17f5 | !StoB_REQ7_p & v8e59be;
assign v85f48a = ENQ_p & v8b5607 | !ENQ_p & v85fac2;
assign v8b5551 = BtoS_ACK0_p & v8e17e8 | !BtoS_ACK0_p & v8b571d;
assign v8b5733 = BtoS_ACK1_p & v8e4632 | !BtoS_ACK1_p & v8575eb;
assign v880b52 = BtoS_ACK0_p & v85e0b0 | !BtoS_ACK0_p & v87c63e;
assign v8e1f85 = BtoS_ACK0_p & v889f3d | !BtoS_ACK0_p & v8e4b0e;
assign v8e5ad2 = ENQ_p & v85e45f | !ENQ_p & v862c12;
assign v8e5a27 = StoB_REQ6_p & v8a5b53 | !StoB_REQ6_p & v8e1b43;
assign v8b5812 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b575f;
assign v856eeb = BtoS_ACK7_p & v8e4235 | !BtoS_ACK7_p & v85dbf8;
assign v85cd17 = BtoS_ACK6_p & v85737f | !BtoS_ACK6_p & v8b578b;
assign v86695b = BtoS_ACK7_p & v8e1933 | !BtoS_ACK7_p & v8e4b9b;
assign v8b5779 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e2060;
assign v8e58d3 = StoB_REQ6_p & v8e16ce | !StoB_REQ6_p & v8e5a68;
assign v85c941 = jx0_p & v844f91 | !jx0_p & !v8b5893;
assign v85f401 = StoB_REQ8_p & v85736b | !StoB_REQ8_p & v8e46fa;
assign v884319 = jx2_p & v8e59de | !jx2_p & v8565fe;
assign v8b5569 = jx1_p & v8be0f9 | !jx1_p & !v844f91;
assign v85c9c5 = jx0_p & v844f91 | !jx0_p & !v8e4831;
assign v8e5a62 = StoB_REQ8_p & v8e5887 | !StoB_REQ8_p & v8cc8ae;
assign v8cc8fa = BtoS_ACK7_p & v8450b6 | !BtoS_ACK7_p & v8b57f3;
assign v8b570c = jx1_p & v85acf3 | !jx1_p & !v8b56c3;
assign v8e4e56 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85bdac;
assign v8e59d4 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b57fc;
assign v8b55d4 = BtoS_ACK3_p & v85dbdd | !BtoS_ACK3_p & v86b9f0;
assign v88934b = EMPTY_p & v8b5506 | !EMPTY_p & v8b54ec;
assign v8e159f = BtoS_ACK0_p & v8e5913 | !BtoS_ACK0_p & v8e56cb;
assign v8b5863 = jx2_p & v856ef1 | !jx2_p & !v85b036;
assign v8b55c5 = jx2_p & v8b560e | !jx2_p & v856801;
assign v8b5679 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e3cd1;
assign v8b5720 = jx2_p & v88460a | !jx2_p & v8e58e0;
assign v8571d6 = jx2_p & v8b55c3 | !jx2_p & v856b8f;
assign v85d382 = BtoS_ACK0_p & v8e4c47 | !BtoS_ACK0_p & v8e4791;
assign v85d475 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85dbb6;
assign v85e332 = StoB_REQ7_p & v86290d | !StoB_REQ7_p & v85e1dd;
assign v8b5891 = RtoB_ACK1_p & v8e3fa0 | !RtoB_ACK1_p & v8e1ed4;
assign v8e4a95 = StoB_REQ1_p & v8e5bb2 | !StoB_REQ1_p & v844f91;
assign v8e48d7 = StoB_REQ0_p & v8dc594 | !StoB_REQ0_p & v8e5917;
assign v8a5bcf = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v85dbdd;
assign v8e5c6a = jx0_p & v8af277 | !jx0_p & v8e5920;
assign v85c7c5 = jx1_p & v8e4574 | !jx1_p & !v8e4c47;
assign v85b09e = StoB_REQ0_p & v882912 | !StoB_REQ0_p & v8b55cb;
assign v8e41a5 = EMPTY_p & v889f94 | !EMPTY_p & v8e14ca;
assign v8b5879 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8a54e5;
assign v8e5a63 = StoB_REQ7_p & v8e3eb2 | !StoB_REQ7_p & v8e4a68;
assign v8b584e = EMPTY_p & v8635e4 | !EMPTY_p & v857056;
assign v8a5b1b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e3cb6;
assign v8b56d2 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85ba51;
assign v8e4432 = BtoS_ACK8_p & v8af325 | !BtoS_ACK8_p & v8e4036;
assign v8dc580 = StoB_REQ1_p & v8a5b4f | !StoB_REQ1_p & v844f91;
assign v8e422f = StoB_REQ7_p & v8567bb | !StoB_REQ7_p & v8e45c6;
assign v8af231 = StoB_REQ8_p & v856eeb | !StoB_REQ8_p & v85a0ae;
assign v85f8fd = jx1_p & v8b560a | !jx1_p & !v8b5827;
assign v86e551 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v89b6ce;
assign v8e164c = jx0_p & v88bcd0 | !jx0_p & !v8e4605;
assign v8e1638 = StoB_REQ0_p & v8e4791 | !StoB_REQ0_p & v85b54e;
assign v8e5a6e = DEQ_p & v85663a | !DEQ_p & v85e81e;
assign v8e5223 = jx2_p & v8cce2b | !jx2_p & v8571db;
assign v861740 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e3bef;
assign v8566f1 = StoB_REQ7_p & v85dee5 | !StoB_REQ7_p & v8e22c7;
assign v8e3d3c = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v86650a;
assign v85722b = BtoS_ACK7_p & v8e594c | !BtoS_ACK7_p & !v8af37d;
assign v85dbad = jx1_p & v85670f | !jx1_p & !v8b56d2;
assign v8e39e1 = RtoB_ACK1_p & v8e431c | !RtoB_ACK1_p & !v856404;
assign v8b582f = StoB_REQ0_p & v856395 | !StoB_REQ0_p & v8b54ea;
assign v8e38cd = BtoS_ACK8_p & v8e15fd | !BtoS_ACK8_p & v8b5842;
assign v85da39 = jx0_p & v86baf9 | !jx0_p & v8e3dcc;
assign v86e4e7 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9d;
assign v85ad62 = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8e3df8;
assign v86cb45 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e1c26;
assign v8893ab = BtoR_REQ0_p & v867a97 | !BtoR_REQ0_p & v8cce0d;
assign v8b5844 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v866544;
assign v8658a0 = ENQ_p & v85ba14 | !ENQ_p & v85fb12;
assign v8e5913 = jx0_p & v8b56ce | !jx0_p & !v844f9d;
assign v8e5aa8 = ENQ_p & v85e45f | !ENQ_p & v85d933;
assign v85b6b5 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85e18a;
assign v8b55cb = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v8e41fc = ENQ_p & v8af46c | !ENQ_p & v8e4b2c;
assign v8e420a = jx2_p & v844f91 | !jx2_p & !v8e238d;
assign v86584f = jx1_p & v8e5bd2 | !jx1_p & v8b55ff;
assign v8b572f = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v867a58;
assign v865770 = DEQ_p & v8e1bda | !DEQ_p & v8b5814;
assign v882156 = StoB_REQ0_p & v8e1084 | !StoB_REQ0_p & v8e10b7;
assign v8e4163 = BtoS_ACK1_p & v8e52b0 | !BtoS_ACK1_p & v8e58d7;
assign v8e19c3 = jx1_p & v8e58e8 | !jx1_p & !v865802;
assign v86f856 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v86f9a1;
assign v85b29f = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v858462;
assign v8e592f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8574d0;
assign v85a07c = jx1_p & v8e1982 | !jx1_p & v844f91;
assign v8e1090 = ENQ_p & v844f91 | !ENQ_p & v8e228f;
assign v8e5510 = RtoB_ACK0_p & v8af3c1 | !RtoB_ACK0_p & !v844f91;
assign v8e4f71 = StoB_REQ1_p & v8e4637 | !StoB_REQ1_p & v844f91;
assign v8b580f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85d9d8;
assign v8b57f2 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v86e8c2;
assign v85a6a9 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8af160;
assign v8e388a = jx1_p & v85dee1 | !jx1_p & !v8dc612;
assign v8b583b = jx2_p & v873e9c | !jx2_p & v86d6bd;
assign v8e58cd = jx1_p & v8e3ae7 | !jx1_p & v8b5538;
assign v85b06b = BtoR_REQ1_p & v88934e | !BtoR_REQ1_p & v8e1c96;
assign v8cc95a = ENQ_p & v8572d0 | !ENQ_p & v88927c;
assign v85665c = StoB_REQ8_p & v8b573e | !StoB_REQ8_p & v8e58f5;
assign v8e4022 = ENQ_p & v8e3a26 | !ENQ_p & v8e4432;
assign v8e3dad = jx1_p & v8e2431 | !jx1_p & !v8e5a63;
assign v8e3c39 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & v85d7b1;
assign v8e39c1 = jx0_p & v844f91 | !jx0_p & v889f3d;
assign v8e58d4 = BtoS_ACK8_p & v8af325 | !BtoS_ACK8_p & v86513d;
assign v8b57e0 = BtoS_ACK6_p & v85ad82 | !BtoS_ACK6_p & v8e4cfc;
assign v856a23 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e509c;
assign v8e47f2 = jx0_p & v844f91 | !jx0_p & !v86f856;
assign v865836 = jx1_p & v85aeb5 | !jx1_p & v844f91;
assign v8e4397 = jx1_p & v8e422f | !jx1_p & v845189;
assign v84521e = RtoB_ACK0_p & v8e5958 | !RtoB_ACK0_p & v8e591c;
assign v856390 = StoB_REQ6_p & v86007f | !StoB_REQ6_p & v8e5085;
assign v856f08 = jx2_p & v8e207d | !jx2_p & v8b5689;
assign v8b55a0 = StoB_REQ8_p & v85e8b5 | !StoB_REQ8_p & v8af2be;
assign v8567d9 = ENQ_p & v85e45f | !ENQ_p & v8665a0;
assign v8665a9 = StoB_REQ3_p & v85ea8d | !StoB_REQ3_p & v8e5a72;
assign v85f1cb = BtoS_ACK0_p & v8e3eb2 | !BtoS_ACK0_p & v8e51f4;
assign v8b56fb = jx2_p & v8b5643 | !jx2_p & v844f91;
assign v8e3cfe = ENQ_p & v8b5607 | !ENQ_p & v844f91;
assign v85e0ba = BtoS_ACK7_p & v85e947 | !BtoS_ACK7_p & v8b588a;
assign v8e589b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e5917;
assign v85dd3e = jx1_p & v8ca185 | !jx1_p & !v8e3b66;
assign v889fde = jx0_p & v8b5856 | !jx0_p & !v8e5977;
assign v856fa4 = jx2_p & v8e54fe | !jx2_p & !v8b5895;
assign v8b5669 = jx0_p & v844f91 | !jx0_p & v856594;
assign v8e5a72 = StoB_REQ5_n & v8b56bd | !StoB_REQ5_n & v85ea8d;
assign v8e1862 = stateG7_1_p & v8dc6bf | !stateG7_1_p & v8e5b16;
assign v8e469a = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v856fe9;
assign v859fe9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b56ce;
assign v85db26 = jx2_p & v8b57e2 | !jx2_p & v8e41d0;
assign v8e1d33 = StoB_REQ5_p & v85ea8d | !StoB_REQ5_p & v844fb7;
assign v844fc9 = ENQ_p & v844f91 | !ENQ_p & !v844f91;
assign v8665a0 = BtoS_ACK8_p & v85a98f | !BtoS_ACK8_p & v8e57d0;
assign v8e3de0 = jx1_p & v8a87cd | !jx1_p & v8b56d6;
assign v85ab77 = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & v899283;
assign v8e45a4 = BtoS_ACK6_p & v8b56ae | !BtoS_ACK6_p & v880b7a;
assign v8e5a1c = jx0_p & v8b588b | !jx0_p & v8dc580;
assign v8b56ec = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8665a9;
assign v85e362 = jx0_p & v85b6b5 | !jx0_p & !v8b5567;
assign v8b5732 = ENQ_p & v844fbf | !ENQ_p & !v8b55a4;
assign v8e1964 = StoB_REQ8_p & v85da27 | !StoB_REQ8_p & v8b5684;
assign v856fdc = BtoS_ACK8_p & v8b56a5 | !BtoS_ACK8_p & v8e2213;
assign v8b57b3 = jx0_p & v8b5807 | !jx0_p & v8569c1;
assign v889350 = BtoS_ACK7_p & v85e947 | !BtoS_ACK7_p & v856473;
assign v856fba = StoB_REQ8_p & v85ad0c | !StoB_REQ8_p & v8e1e31;
assign v8e1ebe = BtoS_ACK6_p & v85bd7c | !BtoS_ACK6_p & v86290d;
assign v8e1961 = BtoS_ACK8_p & v882bc3 | !BtoS_ACK8_p & !v845069;
assign v8e4805 = ENQ_p & v8e4e6e | !ENQ_p & v85d79a;
assign v8e1484 = BtoS_ACK0_p & v899247 | !BtoS_ACK0_p & v85fbed;
assign v8e57a6 = jx1_p & v889f8a | !jx1_p & v85a8af;
assign v8e4468 = jx0_p & v8b56ce | !jx0_p & v844f91;
assign v85d42f = BtoS_ACK2_p & v85dbdd | !BtoS_ACK2_p & !v85ea8d;
assign v85b2e6 = BtoS_ACK0_p & v8b57be | !BtoS_ACK0_p & v8564e9;
assign v8e49d3 = BtoS_ACK1_p & v85c469 | !BtoS_ACK1_p & v8e1756;
assign v8565fe = jx1_p & v85e8bf | !jx1_p & v8e58ce;
assign v8e14dc = jx2_p & v8e1add | !jx2_p & v8e4603;
assign v85d43b = StoB_REQ7_p & v8e209c | !StoB_REQ7_p & v8e2303;
assign v8b5555 = BtoS_ACK6_p & v8e4877 | !BtoS_ACK6_p & v85a9b1;
assign v8e49b1 = StoB_REQ0_p & v8e5033 | !StoB_REQ0_p & v8b55cb;
assign v8565bb = BtoS_ACK6_p & v89924f | !BtoS_ACK6_p & v8566db;
assign v8e4cc7 = BtoS_ACK0_p & v8e5b6b | !BtoS_ACK0_p & v8e4b0e;
assign v85ce72 = RtoB_ACK0_p & v8e2373 | !RtoB_ACK0_p & v8e21d1;
assign v8e5a22 = jx2_p & v8b5793 | !jx2_p & v85dfab;
assign v8e1e6c = DEQ_p & v8b57ae | !DEQ_p & v8e591f;
assign v8e56ef = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8e1810;
assign v845187 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8672b3;
assign v8e5895 = BtoS_ACK6_p & v8568c2 | !BtoS_ACK6_p & v8565ab;
assign v844fbd = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844f91;
assign v86531f = BtoS_ACK8_p & v8b568f | !BtoS_ACK8_p & !v85c1d4;
assign v880b12 = BtoS_ACK0_p & v85aa18 | !BtoS_ACK0_p & v8b578f;
assign v85db5c = RtoB_ACK1_p & v8b57b5 | !RtoB_ACK1_p & v89954f;
assign v8b5609 = BtoS_ACK6_p & v8e5956 | !BtoS_ACK6_p & v8b5727;
assign v8b55b1 = StoB_REQ7_p & v8452dc | !StoB_REQ7_p & v8b5559;
assign v8564c4 = ENQ_p & v8572d0 | !ENQ_p & v8e4235;
assign v856275 = EMPTY_p & v8e5a5f | !EMPTY_p & v857144;
assign v86006a = BtoR_REQ0_p & v8e1862 | !BtoR_REQ0_p & v8601d6;
assign v88924e = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v85c416;
assign v8b5826 = BtoS_ACK7_p & v865862 | !BtoS_ACK7_p & !v8a5b8c;
assign v8e59e6 = RtoB_ACK0_p & v8e4aa2 | !RtoB_ACK0_p & v8e4579;
assign v867a85 = jx1_p & v8e4514 | !jx1_p & v8b5896;
assign v8e4b4d = jx1_p & v85dee1 | !jx1_p & v844f91;
assign v8568a8 = EMPTY_p & v8e5a5f | !EMPTY_p & v8b5846;
assign v8e21da = RtoB_ACK1_p & v8e519d | !RtoB_ACK1_p & v8b56d1;
assign v8af2be = BtoS_ACK7_p & v8e55ef | !BtoS_ACK7_p & v85696d;
assign v85696d = BtoS_ACK6_p & v856f89 | !BtoS_ACK6_p & v8e43dc;
assign v8b56ae = jx2_p & v8af3c9 | !jx2_p & !v844f91;
assign v85aa14 = EMPTY_p & v85f343 | !EMPTY_p & v865770;
assign v8b565b = StoB_REQ2_p & v85ea8d | !StoB_REQ2_p & !v844f91;
assign v8e436f = DEQ_p & v8e1f1b | !DEQ_p & v8e3cfe;
assign v8e473e = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & v8e5a2d;
assign v8650c5 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e5a75;
assign v85c9fb = jx1_p & v8dc673 | !jx1_p & v844f91;
assign jx1_n = !v880bc3;
assign v8e484a = jx1_p & v85dee1 | !jx1_p & !v8e4e95;
assign v85638e = jx2_p & v85ffb2 | !jx2_p & v8e4e45;
assign v882429 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v84513a;
assign v8af26f = FULL_p & v85f2b2 | !FULL_p & v8b553d;
assign v8e1aee = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e10b7;
assign v8b54dc = jx2_p & v856fbd | !jx2_p & v844f91;
assign v85688c = StoB_REQ8_p & v8e3d3c | !StoB_REQ8_p & v8b55bc;
assign v8e5650 = jx2_p & v8e46b2 | !jx2_p & v856386;
assign v85e23a = jx1_p & v85f42f | !jx1_p & v8b5841;
assign v8e1755 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5b48;
assign v856e1f = jx1_p & v86290d | !jx1_p & v8e5a9d;
assign v8e4a8a = StoB_REQ1_p & v861740 | !StoB_REQ1_p & v8be167;
assign v8b55e6 = jx2_p & v8e3f8b | !jx2_p & v85ffcd;
assign v85c93d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8af1a3;
assign v8b5641 = BtoS_ACK0_p & v85a8af | !BtoS_ACK0_p & v8e59d0;
assign v856be5 = BtoR_REQ1_p & v889ec2 | !BtoR_REQ1_p & v85726b;
assign v8e570f = jx2_p & v8b5768 | !jx2_p & v8e1d42;
assign v860551 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4637;
assign v85f814 = jx2_p & v8e39e6 | !jx2_p & v856386;
assign v85724c = jx2_p & v8563a6 | !jx2_p & v8b551c;
assign v85d886 = jx1_p & v85da8e | !jx1_p & v844f91;
assign v8a5c52 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v856bc8;
assign v8b5622 = ENQ_p & v8e1d7d | !ENQ_p & v8e4461;
assign v845373 = jx2_p & v88c2da | !jx2_p & v8e2248;
assign v8b56b6 = jx2_p & v8e2040 | !jx2_p & v8af18f;
assign v8b5842 = StoB_REQ8_p & v8e4ea5 | !StoB_REQ8_p & v8e14ea;
assign v8af0ec = BtoS_ACK2_p & v8e3883 | !BtoS_ACK2_p & v8e4e35;
assign v8a5c02 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v86e8c2;
assign v8af0dc = StoB_REQ7_p & v8af418 | !StoB_REQ7_p & v85e237;
assign v85e99d = ENQ_p & v8e4d59 | !ENQ_p & v85d8e2;
assign v845380 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e2282;
assign v8e520c = BtoS_ACK0_p & v84507a | !BtoS_ACK0_p & !v85ab77;
assign v89b438 = StoB_REQ0_p & v88c2b9 | !StoB_REQ0_p & !v844f91;
assign v8566fa = EMPTY_p & v85d543 | !EMPTY_p & v85a4f0;
assign v865b8f = stateG7_1_p & v8e4f00 | !stateG7_1_p & v85695e;
assign v84507a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8e40a9;
assign v8cce3b = jx2_p & v8e4523 | !jx2_p & v845146;
assign v899247 = jx0_p & v8e5494 | !jx0_p & v844f91;
assign v8e1eb4 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8b572f;
assign v8e4184 = jx1_p & v8e4514 | !jx1_p & v8e4050;
assign v85db04 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e5a8f;
assign v8b5880 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8a8877;
assign v8b5544 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dc552;
assign v8e4f78 = BtoR_REQ0_p & v8e1c7f | !BtoR_REQ0_p & !v856261;
assign v8e41c2 = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v8e22ae;
assign v8e4be1 = jx1_p & v883b69 | !jx1_p & v8e40df;
assign v883cf8 = StoB_REQ6_p & v8e58d2 | !StoB_REQ6_p & v844f91;
assign v8cc95b = ENQ_p & v8af46c | !ENQ_p & v856b71;
assign v8b5548 = jx1_p & v844f91 | !jx1_p & v85a8af;
assign v8b57fb = BtoS_ACK0_p & v8b5554 | !BtoS_ACK0_p & v8b5610;
assign v8e59b1 = StoB_REQ7_p & v85a8af | !StoB_REQ7_p & v8e1701;
assign v85cc2b = BtoR_REQ0_p & v8e5208 | !BtoR_REQ0_p & v8e598b;
assign v8e5a15 = jx1_p & v85c83d | !jx1_p & !v844f91;
assign v8e1956 = jx2_p & v865772 | !jx2_p & v8e41ec;
assign v85ddb7 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v85ea8d;
assign v8dc5b6 = jx2_p & v85a648 | !jx2_p & v8e4fe5;
assign v856261 = EMPTY_p & v8e3ab5 | !EMPTY_p & !v889244;
assign v8e572e = BtoS_ACK8_p & v8b5844 | !BtoS_ACK8_p & v8452da;
assign v8e5a94 = DEQ_p & v85e1a3 | !DEQ_p & v85f2b2;
assign v85aeb5 = BtoS_ACK0_p & v85dbda | !BtoS_ACK0_p & v8e48b6;
assign v8e44d0 = BtoS_ACK7_p & v8b55e6 | !BtoS_ACK7_p & !v856bd5;
assign v85ccf0 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8e3d7b;
assign v889f94 = ENQ_p & v8e4e6e | !ENQ_p & v8af19b;
assign v881ad8 = jx1_p & v8e46de | !jx1_p & !v85cc2a;
assign v88c2f2 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e5b2c;
assign v865261 = jx3_p & v8e4916 | !jx3_p & v8e4096;
assign v8bf8d3 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v88e287;
assign v8a5c49 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8991c0;
assign v89921c = jx1_p & v8e59d1 | !jx1_p & v85d2e2;
assign v8992a4 = jx0_p & v857943 | !jx0_p & !v86f9a1;
assign v8e4b2c = BtoS_ACK8_p & v85b66d | !BtoS_ACK8_p & v85e4d3;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v877314 = StoB_REQ6_p & v85b3a4 | !StoB_REQ6_p & v8e1484;
assign v8b54d4 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v85afc8;
assign v8e4918 = BtoS_ACK6_p & v85a008 | !BtoS_ACK6_p & v8e21c5;
assign v85b400 = StoB_REQ1_p & v86f9a1 | !StoB_REQ1_p & !v856eba;
assign v844fa1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f91;
assign v8b57d0 = jx0_p & v844f97 | !jx0_p & v844f91;
assign v8e428a = StoB_REQ1_p & v85db04 | !StoB_REQ1_p & v8b55dd;
assign v857309 = BtoS_ACK0_p & v8e3eb2 | !BtoS_ACK0_p & v857542;
assign v8e5a5a = EMPTY_p & v8e5a82 | !EMPTY_p & v8dc5e7;
assign v8e47ef = StoB_REQ3_p & v86e8c2 | !StoB_REQ3_p & !v844f91;
assign v8b572c = FULL_p & v85a893 | !FULL_p & v8564c4;
assign v89954f = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8b54d4;
assign v86007f = BtoS_ACK0_p & v8e4c47 | !BtoS_ACK0_p & v85f2c8;
assign v8e4294 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8e4224;
assign v8e4a30 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e428a;
assign v8b54d7 = BtoS_ACK6_p & v8af14f | !BtoS_ACK6_p & v8e59d4;
assign v8b5836 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8af268;
assign v8e5989 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v856594;
assign v8e40ce = jx2_p & v8b5601 | !jx2_p & v86d6bd;
assign v8e1a90 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e5924;
assign v8b56a2 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8af185;
assign v8af185 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8e3a10;
assign v8e15a0 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85626a;
assign v85733c = stateG12_p & v856558 | !stateG12_p & !v8e3f84;
assign v8e10fb = BtoS_ACK8_p & v85d53f | !BtoS_ACK8_p & v8af231;
assign v889ec1 = BtoS_ACK2_p & v8e16ea | !BtoS_ACK2_p & v880dfd;
assign v8b55d7 = ENQ_p & v85ba14 | !ENQ_p & v8b558c;
assign v8dc668 = EMPTY_p & v85f2b2 | !EMPTY_p & v8e18ff;
assign v8e1811 = jx1_p & v8b5630 | !jx1_p & !v8562b8;
assign v858482 = jx1_p & v8a87cd | !jx1_p & !v85f2f8;
assign v8dc6c6 = jx3_p & v86654a | !jx3_p & v8e21da;
assign v8af19b = BtoS_ACK8_p & v8b555a | !BtoS_ACK8_p & v8b55a0;
assign v865121 = jx0_p & v88c324 | !jx0_p & !v8e55c9;
assign v85abee = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85658e;
assign v85b670 = RtoB_ACK0_p & v857107 | !RtoB_ACK0_p & v88bc2b;
assign v85dcd6 = jx1_p & v8e58a0 | !jx1_p & !v844f91;
assign v8e3916 = BtoS_ACK0_p & v85dbda | !BtoS_ACK0_p & v8a5c2b;
assign v85f448 = jx2_p & v8452fa | !jx2_p & v8e15b2;
assign v8e4d7d = BtoS_ACK0_p & v86e347 | !BtoS_ACK0_p & v8cc8c9;
assign v8e3f8b = jx1_p & v8a5c45 | !jx1_p & !v85e259;
assign v8e4aa2 = BtoR_REQ1_p & v8b57bd | !BtoR_REQ1_p & !v844f91;
assign v857549 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e4bb0;
assign v8e1d1f = jx1_p & v8af14f | !jx1_p & v8e59df;
assign v8e21d3 = jx2_p & v8e5060 | !jx2_p & v85b49f;
assign v85f35f = BtoS_ACK0_p & v8e4d7b | !BtoS_ACK0_p & v8b5794;
assign v88bc4c = BtoS_ACK8_p & v8e597f | !BtoS_ACK8_p & v86b0d6;
assign v8b563f = BtoS_ACK1_p & v8e1692 | !BtoS_ACK1_p & v8e566a;
assign v8e193b = BtoS_ACK2_p & v8bf0c7 | !BtoS_ACK2_p & v856556;
assign v8e1106 = RtoB_ACK1_p & v8e4416 | !RtoB_ACK1_p & v8e4ca0;
assign v8e1c52 = StoB_REQ0_p & v8e5033 | !StoB_REQ0_p & v844f97;
assign v8be124 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8b55f8;
assign v889f5a = ENQ_p & v85ba14 | !ENQ_p & v8e3ad8;
assign v8e1f66 = BtoS_ACK0_p & v8cdce6 | !BtoS_ACK0_p & v8e4ffe;
assign v885308 = jx2_p & v8e3dad | !jx2_p & v8b552a;
assign v8e15fd = jx2_p & v85a5e3 | !jx2_p & !v8e238d;
assign v8b5501 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e3899;
assign v8cc8ae = BtoS_ACK7_p & v8e5a5e | !BtoS_ACK7_p & v8e1504;
assign v85c754 = BtoS_ACK7_p & v8e3c83 | !BtoS_ACK7_p & v845047;
assign v8b5645 = jx1_p & v85f5a7 | !jx1_p & v85d6ea;
assign v8562f2 = jx1_p & v844f91 | !jx1_p & v8e1f00;
assign v862719 = ENQ_p & v8b5607 | !ENQ_p & v8e3bee;
assign v8566be = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v8e425a;
assign v8e5977 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8e1d99;
assign v8e1b44 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e5a1c;
assign v8cc8cf = stateG7_1_p & v844f91 | !stateG7_1_p & !v8e3a68;
assign v85ae46 = DEQ_p & v8e240e | !DEQ_p & v8e3cfe;
assign v8b5601 = jx1_p & v8e5be4 | !jx1_p & v8e2267;
assign v8b5578 = BtoS_ACK8_p & v8e420a | !BtoS_ACK8_p & v8e5b23;
assign v8833ba = DEQ_p & v85a34c | !DEQ_p & v8b56c2;
assign SLC1_n = v8dc6c6;
assign v8e1654 = jx0_p & v86baf9 | !jx0_p & v8e4d0c;
assign v8845c4 = BtoR_REQ0_p & v8e3dde | !BtoR_REQ0_p & v8e4416;
assign v8e3e1e = jx0_p & v844f91 | !jx0_p & v88c324;
assign v85fc37 = EMPTY_p & v8e42f6 | !EMPTY_p & v859ffa;
assign v85c96a = jx0_p & v85b1c3 | !jx0_p & !v85abc1;
assign v85e1b8 = StoB_REQ3_p & v85ea8d | !StoB_REQ3_p & !v880dfd;
assign v8b562e = StoB_REQ2_p & v8e4224 | !StoB_REQ2_p & v8b56ec;
assign v8cc909 = BtoS_ACK0_p & v86c74d | !BtoS_ACK0_p & v85d3cc;
assign v8452da = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8e599c;
assign v85fa63 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e5244;
assign v8e1f36 = jx2_p & v881b59 | !jx2_p & !v844f91;
assign v8e5967 = RtoB_ACK1_p & v8e598e | !RtoB_ACK1_p & v85da5d;
assign v856867 = BtoS_ACK7_p & v86290d | !BtoS_ACK7_p & v85da20;
assign v8e4786 = StoB_REQ7_p & v8b5641 | !StoB_REQ7_p & v8dc68b;
assign v85eaf9 = BtoS_ACK0_p & v8e4f71 | !BtoS_ACK0_p & v85f7ea;
assign v8e3a2f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v85c6f5;
assign v8bf293 = BtoS_ACK2_p & v8e2136 | !BtoS_ACK2_p & v8e5708;
assign v8892d9 = jx1_p & v861da7 | !jx1_p & v8e1a78;
assign v86b6cf = StoB_REQ1_p & v85d671 | !StoB_REQ1_p & v85659c;
assign v8b54eb = ENQ_p & v8572d0 | !ENQ_p & v8e58ec;
assign v8e59cc = EMPTY_p & v8b56ab | !EMPTY_p & v8e522a;
assign v867c19 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8a923a;
assign v8b5758 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v856883;
assign v8569ee = jx1_p & v844f91 | !jx1_p & !v8e400a;
assign v8e22b0 = BtoS_ACK8_p & v8e2222 | !BtoS_ACK8_p & !v85f401;
assign v8e4b9f = jx1_p & v8e4514 | !jx1_p & v8b5571;
assign v8892a6 = BtoS_ACK7_p & v8618f2 | !BtoS_ACK7_p & v85cc48;
assign v8e5208 = EMPTY_p & v8e1c59 | !EMPTY_p & v8e3a16;
assign v8e222f = BtoS_ACK6_p & v8450f2 | !BtoS_ACK6_p & v85aad0;
assign v85aeed = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88d5d7;
assign v8dc617 = jx0_p & v8b5600 | !jx0_p & v8e4a95;
assign v8e1d49 = BtoS_ACK6_p & v85724c | !BtoS_ACK6_p & v8e240d;
assign v88c2da = jx1_p & v8e58ad | !jx1_p & v8e59b1;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v8e20a6 = BtoS_ACK7_p & v856f73 | !BtoS_ACK7_p & v866ae1;
assign v85b540 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v856688;
assign v85d860 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85e61d;
assign v8b556d = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85de0b;
assign v8e4be4 = ENQ_p & v8a3c77 | !ENQ_p & v8b55db;
assign v8b5640 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b54de;
assign v8b5889 = StoB_REQ6_p & v8e5982 | !StoB_REQ6_p & v8e22c7;
assign v8e4f2e = ENQ_p & v844fbf | !ENQ_p & !v8b5884;
assign v8e59ec = jx2_p & v8e57a6 | !jx2_p & v844f91;
assign v8e3992 = jx2_p & v85dcf5 | !jx2_p & !v8b5645;
assign v863949 = BtoS_ACK6_p & v85cbd3 | !BtoS_ACK6_p & v85c47a;
assign v8e1b00 = StoB_REQ6_p & v85d382 | !StoB_REQ6_p & v8691fd;
assign v8e1aa8 = stateG7_1_p & v8e59c5 | !stateG7_1_p & v845360;
assign v8e4637 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9b;
assign v85ca46 = EMPTY_p & v8e1d85 | !EMPTY_p & v85740b;
assign v8e46d9 = BtoS_ACK6_p & v85ad82 | !BtoS_ACK6_p & v8672c1;
assign v8e1f8f = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v85e694;
assign v8e5a02 = BtoS_ACK1_p & v8e52b0 | !BtoS_ACK1_p & v8a5c49;
assign v845146 = jx1_p & v8dc594 | !jx1_p & v8e3911;
assign v858462 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v85ea8d;
assign v8e519d = EMPTY_p & v8e1961 | !EMPTY_p & v8b5743;
assign v8e5a48 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88c324;
assign v8e5962 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v85ffcd;
assign v8b5813 = EMPTY_p & v8af461 | !EMPTY_p & v8e5a94;
assign v8e4cb1 = StoB_REQ0_p & v8e56dc | !StoB_REQ0_p & v8e5a80;
assign v85735b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85c895;
assign v8569c1 = BtoS_ACK1_p & v8573f7 | !BtoS_ACK1_p & v8570f0;
assign v85bbe2 = jx2_p & v8e484a | !jx2_p & v8e1811;
assign v85f411 = jx1_p & v8e5a7f | !jx1_p & v86290d;
assign v85e82e = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & v8e4605;
assign v85c971 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8e52b0;
assign v8b569c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e5b0f;
assign v88c352 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v88e4cb;
assign v8451d1 = BtoS_ACK6_p & v86d36d | !BtoS_ACK6_p & v8e444a;
assign v88c326 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4468;
assign v889fca = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v845060;
assign v8e59e5 = StoB_REQ6_p & v8af2e6 | !StoB_REQ6_p & v85e946;
assign v8e3ed3 = jx2_p & v85e355 | !jx2_p & !v844f91;
assign v8e19ae = DEQ_p & v8e5a21 | !DEQ_p & v8601d6;
assign v8b5712 = BtoS_ACK7_p & v858f70 | !BtoS_ACK7_p & v85db87;
assign v8570f0 = StoB_REQ1_p & v85f2ba | !StoB_REQ1_p & v8e415b;
assign v8a5b53 = BtoS_ACK0_p & v8e5a10 | !BtoS_ACK0_p & v8b55ab;
assign v85b642 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fb1;
assign v8e58c1 = BtoR_REQ0_p & v8b5691 | !BtoR_REQ0_p & v8b57a9;
assign v883e72 = StoB_REQ0_p & v8e39cc | !StoB_REQ0_p & v85da39;
assign v8e3dde = stateG7_1_p & v8b55a7 | !stateG7_1_p & v8893a8;
assign v8b5685 = BtoS_ACK6_p & v8b55b0 | !BtoS_ACK6_p & v8b56b6;
assign v85f5e7 = jx2_p & v8e4b4d | !jx2_p & !v85bd67;
assign v85aea7 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4a1f;
assign v85673d = BtoS_ACK0_p & v857540 | !BtoS_ACK0_p & v8be150;
assign v85768f = jx2_p & v8e1d1f | !jx2_p & v8e41ec;
assign v856f73 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85daf5;
assign v8680cc = BtoR_REQ1_p & v8e53d3 | !BtoR_REQ1_p & v8e39bb;
assign v8b5773 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & !v8451c3;
assign v844fb5 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v85eae6 = EMPTY_p & v85dc21 | !EMPTY_p & v8b574f;
assign v8e4e0e = BtoR_REQ0_p & v85d598 | !BtoR_REQ0_p & !v8e2239;
assign v85e0b0 = jx0_p & v844f9f | !jx0_p & !v8b5823;
assign v8dc594 = jx0_p & v844f9b | !jx0_p & v844f99;
assign v8b5805 = jx1_p & v8e509c | !jx1_p & v8af355;
assign v8e240d = jx2_p & v8e5a15 | !jx2_p & v86290f;
assign v899283 = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & !v8e1f7f;
assign v8e1975 = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v8b56b7;
assign v8568c2 = jx2_p & v8b5503 | !jx2_p & !v8e238d;
assign v845026 = jx2_p & v85b421 | !jx2_p & !v85cea0;
assign v8b5873 = BtoR_REQ0_p & v85e618 | !BtoR_REQ0_p & v8e413b;
assign v8b5808 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8b56e1;
assign v8b564c = EMPTY_p & v845027 | !EMPTY_p & v856f27;
assign v8e40af = jx1_p & v8e5a6a | !jx1_p & v85a8af;
assign v8b5790 = BtoS_ACK7_p & v85a894 | !BtoS_ACK7_p & !v8564bf;
assign v8e58d5 = StoB_REQ2_p & v8e3bef | !StoB_REQ2_p & v8e38a7;
assign v8e5946 = jx2_p & v85c7c5 | !jx2_p & !v85dfab;
assign v8e4d75 = jx1_p & v8b56ee | !jx1_p & v8e5bed;
assign v8569a8 = jx1_p & v8e1f02 | !jx1_p & v8e5611;
assign v8e3d36 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v8e4394;
assign v8e5c10 = RtoB_ACK1_p & v8af3c1 | !RtoB_ACK1_p & v8e5510;
assign v85ca3a = jx2_p & v85ccc4 | !jx2_p & v8e4e45;
assign v8ccdf5 = BtoS_ACK8_p & v85a98f | !BtoS_ACK8_p & v8b55fa;
assign v8b5817 = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & !v8e46e5;
assign v85b724 = jx2_p & v8e1d1f | !jx2_p & v8571db;
assign v8e46de = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v865820;
assign v8e5a35 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v856ce2;
assign v85b5fb = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8af15c;
assign v8e47b7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e82e;
assign v8b56c2 = ENQ_p & v85e45f | !ENQ_p & v8dc56c;
assign v845074 = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & !v889f82;
assign v8ce34d = BtoS_ACK0_p & v8e39c1 | !BtoS_ACK0_p & v85ce5c;
assign v8e4d0b = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v85dffb;
assign v8451b6 = BtoS_ACK0_p & v8e4637 | !BtoS_ACK0_p & v8e1667;
assign v8e118d = BtoS_ACK0_p & v8e4637 | !BtoS_ACK0_p & v8e1aee;
assign v8e46fa = BtoS_ACK7_p & v856fa4 | !BtoS_ACK7_p & !v8e4670;
assign v8e214e = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e469a;
assign v8e59c6 = jx2_p & v865810 | !jx2_p & !v870e66;
assign v8b5852 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8e1692;
assign v85e8a6 = BtoS_ACK0_p & v8b55cb | !BtoS_ACK0_p & v85dddb;
assign v8e4c64 = DEQ_p & v85e1a3 | !DEQ_p & v8b553d;
assign v8b5659 = BtoS_ACK6_p & v8e3992 | !BtoS_ACK6_p & v8af12b;
assign v866503 = BtoS_ACK7_p & v85d805 | !BtoS_ACK7_p & v85e1e9;
assign v8e5a2d = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v856951;
assign v8b55ab = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8b553e;
assign v85d917 = StoB_REQ1_p & v8b558d | !StoB_REQ1_p & v889f58;
assign v86f85b = jx0_p & v85e7d3 | !jx0_p & !v85f2cd;
assign v8e1acc = jx1_p & v8e118d | !jx1_p & v8e1bf6;
assign v8e1995 = jx1_p & v85dee1 | !jx1_p & v85ea90;
assign v8b553d = ENQ_p & v8a3c77 | !ENQ_p & v8b565e;
assign v8b57d9 = BtoS_ACK8_p & v85f334 | !BtoS_ACK8_p & v8e3ea1;
assign v8dc68b = StoB_REQ6_p & v8451c4 | !StoB_REQ6_p & v85dac7;
assign v8e3de2 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v85ea8d;
assign v85aad0 = jx2_p & v8b5624 | !jx2_p & v8b5627;
assign v85d2dd = EMPTY_p & v8b54f7 | !EMPTY_p & v8b574f;
assign v8e488c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e233b;
assign v8e3d0c = jx0_p & v8b556f | !jx0_p & !v844f99;
assign v8e56cb = StoB_REQ0_p & v8b56fd | !StoB_REQ0_p & v856a21;
assign v86c65e = jx1_p & v8b57df | !jx1_p & v844f91;
assign v85d5a0 = jx0_p & v85714b | !jx0_p & !v84507a;
assign v8e1f2b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b55c2;
assign v889f88 = jx0_p & v8b56ce | !jx0_p & v85aea7;
assign v85bdb6 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856959;
assign v8e592b = StoB_REQ8_p & v86a790 | !StoB_REQ8_p & v8e23df;
assign v8e58e9 = BtoR_REQ1_p & v867a97 | !BtoR_REQ1_p & v8893ab;
assign v8b55fa = StoB_REQ8_p & v8e41c2 | !StoB_REQ8_p & v8b57c6;
assign v8e51c8 = jx0_p & v85e80e | !jx0_p & !v8b563f;
assign v8af102 = StoB_REQ8_p & v8b572a | !StoB_REQ8_p & v8b55d2;
assign v8b577c = jx0_p & v844f9f | !jx0_p & !v8b581e;
assign v8b5827 = StoB_REQ7_p & v8e59db | !StoB_REQ7_p & v8e460d;
assign v8b5675 = BtoS_ACK1_p & v8b5600 | !BtoS_ACK1_p & v85abc2;
assign v8e1cd3 = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & v88c2b9;
assign v8e59db = BtoS_ACK0_p & v8e3eb2 | !BtoS_ACK0_p & v85acdb;
assign v8e539f = EMPTY_p & v862719 | !EMPTY_p & v8a5bcc;
assign v858ae4 = BtoS_ACK0_p & v8e1e0a | !BtoS_ACK0_p & v8e47b7;
assign v8b5724 = jx2_p & v8e4f3b | !jx2_p & v8e1650;
assign v85ea88 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v85ad35;
assign v8b56d7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85b04f;
assign v8e3a26 = BtoS_ACK8_p & v8af325 | !BtoS_ACK8_p & !v8dc58d;
assign v8e4267 = jx1_p & v8b569c | !jx1_p & v844f91;
assign v85d3e1 = BtoS_ACK6_p & v8cce3b | !BtoS_ACK6_p & v8e4191;
assign v85d59f = jx0_p & v85da91 | !jx0_p & v844f91;
assign v8e1857 = BtoS_ACK0_p & v8e5033 | !BtoS_ACK0_p & !v88d5d7;
assign v8ce3d5 = BtoS_ACK2_p & v85dbdd | !BtoS_ACK2_p & !v8e4224;
assign v8e17f5 = StoB_REQ0_p & v883ca3 | !StoB_REQ0_p & v84520b;
assign v8e5a84 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v85b938;
assign v8e3fe8 = BtoR_REQ0_p & v85c77b | !BtoR_REQ0_p & !v856261;
assign v85cde3 = BtoS_ACK6_p & v85b724 | !BtoS_ACK6_p & v8892a1;
assign v8b5559 = StoB_REQ6_p & v8452dc | !StoB_REQ6_p & v8e5769;
assign v85b238 = BtoS_ACK0_p & v8b585f | !BtoS_ACK0_p & v85e282;
assign v8e2000 = StoB_REQ0_p & v8e4c47 | !StoB_REQ0_p & v8cdce6;
assign v8e57d8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af188;
assign v8e165a = jx2_p & v8e58ac | !jx2_p & !v870e66;
assign v8af383 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e438b;
assign v85e8bf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8e531e;
assign v8587ce = jx1_p & v8451d8 | !jx1_p & !v8b55ca;
assign v8e5ace = jx2_p & v85da55 | !jx2_p & v8e2248;
assign v8e1618 = StoB_REQ7_p & v85b3a4 | !StoB_REQ7_p & v85dbd4;
assign v85b2ae = StoB_REQ0_p & v8dc594 | !StoB_REQ0_p & v8e4637;
assign v85dac7 = BtoS_ACK0_p & v8af327 | !BtoS_ACK0_p & v85f62f;
assign v8e599d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e9c5;
assign v85df05 = BtoS_ACK7_p & v8568c2 | !BtoS_ACK7_p & v8e5895;
assign v8e3c11 = jx0_p & v8e45d6 | !jx0_p & !v86066c;
assign v8e594f = ENQ_p & v844f91 | !ENQ_p & v8e1a97;
assign v86c2ed = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v856951;
assign v85b6c8 = stateG7_1_p & v8e3a68 | !stateG7_1_p & !v844f91;
assign v8e199b = StoB_REQ7_p & v8e4254 | !StoB_REQ7_p & v8e5344;
assign v856443 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85d9d4;
assign v844f91 = 1;
assign v85e340 = StoB_REQ2_p & v8af160 | !StoB_REQ2_p & !v856452;
assign v8e238d = jx1_p & v883ca3 | !jx1_p & !v844f91;
assign v844fbb = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844f91;
assign v8dc639 = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v8b576e;
assign v8cce0d = ENQ_p & v85e3a6 | !ENQ_p & v844f91;
assign v845037 = StoB_REQ5_n & v844f9f | !StoB_REQ5_n & v8af369;
assign v8e5a56 = EMPTY_p & v8e58b8 | !EMPTY_p & v8e1e6c;
assign v8b569b = ENQ_p & v8562d0 | !ENQ_p & !v8af4b7;
assign v8e5960 = BtoS_ACK0_p & v86c74d | !BtoS_ACK0_p & v8e38c7;
assign v8e4877 = jx2_p & v8e415a | !jx2_p & v8b55bf;
assign v85bd68 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e5b63;
assign v889f82 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v856452;
assign v856959 = BtoS_ACK3_p & v8e16ea | !BtoS_ACK3_p & !v8e5bd5;
assign v856474 = jx1_p & v85b073 | !jx1_p & !v845183;
assign v8967e3 = RtoB_ACK1_p & v89a257 | !RtoB_ACK1_p & !v85c6d3;
assign v8e4411 = BtoS_ACK0_p & v8e17e8 | !BtoS_ACK0_p & v8b5837;
assign v8b56a3 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v85cd1f;
assign v856f27 = DEQ_p & v8e41fc | !DEQ_p & v8b57a9;
assign v8b5776 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v866511;
assign v8e5bbe = jx0_p & v85dc0d | !jx0_p & !v85b29f;
assign v85b99e = BtoS_ACK6_p & v857374 | !BtoS_ACK6_p & v8e44d3;
assign v8e5908 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v856452;
assign v85aba0 = BtoS_ACK7_p & v8563e3 | !BtoS_ACK7_p & v8e45b5;
assign v8b5804 = DEQ_p & v8b5814 | !DEQ_p & v8e1e8f;
assign v8563a2 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8e148a;
assign v8af480 = BtoR_REQ0_p & v8e44ed | !BtoR_REQ0_p & v860057;
assign v8b5872 = BtoS_ACK0_p & v85a153 | !BtoS_ACK0_p & v85fc09;
assign v8e181b = BtoS_ACK6_p & v8b583c | !BtoS_ACK6_p & v8e59ec;
assign v86cf33 = BtoR_REQ1_p & v8e583d | !BtoR_REQ1_p & v8e202c;
assign v8dc5ab = BtoS_ACK0_p & v8e400a | !BtoS_ACK0_p & v85d376;
assign v8e44c7 = jx1_p & v8b58bb | !jx1_p & v8a691b;
assign v8e56dc = jx0_p & v88bcd0 | !jx0_p & !v844f91;
assign v8567f9 = EMPTY_p & v8e22b0 | !EMPTY_p & v8e438f;
assign v8574cc = jx0_p & v85b1c3 | !jx0_p & v844f91;
assign v845230 = jx2_p & v845245 | !jx2_p & !v8b568d;
assign BtoS_ACK3_n = !v865dba;
assign v8e4235 = jx2_p & v8569ee | !jx2_p & v844f91;
assign v8e5b68 = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & v85dee3;
assign v85e4d3 = StoB_REQ8_p & v889f0e | !StoB_REQ8_p & v8b55a3;
assign v8dc612 = StoB_REQ7_p & v8e5a9d | !StoB_REQ7_p & v85ca01;
assign v8e1692 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v85f287;
assign v8e59d0 = jx0_p & v844f91 | !jx0_p & !v85b29f;
assign v8b5850 = BtoR_REQ1_p & v8b57bd | !BtoR_REQ1_p & !v8e59f5;
assign v889f3d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e40a9;
assign v856edf = jx1_p & v8e48d7 | !jx1_p & !v844f91;
assign v8e2475 = stateG7_1_p & v8892bc | !stateG7_1_p & v8e5a56;
assign BtoS_ACK6_n = !v8893b1;
assign v856264 = jx2_p & v8e41d9 | !jx2_p & !v844f91;
assign v8e1985 = ENQ_p & v8562d0 | !ENQ_p & !v8b5892;
assign v85dffb = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v8e5a72;
assign v857139 = jx2_p & v8e19c7 | !jx2_p & !v8e4c34;
assign v8a3c77 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e5998;
assign v8e543c = BtoR_REQ1_p & v8e2239 | !BtoR_REQ1_p & !v8e4e0e;
assign v8e5936 = BtoS_ACK6_p & v8e5650 | !BtoS_ACK6_p & v8cafe0;
assign v85a893 = ENQ_p & v8572d0 | !ENQ_p & v844f91;
assign v8e4872 = EMPTY_p & v8b56c2 | !EMPTY_p & v8a5552;
assign v8b5697 = BtoS_ACK7_p & v85bdbc | !BtoS_ACK7_p & v8e590d;
assign v8e3d2a = StoB_REQ0_p & v85c96a | !StoB_REQ0_p & v8e51c8;
assign v8e1480 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85e9ee;
assign v8b5643 = jx1_p & v844f91 | !jx1_p & !v8e59f9;
assign v8e58d2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v889f88;
assign v8a5c15 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v85f8f2;
assign v8e1ea1 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8e4185;
assign v8b5627 = jx1_p & v85e152 | !jx1_p & v856d2f;
assign v8e5950 = ENQ_p & v8b55a4 | !ENQ_p & !v85ccc6;
assign v8b558a = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v857499;
assign v8a5b4f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e2136;
assign v8e1f55 = jx2_p & v8e14ab | !jx2_p & !v85f57e;
assign v8e4c46 = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & !v8b5626;
assign v85655b = BtoS_ACK0_p & v8e5033 | !BtoS_ACK0_p & v85fc09;
assign v86bbca = StoB_REQ6_p & v8e38f1 | !StoB_REQ6_p & v85e60f;
assign v85de51 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f95;
assign v8e3f79 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8e18dd;
assign v8e41db = ENQ_p & v8b5607 | !ENQ_p & v8e5242;
assign v8b554e = EMPTY_p & v885d2d | !EMPTY_p & v8e438f;
assign v8be150 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85a24b;
assign v8e228f = BtoS_ACK8_p & v8b5577 | !BtoS_ACK8_p & !v8e45a8;
assign v880b7a = jx2_p & v85d7a7 | !jx2_p & !v844f91;
assign v85d57d = BtoS_ACK6_p & v8e4f16 | !BtoS_ACK6_p & v8a5b9d;
assign v8e53d3 = stateG7_1_p & v85eae6 | !stateG7_1_p & v85dc22;
assign v8e4e95 = StoB_REQ7_p & v8e23ae | !StoB_REQ7_p & v8b55c0;
assign v8e4943 = BtoS_ACK1_p & v8e4637 | !BtoS_ACK1_p & v8af15c;
assign v8b55d8 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8e20a6;
assign v8e5985 = jx2_p & v856314 | !jx2_p & v844f91;
assign v8601d6 = ENQ_p & v844fbf | !ENQ_p & !v844f91;
assign v889ec0 = BtoS_ACK1_p & v85b938 | !BtoS_ACK1_p & v8892b6;
assign v8b57e2 = jx1_p & v8af29a | !jx1_p & v844f91;
assign v8b555f = BtoS_ACK8_p & v8e55ec | !BtoS_ACK8_p & v8e3bdc;
assign v8a5bcc = DEQ_p & v8e41db | !DEQ_p & v8e3cfe;
assign v86e347 = jx0_p & v85c632 | !jx0_p & !v856594;
assign v8b57b7 = RtoB_ACK0_p & v88934b | !RtoB_ACK0_p & v8e4187;
assign v8e5a71 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8b54e9;
assign v856bc1 = BtoS_ACK7_p & v8e5a5e | !BtoS_ACK7_p & v863949;
assign v8e1718 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e229e;
assign v8e589d = BtoS_ACK0_p & v85c9c5 | !BtoS_ACK0_p & v8b5651;
assign v8e5a98 = stateG7_1_p & v8b5563 | !stateG7_1_p & v8b5667;
assign v85de34 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v844f91;
assign v8dc55f = DEQ_p & v8b57c8 | !DEQ_p & v86c2d3;
assign v8e4c11 = jx2_p & v89921c | !jx2_p & !v8e2355;
assign v85de64 = jx0_p & v8b56ce | !jx0_p & v8e4831;
assign v860007 = StoB_REQ0_p & v8664e6 | !StoB_REQ0_p & v844f91;
assign v8e59ee = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8451a1;
assign v8e41ec = jx1_p & v8b57df | !jx1_p & v8af14f;
assign v8cce1f = jx1_p & v844f91 | !jx1_p & v8dc599;
assign v8e3bda = BtoS_ACK6_p & v8b552b | !BtoS_ACK6_p & v8e4fe5;
assign v85ea90 = StoB_REQ7_p & v8e4c47 | !StoB_REQ7_p & v8e42fe;
assign v8565e5 = jx1_p & v844f91 | !jx1_p & v8e38f1;
assign v8e5a0b = StoB_REQ7_p & v8e3a74 | !StoB_REQ7_p & v844f91;
assign v85b2bc = jx0_p & v8e4d94 | !jx0_p & v8e55c9;
assign v88c355 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4f71;
assign v8af3c9 = jx1_p & v8b56ee | !jx1_p & v85f2f8;
assign v84535e = jx1_p & v88c32e | !jx1_p & v8e40df;
assign v89920a = BtoS_ACK6_p & v85ad82 | !BtoS_ACK6_p & v8e544a;
assign v8e4dcf = StoB_REQ1_p & v85e93d | !StoB_REQ1_p & v8b5817;
assign v8e3e82 = StoB_REQ1_p & v8e3d7b | !StoB_REQ1_p & v8e52b0;
assign v8e58ef = StoB_REQ7_p & v85e652 | !StoB_REQ7_p & v85d7e9;
assign v85d3cc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b57b3;
assign v8e3b66 = StoB_REQ7_p & v8e3eb2 | !StoB_REQ7_p & v8cce20;
assign v85fa64 = StoB_REQ6_p & v8e5212 | !StoB_REQ6_p & v8e42b2;
assign v865862 = jx2_p & v85641f | !jx2_p & !v868a25;
assign v8af4c4 = jx1_p & v8e4fe5 | !jx1_p & v85b512;
assign v8dc5ff = jx2_p & v85e091 | !jx2_p & v85dfab;
assign v8e1d42 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v885341;
assign v8e5a3b = BtoS_ACK1_p & v8573f7 | !BtoS_ACK1_p & v86654f;
assign v85626a = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8b57f2;
assign v8e233b = jx0_p & v8b552d | !jx0_p & v889f3d;
assign v8e2154 = ENQ_p & v8e4e6e | !ENQ_p & v8bf437;
assign v8b54f0 = DEQ_p & v85a277 | !DEQ_p & v862911;
assign v8e509c = StoB_REQ6_p & v8572ac | !StoB_REQ6_p & v8e22c7;
assign v8e197f = StoB_REQ7_p & v8e4c47 | !StoB_REQ7_p & v8452cd;
assign v85b66d = jx2_p & v8e4b2a | !jx2_p & v86d6bd;
assign v8e5a82 = ENQ_p & v8562d0 | !ENQ_p & !v85d6fe;
assign v8e48b6 = jx0_p & v85adf5 | !jx0_p & v844f91;
assign v85ad35 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8af160;
assign v867a75 = StoB_REQ1_p & v86f9a1 | !StoB_REQ1_p & v845074;
assign v8a5b25 = jx0_p & v844f91 | !jx0_p & v86f9a1;
assign v8af3b8 = StoB_REQ8_p & v8e59d6 | !StoB_REQ8_p & v8e3a7c;
assign v8b56a6 = BtoS_ACK7_p & v856255 | !BtoS_ACK7_p & v85744d;
assign v85aa21 = jx0_p & v8e40a9 | !jx0_p & !v84507a;
assign v8e3b74 = BtoR_REQ0_p & v8b54ed | !BtoR_REQ0_p & v8e3cfe;
assign v8572ac = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8e4c9d;
assign v8e3bbb = StoB_REQ8_p & v85df05 | !StoB_REQ8_p & v8e58a1;
assign v85a0d2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85da91;
assign v85cea0 = jx1_p & v8e2470 | !jx1_p & !v8e3ae7;
assign v8e20ff = StoB_REQ1_p & v85c416 | !StoB_REQ1_p & v85e340;
assign BtoS_ACK5_n = !v88c3ad;
assign v85ff96 = EMPTY_p & v85654c | !EMPTY_p & v8e522a;
assign v85d8ae = EMPTY_p & v85bbe5 | !EMPTY_p & v8b5743;
assign v8b57ac = RtoB_ACK0_p & v8e4aa2 | !RtoB_ACK0_p & v8e3e8e;
assign v8b56ab = ENQ_p & v8af46c | !ENQ_p & v8e4668;
assign v8e5098 = jx1_p & v85dee1 | !jx1_p & !v8b5745;
assign v8b5822 = BtoR_REQ0_p & v8e5a9f | !BtoR_REQ0_p & v8b5558;
assign v8e1a8c = jx2_p & v8b57fe | !jx2_p & v856474;
assign v8b56c8 = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & !v844fb7;
assign v85dee3 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v8e2395;
assign v8e14db = jx1_p & v85dee1 | !jx1_p & !v856eca;
assign v8e583f = BtoS_ACK1_p & v8573f7 | !BtoS_ACK1_p & v88424e;
assign v8e59a9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4e2c;
assign v85e5db = ENQ_p & v8e5607 | !ENQ_p & !v844f91;
assign v8e39eb = stateG7_1_p & v85f839 | !stateG7_1_p & v856c6c;
assign v8e4337 = jx1_p & v85acf3 | !jx1_p & v85ad39;
assign v8e4f00 = EMPTY_p & v8e4be4 | !EMPTY_p & v863db8;
assign v8e2040 = jx1_p & v844f91 | !jx1_p & v85f35f;
assign v85f244 = jx0_p & v86baf9 | !jx0_p & !v8b56a8;
assign v8cc8f2 = jx0_p & v8e4a30 | !jx0_p & !v8e59d3;
assign v8e597b = StoB_REQ8_p & v8e16d2 | !StoB_REQ8_p & v856ae7;
assign v8563e3 = jx2_p & v8b5505 | !jx2_p & v86290d;
assign v856725 = EMPTY_p & v8e54de | !EMPTY_p & v8b5809;
assign v8e1b43 = BtoS_ACK0_p & v8e5a10 | !BtoS_ACK0_p & v8b572b;
assign v85fa19 = BtoS_ACK8_p & v8af325 | !BtoS_ACK8_p & v8e4189;
assign v85d7bb = StoB_REQ6_p & v8b5517 | !StoB_REQ6_p & !v8e4662;
assign v85659e = BtoS_ACK6_p & v85cb94 | !BtoS_ACK6_p & v8569c7;
assign v856479 = StoB_REQ2_p & v856598 | !StoB_REQ2_p & v85cb88;
assign v8e59bd = jx1_p & v8e416f | !jx1_p & v8e55a8;
assign v8a880e = StoB_REQ8_p & v8af4a4 | !StoB_REQ8_p & v8e5049;
assign v8e1a9b = jx2_p & v85e23a | !jx2_p & v8b54e6;
assign v85c73b = jx0_p & v8e4832 | !jx0_p & v85e7f0;
assign v85da6c = jx0_p & v85b3fb | !jx0_p & v85f2cd;
assign v85b6b7 = BtoS_ACK2_p & v857499 | !BtoS_ACK2_p & v8e40f6;
assign v8e4514 = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v8e4574;
assign v8e589a = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v856c3d;
assign v8451d8 = StoB_REQ7_p & v845249 | !StoB_REQ7_p & v863e80;
assign v8e1c87 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4d8f;
assign v8af292 = jx2_p & v8be114 | !jx2_p & !v8587ce;
assign v8b57be = StoB_REQ0_p & v8b57a5 | !StoB_REQ0_p & !v8af243;
assign v8e59f9 = BtoS_ACK0_p & v8e400a | !BtoS_ACK0_p & v85d98f;
assign v8b54f4 = jx1_p & v8e46de | !jx1_p & !v8e1c52;
assign v8e1756 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b5764;
assign v8e1c27 = jx2_p & v85a3a4 | !jx2_p & !v85dfab;
assign v8e17a8 = stateG12_p & v8b566d | !stateG12_p & !v85ccc6;
assign v856763 = StoB_REQ7_p & v8b56e5 | !StoB_REQ7_p & v8b54c0;
assign v8e4153 = StoB_REQ8_p & v8e5413 | !StoB_REQ8_p & !v844f91;
assign v8e1a74 = StoB_REQ8_p & v8e15a4 | !StoB_REQ8_p & v8e1abc;
assign v889f78 = StoB_REQ8_p & v85da27 | !StoB_REQ8_p & v86695b;
assign v8e438a = BtoS_ACK7_p & v856264 | !BtoS_ACK7_p & v8565b3;
assign v8e424e = jx2_p & v8e4f56 | !jx2_p & v85dbad;
assign v856919 = BtoS_ACK1_p & v8e4a1f | !BtoS_ACK1_p & v8b565c;
assign v8e19fe = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8e5033;
assign v8e58a0 = BtoS_ACK0_p & v8e4637 | !BtoS_ACK0_p & v882156;
assign v8e48f1 = RtoB_ACK1_p & v86cf33 | !RtoB_ACK1_p & v88bcc9;
assign v8b560e = jx1_p & v85acf3 | !jx1_p & v85b07e;
assign v8e4ed1 = RtoB_ACK1_p & v8e1c89 | !RtoB_ACK1_p & v8b5522;
assign v8b57c1 = jx1_p & v8e589b | !jx1_p & v85dee5;
assign v8b57c6 = BtoS_ACK7_p & v85638e | !BtoS_ACK7_p & v8e10c0;
assign v8dc551 = jx0_p & v85f50b | !jx0_p & v85da56;
assign v8e4142 = StoB_REQ0_p & v8e1084 | !StoB_REQ0_p & v844f91;
assign v8b576a = DEQ_p & v8e17a8 | !DEQ_p & v8e2147;
assign v87aaa9 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v8e5a35;
assign v856878 = jx2_p & v844f91 | !jx2_p & v899197;
assign v8e1969 = jx1_p & v8e1a1d | !jx1_p & v8e1598;
assign v8562d0 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v844fbd;
assign v8b56ba = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85d971;
assign v8e58f5 = BtoS_ACK7_p & v8563e3 | !BtoS_ACK7_p & v8e56a0;
assign v8b5677 = BtoS_ACK0_p & v86972a | !BtoS_ACK0_p & v889fca;
assign v8e4db6 = BtoS_ACK6_p & v85a008 | !BtoS_ACK6_p & v8e1cfb;
assign v856367 = BtoS_ACK2_p & v85725c | !BtoS_ACK2_p & v8e4270;
assign v85e08e = BtoS_ACK7_p & v8e4e4e | !BtoS_ACK7_p & v8e3977;
assign v8e1770 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85b514;
assign v8573c8 = ENQ_p & v85e3a6 | !ENQ_p & v8e55e7;
assign v8672c7 = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & v8846fb;
assign v85d6ab = StoB_REQ3_p & v8b5800 | !StoB_REQ3_p & v844f9f;
assign v85a5eb = EMPTY_p & v889f5a | !EMPTY_p & v8b574f;
assign v8b582a = BtoS_ACK8_p & v8e53a5 | !BtoS_ACK8_p & !v8b573a;
assign v8b54da = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e4b5f;
assign v85c8b5 = jx0_p & v844f91 | !jx0_p & v8b5893;
assign v8e4e81 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v8564e9;
assign v856b8e = BtoR_REQ0_p & v8cce39 | !BtoR_REQ0_p & v856364;
assign v8b55e9 = DEQ_p & v85f27b | !DEQ_p & v8b55ed;
assign v8e5a68 = BtoS_ACK0_p & v8cce79 | !BtoS_ACK0_p & !v8e479e;
assign v898498 = StoB_REQ1_p & v85df40 | !StoB_REQ1_p & v85ba1d;
assign v85e355 = jx1_p & v8cce41 | !jx1_p & v844f91;
assign v8e432e = BtoS_ACK7_p & v8e1f55 | !BtoS_ACK7_p & !v8812e9;
assign v8892c0 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e23ce;
assign v8e55ba = BtoS_ACK8_p & v85d914 | !BtoS_ACK8_p & v85a4be;
assign v8563a9 = BtoS_ACK7_p & v8e2025 | !BtoS_ACK7_p & v85cde3;
assign v8e16ce = BtoS_ACK0_p & v85699e | !BtoS_ACK0_p & !v8564e9;
assign v8b57df = StoB_REQ0_p & v8e388e | !StoB_REQ0_p & v8e3d0c;
assign v8e2416 = jx2_p & v85dcf5 | !jx2_p & !v8e4ac8;
assign v856ec1 = BtoS_ACK8_p & v8e4602 | !BtoS_ACK8_p & !v8e1b23;
assign v84518e = BtoS_ACK7_p & v8b561b | !BtoS_ACK7_p & !v845109;
assign v8e5be4 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5525;
assign v8e4baa = BtoS_ACK6_p & v8e56ac | !BtoS_ACK6_p & v8e240d;
assign v8e4b24 = BtoS_ACK0_p & v856594 | !BtoS_ACK0_p & !v8e47dd;
assign v8e4c04 = StoB_REQ1_p & v899202 | !StoB_REQ1_p & v85e000;
assign v85df70 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85fa6e;
assign v8e501a = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844fb7;
assign v8e5b11 = StoB_REQ6_p & v85b5f6 | !StoB_REQ6_p & v85677f;
assign v85b380 = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & v8e4c73;
assign v85e1a0 = jx1_p & v85ccfd | !jx1_p & v844f91;
assign v880b59 = jx2_p & v856b6d | !jx2_p & v8af213;
assign v8e5957 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5883;
assign v8e4187 = BtoR_REQ1_p & v8e5a98 | !BtoR_REQ1_p & v8892d3;
assign v8b56f8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86d019;
assign v8e45ab = ENQ_p & v8af34b | !ENQ_p & v8e3a58;
assign v85bd7c = jx2_p & v85db32 | !jx2_p & v8b54db;
assign v8e4d72 = BtoS_ACK7_p & v8e2025 | !BtoS_ACK7_p & v8cce49;
assign v8e5799 = jx0_p & v8e49d3 | !jx0_p & !v844f91;
assign v8e5b6d = jx2_p & v8e58b6 | !jx2_p & !v85e895;
assign v8e43ad = jx0_p & v844f9f | !jx0_p & !v85a0f8;
assign v8e544a = jx2_p & v8e5907 | !jx2_p & v856b8f;
assign v85cbd3 = jx2_p & v8e1e0e | !jx2_p & v85dfab;
assign v88c38a = StoB_REQ7_p & v85d382 | !StoB_REQ7_p & v8e1cc4;
assign v85fedf = BtoS_ACK1_p & v8e1eb9 | !BtoS_ACK1_p & v8e1bc1;
assign v8e565f = jx1_p & v85dee1 | !jx1_p & !v8e41a7;
assign v85db1a = BtoS_ACK0_p & v8e3979 | !BtoS_ACK0_p & v8e57a4;
assign v899fb0 = BtoS_ACK6_p & v8b5840 | !BtoS_ACK6_p & v8b5720;
assign v881aaf = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9b;
assign v8b5816 = StoB_REQ6_p & v8e1f00 | !StoB_REQ6_p & v8e159f;
assign v8e54a9 = BtoS_ACK0_p & v8e1c52 | !BtoS_ACK0_p & !v8e5754;
assign v8573f7 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v8b550c;
assign v8b564f = BtoS_ACK7_p & v88928c | !BtoS_ACK7_p & v8e3c65;
assign v8e4d32 = BtoS_ACK0_p & v8b56e6 | !BtoS_ACK0_p & v8e1c07;
assign v8b581e = BtoS_ACK1_p & v8e16ea | !BtoS_ACK1_p & v8e4d85;
assign v856fdd = EMPTY_p & v85ca37 | !EMPTY_p & v865770;
assign v856a1f = jx1_p & v8b56ee | !jx1_p & v8e4c47;
assign v85d6b7 = RtoB_ACK0_p & v856653 | !RtoB_ACK0_p & v8b5585;
assign v8e38a7 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8e417e;
assign v8e4ece = BtoS_ACK1_p & v8e3d7b | !BtoS_ACK1_p & v8e4c46;
assign v85a622 = StoB_REQ7_p & v8b5641 | !StoB_REQ7_p & v8e242d;
assign v8af14f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v86dabf;
assign v89a257 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8b57bd;
assign v883566 = jx0_p & v86baf9 | !jx0_p & v844f91;
assign v8e5a6a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85c93d;
assign v8af40a = BtoS_ACK8_p & v8b562f | !BtoS_ACK8_p & v8af102;
assign v85b07e = BtoS_ACK0_p & v85ad39 | !BtoS_ACK0_p & v8b55e1;
assign v86582f = jx2_p & v8e5906 | !jx2_p & v86290d;
assign v8b587d = StoB_REQ7_p & v85f1cb | !StoB_REQ7_p & v8e59e4;
assign v8e5a9f = stateG7_1_p & v8b5649 | !stateG7_1_p & v8e4872;
assign v8e5242 = BtoS_ACK8_p & v8b55a6 | !BtoS_ACK8_p & v85c47d;
assign v8a6915 = jx1_p & v867a93 | !jx1_p & v85d2e2;
assign v85da91 = BtoS_ACK1_p & v8e2265 | !BtoS_ACK1_p & v85e548;
assign v8e1c96 = EMPTY_p & v8e44d9 | !EMPTY_p & v8563b6;
assign v8b5630 = BtoS_ACK0_p & v85dbda | !BtoS_ACK0_p & v8e508f;
assign v8e4a57 = jx0_p & v844f91 | !jx0_p & v85da91;
assign v8562ab = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b56a0;
assign v8b573e = BtoS_ACK7_p & v86290d | !BtoS_ACK7_p & v8e1ebe;
assign v88c31b = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e4a06;
assign v8e56dd = ENQ_p & v8e4e6e | !ENQ_p & v8e4b6f;
assign v8e1abc = BtoS_ACK7_p & v85c80b | !BtoS_ACK7_p & v8e597e;
assign v8e1d85 = ENQ_p & v8af46c | !ENQ_p & v85d701;
assign v880bdf = StoB_REQ7_p & v85e0a1 | !StoB_REQ7_p & v84523b;
assign v857499 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f9f;
assign v8e5883 = StoB_REQ6_p & v8e3cb6 | !StoB_REQ6_p & v85673d;
assign v8cce52 = StoB_REQ7_p & v8e4c47 | !StoB_REQ7_p & v8e2000;
assign v85e7be = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8573b2;
assign v8e57d3 = BtoS_ACK0_p & v8e4d7b | !BtoS_ACK0_p & v8e58f9;
assign v85b0a3 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b54fc;
assign v8b55ef = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v8e4345;
assign v889e03 = BtoS_ACK2_p & v8bf0c7 | !BtoS_ACK2_p & v8e5259;
assign v8e49eb = ENQ_p & v85e45f | !ENQ_p & v88c2fb;
assign v8e5259 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856c62;
assign v8b57d3 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e5a66;
assign v85f62f = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v85705c;
assign v8e598e = EMPTY_p & v8b5798 | !EMPTY_p & v8e17ae;
assign v889f96 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e4eb5;
assign v8e42dc = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v86349c;
assign v85b49f = jx1_p & v8e59d5 | !jx1_p & v8e58ce;
assign v85697c = jx1_p & v8e3f65 | !jx1_p & v844f91;
assign v8e55a6 = BtoS_ACK7_p & v889f6d | !BtoS_ACK7_p & !v85659e;
assign v8e59e7 = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & !v8e199a;
assign v8e5a39 = StoB_REQ0_p & v8e5a9d | !StoB_REQ0_p & v899247;
assign v85eb04 = BtoS_ACK7_p & v85a894 | !BtoS_ACK7_p & !v8e45a4;
assign v8e47dd = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8af44d;
assign v8e58d7 = StoB_REQ1_p & v8e4c46 | !StoB_REQ1_p & v85679b;
assign v859ffa = DEQ_p & v8e2429 | !DEQ_p & v85f2b2;
assign v8e3dec = StoB_REQ2_p & v85ea8d | !StoB_REQ2_p & v8665a9;
assign v85dcf5 = jx1_p & v844fa3 | !jx1_p & !v85e2b5;
assign v8b584c = jx2_p & v8e565f | !jx2_p & v85b5d9;
assign v8e21b3 = stateG7_1_p & v844f91 | !stateG7_1_p & !v856725;
assign v8e3e4b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e58cc;
assign v885fa8 = BtoS_ACK0_p & v8e466b | !BtoS_ACK0_p & v8e3e3a;
assign v85d6fe = BtoS_ACK8_p & v8b5863 | !BtoS_ACK8_p & !v8b55a5;
assign v85f2f8 = jx0_p & v8e4f80 | !jx0_p & v844f9d;
assign v856b08 = StoB_REQ1_p & v85c416 | !StoB_REQ1_p & v8af160;
assign v8e56ac = jx2_p & v8563a6 | !jx2_p & v8e3e49;
assign v8e3b88 = BtoS_ACK7_p & v8b55e6 | !BtoS_ACK7_p & !v8565bb;
assign v85d7e9 = StoB_REQ6_p & v8cc909 | !StoB_REQ6_p & v8b56c3;
assign v85df2b = BtoS_ACK0_p & v8e58d6 | !BtoS_ACK0_p & !v85d2bd;
assign v85ad82 = jx2_p & v856a1f | !jx2_p & v85dfab;
assign v8564db = jx1_p & v8e469f | !jx1_p & v85df0b;
assign v85dc22 = EMPTY_p & v8e20ac | !EMPTY_p & v8b574f;
assign v8e1bc1 = StoB_REQ1_p & v88924e | !StoB_REQ1_p & v8e56d9;
assign v856afe = EMPTY_p & v8569df | !EMPTY_p & v8e58b0;
assign v8e38ea = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v8e3b4b;
assign v8451f9 = BtoS_ACK6_p & v8b55b0 | !BtoS_ACK6_p & v8e3f7f;
assign v8a555c = BtoR_REQ1_p & v8b54f9 | !BtoR_REQ1_p & v8e58c1;
assign v8e51d0 = jx1_p & v8e4574 | !jx1_p & !v844f91;
assign v8e5266 = StoB_REQ8_p & v8e57dd | !StoB_REQ8_p & v85ddc7;
assign v85f567 = StoB_REQ8_p & v8e5a61 | !StoB_REQ8_p & v8e3fca;
assign v85cd1c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8af160;
assign v856575 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87c63a;
assign v8b565c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8566f3;
assign v8af29a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8af46d;
assign v8b5897 = BtoS_ACK6_p & v8e4235 | !BtoS_ACK6_p & v8b56fb;
assign v85761b = jx1_p & v8e59f6 | !jx1_p & !v8e400a;
assign v8e42a4 = jx2_p & v85db32 | !jx2_p & v868a25;
assign v85dd64 = StoB_REQ7_p & v86290d | !StoB_REQ7_p & v865d5b;
assign v8e5889 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e1f85;
assign v8e4ba8 = BtoS_ACK8_p & v8e176c | !BtoS_ACK8_p & v85ad1a;
assign v8a5561 = BtoS_ACK1_p & v8e519b | !BtoS_ACK1_p & v867a75;
assign v8574ed = BtoS_ACK0_p & v8e388e | !BtoS_ACK0_p & v8e47f2;
assign v8e590b = BtoS_ACK0_p & v8e5048 | !BtoS_ACK0_p & v8b55e4;
assign v8e18dd = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & v844f9f;
assign v8e58cc = StoB_REQ6_p & v85dff8 | !StoB_REQ6_p & v844f91;
assign v8564f5 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v845037;
assign v8af21d = BtoS_ACK6_p & v885308 | !BtoS_ACK6_p & v8b56be;
assign v8e2288 = BtoS_ACK7_p & v85a008 | !BtoS_ACK7_p & v8e4918;
assign v84501d = FULL_p & v860057 | !FULL_p & v86c2d3;
assign v8e4996 = BtoS_ACK6_p & v85cb94 | !BtoS_ACK6_p & v8e1fa5;
assign v856902 = jx2_p & v8e1730 | !jx2_p & v8b553b;
assign v85e000 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8e519b;
assign v8b582d = BtoS_ACK8_p & v86290d | !BtoS_ACK8_p & v8e4959;
assign v85d3c7 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8e5b68;
assign v85dcb5 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856b4b;
assign v8dc5b0 = RtoB_ACK1_p & v856653 | !RtoB_ACK1_p & v85d6b7;
assign v856dbe = EMPTY_p & v8b561f | !EMPTY_p & v8e5a6e;
assign v85e272 = StoB_REQ8_p & v856466 | !StoB_REQ8_p & v8e3b2f;
assign v8e1d76 = BtoS_ACK7_p & v8e516c | !BtoS_ACK7_p & v8e3a6a;
assign v8e4461 = BtoS_ACK8_p & v8e1e59 | !BtoS_ACK8_p & v8e4d9f;
assign v8e1d7d = BtoS_ACK8_p & v8e1e59 | !BtoS_ACK8_p & !v8b55f7;
assign v8e58b3 = StoB_REQ8_p & v8b5621 | !StoB_REQ8_p & v8e2177;
assign v8984af = jx1_p & v85ccfd | !jx1_p & v85e8a6;
assign v8e46a3 = BtoS_ACK0_p & v8e17e8 | !BtoS_ACK0_p & v8b57bb;
assign v8e5a2c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5722;
assign v8e464c = jx0_p & v8e4831 | !jx0_p & v844f91;
assign v8e479e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8e59b7;
assign v845064 = StoB_REQ8_p & v8b5621 | !StoB_REQ8_p & v8e59ae;
assign v8b55ac = ENQ_p & v8b5607 | !ENQ_p & v8e1d09;
assign v8e503a = BtoS_ACK7_p & v8a5cb5 | !BtoS_ACK7_p & !v8e5959;
assign v8a5c2d = StoB_REQ7_p & v8a5bfd | !StoB_REQ7_p & v8e53be;
assign v85b2a9 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8e4f80;
assign v8b5763 = jx0_p & v8b54d3 | !jx0_p & v856919;
assign v8dc6bf = EMPTY_p & v85b9a7 | !EMPTY_p & v8e588f;
assign DEQ_n = !v8967e3;
assign v8e4416 = EMPTY_p & v856ff6 | !EMPTY_p & v8893a8;
assign v85c435 = jx0_p & v85e7ea | !jx0_p & !v8b55cb;
assign v85736b = BtoS_ACK7_p & v865862 | !BtoS_ACK7_p & !v899fb0;
assign v8dc5fb = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8af0ec;
assign v867a58 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9d;
assign v8af327 = jx0_p & v8e4c04 | !jx0_p & !v8dc5ec;
assign v8e58e6 = jx1_p & v8b563d | !jx1_p & v85a8af;
assign v85cc2a = StoB_REQ7_p & v8e5033 | !StoB_REQ7_p & v8e1c52;
assign v860057 = ENQ_p & v8562d0 | !ENQ_p & v844f91;
assign v8b568e = jx1_p & v844f91 | !jx1_p & v85727c;
assign v8565cc = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v856c55;
assign v8e18bd = StoB_REQ6_p & v8caede | !StoB_REQ6_p & v8af3cb;
assign v8b554a = EMPTY_p & v8e3f84 | !EMPTY_p & v8b5796;
assign v8e39bb = BtoR_REQ0_p & v8b5545 | !BtoR_REQ0_p & v8569df;
assign v8e58ae = DEQ_p & v85d2c4 | !DEQ_p & v8cce0d;
assign v8cce02 = BtoS_ACK2_p & v8e16ea | !BtoS_ACK2_p & v8e17e6;
assign v8e1f00 = BtoS_ACK0_p & v85a8af | !BtoS_ACK0_p & v8b56fd;
assign v8dc554 = BtoS_ACK6_p & v8b55b0 | !BtoS_ACK6_p & v8e5942;
assign v8b5884 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v85ce79;
assign v8e1f2f = BtoS_ACK1_p & v8e52f8 | !BtoS_ACK1_p & v85c4c3;
assign v8af40e = BtoS_ACK0_p & v8e3d0c | !BtoS_ACK0_p & v8b56f5;
assign v85e0a1 = BtoS_ACK0_p & v865820 | !BtoS_ACK0_p & v8e59fb;
assign v8e3fce = FULL_p & v8e3cfe | !FULL_p & v85d8ad;
assign v8e5a21 = stateG12_p & v8b5732 | !stateG12_p & !v8b55a4;
assign v8e44b5 = BtoS_ACK2_p & v8e2136 | !BtoS_ACK2_p & v899219;
assign v8e17d6 = jx2_p & v856765 | !jx2_p & v844f91;
assign v8af213 = jx1_p & v8e3916 | !jx1_p & v8e23a9;
assign v8e58c2 = jx2_p & v8e1969 | !jx2_p & v8e2248;
assign v8e1823 = BtoR_REQ0_p & v85ddb8 | !BtoR_REQ0_p & v8b567f;
assign v85f8da = BtoR_REQ1_p & v8b58b1 | !BtoR_REQ1_p & v8e197c;
assign v85ce79 = StoB_REQ8_p & v8e3dd3 | !StoB_REQ8_p & v844f91;
assign v8e1a88 = EMPTY_p & v85da46 | !EMPTY_p & v863db8;
assign v8b35e8 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8e4f80;
assign v8b5691 = stateG7_1_p & v8e59cc | !stateG7_1_p & v85ff96;
assign v8b560a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v882429;
assign v85a9b1 = jx2_p & v85c7af | !jx2_p & v8564ef;
assign v8b55dd = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e1c1c;
assign v8e5ba4 = ENQ_p & v8af46c | !ENQ_p & v8b57d9;
assign v8e570e = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & !v85e340;
assign v8e1764 = jx2_p & v8e4b4d | !jx2_p & !v85e4ac;
assign v85e9b9 = jx0_p & v87aaa9 | !jx0_p & v8e45f5;
assign v85aa18 = jx0_p & v8a87b4 | !jx0_p & v8e3d7b;
assign v856c71 = StoB_REQ7_p & v85f646 | !StoB_REQ7_p & v8b54f5;
assign v8e239b = jx0_p & v85d314 | !jx0_p & v844f91;
assign v8e425a = StoB_REQ8_p & v8e55a6 | !StoB_REQ8_p & !v844f91;
assign v85b5c5 = jx1_p & v85acf3 | !jx1_p & v8e46a3;
assign v85ccec = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85e887;
assign v8cc9b5 = jx3_p & v8e572f | !jx3_p & v8563cb;
assign v889f95 = jx0_p & v8b556d | !jx0_p & v844f91;
assign v880b6e = jx1_p & v85d8ba | !jx1_p & !v844f91;
assign v8e4d5c = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v86582c;
assign v856bd4 = DEQ_p & v85a34c | !DEQ_p & v8e5aa8;
assign v8e53b1 = StoB_REQ6_p & v8a6968 | !StoB_REQ6_p & v8e1f85;
assign v8b561f = ENQ_p & v8e3f4c | !ENQ_p & !v8b569a;
assign v8b55f2 = DEQ_p & v8e45ab | !DEQ_p & v85e99d;
assign v8842d0 = BtoS_ACK6_p & v8cce3b | !BtoS_ACK6_p & v8b55c5;
assign v8e4217 = StoB_REQ0_p & v8dc594 | !StoB_REQ0_p & v8e4f71;
assign v8e572f = RtoB_ACK1_p & v85ca46 | !RtoB_ACK1_p & v860053;
assign v85ca40 = StoB_REQ1_p & v8e1ead | !StoB_REQ1_p & v844f91;
assign v88928c = jx2_p & v8892d9 | !jx2_p & v8e436b;
assign v8af46c = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e2158;
assign v8e41c1 = jx1_p & v880bdf | !jx1_p & !v85b2d5;
assign v85b5f3 = stateG7_1_p & v8db551 | !stateG7_1_p & v8e40eb;
assign v8e3979 = jx0_p & v844f91 | !jx0_p & v8b56ce;
assign v885d2d = BtoS_ACK8_p & v8af2e0 | !BtoS_ACK8_p & !v87f6a7;
assign v8e5a01 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b55fc;
assign v8e22f8 = StoB_REQ7_p & v8e1f00 | !StoB_REQ7_p & v8b5816;
assign v870e66 = jx1_p & v8dc6a0 | !jx1_p & v8e1d73;
assign v85c73e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v85fc09;
assign v8b57b8 = jx1_p & v844f91 | !jx1_p & v8b42e8;
assign v856c2e = jx1_p & v8e3f6f | !jx1_p & v8b5538;
assign v8e4d04 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8be0f9;
assign v8b55f7 = BtoS_ACK7_p & v8e1c8a | !BtoS_ACK7_p & !v8e1e59;
assign v86658f = BtoS_ACK2_p & v8b5875 | !BtoS_ACK2_p & v889f3b;
assign v85672e = jx0_p & v8e3c39 | !jx0_p & v8e59c0;
assign v856fe9 = BtoS_ACK5_p & v8b56c8 | !BtoS_ACK5_p & v844f9f;
assign v8e4603 = jx1_p & v8e58c9 | !jx1_p & !v8e199b;
assign v861611 = BtoS_ACK8_p & v8b5696 | !BtoS_ACK8_p & !v8b5621;
assign v87ee2b = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v8568f6;
assign v8cce31 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8e59c0;
assign v856354 = jx1_p & v844f91 | !jx1_p & v85aeed;
assign v84523b = StoB_REQ6_p & v85e0a1 | !StoB_REQ6_p & v8e3b75;
assign v8b5807 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8dc59e;
assign v8b5823 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4632;
assign v85d434 = jx1_p & v8a87cd | !jx1_p & v8e4c47;
assign v8b573a = StoB_REQ8_p & v8b5790 | !StoB_REQ8_p & v8e5a2b;
assign v865d55 = StoB_REQ8_p & v866503 | !StoB_REQ8_p & !v88486d;
assign v889f0e = BtoS_ACK7_p & v85a008 | !BtoS_ACK7_p & v8e4db6;
assign v85ad8b = StoB_REQ8_p & v8e5707 | !StoB_REQ8_p & v8563a9;
assign v8af2da = jx1_p & v85dee1 | !jx1_p & !v85a1f0;
assign v856481 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8567a3;
assign v85679b = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8b5626;
assign v8b58ad = BtoS_ACK6_p & v85d805 | !BtoS_ACK6_p & v8e5b7d;
assign v8b5681 = BtoS_ACK7_p & v8a5c84 | !BtoS_ACK7_p & !v8e14e0;
assign v8b5610 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v856b4f;
assign v856799 = jx1_p & v85b4ff | !jx1_p & !v85d52e;
assign v8b563d = StoB_REQ6_p & v88c326 | !StoB_REQ6_p & v8b5806;
assign v8e59c5 = EMPTY_p & v8cc95a | !EMPTY_p & v8e5880;
assign v8b57ea = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8af18b;
assign v85d8f4 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85b2d3;
assign jx2_n = !v8b3618;
assign v8e5a75 = BtoS_ACK3_p & v8b5875 | !BtoS_ACK3_p & v85dffb;
assign v85ceaf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8451d7;
assign v8e3a36 = jx2_p & v8a54eb | !jx2_p & !v8b57c1;
assign v8e59d5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8e4142;
assign v87f6a7 = StoB_REQ8_p & v8e3972 | !StoB_REQ8_p & v8e503a;
assign v85ad39 = jx0_p & v844fa0 | !jx0_p & v85dbdd;
assign v8e3af1 = StoB_REQ0_p & v8e5033 | !StoB_REQ0_p & v84507a;
assign v8e59f0 = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v8e5778;
assign v8b5721 = jx0_p & v8b587e | !jx0_p & v8e4ece;
assign v8e50df = BtoS_ACK0_p & v8b56e6 | !BtoS_ACK0_p & v8e22fd;
assign v8e5a64 = BtoS_ACK0_p & v8b585f | !BtoS_ACK0_p & v8e1fdc;
assign v8e595d = jx2_p & v865131 | !jx2_p & v8e58b4;
assign v8b57ce = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8e593b;
assign v8b56be = jx2_p & v8e46b8 | !jx2_p & v8564db;
assign v85e951 = StoB_REQ6_p & v8e59f9 | !StoB_REQ6_p & v8dc5ab;
assign v8b5527 = BtoS_ACK8_p & v8af186 | !BtoS_ACK8_p & !v85e858;
assign v8e5606 = jx1_p & v8e596c | !jx1_p & v85dba0;
assign v8af419 = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8e20f6;
assign v845360 = EMPTY_p & v8b54eb | !EMPTY_p & v8e5880;
assign v8b5749 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v889f4f;
assign v85663a = stateG12_p & v844f91 | !stateG12_p & !v8b569a;
assign v85f53b = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8af327;
assign v8e2045 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v845351;
assign v8e55ef = jx2_p & v8b587b | !jx2_p & v844f91;
assign v856b48 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v844f91;
assign v856386 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5a2c;
assign v8b54d8 = jx0_p & v856960 | !jx0_p & v8e1c5f;
assign v866812 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v85c986;
assign v8e2158 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e4086;
assign v8991c0 = StoB_REQ2_p & v8db8b5 | !StoB_REQ2_p & v844f91;
assign v8b569f = BtoR_REQ0_p & v8b57bd | !BtoR_REQ0_p & !v8b554a;
assign v8e52a2 = BtoR_REQ1_p & v8b55a7 | !BtoR_REQ1_p & v8845c4;
assign v8e1664 = StoB_REQ0_p & v8e3979 | !StoB_REQ0_p & v85db39;
assign v85e33b = jx1_p & v8e5a64 | !jx1_p & !v8e1f85;
assign v8e56a0 = BtoS_ACK6_p & v856b36 | !BtoS_ACK6_p & v85fabb;
assign v8e3a68 = EMPTY_p & v8e594f | !EMPTY_p & v8b55d5;
assign v8be142 = BtoS_ACK0_p & v8e4637 | !BtoS_ACK0_p & v8a881f;
assign v85afea = jx1_p & v88924d | !jx1_p & !v85e237;
assign v8e59d6 = BtoS_ACK7_p & v8a5c58 | !BtoS_ACK7_p & v8572b6;
assign v85f123 = BtoS_ACK0_p & v85ad39 | !BtoS_ACK0_p & v8e1f19;
assign v8b54c4 = BtoS_ACK2_p & v8bf0c7 | !BtoS_ACK2_p & v8e1934;
assign v8b5793 = jx1_p & v8e4514 | !jx1_p & v8e477d;
assign v844fa0 = StoB_REQ5_n & v844f91 | !StoB_REQ5_n & !v844f91;
assign v8e3911 = StoB_REQ0_p & v8b57d0 | !StoB_REQ0_p & v8e5033;
assign v8892a1 = jx2_p & v856ad9 | !jx2_p & v8984af;
assign v8e3ea2 = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v8e4c41;
assign v8e5900 = EMPTY_p & v8b5887 | !EMPTY_p & v85af2b;
assign v8b566c = BtoS_ACK0_p & v85b09e | !BtoS_ACK0_p & v8984d7;
assign v856406 = jx2_p & v844f91 | !jx2_p & v8e45e3;
assign v861ed7 = BtoS_ACK6_p & v85f814 | !BtoS_ACK6_p & v8e5a5c;
assign v8b5757 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v8b550c = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v8b5875;
assign v8e522a = DEQ_p & v85654c | !DEQ_p & v8e59fd;
assign v8e4fc9 = BtoS_ACK0_p & v889f88 | !BtoS_ACK0_p & v8b56a4;
assign v87c63a = jx0_p & v85d433 | !jx0_p & !v8e5a33;
assign v85f133 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v865f86;
assign v85a10a = jx2_p & v865772 | !jx2_p & v8571db;
assign v85a3a4 = jx1_p & v8e4574 | !jx1_p & !v8b56d6;
assign v867398 = EMPTY_p & v8dc60e | !EMPTY_p & v8833ba;
assign v899550 = StoB_REQ3_p & v856fe9 | !StoB_REQ3_p & v8e18dd;
assign v8e23ce = BtoS_ACK0_p & v8cf0f4 | !BtoS_ACK0_p & v85735b;
assign v8e3a6a = BtoS_ACK6_p & v8e5ace | !BtoS_ACK6_p & v86582f;
assign v8e19b2 = stateG7_1_p & v8e4a83 | !stateG7_1_p & v8b5649;
assign v8b5500 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85ba36;
assign v85b906 = RtoB_ACK0_p & v8b54fa | !RtoB_ACK0_p & v85666e;
assign v8e2060 = StoB_REQ6_p & v8b5677 | !StoB_REQ6_p & v857558;
assign v8e19a8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5693;
assign v8a5cb3 = BtoS_ACK2_p & v85725c | !BtoS_ACK2_p & v8af330;
assign v8b551c = jx1_p & v8b5508 | !jx1_p & !v8566f1;
assign v8b574f = DEQ_p & v889f5a | !DEQ_p & v8af41e;
assign v8e1d5f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e2436;
assign v8b5672 = jx2_p & v8e14ab | !jx2_p & !v856edf;
assign v8b55a6 = jx2_p & v8e4be1 | !jx2_p & v8b55bf;
assign v8e599c = BtoS_ACK7_p & v866544 | !BtoS_ACK7_p & v8b54d7;
assign v8e4ad3 = StoB_REQ8_p & v8a8822 | !StoB_REQ8_p & v8892a6;
assign v85ccc4 = jx1_p & v844f91 | !jx1_p & !v8e5a9d;
assign v863e80 = StoB_REQ6_p & v8e559d | !StoB_REQ6_p & v8e5171;
assign v85f52f = BtoS_ACK7_p & v85de51 | !BtoS_ACK7_p & v8b5666;
assign v8451d7 = jx0_p & v8e4943 | !jx0_p & v8cce31;
assign v8b562a = jx0_p & v857549 | !jx0_p & v8b5533;
assign v8e1ec6 = BtoS_ACK8_p & v8dc5ff | !BtoS_ACK8_p & v8e5887;
assign v856fbd = jx1_p & v8e1718 | !jx1_p & !v8e400a;
assign v8e4e6e = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8b5880;
assign v8af0f7 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v86e720;
assign v8e243e = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v85ddb7;
assign v8dc5ec = StoB_REQ1_p & v86e4e7 | !StoB_REQ1_p & v8e56eb;
assign v8567a3 = StoB_REQ2_p & v8e469a | !StoB_REQ2_p & v8b57ef;
assign v8b588e = BtoS_ACK7_p & v8e594c | !BtoS_ACK7_p & !v8e5a43;
assign v85631f = jx2_p & v85f4e0 | !jx2_p & !v8e5606;
assign v865820 = jx0_p & v8e4f71 | !jx0_p & v8dc58b;
assign v867a71 = StoB_REQ1_p & v8dc67d | !StoB_REQ1_p & v85f386;
assign v8e59df = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8dc599;
assign v8e4617 = jx0_p & v844f9f | !jx0_p & v8b5857;
assign v8e5943 = BtoS_ACK7_p & v8a5c84 | !BtoS_ACK7_p & !v8842d0;
assign v8e415a = jx1_p & v8e5753 | !jx1_p & v8e40df;
assign v8b57fe = jx1_p & v8e58d8 | !jx1_p & !v8b5795;
assign v8b578f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85c73b;
assign v8672c1 = jx2_p & v8b35f5 | !jx2_p & v856a93;
assign v8af369 = StoB_REQ5_p & v844fb7 | !StoB_REQ5_p & !v844f91;
assign v8b5698 = BtoS_ACK1_p & v8e213d | !BtoS_ACK1_p & v8847b9;
assign v8a54eb = jx1_p & v8a87cd | !jx1_p & !v8e1841;
assign v8a5552 = DEQ_p & v8b56c2 | !DEQ_p & v8e5aa8;
assign v8e4071 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8b574d;
assign v85ae84 = stateG7_1_p & v85c6f0 | !stateG7_1_p & v8db551;
assign v8b54fa = BtoR_REQ0_p & v8e539f | !BtoR_REQ0_p & v85dcb9;
assign v8e5171 = BtoS_ACK0_p & v8e4831 | !BtoS_ACK0_p & v85ceaf;
assign v8b54c7 = StoB_REQ0_p & v85f2f8 | !StoB_REQ0_p & v85e4fc;
assign v856ca7 = jx2_p & v8e21d0 | !jx2_p & v8e4e45;
assign v8e1c72 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5501;
assign v8e4f80 = StoB_REQ5_n & v844f9f | !StoB_REQ5_n & !v844f91;
assign v8563b6 = DEQ_p & v8e45ab | !DEQ_p & v8e591f;
assign v8e202c = EMPTY_p & v85d812 | !EMPTY_p & v856b8b;
assign v856653 = EMPTY_p & v8e4805 | !EMPTY_p & v8af457;
assign v85f2f0 = BtoS_ACK8_p & v8e3ed3 | !BtoS_ACK8_p & v85bd37;
assign v870cce = StoB_REQ7_p & v8567bb | !StoB_REQ7_p & v8b577d;
assign v8b569a = BtoS_ACK8_p & v86290d | !BtoS_ACK8_p & v86ed0b;
assign v8e1933 = jx2_p & v85b9de | !jx2_p & v885341;
assign v8e5896 = jx2_p & v8e5a59 | !jx2_p & v8e1ffd;
assign v8e4c41 = StoB_REQ2_p & v845268 | !StoB_REQ2_p & v8dc593;
assign v856c90 = BtoS_ACK7_p & v8b56f7 | !BtoS_ACK7_p & v8b5546;
assign v85d3cb = StoB_REQ7_p & v85dee5 | !StoB_REQ7_p & v85ffcd;
assign v88c2b9 = jx0_p & v8b5757 | !jx0_p & !v844f91;
assign v8dc673 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b569c;
assign v864971 = BtoS_ACK6_p & v85737f | !BtoS_ACK6_p & v85fc4e;
assign v85aaed = BtoS_ACK8_p & v85df15 | !BtoS_ACK8_p & v8e4ad3;
assign v856c3c = jx2_p & v85f43b | !jx2_p & !v8e19c3;
assign v85d90a = jx0_p & v844f9f | !jx0_p & !v8b5852;
assign v8cc8b1 = BtoS_ACK8_p & v8af325 | !BtoS_ACK8_p & v8e20d0;
assign v85a51c = BtoS_ACK1_p & v899202 | !BtoS_ACK1_p & v8dc67d;
assign v8831e7 = jx1_p & v8e1c72 | !jx1_p & v8e1765;
assign v844fb1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v889f6d = jx2_p & v8a54eb | !jx2_p & !v8b553b;
assign v8569ce = jx1_p & v85f4ff | !jx1_p & v8e1d5f;
assign v8b552a = jx1_p & v8af1e3 | !jx1_p & !v8e4589;
assign v8b58b2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5889;
assign v8b5649 = EMPTY_p & v856ba0 | !EMPTY_p & v8a5552;
assign v8af402 = jx1_p & v85da38 | !jx1_p & v8e2267;
assign v8e5a19 = EMPTY_p & v8af2f2 | !EMPTY_p & v8e3d66;
assign v8563e4 = BtoS_ACK7_p & v86c874 | !BtoS_ACK7_p & v8e222f;
assign v8e5708 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85ddb7;
assign v85653c = jx1_p & v844f91 | !jx1_p & !v8e5033;
assign v8e589c = BtoR_REQ1_p & v881b42 | !BtoR_REQ1_p & v85f12d;
assign v8e3e8e = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8e392a;
assign v88d5d7 = jx0_p & v8b5757 | !jx0_p & v844f91;
assign v8b5508 = StoB_REQ7_p & v85b5f6 | !StoB_REQ7_p & v85677f;
assign v856801 = jx1_p & v8e3c81 | !jx1_p & !v8e5298;
assign v899261 = BtoR_REQ1_p & v85d598 | !BtoR_REQ1_p & !v8e2239;
assign v86290f = jx1_p & v844f91 | !jx1_p & !v844f91;
assign v845101 = EMPTY_p & v85ce6f | !EMPTY_p & v85a4f0;
assign v8e591c = BtoR_REQ1_p & v8e5a19 | !BtoR_REQ1_p & v8af480;
assign v8e3c8e = DEQ_p & v856ec1 | !DEQ_p & !v844f91;
assign v8e19c4 = jx1_p & v8e501b | !jx1_p & v844f91;
assign v8e3f7f = jx2_p & v8b5518 | !jx2_p & v8e5a1f;
assign v8b42e6 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8b5699;
assign v85f386 = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v85d9cc;
assign v8b5515 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85c7b4;
assign v8e5048 = jx0_p & v844f9b | !jx0_p & !v889f3d;
assign v8e549e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8e5861;
assign v8e4764 = jx2_p & v844f91 | !jx2_p & !v8e16f6;
assign v8e58f9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dc5d5;
assign v8e2265 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v857499;
assign v8b55e8 = jx0_p & v8b5686 | !jx0_p & !v8e1f74;
assign v8af330 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e1f8f;
assign v8e5b8b = stateG7_1_p & v845101 | !stateG7_1_p & v85dfaa;
assign v85d971 = BtoS_ACK2_p & v8e16ea | !BtoS_ACK2_p & v8e1f76;
assign v85660c = BtoS_ACK0_p & v8e4f71 | !BtoS_ACK0_p & v84515d;
assign v8e4e25 = BtoS_ACK6_p & v8af325 | !BtoS_ACK6_p & v8b5615;
assign v8e5433 = jx2_p & v8e1bf9 | !jx2_p & !v85cea0;
assign v8e520d = StoB_REQ8_p & v88bcc8 | !StoB_REQ8_p & v8563e4;
assign v8e3ab5 = ENQ_p & v8a5b9b | !ENQ_p & v8e38c8;
assign v8af18f = jx1_p & v8af40e | !jx1_p & v844f91;
assign v8b57a5 = jx0_p & v844f91 | !jx0_p & v844f97;
assign v8e4800 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v881aaf;
assign v8cc8e8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v86f9a1;
assign v8e3a7c = BtoS_ACK7_p & v85d3d0 | !BtoS_ACK7_p & v8e21a2;
assign v8e5600 = StoB_REQ0_p & v85c96a | !StoB_REQ0_p & v8b54d1;
assign v8573b2 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v8af160;
assign v8565a3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844f95;
assign v8b54e6 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88d6ad;
assign v885f57 = BtoS_ACK0_p & v8e5a1c | !BtoS_ACK0_p & v85f133;
assign v864a5d = RtoB_ACK1_p & v8e455f | !RtoB_ACK1_p & v85b670;
assign v8b5875 = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & v844f9d;
assign v85e7ea = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v8e2451;
assign v8e212b = BtoS_ACK7_p & v8e5a5e | !BtoS_ACK7_p & v8b5847;
assign v881da6 = BtoS_ACK0_p & v8b5722 | !BtoS_ACK0_p & v85a0d2;
assign v8a6968 = BtoS_ACK0_p & v889f3d | !BtoS_ACK0_p & v8e47b7;
assign v85fc5a = jx0_p & v85f689 | !jx0_p & v867a75;
assign v8e2381 = jx0_p & v844f9f | !jx0_p & v844f9d;
assign v8dc555 = jx0_p & v86c57a | !jx0_p & v8e5569;
assign v8e18fe = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b586a;
assign v8e1ead = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v8b5543;
assign v8e49ee = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v85c632;
assign v8e4ca6 = jx1_p & v85680b | !jx1_p & v8e59b1;
assign v8ccdf7 = BtoS_ACK1_p & v8e52f8 | !BtoS_ACK1_p & v856f22;
assign v8e593b = jx0_p & v8e59ca | !jx0_p & !v844f91;
assign v8e46e5 = StoB_REQ2_p & v8af389 | !StoB_REQ2_p & !v8e2395;
assign v8b5851 = jx1_p & v889f73 | !jx1_p & !v844f91;
assign v8e1eb3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b5776;
assign v8b57f5 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v8e4637;
assign v8e4ea5 = BtoS_ACK7_p & v8e420a | !BtoS_ACK7_p & v85e545;
assign v8e3df8 = jx0_p & v85b6b5 | !jx0_p & v844f91;
assign v845189 = StoB_REQ7_p & v8e1d94 | !StoB_REQ7_p & v85ea86;
assign v85dc95 = BtoS_ACK7_p & v8b55b0 | !BtoS_ACK7_p & v8451f9;
assign v88c2fb = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & v8e41c2;
assign v8e5c69 = StoB_REQ0_p & v8564b7 | !StoB_REQ0_p & v865121;
assign v85695e = EMPTY_p & v85696e | !EMPTY_p & v863db8;
assign v8562b6 = jx1_p & v8574ed | !jx1_p & v844f91;
assign v8caede = BtoS_ACK0_p & v8568a1 | !BtoS_ACK0_p & v8e4cb1;
assign v8e3db0 = jx1_p & v8b56ee | !jx1_p & !v8e4a68;
assign v8e16d2 = BtoS_ACK7_p & v8e3bf7 | !BtoS_ACK7_p & v8e1088;
assign v8e441a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85c718;
assign v856eb9 = jx1_p & v8e38b1 | !jx1_p & v856345;
assign v8e3d83 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85a05d;
assign v8e5a09 = jx0_p & v85fedf | !jx0_p & v8a5561;
assign v8b5796 = DEQ_p & v844f91 | !DEQ_p & !v85733c;
assign v85e0e3 = BtoS_ACK0_p & v8e3eb2 | !BtoS_ACK0_p & v8e4617;
assign v880b9c = jx1_p & v86c2ed | !jx1_p & v8e59b1;
assign v85f3b1 = ENQ_p & v844fbf | !ENQ_p & !v8566be;
assign v8e3e49 = jx1_p & v8af1e3 | !jx1_p & !v8566f1;
assign v86d36d = jx2_p & v8e58cd | !jx2_p & !v8cb249;
assign v8e5897 = jx1_p & v85dee1 | !jx1_p & !v8e5212;
assign v85d42c = BtoS_ACK8_p & v8b582b | !BtoS_ACK8_p & v8e1964;
assign v8b5579 = stateG12_p & v8601d6 | !stateG12_p & !v844f91;
assign v88e4cb = jx2_p & v8e482a | !jx2_p & v8e1ffd;
assign v85da27 = BtoS_ACK7_p & v8e17d6 | !BtoS_ACK7_p & v85e4bb;
assign v8e192f = BtoS_ACK2_p & v8b5875 | !BtoS_ACK2_p & v8e1f43;
assign v8b5848 = EMPTY_p & v8b5732 | !EMPTY_p & v8a552d;
assign v8af277 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v8e1ead;
assign v8e409a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8992a4;
assign v8b56ed = StoB_REQ0_p & v8e56dc | !StoB_REQ0_p & v8e19e8;
assign v85b9a7 = ENQ_p & v844fbf | !ENQ_p & !v8e4236;
assign v856b6d = jx1_p & v85dee1 | !jx1_p & !v8e23ae;
assign v8e4976 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8a554b;
assign v857558 = BtoS_ACK0_p & v8dc617 | !BtoS_ACK0_p & v8e441a;
assign v85f343 = ENQ_p & v85e3a6 | !ENQ_p & v8e3cda;
assign v8e21d1 = BtoR_REQ1_p & v8e19b2 | !BtoR_REQ1_p & v8b5822;
assign v85dbef = BtoS_ACK0_p & v85dbda | !BtoS_ACK0_p & v8b584a;
assign v8e4003 = BtoS_ACK1_p & v85e000 | !BtoS_ACK1_p & v89925a;
assign v8b54d3 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v85cdc5;
assign v8e5350 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v881aaf;
assign v8852fd = jx1_p & v870cce | !jx1_p & v864623;
assign v85dbd4 = StoB_REQ6_p & v85b3a4 | !StoB_REQ6_p & v8e3e0e;
assign v8e38b1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5806;
assign v85fbec = BtoS_ACK7_p & v8a87fd | !BtoS_ACK7_p & v8dc571;
assign v8b55c6 = jx2_p & v85708d | !jx2_p & !v85e4af;
assign v85db87 = BtoS_ACK6_p & v85f814 | !BtoS_ACK6_p & v8e229f;
assign v8e4e35 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85dffb;
assign v8e56e1 = RtoB_ACK1_p & v85fc37 | !RtoB_ACK1_p & v8e1f59;
assign v8b56f5 = StoB_REQ0_p & v8a5b25 | !StoB_REQ0_p & v8e3c73;
assign v8e3dcc = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8e19fd;
assign v8b57da = BtoS_ACK0_p & v86290d | !BtoS_ACK0_p & v85fc09;
assign v8e45f1 = BtoS_ACK6_p & v8e5433 | !BtoS_ACK6_p & v8a5b9d;
assign v8e3c73 = jx0_p & v85fb40 | !jx0_p & v86f9a1;
assign v85f223 = StoB_REQ1_p & v88924e | !StoB_REQ1_p & v8e570e;
assign v8b55e1 = jx0_p & v85ad10 | !jx0_p & v8e19b1;
assign v8b5545 = stateG7_1_p & v85d2dd | !stateG7_1_p & v85a5eb;
assign v8e58ec = BtoS_ACK8_p & v8b54dc | !BtoS_ACK8_p & v8e5a11;
assign v8b5565 = EMPTY_p & v8b5527 | !EMPTY_p & v8af36d;
assign v86baf9 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v85a6a9;
assign v8a5c04 = RtoB_ACK1_p & v8b554e | !RtoB_ACK1_p & v856819;
assign v845351 = jx0_p & v8564de | !jx0_p & v85e548;
assign v8b56cf = jx2_p & v8e1542 | !jx2_p & v856799;
assign v8b55a3 = BtoS_ACK7_p & v880b8e | !BtoS_ACK7_p & v8e19b0;
assign v8b57b2 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v857625;
assign v8e1504 = BtoS_ACK6_p & v8e4f37 | !BtoS_ACK6_p & v8450f8;
assign v8e4885 = StoB_REQ1_p & v8e407e | !StoB_REQ1_p & v86ae81;
assign v8a554b = BtoS_ACK0_p & v8b56ce | !BtoS_ACK0_p & v8562ab;
assign v85da2e = jx0_p & v844f9f | !jx0_p & v883cc4;
assign v85d671 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e3f79;
assign v85f287 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v8e16ea;
assign v85dd9f = StoB_REQ1_p & v88924e | !StoB_REQ1_p & v8573b2;
assign v88173a = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & v8e592f;
assign v8e44a1 = BtoS_ACK6_p & v864f49 | !BtoS_ACK6_p & v8e1a90;
assign v85f689 = BtoS_ACK1_p & v8e1eb9 | !BtoS_ACK1_p & !v8e20ff;
assign v8b588b = StoB_REQ1_p & v8e19f0 | !StoB_REQ1_p & v844f91;
assign v85ca8a = RtoB_ACK1_p & v8e5900 | !RtoB_ACK1_p & v845235;
assign v899224 = jx2_p & v8e2079 | !jx2_p & v856edf;
assign v8e5c47 = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v85adaf;
assign v85dbe7 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8984a8;
assign v8e5a6f = StoB_REQ8_p & v8b5605 | !StoB_REQ8_p & v8e212b;
assign v8b57c8 = ENQ_p & v8562d0 | !ENQ_p & !v86531f;
assign v8b56ff = FULL_p & v8b55ed | !FULL_p & v85e0c2;
assign v85dda8 = BtoS_ACK0_p & v8a87ae | !BtoS_ACK0_p & !v8b5750;
assign v8b5800 = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & v844fb7;
assign v85f646 = BtoS_ACK0_p & v8e3d0c | !BtoS_ACK0_p & v8e179a;
assign v85ba99 = BtoS_ACK0_p & v85d90a | !BtoS_ACK0_p & v8e1638;
assign v8e188a = jx1_p & v8e4d32 | !jx1_p & v85655b;
assign v845222 = jx1_p & v8a87cd | !jx1_p & !v85ad39;
assign v86d6bd = jx1_p & v88c355 | !jx1_p & !v8e1c52;
assign v8b568d = StoB_REQ7_p & v85e5cf | !StoB_REQ7_p & v844f91;
assign v8af41c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e9b9;
assign v8892a8 = BtoS_ACK8_p & v8e4792 | !BtoS_ACK8_p & v8b5801;
assign v85cb89 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v885f57;
assign v885455 = jx0_p & v8b5757 | !jx0_p & !v856594;
assign v85c5cf = jx2_p & v8e19c2 | !jx2_p & !v8b5829;
assign v85cd1f = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v865125;
assign v8b580b = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v8b573f;
assign v8b56a0 = jx0_p & v85f647 | !jx0_p & v8b54e8;
assign v8e5646 = jx1_p & v8e473e | !jx1_p & v86290d;
assign v845245 = jx1_p & v85d8ba | !jx1_p & !v8e5a0b;
assign v856eca = StoB_REQ7_p & v8e5a9d | !StoB_REQ7_p & v8e5a39;
assign v8be0ec = StoB_REQ6_p & v8e19fe | !StoB_REQ6_p & v85daf5;
assign v85bbb6 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e4224;
assign v8892cb = StoB_REQ8_p & v85737f | !StoB_REQ8_p & v8e58b7;
assign v8b5626 = StoB_REQ2_p & v85ea8d | !StoB_REQ2_p & v8e4caf;
assign v8e22bd = StoB_REQ1_p & v8e1eb4 | !StoB_REQ1_p & v856cb3;
assign v8e5b0d = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85b540;
assign v8e5698 = EMPTY_p & v8dc606 | !EMPTY_p & v8e5880;
assign v8cce41 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e53e7;
assign v8e15a4 = BtoS_ACK7_p & v8e1a5a | !BtoS_ACK7_p & v8b57e0;
assign v8451a1 = StoB_REQ6_p & v84530b | !StoB_REQ6_p & v86dabf;
assign v8e5769 = BtoS_ACK0_p & v85d90a | !BtoS_ACK0_p & v8e1bf5;
assign v8af432 = EMPTY_p & v8b566b | !EMPTY_p & v85dcb8;
assign v8be147 = BtoS_ACK0_p & v85dd89 | !BtoS_ACK0_p & v8e488c;
assign v85a4fc = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e56eb;
assign v8b55c1 = BtoS_ACK0_p & v865820 | !BtoS_ACK0_p & v856575;
assign v8e3b2b = jx1_p & v8563df | !jx1_p & v8e5949;
assign v866544 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v86dabf;
assign v8991aa = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b555e;
assign v8b55b0 = jx2_p & v8cce1f | !jx2_p & v86c65e;
assign v85dfab = jx1_p & v8b56e6 | !jx1_p & v85de53;
assign v8e10f9 = jx2_p & v856b6d | !jx2_p & v8e1811;
assign v8e1f0d = BtoR_REQ0_p & v8b5813 | !BtoR_REQ0_p & v8573cf;
assign v8e14ca = DEQ_p & v8e56dd | !DEQ_p & v8b56ff;
assign v8b577f = StoB_REQ2_p & v8e4224 | !StoB_REQ2_p & !v844f91;
assign v8b5892 = BtoS_ACK8_p & v8b5863 | !BtoS_ACK8_p & !v8e58b3;
assign v8e5a5c = jx2_p & v8be0ea | !jx2_p & v844f91;
assign v8e5965 = StoB_REQ3_p & v8e4f80 | !StoB_REQ3_p & v844f91;
assign v8893a8 = ENQ_p & v8e3a26 | !ENQ_p & v85fa19;
assign v8e4255 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8e1c12;
assign v8e14ea = BtoS_ACK7_p & v8b54f2 | !BtoS_ACK7_p & v8e45f1;
assign v8e19fd = StoB_REQ1_p & v8e1e8c | !StoB_REQ1_p & !v85ea88;
assign v8b555e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844fa1;
assign v85649c = BtoS_ACK0_p & v86c74d | !BtoS_ACK0_p & v8b5836;
assign v8e18e6 = BtoS_ACK7_p & v8a5c84 | !BtoS_ACK7_p & !v85d3e1;
assign v8b567f = EMPTY_p & v85ffb3 | !EMPTY_p & v8b5846;
assign v85db08 = jx2_p & v8831e7 | !jx2_p & v8565fe;
assign v88bbf7 = jx1_p & v844f91 | !jx1_p & !v8e1857;
assign v85f218 = jx1_p & v85df5a | !jx1_p & v8e51d9;
assign v8af31b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b5543;
assign v8e2248 = jx1_p & v870cce | !jx1_p & v8b57d1;
assign v8a87f0 = BtoS_ACK0_p & v84520b | !BtoS_ACK0_p & v85df7f;
assign v8892b6 = StoB_REQ1_p & v8e1d99 | !StoB_REQ1_p & v8cce02;
assign v8e3a67 = EMPTY_p & v8b5732 | !EMPTY_p & v8e19ae;
assign v8b5542 = jx1_p & v844f91 | !jx1_p & v8b5641;
assign v8e5069 = BtoS_ACK6_p & v857139 | !BtoS_ACK6_p & v8a5b9d;
assign v8e5979 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5721;
assign v85654c = ENQ_p & v8af46c | !ENQ_p & v8af0dd;
assign v8b5814 = ENQ_p & v85e3a6 | !ENQ_p & v8e1852;
assign v8bf0c7 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v844f91;
assign v85f2a6 = ENQ_p & v8e4e6e | !ENQ_p & v85c436;
assign v8b5684 = BtoS_ACK7_p & v8e1933 | !BtoS_ACK7_p & v88c352;
assign v8e10c3 = jx2_p & v8e1995 | !jx2_p & v85dfab;
assign v866511 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8e57a1;
assign v8967e2 = jx0_p & v85e7d3 | !jx0_p & !v85aab4;
assign v844f9d = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v844f91;
assign v8b58b3 = BtoS_ACK0_p & v8e4913 | !BtoS_ACK0_p & v8e51ad;
assign v8b57e3 = BtoS_ACK2_p & v8b5875 | !BtoS_ACK2_p & !v8e5a72;
assign v85bbe5 = BtoS_ACK8_p & v8e1a8c | !BtoS_ACK8_p & !v8b56e0;
assign v8e392a = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8cc8cf;
assign v8e3af6 = jx0_p & v844f91 | !jx0_p & !v86d0c6;
assign v8b5719 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b57ea;
assign v8e2144 = StoB_REQ8_p & v8e5a61 | !StoB_REQ8_p & v8e3926;
assign v8e3b4b = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v8e5a78;
assign v85e66e = jx1_p & v844f91 | !jx1_p & v8e4040;
assign v8b57a8 = jx2_p & v880b9c | !jx2_p & v8852fd;
assign v8e57c2 = BtoS_ACK8_p & v8b5820 | !BtoS_ACK8_p & v85665c;
assign v860037 = jx2_p & v8e58cd | !jx2_p & !v8e4c34;
assign v8e4fa6 = StoB_REQ6_p & v8e198d | !StoB_REQ6_p & v85e5cf;
assign v889f58 = BtoS_ACK2_p & v8e16ea | !BtoS_ACK2_p & v863b40;
assign v8e438b = BtoS_ACK0_p & v8b5722 | !BtoS_ACK0_p & v8e2045;
assign v8e5569 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v856e07;
assign v8e4ca0 = RtoB_ACK0_p & v8e5372 | !RtoB_ACK0_p & v8e52a2;
assign v8dc606 = ENQ_p & v8572d0 | !ENQ_p & v85f427;
assign v85da46 = ENQ_p & v8a3c77 | !ENQ_p & v8892a8;
assign v85e237 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v85e0b0;
assign v8af47b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v86f9a1;
assign v8e200b = StoB_REQ0_p & v8574cc | !StoB_REQ0_p & v8e152b;
assign v85e7f0 = BtoS_ACK1_p & v8e3d7b | !BtoS_ACK1_p & v8e59e7;
assign v85ce6f = BtoS_ACK8_p & v8e4e15 | !BtoS_ACK8_p & v8b57f9;
assign v8563be = jx2_p & v8e20e3 | !jx2_p & v844f91;
assign v8e1be3 = StoB_REQ6_p & v85e259 | !StoB_REQ6_p & v8e42c6;
assign v8e5b6b = StoB_REQ0_p & v8e39c1 | !StoB_REQ0_p & v8e233b;
assign v8e17c4 = jx1_p & v86cb45 | !jx1_p & v85cb89;
assign v8e5bd2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8a5c45;
assign v8e1ed4 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8b56a2;
assign v8e44d9 = ENQ_p & v8af34b | !ENQ_p & v85d533;
assign v8b557e = jx0_p & v844f9f | !jx0_p & !v85a4fc;
assign v8e516c = jx2_p & v856813 | !jx2_p & v86290d;
assign v8db551 = EMPTY_p & v8e57c2 | !EMPTY_p & v899fe9;
assign v8b578b = jx2_p & v8562f2 | !jx2_p & v844f91;
assign v8e595c = StoB_REQ1_p & v8e44b5 | !StoB_REQ1_p & v844f91;
assign v8af190 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & !v88d5d7;
assign v8e4aec = jx2_p & v8b5542 | !jx2_p & v844f91;
assign v8e5924 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8e4b24;
assign v856f89 = jx2_p & v8e511b | !jx2_p & v8b552b;
assign v865827 = StoB_REQ0_p & v84523d | !StoB_REQ0_p & v8b5893;
assign v8e4270 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e5692;
assign v8e5c2a = BtoS_ACK0_p & v85d90a | !BtoS_ACK0_p & v8e5600;
assign v8e4cfc = jx2_p & v856663 | !jx2_p & v8e53c6;
assign v86b0d6 = StoB_REQ8_p & v85ba47 | !StoB_REQ8_p & v8b5697;
assign v8e469f = StoB_REQ7_p & v8e1199 | !StoB_REQ7_p & v8b56fe;
assign v8840fd = StoB_REQ1_p & v8e40a9 | !StoB_REQ1_p & v844f91;
assign v8e3e83 = EMPTY_p & v85e68a | !EMPTY_p & v8b55f2;
assign v8e59c7 = BtoS_ACK0_p & v8af418 | !BtoS_ACK0_p & v8e43ad;
assign v85ba2f = BtoS_ACK1_p & v8e52b0 | !BtoS_ACK1_p & v85f3fb;
assign v8e5a3c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v85ffcd;
assign v85c6d3 = RtoB_ACK0_p & v8b5850 | !RtoB_ACK0_p & !v844f91;
assign v8e43fa = jx1_p & v8e4514 | !jx1_p & v8b55b1;
assign v8af37f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e589d;
assign v8b5644 = StoB_REQ2_p & v8e469a | !StoB_REQ2_p & v856cd5;
assign v8e1c07 = jx0_p & v856dc8 | !jx0_p & !v86bf1f;
assign v883ca1 = jx0_p & v85d45f | !jx0_p & v844f91;
assign v8575ef = BtoS_ACK0_p & v85f59b | !BtoS_ACK0_p & v8e4f28;
assign v883cc4 = BtoS_ACK1_p & v8b5875 | !BtoS_ACK1_p & v86658f;
assign v85e3a6 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e58fd;
assign v8e4fe5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b56d7;
assign v8b556f = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v8e413b = EMPTY_p & v85b6e3 | !EMPTY_p & v856b8b;
assign v8e15cb = stateG12_p & v8e1d85 | !stateG12_p & v85d701;
assign v85aa15 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e5a72;
assign v8cc8ad = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5719;
assign v8b5530 = jx1_p & v8e5bd2 | !jx1_p & v844f91;
assign v8e4670 = BtoS_ACK6_p & v845373 | !BtoS_ACK6_p & v8e5723;
assign v8e51ad = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8e5799;
assign v8e3ac5 = StoB_REQ0_p & v85c8b5 | !StoB_REQ0_p & !v8e1810;
assign v856809 = BtoS_ACK1_p & v8e52b0 | !BtoS_ACK1_p & v8e597a;
assign v845268 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v867a58;
assign v8e3eb2 = jx0_p & v844f9f | !jx0_p & v8b5875;
assign v8e10ed = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v881a3e;
assign v85eb45 = BtoS_ACK2_p & v8e2136 | !BtoS_ACK2_p & v8b54da;
assign v8e1c89 = EMPTY_p & v8658a0 | !EMPTY_p & v8b54cb;
assign v8e4574 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v86290d;
assign v8e4c34 = jx1_p & v8e3c25 | !jx1_p & !v8e3ae7;
assign v8e3fca = BtoS_ACK7_p & v85d3d0 | !BtoS_ACK7_p & v8e1d49;
assign v8e1730 = jx1_p & v86290d | !jx1_p & v8e1841;
assign v8e199a = StoB_REQ2_p & v8e4224 | !StoB_REQ2_p & !v8574d0;
assign v8e598d = StoB_REQ0_p & v86290d | !StoB_REQ0_p & !v844f91;
assign v8e5413 = BtoS_ACK7_p & v8e3a36 | !BtoS_ACK7_p & !v8e5a60;
assign v856901 = EMPTY_p & v8b5682 | !EMPTY_p & v8e4c64;
assign v8e396e = BtoS_ACK0_p & v8b56e6 | !BtoS_ACK0_p & v8e1654;
assign v8a9208 = jx0_p & v8e4637 | !jx0_p & v8b57f5;
assign v8b589d = StoB_REQ0_p & v85db90 | !StoB_REQ0_p & v8e4d0d;
assign v8b5743 = DEQ_p & v85dd7f | !DEQ_p & v86290f;
assign v87d771 = jx2_p & v8e4eef | !jx2_p & v8b567a;
assign v8e5b16 = EMPTY_p & v8e4f2e | !EMPTY_p & v8e588f;
assign v8e1f7e = StoB_REQ6_p & v8e4050 | !StoB_REQ6_p & v8e5c2a;
assign v8dc59e = StoB_REQ1_p & v8e193b | !StoB_REQ1_p & v8e4bb0;
assign v856d2f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v86e551;
assign v8e5949 = BtoS_ACK0_p & v8af190 | !BtoS_ACK0_p & v8b56e1;
assign v8e4d0c = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v86f9a1;
assign v8e5907 = jx1_p & v8e4514 | !jx1_p & v85d382;
assign v85c986 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8db8b5;
assign v88424e = StoB_REQ1_p & v8e4c46 | !StoB_REQ1_p & v8e5173;
assign v86b9f0 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v88c2d2;
assign v857578 = StoB_REQ2_p & v857010 | !StoB_REQ2_p & v8b5754;
assign v8b56e1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v88d5d7;
assign v8e1f73 = BtoS_ACK7_p & v8e5946 | !BtoS_ACK7_p & !v85f594;
assign v86d1ff = BtoS_ACK1_p & v8e52f8 | !BtoS_ACK1_p & v8e4885;
assign v8e5952 = BtoS_ACK2_p & v856b48 | !BtoS_ACK2_p & v8e3d7b;
assign v8e160f = StoB_REQ2_p & v8db8b5 | !StoB_REQ2_p & v8b54c1;
assign v8db83f = StoB_REQ7_p & v86290d | !StoB_REQ7_p & v86299d;
assign v857037 = StoB_REQ1_p & v8e5b0d | !StoB_REQ1_p & v856be2;
assign v8e4172 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88c2e1;
assign v8b5775 = BtoS_ACK7_p & v85d3d0 | !BtoS_ACK7_p & v85b6c9;
assign v8b57d1 = StoB_REQ7_p & v8e1d94 | !StoB_REQ7_p & v8e3bf3;
assign v8e3ec6 = jx1_p & v8b56ee | !jx1_p & v85ea90;
assign v8e436c = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v857010;
assign v8e47f9 = StoB_REQ7_p & v857309 | !StoB_REQ7_p & v844f91;
assign v85f422 = BtoS_ACK0_p & v8e400a | !BtoS_ACK0_p & v85db90;
assign v88bcc9 = RtoB_ACK0_p & v8b5873 | !RtoB_ACK0_p & v8680cc;
assign v8b54d9 = BtoS_ACK1_p & v8b5875 | !BtoS_ACK1_p & v8b57e3;
assign v86ed0b = StoB_REQ8_p & v86290d | !StoB_REQ8_p & !v844f91;
assign v8e1fe7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8564e9;
assign v85b2d3 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8a5c02;
assign v85e7d3 = BtoS_ACK1_p & v85e000 | !BtoS_ACK1_p & v86653e;
assign v85df25 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v845268;
assign v8b553c = jx0_p & v844f9f | !jx0_p & !v8e201e;
assign v8565ab = jx2_p & v8e3917 | !jx2_p & !v8e484f;
assign v870b4c = jx2_p & v8e58ac | !jx2_p & !v85ffcd;
assign v8af186 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e5a3c;
assign v856951 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8b5669;
assign v8e2059 = BtoS_ACK8_p & v8b5577 | !BtoS_ACK8_p & !v8e5943;
assign v8e4a6c = jx1_p & v8af40e | !jx1_p & v85c120;
assign v85c6ec = StoB_REQ6_p & v8e3a2f | !StoB_REQ6_p & v8b5687;
assign v8e22de = StoB_REQ1_p & v866812 | !StoB_REQ1_p & v8b577b;
assign v8b3615 = jx0_p & v8e4212 | !jx0_p & v85b5db;
assign v8e576d = BtoS_ACK3_p & v8e16ea | !BtoS_ACK3_p & !v85e1b8;
assign v857625 = StoB_REQ5_n & v867a58 | !StoB_REQ5_n & !v85ea8d;
assign v8b56d6 = StoB_REQ6_p & v8e4c47 | !StoB_REQ6_p & v8e42fe;
assign v85b5bc = jx1_p & v8e57d8 | !jx1_p & !v8a5c2d;
assign v856960 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v8b55ef;
assign v8e5486 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a5bd1;
assign v8e19f0 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e519b;
assign v8a87d6 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v856b08;
assign v85e1e9 = BtoS_ACK6_p & v85d805 | !BtoS_ACK6_p & v8b5860;
assign v85ca37 = ENQ_p & v85e3a6 | !ENQ_p & v85d42c;
assign v85cdc5 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v84507b;
assign v85b6c9 = BtoS_ACK6_p & v84507d | !BtoS_ACK6_p & v8e240d;
assign v858f70 = jx2_p & v85cccf | !jx2_p & v844f91;
assign v8e55cf = jx1_p & v8451b6 | !jx1_p & !v844f91;
assign v8e4f0c = BtoS_ACK7_p & v880b8e | !BtoS_ACK7_p & v8e58b1;
assign v8b5567 = BtoS_ACK1_p & v8e1692 | !BtoS_ACK1_p & v856705;
assign v8b577b = BtoS_ACK2_p & v85f287 | !BtoS_ACK2_p & v85e111;
assign v8b582b = jx2_p & v85767f | !jx2_p & v8e1d42;
assign v8b5760 = ENQ_p & v844fbf | !ENQ_p & !v8e3d36;
assign v8dc6a0 = StoB_REQ7_p & v8b5812 | !StoB_REQ7_p & v85ffcd;
assign v8e465f = BtoS_ACK7_p & v8b54f2 | !BtoS_ACK7_p & v8e5069;
assign v8e5a60 = BtoS_ACK6_p & v8e4131 | !BtoS_ACK6_p & v8e59d8;
assign v889fea = jx3_p & v8e56e1 | !jx3_p & v85dbf1;
assign v85a008 = jx2_p & v844f91 | !jx2_p & v85653c;
assign v866ae1 = BtoS_ACK6_p & v85d3e9 | !BtoS_ACK6_p & v86cb45;
assign v8e54e0 = jx2_p & v88c39f | !jx2_p & v8a747c;
assign v8e5753 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af46d;
assign v8e3972 = BtoS_ACK7_p & v85df78 | !BtoS_ACK7_p & !v8a5bca;
assign v8e5a55 = BtoS_ACK3_p & v8e16ea | !BtoS_ACK3_p & v85e694;
assign v8e4236 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e4f0b;
assign v8b54db = jx1_p & v883ca3 | !jx1_p & v8e5033;
assign v88e277 = EMPTY_p & v845027 | !EMPTY_p & v8e5a08;
assign v85dcee = EMPTY_p & v85f48a | !EMPTY_p & v8a5bcc;
assign v88934d = DEQ_p & v8b571f | !DEQ_p & v8b57a9;
assign v85f49e = StoB_REQ8_p & v8b5662 | !StoB_REQ8_p & v8dc5be;
assign v88bc2b = BtoR_REQ1_p & v8e5208 | !BtoR_REQ1_p & v85cc2b;
assign v8b54c5 = BtoS_ACK8_p & v85e565 | !BtoS_ACK8_p & v8e1a74;
assign v8af493 = StoB_REQ8_p & v8e4235 | !StoB_REQ8_p & v8e57e7;
assign v8e388e = jx0_p & v844f91 | !jx0_p & !v844f99;
assign v8e4059 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8e44eb;
assign v85dcb8 = DEQ_p & v8e59a8 | !DEQ_p & v85a893;
assign v86349c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e4f40;
assign v8e1cfb = jx2_p & v844f91 | !jx2_p & v88bbf7;
assign v8e5a33 = StoB_REQ1_p & v86f9a1 | !StoB_REQ1_p & !v844f91;
assign v85696e = ENQ_p & v8a3c77 | !ENQ_p & v8b57fa;
assign v8e3ae7 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85fc4d;
assign v8b587a = jx2_p & v8e1730 | !jx2_p & v8b57c1;
assign v8e56eb = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e16ea;
assign v8b54d6 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8e4d0b;
assign v8e59f5 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v8b57bd;
assign v8e519b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9f;
assign v87c649 = jx3_p & v85a990 | !jx3_p & v8b5622;
assign v8b5887 = ENQ_p & v844fbf | !ENQ_p & !v85d73d;
assign v8e59d1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5517;
assign v867a97 = EMPTY_p & v8b5814 | !EMPTY_p & v8b5804;
assign v8af1e3 = StoB_REQ7_p & v8e4217 | !StoB_REQ7_p & v85b2ae;
assign v8b550b = jx1_p & v85acf3 | !jx1_p & v8e4411;
assign v85e9ee = BtoS_ACK3_p & v8e16ea | !BtoS_ACK3_p & v8e5692;
assign v85af2b = DEQ_p & v85f3b1 | !DEQ_p & v8601d6;
assign v889f4f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8ce34d;
assign v8e548f = StoB_REQ0_p & v85a8af | !StoB_REQ0_p & v8e5913;
assign v8b5701 = BtoS_ACK6_p & v8e5962 | !BtoS_ACK6_p & v8e1f02;
assign v8e3f84 = ENQ_p & v865764 | !ENQ_p & v844f91;
assign v8b5696 = jx2_p & v85dd7c | !jx2_p & !v844f91;
assign v8b586b = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v8e57c9;
assign v8e4f40 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e519b;
assign v8b5736 = BtoS_ACK6_p & v8845b3 | !BtoS_ACK6_p & v85ba35;
assign v8b576f = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8db8b5;
assign v85668b = stateG7_1_p & v8e1778 | !stateG7_1_p & v8b54ed;
assign v8b56bd = StoB_REQ5_p & v844fb7 | !StoB_REQ5_p & v85ea8d;
assign v85ddb8 = EMPTY_p & v85ffb3 | !EMPTY_p & v857144;
assign v85705c = jx0_p & v8e4003 | !jx0_p & !v889f6b;
assign v856ba0 = ENQ_p & v85e45f | !ENQ_p & v8672c7;
assign v8af12b = jx2_p & v880b6e | !jx2_p & !v844f91;
assign v8e1c84 = jx2_p & v8e484a | !jx2_p & v8af213;
assign v85ad92 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4d5c;
assign v859ffb = jx0_p & v85acfd | !jx0_p & !v844f91;
assign v88c324 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v8b54e8;
assign v8e198d = BtoS_ACK0_p & v8e4831 | !BtoS_ACK0_p & v856eb7;
assign v8e58b4 = jx1_p & v8e396e | !jx1_p & !v85e8fd;
assign v8b5722 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e2265;
assign v8e59b9 = BtoS_ACK6_p & v85faba | !BtoS_ACK6_p & v8b55ea;
assign v8b5611 = EMPTY_p & v8dc60e | !EMPTY_p & v856bd4;
assign v8e58aa = jx1_p & v8b576c | !jx1_p & !v845183;
assign v8e1e6a = StoB_REQ1_p & v8b556f | !StoB_REQ1_p & v844f9b;
assign v85d314 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v8b57de = StoB_REQ0_p & v8e59d0 | !StoB_REQ0_p & v8e5bbe;
assign v8e5930 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b42e8;
assign v8b5667 = EMPTY_p & v85f2f0 | !EMPTY_p & v8b54f0;
assign v86d72e = jx0_p & v857943 | !jx0_p & !v85b400;
assign v8b572d = StoB_REQ7_p & v8e1f00 | !StoB_REQ7_p & v8e5a27;
assign v865897 = jx2_p & v8b57cc | !jx2_p & v856386;
assign v8b5784 = jx1_p & v8e1f02 | !jx1_p & v8af0f7;
assign v856a2e = BtoS_ACK6_p & v8b55b0 | !BtoS_ACK6_p & v856fe8;
assign v8a5c22 = jx2_p & v8566b6 | !jx2_p & !v8b57ec;
assign v8e4cae = BtoS_ACK6_p & v8af325 | !BtoS_ACK6_p & v8e1764;
assign v856312 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8e501a;
assign v8af3f2 = BtoS_ACK0_p & v889f88 | !BtoS_ACK0_p & v8e1f2b;
assign v8e58cb = StoB_REQ0_p & v89920d | !StoB_REQ0_p & !v85c435;
assign v8e3ca1 = jx2_p & v8a5bf8 | !jx2_p & v8e16f6;
assign v865d5b = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8e4913;
assign v85ccdf = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85bdac;
assign v86c874 = jx2_p & v8e58e6 | !jx2_p & v8e436b;
assign v85680b = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v8e4636;
assign v8e3a58 = BtoS_ACK8_p & v8e5a22 | !BtoS_ACK8_p & v8b5648;
assign v8b5859 = jx2_p & v85b5bc | !jx2_p & v8e57d8;
assign v85f427 = BtoS_ACK8_p & v8cce37 | !BtoS_ACK8_p & v8b579c;
assign v8e57ab = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e15b2;
assign v85a4be = StoB_REQ8_p & v8e44f7 | !StoB_REQ8_p & v8b564f;
assign v8e21a2 = BtoS_ACK6_p & v8e5252 | !BtoS_ACK6_p & v8e240d;
assign v8e4e9e = BtoS_ACK6_p & v8e4e0b | !BtoS_ACK6_p & v85f3dd;
assign v85e93d = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8af389;
assign v8e41a7 = StoB_REQ7_p & v8e23ae | !StoB_REQ7_p & v8e1893;
assign v88926c = jx0_p & v85da91 | !jx0_p & v8b5722;
assign v8e109f = BtoS_ACK8_p & v8e57ab | !BtoS_ACK8_p & v8e3eb5;
assign v8e5678 = StoB_REQ6_p & v8e4217 | !StoB_REQ6_p & v85b2ae;
assign v8451c4 = BtoS_ACK0_p & v8e5a10 | !BtoS_ACK0_p & v857615;
assign v8e58a6 = jx1_p & v85dee1 | !jx1_p & !v85ad62;
assign v8e3bef = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v85c4b8;
assign v8562ad = jx0_p & v844f91 | !jx0_p & !v84507a;
assign v8e242d = StoB_REQ6_p & v8b5641 | !StoB_REQ6_p & v8af147;
assign v85dd8c = jx1_p & v85eaf9 | !jx1_p & v8e56ca;
assign v85c771 = StoB_REQ0_p & v85f2f8 | !StoB_REQ0_p & v8e5aa4;
assign v8e3d4a = BtoS_ACK8_p & v8b582b | !BtoS_ACK8_p & v889f78;
assign v8e23c6 = jx1_p & v8e57ab | !jx1_p & !v8af0dc;
assign v8e4050 = BtoS_ACK0_p & v8e4c47 | !BtoS_ACK0_p & v85c96a;
assign v8a8822 = BtoS_ACK7_p & v85a008 | !BtoS_ACK7_p & v86bc13;
assign v85bdac = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e39c1;
assign v8e44a9 = ENQ_p & v8af34b | !ENQ_p & v87356b;
assign v8e57ee = StoB_REQ6_p & v880b52 | !StoB_REQ6_p & v85afbc;
assign v861ca6 = RtoB_ACK1_p & v88c2c2 | !RtoB_ACK1_p & v85cdde;
assign v89929e = jx1_p & v8b5630 | !jx1_p & v844f91;
assign v8e4761 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v856443;
assign v8e1a1d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e588e;
assign v8e531e = StoB_REQ0_p & v8991c9 | !StoB_REQ0_p & v844f91;
assign v8b58bb = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e436b;
assign v8e51cf = jx0_p & v844f9f | !jx0_p & !v860064;
assign jx3_n = !v87c649;
assign v883d05 = jx3_p & v8e52f2 | !jx3_p & v86f694;
assign v8e474f = StoB_REQ1_p & v856e07 | !StoB_REQ1_p & !v844f91;
assign v8e1c8a = jx2_p & v8a5bf8 | !jx2_p & !v844f91;
assign v8cce8a = jx3_p & v8e5967 | !jx3_p & v8b5613;
assign v85d53f = jx2_p & v8e23c6 | !jx2_p & v8e57ab;
assign v8b5595 = StoB_REQ6_p & v8e1a2e | !StoB_REQ6_p & v8e44c8;
assign v8e4e02 = jx2_p & v8b35f0 | !jx2_p & v8562b6;
assign v86ce9d = BtoS_ACK0_p & v865827 | !BtoS_ACK0_p & v8e56ef;
assign v8af4b7 = BtoS_ACK8_p & v8af12b | !BtoS_ACK8_p & !v85e1fe;
assign v8e16ea = StoB_REQ5_p & v844f9d | !StoB_REQ5_p & v844f91;
assign v856913 = DEQ_p & v8b5579 | !DEQ_p & !v8b585b;
assign v8dc5d5 = jx0_p & v8e1b02 | !jx0_p & v85d792;
assign v85643a = StoB_REQ8_p & v889f0e | !StoB_REQ8_p & v8b55cf;
assign v856558 = ENQ_p & v8b554b | !ENQ_p & v8b56e8;
assign v8e46b8 = jx1_p & v8b560a | !jx1_p & !v8b587d;
assign v8564b7 = jx0_p & v844f91 | !jx0_p & !v8e55c9;
assign v85d2e8 = jx1_p & v8e58cf | !jx1_p & !v8e1931;
assign v85f4e0 = jx1_p & v85d8ba | !jx1_p & !v85f816;
assign v8cafe0 = jx2_p & v85ace0 | !jx2_p & v8e57d8;
assign v8b5846 = DEQ_p & v8e2154 | !DEQ_p & v85e0c2;
assign v8dc56c = BtoS_ACK8_p & v856ca7 | !BtoS_ACK8_p & v8b56b3;
assign v8b579c = StoB_REQ8_p & v8e4235 | !StoB_REQ8_p & v8e595b;
assign v8a881f = StoB_REQ0_p & v8991c9 | !StoB_REQ0_p & v8e4eba;
assign v85c6f0 = EMPTY_p & v8b56b2 | !EMPTY_p & v899fe9;
assign v8bf8d8 = jx1_p & v8b5879 | !jx1_p & v844f91;
assign v8e552e = StoB_REQ7_p & v8e3eb2 | !StoB_REQ7_p & v8e4051;
assign v8e20ac = ENQ_p & v85ba14 | !ENQ_p & v85d507;
assign v8e4497 = DEQ_p & v8e1bda | !DEQ_p & v8cce0d;
assign v8e4eba = jx0_p & v86c57a | !jx0_p & v8a5c52;
assign v8e4b9b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8e1a9b;
assign v8e5372 = EMPTY_p & v8e5a07 | !EMPTY_p & v8893a8;
assign v8e1c1c = StoB_REQ2_p & v8e5a8f | !StoB_REQ2_p & v8b5883;
assign v8e597a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8b565b;
assign v8a5b9b = BtoS_ACK8_p & v86290d | !BtoS_ACK8_p & v8e463e;
assign v85a0bf = StoB_REQ1_p & v85a05d | !StoB_REQ1_p & v85cc56;
assign v85db90 = jx0_p & v8e4d94 | !jx0_p & !v844f91;
assign v8569df = ENQ_p & v85ba14 | !ENQ_p & v844f91;
assign v8b57ab = BtoS_ACK6_p & v8e4f36 | !BtoS_ACK6_p & v8dc5b6;
assign v8e59a8 = stateG12_p & v8b566b | !stateG12_p & v8e109f;
assign v8e55c9 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8e4294;
assign v856813 = jx1_p & v87ee2b | !jx1_p & v86290d;
assign v85641f = jx1_p & v844f91 | !jx1_p & !v8e5bed;
assign v85fb40 = BtoS_ACK1_p & v8b556f | !BtoS_ACK1_p & !v85c416;
assign v8e1f43 = BtoS_ACK3_p & v8b5875 | !BtoS_ACK3_p & !v8e5a72;
assign v85b512 = StoB_REQ7_p & v8e38f1 | !StoB_REQ7_p & v86bbca;
assign v8e44ed = stateG7_1_p & v8e5a19 | !stateG7_1_p & v85d3b1;
assign v84515d = StoB_REQ0_p & v8e1084 | !StoB_REQ0_p & v85df70;
assign v8e4f56 = jx1_p & v85acf3 | !jx1_p & v85f123;
assign v856cac = jx2_p & v8e40af | !jx2_p & v844f91;
assign v8b555a = jx2_p & v8e1b05 | !jx2_p & v844f91;
assign v8e1b05 = jx1_p & v8e5939 | !jx1_p & v85a8af;
assign v8be114 = jx1_p & v8e1f02 | !jx1_p & v8b564d;
assign v8e59fb = StoB_REQ0_p & v8a54f3 | !StoB_REQ0_p & v87c63a;
assign v8e58f8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85d757;
assign v8b565d = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8967e2;
assign v8b54ec = DEQ_p & v8af1a0 | !DEQ_p & v862911;
assign v8b55e4 = StoB_REQ0_p & v8e56dc | !StoB_REQ0_p & v8e164c;
assign v8e1e8f = FULL_p & v8cce0d | !FULL_p & v8b5814;
assign v8e5a7f = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & !v85c6ec;
assign v85e942 = StoB_REQ0_p & v8a54f3 | !StoB_REQ0_p & v8992a4;
assign v8e400a = jx0_p & v844f9f | !jx0_p & !v844f91;
assign v8b550e = BtoS_ACK7_p & v8b54f2 | !BtoS_ACK7_p & v85d57d;
assign v8a8877 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8e1eb3;
assign v85a0f3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af271;
assign v856c62 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8bf0c7;
assign v8b585f = jx0_p & v844f9b | !jx0_p & !v8e40a9;
assign v8e3ff2 = StoB_REQ3_p & v856688 | !StoB_REQ3_p & !v844f9f;
assign v85f12d = EMPTY_p & v8e5ba4 | !EMPTY_p & v8e5a08;
assign v8bf339 = jx2_p & v8e1813 | !jx2_p & v8b5851;
assign v8e1fdc = StoB_REQ0_p & v8e57b4 | !StoB_REQ0_p & v8b55a2;
assign v8e3d40 = jx0_p & v8e4003 | !jx0_p & !v8e1f2f;
assign v8e599e = jx2_p & v8e4b4d | !jx2_p & !v8e4a14;
assign v86c74d = jx0_p & v8af226 | !jx0_p & v8e5971;
assign v85767e = ENQ_p & v8e4d59 | !ENQ_p & v85d533;
assign v8b54f7 = ENQ_p & v85ba14 | !ENQ_p & v8e38cd;
assign v8892c1 = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v85b979;
assign v8e3a0e = StoB_REQ1_p & v86f9a1 | !StoB_REQ1_p & !v8e1e8c;
assign v8b57fc = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85e8a6;
assign v856895 = StoB_REQ0_p & v8e39cc | !StoB_REQ0_p & v8e4bdc;
assign v845060 = jx0_p & v85b3fb | !jx0_p & v85aab4;
assign v8e585b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5757;
assign v85714b = BtoS_ACK1_p & v8e40a9 | !BtoS_ACK1_p & !v856edd;
assign v8e4a68 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85aa18;
assign v85ace0 = jx1_p & v8e57d8 | !jx1_p & !v8e2091;
assign v85ba36 = StoB_REQ1_p & v8b55ef | !StoB_REQ1_p & v844f91;
assign v8e51cd = BtoS_ACK1_p & v8e3d7b | !BtoS_ACK1_p & v8e4dcf;
assign v8b56a4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5763;
assign v8a5bbf = BtoS_ACK0_p & v8e4913 | !BtoS_ACK0_p & v8b57ce;
assign v889f6b = BtoS_ACK1_p & v8e56eb | !BtoS_ACK1_p & v85d917;
assign v85ccc2 = jx0_p & v844f9f | !jx0_p & v8b5516;
assign v8e48d8 = StoB_REQ8_p & v86290d | !StoB_REQ8_p & v8b56a6;
assign v8e508f = jx0_p & v856dc8 | !jx0_p & v844f91;
assign v8e5973 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v8b57d3;
assign v8e5426 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e5965;
assign v8e2136 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9d;
assign v8af0de = jx2_p & v8b57b8 | !jx2_p & !v8e5903;
assign v8e501b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85c8f2;
assign v8af418 = jx0_p & v844f9f | !jx0_p & !v8e16ea;
assign v8e3e3a = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & v85714b;
assign v8e57f0 = BtoS_ACK6_p & v85ad82 | !BtoS_ACK6_p & v8e38c3;
assign v8e1701 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v8e5a10;
assign v8b55d1 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b55e7;
assign v8e5a69 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e20a2;
assign v85d9d4 = BtoS_ACK0_p & v8e40a5 | !BtoS_ACK0_p & v85a0d2;
assign v85a51b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e40f6;
assign v85f816 = StoB_REQ7_p & v85e0e3 | !StoB_REQ7_p & v844f91;
assign v8e5a78 = jx2_p & v8af2da | !jx2_p & v8e1811;
assign v8e1a2e = BtoS_ACK0_p & v85e0b0 | !BtoS_ACK0_p & v8e10ed;
assign v8568a1 = jx0_p & v8e1e6a | !jx0_p & !v88475f;
assign v8e499d = jx2_p & v8e1800 | !jx2_p & v85ffcd;
assign v856eba = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v85cd1c;
assign v8af461 = ENQ_p & v8a3c77 | !ENQ_p & v8b555f;
assign v8e1d80 = EMPTY_p & v8b57ae | !EMPTY_p & v8e1e6c;
assign v8e42b2 = BtoS_ACK0_p & v8e5a9d | !BtoS_ACK0_p & v8e200b;
assign v8e572b = BtoS_ACK7_p & v85ca3a | !BtoS_ACK7_p & v8b5761;
assign v8984d7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v85c435;
assign v85cdc8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v845074;
assign v8b5621 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v8b5696;
assign v8a5bf8 = jx1_p & v86290d | !jx1_p & !v844f91;
assign v8e4e0b = jx2_p & v8a6915 | !jx2_p & !v870e66;
assign v85ab00 = BtoR_REQ1_p & v8565a2 | !BtoR_REQ1_p & v85aa14;
assign v8e438d = StoB_REQ8_p & v85eb04 | !StoB_REQ8_p & v8e44d0;
assign v8b56fa = BtoS_ACK2_p & v8e5965 | !BtoS_ACK2_p & v88c32b;
assign v8e5a73 = StoB_REQ7_p & v8a87cd | !StoB_REQ7_p & v8e59f0;
assign v86bf1f = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v8b586a;
assign v8b55ca = StoB_REQ7_p & v8e1fe7 | !StoB_REQ7_p & !v8e4fa6;
assign v8e570a = StoB_REQ1_p & v85eb45 | !StoB_REQ1_p & v844f91;
assign v8e1d32 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e4588;
assign v88c2be = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b56f8;
assign v8892d3 = stateG7_1_p & v8b5667 | !stateG7_1_p & v85d35a;
assign v8e3d7b = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v856b48;
assign v8e3a74 = BtoS_ACK0_p & v8e3eb2 | !BtoS_ACK0_p & v85da2e;
assign v8b575f = jx0_p & v8e4831 | !jx0_p & v8e1a00;
assign v85acdb = jx0_p & v857549 | !jx0_p & v8b54d9;
assign v8e583d = EMPTY_p & v85d812 | !EMPTY_p & v8e5625;
assign v881bc6 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b58ab;
assign v8e3d91 = jx2_p & v8b5530 | !jx2_p & !v844f91;
assign v8af3e3 = RtoB_ACK0_p & v85b06b | !RtoB_ACK0_p & v8b5858;
assign v8e4c29 = jx2_p & v8e2079 | !jx2_p & v85f57e;
assign v8e4b6f = BtoS_ACK8_p & v856cac | !BtoS_ACK8_p & v8892cb;
assign v8584f3 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e5973;
assign v8e4d7b = jx0_p & v899202 | !jx0_p & v8e52b0;
assign v85fc19 = StoB_REQ0_p & v8e57b4 | !StoB_REQ0_p & v85e566;
assign v8b566d = ENQ_p & v865764 | !ENQ_p & v8b582d;
assign v8e47d6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85d860;
assign v85c77b = EMPTY_p & v8e5950 | !EMPTY_p & v8b576a;
assign v85f59c = ENQ_p & v8af46c | !ENQ_p & v85aaed;
assign v862911 = jx2_p & v844f91 | !jx2_p & !v844f91;
assign v85e81e = stateG12_p & v844f91 | !stateG12_p & !v86290d;
assign v868a25 = jx1_p & v8e59be | !jx1_p & v8e5033;
assign v856656 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e1d5c;
assign v8b3618 = jx3_p & v844f91 | !jx3_p & !v8e1106;
assign v8e4a83 = EMPTY_p & v8567d9 | !EMPTY_p & v8a5552;
assign v8b58b7 = BtoS_ACK0_p & v86290d | !BtoS_ACK0_p & v88c2b9;
assign v8e3cda = BtoS_ACK8_p & v8e570f | !BtoS_ACK8_p & v8e59c9;
assign v85acf3 = StoB_REQ7_p & v8e4574 | !StoB_REQ7_p & !v8a87cd;
assign v8e444a = jx2_p & v8e5a18 | !jx2_p & !v85e33b;
assign v85f57e = jx1_p & v85b2ae | !jx1_p & !v844f91;
assign v856f22 = StoB_REQ1_p & v866812 | !StoB_REQ1_p & v876a22;
assign v89925a = StoB_REQ1_p & v8dc67d | !StoB_REQ1_p & v86653e;
assign v85e61d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85b0a3;
assign v8635e4 = ENQ_p & v8572d0 | !ENQ_p & v845039;
assign v85ada7 = jx0_p & v86baf9 | !jx0_p & v85b9a9;
assign v881baf = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e14bc;
assign v8b5792 = jx1_p & v844f91 | !jx1_p & v8b56f8;
assign v8e5075 = BtoS_ACK3_p & v8e16ea | !BtoS_ACK3_p & v880dfd;
assign v85660f = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8e50c2;
assign v8b571e = BtoS_ACK7_p & v8e1c27 | !BtoS_ACK7_p & !v8b5832;
assign v8572f7 = BtoS_ACK0_p & v883ca3 | !BtoS_ACK0_p & v8e56dc;
assign v865131 = jx1_p & v8e4514 | !jx1_p & v86007f;
assign v8a6914 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v85c941;
assign v844fa3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844f91;
assign v85f334 = jx2_p & v8af47a | !jx2_p & v8b54f4;
assign v856669 = DEQ_p & v8e1651 | !DEQ_p & !v844f91;
assign v8618f2 = jx2_p & v85d886 | !jx2_p & v85653c;
assign v8e1cd8 = stateG12_p & v860057 | !stateG12_p & v844f91;
assign v86653e = BtoS_ACK2_p & v8e519b | !BtoS_ACK2_p & v8e5908;
assign v8e1f59 = RtoB_ACK0_p & v85fc37 | !RtoB_ACK0_p & v8dc668;
assign v8b55d5 = DEQ_p & v8e1090 | !DEQ_p & v844f91;
assign v85ae38 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8cc8e8;
assign v8e59ca = BtoS_ACK1_p & v85c469 | !BtoS_ACK1_p & v85e836;
assign v8b5756 = BtoS_ACK7_p & v8e3c83 | !BtoS_ACK7_p & v8b585a;
assign v8e4bdc = jx0_p & v8b56ef | !jx0_p & v85c433;
assign v87356b = BtoS_ACK8_p & v8e5a22 | !BtoS_ACK8_p & v8b586c;
assign v8e4caf = StoB_REQ3_p & v85ea8d | !StoB_REQ3_p & !v844f91;
assign v8e1813 = jx1_p & v85acf3 | !jx1_p & !v8b55a1;
assign v8e55a3 = BtoS_ACK1_p & v8a87b4 | !BtoS_ACK1_p & v86b6cf;
assign v8e1590 = jx0_p & v85adf5 | !jx0_p & !v8e18fe;
assign v85d34c = BtoS_ACK6_p & v880bc4 | !BtoS_ACK6_p & v8563be;
assign v8e52f8 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85f287;
assign v85ccc6 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v844fa5;
assign v8b55bd = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844faf;
assign v8e5bb2 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856b48;
assign v85f7ea = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b56a9;
assign v8e3db6 = StoB_REQ8_p & v8e2288 | !StoB_REQ8_p & v8e4f0c;
assign v85e5cf = BtoS_ACK0_p & v8e4831 | !BtoS_ACK0_p & v8b5544;
assign v8e45e3 = jx1_p & v844f91 | !jx1_p & !v8e5a2f;
assign v8dc58d = BtoS_ACK7_p & v8e3ca1 | !BtoS_ACK7_p & !v856803;
assign v8b5668 = BtoS_ACK8_p & v8e3d91 | !BtoS_ACK8_p & v85f49e;
assign v8e5344 = StoB_REQ6_p & v885fa8 | !StoB_REQ6_p & v8a5bb4;
assign v866593 = BtoS_ACK8_p & v845026 | !BtoS_ACK8_p & v8e3bbb;
assign v8e162c = jx2_p & v8b5765 | !jx2_p & v8b55bf;
assign v85bbcc = BtoS_ACK8_p & v8be11a | !BtoS_ACK8_p & !v8e4a48;
assign v8564fa = BtoS_ACK7_p & v8e1933 | !BtoS_ACK7_p & v85d69a;
assign v8e5a9d = jx0_p & v844f9f | !jx0_p & v844f91;
assign v86f9a1 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f99;
assign v8e5a13 = ENQ_p & v8af34b | !ENQ_p & v85cbe8;
assign v8e1f47 = StoB_REQ0_p & v85db90 | !StoB_REQ0_p & v8cc8f2;
assign v85de0b = StoB_REQ1_p & v861740 | !StoB_REQ1_p & v8b567b;
assign v86d0c6 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8e1d21;
assign v8e53a5 = jx2_p & v86584f | !jx2_p & !v870e66;
assign v8e5252 = jx2_p & v8563a6 | !jx2_p & v8b552a;
assign v8af11e = jx2_p & v8e5b58 | !jx2_p & v8e41ec;
assign v8cce49 = BtoS_ACK6_p & v85768f | !BtoS_ACK6_p & v8b5724;
assign v85da20 = BtoS_ACK6_p & v8e42a4 | !BtoS_ACK6_p & v86290d;
assign v8e4d85 = BtoS_ACK2_p & v8e16ea | !BtoS_ACK2_p & v8e5075;
assign v85cccf = jx1_p & v8e229e | !jx1_p & !v8e400a;
assign v8b58aa = StoB_REQ7_p & v845249 | !StoB_REQ7_p & v844f91;
assign v85708d = jx1_p & v85c8f2 | !jx1_p & v8e17b8;
assign v8b56db = jx2_p & v8565e5 | !jx2_p & v844f91;
assign v8be143 = BtoS_ACK7_p & v856264 | !BtoS_ACK7_p & v85c593;
assign v856f8d = jx1_p & v8e549e | !jx1_p & !v8e4254;
assign v85ccc3 = jx0_p & v8b5757 | !jx0_p & !v84507a;
assign v8e4916 = RtoB_ACK1_p & v8b5565 | !RtoB_ACK1_p & v888cd4;
assign v8b572a = BtoS_ACK7_p & v8e176c | !BtoS_ACK7_p & v8b58ad;
assign v85d812 = ENQ_p & v85ba14 | !ENQ_p & v866593;
assign v859fe4 = jx0_p & v85e50d | !jx0_p & !v844f91;
assign v8b55c2 = jx0_p & v85b898 | !jx0_p & v8451cf;
assign v85e946 = BtoS_ACK0_p & v8b5663 | !BtoS_ACK0_p & v8e5c0a;
assign v8b588f = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v85bbe2;
assign v844fb7 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f91;
assign v856255 = StoB_REQ6_p & v86290d | !StoB_REQ6_p & v865d5b;
assign v8b5771 = BtoS_ACK0_p & v85f2f8 | !BtoS_ACK0_p & v8e38b0;
assign v8e19b1 = BtoS_ACK1_p & v85dbdd | !BtoS_ACK1_p & v85d42f;
assign v8e4391 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v856eba;
assign v889290 = BtoS_ACK7_p & v85e947 | !BtoS_ACK7_p & v8dc554;
assign v8575eb = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v856367;
assign v84514a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8860f1;
assign v845160 = StoB_REQ8_p & v856867 | !StoB_REQ8_p & v85aba0;
assign v8dc5d8 = BtoS_ACK0_p & v899247 | !BtoS_ACK0_p & v8b5839;
assign v8e5a2b = BtoS_ACK7_p & v8e499d | !BtoS_ACK7_p & !v8e4e9e;
assign v85f2cd = BtoS_ACK1_p & v8e5bb2 | !BtoS_ACK1_p & v88173a;
assign v8e3c9e = StoB_REQ1_p & v88924e | !StoB_REQ1_p & !v85a6a9;
assign v8bf910 = jx3_p & v864a5d | !jx3_p & v85ca8a;
assign v85d9d8 = jx0_p & v844f91 | !jx0_p & !v85e7ea;
assign v85c4c3 = StoB_REQ1_p & v8e407e | !StoB_REQ1_p & v8b580b;
assign v8e4f37 = jx2_p & v8e3ec6 | !jx2_p & v85dfab;
assign v8e59de = jx1_p & v844f91 | !jx1_p & v8e22d4;
assign v8af47a = jx1_p & v8e5aa3 | !jx1_p & v8e2267;
assign v8e3ea1 = StoB_REQ8_p & v8a5cca | !StoB_REQ8_p & v8e162b;
assign v8e466b = StoB_REQ0_p & v85ccc3 | !StoB_REQ0_p & v85d5a0;
assign BtoS_ACK1_n = !v8cc9b5;
assign v8e1e59 = jx2_p & v8e4b4d | !jx2_p & v844f91;
assign v8b5731 = BtoS_ACK6_p & v8e3bf7 | !BtoS_ACK6_p & v8af0de;
assign v8af34f = BtoS_ACK7_p & v8e4636 | !BtoS_ACK7_p & !v8e44a1;
assign v8452dc = BtoS_ACK0_p & v8e4c47 | !BtoS_ACK0_p & v8e22c3;
assign v8e38c3 = jx2_p & v8e4184 | !jx2_p & v8e188a;
assign v88c339 = BtoS_ACK6_p & v8e4c11 | !BtoS_ACK6_p & v85d6a8;
assign v8e2440 = jx1_p & v85acf3 | !jx1_p & !v880b12;
assign v85abc2 = BtoS_ACK2_p & v8bf0c7 | !BtoS_ACK2_p & v85bd68;
assign v85d9cc = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v856f79;
assign v85f33d = StoB_REQ1_p & v8e1e8c | !StoB_REQ1_p & v844f91;
assign v85cc56 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856479;
assign v8b5516 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b576f;
assign v8e5a51 = StoB_REQ1_p & v8e4f80 | !StoB_REQ1_p & v8e213d;
assign v85afbc = BtoS_ACK0_p & v85e0b0 | !BtoS_ACK0_p & v859fe5;
assign v8e5049 = BtoS_ACK7_p & v88928c | !BtoS_ACK7_p & v8b57ab;
assign v85d35a = EMPTY_p & v85a277 | !EMPTY_p & v8b54f0;
assign v8b5689 = jx1_p & v8b5862 | !jx1_p & v8e4761;
assign v8b5674 = jx0_p & v85da91 | !jx0_p & v8e47d6;
assign v85b60a = jx2_p & v85cb8e | !jx2_p & !v844f91;
assign v8e1931 = StoB_REQ7_p & v8e4e81 | !StoB_REQ7_p & v8b5658;
assign v856e07 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v85cd1c;
assign v8e5194 = BtoS_ACK8_p & v8e5833 | !BtoS_ACK8_p & v8e4ad3;
assign v8a5b9d = jx2_p & v8e4e99 | !jx2_p & !v8e21cf;
assign v8b568f = jx2_p & v856ef1 | !jx2_p & !v8e4ac8;
assign v8e460c = BtoS_ACK1_p & v8e4632 | !BtoS_ACK1_p & v8e1c87;
assign v8e4959 = StoB_REQ8_p & v86290d | !StoB_REQ8_p & v844f91;
assign v88bcd0 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8af160;
assign v8573cf = EMPTY_p & v8af461 | !EMPTY_p & v8e4c64;
assign v8e3a10 = stateG7_1_p & v856725 | !stateG7_1_p & !v844f91;
assign v857010 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v867a58;
assign v8e20a4 = ENQ_p & v8572d0 | !ENQ_p & v8e10fb;
assign v857542 = jx0_p & v8e4d94 | !jx0_p & v8e3bba;
assign v8e4261 = jx0_p & v8b5698 | !jx0_p & v8e51cd;
assign v85e994 = jx1_p & v8e5a64 | !jx1_p & v8e1857;
assign SLC0_n = v8a5564;
assign v8e59c0 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v856eba;
assign v8b56e5 = BtoS_ACK0_p & v8b575f | !BtoS_ACK0_p & v84514a;
assign v85e664 = BtoS_ACK8_p & v8e5223 | !BtoS_ACK8_p & v85ad8b;
assign v8e453e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e57d3;
assign v85b979 = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v8e5468;
assign v8b554b = BtoS_ACK8_p & v8e4b00 | !BtoS_ACK8_p & v8a5c15;
assign v8e1b90 = BtoS_ACK7_p & v85d805 | !BtoS_ACK7_p & v8e58e4;
assign v85c639 = jx1_p & v8e4514 | !jx1_p & v8e5366;
assign v8b5858 = BtoR_REQ1_p & v8e2475 | !BtoR_REQ1_p & v856b8e;
assign v85f6bc = jx0_p & v85e000 | !jx0_p & !v8e5bb2;
assign v8b57bd = EMPTY_p & v844fc9 | !EMPTY_p & !v844fcb;
assign v8b58a7 = jx1_p & v8b56ee | !jx1_p & v8e1841;
assign v8e1c26 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8b5526;
assign v8e1982 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af37f;
assign v8e535e = jx2_p & v8e2440 | !jx2_p & v8e55cf;
assign v8e51d9 = BtoS_ACK0_p & v8e5033 | !BtoS_ACK0_p & !v85ba51;
assign v866529 = jx1_p & v8b56ca | !jx1_p & v844f91;
assign v8b57ae = ENQ_p & v8af34b | !ENQ_p & v85d8e2;
assign v8e44a2 = EMPTY_p & v85f59c | !EMPTY_p & v8e522a;
assign v8e55e7 = BtoS_ACK8_p & v8b555e | !BtoS_ACK8_p & v8b5773;
assign v8e3a16 = DEQ_p & v8e3af2 | !DEQ_p & v8b589f;
assign v860064 = BtoS_ACK1_p & v8e4632 | !BtoS_ACK1_p & v8e1d32;
assign v856bd5 = BtoS_ACK6_p & v8e59c6 | !BtoS_ACK6_p & v8af292;
assign v8e4d0d = jx0_p & v8e4d94 | !jx0_p & !v85db0d;
assign v8be167 = BtoS_ACK2_p & v8bf0c7 | !BtoS_ACK2_p & v8b58ae;
assign v8e46da = jx0_p & v844f91 | !jx0_p & v84507a;
assign v8566f3 = BtoS_ACK2_p & v8e3883 | !BtoS_ACK2_p & v8b54d6;
assign v8e207d = jx1_p & v85ccec | !jx1_p & !v8dc5cb;
assign v85e111 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8e576d;
assign v866552 = BtoS_ACK1_p & v8e3d7b | !BtoS_ACK1_p & v85d3c7;
assign v899197 = jx1_p & v844f91 | !jx1_p & v88d5d7;
assign v8e58fd = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844fbb;
assign v85a863 = jx1_p & v8b56ee | !jx1_p & v8e45fa;
assign v8e5a00 = BtoS_ACK1_p & v8e16ea | !BtoS_ACK1_p & v85e0b5;
assign v85bd37 = StoB_REQ8_p & v8b5662 | !StoB_REQ8_p & v8e438a;
assign v8e4212 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85ca40;
assign v8e42ab = EMPTY_p & v84510d | !EMPTY_p & v85a4f0;
assign v85fa42 = StoB_REQ8_p & v889290 | !StoB_REQ8_p & v85c754;
assign v85c73d = EMPTY_p & v8e3cfe | !EMPTY_p & v85ae46;
assign v8e5173 = BtoS_ACK2_p & v8b550c | !BtoS_ACK2_p & !v8e3dec;
assign v8e5033 = jx0_p & v844f97 | !jx0_p & !v844f91;
assign v85a98f = jx2_p & v8e388a | !jx2_p & v8e4e45;
assign v8b56cd = StoB_REQ6_p & v85bdac | !StoB_REQ6_p & v8be147;
assign v85726b = BtoR_REQ0_p & v8e1aa8 | !BtoR_REQ0_p & v85a893;
assign v85b739 = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & v8b5757;
assign v8e4a06 = StoB_REQ3_p & v8e18dd | !StoB_REQ3_p & v844f9f;
assign v8dc65c = BtoS_ACK0_p & v85e0b0 | !BtoS_ACK0_p & v8b589d;
assign v8e5468 = jx2_p & v8e5897 | !jx2_p & v8e1811;
assign v8e4602 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e4636;
assign v8e1852 = BtoS_ACK8_p & v8e17d6 | !BtoS_ACK8_p & v85da27;
assign v880b8e = jx2_p & v88c371 | !jx2_p & v86d6bd;
assign v8e1b02 = BtoS_ACK1_p & v899202 | !BtoS_ACK1_p & v8dc5ad;
assign v8e1a00 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v844f99;
assign v8e48a0 = StoB_REQ6_p & v85b238 | !StoB_REQ6_p & v856c6d;
assign v8af243 = jx0_p & v8b5757 | !jx0_p & !v844f97;
assign v8e2121 = StoB_REQ6_p & v86290d | !StoB_REQ6_p & !v844f91;
assign jx0_n = !v8992c3;
assign v8e417e = StoB_REQ3_p & v85c4b8 | !StoB_REQ3_p & v8e18dd;
assign v8b56ee = StoB_REQ7_p & v86290d | !StoB_REQ7_p & !v844f91;
assign v8e5aa3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8be0ec;
assign v85e103 = StoB_REQ7_p & v85b3c3 | !StoB_REQ7_p & v8af176;
assign v85dbda = jx0_p & v844f9b | !jx0_p & v844f91;
assign v856ad9 = jx1_p & v8e59d4 | !jx1_p & v8803e2;
assign v8e4eef = jx1_p & v85dee1 | !jx1_p & !v8e1618;
assign v8e597e = BtoS_ACK6_p & v85cbd3 | !BtoS_ACK6_p & v8e50a2;
assign v8e45a8 = BtoS_ACK7_p & v8a5c84 | !BtoS_ACK7_p & !v8ca6f1;
assign v857144 = DEQ_p & v8e2154 | !DEQ_p & v8b55ed;
assign v856705 = StoB_REQ1_p & v8e4294 | !StoB_REQ1_p & v8e3c75;
assign SLC2_n = v865261;
assign v85ba51 = StoB_REQ0_p & v88c2b9 | !StoB_REQ0_p & v88d5d7;
assign v8e17e8 = jx0_p & v8e19f0 | !jx0_p & v8a5b4f;
assign v8e46ed = StoB_REQ7_p & v8af418 | !StoB_REQ7_p & v8e3c2f;
assign v86e8c2 = StoB_REQ5_n & v8e5000 | !StoB_REQ5_n & v844f91;
assign v8e3926 = BtoS_ACK7_p & v85d3d0 | !BtoS_ACK7_p & v8e4baa;
assign v865764 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8e4959;
assign v856c6c = EMPTY_p & v8e56dd | !EMPTY_p & v8e14ca;
assign v856598 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8b5800;
assign v8e503e = DEQ_p & v8e4103 | !DEQ_p & v85a893;
assign v8cce14 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v861740;
assign v8e5906 = jx1_p & v8e5a73 | !jx1_p & v86290d;
assign v856bc8 = StoB_REQ1_p & v856e07 | !StoB_REQ1_p & !v856eba;
assign v85cc98 = DEQ_p & v8e1dbf | !DEQ_p & v85a893;
assign v85da9f = BtoS_ACK7_p & v8618f2 | !BtoS_ACK7_p & v8b5736;
assign v8b561b = jx2_p & v8b5805 | !jx2_p & !v845136;
assign v8e15ab = BtoS_ACK0_p & v8e3d0c | !BtoS_ACK0_p & v8b582f;
assign v85f2c8 = jx0_p & v85b6b5 | !jx0_p & !v8e55c9;
assign v8a87b4 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8bf0c7;
assign v8b5624 = jx1_p & v8e4172 | !jx1_p & v85a622;
assign v889f9b = stateG12_p & v8658a0 | !stateG12_p & v85fb12;
assign v8b55c7 = EMPTY_p & v8e20a4 | !EMPTY_p & v857056;
assign v8b57b5 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8e4638;
assign v8e3dc6 = StoB_REQ0_p & v883ca3 | !StoB_REQ0_p & v8568a1;
assign v85cb94 = jx2_p & v8b58a7 | !jx2_p & v8b553b;
assign v8cc8e9 = jx2_p & v85f411 | !jx2_p & v86290d;
assign v8e53c6 = jx1_p & v8e50df | !jx1_p & v8b5872;
assign v8cce2b = jx1_p & v8b5844 | !jx1_p & v8e59df;
assign v8b35f5 = jx1_p & v8e4514 | !jx1_p & v8452dc;
assign v85fbed = StoB_REQ0_p & v8e42b6 | !StoB_REQ0_p & v883ca1;
assign v8e48fc = EMPTY_p & v8b55ac | !EMPTY_p & v8e436f;
assign v85d794 = StoB_REQ1_p & v85cd1c | !StoB_REQ1_p & v844f91;
assign v8b552b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v859fe9;
assign v85dddb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v85e7ea;
assign v8e58e4 = BtoS_ACK6_p & v85d805 | !BtoS_ACK6_p & v8e1ccb;
assign v8e1579 = jx2_p & v8e3db0 | !jx2_p & v856edf;
assign v8e1ccb = jx2_p & v8b5792 | !jx2_p & v85b49f;
assign v85ea8d = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9d;
assign v856fe8 = jx2_p & v8b568e | !jx2_p & v85e1a0;
assign v8e5a8f = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v8e5000;
assign v8a5c58 = jx2_p & v8e51d0 | !jx2_p & v86290f;
assign v857615 = StoB_REQ0_p & v8e400a | !StoB_REQ0_p & v867b8d;
assign v8b5799 = jx0_p & v8e3c39 | !jx0_p & v8af15c;
assign v8b54c1 = BtoS_ACK3_p & v8b5875 | !BtoS_ACK3_p & !v8665a9;
assign v85e27e = StoB_REQ7_p & v8e4050 | !StoB_REQ7_p & v884bb3;
assign v8b588a = BtoS_ACK6_p & v85e947 | !BtoS_ACK6_p & v8e5942;
assign v8e17b8 = StoB_REQ6_p & v85aea9 | !StoB_REQ6_p & v8e2436;
assign v8b584a = jx0_p & v8e4fad | !jx0_p & v844f91;
assign v85f647 = BtoS_ACK1_p & v8e19f0 | !BtoS_ACK1_p & v8af31b;
assign v85fb12 = BtoS_ACK8_p & v8e3f6f | !BtoS_ACK8_p & v8b5614;
assign v8b56f7 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85fc4d;
assign v85ba14 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v8b56a3;
assign v8e1542 = jx1_p & v86cb45 | !jx1_p & v85abee;
assign v8b56fd = jx0_p & v844f91 | !jx0_p & !v8b5516;
assign v85cb88 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v85d6ab;
assign v8563a6 = jx1_p & v8ca185 | !jx1_p & !v8e5a63;
assign v85e9c5 = jx0_p & v844f91 | !jx0_p & v8b5757;
assign v8b55a2 = jx0_p & v85e7be | !jx0_p & !v85cb96;
assign v8af36d = DEQ_p & v8b5527 | !DEQ_p & !v844f91;
assign v8b5893 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8e4637;
assign v8e2239 = EMPTY_p & v86290d | !EMPTY_p & !v85e81e;
assign v8b576e = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v8e1aea;
assign v85a600 = BtoS_ACK8_p & v8b5820 | !BtoS_ACK8_p & v845160;
assign v8b5840 = jx2_p & v8e4d75 | !jx2_p & v868a25;
assign v8e5494 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v8a87b4;
assign v8dc5cb = StoB_REQ7_p & v8e59c7 | !StoB_REQ7_p & v8b5595;
assign v8b5687 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8e58d6;
assign v8566b6 = jx1_p & v8b58b2 | !jx1_p & v8b5779;
assign v86cbc7 = BtoS_ACK8_p & v865856 | !BtoS_ACK8_p & v8e592b;
assign v8b5862 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af383;
assign v85f34e = BtoS_ACK6_p & v8e176c | !BtoS_ACK6_p & v8e5b7d;
assign v85d3e9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85daf5;
assign v8e484f = jx1_p & v8572f7 | !jx1_p & !v844f91;
assign v8e58b0 = DEQ_p & v8b57a6 | !DEQ_p & v8569df;
assign v85744d = BtoS_ACK6_p & v85dd64 | !BtoS_ACK6_p & v8db83f;
assign v8e1eb9 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v8e519b;
assign v8e502c = BtoS_ACK6_p & v8e1579 | !BtoS_ACK6_p & v8bf339;
assign v8e4131 = jx2_p & v8b58a7 | !jx2_p & v8b57c1;
assign v8e455f = BtoR_REQ1_p & v8e3a67 | !BtoR_REQ1_p & v8b5848;
assign v8b55a7 = EMPTY_p & v8e4022 | !EMPTY_p & v8893a8;
assign v856b36 = jx2_p & v880b9c | !jx2_p & v8e2248;
assign v8e1f02 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b56eb;
assign v8e1893 = StoB_REQ6_p & v8e23ae | !StoB_REQ6_p & v8dc5d8;
assign v85d7c8 = BtoS_ACK7_p & v85638e | !BtoS_ACK7_p & v8e58a7;
assign v8e59f6 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v867aa7;
assign v8b5663 = jx0_p & v8e5996 | !jx0_p & !v8e49ee;
assign v8452fa = jx1_p & v867aa7 | !jx1_p & !v889264;
assign v85f697 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e417e;
assign v88e287 = BtoS_ACK0_p & v8e550e | !BtoS_ACK0_p & v84521c;
assign v84521c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85d59f;
assign v8b5764 = BtoS_ACK2_p & v8a5bcf | !BtoS_ACK2_p & v8e58c4;
assign v8e4ffe = StoB_REQ0_p & v889fde | !StoB_REQ0_p & v8e51e4;
assign v8e5a11 = StoB_REQ8_p & v8e4235 | !StoB_REQ8_p & v8e2229;
assign v8e4d94 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85db04;
assign v8b57e9 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8e5aa0;
assign v8e41d9 = jx1_p & v8e53e7 | !jx1_p & v844f91;
assign v8e5bd5 = StoB_REQ3_p & v85ea8d | !StoB_REQ3_p & v8e1d33;
assign v85e60f = BtoS_ACK0_p & v8e5913 | !BtoS_ACK0_p & v8e5c69;
assign v8e1934 = StoB_REQ2_p & v8b57f2 | !StoB_REQ2_p & v8e3b0a;
assign v85adaf = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v85e1b8;
assign v8cce20 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b5554;
assign v8e5b2c = BtoS_ACK0_p & v85c941 | !BtoS_ACK0_p & v8e5a71;
assign v85da8e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b5525;
assign v8b57ff = BtoS_ACK0_p & v8e3d0c | !BtoS_ACK0_p & v8e587f;
assign v856345 = StoB_REQ7_p & v85a8af | !StoB_REQ7_p & v8e548f;
assign v85f2aa = BtoS_ACK6_p & v85f6b4 | !BtoS_ACK6_p & v8e4d29;
assign v8e2035 = StoB_REQ0_p & v88d5d7 | !StoB_REQ0_p & !v844f91;
assign v8b5651 = StoB_REQ0_p & v86290d | !StoB_REQ0_p & v8626fe;
assign v8b5699 = jx0_p & v8e4831 | !jx0_p & !v844f91;
assign v8e4229 = jx0_p & v844f9f | !jx0_p & !v8e460c;
assign v8e4579 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v860886;
assign v8e10c0 = BtoS_ACK6_p & v85f64e | !BtoS_ACK6_p & v8b584c;
assign v856a21 = jx0_p & v88c324 | !jx0_p & !v8b5516;
assign v85c120 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85e006;
assign v8e564d = StoB_REQ0_p & v883ca3 | !StoB_REQ0_p & v8e5048;
assign v8b575b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v85db1a;
assign v85a25b = jx2_p & v8cce04 | !jx2_p & v88bbf7;
assign v8e3cf8 = StoB_REQ0_p & v8e464c | !StoB_REQ0_p & v8e4831;
assign v8e1e94 = RtoB_ACK1_p & v8b557d | !RtoB_ACK1_p & v85ce72;
assign v84510d = BtoS_ACK8_p & v863508 | !BtoS_ACK8_p & v8af3b8;
assign v8e597f = jx2_p & v856c2e | !jx2_p & !v8e4c34;
assign v8e44dd = BtoS_ACK0_p & v8b56e6 | !BtoS_ACK0_p & v8e1590;
assign v856358 = jx1_p & v8991fe | !jx1_p & v856345;
assign v8e5707 = BtoS_ACK7_p & v8b55b0 | !BtoS_ACK7_p & v856a2e;
assign v8b55e7 = StoB_REQ1_p & v85d671 | !StoB_REQ1_p & v8b5515;
assign v8e20fa = BtoS_ACK3_p & v844fa0 | !BtoS_ACK3_p & !v844f91;
assign v8b58b1 = stateG7_1_p & v8e41a5 | !stateG7_1_p & v85f839;
assign v85bd67 = jx1_p & v85e383 | !jx1_p & v844f91;
assign v8e5a18 = jx1_p & v8b58b2 | !jx1_p & v85a0f3;
assign v863db8 = DEQ_p & v85696e | !DEQ_p & v8af26f;
assign v8e47f8 = StoB_REQ7_p & v8e59f9 | !StoB_REQ7_p & v85e951;
assign v8e4118 = StoB_REQ0_p & v85f2c8 | !StoB_REQ0_p & v85e362;
assign v8b5607 = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & v85afc0;
assign v8564de = BtoS_ACK1_p & v8e2265 | !BtoS_ACK1_p & v85a51b;
assign v85a24b = jx0_p & v88c324 | !jx0_p & v8e4831;
assign v844fbf = BtoS_ACK8_p & v844f91 | !BtoS_ACK8_p & !v844f91;
assign v85fa3e = StoB_REQ2_p & v8db8b5 | !StoB_REQ2_p & v8574d0;
assign v8567bb = StoB_REQ0_p & v883ca3 | !StoB_REQ0_p & v8e3d0c;
assign v85de73 = BtoS_ACK7_p & v8e5a5e | !BtoS_ACK7_p & v8566fb;
assign v85acfd = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85a0bf;
assign v8e1f1b = stateG12_p & v8b55ac | !stateG12_p & v8e1d09;
assign v8b5543 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856452;
assign v8819a3 = jx0_p & v845380 | !jx0_p & !v85724d;
assign v85b3c3 = BtoS_ACK0_p & v88d5d7 | !BtoS_ACK0_p & v85b739;
assign v8b57a6 = stateG12_p & v8569df | !stateG12_p & v844f91;
assign v85fb1e = jx2_p & v8e4b9f | !jx2_p & v8e58b4;
assign v85b863 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v856312;
assign v8af1a0 = BtoS_ACK8_p & v870b4c | !BtoS_ACK8_p & !v8e238b;
assign v8e58cf = StoB_REQ7_p & v85660c | !StoB_REQ7_p & v8e4b4e;
assign v8e42b6 = jx0_p & v8cce14 | !jx0_p & v844f91;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v8b5728 = DEQ_p & v844f91 | !DEQ_p & !v85e5db;
assign v8e229e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b5838;
assign v86dabf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b55cb;
assign v8e22ae = BtoS_ACK6_p & v856ca7 | !BtoS_ACK6_p & v85d539;
assign v88460a = jx1_p & v8b56ee | !jx1_p & v8e593d;
assign v8b5614 = StoB_REQ8_p & v844f91 | !StoB_REQ8_p & v856c90;
assign v889f0f = EMPTY_p & v8573c8 | !EMPTY_p & v8e58ae;
assign v856be2 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8e1abe;
assign v8b54de = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8e5692;
assign v85d376 = StoB_REQ0_p & v85d98f | !StoB_REQ0_p & v859ffb;
assign v8e21c8 = StoB_REQ8_p & v8e1f73 | !StoB_REQ8_p & v8b571e;
assign v8a887e = jx3_p & v8dc5b0 | !jx3_p & v861ca6;
assign v85c895 = jx0_p & v844f91 | !jx0_p & v86ea54;
assign v85664e = BtoS_ACK8_p & v8af12b | !BtoS_ACK8_p & !v845064;
assign v864f49 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8e5989;
assign v8e17ae = DEQ_p & v860006 | !DEQ_p & v860057;
assign v85d5b1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8bf8d3;
assign v8e4b2a = jx1_p & v8e4988 | !jx1_p & v8e2267;
assign v85d750 = BtoR_REQ1_p & v8e5b8b | !BtoR_REQ1_p & v8e20ba;
assign v86a790 = BtoS_ACK7_p & v8b55b0 | !BtoS_ACK7_p & v8b5685;
assign v8e420f = jx2_p & v8e43fa | !jx2_p & v856a93;
assign v8b585b = stateG12_p & v8e1695 | !stateG12_p & !v8601d6;
assign v85dcb9 = EMPTY_p & v862719 | !EMPTY_p & v8e1eab;
assign v8b56a8 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85f33d;
assign v8e594c = jx2_p & v8be0f6 | !jx2_p & !v8b55bf;
assign v8664e6 = jx0_p & v844f9f | !jx0_p & v85b29f;
assign v8e5a7e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85f35f;
assign v85666e = BtoR_REQ1_p & v85668b | !BtoR_REQ1_p & v8e3b74;
assign v8e4c6e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e4040;
assign v8e38b0 = jx0_p & v8e4f80 | !jx0_p & v8e4b64;
assign v8e4224 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v85ea8d;
assign v85f9b8 = BtoS_ACK8_p & v844fa3 | !BtoS_ACK8_p & !v8cc8c3;
assign v8dc60e = ENQ_p & v85e45f | !ENQ_p & v8ccdf5;
assign v856688 = BtoS_ACK5_p & v844fb7 | !BtoS_ACK5_p & v8e5000;
assign v8b55f8 = StoB_REQ2_p & v8e3f79 | !StoB_REQ2_p & v88c31b;
assign v8e57a4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e3e1e;
assign v85d69a = BtoS_ACK6_p & v8e3b37 | !BtoS_ACK6_p & v8e5896;
assign v85e566 = jx0_p & v8e4b93 | !jx0_p & !v8e111b;
assign v85deb3 = BtoS_ACK6_p & v85d805 | !BtoS_ACK6_p & v884319;
assign v8e5a08 = DEQ_p & v8e41fc | !DEQ_p & v8cc95b;
assign v8e5723 = jx2_p & v8e59bd | !jx2_p & v8b55f4;
assign v8e58f1 = StoB_REQ0_p & v8991c9 | !StoB_REQ0_p & v8b56a9;
assign v85d9f0 = BtoS_ACK6_p & v8e4f37 | !BtoS_ACK6_p & v8571d6;
assign v883b69 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v85de51;
assign v856c3d = StoB_REQ3_p & v85ea8d | !StoB_REQ3_p & v844fb7;
assign v84530b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v882912;
assign v8b55b8 = StoB_REQ0_p & v8a54f3 | !StoB_REQ0_p & v86d72e;
assign v8e1ee5 = BtoS_ACK0_p & v8e5048 | !BtoS_ACK0_p & v8b56ed;
assign v85650e = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8b58ae;
assign v856fc9 = jx2_p & v85a23c | !jx2_p & v8b55bf;
assign v8e3d66 = DEQ_p & v8b569b | !DEQ_p & v84501d;
assign v86513d = BtoS_ACK7_p & v8e4764 | !BtoS_ACK7_p & v89928e;
assign v8565a2 = EMPTY_p & v85f343 | !EMPTY_p & v8e4497;
assign v85f6b4 = jx2_p & v8e1bf9 | !jx2_p & !v8cb249;
assign v88c2e1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8e1da5;
assign v8e1678 = StoB_REQ6_p & v8e157d | !StoB_REQ6_p & v85ea99;
assign v85da5d = RtoB_ACK0_p & v8e598e | !RtoB_ACK0_p & v8e4fe9;
assign v8e45d6 = BtoS_ACK1_p & v8e1eb9 | !BtoS_ACK1_p & v85f223;
assign ENQ_n = (BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!SLC0_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!SLC0_n & ((BtoS_ACK2_n))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((RtoB_ACK0_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((EMPTY_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((BtoR_REQ0_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((EMPTY_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((EMPTY_n & ((stateG7_1_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n & ((!StoB_REQ4_n))))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((EMPTY_n & ((stateG7_0_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!SLC0_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!SLC0_n & ((BtoS_ACK2_n))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))) | (!SLC1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!stateG7_0_n & ((BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n))))))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))) | (!jx0_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((!jx0_n))))) | (!jx3_n & ((StoB_REQ8_n))))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((!jx0_n))))) | (!jx3_n & ((StoB_REQ8_n))))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((!jx0_n))))) | (!jx3_n & ((StoB_REQ8_n))))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK8_n & ((StoB_REQ8_n))) | (!BtoS_ACK8_n & ((jx3_n & ((StoB_REQ8_n & ((BtoS_ACK7_n & ((jx0_n & ((StoB_REQ7_n))))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ8_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))) | (!jx3_n & ((StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!jx1_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))) | (!StoB_REQ0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))))))) | (!StoB_REQ8_n & ((jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((jx0_n & ((jx1_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((!StoB_REQ5_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC2_n & ((!SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK5_n & ((StoB_REQ5_n & ((!BtoS_ACK4_n))))))))))) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!SLC2_n & ((SLC1_n & ((!BtoS_ACK1_n & ((SLC0_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))) | (!SLC1_n & ((StoB_REQ1_n & ((BtoS_ACK1_n & ((SLC0_n)))))))))))))))))))))))))))))))))))))));
assign SLC3_n = (BtoR_REQ1_n & ((EMPTY_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))))))) | (!RtoB_ACK1_n & ((BtoR_REQ0_n & ((EMPTY_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((EMPTY_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))))))) | (!RtoB_ACK0_n & ((EMPTY_n & ((stateG7_0_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG7_0_n & ((BtoS_ACK8_n & ((jx3_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx3_n & ((jx2_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx2_n & ((ENQ_n))))))) | (!BtoS_ACK8_n & ((jx3_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx3_n & ((jx2_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((BtoS_ACK8_n & ((jx3_n & ((ENQ_n & ((!jx0_n))) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx3_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!stateG7_1_n & ((stateG12_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!DEQ_n & ((stateG12_n & ((BtoS_ACK8_n & ((jx3_n & ((ENQ_n & ((!jx0_n))) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx3_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))))) | (!stateG12_n & ((BtoS_ACK8_n & ((ENQ_n) | (!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK8_n & ((!ENQ_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n)))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  StoB_REQ4_p = 0;
  StoB_REQ5_p = 0;
  StoB_REQ6_p = 0;
  StoB_REQ7_p = 0;
  StoB_REQ8_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoS_ACK4_p = 0;
  BtoS_ACK5_p = 0;
  BtoS_ACK6_p = 0;
  BtoS_ACK7_p = 0;
  BtoS_ACK8_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  SLC2_p = 0;
  SLC3_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
  jx3_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  StoB_REQ4_p = StoB_REQ4_n;
  StoB_REQ5_p = StoB_REQ5_n;
  StoB_REQ6_p = StoB_REQ6_n;
  StoB_REQ7_p = StoB_REQ7_n;
  StoB_REQ8_p = StoB_REQ8_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoS_ACK4_p = BtoS_ACK4_n;
  BtoS_ACK5_p = BtoS_ACK5_n;
  BtoS_ACK6_p = BtoS_ACK6_n;
  BtoS_ACK7_p = BtoS_ACK7_n;
  BtoS_ACK8_p = BtoS_ACK8_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  SLC2_p = SLC2_n;
  SLC3_p = SLC3_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
  jx3_p = jx3_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
