module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hbusreq2, hlock2, hbusreq3, hlock3, hbusreq4, hlock4, hbusreq5, hlock5, hburst0, hburst1, hmaster0, hmaster1, hmaster2, hmastlock, start, decide, locked, hgrant0, hgrant1, hgrant2, hgrant3, hgrant4, hgrant5, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, stateG10_2, stateG10_3, stateG10_4, stateG10_5, jx0, jx1, jx2);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v845542;
  wire v84557e;
  wire v845560;
  wire v88d3e4;
  wire v10d3fd2;
  wire v10d3fd3;
  wire v10d3fd4;
  wire v10d3fd5;
  wire v10d3fd6;
  wire v10d3fd7;
  wire v845580;
  wire v10d3fd8;
  wire v10d3fd9;
  wire v10d3fda;
  wire v10d3fdb;
  wire v10d3fdc;
  wire v10d3fdd;
  wire v10d3fde;
  wire v10d3fdf;
  wire v10d3fe0;
  wire v10d3fe1;
  wire v10d3fe2;
  wire v10d3fe3;
  wire v10d3fe4;
  wire v10d3fe5;
  wire v10d3fe6;
  wire v10d3fe7;
  wire v10d3fe8;
  wire v10d3fe9;
  wire v10d3fea;
  wire v10d3feb;
  wire v10d3fec;
  wire v10d3fed;
  wire v10d3fee;
  wire v10d3fef;
  wire v10d3ff0;
  wire v10d3ff1;
  wire v10d3ff2;
  wire v10d3ff3;
  wire v10d3ff4;
  wire v10d3ff5;
  wire v10d3ff6;
  wire v10d3ff7;
  wire v10d3ff8;
  wire v10d3ff9;
  wire v10d3ffa;
  wire v10d3ffb;
  wire v10d3ffc;
  wire v10d3ffd;
  wire v10d3ffe;
  wire v10d3fff;
  wire v10d4000;
  wire v10d4001;
  wire v10d4002;
  wire v10d4006;
  wire v10d4007;
  wire v10d4008;
  wire v10d4009;
  wire v10d400a;
  wire v10d400b;
  wire v10d400c;
  wire v10d400d;
  wire v10d400e;
  wire v10d400f;
  wire v10d4010;
  wire v10d4011;
  wire v10d4012;
  wire v10d4013;
  wire v10d4014;
  wire v10d4015;
  wire v10d4016;
  wire v10d4017;
  wire v10d4018;
  wire v10d4019;
  wire v10d401a;
  wire v10d401b;
  wire v10d401c;
  wire v10d401d;
  wire v10d401e;
  wire v10d401f;
  wire v10d4020;
  wire v10d4021;
  wire v10d4022;
  wire v10d4023;
  wire v10d4024;
  wire v10d4025;
  wire v10d4026;
  wire v10d4027;
  wire v10d4028;
  wire v10d4029;
  wire v10d402a;
  wire v10d402b;
  wire v10d402c;
  wire v10d402d;
  wire v10d402e;
  wire v10d402f;
  wire v10d4030;
  wire v10d4031;
  wire v10d4032;
  wire v10d4033;
  wire v10d4034;
  wire v10d4035;
  wire v10d4036;
  wire v10d4037;
  wire v10d4038;
  wire v10d4039;
  wire v10d403a;
  wire v10d403b;
  wire v10d403c;
  wire v10d403d;
  wire v10d403e;
  wire v10d403f;
  wire v10d4040;
  wire v10d4041;
  wire v10d4042;
  wire v10d4043;
  wire v10d4044;
  wire v10d4045;
  wire v10d4046;
  wire v10d4047;
  wire v10d4048;
  wire v10d4049;
  wire v10d404a;
  wire v10d404b;
  wire v10d404c;
  wire v10d404d;
  wire v10d404e;
  wire v10d404f;
  wire v10d4050;
  wire v10d4051;
  wire v10d4052;
  wire v10d4053;
  wire v10d4054;
  wire v10d4055;
  wire v10d4056;
  wire v10d4057;
  wire v10d4058;
  wire v10d4059;
  wire v10d405a;
  wire v10d405b;
  wire v10d405c;
  wire v10d405d;
  wire v10d405e;
  wire v10d405f;
  wire v10d4060;
  wire v10d4061;
  wire v10d4062;
  wire v10d4063;
  wire v10d4064;
  wire v10d4065;
  wire v10d4066;
  wire v10d4067;
  wire v10d4068;
  wire v10d4069;
  wire v10d406a;
  wire v10d406b;
  wire v10d406c;
  wire v10d406d;
  wire v10d406e;
  wire v10d406f;
  wire v10d4070;
  wire v10d4071;
  wire v10d4072;
  wire v10d4073;
  wire v10d4074;
  wire v10d4075;
  wire v10d4076;
  wire v10d4077;
  wire v10d4078;
  wire v10d4079;
  wire v10d407a;
  wire v10d407b;
  wire v10d407c;
  wire v10d407d;
  wire v10d407e;
  wire v10d407f;
  wire v10d4080;
  wire v10d4081;
  wire v10d4082;
  wire v10d4083;
  wire v10d4084;
  wire v10d4085;
  wire v10d4086;
  wire v10d4087;
  wire v10d4088;
  wire v10d4089;
  wire v10d408a;
  wire v10d408b;
  wire v10d408c;
  wire v10d408d;
  wire v10d408e;
  wire v10d408f;
  wire v10d4090;
  wire v10d4091;
  wire v10d4092;
  wire v10d4093;
  wire v10d4094;
  wire v10d4095;
  wire v10d4096;
  wire v10d4097;
  wire v10d4098;
  wire v10d4099;
  wire v10d409a;
  wire v10d409b;
  wire v10d409c;
  wire v10d409d;
  wire v10d409e;
  wire v10d409f;
  wire v10d40a0;
  wire v10d40a1;
  wire v10d40a2;
  wire v10d40a3;
  wire v10d40a4;
  wire v10d40a5;
  wire v10d40a6;
  wire v10d40a7;
  wire v10d40a8;
  wire v10d40a9;
  wire v10d40aa;
  wire v10d40ab;
  wire v10d40ac;
  wire v10d40ad;
  wire v10d40ae;
  wire v10d40af;
  wire v10d40b0;
  wire v10d40b1;
  wire v10d40b2;
  wire v10d40b3;
  wire v10d40b4;
  wire v10d40b5;
  wire v10d40b6;
  wire v10d40b7;
  wire v10d40b8;
  wire v10d40b9;
  wire v10d40ba;
  wire v10d40bb;
  wire v10d40bc;
  wire v10d40bd;
  wire v10d40be;
  wire v10d40bf;
  wire v10d40c0;
  wire v10d40c1;
  wire v10d40c2;
  wire v10d40c3;
  wire v10d40c4;
  wire v10d40c5;
  wire v10d40c6;
  wire v10d40c7;
  wire v10d40c8;
  wire v10d40c9;
  wire v10d40ca;
  wire v10d40cb;
  wire v10d40cc;
  wire v10d40cd;
  wire v10d40ce;
  wire v10d40cf;
  wire v10d40d0;
  wire v10d40d1;
  wire v10d40d2;
  wire v10d40d3;
  wire v10d40d4;
  wire v10d40d5;
  wire v10d40d6;
  wire v10d40d7;
  wire v10d40d8;
  wire v10d40d9;
  wire v10d40da;
  wire v10d40db;
  wire v10d40dc;
  wire v10d40dd;
  wire v10d40de;
  wire v10d4264;
  wire v10d4265;
  wire v10d4266;
  wire v10d4267;
  wire v10d4268;
  wire v10d4269;
  wire v10d426a;
  wire v10d426b;
  wire v10d426c;
  wire v10d426d;
  wire v10d426e;
  wire v10d426f;
  wire v10d4270;
  wire v10d4271;
  wire v10d4272;
  wire v10d4273;
  wire v10d4274;
  wire v10d4275;
  wire v10d4276;
  wire v10d4277;
  wire v10d4278;
  wire v10d4279;
  wire v10d427a;
  wire v10d427b;
  wire v10d427c;
  wire v10d427d;
  wire v10d427e;
  wire v10d427f;
  wire v10d4280;
  wire v10d4281;
  wire v10d4282;
  wire v10d4283;
  wire v10d4284;
  wire v10d4285;
  wire v10d4286;
  wire v10d4287;
  wire v10d4288;
  wire v10d4289;
  wire v10d428a;
  wire v10d428b;
  wire v10d428c;
  wire v10d428d;
  wire v10d428e;
  wire v10d428f;
  wire v10d4290;
  wire v10d4291;
  wire v10d4292;
  wire v10d4293;
  wire v10d4294;
  wire v10d4295;
  wire v10d4296;
  wire v10d4297;
  wire v10d4298;
  wire v10d4299;
  wire v10d429a;
  wire v10d429b;
  wire v10d429c;
  wire v10d429d;
  wire v10d429e;
  wire v10d429f;
  wire v10d42a0;
  wire v10d42a1;
  wire v10d42a2;
  wire v10d42a3;
  wire v10d42a4;
  wire v10d42a5;
  wire v10d42a6;
  wire v10d42a7;
  wire v10d42a8;
  wire v10d42a9;
  wire v10d42aa;
  wire v10d42ae;
  wire v10d42af;
  wire v10d42b0;
  wire v10d42b1;
  wire v10d42b2;
  wire v10d42b3;
  wire v10d42b4;
  wire v10d42b5;
  wire v10d42b6;
  wire v10d42b7;
  wire v10d42b8;
  wire v10d42b9;
  wire v10d42ba;
  wire v10d42bb;
  wire v10d42bc;
  wire v10d42bd;
  wire v10d42be;
  wire v10d42bf;
  wire v10d42c0;
  wire v10d42c1;
  wire v10d42c2;
  wire v10d42c3;
  wire v10d42c4;
  wire v10d42c5;
  wire v10d42c6;
  wire v10d42c7;
  wire v10d42c8;
  wire v10d42c9;
  wire v10d42ca;
  wire v10d42cb;
  wire v10d42cc;
  wire v10d42cd;
  wire v10d42ce;
  wire v10d42cf;
  wire v10d42d0;
  wire v10d42d1;
  wire v10d42d2;
  wire v10d42d3;
  wire v10d42d4;
  wire v10d42d5;
  wire v10d42d6;
  wire v10d42d7;
  wire v10d42d8;
  wire v10d42d9;
  wire v10d42da;
  wire v10d42db;
  wire v10d42dc;
  wire v10d42dd;
  wire v10d42de;
  wire v10d42df;
  wire v10d42e0;
  wire v10d42e1;
  wire v10d4304;
  wire v10d4305;
  wire v84554c;
  wire v11ac602;
  wire v11ac67a;
  wire v11ac67b;
  wire v11ac67c;
  wire v11ac6a3;
  wire v11ac6c8;
  wire v11ac6c9;
  wire v11ac6ca;
  wire v845550;
  wire v845576;
  wire c50efb;
  wire c50efc;
  wire c50efd;
  wire c50efe;
  wire v84555c;
  wire v845568;
  wire b09421;
  wire v90d5cd;
  wire v85e75f;
  wire v9dde65;
  wire ae2496;
  wire v85e749;
  wire v11f33c5;
  wire v8b6f6c;
  wire v11f33c6;
  wire v11f3405;
  wire v845586;
  wire v155392f;
  wire v84556c;
  wire acd334;
  wire v1553930;
  wire v1553931;
  wire v1553932;
  wire v1553933;
  wire v1553934;
  wire v1553137;
  wire v1553138;
  wire v1553139;
  wire v155313a;
  wire v155313b;
  wire v155313c;
  wire v155313d;
  wire v155313e;
  wire v155313f;
  wire v1553140;
  wire v1553141;
  wire v1553142;
  wire v1553143;
  wire v1553144;
  wire v1553145;
  wire v1553146;
  wire v1553147;
  wire v1553148;
  wire v155314c;
  wire v155314d;
  wire v155314e;
  wire v155314f;
  wire v1553150;
  wire v1553151;
  wire v1553152;
  wire v1553153;
  wire v1553154;
  wire v1553155;
  wire v1553156;
  wire v1553157;
  wire v1553158;
  wire v1553215;
  wire v1553216;
  wire v1553217;
  wire v1553218;
  wire v1553219;
  wire v155321a;
  wire v155321b;
  wire v155321c;
  wire v155321d;
  wire v155321e;
  wire v155321f;
  wire v1553220;
  wire v1553221;
  wire v1553222;
  wire v1553223;
  wire v1553224;
  wire v1553225;
  wire v1553226;
  wire v1553227;
  wire v1553228;
  wire v1553229;
  wire v155322a;
  wire v155322b;
  wire v155322c;
  wire v155322d;
  wire v155322e;
  wire v155322f;
  wire v1553230;
  wire v1553231;
  wire v1553232;
  wire v1553233;
  wire v1553234;
  wire v1553235;
  wire v1553236;
  wire v1553237;
  wire v1553238;
  wire v1553239;
  wire v155323a;
  wire v15532be;
  wire v15532bf;
  wire v15532c1;
  wire v15532c2;
  wire v15532c3;
  wire v15532c4;
  wire v15532c5;
  wire v15532c6;
  wire v15532c7;
  wire v15532c8;
  wire v15532c9;
  wire v15532ca;
  wire v15532cb;
  wire v15532cc;
  wire v15532cd;
  wire v1553306;
  wire v155337f;
  wire v1553380;
  wire v1553381;
  wire v1553382;
  wire v1553383;
  wire v1553384;
  wire v1553385;
  wire v1553386;
  wire v1553387;
  wire v1553388;
  wire v1553389;
  wire v155338a;
  wire v155338b;
  wire v155338c;
  wire v155338d;
  wire v155338e;
  wire v155338f;
  wire v1553390;
  wire v1553391;
  wire v1553392;
  wire v1553393;
  wire v1553394;
  wire v1553395;
  wire v1553396;
  wire v1553397;
  wire v1553398;
  wire v1553399;
  wire v155339a;
  wire v155339b;
  wire v155339c;
  wire v155339d;
  wire v155339e;
  wire v155339f;
  wire v15533a0;
  wire v15533a1;
  wire v15533a2;
  wire v15533a3;
  wire v15533a4;
  wire v15533a5;
  wire v15533a6;
  wire v15533a7;
  wire v15533a8;
  wire v15533a9;
  wire v15533aa;
  wire v15533ab;
  wire v15533ac;
  wire v15533ad;
  wire v15533ae;
  wire v15533af;
  wire v15533b0;
  wire v15533b1;
  wire v15533b2;
  wire v15533b3;
  wire v15533b4;
  wire v15533b5;
  wire v15533b6;
  wire v15533b7;
  wire v15533b8;
  wire v1553412;
  wire v1553413;
  wire v1553414;
  wire v1553415;
  wire v1553416;
  wire v1553417;
  wire v1553418;
  wire v1553419;
  wire v155341a;
  wire v155341b;
  wire v155341c;
  wire v155341d;
  wire v155341e;
  wire v155341f;
  wire v1553420;
  wire v1553421;
  wire v1553422;
  wire v1553423;
  wire v1553424;
  wire v1553425;
  wire v1553426;
  wire v1553427;
  wire v1553428;
  wire v1553429;
  wire v155342a;
  wire v155342b;
  wire v155342c;
  wire v155342d;
  wire v155342e;
  wire v155342f;
  wire v1553430;
  wire v1553431;
  wire v1553432;
  wire v1553433;
  wire v1553434;
  wire v1553435;
  wire v1553436;
  wire v1553437;
  wire v1553438;
  wire v1553439;
  wire v155343a;
  wire v155343b;
  wire v155343c;
  wire v155343d;
  wire v155343e;
  wire v155343f;
  wire v1553440;
  wire v1553441;
  wire v1553442;
  wire v1553443;
  wire v1553444;
  wire v1553445;
  wire v1553446;
  wire v1553447;
  wire v1553448;
  wire v15534ce;
  wire v15534cf;
  wire v15534d0;
  wire v15534d1;
  wire v15534d2;
  wire v15534d3;
  wire v15534d4;
  wire v15534d5;
  wire v15534d6;
  wire v15534d7;
  wire v15534d8;
  wire v15534d9;
  wire v15534da;
  wire v15534db;
  wire v15534dc;
  wire v15534dd;
  wire v15534eb;
  wire v15534ec;
  wire v15534ed;
  wire v15534ee;
  wire v15534ef;
  wire v15534f0;
  wire v15534f1;
  wire v15534f2;
  wire v15534f3;
  wire v15534f4;
  wire v15534f5;
  wire v15534f6;
  wire v15534f7;
  wire v15534f8;
  wire v15534f9;
  wire v15534fa;
  wire v15534fb;
  wire v15534fc;
  wire v15534fd;
  wire v15534fe;
  wire v15534ff;
  wire v1553500;
  wire v1553501;
  wire v1553502;
  wire v1553503;
  wire v1553504;
  wire v1553505;
  wire v1553506;
  wire v1553507;
  wire v1553508;
  wire v1553509;
  wire v155350a;
  wire v155350b;
  wire v155350c;
  wire v155350d;
  wire v155350e;
  wire v155350f;
  wire v1553510;
  wire v1553511;
  wire v1553512;
  wire v1553513;
  wire v1553514;
  wire v1553515;
  wire v1553516;
  wire v1553517;
  wire v1553518;
  wire v1553519;
  wire v155351a;
  wire v155351b;
  wire v155351c;
  wire v1552d47;
  wire v1552d48;
  wire v1552d49;
  wire v1552d4a;
  wire v1552d4b;
  wire v1552d4c;
  wire v1552d4d;
  wire v1552d4e;
  wire v1552d51;
  wire v1552d52;
  wire v1552d53;
  wire v1552d54;
  wire v1552d55;
  wire v1552d56;
  wire v1552d57;
  wire v1552d58;
  wire v1552d59;
  wire v1552d5a;
  wire v1552d5b;
  wire v1552d5c;
  wire v1552d5d;
  wire v1552d5e;
  wire v1552d5f;
  wire v1552d60;
  wire v1552d61;
  wire v1552d62;
  wire v1552d63;
  wire v1552d64;
  wire v1552d65;
  wire v1552d66;
  wire v1552d67;
  wire v1552d68;
  wire v1552d69;
  wire v1552d6a;
  wire v1552d6b;
  wire v1552d6c;
  wire v1552d6d;
  wire v1552d6e;
  wire v1552d74;
  wire v1552d75;
  wire v1552d76;
  wire v1552d77;
  wire v1552d78;
  wire v1552d79;
  wire v1552d7a;
  wire v1552d7b;
  wire v1552d7c;
  wire v1552d7d;
  wire v1552d7e;
  wire v1552d7f;
  wire v1552d80;
  wire v1552d81;
  wire v1552d82;
  wire v1552d83;
  wire v1552d84;
  wire v1552d85;
  wire v1552d86;
  wire v1552d87;
  wire v1552d88;
  wire v1552d89;
  wire v1552d8a;
  wire v1552d8b;
  wire v1552d8c;
  wire v1552d8d;
  wire v1552d8e;
  wire v1552d8f;
  wire v1552d90;
  wire v1552d91;
  wire v1552d92;
  wire v1552d93;
  wire v1552d94;
  wire v1552d95;
  wire v1552d96;
  wire v1552d97;
  wire v1552d98;
  wire v1552d99;
  wire v1552d9a;
  wire v1552d9b;
  wire v1552d9c;
  wire v1552d9d;
  wire v1552d9e;
  wire v1552d9f;
  wire v1552da0;
  wire v1552da1;
  wire v1552da2;
  wire v1552da3;
  wire v1552f53;
  wire v1552f54;
  wire v1552f55;
  wire v1552f56;
  wire v1552f57;
  wire v1552f58;
  wire v1552f59;
  wire v1552f5a;
  wire v1552f5b;
  wire v1552f5c;
  wire v1552f5d;
  wire v1552f5e;
  wire v1552f5f;
  wire v1552f60;
  wire v1552f61;
  wire v1552f62;
  wire v1552f63;
  wire v1552f64;
  wire v1552f65;
  wire v1552f66;
  wire v1552f67;
  wire v1552f68;
  wire v1552f69;
  wire v1552f6a;
  wire v1552f6b;
  wire v1552f6c;
  wire v1552f6d;
  wire v1552f6e;
  wire v1552f6f;
  wire v1552f70;
  wire v1552f71;
  wire v1552f72;
  wire v1552f73;
  wire v1552f74;
  wire v1552f75;
  wire v1552f76;
  wire v1552f77;
  wire v1552f78;
  wire v1552f79;
  wire v1552f7a;
  wire v1552f7b;
  wire v1552f7c;
  wire v1552f7d;
  wire v1552f7e;
  wire v1552f7f;
  wire v1552f80;
  wire v1552f81;
  wire v1552f82;
  wire v1552f83;
  wire v1552f84;
  wire v1552f85;
  wire v1552f86;
  wire v1552f87;
  wire v1552f88;
  wire v1552f89;
  wire v1552f8a;
  wire v1552f8b;
  wire v1552f8c;
  wire v1552f8d;
  wire v1552fcb;
  wire v1552fcc;
  wire v1552fcd;
  wire v1552fce;
  wire v1552fcf;
  wire v1552fd0;
  wire v1552fd1;
  wire v1552fd2;
  wire v1552fd3;
  wire v1552fd4;
  wire v1552fd5;
  wire v1552fd6;
  wire v1552fd7;
  wire v1552fd8;
  wire v155304c;
  wire v155304d;
  wire v155304e;
  wire v155304f;
  wire v1553050;
  wire v1553051;
  wire v1553052;
  wire v1553053;
  wire v1553054;
  wire v1553055;
  wire v1553056;
  wire v1553057;
  wire v1553058;
  wire v1553059;
  wire v155305a;
  wire v155305b;
  wire v155305c;
  wire v155305d;
  wire v155305e;
  wire v155305f;
  wire v1553060;
  wire v1553061;
  wire v1553089;
  wire v155308a;
  wire v155308b;
  wire v155308c;
  wire v155308d;
  wire v155308e;
  wire v155308f;
  wire v1553090;
  wire v1553091;
  wire v1553092;
  wire v1553093;
  wire v1553094;
  wire v1553095;
  wire v1553096;
  wire v1553097;
  wire v1553098;
  wire v1553099;
  wire v155309a;
  wire v155309b;
  wire v155309c;
  wire v155309d;
  wire v155309e;
  wire v155309f;
  wire v15530a0;
  wire v15530a1;
  wire v15530a2;
  wire v15530a3;
  wire v15530a4;
  wire v15530a5;
  wire v15530a6;
  wire v15530a7;
  wire v15530a8;
  wire v15530a9;
  wire v15530aa;
  wire v15530ab;
  wire v15530ac;
  wire v15530ad;
  wire v15530ae;
  wire v15530af;
  wire v15530b0;
  wire v15530b1;
  wire v15530b2;
  wire v15530b3;
  wire v15530b4;
  wire v15530b5;
  wire v15530b6;
  wire v15530b7;
  wire v15530e8;
  wire v15530e9;
  wire v15530ea;
  wire v15530eb;
  wire v15530ec;
  wire v15530ed;
  wire v15530ee;
  wire v15530ef;
  wire v15530f0;
  wire v15530f1;
  wire v15530f2;
  wire v15530f3;
  wire v15530f4;
  wire v15530f5;
  wire v15530fd;
  wire v15530fe;
  wire v15530ff;
  wire v1553100;
  wire v1553101;
  wire v1553102;
  wire v1553103;
  wire v1553104;
  wire v1553105;
  wire v1553106;
  wire v1552960;
  wire v1552961;
  wire v1552962;
  wire v1552963;
  wire v155298b;
  wire v155298c;
  wire v155298d;
  wire v155298e;
  wire v155298f;
  wire v1552990;
  wire v845564;
  wire v10a153f;
  wire v845574;
  wire v10a1540;
  wire v10a1541;
  wire v10a1542;
  wire v10a1543;
  wire a81304;
  wire v87abb5;
  wire v8dfa41;
  wire v86ab0d;
  wire v936735;
  wire d80730;
  wire d80731;
  wire d80732;
  wire d80733;
  wire d80734;
  wire d80735;
  wire d80736;
  wire d80737;
  wire d80738;
  wire v8b8a8c;
  wire d80739;
  wire d8073a;
  wire d8073b;
  wire d8073c;
  wire d8073d;
  wire d8073e;
  wire d8073f;
  wire d80740;
  wire d80741;
  wire d80742;
  wire d80743;
  wire d80744;
  wire d80745;
  wire d80746;
  wire d80747;
  wire d80748;
  wire d80749;
  wire d8074a;
  wire d8074b;
  wire d8074c;
  wire d8074d;
  wire d8074e;
  wire d8074f;
  wire d80750;
  wire d80751;
  wire d80752;
  wire d80753;
  wire d80754;
  wire d80755;
  wire d80756;
  wire d80757;
  wire d80758;
  wire d80759;
  wire d8075a;
  wire d8075b;
  wire d8075c;
  wire d8075d;
  wire d8075e;
  wire d8075f;
  wire d80760;
  wire d80761;
  wire d80762;
  wire d80763;
  wire d80764;
  wire d80765;
  wire d80766;
  wire d80767;
  wire d80768;
  wire d80769;
  wire d8076a;
  wire d8076b;
  wire d8076c;
  wire d8076d;
  wire d8076e;
  wire d8076f;
  wire d80770;
  wire d80771;
  wire d80772;
  wire d80773;
  wire d80774;
  wire d80775;
  wire d80776;
  wire d80777;
  wire d80778;
  wire d80779;
  wire d8077a;
  wire d8077b;
  wire d8077c;
  wire d8077d;
  wire d8077e;
  wire d8077f;
  wire d80780;
  wire d80781;
  wire d80782;
  wire d80783;
  wire d80784;
  wire d80785;
  wire d80786;
  wire d80787;
  wire d80788;
  wire d80789;
  wire d8078a;
  wire d8078b;
  wire d8078c;
  wire d8078d;
  wire d8078e;
  wire d8078f;
  wire d80790;
  wire d80791;
  wire d80792;
  wire d80793;
  wire d80794;
  wire d80795;
  wire d80796;
  wire d80797;
  wire d80798;
  wire d80799;
  wire d8079a;
  wire d8079b;
  wire d8079c;
  wire d8079d;
  wire d8079e;
  wire d8079f;
  wire d807a0;
  wire d807a1;
  wire d807a2;
  wire d807a3;
  wire d807a4;
  wire d807a5;
  wire d807a6;
  wire d807a7;
  wire d807a8;
  wire d807a9;
  wire d807aa;
  wire d807ab;
  wire d807ac;
  wire d807ad;
  wire d807ae;
  wire d807af;
  wire d807b0;
  wire d807b1;
  wire d807b2;
  wire d807b3;
  wire d807b4;
  wire d807b5;
  wire d807b6;
  wire d807b7;
  wire d807b8;
  wire d807b9;
  wire d807ba;
  wire d807bb;
  wire d807bc;
  wire d807bd;
  wire d807be;
  wire d807bf;
  wire d807c0;
  wire v893df7;
  wire v8a9c96;
  wire v906a5a;
  wire v156645f;
  wire a66272;
  wire a66273;
  wire a66275;
  wire a66276;
  wire a66278;
  wire a6627a;
  wire v84556a;
  wire a6627b;
  wire a6627c;
  wire a6627d;
  wire a6627e;
  wire a6627f;
  wire a66280;
  wire a66281;
  wire v845570;
  wire a66283;
  wire a66284;
  wire a66285;
  wire a66286;
  wire a66287;
  wire a66289;
  wire a6628b;
  wire a6628c;
  wire a6628e;
  wire a6628f;
  wire a66290;
  wire a66291;
  wire a66292;
  wire a66293;
  wire a66294;
  wire a66295;
  wire a66296;
  wire a66297;
  wire a66298;
  wire a66299;
  wire a6629a;
  wire a6629b;
  wire a6629c;
  wire a6629d;
  wire a6629e;
  wire a6629f;
  wire v84557a;
  wire a662a0;
  wire a662a1;
  wire a662a2;
  wire a662a3;
  wire a662a4;
  wire a662a6;
  wire a662a7;
  wire a662a9;
  wire a662aa;
  wire a662ab;
  wire a662ac;
  wire a662ad;
  wire a662ae;
  wire a662b2;
  wire a662b4;
  wire a662b7;
  wire a662b8;
  wire a662b9;
  wire a662ba;
  wire a662bb;
  wire a662bc;
  wire a662bd;
  wire a662be;
  wire a662c0;
  wire a662c1;
  wire a662c2;
  wire a662c3;
  wire a662c5;
  wire a662c6;
  wire a662c7;
  wire a662ca;
  wire a662cb;
  wire a662cc;
  wire a662cd;
  wire a662cf;
  wire a662d0;
  wire a662d2;
  wire a65ad6;
  wire a65ad7;
  wire a65ada;
  wire a65adb;
  wire a65adc;
  wire a65add;
  wire a65ae0;
  wire a65ae1;
  wire a65ae2;
  wire a65ae4;
  wire a65ae5;
  wire a65ae6;
  wire a65ae7;
  wire a65ae8;
  wire a65ae9;
  wire a65aea;
  wire a65aeb;
  wire a65aed;
  wire a65aee;
  wire a65af0;
  wire a65af1;
  wire a65af2;
  wire a65af3;
  wire a65af4;
  wire a65af5;
  wire a65af6;
  wire a65af7;
  wire a65af8;
  wire a65af9;
  wire a65afe;
  wire a65aff;
  wire a65b06;
  wire a65b07;
  wire a65b09;
  wire a65b0a;
  wire a65b0d;
  wire a65b12;
  wire a65b13;
  wire a65b14;
  wire a65b17;
  wire a65b18;
  wire a65b19;
  wire a65b1a;
  wire a65b20;
  wire a65b21;
  wire a65b23;
  wire a65b25;
  wire a65b26;
  wire a65b27;
  wire a65b28;
  wire a65b29;
  wire a65b2b;
  wire a65b2c;
  wire a65b2e;
  wire a65b2f;
  wire a65b30;
  wire a65b31;
  wire a65b32;
  wire a65b38;
  wire a65b3a;
  wire a65b3b;
  wire a65b3c;
  wire a65b3d;
  wire a65b3f;
  wire a65b40;
  wire a65851;
  wire a65852;
  wire a65853;
  wire a65854;
  wire a65856;
  wire a65857;
  wire a65858;
  wire a65859;
  wire a6585b;
  wire a6585c;
  wire a6585d;
  wire a6585e;
  wire a6585f;
  wire a65861;
  wire a65862;
  wire a65863;
  wire a65864;
  wire a65866;
  wire a65867;
  wire a65869;
  wire a6586a;
  wire a6586b;
  wire a6586c;
  wire a6586d;
  wire a6586e;
  wire a65873;
  wire a65878;
  wire a65879;
  wire a6587a;
  wire a6587b;
  wire a6587e;
  wire a6587f;
  wire a65883;
  wire a65884;
  wire a65885;
  wire a65886;
  wire a65888;
  wire a6588a;
  wire a6588d;
  wire a6588f;
  wire a65890;
  wire a65891;
  wire a65892;
  wire a65893;
  wire a65894;
  wire a65896;
  wire a65898;
  wire v9a051b;
  wire a658a3;
  wire a658a5;
  wire a658a7;
  wire v8af912;
  wire afe156;
  wire a658a8;
  wire a658a9;
  wire a658aa;
  wire a658ab;
  wire a658ac;
  wire a658ad;
  wire a658b0;
  wire ab8d68;
  wire a658b2;
  wire a658b3;
  wire a658b4;
  wire a658b5;
  wire a658b6;
  wire a658b7;
  wire a67ea5;
  wire v9f3194;
  wire v110b6cc;
  wire a658ba;
  wire a658bb;
  wire a658bc;
  wire a658bd;
  wire a658be;
  wire a658bf;
  wire a658c1;
  wire a658c3;
  wire a658c6;
  wire a658c7;
  wire a658c8;
  wire a658c9;
  wire a658ca;
  wire a658cb;
  wire a658cc;
  wire a658ce;
  wire a658cf;
  wire a658d0;
  wire a658d1;
  wire a658d2;
  wire a658d3;
  wire a658d4;
  wire a658d5;
  wire a658d6;
  wire a658d7;
  wire a658d8;
  wire a658da;
  wire a658db;
  wire a658dc;
  wire a658de;
  wire a658e0;
  wire a658e1;
  wire a658e2;
  wire a658e3;
  wire a658e5;
  wire a658e7;
  wire a658e8;
  wire a658ea;
  wire a658eb;
  wire a658ed;
  wire a658ee;
  wire a658ef;
  wire a658f0;
  wire a658f1;
  wire a658f2;
  wire a658f4;
  wire a658f6;
  wire a658f9;
  wire a658fb;
  wire a658fc;
  wire a658fd;
  wire a658fe;
  wire a658ff;
  wire a65909;
  wire a6590b;
  wire a6590e;
  wire a6590f;
  wire a65910;
  wire a65911;
  wire a65912;
  wire a65913;
  wire a65915;
  wire a65916;
  wire a65917;
  wire a65919;
  wire a6591b;
  wire a6591c;
  wire a6591e;
  wire a6591f;
  wire a65920;
  wire a65921;
  wire a65922;
  wire a65923;
  wire a65924;
  wire a65925;
  wire a65926;
  wire a65927;
  wire a65928;
  wire a65929;
  wire a6592a;
  wire a6592b;
  wire a6535b;
  wire a6535d;
  wire a6535e;
  wire a65360;
  wire v845558;
  wire a65361;
  wire a65362;
  wire a65363;
  wire a65364;
  wire a65365;
  wire a65366;
  wire a65367;
  wire a65368;
  wire a65369;
  wire a6536d;
  wire a6536e;
  wire a65370;
  wire a65371;
  wire a65372;
  wire a65376;
  wire a65377;
  wire a65378;
  wire a65379;
  wire a6537a;
  wire a6537b;
  wire a6537d;
  wire a6537e;
  wire a6537f;
  wire a65380;
  wire a65381;
  wire a65382;
  wire a65384;
  wire a65387;
  wire a65389;
  wire a6538a;
  wire a6538b;
  wire a6538d;
  wire a6538e;
  wire a6538f;
  wire a65390;
  wire a65391;
  wire a65392;
  wire a65393;
  wire a65394;
  wire a65395;
  wire a65396;
  wire a65399;
  wire a6539a;
  wire a6539b;
  wire a653a1;
  wire a653a2;
  wire a653a3;
  wire a653a7;
  wire a653a8;
  wire a653a9;
  wire a653aa;
  wire a653ab;
  wire a653ac;
  wire a653ad;
  wire a653ae;
  wire a653b4;
  wire a653b5;
  wire a653b6;
  wire a653b7;
  wire a653b8;
  wire a653b9;
  wire a653ba;
  wire a653bb;
  wire a653bc;
  wire a653bd;
  wire a653bf;
  wire a653c0;
  wire a653c2;
  wire a653c3;
  wire a653c4;
  wire a653c5;
  wire a653c6;
  wire a653c7;
  wire a653c8;
  wire a653c9;
  wire a653cb;
  wire a653cc;
  wire a653cd;
  wire a653cf;
  wire a653d0;
  wire a653d1;
  wire a653d3;
  wire a653d4;
  wire a653d5;
  wire a653d6;
  wire a653d7;
  wire a653d8;
  wire a653d9;
  wire a653da;
  wire a653dc;
  wire a653dd;
  wire a653de;
  wire a653df;
  wire a653e0;
  wire a653e2;
  wire a653e3;
  wire a653e4;
  wire a653e5;
  wire a653e6;
  wire a653e7;
  wire a653e8;
  wire a653e9;
  wire a653ea;
  wire a653ec;
  wire a653ed;
  wire a653ef;
  wire a653f0;
  wire a653f3;
  wire a653f4;
  wire a653f5;
  wire a653f8;
  wire a653f9;
  wire a653fa;
  wire a653fc;
  wire a653fd;
  wire a653fe;
  wire a653ff;
  wire a65400;
  wire a65401;
  wire a65403;
  wire a65405;
  wire a65407;
  wire a65408;
  wire a65409;
  wire a6540a;
  wire a6540b;
  wire a6540c;
  wire a6540d;
  wire v949cd9;
  wire a1db63;
  wire a6540e;
  wire a6540f;
  wire a65410;
  wire a65412;
  wire a65414;
  wire a65416;
  wire a65418;
  wire a65419;
  wire a6541b;
  wire a6541d;
  wire a6541e;
  wire a6541f;
  wire a65422;
  wire a65424;
  wire a65426;
  wire a65427;
  wire a65429;
  wire a6542b;
  wire a6542d;
  wire a6542e;
  wire a6542f;
  wire a65431;
  wire a65433;
  wire a65434;
  wire a65436;
  wire a65437;
  wire a65438;
  wire a65439;
  wire a6543a;
  wire a6543c;
  wire a6543d;
  wire a6543e;
  wire a6543f;
  wire a65440;
  wire a65441;
  wire a65443;
  wire a65444;
  wire a65445;
  wire a65446;
  wire a65449;
  wire a6544b;
  wire a6544c;
  wire a65450;
  wire a65451;
  wire a65452;
  wire a65454;
  wire a65455;
  wire a65456;
  wire a65457;
  wire a65458;
  wire a65459;
  wire a6545a;
  wire a6545b;
  wire a6545c;
  wire a6545d;
  wire a65460;
  wire a65461;
  wire a65463;
  wire a65464;
  wire a65465;
  wire v1566987;
  wire a65466;
  wire a65467;
  wire a65468;
  wire a65469;
  wire a6546a;
  wire a6546c;
  wire a6546d;
  wire a6546f;
  wire a65470;
  wire a65471;
  wire a65472;
  wire a65473;
  wire a65474;
  wire a65475;
  wire a65476;
  wire a65478;
  wire a65479;
  wire a6548a;
  wire a6548b;
  wire a6548c;
  wire a6548d;
  wire a6548f;
  wire a65490;
  wire a65491;
  wire a65492;
  wire a65493;
  wire a65494;
  wire a65495;
  wire a65496;
  wire a65498;
  wire a65499;
  wire a6549a;
  wire a6549b;
  wire a654a9;
  wire a654ab;
  wire a654ac;
  wire a654ad;
  wire a654ae;
  wire a654af;
  wire a654b0;
  wire a654b1;
  wire a654b2;
  wire a654b4;
  wire a654b5;
  wire a654b6;
  wire a654b8;
  wire a654b9;
  wire a654ba;
  wire a654bb;
  wire a654bc;
  wire a654bd;
  wire a654be;
  wire a654c0;
  wire a654c3;
  wire a654c5;
  wire a654c6;
  wire a654c9;
  wire a654cb;
  wire a65613;
  wire a65614;
  wire a65615;
  wire a65616;
  wire a65619;
  wire a6561a;
  wire a6561c;
  wire a6561d;
  wire a6561f;
  wire a65620;
  wire a65621;
  wire a65622;
  wire a65623;
  wire a65624;
  wire a65625;
  wire a65626;
  wire a65627;
  wire a65628;
  wire a6562a;
  wire a6562c;
  wire a6562d;
  wire a6562e;
  wire a65630;
  wire a65632;
  wire a65634;
  wire a65635;
  wire a65636;
  wire a65637;
  wire a65638;
  wire a65639;
  wire a6563a;
  wire a6563b;
  wire a6563c;
  wire a6563e;
  wire a6563f;
  wire a65640;
  wire a65643;
  wire a65644;
  wire a65645;
  wire a65646;
  wire a65647;
  wire a65648;
  wire a6564a;
  wire a6564b;
  wire a6564c;
  wire a6564d;
  wire a6564e;
  wire a6564f;
  wire a65650;
  wire a65652;
  wire a65653;
  wire a65655;
  wire a65656;
  wire a65658;
  wire a6565a;
  wire a6565c;
  wire a6565f;
  wire a65661;
  wire a65663;
  wire a65665;
  wire a65666;
  wire a65667;
  wire a65669;
  wire a6566a;
  wire a6566b;
  wire a6566c;
  wire a6566d;
  wire a6566e;
  wire a6566f;
  wire a65670;
  wire a65671;
  wire a65672;
  wire a65674;
  wire a65676;
  wire a65677;
  wire a65678;
  wire a6567a;
  wire a6567b;
  wire a6567c;
  wire a6567d;
  wire a6567e;
  wire a6567f;
  wire a65680;
  wire a65681;
  wire a65682;
  wire a65684;
  wire a65685;
  wire a65686;
  wire a65687;
  wire a65688;
  wire a6568a;
  wire a6568b;
  wire a6568d;
  wire a6568e;
  wire a6568f;
  wire a65690;
  wire a65691;
  wire a65692;
  wire a65693;
  wire a65698;
  wire a65699;
  wire a6569a;
  wire a6569c;
  wire a6569e;
  wire a656a0;
  wire a656a1;
  wire a656a2;
  wire a656a3;
  wire a656a4;
  wire a656a5;
  wire a656a9;
  wire a656ab;
  wire a656ac;
  wire a656ad;
  wire a656ae;
  wire a656b0;
  wire a656b1;
  wire a656b2;
  wire a656b4;
  wire a656b6;
  wire a656b8;
  wire a656b9;
  wire a656bc;
  wire a656bd;
  wire a656be;
  wire a656c0;
  wire a656c1;
  wire a656c2;
  wire a656c3;
  wire a656c4;
  wire a656c5;
  wire a656c8;
  wire a656c9;
  wire a656ca;
  wire a656cb;
  wire a656cd;
  wire a656ce;
  wire a656cf;
  wire a656d0;
  wire a656d1;
  wire a656d2;
  wire a656d3;
  wire a646d8;
  wire a646d9;
  wire a646da;
  wire a646db;
  wire a646dc;
  wire a64704;
  wire a64705;
  wire a64707;
  wire a64708;
  wire a64709;
  wire a6470a;
  wire a6470b;
  wire a6470c;
  wire a6470d;
  wire a6470e;
  wire a6470f;
  wire a64712;
  wire a64713;
  wire a64714;
  wire a64715;
  wire a64716;
  wire a64717;
  wire a64719;
  wire v1668c17;
  wire v1668c18;
  wire v1668c19;
  wire v1668c1a;
  wire v1668c1b;
  wire v1668c1c;
  wire v1668c1d;
  wire v1668c1e;
  wire v1668c1f;
  wire v1668c20;
  wire v1668c21;
  wire v1668c22;
  wire v1668c23;
  wire v1668c24;
  wire v1668c25;
  wire v1668c26;
  wire v1668c27;
  wire v1668c28;
  wire v1668c29;
  wire v1668c2a;
  wire v1668c2b;
  wire v1668c2c;
  wire v1668c2d;
  wire v1668c2e;
  wire v1668c2f;
  wire v1668c30;
  wire v1668c31;
  wire v1668c32;
  wire v1668c33;
  wire v1668c34;
  wire v1668c35;
  wire v1668c36;
  wire v1668c37;
  wire v1668c38;
  wire v84556e;
  wire v1668c39;
  wire v1668c3a;
  wire v1668c3b;
  wire v1668c3c;
  wire v1668c3d;
  wire v1668c3e;
  wire v1668c3f;
  wire v1668c40;
  wire v1668c41;
  wire v1668c42;
  wire v1668c43;
  wire v1668c44;
  wire v1668c45;
  wire v1668c46;
  wire v1668c47;
  wire v1668c48;
  wire v1668c49;
  wire v1668c4a;
  wire v1668c4b;
  wire v1668c4c;
  wire v1668c4d;
  wire v1668c4e;
  wire v1668c4f;
  wire v1668c50;
  wire v1668c51;
  wire v1668c52;
  wire v1668c53;
  wire v1668c54;
  wire v1668c55;
  wire v1668c56;
  wire v1668c57;
  wire v1668c58;
  wire v1668c59;
  wire v1668c5a;
  wire v1668c5b;
  wire v1668c5f;
  wire v1668c60;
  wire v1668c61;
  wire v1668c62;
  wire v1668c63;
  wire v1668c64;
  wire v1668c65;
  wire v1668c66;
  wire v1668c67;
  wire v960a34;
  wire v92fc87;
  wire ab83a0;
  wire v1668c68;
  wire v1668c69;
  wire v1668c6a;
  wire v1668c6b;
  wire v1668c6c;
  wire v1668c6d;
  wire v1668c6e;
  wire v1668c6f;
  wire v1668c70;
  wire v1668c71;
  wire v1668c72;
  wire v1668c73;
  wire v1668c74;
  wire v1668c75;
  wire v1668c76;
  wire v1668c77;
  wire v1668c78;
  wire v1668c79;
  wire v1668c7a;
  wire v1668c7b;
  wire v1668c7c;
  wire v1668c7d;
  wire v1668c7e;
  wire v1668c81;
  wire v1668c82;
  wire v1668c83;
  wire v1668c86;
  wire v1668c87;
  wire v1668c88;
  wire v1668c89;
  wire v1668c8a;
  wire v1668c8b;
  wire v1668c8c;
  wire v1668c8d;
  wire v1668c8e;
  wire v1668c8f;
  wire v9337f3;
  wire a7c7c1;
  wire v1668c95;
  wire v1668c99;
  wire v1668c9a;
  wire v1668c9b;
  wire v1668c9c;
  wire v1668c9d;
  wire v1668c9e;
  wire v1668c9f;
  wire v1668ca0;
  wire v1668ca1;
  wire v1668ca2;
  wire v1668ca5;
  wire v1668ca6;
  wire v1668ca7;
  wire v1668caa;
  wire v1668cab;
  wire v1668cac;
  wire v1668cad;
  wire v1668cae;
  wire v1668caf;
  wire v1668cb5;
  wire v1668cb6;
  wire v1668cba;
  wire v1668cbb;
  wire v1668cbc;
  wire v1668cbd;
  wire v1668cbe;
  wire v1668cbf;
  wire v1668cc0;
  wire v1668cc1;
  wire v1668cc2;
  wire v1668cc3;
  wire v1668cc4;
  wire v1668cc5;
  wire v1668cc6;
  wire v1668cc7;
  wire v1668cc8;
  wire v1668cc9;
  wire v1668cca;
  wire v1668ccb;
  wire v1668ccc;
  wire v1668ccd;
  wire v1668cce;
  wire v1668ccf;
  wire v1668cd0;
  wire v1668cd1;
  wire v1668cd2;
  wire v1668cd3;
  wire v1668cd4;
  wire v1668cd5;
  wire v1668cd6;
  wire v1668cd7;
  wire v1668cd8;
  wire v1668cd9;
  wire v1668cda;
  wire v1668cdb;
  wire v1668cdc;
  wire v1668cdd;
  wire v1668cde;
  wire v1668cdf;
  wire v1668ce0;
  wire v1668ce1;
  wire v1668ce2;
  wire v1668ce3;
  wire v1668ce4;
  wire v1668ce5;
  wire v1668ce6;
  wire v1668ce7;
  wire v1668cea;
  wire v1668ceb;
  wire v1668cec;
  wire v1668cf0;
  wire v1668cf1;
  wire v1668cf2;
  wire v1668cf5;
  wire v1668cf6;
  wire v1668cf7;
  wire v1668cfb;
  wire v1668cfc;
  wire v1668cfd;
  wire v1668cfe;
  wire v1668cff;
  wire v1668d00;
  wire v1668d01;
  wire v1668d02;
  wire v1668d05;
  wire v1668d06;
  wire v1668d07;
  wire v1668d0b;
  wire v1668d0e;
  wire v1668d0f;
  wire v1668d10;
  wire v1668d11;
  wire v1668d12;
  wire v1668d13;
  wire v1668d14;
  wire v1668d15;
  wire v1668d16;
  wire v1668d17;
  wire v1668d18;
  wire v1668d19;
  wire v1668d1a;
  wire v1668d1b;
  wire v1668d1c;
  wire v1668d1d;
  wire v1668d1e;
  wire v1668d1f;
  wire v1668d21;
  wire v1668d22;
  wire v1668d23;
  wire v1668d24;
  wire v1668d25;
  wire v1668d26;
  wire v1668d27;
  wire v1668d28;
  wire v1668d29;
  wire v1668d2a;
  wire v1668d2b;
  wire v1668d2c;
  wire v1668d2d;
  wire v1668d2e;
  wire v1668d2f;
  wire v1668d30;
  wire v1668d31;
  wire v1668d32;
  wire v1668d33;
  wire v1668d34;
  wire v1668d35;
  wire v1668d36;
  wire v1668d37;
  wire v1668d38;
  wire v1668d39;
  wire v1668d3a;
  wire v1668d3b;
  wire v1668d3c;
  wire v1668d3d;
  wire v1668d3e;
  wire v1668d3f;
  wire v1668d40;
  wire v1668d41;
  wire v1668d42;
  wire v1668d43;
  wire v1668d44;
  wire v1668d45;
  wire v1668d46;
  wire v1668d47;
  wire v1668d48;
  wire v1668d49;
  wire v1668d4a;
  wire v1668d4b;
  wire v1668d4c;
  wire v1668d4d;
  wire v1668d4e;
  wire v1668d4f;
  wire v1668d50;
  wire v1668d51;
  wire v1668d52;
  wire v1668d53;
  wire v1668d54;
  wire v1668d55;
  wire v1668d56;
  wire v1668d57;
  wire v1668d58;
  wire v1668d59;
  wire v1668d5a;
  wire v1668d5b;
  wire v1668d5c;
  wire v1668d5d;
  wire v1668d5e;
  wire v1668d5f;
  wire v1668d60;
  wire v1668d61;
  wire v1668d62;
  wire v1668d63;
  wire v1668d64;
  wire v1668d65;
  wire v1668d66;
  wire v1668d67;
  wire v1668d68;
  wire v1668d69;
  wire v1668d6a;
  wire v1668d6b;
  wire v1668d6c;
  wire v1668d6d;
  wire v1668d6e;
  wire v1668d6f;
  wire v1668d70;
  wire v1668d71;
  wire v1668d72;
  wire v1668d73;
  wire v1668d74;
  wire v1668d75;
  wire v1668d76;
  wire v1668d77;
  wire v1668d78;
  wire v1668d79;
  wire v1668d7a;
  wire v1668d7b;
  wire v1668d7c;
  wire v1668d7d;
  wire v1668d7e;
  wire v1668d7f;
  wire v1668d80;
  wire v1668d81;
  wire v1668d82;
  wire v1668d83;
  wire v1668d84;
  wire v1668d85;
  wire v1668d86;
  wire v1668d87;
  wire v1668d88;
  wire v1668d89;
  wire v1668d8a;
  wire v1668d8b;
  wire v1668d8c;
  wire v1668d8d;
  wire v1668d8e;
  wire v1668d8f;
  wire v1668d90;
  wire v1668d91;
  wire v1668d92;
  wire v1668d93;
  wire v1668d94;
  wire v1668d97;
  wire v1668d98;
  wire v1668d99;
  wire v1668d9a;
  wire v1668d9b;
  wire v1668d9c;
  wire v1668d9d;
  wire v1668d9e;
  wire v1668d9f;
  wire v1668da0;
  wire v1668da1;
  wire v1668da2;
  wire v1668da3;
  wire v1668da4;
  wire v1668da5;
  wire v1668da6;
  wire v1668da7;
  wire v1668da8;
  wire v1668da9;
  wire v1668daa;
  wire v1668dab;
  wire v1668dac;
  wire v1668dad;
  wire v1668dae;
  wire v1668daf;
  wire v1668db0;
  wire v1668db1;
  wire v1668db3;
  wire v1668db4;
  wire v1668db5;
  wire v1668db6;
  wire v1668db7;
  wire v1668db8;
  wire v1668db9;
  wire v1668dba;
  wire v1668dbb;
  wire v1668dbc;
  wire v1668dbd;
  wire v1668dbe;
  wire v1668dbf;
  wire v1668dc0;
  wire v1668dc1;
  wire v1668dc2;
  wire v1668dc3;
  wire v1668dc4;
  wire v1668dc5;
  wire v1668dc6;
  wire v1668dc7;
  wire v1668dc8;
  wire v1668dc9;
  wire v1668dca;
  wire v1668dcb;
  wire v1668dcc;
  wire v1668dcd;
  wire v1668dce;
  wire v1668dcf;
  wire v1668dd0;
  wire v1668dd1;
  wire v1668dd2;
  wire v1668dd3;
  wire v1668dd4;
  wire v1668dd7;
  wire v1668dd8;
  wire v1668dd9;
  wire v1668dda;
  wire v1668ddb;
  wire v1668ddc;
  wire v1668ddd;
  wire v1668dde;
  wire v1668ddf;
  wire v1668de0;
  wire v1668de1;
  wire v1668de2;
  wire v1668de3;
  wire v1668de4;
  wire v1668de5;
  wire v1668de6;
  wire v1668de7;
  wire v1668de8;
  wire v1668e01;
  wire v1668e02;
  wire v1668e03;
  wire v1668e04;
  wire v1668e05;
  wire v1668e06;
  wire v1668e07;
  wire v1668e08;
  wire v1668e09;
  wire v1668e0a;
  wire v1668e0b;
  wire v1668e0c;
  wire v1668e0d;
  wire v1668e0e;
  wire v1668e0f;
  wire v1668e10;
  wire v166939b;
  wire v166939c;
  wire v166939d;
  wire v166939e;
  wire v166939f;
  wire v16693a0;
  wire v16693a1;
  wire v16693a2;
  wire v16693a3;
  wire v16693a4;
  wire v16693a5;
  wire v16693a6;
  wire v16693a7;
  wire v16693a8;
  wire v16693a9;
  wire v16693aa;
  wire v16693ab;
  wire v16693ac;
  wire v16693ad;
  wire v16693ae;
  wire v16693af;
  wire v16693b0;
  wire v16693b1;
  wire v16693b2;
  wire v1669591;
  wire v1669592;
  wire v1669593;
  wire v1669594;
  wire v1669595;
  wire v1669596;
  wire v1669598;
  wire v1669599;
  wire v166959a;
  wire v166959b;
  wire v166959c;
  wire v166959d;
  wire v166959e;
  wire v166959f;
  wire v16695a0;
  wire v16695a1;
  wire v16695a2;
  wire v16695a3;
  wire v16695a4;
  wire v16695a5;
  wire v16695a6;
  wire v16695a7;
  wire v16695a8;
  wire v16695a9;
  wire v16695aa;
  wire v16695ab;
  wire v16695ac;
  wire v16695ad;
  wire v16695ae;
  wire v16695af;
  wire v16695b0;
  wire v16695b1;
  wire v16695b2;
  wire v16695b9;
  wire v16695ba;
  wire v16695bb;
  wire v16695bc;
  wire v16695bd;
  wire v16695c4;
  wire v16695c5;
  wire v16695c6;
  wire v16695c7;
  wire v16695c8;
  wire v16695c9;
  wire v16695ca;
  wire v1446394;
  wire v1446395;
  wire v1446396;
  wire v1446397;
  wire v1446398;
  wire v1446399;
  wire v144639a;
  wire v144639b;
  wire v845588;
  wire v146d169;
  wire v144639c;
  wire v144639d;
  wire v144639e;
  wire v144639f;
  wire v14463a0;
  wire v14463a1;
  wire v14463a2;
  wire v14463a3;
  wire v14463a4;
  wire v14463a5;
  wire v14463a6;
  wire v14463a7;
  wire v14463a8;
  wire v14463a9;
  wire v14463aa;
  wire v14463ab;
  wire v14463ac;
  wire v14463ad;
  wire v14463b1;
  wire v14463b2;
  wire v14463b3;
  wire v14463b4;
  wire v14463b5;
  wire v14463b6;
  wire v14463b7;
  wire v14463b8;
  wire v14463b9;
  wire v14463ba;
  wire v14463bb;
  wire v14463bc;
  wire v14463bd;
  wire v14463be;
  wire v14463bf;
  wire v14463c0;
  wire v14463c1;
  wire v14463c2;
  wire v14463c3;
  wire v14463c4;
  wire v14463c5;
  wire v14463c6;
  wire v14463c7;
  wire v14463c8;
  wire v14463c9;
  wire v14463ca;
  wire v14463cb;
  wire v14463cc;
  wire v14463cd;
  wire v14463ce;
  wire v14463cf;
  wire v14463d0;
  wire v14463d1;
  wire v14463d2;
  wire v14463d3;
  wire v14463d4;
  wire v14463d5;
  wire v14463d6;
  wire v14463d7;
  wire v14463d8;
  wire v14463d9;
  wire v14463da;
  wire v14463db;
  wire v14463dc;
  wire v14463dd;
  wire v14463de;
  wire v14463df;
  wire v14463e0;
  wire v14463e1;
  wire v14463e2;
  wire v14463e3;
  wire v14463e4;
  wire v14463e5;
  wire v14463e6;
  wire v14463e7;
  wire v14463e8;
  wire v14463e9;
  wire v14463ea;
  wire v14463eb;
  wire v14463ec;
  wire v14463ed;
  wire v14463ee;
  wire v14463ef;
  wire v14463f0;
  wire v14463f1;
  wire v14463f2;
  wire v14463f3;
  wire v14463f4;
  wire v14463f5;
  wire v14463f6;
  wire v14463f7;
  wire v14463f8;
  wire v14463f9;
  wire v14463fa;
  wire v14463fb;
  wire v14463fc;
  wire v14463fd;
  wire v14463fe;
  wire v14463ff;
  wire v1446400;
  wire v1446401;
  wire v1446402;
  wire v1446403;
  wire v1446404;
  wire v1446405;
  wire v1446406;
  wire v1446407;
  wire v1446408;
  wire v1446409;
  wire v144640a;
  wire v144640b;
  wire v144640c;
  wire v144640d;
  wire v144640e;
  wire v144640f;
  wire v1446410;
  wire v1446411;
  wire v1446412;
  wire v1446413;
  wire v1446414;
  wire v1446415;
  wire v1446416;
  wire v1446417;
  wire v1446418;
  wire v1446419;
  wire v144641a;
  wire v144641b;
  wire v144641c;
  wire v144641d;
  wire v144641e;
  wire v144641f;
  wire v1446420;
  wire v1446421;
  wire v1446422;
  wire v1446423;
  wire v1446424;
  wire v1446425;
  wire v1446426;
  wire v1446427;
  wire v1446428;
  wire v1446429;
  wire v144642a;
  wire v144642b;
  wire v144642c;
  wire v144642d;
  wire v144642e;
  wire v144642f;
  wire v1446430;
  wire v1446431;
  wire v1446432;
  wire v1446433;
  wire v1446434;
  wire v1446435;
  wire v1446436;
  wire v1446437;
  wire v1446438;
  wire v1446439;
  wire v144643a;
  wire v144643b;
  wire v144643c;
  wire v144643d;
  wire v144643e;
  wire v144643f;
  wire v1446440;
  wire v1446441;
  wire v1446442;
  wire v1446443;
  wire v1446444;
  wire v1446445;
  wire v1446446;
  wire v1446447;
  wire v1446448;
  wire v1446449;
  wire v144644a;
  wire v144644b;
  wire v144644c;
  wire v144644d;
  wire v144644e;
  wire v144644f;
  wire v1446450;
  wire v1446455;
  wire v1446456;
  wire v1446457;
  wire v1446459;
  wire v144645a;
  wire v144645b;
  wire v144645d;
  wire v144645e;
  wire v144645f;
  wire v1446460;
  wire v1446461;
  wire v1446462;
  wire v1446463;
  wire v1446464;
  wire v1446465;
  wire v1446466;
  wire v1446467;
  wire v845584;
  wire v1446468;
  wire v144646d;
  wire v144646e;
  wire v144646f;
  wire v1446471;
  wire v1446472;
  wire v1446473;
  wire v1446475;
  wire v1446476;
  wire v1446477;
  wire v1446478;
  wire v1446479;
  wire v144647a;
  wire v144647b;
  wire v144647c;
  wire v144647d;
  wire v144647e;
  wire v144647f;
  wire v1446480;
  wire v1446481;
  wire v1446482;
  wire v1446483;
  wire v1446484;
  wire v1446485;
  wire v144648a;
  wire v144648b;
  wire v144648c;
  wire v144648d;
  wire v1446493;
  wire v1446494;
  wire v144649a;
  wire v144649b;
  wire v144649c;
  wire v144649d;
  wire v144649e;
  wire v144649f;
  wire v14464a0;
  wire v14464a1;
  wire v14464a2;
  wire v14464a3;
  wire v14464a4;
  wire v14464a5;
  wire v14464a6;
  wire v14464a7;
  wire v14464a8;
  wire v1446555;
  wire v1446556;
  wire v1446558;
  wire v1446559;
  wire v144655a;
  wire v144655b;
  wire v144655c;
  wire v144655d;
  wire v144655e;
  wire v144655f;
  wire v1446560;
  wire v1446561;
  wire v1446562;
  wire v1446563;
  wire v1446564;
  wire v14465a9;
  wire v14465aa;
  wire v14465ab;
  wire v14465ac;
  wire v14465ad;
  wire v14465ae;
  wire v14465af;
  wire v14465b0;
  wire v14465b1;
  wire v14465b2;
  wire v14465b3;
  wire v14465b4;
  wire v14465b5;
  wire v14465b6;
  wire v14465b7;
  wire v14465b8;
  wire v14465b9;
  wire v14465ba;
  wire v14465bb;
  wire v14465bc;
  wire v14465bd;
  wire v14465be;
  wire v14465bf;
  wire v14465c0;
  wire v14465c1;
  wire v14465c2;
  wire v14465c3;
  wire v14465c4;
  wire v14465c5;
  wire v14465c6;
  wire v14465c7;
  wire v14465c8;
  wire v14465c9;
  wire v14465ca;
  wire v14465cb;
  wire v14465cc;
  wire v14465cd;
  wire v14465ce;
  wire v14465cf;
  wire v14465d0;
  wire v14465d1;
  wire v14465d2;
  wire v14465d3;
  wire v14465d4;
  wire v14465d5;
  wire v14465d6;
  wire v14465d7;
  wire v14465d8;
  wire v14465d9;
  wire v14465da;
  wire v14465db;
  wire v14465dc;
  wire v14465dd;
  wire v14465de;
  wire v14465df;
  wire v14465e0;
  wire v14465e1;
  wire v14465e2;
  wire v14465e3;
  wire v14465e4;
  wire v14465e5;
  wire v14465e6;
  wire v14465e7;
  wire v14465e8;
  wire v14465e9;
  wire v14465ea;
  wire v14465eb;
  wire v14465ec;
  wire v14465ed;
  wire v14465ee;
  wire v14465ef;
  wire v14465f0;
  wire v14465f1;
  wire v14465f2;
  wire v14465f3;
  wire v14465f4;
  wire v14465f5;
  wire v14465f6;
  wire v14465f7;
  wire v14465f8;
  wire v14465f9;
  wire v14465fa;
  wire v1446600;
  wire v1446601;
  wire v1446602;
  wire v1446603;
  wire v1446604;
  wire v1446605;
  wire v1446606;
  wire v1446607;
  wire v1446608;
  wire v1446609;
  wire v144660a;
  wire v144660b;
  wire v144660c;
  wire v144660d;
  wire v144660e;
  wire v144660f;
  wire v1446610;
  wire v1446611;
  wire v1446612;
  wire v1446613;
  wire v1446614;
  wire v1446615;
  wire v1446616;
  wire v1446617;
  wire v1446618;
  wire v1446619;
  wire v144661a;
  wire v144661b;
  wire v144661c;
  wire v144661d;
  wire v144661e;
  wire v144661f;
  wire v1446620;
  wire v1446621;
  wire v1446622;
  wire v1446623;
  wire v1446624;
  wire v1446625;
  wire v1446626;
  wire v1446627;
  wire v1446628;
  wire v1446629;
  wire v144662a;
  wire v144662b;
  wire v144662c;
  wire v144662d;
  wire v144662e;
  wire v144662f;
  wire v1446630;
  wire v1446631;
  wire v1446632;
  wire v1446633;
  wire v1446634;
  wire v1446635;
  wire v1446636;
  wire v1446637;
  wire v1446638;
  wire v1446639;
  wire v144663a;
  wire v144663b;
  wire v144663c;
  wire v144663d;
  wire v144663e;
  wire v144663f;
  wire v1446640;
  wire v1446641;
  wire v1446642;
  wire v1446643;
  wire v1446644;
  wire v1446645;
  wire v1446646;
  wire v1446647;
  wire v1446648;
  wire v1446649;
  wire v144664a;
  wire v144664b;
  wire v144664c;
  wire v144664d;
  wire v1446651;
  wire v1446652;
  wire v1446653;
  wire v1446654;
  wire v1446655;
  wire v1446656;
  wire v1446657;
  wire v1446658;
  wire v1446659;
  wire v144665a;
  wire v144665b;
  wire v144665f;
  wire v1446660;
  wire v1446661;
  wire v1446662;
  wire v1446663;
  wire v1446664;
  wire v1446665;
  wire v1446666;
  wire v1446667;
  wire v1446668;
  wire v1446669;
  wire v144666a;
  wire v144666f;
  wire v1446670;
  wire v1446671;
  wire v1446672;
  wire v1446673;
  wire v1446674;
  wire v1446675;
  wire v1446676;
  wire v1446677;
  wire v1446678;
  wire v144667d;
  wire v144667e;
  wire v144667f;
  wire v1446680;
  wire v1446681;
  wire v1446682;
  wire v1446683;
  wire v1446684;
  wire v1446685;
  wire v1446686;
  wire v1446687;
  wire v1446688;
  wire v1446689;
  wire v144668a;
  wire v144668b;
  wire v144668c;
  wire v144668d;
  wire v144668e;
  wire v1446693;
  wire v1446694;
  wire v1446695;
  wire v1446696;
  wire v1446697;
  wire v1446698;
  wire v1446699;
  wire v144669a;
  wire v144669b;
  wire v144669c;
  wire v14466a1;
  wire v14466a2;
  wire v14466a3;
  wire v14466a4;
  wire v14466a5;
  wire v14466a6;
  wire v14466a7;
  wire v14466a8;
  wire v14466a9;
  wire v14466aa;
  wire v14466ab;
  wire v14466ac;
  wire v14466ad;
  wire v14466ae;
  wire v14466af;
  wire v14466b0;
  wire v14466b1;
  wire v14466b6;
  wire v14466b7;
  wire v14466b8;
  wire v14466b9;
  wire v14466ba;
  wire v14466bb;
  wire v14466bc;
  wire v14466bd;
  wire v14466be;
  wire v14466bf;
  wire v14466c4;
  wire v14466c5;
  wire v14466c6;
  wire v14466c7;
  wire v14466c8;
  wire v14466c9;
  wire v14466ca;
  wire v14466cb;
  wire v14466cc;
  wire v14466cd;
  wire v14466ce;
  wire v14466cf;
  wire v14466d0;
  wire v14466d1;
  wire v14466d2;
  wire v14466d3;
  wire v14466d4;
  wire v14466d5;
  wire v14466d6;
  wire v14466d7;
  wire v14466d8;
  wire v14466d9;
  wire v14466da;
  wire v14466db;
  wire v14466dc;
  wire v14466dd;
  wire v14466de;
  wire v14466df;
  wire v14466e0;
  wire v14466e1;
  wire v14466e2;
  wire v14466e3;
  wire v14466e4;
  wire v14466e5;
  wire v14466e6;
  wire v14466e7;
  wire v14466e8;
  wire v14466e9;
  wire v14466ea;
  wire v14466eb;
  wire v14466ec;
  wire v14466ed;
  wire v14466ee;
  wire v14466ef;
  wire v14466f0;
  wire v14466f1;
  wire v14466f2;
  wire v14466f3;
  wire v14466f4;
  wire v14466f5;
  wire v14466f6;
  wire v14466f7;
  wire v14466f8;
  wire v14466f9;
  wire v14466fd;
  wire v14466fe;
  wire v14466ff;
  wire v1446700;
  wire v1446701;
  wire v1446702;
  wire v1446703;
  wire v1446704;
  wire v1446705;
  wire v1446706;
  wire v1446707;
  wire v144670b;
  wire v144670c;
  wire v144670d;
  wire v144670e;
  wire v144670f;
  wire v1446710;
  wire v1446711;
  wire v1446712;
  wire v1446713;
  wire v1446714;
  wire v1446715;
  wire v1446716;
  wire v1446717;
  wire v1446718;
  wire v1446719;
  wire v144671a;
  wire v144671b;
  wire v144671c;
  wire v144671d;
  wire v144671e;
  wire v144671f;
  wire v1446720;
  wire v1446721;
  wire v1446722;
  wire v1446723;
  wire v1446724;
  wire v1446725;
  wire v1446726;
  wire v1446727;
  wire v1446728;
  wire v1446729;
  wire v144672a;
  wire v144672b;
  wire v144672c;
  wire v144672d;
  wire v144672e;
  wire v144672f;
  wire v1446730;
  wire v1446731;
  wire v1446732;
  wire v1446733;
  wire v1446734;
  wire v1446735;
  wire v1446736;
  wire v1446737;
  wire v1446738;
  wire v1446739;
  wire v144673a;
  wire v144673b;
  wire v144673c;
  wire v144673d;
  wire v144673e;
  wire v144673f;
  wire v1446740;
  wire v1446741;
  wire v1446742;
  wire v1446743;
  wire v1446744;
  wire v1446745;
  wire v1446746;
  wire v1446747;
  wire v1446748;
  wire v1446749;
  wire v144674a;
  wire v144674b;
  wire v144674c;
  wire v144674d;
  wire v144674e;
  wire v1445f52;
  wire v1445f53;
  wire v1445f54;
  wire v1445f55;
  wire v1445f56;
  wire v1445f57;
  wire v1445f58;
  wire v1445f59;
  wire v1445f5a;
  wire v1445f5b;
  wire v1445f5c;
  wire v1445f5d;
  wire v1445f5e;
  wire v1445f5f;
  wire v1445f60;
  wire v1445f61;
  wire v1445f62;
  wire v1445f63;
  wire v1445f64;
  wire v1445f65;
  wire v1445f66;
  wire v1445f67;
  wire v1445f68;
  wire v1445f69;
  wire v1445f6a;
  wire v1445f6b;
  wire v1445f6c;
  wire v1445f6d;
  wire v1445f6e;
  wire v1445f6f;
  wire v1445f70;
  wire v1445f71;
  wire v1445f72;
  wire v1445f73;
  wire v1445f74;
  wire v1445f75;
  wire v1445f76;
  wire v1445f77;
  wire v1445f78;
  wire v1445f79;
  wire v1445f7a;
  wire v1445f7b;
  wire v1445f7c;
  wire v1445f7d;
  wire v1445f7e;
  wire v1445f7f;
  wire v1445f80;
  wire v1445f81;
  wire v1445f82;
  wire v1445f83;
  wire v1445f84;
  wire v1445f85;
  wire v1445f86;
  wire v1445f87;
  wire v1445f88;
  wire v1445f89;
  wire v1445f8a;
  wire v1445f8b;
  wire v1445f8c;
  wire v1445f8d;
  wire v1445f8e;
  wire v1445f8f;
  wire v1445f90;
  wire v1445f91;
  wire v1445f92;
  wire v1445f93;
  wire v1445f94;
  wire v1445f95;
  wire v1445f96;
  wire v1445f97;
  wire v1445f98;
  wire v1445f99;
  wire v1445f9a;
  wire v1445f9b;
  wire v1445f9c;
  wire v1445f9d;
  wire v1445f9e;
  wire v1445f9f;
  wire v1445fa0;
  wire v1445fa1;
  wire v1445fa2;
  wire v1445fa3;
  wire v1445fa4;
  wire v1445fa5;
  wire v1445fa6;
  wire v1445fa7;
  wire v1445fa8;
  wire v1445fa9;
  wire v1445faa;
  wire v1445fab;
  wire v1445fac;
  wire v1445fad;
  wire v1445fae;
  wire v1445faf;
  wire v1445fb0;
  wire v1445fb1;
  wire v1445fb2;
  wire v1445fb3;
  wire v1445fb4;
  wire v1445fb5;
  wire v1445fb6;
  wire v1445fb7;
  wire v1445fb8;
  wire v1445fb9;
  wire v1445fba;
  wire v1445fbb;
  wire v1445fbc;
  wire v1445fbd;
  wire v1445fbe;
  wire v1445fbf;
  wire v1445fc0;
  wire v1445fc1;
  wire v1445fc2;
  wire v1445fc3;
  wire v1445fc4;
  wire v1445fc5;
  wire v1445fc6;
  wire v1445fc7;
  wire v1445fc8;
  wire v1445fc9;
  wire v1445fca;
  wire v1445fcb;
  wire v1445fcc;
  wire v1445fcd;
  wire v1445fce;
  wire v1445fcf;
  wire v1445fd0;
  wire v1445fd1;
  wire v1445fd2;
  wire v1445fd3;
  wire v1445fd4;
  wire v1445fd5;
  wire v1445fd6;
  wire v1445fd7;
  wire v1445fd8;
  wire v1445fd9;
  wire v1445fda;
  wire v1445fdb;
  wire v1445fdc;
  wire v1445fdd;
  wire v1445fde;
  wire v1445fdf;
  wire v1445fe0;
  wire v1445fe1;
  wire v1445fe2;
  wire v1445fe3;
  wire v1445fe4;
  wire v1445fe5;
  wire v1445fe6;
  wire v1445fe7;
  wire v1445fe8;
  wire v1445fe9;
  wire v1445fea;
  wire v1445feb;
  wire v1445fec;
  wire v1445fed;
  wire v1445fee;
  wire v1445fef;
  wire v1445ff0;
  wire v1445ff1;
  wire v1445ff2;
  wire v1445ff3;
  wire v1445ff4;
  wire v1445ff5;
  wire v1445ff6;
  wire v1445ff7;
  wire v1445ff8;
  wire v1445ff9;
  wire v1445ffa;
  wire v1445ffb;
  wire v1445ffc;
  wire v1445ffd;
  wire v1445ffe;
  wire v1445fff;
  wire v1446000;
  wire v1446001;
  wire v1446002;
  wire v1446003;
  wire v1446004;
  wire v1446005;
  wire v1446006;
  wire v1446007;
  wire v1446008;
  wire v1446009;
  wire v144600a;
  wire v144600b;
  wire v144600c;
  wire v144600d;
  wire v144600e;
  wire v144600f;
  wire v1446010;
  wire v1446011;
  wire v1446012;
  wire v1446013;
  wire v1446014;
  wire v1446015;
  wire v1446016;
  wire v1446017;
  wire v1446018;
  wire v1446019;
  wire v144601a;
  wire v144601b;
  wire v144601c;
  wire v144602b;
  wire v144602c;
  wire v1446038;
  wire v1446039;
  wire v144603a;
  wire v144603b;
  wire v144603c;
  wire v144603d;
  wire v144603e;
  wire v144603f;
  wire v1446040;
  wire v1446041;
  wire v1446042;
  wire v1446043;
  wire v1446044;
  wire v1446045;
  wire v1446046;
  wire v1446047;
  wire v1446048;
  wire v1446049;
  wire v144604a;
  wire v144604b;
  wire v144604c;
  wire v144604d;
  wire v144604e;
  wire v144604f;
  wire v1446050;
  wire v1446051;
  wire v1446052;
  wire v1446053;
  wire v1446054;
  wire v1446055;
  wire v1446056;
  wire v1446057;
  wire v1446058;
  wire v1446059;
  wire v144605a;
  wire v144605b;
  wire v144605c;
  wire v144605d;
  wire v144605e;
  wire v144605f;
  wire v1446060;
  wire v1446061;
  wire v1446062;
  wire v1446063;
  wire v1446064;
  wire v1446065;
  wire v1446066;
  wire v1446067;
  wire v1446068;
  wire v1446069;
  wire v144606a;
  wire v144606b;
  wire v144606c;
  wire v144606d;
  wire v144606e;
  wire v144606f;
  wire v1446070;
  wire v1446071;
  wire v1446072;
  wire v1446073;
  wire v1446074;
  wire v1446075;
  wire v1446076;
  wire v1446077;
  wire v1446078;
  wire v1446079;
  wire v144607a;
  wire v144607b;
  wire v144607c;
  wire v144607d;
  wire v144607e;
  wire v144607f;
  wire v1446080;
  wire v1446081;
  wire v1446082;
  wire v1446083;
  wire v1446084;
  wire v1446085;
  wire v1446086;
  wire v1446087;
  wire v1446088;
  wire v1446089;
  wire v144608a;
  wire v144608b;
  wire v144608c;
  wire v144608d;
  wire v144608e;
  wire v144608f;
  wire v1446090;
  wire v1446091;
  wire v1446092;
  wire v1446093;
  wire v1446094;
  wire v1446095;
  wire v1446096;
  wire v1446097;
  wire v1446098;
  wire v1446099;
  wire v144609a;
  wire v144609b;
  wire v144609c;
  wire v144609d;
  wire v144609e;
  wire v144609f;
  wire v14460a0;
  wire v14460a1;
  wire v14460a2;
  wire v14460a3;
  wire v14460a4;
  wire v14460a5;
  wire v14460a6;
  wire v14460a7;
  wire v14460a8;
  wire v14460a9;
  wire v14460aa;
  wire v14460ab;
  wire v14460ac;
  wire v14460ad;
  wire v14460ae;
  wire v14460af;
  wire v14460b0;
  wire v14460b1;
  wire v14460b2;
  wire v14460b3;
  wire v14460b4;
  wire v14460b5;
  wire v14460b6;
  wire v14460b7;
  wire v14460b8;
  wire v14460b9;
  wire v14460ba;
  wire v14460bb;
  wire v14460bc;
  wire v14460bd;
  wire v14460be;
  wire v14460bf;
  wire v14460c0;
  wire v14460c1;
  wire v14460c2;
  wire v14460c3;
  wire v14460c4;
  wire v14460c5;
  wire v14460c6;
  wire v14460c7;
  wire v14460c8;
  wire v14460c9;
  wire v14460ca;
  wire v14460cb;
  wire v14460cc;
  wire v14460cd;
  wire v14460ce;
  wire v14460cf;
  wire v14460d0;
  wire v14460d1;
  wire v14460d2;
  wire v14460d3;
  wire v14460d4;
  wire v14460d5;
  wire v14460d6;
  wire v14460d7;
  wire v14460d8;
  wire v14460d9;
  wire v14460da;
  wire v14460db;
  wire v14460dc;
  wire v14460dd;
  wire v14460de;
  wire v14460df;
  wire v14460e0;
  wire v14460e1;
  wire v14460e2;
  wire v14460e3;
  wire v14460e4;
  wire v14460e5;
  wire v14460e6;
  wire v14460e7;
  wire v14460e8;
  wire v14460e9;
  wire v14460ea;
  wire v14460eb;
  wire v14460ec;
  wire v14460ed;
  wire v14460ee;
  wire v14460ef;
  wire v14460f0;
  wire v14460f1;
  wire v14460f2;
  wire v14460f3;
  wire v14460f4;
  wire v14460f5;
  wire v14460f6;
  wire v14460f7;
  wire v14460f8;
  wire v14460f9;
  wire v14460fa;
  wire v14460fb;
  wire v14460fc;
  wire v14460fd;
  wire v14460fe;
  wire v14460ff;
  wire v1446100;
  wire v1446101;
  wire v1446102;
  wire v1446103;
  wire v1446104;
  wire v1446105;
  wire v1446106;
  wire v1446107;
  wire v1446108;
  wire v1446109;
  wire v144610a;
  wire v144610b;
  wire v144610c;
  wire v144610d;
  wire v144610e;
  wire v144610f;
  wire v1446110;
  wire v1446111;
  wire v1446112;
  wire v1446113;
  wire v1446114;
  wire v1446115;
  wire v1446116;
  wire v1446117;
  wire v1446118;
  wire v1446119;
  wire v144611a;
  wire v144611b;
  wire v144611c;
  wire v144611d;
  wire v144611e;
  wire v144611f;
  wire v1446120;
  wire v1446121;
  wire v1446122;
  wire v1446123;
  wire v1446124;
  wire v1446125;
  wire v1446126;
  wire v1446127;
  wire v1446128;
  wire v1446129;
  wire v144612a;
  wire v144612b;
  wire v144612c;
  wire v144612d;
  wire v144612e;
  wire v144612f;
  wire v1446130;
  wire v1446131;
  wire v1446132;
  wire v1446133;
  wire v1446134;
  wire v1446135;
  wire v1446136;
  wire v1446137;
  wire v1446138;
  wire v1446139;
  wire v144613a;
  wire v144613b;
  wire v144613c;
  wire v144613d;
  wire v144613e;
  wire v144613f;
  wire v1446140;
  wire v1446141;
  wire v1446142;
  wire v1446143;
  wire v1446144;
  wire v1446145;
  wire v1446146;
  wire v1446147;
  wire v1446148;
  wire v1446149;
  wire v144614a;
  wire v144614b;
  wire v144614c;
  wire v144614d;
  wire v144614e;
  wire v144614f;
  wire v1446150;
  wire v1446151;
  wire v1446152;
  wire v1446153;
  wire v1446154;
  wire v1446155;
  wire v1446156;
  wire v1446157;
  wire v1446158;
  wire v1446159;
  wire v144615a;
  wire v144615b;
  wire v144615c;
  wire v144615d;
  wire v144615e;
  wire v144615f;
  wire v1446160;
  wire v1446161;
  wire v1446162;
  wire v1446163;
  wire v1446164;
  wire v1446165;
  wire v1446166;
  wire v1446167;
  wire v1446168;
  wire v1446169;
  wire v144616a;
  wire v144616b;
  wire v144616c;
  wire v144616d;
  wire v144616e;
  wire v144616f;
  wire v1446170;
  wire v1446171;
  wire v1446172;
  wire v1446173;
  wire v1446174;
  wire v1446175;
  wire v1446176;
  wire v1446177;
  wire v1446178;
  wire v1446179;
  wire v144617a;
  wire v144617b;
  wire v144617c;
  wire v144617d;
  wire v144617e;
  wire v144617f;
  wire v1446180;
  wire v1446181;
  wire v1446182;
  wire v1446183;
  wire v1446184;
  wire v1446185;
  wire v1446186;
  wire v1446187;
  wire v1446188;
  wire v1446189;
  wire v144618a;
  wire v144618b;
  wire v144618c;
  wire v144618d;
  wire v144618e;
  wire v144618f;
  wire v1446190;
  wire v1446191;
  wire v1446192;
  wire v1446193;
  wire v1446194;
  wire v1446195;
  wire v1446196;
  wire v1446197;
  wire v1446198;
  wire v1446199;
  wire v144619a;
  wire v144619b;
  wire v144619c;
  wire v144619d;
  wire v144619e;
  wire v14461b0;
  wire v14461b1;
  wire v14461b2;
  wire v14461b3;
  wire v14461b8;
  wire v14461b9;
  wire v14461ba;
  wire v14461bb;
  wire v14461bc;
  wire v14461bd;
  wire v14461be;
  wire v14461bf;
  wire v14461c0;
  wire v14461c1;
  wire v14461c2;
  wire v14461c3;
  wire v14461c4;
  wire v14461c5;
  wire v14461c6;
  wire v14461cc;
  wire v14461cd;
  wire v14461ce;
  wire v14461cf;
  wire v14461d4;
  wire v14461d5;
  wire v14461d6;
  wire v14461d7;
  wire v14461d8;
  wire v14461d9;
  wire v14461da;
  wire v14461db;
  wire v14461dc;
  wire v14461dd;
  wire v14461de;
  wire v14461df;
  wire v14461e0;
  wire v14461e1;
  wire v14461e2;
  wire v14461e3;
  wire v14461e4;
  wire v14461e5;
  wire v14461e6;
  wire v14461e7;
  wire v14461e8;
  wire v14461e9;
  wire v14461ea;
  wire v14461eb;
  wire v14461ec;
  wire v14461ed;
  wire v14461ee;
  wire v14461ef;
  wire v14461f0;
  wire v14461f1;
  wire v14461f2;
  wire v14461f3;
  wire v14461f4;
  wire v14461f5;
  wire v14461fa;
  wire v14461fb;
  wire v14461fc;
  wire v14461fd;
  wire v14461fe;
  wire v14461ff;
  wire v1446200;
  wire v1446201;
  wire v1446202;
  wire v1446203;
  wire v1446208;
  wire v1446209;
  wire v144620a;
  wire v144620b;
  wire v144620c;
  wire v144620d;
  wire v144620e;
  wire v144620f;
  wire v1446210;
  wire v1446211;
  wire v1446212;
  wire v1446213;
  wire v1446214;
  wire v1446215;
  wire v1446216;
  wire v1446217;
  wire v1446218;
  wire v1446219;
  wire v144621a;
  wire v144621b;
  wire v144621c;
  wire v144621d;
  wire v1446221;
  wire v1446222;
  wire v1446223;
  wire v1446224;
  wire v1446228;
  wire v1446229;
  wire v144622a;
  wire v144622b;
  wire v144622c;
  wire v144622d;
  wire v144622e;
  wire v1446232;
  wire v1446233;
  wire v1446234;
  wire v1446235;
  wire v1446236;
  wire v1446237;
  wire v1446238;
  wire v1446239;
  wire v144623a;
  wire v144623b;
  wire v144623c;
  wire v144623d;
  wire v144623e;
  wire v144623f;
  wire v1446243;
  wire v1446244;
  wire v1446245;
  wire v1446246;
  wire v144624a;
  wire v144624b;
  wire v144624c;
  wire v144624d;
  wire v144624e;
  wire v144624f;
  wire v1446250;
  wire v1446254;
  wire v1446255;
  wire v1446256;
  wire v1446257;
  wire v1446258;
  wire v1446259;
  wire v144625a;
  wire v144625b;
  wire v144625c;
  wire v144625d;
  wire v144625e;
  wire v144625f;
  wire v1446260;
  wire v1446261;
  wire v1446262;
  wire v1446263;
  wire v1446264;
  wire v1446265;
  wire v1446266;
  wire v1446267;
  wire v1446268;
  wire v1446269;
  wire v144626a;
  wire v144626b;
  wire v144626c;
  wire v144626d;
  wire v144626e;
  wire v144626f;
  wire v1446270;
  wire v1446271;
  wire v1446272;
  wire v1446273;
  wire v1446274;
  wire v1446275;
  wire v1446276;
  wire v1446277;
  wire v1446278;
  wire v1446279;
  wire v144627a;
  wire v144627b;
  wire v144627c;
  wire v144627d;
  wire v144627e;
  wire v144627f;
  wire v1446280;
  wire v1446281;
  wire v1446282;
  wire v1446283;
  wire v1446284;
  wire v1446285;
  wire v1446286;
  wire v1446287;
  wire v1446288;
  wire v1446289;
  wire v144628a;
  wire v144628b;
  wire v144628c;
  wire v144628d;
  wire v144628e;
  wire v144628f;
  wire v1446290;
  wire v1446291;
  wire v1446292;
  wire v1446293;
  wire v1446294;
  wire v1446298;
  wire v1446299;
  wire v144629a;
  wire v144629b;
  wire v144629f;
  wire v14462a0;
  wire v14462a1;
  wire v14462a2;
  wire v14462a3;
  wire v14462a4;
  wire v14462a5;
  wire v14462e6;
  wire v14462e7;
  wire v14462e8;
  wire v14462e9;
  wire v14462ea;
  wire v14462eb;
  wire v14462ec;
  wire v14462ed;
  wire v14462ee;
  wire v14462ef;
  wire v14462f0;
  wire v14462f1;
  wire v14462f2;
  wire v14462f3;
  wire v14462f4;
  wire v14462f5;
  wire v14462f6;
  wire v14462f7;
  wire v14462f8;
  wire v14462f9;
  wire v14462fa;
  wire v14462fe;
  wire v14462ff;
  wire v1446300;
  wire v1446301;
  wire v1446302;
  wire v1446303;
  wire v1446304;
  wire v1446308;
  wire v1446309;
  wire v144630a;
  wire v144630b;
  wire v144630c;
  wire v1446310;
  wire v1446311;
  wire v1446312;
  wire v1446313;
  wire v1446314;
  wire v1446315;
  wire v1446316;
  wire v144631a;
  wire v144631b;
  wire v144631c;
  wire v144631d;
  wire v144631e;
  wire v144631f;
  wire v1446320;
  wire v1446321;
  wire v1446322;
  wire v1446323;
  wire v1446324;
  wire v1446325;
  wire v1446326;
  wire v1446327;
  wire v1446328;
  wire v1446329;
  wire v144632a;
  wire v144632b;
  wire v144632c;
  wire v144632d;
  wire v144632e;
  wire v144632f;
  wire v1446330;
  wire v1446331;
  wire v1446332;
  wire v1446333;
  wire v1446334;
  wire v1446335;
  wire v1446336;
  wire v1446337;
  wire v1446338;
  wire v1446339;
  wire v144633a;
  wire v144633b;
  wire v144633c;
  wire v144633d;
  wire v144633e;
  wire v144633f;
  wire v1446340;
  wire v1446341;
  wire v1446342;
  wire v1446343;
  wire v1446344;
  wire v1446345;
  wire v1446346;
  wire v1446347;
  wire v1446348;
  wire v1446349;
  wire v144634a;
  wire v144634b;
  wire v144634c;
  wire v144634d;
  wire v144634e;
  wire v144634f;
  wire v1445b55;
  wire v1445b56;
  wire v1445b57;
  wire v1445b58;
  wire v1445b5c;
  wire v1445b5d;
  wire v1445b5e;
  wire v1445b5f;
  wire v1445b60;
  wire v1445b64;
  wire v1445b65;
  wire v1445b66;
  wire v1445b67;
  wire v1445b68;
  wire v1445b69;
  wire v1445b6a;
  wire v1445b6b;
  wire v1445b6c;
  wire v1445b6d;
  wire v1445b6e;
  wire v1445b6f;
  wire v1445b70;
  wire v1445b71;
  wire v1445b72;
  wire v1445b73;
  wire v1445b74;
  wire v1445b75;
  wire v1445b76;
  wire v1445b77;
  wire v1445b78;
  wire v1445b79;
  wire v1445b7a;
  wire v1445b7b;
  wire v1445b7c;
  wire v1445b7d;
  wire v1445b7e;
  wire v1445b7f;
  wire v1445b80;
  wire v1445b81;
  wire v1445b82;
  wire v1445b83;
  wire v1445b84;
  wire v1445b85;
  wire v1445b86;
  wire v1445b87;
  wire v1445b88;
  wire v1445b89;
  wire v1445b8a;
  wire v1445b8b;
  wire v1445b8c;
  wire v1445b8d;
  wire v1445b8e;
  wire v1445b8f;
  wire v1445b90;
  wire v1445b91;
  wire v1445b92;
  wire v1445b93;
  wire v1445b94;
  wire v1445b95;
  wire v1445b9b;
  wire v1445b9c;
  wire v1445b9d;
  wire v1445b9e;
  wire v1445ba3;
  wire v1445ba4;
  wire v1445ba5;
  wire v1445ba6;
  wire v1445ba7;
  wire v1445ba8;
  wire v1445ba9;
  wire v1445baa;
  wire v1445bab;
  wire v1445bac;
  wire v1445bad;
  wire v1445bae;
  wire v1445baf;
  wire v1445bb0;
  wire v1445bb1;
  wire v1445bb2;
  wire v1445bb3;
  wire v1445bb4;
  wire v1445bb5;
  wire v1445bb6;
  wire v1445bb7;
  wire v1445bb8;
  wire v1445bb9;
  wire v1445bba;
  wire v1445bbb;
  wire v1445bbc;
  wire v1445bbd;
  wire v1445bc2;
  wire v1445bc3;
  wire v1445bc4;
  wire v1445bc5;
  wire v1445bc6;
  wire v1445bc7;
  wire v1445bc8;
  wire v1445bc9;
  wire v1445bca;
  wire v1445bcb;
  wire v1445bcc;
  wire v1445bd1;
  wire v1445bd2;
  wire v1445bd3;
  wire v1445bd4;
  wire v1445bd5;
  wire v1445bd6;
  wire v1445bd7;
  wire v1445bd8;
  wire v1445bd9;
  wire v1445bda;
  wire v1445bdb;
  wire v1445bdc;
  wire v1445bdd;
  wire v1445bde;
  wire v1445bdf;
  wire v1445be0;
  wire v1445be1;
  wire v1445be2;
  wire v1445be3;
  wire v1445be4;
  wire v1445be5;
  wire v1445be6;
  wire v1445be7;
  wire v1445be8;
  wire v1445be9;
  wire v1445bea;
  wire v1445beb;
  wire v1445bec;
  wire v1445bed;
  wire v1445bee;
  wire v1445bef;
  wire v1445bf0;
  wire v1445bf1;
  wire v1445bf2;
  wire v1445bf3;
  wire v1445bf7;
  wire v1445bf8;
  wire v1445bf9;
  wire v1445bfa;
  wire v1445bfe;
  wire v1445d7f;
  wire v1445d80;
  wire v1445d81;
  wire v1445d82;
  wire v1445d83;
  wire v1445d84;
  wire v1445d85;
  wire v1445d86;
  wire v1445d87;
  wire v1445d88;
  wire v1445d89;
  wire v1445d8a;
  wire v1445d8b;
  wire v1445d8c;
  wire v1445d8d;
  wire v1445d8e;
  wire v1445d8f;
  wire v1445d90;
  wire v1445d91;
  wire v1445d92;
  wire v1445d93;
  wire v1445d94;
  wire v1445d95;
  wire v1445d96;
  wire v1445d97;
  wire v1445d98;
  wire v1445d99;
  wire v1445d9a;
  wire v1445d9b;
  wire v1445d9c;
  wire v1445d9d;
  wire v1445d9e;
  wire v1445d9f;
  wire v1445da0;
  wire v1445da1;
  wire v1445da2;
  wire v1445da3;
  wire v1445da4;
  wire v1445da5;
  wire v1445da6;
  wire v1445da7;
  wire v1445da8;
  wire v1445da9;
  wire v1445db2;
  wire v1445db3;
  wire v1445db4;
  wire v1445db5;
  wire v1445db6;
  wire v1445db7;
  wire v1445db8;
  wire v1445db9;
  wire v1445dba;
  wire v1445dbb;
  wire v1445dc1;
  wire v1445dc2;
  wire v1445dc3;
  wire v1445dc4;
  wire v1445dc5;
  wire v1445dc6;
  wire v1445dc7;
  wire v1445dc8;
  wire v1445dc9;
  wire v1445dca;
  wire v1445dcb;
  wire v1445dcc;
  wire v1445dcd;
  wire v1445dce;
  wire v1445dcf;
  wire v1445dd0;
  wire v1445dd1;
  wire v1445dd2;
  wire v1445dd3;
  wire v1445dd7;
  wire v1445dd8;
  wire v1445dd9;
  wire v1445dda;
  wire v1445ddb;
  wire v1445ddc;
  wire v1445ddd;
  wire v1445dde;
  wire v1445ddf;
  wire v1445de0;
  wire v1445de1;
  wire v1445de5;
  wire v1445de6;
  wire v1445de7;
  wire v1445de8;
  wire v1445de9;
  wire v1445dea;
  wire v1445deb;
  wire v1445dec;
  wire v1445ded;
  wire v1445dee;
  wire v1445def;
  wire v1445df0;
  wire v1445df1;
  wire v1445df2;
  wire v1445df3;
  wire v1445df4;
  wire v1445df5;
  wire v1445df6;
  wire v1445df7;
  wire v1445df8;
  wire v1445df9;
  wire v1445dfa;
  wire v1445dfb;
  wire v1445dfc;
  wire v1445dfd;
  wire v1445dfe;
  wire v1445dff;
  wire v1445e00;
  wire v1445e01;
  wire v1445e02;
  wire v1445e03;
  wire v1445e04;
  wire v1445e05;
  wire v1445e06;
  wire v1445e07;
  wire v1445e08;
  wire v1445e09;
  wire v1445e0a;
  wire v1445e0b;
  wire v1445e0c;
  wire v1445e0d;
  wire v1445e0e;
  wire v1445e0f;
  wire v1445e10;
  wire v1445e11;
  wire v1445e12;
  wire v1445e13;
  wire v1445e17;
  wire v1445e18;
  wire v1445e19;
  wire v1445e1a;
  wire v1445e1b;
  wire v1445e1c;
  wire v1445e1d;
  wire v1445e1e;
  wire v1445e1f;
  wire v1445e20;
  wire v1445e21;
  wire v1445e22;
  wire v1445e23;
  wire v1445e24;
  wire v1445e25;
  wire v1445e26;
  wire v1445e27;
  wire v1445e28;
  wire v1445e29;
  wire v1445e2a;
  wire v1445e2b;
  wire v1445e2c;
  wire v1445e2d;
  wire v1445e2e;
  wire v1445e2f;
  wire v1445e30;
  wire v1445e31;
  wire v1445e32;
  wire v1445e33;
  wire v1445e34;
  wire v1445e35;
  wire v1445e36;
  wire v1445e37;
  wire v1445e38;
  wire v1445e39;
  wire v1445e3a;
  wire v1445e3b;
  wire v1445e3c;
  wire v1445e3d;
  wire v1445e3e;
  wire v1445e3f;
  wire v1445e45;
  wire v1445e46;
  wire v1445e47;
  wire v1445e48;
  wire v1445e49;
  wire v1445e4a;
  wire v1445e4b;
  wire v1445e4c;
  wire v1445e4d;
  wire v1445e4e;
  wire v1445e4f;
  wire v1445e50;
  wire v1445e51;
  wire v1445e52;
  wire v1445e53;
  wire v1445e54;
  wire v1445e55;
  wire v1445e56;
  wire v1445e57;
  wire v1445e58;
  wire v1445e59;
  wire v1445e5a;
  wire v1445e5b;
  wire v1445e5c;
  wire v1445e5d;
  wire v1445e5e;
  wire v1445e5f;
  wire v1445e60;
  wire v1445e64;
  wire v1445e65;
  wire v1445e66;
  wire v1445e67;
  wire v1445e68;
  wire v1445e69;
  wire v1445e6a;
  wire v1445e6b;
  wire v1445e6c;
  wire v1445e6d;
  wire v1445e6e;
  wire v1445e6f;
  wire v1445e70;
  wire v1445e71;
  wire v1445e72;
  wire v1445e73;
  wire v1445e74;
  wire v1445e75;
  wire v1445e76;
  wire v1445e77;
  wire v1445e78;
  wire v1445e79;
  wire v1445e7a;
  wire v1445e7b;
  wire v1445e7c;
  wire v1445e7d;
  wire v1445e7e;
  wire v1445e7f;
  wire v1445e80;
  wire v1445e81;
  wire v1445e82;
  wire v1445e83;
  wire v1445e84;
  wire v1445e85;
  wire v1445e86;
  wire v1445e87;
  wire v1445e88;
  wire v1445e89;
  wire v1445e8a;
  wire v1445e8b;
  wire v1445e8c;
  wire v1445e8d;
  wire v1445e8e;
  wire v1445e8f;
  wire v1445e90;
  wire v1445e91;
  wire v1445e92;
  wire v1445e93;
  wire v1445e94;
  wire v1445e95;
  wire v1445e96;
  wire v1445e97;
  wire v1445e98;
  wire v1445e99;
  wire v1445e9a;
  wire v1445e9b;
  wire v1445e9c;
  wire v1445e9d;
  wire v1445e9e;
  wire v1445e9f;
  wire v1445ea0;
  wire v1445ea1;
  wire v1445ea2;
  wire v1445ea3;
  wire v1445ea4;
  wire v1445ea5;
  wire v1445ea6;
  wire v1445ea7;
  wire v1445ea8;
  wire v1445ea9;
  wire v1445eaa;
  wire v1445eab;
  wire v1445eac;
  wire v1445ead;
  wire v1445eae;
  wire v1445eaf;
  wire v1445eb0;
  wire v1445eb1;
  wire v1445eb2;
  wire v1445eb3;
  wire v1445eb4;
  wire v1445eb5;
  wire v1445eb6;
  wire v1445eb7;
  wire v1445eb8;
  wire v1445eb9;
  wire v1445eba;
  wire v1445ebb;
  wire v1445ebc;
  wire v1445ebd;
  wire v1445ebe;
  wire v1445ebf;
  wire v1445ec0;
  wire v1445ec1;
  wire v1445ec2;
  wire v1445ec3;
  wire v1445ec4;
  wire v1445ec5;
  wire v1445ec6;
  wire v1445ec7;
  wire v1445ec8;
  wire v1445ec9;
  wire v1445eca;
  wire v1445ecb;
  wire v1445ecc;
  wire v1445ecd;
  wire v1445ece;
  wire v1445ecf;
  wire v1445ed0;
  wire v1445ed1;
  wire v1445ed2;
  wire v1445ed3;
  wire v1445ed4;
  wire v1445ed5;
  wire v1445ed6;
  wire v1445ed7;
  wire v1445ed8;
  wire v1445ed9;
  wire v1445eda;
  wire v1445edb;
  wire v1445edc;
  wire v1445edd;
  wire v1445ede;
  wire v1445edf;
  wire v1445ee0;
  wire v1445ee1;
  wire v1445ee2;
  wire v1445ee3;
  wire v1445ee4;
  wire v1445ee5;
  wire v1445ee6;
  wire v1445ee7;
  wire v1445ee8;
  wire v1445ee9;
  wire v1445eea;
  wire v1445eeb;
  wire v1445eec;
  wire v1445eed;
  wire v1445eee;
  wire v1445eef;
  wire v1445ef0;
  wire v1445ef1;
  wire v1445ef2;
  wire v1445ef3;
  wire v1445ef4;
  wire v1445ef5;
  wire v1445ef6;
  wire v1445ef7;
  wire v1445ef8;
  wire v1445ef9;
  wire v1445efa;
  wire v1445efb;
  wire v1445efc;
  wire v1445efd;
  wire v1445efe;
  wire v1445eff;
  wire v1445f00;
  wire v1445f01;
  wire v1445f02;
  wire v1445f03;
  wire v1445f04;
  wire v1445f05;
  wire v1445f06;
  wire v1445f07;
  wire v1445f08;
  wire v1445f09;
  wire v1445f0a;
  wire v1445f0b;
  wire v1445f0c;
  wire v1445f0d;
  wire v1445f11;
  wire v1445f12;
  wire v1445f13;
  wire v1445f14;
  wire v1445f15;
  wire v1445f16;
  wire v1445f17;
  wire v1445f18;
  wire v1445f19;
  wire v1445f1a;
  wire v1445f1b;
  wire v1445f1c;
  wire v1445f1d;
  wire v1445f1e;
  wire v1445f1f;
  wire v1445f20;
  wire v1445f21;
  wire v1445f25;
  wire v1445f26;
  wire v1445f27;
  wire v1445f28;
  wire v1445f29;
  wire v1445f34;
  wire v1445f35;
  wire v1445f36;
  wire v1445f37;
  wire v1445f38;
  wire v1445f39;
  wire v1445f3a;
  wire v1445f3f;
  wire v1445f40;
  wire v1445f41;
  wire v1445f42;
  wire v1445f47;
  wire v1445f48;
  wire v1445f49;
  wire v1445f4a;
  wire v1445f4b;
  wire v1445f4c;
  wire v1445f4d;
  wire v1445f4e;
  wire v1445f4f;
  wire v1445753;
  wire v1445754;
  wire v1445755;
  wire v1445756;
  wire v1445757;
  wire v1445758;
  wire v1445759;
  wire v144575e;
  wire v144575f;
  wire v1445760;
  wire v1445761;
  wire v1445766;
  wire v1445767;
  wire v1445768;
  wire v1445769;
  wire v144576a;
  wire v144576b;
  wire v144576c;
  wire v144576d;
  wire v144576e;
  wire v144576f;
  wire v1445770;
  wire v1445771;
  wire v1445772;
  wire v1445773;
  wire v1445774;
  wire v1445775;
  wire v1445776;
  wire v1445777;
  wire v1445778;
  wire v1445779;
  wire v144577a;
  wire v144577b;
  wire v144577c;
  wire v144577d;
  wire v144577e;
  wire v144577f;
  wire v1445780;
  wire v1445781;
  wire v1445782;
  wire v1445783;
  wire v1445784;
  wire v1445785;
  wire v1445786;
  wire v1445787;
  wire v1445788;
  wire v1445789;
  wire v144578a;
  wire v144578b;
  wire v144578c;
  wire v144578d;
  wire v144578e;
  wire v144578f;
  wire v1445790;
  wire v1445791;
  wire v1445795;
  wire v1445796;
  wire v1445797;
  wire v1445798;
  wire v1445799;
  wire v144579a;
  wire v144579b;
  wire v144579c;
  wire v144579d;
  wire v144579e;
  wire v144579f;
  wire v14457a3;
  wire v14457a4;
  wire v14457a5;
  wire v14457a6;
  wire v14457a7;
  wire v14457a8;
  wire v14457a9;
  wire v14457aa;
  wire v14457ab;
  wire v14457ac;
  wire v14457ad;
  wire v14457ae;
  wire v14457af;
  wire v14457b0;
  wire v14457b1;
  wire v14457b2;
  wire v14457b3;
  wire v14457b4;
  wire v14457b9;
  wire v14457ba;
  wire v14457bb;
  wire v14457bc;
  wire v14457bd;
  wire v14457be;
  wire v14457bf;
  wire v14457c0;
  wire v14457c1;
  wire v14457c2;
  wire v14457c3;
  wire v14457c4;
  wire v14457c5;
  wire v14457c6;
  wire v14457c7;
  wire v14457c8;
  wire v14457cd;
  wire v14457ce;
  wire v14457cf;
  wire v14457d0;
  wire v14457d1;
  wire v14457d2;
  wire v14457d3;
  wire v14457d4;
  wire v14457d5;
  wire v14457d6;
  wire v14457d7;
  wire v14457d8;
  wire v14457d9;
  wire v14457da;
  wire v14457db;
  wire v14457dc;
  wire v14457dd;
  wire v14457de;
  wire v14457df;
  wire v14457e0;
  wire v14457e1;
  wire v14457e2;
  wire v14457e3;
  wire v14457e4;
  wire v14457e9;
  wire v14457ea;
  wire v14457eb;
  wire v14457ec;
  wire v14457ed;
  wire v14457ee;
  wire v14457ef;
  wire v14457f0;
  wire v14457f1;
  wire v14457f2;
  wire v14457f3;
  wire v14457f4;
  wire v14457f5;
  wire v14457f6;
  wire v14457f7;
  wire v14457f8;
  wire v14457fd;
  wire v14457fe;
  wire v14457ff;
  wire v1445800;
  wire v1445801;
  wire v1445802;
  wire v1445803;
  wire v1445804;
  wire v1445805;
  wire v1445806;
  wire v1445807;
  wire v1445808;
  wire v1445809;
  wire v144580a;
  wire v144580b;
  wire v144580c;
  wire v144580d;
  wire v144580e;
  wire v144580f;
  wire v1445810;
  wire v1445811;
  wire v1445812;
  wire v1445813;
  wire v1445814;
  wire v1445815;
  wire v1445816;
  wire v1445817;
  wire v1445818;
  wire v1445819;
  wire v144581a;
  wire v144581b;
  wire v144581c;
  wire v144581d;
  wire v144581e;
  wire v144581f;
  wire v1445820;
  wire v1445821;
  wire v1445822;
  wire v1445823;
  wire v1445824;
  wire v1445825;
  wire v1445826;
  wire v1445827;
  wire v1445828;
  wire v1445829;
  wire v144582a;
  wire v144582b;
  wire v144582c;
  wire v144582d;
  wire v144582e;
  wire v144582f;
  wire v1445830;
  wire v1445831;
  wire v1445832;
  wire v1445833;
  wire v1445834;
  wire v1445835;
  wire v1445836;
  wire v1445837;
  wire v1445838;
  wire v1445839;
  wire v144583a;
  wire v144583b;
  wire v144583c;
  wire v144583d;
  wire v144583e;
  wire v144583f;
  wire v1445840;
  wire v1445841;
  wire v1445842;
  wire v1445843;
  wire v1445844;
  wire v1445845;
  wire v1445846;
  wire v1445847;
  wire v1445848;
  wire v144584c;
  wire v144584d;
  wire v144584e;
  wire v144584f;
  wire v1445850;
  wire v1445851;
  wire v1445852;
  wire v1445853;
  wire v1445854;
  wire v1445855;
  wire v1445856;
  wire v1445857;
  wire v1445858;
  wire v1445859;
  wire v144585a;
  wire v144585b;
  wire v144585c;
  wire v1445860;
  wire v1445861;
  wire v1445862;
  wire v1445863;
  wire v1445864;
  wire v1445865;
  wire v1445866;
  wire v1445867;
  wire v1445868;
  wire v1445869;
  wire v144586a;
  wire v144586b;
  wire v144586c;
  wire v144586d;
  wire v144586e;
  wire v144586f;
  wire v1445870;
  wire v1445871;
  wire v1445872;
  wire v1445873;
  wire v1445874;
  wire v1445875;
  wire v1445876;
  wire v1445877;
  wire v1445878;
  wire v1445879;
  wire v144587a;
  wire v144587b;
  wire v144587c;
  wire v144587d;
  wire v144587e;
  wire v144587f;
  wire v1445880;
  wire v1445881;
  wire v1445882;
  wire v1445883;
  wire v1445884;
  wire v1445885;
  wire v1445886;
  wire v1445887;
  wire v1445888;
  wire v1445889;
  wire v144588a;
  wire v144588b;
  wire v144588c;
  wire v144588d;
  wire v144588e;
  wire v144588f;
  wire v1445890;
  wire v1445891;
  wire v1445892;
  wire v1445893;
  wire v1445894;
  wire v1445895;
  wire v1445896;
  wire v1445897;
  wire v1445898;
  wire v1445899;
  wire v144589a;
  wire v144589b;
  wire v144589c;
  wire v144589d;
  wire v144589e;
  wire v144589f;
  wire v14458a0;
  wire v14458a1;
  wire v14458a2;
  wire v14458a3;
  wire v14458a4;
  wire v14458a5;
  wire v14458a6;
  wire v14458a7;
  wire v14458a8;
  wire v14458a9;
  wire v14458aa;
  wire v14458ab;
  wire v14458ac;
  wire v14458ad;
  wire v14458ae;
  wire v14458af;
  wire v14458b0;
  wire v14458b1;
  wire v14458b2;
  wire v14458b3;
  wire v14458b4;
  wire v14458b5;
  wire v14458b6;
  wire v14458b7;
  wire v14458b8;
  wire v14458b9;
  wire v14458bd;
  wire v14458be;
  wire v14458bf;
  wire v14458c0;
  wire v14458c1;
  wire v14458c2;
  wire v14458c3;
  wire v14458c4;
  wire v14458c5;
  wire v14458c6;
  wire v14458c7;
  wire v14458cb;
  wire v14458cc;
  wire v14458cd;
  wire v14458ce;
  wire v14458cf;
  wire v14458d0;
  wire v14458d1;
  wire v14458d2;
  wire v14458d3;
  wire v14458d4;
  wire v14458d5;
  wire v14458d6;
  wire v14458d7;
  wire v14458d8;
  wire v14458d9;
  wire v14458da;
  wire v14458db;
  wire v14458dc;
  wire v14458dd;
  wire v14458de;
  wire v14458df;
  wire v14458e0;
  wire v14458e1;
  wire v14458e2;
  wire v14458e3;
  wire v14458e4;
  wire v14458e5;
  wire v14458e6;
  wire v14458e7;
  wire v14458e8;
  wire v14458e9;
  wire v14458ea;
  wire v14458eb;
  wire v14458ec;
  wire v14458ed;
  wire v14458ee;
  wire v14458ef;
  wire v14458f0;
  wire v14458f1;
  wire v14458f2;
  wire v14458f3;
  wire v14458f4;
  wire v14458f5;
  wire v14458f6;
  wire v14458f7;
  wire v14458f8;
  wire v14458f9;
  wire v14458fa;
  wire v14458fb;
  wire v14458fc;
  wire v14458fd;
  wire v14458fe;
  wire v14458ff;
  wire v1445900;
  wire v1445901;
  wire v1445902;
  wire v1445903;
  wire v1445904;
  wire v1445905;
  wire v1445906;
  wire v1445907;
  wire v1445908;
  wire v1445909;
  wire v144590a;
  wire v144590b;
  wire v144590c;
  wire v144590d;
  wire v144590e;
  wire v144590f;
  wire v1445910;
  wire v1445911;
  wire v1445912;
  wire v1445913;
  wire v1445914;
  wire v1445915;
  wire v1445916;
  wire v1445917;
  wire v1445918;
  wire v1445919;
  wire v144591a;
  wire v144591b;
  wire v144591c;
  wire v144591d;
  wire v144591e;
  wire v144591f;
  wire v1445920;
  wire v1445921;
  wire v1445922;
  wire v1445923;
  wire v1445924;
  wire v1445925;
  wire v1445926;
  wire v1445927;
  wire v1445928;
  wire v1445929;
  wire v144592a;
  wire v144598e;
  wire v144598f;
  wire v1445990;
  wire v1445991;
  wire v1445992;
  wire v1445993;
  wire v1445994;
  wire v1445995;
  wire v1445996;
  wire v1445997;
  wire v1445998;
  wire v1445999;
  wire v144599a;
  wire v144599b;
  wire v144599c;
  wire v144599d;
  wire v144599e;
  wire v144599f;
  wire v14459a0;
  wire v14459a1;
  wire v14459a2;
  wire v14459a3;
  wire v14459a4;
  wire v14459a5;
  wire v14459a6;
  wire v14459a7;
  wire v14459a8;
  wire v14459a9;
  wire v14459aa;
  wire v14459ab;
  wire v14459ac;
  wire v14459ad;
  wire v14459ae;
  wire v14459af;
  wire v14459b0;
  wire v14459b1;
  wire v14459b2;
  wire v14459b3;
  wire v14459b4;
  wire v14459b5;
  wire v14459b6;
  wire v14459b7;
  wire v14459b8;
  wire v14459b9;
  wire v14459ba;
  wire v14459bb;
  wire v14459bc;
  wire v14459bd;
  wire v14459be;
  wire v14459bf;
  wire v14459c0;
  wire v14459c1;
  wire v14459c2;
  wire v14459c3;
  wire v14459c4;
  wire v14459c5;
  wire v14459c6;
  wire v14459c7;
  wire v14459c8;
  wire v14459c9;
  wire v14459ca;
  wire v14459cb;
  wire v14459cc;
  wire v14459cd;
  wire v14459ce;
  wire v14459cf;
  wire v14459d0;
  wire v14459d1;
  wire v14459d2;
  wire v14459d3;
  wire v14459d4;
  wire v14459d5;
  wire v14459d6;
  wire v14459d7;
  wire v14459d8;
  wire v14459d9;
  wire v14459da;
  wire v14459db;
  wire v14459dc;
  wire v14459dd;
  wire v14459de;
  wire v14459df;
  wire v14459e0;
  wire v14459e1;
  wire v14459e2;
  wire v14459e3;
  wire v14459e4;
  wire v14459e5;
  wire v14459e6;
  wire v14459e7;
  wire v14459e8;
  wire v14459e9;
  wire v14459ea;
  wire v14459eb;
  wire v14459ec;
  wire v14459ed;
  wire v14459ee;
  wire v14459ef;
  wire v14459f0;
  wire v14459f1;
  wire v14459f2;
  wire v14459f3;
  wire v14459f4;
  wire v14459f5;
  wire v14459f6;
  wire v14459f7;
  wire v14459f8;
  wire v14459f9;
  wire v14459fa;
  wire v14459fb;
  wire v14459fc;
  wire v14459fd;
  wire v14459fe;
  wire v14459ff;
  wire v1445a00;
  wire v1445a01;
  wire v1445a02;
  wire v1445a03;
  wire v1445a04;
  wire v1445a05;
  wire v1445a06;
  wire v1445a07;
  wire v1445a08;
  wire v1445a09;
  wire v1445a0a;
  wire v1445a0b;
  wire v1445a0c;
  wire v1445a0d;
  wire v1445a0e;
  wire v1445a0f;
  wire v1445a10;
  wire v1445a11;
  wire v1445a12;
  wire v1445a13;
  wire v1445a14;
  wire v1445a15;
  wire v1445a16;
  wire v1445a17;
  wire v1445a18;
  wire v1445a19;
  wire v1445a1a;
  wire v1445a1b;
  wire v1445a1c;
  wire v1445a1d;
  wire v1445a1e;
  wire v1445a1f;
  wire v1445a20;
  wire v1445a21;
  wire v1445a22;
  wire v1445a23;
  wire v1445a24;
  wire v1445a25;
  wire v1445a26;
  wire v1445a27;
  wire v1445a28;
  wire v1445a29;
  wire v1445a2a;
  wire v1445a2b;
  wire v1445a2c;
  wire v1445a2d;
  wire v1445a2e;
  wire v1445a2f;
  wire v1445a30;
  wire v1445a31;
  wire v1445a32;
  wire v1445a33;
  wire v1445a34;
  wire v1445a35;
  wire v1445a36;
  wire v1445a37;
  wire v1445a38;
  wire v1445a39;
  wire v1445a3a;
  wire v1445a3b;
  wire v1445a3c;
  wire v1445a3d;
  wire v1445a3e;
  wire v1445a3f;
  wire v1445a40;
  wire v1445a41;
  wire v1445a42;
  wire v1445a43;
  wire v1445a44;
  wire v1445a45;
  wire v1445a46;
  wire v1445a47;
  wire v1445a48;
  wire v1445a49;
  wire v1445a4a;
  wire v1445a4b;
  wire v1445a4c;
  wire v1445a4d;
  wire v1445a4e;
  wire v1445a4f;
  wire v1445a50;
  wire v1445a51;
  wire v1445a52;
  wire v1445a53;
  wire v1445a54;
  wire v1445a55;
  wire v1445a56;
  wire v1445a57;
  wire v1445a58;
  wire v1445a59;
  wire v1445a5a;
  wire v1445a5b;
  wire v1445a5c;
  wire v1445a5d;
  wire v1445a5e;
  wire v1445a5f;
  wire v1445a60;
  wire v1445a61;
  wire v1445a62;
  wire v1445a63;
  wire v1445a64;
  wire v1445a65;
  wire v1445a66;
  wire v1445a67;
  wire v1445a68;
  wire v1445a69;
  wire v1445a6a;
  wire v1445a6b;
  wire v1445a6c;
  wire v1445a6d;
  wire v1445a6e;
  wire v1445a6f;
  wire v1445a70;
  wire v1445a71;
  wire v1445a72;
  wire v1445a73;
  wire v1445a74;
  wire v1445a75;
  wire v1445a76;
  wire v1445a77;
  wire v1445a78;
  wire v1445a79;
  wire v1445a7a;
  wire v1445a7b;
  wire v1445a7c;
  wire v1445a7d;
  wire v1445a7e;
  wire v1445a7f;
  wire v1445a80;
  wire v1445a81;
  wire v1445a82;
  wire v1445a83;
  wire v1445a84;
  wire v1445a85;
  wire v1445a86;
  wire v1445a87;
  wire v1445a88;
  wire v1445a89;
  wire v1445a8a;
  wire v1445a8b;
  wire v1445a8c;
  wire v1445a8d;
  wire v1445a8e;
  wire v1445a8f;
  wire v1445a90;
  wire v1445a91;
  wire v1445a92;
  wire v1445a93;
  wire v1445a94;
  wire v1445a95;
  wire v1445a96;
  wire v1445a97;
  wire v1445a98;
  wire v1445a99;
  wire v1445a9a;
  wire v1445a9b;
  wire v1445a9c;
  wire v1445a9d;
  wire v1445a9e;
  wire v1445a9f;
  wire v1445aa0;
  wire v1445aa1;
  wire v1445aa2;
  wire v1445aa3;
  wire v1445aa4;
  wire v1445aa5;
  wire v1445aa6;
  wire v1445aa7;
  wire v1445aa8;
  wire v1445aa9;
  wire v1445aaa;
  wire v1445aab;
  wire v1445aac;
  wire v1445aad;
  wire v1445aae;
  wire v1445aaf;
  wire v1445ab0;
  wire v1445ab1;
  wire v1445ab6;
  wire v1445ab7;
  wire v1445ab8;
  wire v1445ab9;
  wire v1445aba;
  wire v1445abb;
  wire v1445abc;
  wire v1445abd;
  wire v1445abe;
  wire v1445abf;
  wire v1445ac0;
  wire v1445ac1;
  wire v1445ac2;
  wire v1445ac3;
  wire v1445ac4;
  wire v1445ac5;
  wire v1445ac6;
  wire v1445ac7;
  wire v1445ac8;
  wire v1445ac9;
  wire v1445aca;
  wire v1445acb;
  wire v1445acc;
  wire v1445acd;
  wire v1445ace;
  wire v1445acf;
  wire v1445ad0;
  wire v1445ad1;
  wire v1445ad2;
  wire v1445ad3;
  wire v1445ad4;
  wire v1445ad5;
  wire v1445ad6;
  wire v1445ad7;
  wire v1445ad8;
  wire v1445ad9;
  wire v1445ada;
  wire v1445adb;
  wire v1445adc;
  wire v1445add;
  wire v1445ade;
  wire v1445adf;
  wire v1445ae0;
  wire v1445ae1;
  wire v1445ae2;
  wire v1445ae3;
  wire v1445ae4;
  wire v1445ae5;
  wire v1445ae6;
  wire v1445ae7;
  wire v1445ae8;
  wire v1445ae9;
  wire v1445aea;
  wire v1445aeb;
  wire v1445aec;
  wire v1445aed;
  wire v1445aee;
  wire v1445aef;
  wire v1445af0;
  wire v1445af1;
  wire v1445af2;
  wire v1445af3;
  wire v1445af4;
  wire v1445af5;
  wire v1445af6;
  wire v1445af7;
  wire v1445af8;
  wire v1445af9;
  wire v1445afa;
  wire v1445afb;
  wire v1445afc;
  wire v1445afd;
  wire v1445afe;
  wire v1445aff;
  wire v1445b00;
  wire v1445b01;
  wire v1445b02;
  wire v1445b03;
  wire v1445b04;
  wire v1445b05;
  wire v1445b06;
  wire v1445b07;
  wire v1445b08;
  wire v1445b09;
  wire v1445b0a;
  wire v1445b0b;
  wire v1445b0c;
  wire v1445b0d;
  wire v1445b0e;
  wire v1445b0f;
  wire v1445b10;
  wire v1445b11;
  wire v1445b12;
  wire v1445b13;
  wire v1445b14;
  wire v1445b15;
  wire v1445b16;
  wire v1445b17;
  wire v1445b18;
  wire v1445b19;
  wire v1445b1a;
  wire v1445b1b;
  wire v1445b1c;
  wire v1445b1d;
  wire v1445b1e;
  wire v1445b1f;
  wire v1445b20;
  wire v1445b21;
  wire v1445b22;
  wire v1445b23;
  wire v1445b24;
  wire v1445b25;
  wire v1445b26;
  wire v1445b27;
  wire v1445b28;
  wire v1445b29;
  wire v1445b2a;
  wire v1445b2b;
  wire v1445b2f;
  wire v1445b30;
  wire v1445b31;
  wire v1445b32;
  wire v1445b33;
  wire v1445b34;
  wire v1445b35;
  wire v1445b36;
  wire v1445b37;
  wire v1445b38;
  wire v1445b39;
  wire v1445b3d;
  wire v1445b3e;
  wire v1445b3f;
  wire v1445b40;
  wire v1445b41;
  wire v1445b42;
  wire v1445b43;
  wire v1445b44;
  wire v1445b45;
  wire v1445b46;
  wire v1445b47;
  wire v1445b48;
  wire v1445b4d;
  wire v1445b4e;
  wire v1445b4f;
  wire v1445b50;
  wire v1445353;
  wire v1445354;
  wire v1445355;
  wire v1445356;
  wire v1445357;
  wire v1445358;
  wire v144535d;
  wire v144535e;
  wire v144535f;
  wire v1445360;
  wire v1445361;
  wire v1445362;
  wire v1445363;
  wire v1445364;
  wire v1445365;
  wire v1445366;
  wire v1445367;
  wire v1445368;
  wire v1445369;
  wire v144536a;
  wire v144536b;
  wire v144536c;
  wire v144536d;
  wire v144536e;
  wire v144536f;
  wire v1445370;
  wire v1445371;
  wire v1445372;
  wire v1445373;
  wire v1445374;
  wire v1445375;
  wire v1445376;
  wire v1445377;
  wire v1445378;
  wire v1445379;
  wire v144537a;
  wire v144537b;
  wire v144537c;
  wire v144537d;
  wire v144537e;
  wire v144537f;
  wire v1445383;
  wire v1445384;
  wire v1445385;
  wire v1445386;
  wire v1445387;
  wire v1445388;
  wire v1445389;
  wire v144538a;
  wire v144538b;
  wire v144538c;
  wire v144538d;
  wire v1445391;
  wire v1445392;
  wire v1445393;
  wire v1445394;
  wire v1445395;
  wire v1445396;
  wire v1445397;
  wire v1445398;
  wire v1445399;
  wire v144539a;
  wire v144539b;
  wire v144539c;
  wire v144539d;
  wire v144539e;
  wire v144539f;
  wire v14453a0;
  wire v14453a1;
  wire v14453a2;
  wire v14453a3;
  wire v14453a4;
  wire v14453a5;
  wire v14453a6;
  wire v14453a7;
  wire v14453a8;
  wire v14453a9;
  wire v14453aa;
  wire v14453ab;
  wire v14453ac;
  wire v14453ad;
  wire v14453ae;
  wire v14453af;
  wire v14453b0;
  wire v14453b1;
  wire v14453b2;
  wire v14453b3;
  wire v14453b4;
  wire v14453b5;
  wire v14453b6;
  wire v14453b7;
  wire v14453b8;
  wire v14453b9;
  wire v14453ba;
  wire v14453bb;
  wire v14453bc;
  wire v14453bd;
  wire v14453be;
  wire v14453bf;
  wire v14453c0;
  wire v14453c1;
  wire v14453c2;
  wire v14453c3;
  wire v14453c4;
  wire v14453c5;
  wire v14453c6;
  wire v14453c7;
  wire v14453c8;
  wire v14453e1;
  wire v14453e2;
  wire v14453e3;
  wire v14453e4;
  wire v14453e5;
  wire v14453e6;
  wire v14453e7;
  wire v14453e8;
  wire v14453e9;
  wire v14453ea;
  wire v14453eb;
  wire v14453ec;
  wire v14453ed;
  wire v14453ee;
  wire v14453ef;
  wire v14453f0;
  wire v14453f1;
  wire v14453f2;
  wire v14453f3;
  wire v14453f4;
  wire v14453f5;
  wire v14453f6;
  wire v14453f7;
  wire v14453f8;
  wire v14453f9;
  wire v14453fa;
  wire v14453fb;
  wire v14453fc;
  wire v14453fd;
  wire v14453fe;
  wire v14453ff;
  wire v1445400;
  wire v1445401;
  wire v1445402;
  wire v1445403;
  wire v1445404;
  wire v1445405;
  wire v1445406;
  wire v1445407;
  wire v1445408;
  wire v1445409;
  wire v144540a;
  wire v144540b;
  wire v1445411;
  wire v1445412;
  wire v1445413;
  wire v1445414;
  wire v1445415;
  wire v1445416;
  wire v1445417;
  wire v1445418;
  wire v1445419;
  wire v144541a;
  wire v144541b;
  wire v144541c;
  wire v144541d;
  wire v144541e;
  wire v144541f;
  wire v1445420;
  wire v1445421;
  wire v1445422;
  wire v1445423;
  wire v1445424;
  wire v1445425;
  wire v1445426;
  wire v1445427;
  wire v1445428;
  wire v1445429;
  wire v144542a;
  wire v144542b;
  wire v144542c;
  wire v144542d;
  wire v144542e;
  wire v144542f;
  wire v1445430;
  wire v1445431;
  wire v1445432;
  wire v1445433;
  wire v1445434;
  wire v1445435;
  wire v1445436;
  wire v1445437;
  wire v1445438;
  wire v1445439;
  wire v144543a;
  wire v144543b;
  wire v144543c;
  wire v144543d;
  wire v144543e;
  wire v144543f;
  wire v1445440;
  wire v1445441;
  wire v1445442;
  wire v1445443;
  wire v1445444;
  wire v1445445;
  wire v1445446;
  wire v1445447;
  wire v1445448;
  wire v1445449;
  wire v144544a;
  wire v144544b;
  wire v144544c;
  wire v144544d;
  wire v144544e;
  wire v144544f;
  wire v1445450;
  wire v1445451;
  wire v1445452;
  wire v1445453;
  wire v1445454;
  wire v1445455;
  wire v1445456;
  wire v1445457;
  wire v1445458;
  wire v1445459;
  wire v144545a;
  wire v144545b;
  wire v144545c;
  wire v144545d;
  wire v144545e;
  wire v144545f;
  wire v1445468;
  wire v1445469;
  wire v144546b;
  wire v144546c;
  wire v144546d;
  wire v144546e;
  wire v144546f;
  wire v1445470;
  wire v1445471;
  wire v1445472;
  wire v1445473;
  wire v1445479;
  wire v144547a;
  wire v144547c;
  wire v144547d;
  wire v144547e;
  wire v144547f;
  wire v1445480;
  wire v1445481;
  wire v1445482;
  wire v1445489;
  wire v144548a;
  wire v144548c;
  wire v144548d;
  wire v144548e;
  wire v144548f;
  wire v1445490;
  wire v1445491;
  wire v1445492;
  wire v1445493;
  wire v1445494;
  wire v1445498;
  wire v1445499;
  wire v144549a;
  wire v144549b;
  wire v144549c;
  wire v144549d;
  wire v144549e;
  wire v144549f;
  wire v14454a3;
  wire v14454a4;
  wire v14454a6;
  wire v14454a7;
  wire v14454a8;
  wire v14454e8;
  wire v14454e9;
  wire v14454ea;
  wire v14454eb;
  wire v14454ec;
  wire v14454ed;
  wire v14454ee;
  wire v14454ef;
  wire v14454f0;
  wire v14454f1;
  wire v14454f2;
  wire v14454f3;
  wire v14454f7;
  wire v14454f8;
  wire v14454f9;
  wire v14454fa;
  wire v14454fb;
  wire v14454fc;
  wire v14454fd;
  wire v14454fe;
  wire v14454ff;
  wire v1445500;
  wire v1445501;
  wire v1445502;
  wire v1445503;
  wire v1445504;
  wire v1445505;
  wire v1445506;
  wire v1445507;
  wire v1445508;
  wire v1445509;
  wire v144550a;
  wire v144550b;
  wire v144550c;
  wire v144550d;
  wire v144550e;
  wire v144550f;
  wire v1445510;
  wire v1445511;
  wire v1445512;
  wire v1445513;
  wire v1445514;
  wire v1445515;
  wire v1445516;
  wire v1445517;
  wire v1445518;
  wire v1445519;
  wire v144551a;
  wire v144551b;
  wire v144551c;
  wire v144551d;
  wire v144551e;
  wire v144551f;
  wire v1445520;
  wire v1445521;
  wire v1445522;
  wire v1445523;
  wire v1445524;
  wire v1445527;
  wire v1445528;
  wire v1445529;
  wire v144552a;
  wire v144552b;
  wire v144552c;
  wire v144552d;
  wire v144552e;
  wire v144552f;
  wire v1445530;
  wire v1445531;
  wire v1445532;
  wire v1445533;
  wire v1445534;
  wire v1445535;
  wire v1445536;
  wire v1445537;
  wire v1445538;
  wire v144553b;
  wire v144553c;
  wire v144553d;
  wire v144553e;
  wire v144553f;
  wire v1445540;
  wire v1445541;
  wire v1445542;
  wire v1445543;
  wire v1445544;
  wire v1445545;
  wire v1445546;
  wire v1445547;
  wire v1445548;
  wire v1445549;
  wire v144554a;
  wire v144554b;
  wire v144554c;
  wire v144554d;
  wire v144554e;
  wire v144554f;
  wire v1445550;
  wire v1445551;
  wire v1445552;
  wire v1445553;
  wire v1445554;
  wire v1445555;
  wire v1445556;
  wire v1445557;
  wire v1445558;
  wire v114a22f;
  wire v845572;
  wire v114a230;
  wire v114a231;
  wire v114a232;
  wire v114a233;
  wire v114a3be;
  wire v114a3bf;
  wire f2f21a;
  wire f2f21b;
  wire f2f21c;
  wire f2f21d;
  wire f2f21e;
  wire f2f21f;
  wire f2f220;
  wire f2f221;
  wire f2f222;
  wire f2f223;
  wire f2f224;
  wire f2f225;
  wire f2f226;
  wire f2f227;
  wire f2f228;
  wire f2f229;
  wire f2f22a;
  wire f2f22b;
  wire f2f22c;
  wire f2f22d;
  wire f2f22e;
  wire f2f22f;
  wire f2f230;
  wire f2f231;
  wire f2f232;
  wire f2f233;
  wire f2f234;
  wire f2f235;
  wire f2f236;
  wire f2f237;
  wire f2f238;
  wire f2f239;
  wire f2f23a;
  wire f2f23b;
  wire f2f23c;
  wire f2f23d;
  wire f2f27e;
  wire f2f27f;
  wire f2f280;
  wire f2f281;
  wire f2f282;
  wire f2f283;
  wire f2f284;
  wire f2f285;
  wire f2f286;
  wire f2f287;
  wire f2f288;
  wire f2f289;
  wire f2f28a;
  wire f2f28b;
  wire f2f28c;
  wire f2f28d;
  wire f2f28e;
  wire f2f28f;
  wire f2f290;
  wire f2f291;
  wire f2f292;
  wire f2f293;
  wire f2f294;
  wire f2f295;
  wire f2f296;
  wire f2f297;
  wire f2f298;
  wire f2f299;
  wire f2f29a;
  wire f2f29b;
  wire f2f29c;
  wire f2f29d;
  wire f2f29e;
  wire f2f29f;
  wire f2f2a0;
  wire f2f2a1;
  wire f2f2a2;
  wire f2f2a3;
  wire f2f2a4;
  wire f2f2a5;
  wire f2f2a6;
  wire f2f2a7;
  wire f2f2a8;
  wire f2f2a9;
  wire f2f2aa;
  wire f2f2ab;
  wire f2f2ac;
  wire f2f2ad;
  wire f2f2ae;
  wire f2f2af;
  wire f2f2b0;
  wire f2f2b1;
  wire f2f2c8;
  wire f2f2c9;
  wire f2f2ca;
  wire f2f2cb;
  wire f2f2cc;
  wire f2f2cd;
  wire f2f2ce;
  wire f2f2cf;
  wire f2f2d0;
  wire f2f2d1;
  wire f2f2d2;
  wire f2f2d3;
  wire f2f2d4;
  wire f2f2d5;
  wire f2f2d6;
  wire f2f2d7;
  wire f2f2d8;
  wire f2f2d9;
  wire f2f2da;
  wire f2f2db;
  wire f2f2dc;
  wire f2f2dd;
  wire f2f2de;
  wire f2f2df;
  wire f2f2e0;
  wire f2f2e1;
  wire f2f2e2;
  wire f2f2e3;
  wire f2f2e4;
  wire f2f2e5;
  wire f2f2e6;
  wire f2f2e7;
  wire f2f2e8;
  wire f2f2e9;
  wire f2f2ea;
  wire f2f2eb;
  wire f2f2ec;
  wire f2f2ed;
  wire f2f2ee;
  wire f2f2ef;
  wire f2f2f0;
  wire f2f2f1;
  wire f2f327;
  wire f2f328;
  wire f2f329;
  wire f2f32a;
  wire f2f32b;
  wire f2f32c;
  wire f2f32d;
  wire f2f32e;
  wire f2f32f;
  wire f2f330;
  wire f2f331;
  wire f2f332;
  wire f2f333;
  wire f2f334;
  wire f2f335;
  wire f2f336;
  wire f2f337;
  wire f2f338;
  wire f2f339;
  wire f2f33a;
  wire f2f33b;
  wire f2f33c;
  wire f2f33d;
  wire f2f33e;
  wire f2f33f;
  wire f2f340;
  wire f2f341;
  wire f2f342;
  wire f2f343;
  wire f2f344;
  wire f2f345;
  wire f2f346;
  wire f2f347;
  wire f2f34a;
  wire f2f34b;
  wire f2f34c;
  wire f2f34d;
  wire f2f34e;
  wire f2f34f;
  wire f2f350;
  wire f2f351;
  wire f2f352;
  wire f2f353;
  wire f2f354;
  wire f2f355;
  wire f2f356;
  wire f2f357;
  wire f2f358;
  wire f2f359;
  wire f2f35a;
  wire f2f35b;
  wire f2f35c;
  wire f2f35d;
  wire f2f35e;
  wire f2f35f;
  wire f2f360;
  wire f2f361;
  wire f2f362;
  wire f2f363;
  wire f2f367;
  wire f2f368;
  wire f2f369;
  wire f2f36a;
  wire f2f36e;
  wire f2f36f;
  wire f2f370;
  wire f2f371;
  wire f2f372;
  wire f2f373;
  wire f2f374;
  wire f2f375;
  wire f2f376;
  wire f2f377;
  wire f2f378;
  wire f2f379;
  wire f2f37a;
  wire f2f37b;
  wire f2f37c;
  wire f2f37d;
  wire f2f37e;
  wire f2f37f;
  wire f2f380;
  wire f2f381;
  wire f2f382;
  wire f2f383;
  wire f2f384;
  wire f2f385;
  wire f2f386;
  wire f2f387;
  wire f2f388;
  wire f2f389;
  wire f2f38a;
  wire f2f38b;
  wire f2f38c;
  wire f2f38d;
  wire f2f38e;
  wire f2f38f;
  wire f2f390;
  wire f2f391;
  wire f2f392;
  wire f2f393;
  wire f2f394;
  wire f2f395;
  wire f2f396;
  wire f2f397;
  wire f2f398;
  wire f2f399;
  wire f2f39a;
  wire f2f39b;
  wire f2f39c;
  wire f2f39d;
  wire f2f39e;
  wire f2f39f;
  wire f2f3a0;
  wire f2f3a1;
  wire f2f3a2;
  wire f2f3a3;
  wire f2f3a4;
  wire f2f3a5;
  wire f2f3a6;
  wire f2f3a7;
  wire f2f3a8;
  wire f2f3a9;
  wire f2f3aa;
  wire f2f3ab;
  wire f2f3ac;
  wire f2f3ad;
  wire f2f3ae;
  wire f2f3af;
  wire f2f3b0;
  wire f2f3b1;
  wire f2f3b2;
  wire f2f3b3;
  wire f2f3b4;
  wire f2f3b5;
  wire f2f3b6;
  wire f2f3b7;
  wire f2f3b8;
  wire f2f3b9;
  wire f2f3ba;
  wire f2f3bb;
  wire f2f3bc;
  wire f2f3bd;
  wire f2f3be;
  wire f2f3bf;
  wire f2f3c0;
  wire f2f3c1;
  wire f2f3c2;
  wire f2f3c3;
  wire f2f3c4;
  wire f2f3c5;
  wire f2f3c6;
  wire f2f3c7;
  wire f2f3c8;
  wire f2f3c9;
  wire f2f3ca;
  wire f2f3cb;
  wire f2f3cc;
  wire f2f3cd;
  wire f2f3ce;
  wire f2f3cf;
  wire f2f3d0;
  wire f2f3d1;
  wire f2f3d2;
  wire f2f3d3;
  wire f2f3d4;
  wire f2f3d5;
  wire f2f3d6;
  wire f2f3d7;
  wire f2f3d8;
  wire f2f3d9;
  wire f2f3da;
  wire f2f3db;
  wire f2f3dc;
  wire f2f3dd;
  wire f2f3de;
  wire f2f3df;
  wire f2f3e0;
  wire f2f3e1;
  wire f2f3e2;
  wire f2f3e3;
  wire f2f3e4;
  wire f2f3e5;
  wire f2f3e6;
  wire f2f3e7;
  wire f2f3e8;
  wire f2f3e9;
  wire f2f3ea;
  wire f2f3eb;
  wire f2f3ec;
  wire f2f3ed;
  wire f2f3ee;
  wire f2f3ef;
  wire f2f3f0;
  wire f2f3f1;
  wire f2f3f2;
  wire f2f3f3;
  wire f2f3f4;
  wire f2f3f5;
  wire f2f3f6;
  wire f2f3f7;
  wire f2f3f8;
  wire f2f3f9;
  wire f2f3fa;
  wire f2f3fb;
  wire f2f3fc;
  wire f2f3fd;
  wire f2f3fe;
  wire f2f3ff;
  wire f2f400;
  wire f2f401;
  wire f2f402;
  wire f2f403;
  wire f2f404;
  wire f2f405;
  wire f2f406;
  wire f2f407;
  wire f2f408;
  wire f2f409;
  wire f2f40a;
  wire f2f40b;
  wire f2f40c;
  wire f2f40d;
  wire f2f40e;
  wire f2f40f;
  wire f2f410;
  wire f2f411;
  wire f2f412;
  wire f2f413;
  wire f2f414;
  wire f2f415;
  wire f2f416;
  wire f2f417;
  wire f2f418;
  wire f2f419;
  wire f2f41a;
  wire f2f41b;
  wire f2f41c;
  wire f2f41d;
  wire f2f41e;
  wire f2f41f;
  wire f2f420;
  wire f2f421;
  wire f2f422;
  wire f2f423;
  wire f2f424;
  wire f2f425;
  wire f2f426;
  wire f2f427;
  wire f2f428;
  wire f2f429;
  wire f2f42a;
  wire f2f42b;
  wire f2f42c;
  wire f2f42d;
  wire f2f42e;
  wire f2f42f;
  wire f2f430;
  wire f2f431;
  wire f2f432;
  wire f2f433;
  wire f2f434;
  wire f2f435;
  wire f2f436;
  wire f2f437;
  wire f2f438;
  wire f2f439;
  wire f2f43a;
  wire f2f43b;
  wire f2f43c;
  wire f2f43d;
  wire f2f43e;
  wire f2f43f;
  wire f2f440;
  wire f2f441;
  wire f2f442;
  wire f2f443;
  wire f2f444;
  wire f2f445;
  wire f2f446;
  wire f2f447;
  wire f2f448;
  wire f2f449;
  wire f2f44a;
  wire f2f44b;
  wire f2f44c;
  wire f2f44d;
  wire f2f44e;
  wire f2f44f;
  wire f2f450;
  wire f2f451;
  wire f2f452;
  wire f2f453;
  wire f2f454;
  wire f2f455;
  wire f2f456;
  wire f2f457;
  wire f2f458;
  wire f2f459;
  wire f2f45a;
  wire f2f45b;
  wire f2f45c;
  wire f2f45d;
  wire f2f45e;
  wire f2f45f;
  wire f2f460;
  wire f2f461;
  wire f2f462;
  wire f2f4a7;
  wire f2f4a8;
  wire f2f4a9;
  wire f2f4aa;
  wire f2f4ab;
  wire f2f4ac;
  wire v146af2e;
  wire f2f4ad;
  wire f2f4ae;
  wire f2f4af;
  wire f2f4b0;
  wire f2f4b1;
  wire f2f4b2;
  wire f2f4b3;
  wire f2f4b4;
  wire f2f4b5;
  wire f2f4b6;
  wire f2f4b9;
  wire f2f4ba;
  wire f2f4be;
  wire f2f4bf;
  wire f2f4c2;
  wire f2f4c3;
  wire f2f4c4;
  wire f2f519;
  wire f2f51a;
  wire f2f52c;
  wire f2f52d;
  wire f2f52e;
  wire f2f538;
  wire f2f539;
  wire f2f53a;
  wire f2f53b;
  wire f2f53c;
  wire f2f53d;
  wire f2f53e;
  wire f2ed8d;
  wire f2ed8e;
  wire f2ed8f;
  wire f2ed90;
  wire f2ed91;
  wire f2ed92;
  wire f2ed93;
  wire f2ed94;
  wire f2ed95;
  wire f2ed96;
  wire f2ed97;
  wire f2ed98;
  wire f2ed99;
  wire f2ed9a;
  wire f2ed9b;
  wire f2ed9c;
  wire f2ed9d;
  wire f2ed9e;
  wire f2ed9f;
  wire f2eda0;
  wire f2eda1;
  wire f2eda2;
  wire f2eda3;
  wire f2eda4;
  wire f2eda5;
  wire f2ec20;
  wire f2ec21;
  wire f2ec22;
  wire f2ec23;
  wire f2ec24;
  wire f2ec25;
  wire f2ec26;
  wire f2ec27;
  wire f2e710;
  wire f2e711;
  wire f2e712;
  wire f2e713;
  wire f2e714;
  wire f2e715;
  wire f2e730;
  wire f2e731;
  wire f2e732;
  wire f2e733;
  wire f2e734;
  wire f2e73c;
  wire f2e882;
  wire f2e883;
  wire f2e884;
  wire f2e273;
  wire f2e274;
  wire f2e275;
  wire f2e276;
  wire f2e277;
  wire f2e278;
  wire f2e279;
  wire f2e27a;
  wire f2e27b;
  wire f2e3f6;
  wire f2e3f7;
  wire f2e3f8;
  wire f2e3f9;
  wire f2e3fa;
  wire f2e3fb;
  wire f2e3fc;
  wire f2e3fd;
  wire f2e4c7;
  wire f2e4c8;
  wire f2e4c9;
  wire f2e4ca;
  wire f2e4cb;
  wire f2e4cc;
  wire f2e4cd;
  wire f2e4cf;
  wire f2e4d0;
  wire f2e4d1;
  wire f2e4d2;
  wire f2e4d3;
  wire f2e4d4;
  wire f2e4d5;
  wire f2e4d6;
  wire f2e4d7;
  wire f2e4d8;
  wire f2e4d9;
  wire f2e4da;
  wire f2e4db;
  wire f2e4dc;
  wire f2e4dd;
  wire f2e4de;
  wire f2e4df;
  wire f2e4e0;
  wire f2e4e1;
  wire f2e4e2;
  wire f2e4e3;
  wire f2e4e7;
  wire f2e4e8;
  wire f2e4e9;
  wire f2e4f2;
  wire f2e4f3;
  wire f2e4f4;
  wire f2e4f8;
  wire f2e4f9;
  wire f2e4fa;
  wire f2e4fb;
  wire f2e4fc;
  wire f2e4fd;
  wire f2e4fe;
  wire f2e4ff;
  wire f2e500;
  wire f2e501;
  wire f2e502;
  wire f2e503;
  wire f2e504;
  wire f2e505;
  wire f2e506;
  wire d305d4;
  wire d305d5;
  wire d305d6;
  wire d305d7;
  wire d305d8;
  wire d305d9;
  wire d305da;
  wire d305db;
  wire d305dc;
  wire d305dd;
  wire d305de;
  wire d305df;
  wire d305e0;
  wire d305e1;
  wire d305e2;
  wire d305e3;
  wire d305e4;
  wire d305e5;
  wire v84555e;
  wire d305e6;
  wire d305e7;
  wire d305e9;
  wire d305ea;
  wire d305eb;
  wire d305ec;
  wire d305ed;
  wire d305ee;
  wire d305ef;
  wire d305f0;
  wire d305f1;
  wire d305f2;
  wire d305f3;
  wire d305f4;
  wire d305f5;
  wire d305f6;
  wire v84554e;
  wire d305f7;
  wire d305fb;
  wire d305fc;
  wire d305fd;
  wire v84555a;
  wire d305fe;
  wire d305ff;
  wire d30603;
  wire d30604;
  wire d30605;
  wire d30606;
  wire d30607;
  wire d30608;
  wire d30609;
  wire d3060a;
  wire d3060b;
  wire d3060c;
  wire d3060d;
  wire d3060e;
  wire d3060f;
  wire d30610;
  wire d30611;
  wire d30612;
  wire d30613;
  wire d30614;
  wire d30615;
  wire d30616;
  wire d30617;
  wire d30618;
  wire d30619;
  wire d3061a;
  wire d3061b;
  wire d3061c;
  wire d3061d;
  wire d3061e;
  wire d3061f;
  wire d30620;
  wire d30621;
  wire d30622;
  wire d30623;
  wire d30624;
  wire d30625;
  wire d30626;
  wire d30627;
  wire d30628;
  wire d3062c;
  wire d30630;
  wire d30631;
  wire d30632;
  wire d30633;
  wire d30634;
  wire d30635;
  wire d30636;
  wire d30637;
  wire d30638;
  wire d30639;
  wire d3063a;
  wire d3063b;
  wire d3063c;
  wire d3063d;
  wire d3063e;
  wire d3063f;
  wire d30640;
  wire d30641;
  wire d30642;
  wire d30643;
  wire d30644;
  wire d30645;
  wire d30646;
  wire d30647;
  wire d30648;
  wire d30649;
  wire d3064a;
  wire d3064b;
  wire d3064c;
  wire d3064d;
  wire d3064e;
  wire d3064f;
  wire d30650;
  wire d30651;
  wire d30652;
  wire d30653;
  wire d30654;
  wire d30655;
  wire d30656;
  wire d30657;
  wire d30658;
  wire d30659;
  wire d3065a;
  wire d3065b;
  wire d3065c;
  wire d3065d;
  wire d3065e;
  wire d3065f;
  wire d30660;
  wire d30661;
  wire d30662;
  wire d30663;
  wire d30664;
  wire d30665;
  wire d30666;
  wire d30667;
  wire d30668;
  wire d30669;
  wire d3066a;
  wire d3066b;
  wire d3066c;
  wire d3066d;
  wire d3066e;
  wire d3066f;
  wire d30670;
  wire d30671;
  wire d30672;
  wire d30673;
  wire d30674;
  wire d30675;
  wire d30676;
  wire d30677;
  wire d30678;
  wire d30679;
  wire d3067a;
  wire d3067b;
  wire d3067c;
  wire d3067d;
  wire d3067e;
  wire d3067f;
  wire d30680;
  wire d30681;
  wire d30682;
  wire d30683;
  wire d30684;
  wire d30685;
  wire d30686;
  wire d30687;
  wire v845548;
  wire d30688;
  wire d30689;
  wire d3068a;
  wire d3068b;
  wire d3068c;
  wire d3068d;
  wire d3068e;
  wire v84554a;
  wire d3068f;
  wire d30690;
  wire d30691;
  wire d30692;
  wire d30693;
  wire d30694;
  wire d30695;
  wire d30696;
  wire d30697;
  wire d30698;
  wire d30699;
  wire d3069a;
  wire d3069b;
  wire d3069c;
  wire d3069d;
  wire d3069e;
  wire d3069f;
  wire d306a0;
  wire d306a1;
  wire d306a2;
  wire d306a3;
  wire d306a4;
  wire d306a5;
  wire d306a6;
  wire d306a7;
  wire d306a8;
  wire d306a9;
  wire d306aa;
  wire d306ab;
  wire d306ac;
  wire d306ad;
  wire d306ae;
  wire d306af;
  wire d306b0;
  wire d306b1;
  wire d306b2;
  wire d306b3;
  wire d306b4;
  wire d306b5;
  wire d306b6;
  wire d306b7;
  wire d306b8;
  wire d306b9;
  wire d306ba;
  wire d306bb;
  wire d306bc;
  wire d306bd;
  wire d306be;
  wire d306bf;
  wire d306c0;
  wire d306c1;
  wire d306c2;
  wire d306c3;
  wire d306c4;
  wire d306c5;
  wire d306c6;
  wire d306c7;
  wire d306c8;
  wire d306c9;
  wire d306ca;
  wire d306cb;
  wire d306cc;
  wire d306cd;
  wire d306ce;
  wire d306cf;
  wire d306d0;
  wire d306d1;
  wire d306d2;
  wire d306d3;
  wire d306d4;
  wire d306d5;
  wire d306d6;
  wire d306d7;
  wire d306d8;
  wire d306d9;
  wire d306da;
  wire d306db;
  wire d306dc;
  wire d306dd;
  wire d306de;
  wire d306df;
  wire d306e0;
  wire d306e1;
  wire d306e2;
  wire d306e3;
  wire d306e4;
  wire d306e5;
  wire d306e6;
  wire d306e7;
  wire d306e8;
  wire d306e9;
  wire d306ea;
  wire d306eb;
  wire d306ec;
  wire d306ed;
  wire d306ee;
  wire d306ef;
  wire d306f0;
  wire d306f1;
  wire d306f2;
  wire d306f3;
  wire d306f4;
  wire d306f5;
  wire d306f6;
  wire d306f7;
  wire d306f8;
  wire d306f9;
  wire d306fa;
  wire d306fb;
  wire d306fc;
  wire d306fd;
  wire d306fe;
  wire d306ff;
  wire d30700;
  wire d30701;
  wire d30702;
  wire d30703;
  wire d30704;
  wire d30705;
  wire d30706;
  wire d30707;
  wire d30708;
  wire d30709;
  wire d3070a;
  wire d3070b;
  wire d3070c;
  wire d3070d;
  wire d3070e;
  wire d3070f;
  wire d30710;
  wire d30711;
  wire d30712;
  wire d30713;
  wire d30714;
  wire d30715;
  wire d30716;
  wire d30717;
  wire d30718;
  wire d30719;
  wire d3071a;
  wire d3071b;
  wire d3071c;
  wire d3071d;
  wire d3071e;
  wire d3071f;
  wire d30720;
  wire d30721;
  wire d30722;
  wire d30723;
  wire d30724;
  wire d30725;
  wire d30726;
  wire d30727;
  wire d30728;
  wire d30729;
  wire d3072a;
  wire d3072b;
  wire d3072c;
  wire d3072d;
  wire d3072e;
  wire d3072f;
  wire d30730;
  wire d30731;
  wire d30732;
  wire d30733;
  wire d30734;
  wire d30735;
  wire d30736;
  wire d30737;
  wire d30738;
  wire d30739;
  wire d3073a;
  wire d3073b;
  wire d3073c;
  wire d3073d;
  wire d3073e;
  wire d3073f;
  wire d30740;
  wire d30741;
  wire d30742;
  wire d30743;
  wire d30744;
  wire d30745;
  wire d30746;
  wire d30747;
  wire d30748;
  wire d30749;
  wire d3074a;
  wire d3074b;
  wire d3074c;
  wire d3074d;
  wire d3074e;
  wire d3074f;
  wire d30750;
  wire d30751;
  wire d30752;
  wire d30753;
  wire d30754;
  wire d30755;
  wire d30756;
  wire d30757;
  wire d30758;
  wire d30759;
  wire d3075a;
  wire d3075b;
  wire d3075c;
  wire d3075d;
  wire d3075e;
  wire d3075f;
  wire d30760;
  wire d30761;
  wire d30762;
  wire d30763;
  wire d30764;
  wire d30765;
  wire d30766;
  wire d30767;
  wire d30768;
  wire d30769;
  wire d3076a;
  wire d3076b;
  wire d3076c;
  wire d3076d;
  wire d3076e;
  wire d3076f;
  wire d30770;
  wire d30771;
  wire d30772;
  wire d30773;
  wire d30774;
  wire d30775;
  wire d30776;
  wire d30777;
  wire d30778;
  wire d30779;
  wire d3077a;
  wire d3077b;
  wire d3077c;
  wire d3077d;
  wire d3077e;
  wire d3077f;
  wire d30780;
  wire d30781;
  wire d30782;
  wire d30783;
  wire d30784;
  wire d30785;
  wire d30786;
  wire d30787;
  wire d30788;
  wire d30789;
  wire d3078a;
  wire d3078b;
  wire d3078c;
  wire d3078d;
  wire d3078e;
  wire d3078f;
  wire d30790;
  wire d30791;
  wire d30792;
  wire d30793;
  wire d30794;
  wire d30795;
  wire d30796;
  wire d30797;
  wire d30798;
  wire d30799;
  wire d3079a;
  wire d3079b;
  wire d3079c;
  wire d3079d;
  wire d3079e;
  wire d3079f;
  wire d307a0;
  wire d307a1;
  wire d307a2;
  wire d307a3;
  wire d307a4;
  wire d307a5;
  wire d307a6;
  wire d307a7;
  wire d307a8;
  wire d307a9;
  wire d307aa;
  wire d307ab;
  wire d307ac;
  wire d307ad;
  wire d307ae;
  wire d307af;
  wire d307b0;
  wire d307b1;
  wire d307b2;
  wire d307b3;
  wire d307b4;
  wire d307b5;
  wire d307b6;
  wire d307b7;
  wire d307b8;
  wire d307b9;
  wire d307ba;
  wire d307bb;
  wire d307bc;
  wire d307bd;
  wire d307be;
  wire d307bf;
  wire d307c0;
  wire d307c1;
  wire d307c2;
  wire d307c3;
  wire d307c4;
  wire d307c5;
  wire d307c6;
  wire d307c7;
  wire d307c8;
  wire d307c9;
  wire d307ca;
  wire d307cb;
  wire d307cc;
  wire d307cd;
  wire d307ce;
  wire d307cf;
  wire d307d0;
  wire d307d1;
  wire d307d2;
  wire d307d3;
  wire d307d4;
  wire d307d5;
  wire d307d6;
  wire d307d7;
  wire d307d8;
  wire d307d9;
  wire d307da;
  wire d307db;
  wire d307dc;
  wire d307dd;
  wire d307de;
  wire d307df;
  wire d307e0;
  wire d307e1;
  wire d307e2;
  wire d307e3;
  wire d307e4;
  wire d307e5;
  wire d307e6;
  wire d307e7;
  wire d307e8;
  wire d307e9;
  wire d307ea;
  wire d307eb;
  wire d307ec;
  wire d307ed;
  wire d307ee;
  wire d307ef;
  wire d307f0;
  wire d307f1;
  wire d307f2;
  wire d307f3;
  wire d307f4;
  wire d307f5;
  wire d307f6;
  wire d307f7;
  wire d307f8;
  wire d307f9;
  wire d307fa;
  wire d307fb;
  wire d307fc;
  wire d307fd;
  wire d307fe;
  wire d307ff;
  wire d30800;
  wire d30801;
  wire d30802;
  wire d30803;
  wire d30804;
  wire d30805;
  wire d30806;
  wire d30807;
  wire d30808;
  wire d30809;
  wire d3080a;
  wire d3080b;
  wire d3080c;
  wire d3080d;
  wire d3080e;
  wire d3080f;
  wire d30810;
  wire d30811;
  wire d30812;
  wire d30813;
  wire d30814;
  wire d30815;
  wire d30816;
  wire d30817;
  wire d30818;
  wire d30819;
  wire d3081a;
  wire d3081b;
  wire d3081c;
  wire d3081d;
  wire d3081e;
  wire d3081f;
  wire d30820;
  wire d30821;
  wire d30822;
  wire d30823;
  wire d30824;
  wire d30825;
  wire d30826;
  wire d30827;
  wire d30828;
  wire d30829;
  wire d3082a;
  wire d3082b;
  wire d3082c;
  wire d3082d;
  wire d3082e;
  wire d3082f;
  wire d30830;
  wire d30831;
  wire d30832;
  wire d30833;
  wire d30834;
  wire d30835;
  wire d30836;
  wire d30837;
  wire d30838;
  wire d30839;
  wire d3083a;
  wire d3083b;
  wire d3083c;
  wire d3083d;
  wire d3083e;
  wire d3083f;
  wire d30840;
  wire d30841;
  wire d30842;
  wire d30843;
  wire d30844;
  wire d30845;
  wire d30846;
  wire d30847;
  wire d30848;
  wire d30849;
  wire d3084a;
  wire d3084b;
  wire d3084c;
  wire d3084d;
  wire d3084e;
  wire d3084f;
  wire d30850;
  wire d30851;
  wire d30852;
  wire d30853;
  wire d30854;
  wire d30855;
  wire d30856;
  wire d30857;
  wire d30858;
  wire d30859;
  wire d3085a;
  wire d3085b;
  wire d3085c;
  wire d3085d;
  wire d3085e;
  wire d3085f;
  wire d30860;
  wire d30861;
  wire d30862;
  wire d30863;
  wire d30864;
  wire d30865;
  wire d30866;
  wire d30867;
  wire d30868;
  wire d30869;
  wire d3086a;
  wire d3086b;
  wire d3086c;
  wire d3086d;
  wire d3086e;
  wire d3086f;
  wire d30870;
  wire d30871;
  wire d30872;
  wire d30873;
  wire d30874;
  wire d30875;
  wire d30876;
  wire d30877;
  wire d30878;
  wire d30879;
  wire d3087a;
  wire d3087b;
  wire d3087c;
  wire d3087d;
  wire d3087e;
  wire d3087f;
  wire d30880;
  wire d30881;
  wire d30882;
  wire d30883;
  wire d30884;
  wire d30885;
  wire d30886;
  wire d30887;
  wire d30888;
  wire d30889;
  wire d3088a;
  wire d3088b;
  wire d3088c;
  wire d3088d;
  wire d3088e;
  wire d3088f;
  wire d30890;
  wire d30891;
  wire d30892;
  wire d30893;
  wire d30894;
  wire d30895;
  wire d30896;
  wire d30897;
  wire d30898;
  wire d30899;
  wire d3089a;
  wire d3089b;
  wire d3089c;
  wire d3089d;
  wire d3089e;
  wire d3089f;
  wire d308a0;
  wire d308a1;
  wire d308a2;
  wire d308a3;
  wire d308a4;
  wire d308a5;
  wire d308a6;
  wire d308a7;
  wire d308a8;
  wire d308a9;
  wire d308aa;
  wire d308ab;
  wire d308ac;
  wire d308ad;
  wire d308ae;
  wire d308af;
  wire d308b0;
  wire d308b1;
  wire d308b2;
  wire d308b3;
  wire d308b4;
  wire d308b5;
  wire d308b6;
  wire d308b7;
  wire d308b8;
  wire d308b9;
  wire d308ba;
  wire d308bb;
  wire d308bc;
  wire d308bd;
  wire d308be;
  wire d308bf;
  wire d308c0;
  wire d308c1;
  wire d308c2;
  wire d308c3;
  wire d308c4;
  wire d308c5;
  wire d308c6;
  wire d308c7;
  wire d308c8;
  wire d308c9;
  wire d308ca;
  wire d308cb;
  wire d308cc;
  wire d308cd;
  wire d308ce;
  wire d308cf;
  wire d308d0;
  wire d308d1;
  wire d308d2;
  wire d308d3;
  wire d308d4;
  wire v845556;
  wire d308d5;
  wire d308d9;
  wire d308da;
  wire d308db;
  wire d308dc;
  wire d308dd;
  wire d308de;
  wire d308df;
  wire d308e0;
  wire d308e1;
  wire d308e2;
  wire d308e3;
  wire d308e4;
  wire d308e5;
  wire d308e6;
  wire d308e7;
  wire d308ea;
  wire d308eb;
  wire d308f3;
  wire d308f4;
  wire d308f5;
  wire d308f6;
  wire d308f7;
  wire d308fa;
  wire d3090c;
  wire d3090d;
  wire d3090e;
  wire d3090f;
  wire d30910;
  wire d30911;
  wire d30912;
  wire d30913;
  wire d30914;
  wire d30915;
  wire d30916;
  wire d30917;
  wire d30918;
  wire d30919;
  wire d3091a;
  wire d3091b;
  wire d3094a;
  wire d3094b;
  wire d3094c;
  wire d3094d;
  wire d3094e;
  wire d3094f;
  wire d30950;
  wire d30951;
  wire d30952;
  wire d30953;
  wire d30954;
  wire d30955;
  wire d30956;
  wire d30957;
  wire d30958;
  wire d30959;
  wire d3095a;
  wire d3095b;
  wire d30188;
  wire d30189;
  wire d3018d;
  wire d3018e;
  wire d3018f;
  wire d30190;
  wire d30191;
  wire d30192;
  wire d30197;
  wire d3019b;
  wire d3019c;
  wire d3019d;
  wire d3019e;
  wire d3019f;
  wire d301a0;
  wire d301a1;
  wire d301a2;
  wire d301a3;
  wire d301a4;
  wire d301a5;
  wire d301a6;
  wire d301a9;
  wire d301aa;
  wire d301ae;
  wire d301af;
  wire d301b0;
  wire d301b1;
  wire d301b6;
  wire d301b7;
  wire d301b8;
  wire d301b9;
  wire d301ba;
  wire d301bb;
  wire d301bc;
  wire d301bd;
  wire d301be;
  wire d301bf;
  wire d301c0;
  wire d301c1;
  wire d301c2;
  wire d301c3;
  wire d301c4;
  wire d301c5;
  wire d301c6;
  wire d301c7;
  wire d301c8;
  wire d301c9;
  wire d301ca;
  wire d301cb;
  wire d301cc;
  wire d301ce;
  wire d301cf;
  wire d301d0;
  wire d301d1;
  wire d301d2;
  wire d301d3;
  wire d301d4;
  wire d301d5;
  wire d301d6;
  wire d301d7;
  wire d301d8;
  wire d301d9;
  wire d301da;
  wire d301db;
  wire d301dc;
  wire d301dd;
  wire d301de;
  wire d301df;
  wire d301e0;
  wire d301e1;
  wire d301e2;
  wire d301e3;
  wire d301e4;
  wire d301e5;
  wire d301e6;
  wire d301e7;
  wire d301e8;
  wire d301e9;
  wire d301ea;
  wire d301eb;
  wire d301ec;
  wire d301ed;
  wire d301ee;
  wire d301ef;
  wire d301f0;
  wire d301f1;
  wire d301f2;
  wire d301f3;
  wire d301f4;
  wire d301f5;
  wire d301f6;
  wire d301f7;
  wire d301f8;
  wire d301f9;
  wire d301fa;
  wire d301fb;
  wire d301fc;
  wire d301fd;
  wire d301fe;
  wire d301ff;
  wire d30200;
  wire d30201;
  wire d30202;
  wire d30203;
  wire d30204;
  wire d30205;
  wire d30206;
  wire d30207;
  wire d30208;
  wire d30209;
  wire d3020a;
  wire d3020b;
  wire d3020c;
  wire d3020d;
  wire d3020e;
  wire d3020f;
  wire d30210;
  wire d30211;
  wire d30212;
  wire d30213;
  wire d30214;
  wire d30215;
  wire d30216;
  wire d30217;
  wire d30218;
  wire d30219;
  wire d3021a;
  wire d3021b;
  wire d3021c;
  wire d3021d;
  wire d30220;
  wire d30221;
  wire d30222;
  wire d30223;
  wire d30224;
  wire d30225;
  wire d30226;
  wire d30227;
  wire d30228;
  wire d30229;
  wire d3022a;
  wire d3022b;
  wire d3022c;
  wire d3022d;
  wire d3022e;
  wire d3022f;
  wire d30230;
  wire d30231;
  wire d30232;
  wire d30233;
  wire d30234;
  wire d30235;
  wire d30236;
  wire d30237;
  wire d30238;
  wire d3023c;
  wire d3023e;
  wire d3023f;
  wire d30240;
  wire d30241;
  wire d30242;
  wire d30243;
  wire d30244;
  wire d30245;
  wire d30246;
  wire d30247;
  wire d30248;
  wire d30249;
  wire d3024a;
  wire d3024b;
  wire d3024c;
  wire d3024d;
  wire d3024e;
  wire d3024f;
  wire d30250;
  wire d30251;
  wire d30252;
  wire d30255;
  wire d30256;
  wire d30257;
  wire d30258;
  wire d30259;
  wire d3025a;
  wire d3025b;
  wire d3025c;
  wire d3025d;
  wire d3025e;
  wire d3025f;
  wire d30263;
  wire d30264;
  wire d30265;
  wire d30266;
  wire d30267;
  wire d30268;
  wire d30269;
  wire d3026a;
  wire d3026b;
  wire d3026c;
  wire d3026d;
  wire d3026e;
  wire d3026f;
  wire d30270;
  wire d30271;
  wire d30272;
  wire d30273;
  wire d30274;
  wire d30275;
  wire d30276;
  wire d30277;
  wire d30278;
  wire d30279;
  wire d3027a;
  wire d3027b;
  wire d3027c;
  wire d3027d;
  wire d3027e;
  wire d3027f;
  wire d30280;
  wire d30281;
  wire d30282;
  wire d30283;
  wire d30284;
  wire d30285;
  wire d30286;
  wire d30287;
  wire d30288;
  wire d30289;
  wire d3028a;
  wire d3028b;
  wire d3028c;
  wire d3028d;
  wire d3028e;
  wire d3028f;
  wire d30290;
  wire d30291;
  wire d30292;
  wire d30293;
  wire d30294;
  wire d30295;
  wire d30296;
  wire d30297;
  wire d30298;
  wire d30299;
  wire d3029a;
  wire d3029b;
  wire d3029c;
  wire d3029d;
  wire d3029e;
  wire d302d2;
  wire d302d3;
  wire d302d4;
  wire d302d5;
  wire d302d6;
  wire d302d7;
  wire d302d8;
  wire d302d9;
  wire d302da;
  wire d302db;
  wire d302dc;
  wire d302dd;
  wire d302de;
  wire d302df;
  wire d302e0;
  wire d302e1;
  wire d302e2;
  wire d302e3;
  wire d302e4;
  wire d302e5;
  wire d302e6;
  wire d302e7;
  wire d302e8;
  wire d302e9;
  wire d302ea;
  wire d302eb;
  wire d302ec;
  wire d302ed;
  wire d302ee;
  wire d302ef;
  wire d302f0;
  wire d302f1;
  wire d302f2;
  wire d302f3;
  wire d302f4;
  wire d302f5;
  wire d302f6;
  wire d302f7;
  wire d302f8;
  wire d302f9;
  wire d2fe7a;
  wire d2fe7b;
  wire d2fe7c;
  wire d2fe7d;
  wire d2fe7e;
  wire d2fe7f;
  wire d2fe80;
  wire d2fe81;
  wire d2fe82;
  wire d2fe83;
  wire d2fe84;
  wire d2fe85;
  wire d2fe86;
  wire d2fe87;
  wire d2fe88;
  wire d2fe89;
  wire d2fe8a;
  wire d2fe8b;
  wire d2fe8c;
  wire d2fe8d;
  wire d2fe8e;
  wire d2fe8f;
  wire d2fe90;
  wire d2fe91;
  wire d2fe92;
  wire d2fe93;
  wire d2fe94;
  wire d2fe95;
  wire d2fe96;
  wire d2fe97;
  wire d2fe98;
  wire d2fe99;
  wire d2fe9a;
  wire d2fe9b;
  wire d2fe9c;
  wire d2fe9d;
  wire d2fe9e;
  wire d2fe9f;
  wire d2fea0;
  wire d2fea1;
  wire d2fea2;
  wire d2fea3;
  wire d2fea4;
  wire d2fea5;
  wire d2fea6;
  wire d2fea7;
  wire d2fea8;
  wire d2fea9;
  wire d2feaa;
  wire d2feab;
  wire d2feac;
  wire d2fead;
  wire d2feae;
  wire d2feb0;
  wire d2feb1;
  wire d2feb2;
  wire d2feb3;
  wire d2feb4;
  wire d2feb5;
  wire d2feb6;
  wire d2feb7;
  wire d2feb8;
  wire d2feb9;
  wire d2feba;
  wire d2febb;
  wire d2febc;
  wire d2febd;
  wire d2febe;
  wire d2febf;
  wire d2fec0;
  wire d2fec1;
  wire d2fec2;
  wire d2fec3;
  wire d2fec4;
  wire d2fec5;
  wire d2fec6;
  wire d2fec7;
  wire d2fec8;
  wire d2fec9;
  wire d2feca;
  wire d2fecb;
  wire d2fecc;
  wire d2fecd;
  wire d2fece;
  wire d2fecf;
  wire d2fed0;
  wire d2fed1;
  wire d2fed2;
  wire d2fed3;
  wire d2fed4;
  wire d2fed5;
  wire d2fed6;
  wire d2fed7;
  wire d2fed8;
  wire d2fed9;
  wire d2feda;
  wire d2fedb;
  wire d2fedc;
  wire d2fedd;
  wire d2fede;
  wire d2fedf;
  wire d2fee0;
  wire d2fee1;
  wire d2fee2;
  wire d2fee3;
  wire d2fee4;
  wire d2fee5;
  wire d2fee6;
  wire d2fee7;
  wire d2fee8;
  wire d2fee9;
  wire d2feea;
  wire d2feeb;
  wire d2feec;
  wire d2feed;
  wire d2feee;
  wire d2feef;
  wire d2fef0;
  wire d2fef1;
  wire d2fef2;
  wire d2fef3;
  wire d2fef4;
  wire d2fef5;
  wire d2fef6;
  wire d2fef7;
  wire d2fef8;
  wire d2fef9;
  wire d2fefa;
  wire d2fefb;
  wire d2fefc;
  wire d2fefd;
  wire d2fefe;
  wire d2feff;
  wire d2ff00;
  wire d2ff01;
  wire d2ff02;
  wire d2ff03;
  wire d2ff04;
  wire d2ff05;
  wire d2ff06;
  wire d2ff07;
  wire d2ff08;
  wire d2ff09;
  wire d2ff0a;
  wire d2ff0b;
  wire d2ff0c;
  wire d2ff0d;
  wire d300b2;
  wire d300b3;
  wire d300b4;
  wire d300b5;
  wire d300b6;
  wire d300b7;
  wire d300b8;
  wire d300b9;
  wire d300ba;
  wire d300bb;
  wire d300bc;
  wire d300bd;
  wire d300be;
  wire d300bf;
  wire d300c0;
  wire d300c1;
  wire d300c2;
  wire d300c3;
  wire d300c4;
  wire d300c5;
  wire d300c6;
  wire d300c7;
  wire d300c8;
  wire d300c9;
  wire d300ca;
  wire d300cb;
  wire d300cc;
  wire d300cd;
  wire d300ce;
  wire d300cf;
  wire d300d0;
  wire d300d1;
  wire d300d2;
  wire d300d3;
  wire d300d4;
  wire d300d5;
  wire d300d6;
  wire d300d7;
  wire d300d8;
  wire d300d9;
  wire d300da;
  wire d300db;
  wire d300dc;
  wire d300dd;
  wire d300de;
  wire d300df;
  wire d300e0;
  wire d300e1;
  wire d300e2;
  wire d300e3;
  wire d300e4;
  wire d300e5;
  wire d300e6;
  wire d300e7;
  wire d300e8;
  wire d300e9;
  wire d300ea;
  wire d300eb;
  wire d300ec;
  wire d300ed;
  wire d300ee;
  wire d300ef;
  wire d300f0;
  wire d300f1;
  wire d300f2;
  wire d300f3;
  wire d300f4;
  wire d300f5;
  wire d300f6;
  wire d300f7;
  wire d300f8;
  wire d300f9;
  wire d300fa;
  wire d300fb;
  wire d300fc;
  wire d300fd;
  wire d300fe;
  wire d300ff;
  wire d30100;
  wire d30101;
  wire d30102;
  wire d30103;
  wire d30104;
  wire d30105;
  wire d30106;
  wire d30107;
  wire d30108;
  wire d30109;
  wire d3010a;
  wire d3010b;
  wire d3010c;
  wire d3010d;
  wire d3010e;
  wire d3010f;
  wire d30110;
  wire d30111;
  wire d30112;
  wire d30113;
  wire d30114;
  wire d30115;
  wire d30116;
  wire d30117;
  wire d30118;
  wire d30119;
  wire d3011a;
  wire d3011b;
  wire d3011c;
  wire d3011d;
  wire d3011e;
  wire d3011f;
  wire d30120;
  wire d30121;
  wire d30122;
  wire d30123;
  wire d30124;
  wire d30125;
  wire d30126;
  wire d30127;
  wire d30128;
  wire d30129;
  wire d3012a;
  wire d3012b;
  wire d3012c;
  wire d3012d;
  wire d3012e;
  wire d3012f;
  wire d30130;
  wire d30131;
  wire d30132;
  wire d30133;
  wire d30134;
  wire d30135;
  wire d30136;
  wire d30137;
  wire d30138;
  wire d30139;
  wire d3013a;
  wire d3013b;
  wire d3013c;
  wire d3013d;
  wire d3013e;
  wire d3013f;
  wire d30140;
  wire d30141;
  wire d30142;
  wire d30143;
  wire d30144;
  wire d30145;
  wire d30146;
  wire d30147;
  wire d30148;
  wire d30149;
  wire d3014a;
  wire d3014b;
  wire d3014c;
  wire d3014d;
  wire d3014e;
  wire d3014f;
  wire d30150;
  wire d30151;
  wire d30152;
  wire d30153;
  wire d30154;
  wire d30155;
  wire d30156;
  wire d30157;
  wire d30158;
  wire d30159;
  wire d3015a;
  wire d3015b;
  wire d3015c;
  wire d3015d;
  wire d3015e;
  wire d3015f;
  wire d30160;
  wire d30161;
  wire d30162;
  wire d30163;
  wire d30164;
  wire d30165;
  wire d30166;
  wire d30167;
  wire d2f96b;
  wire d2f96c;
  wire d2f96d;
  wire d2f96e;
  wire d2f96f;
  wire d2f970;
  wire d2f971;
  wire d2f972;
  wire d2f973;
  wire d2f974;
  wire d2f975;
  wire d2f976;
  wire d2f977;
  wire d2f978;
  wire d2f979;
  wire d2f97a;
  wire d2f97b;
  wire d2f97c;
  wire d2f97d;
  wire d2f97e;
  wire d2f97f;
  wire d2f980;
  wire d2f981;
  wire d2f982;
  wire d2f983;
  wire d2f984;
  wire d2f985;
  wire d2f986;
  wire d2f987;
  wire d2f988;
  wire d2f989;
  wire d2f98a;
  wire d2f98b;
  wire d2f98c;
  wire d2f98d;
  wire d2f98e;
  wire d2f98f;
  wire d2f990;
  wire d2f991;
  wire d2f992;
  wire d2f993;
  wire d2f994;
  wire d2f995;
  wire d2f996;
  wire d2f997;
  wire d2f998;
  wire d2f999;
  wire d2f99a;
  wire d2f99b;
  wire d2f99c;
  wire d2f99d;
  wire d2f99e;
  wire d2f99f;
  wire d2f9a0;
  wire d2f9a1;
  wire d2f9a2;
  wire d2f9a3;
  wire d2f9a4;
  wire d2f9a5;
  wire d2f9a6;
  wire d2f9a7;
  wire d2f9a8;
  wire d2f9a9;
  wire d2f9aa;
  wire d2f9b5;
  wire d2f9b6;
  wire d2f9b7;
  wire d2f9b8;
  wire d2f9b9;
  wire d2f9ba;
  wire d2f9bb;
  wire d2f9bc;
  wire d2f9bd;
  wire d2f9c8;
  wire d2f9c9;
  wire d2f9ca;
  wire d2f9cb;
  wire d2f9cc;
  wire d2f9cd;
  wire d2f9ce;
  wire d2f9cf;
  wire d2f9d0;
  wire d2f9d1;
  wire d2f9d2;
  wire d2f9d3;
  wire d2f9d4;
  wire d2f9d5;
  wire d2f9d6;
  wire d2f9d7;
  wire d2f9d8;
  wire d2f9d9;
  wire d2facd;
  wire d2face;
  wire d2facf;
  wire d2fad0;
  wire d2fad1;
  wire d2fad2;
  wire d2fad3;
  wire d2fad4;
  wire d2fad5;
  wire d2fad6;
  wire d2fad7;
  wire d2fad8;
  wire d2fad9;
  wire d2fada;
  wire d2fadb;
  wire d2fadc;
  wire d2fadd;
  wire d2fade;
  wire d2fadf;
  wire d2fae0;
  wire d2fae1;
  wire d2fae2;
  wire d2fae3;
  wire d2fae4;
  wire d2fae5;
  wire d2fae6;
  wire d2fae7;
  wire d2fae8;
  wire d2fae9;
  wire d2faea;
  wire d2faeb;
  wire d2faec;
  wire d2faed;
  wire d2faee;
  wire d2faef;
  wire d2faf0;
  wire d2faf1;
  wire d2faf2;
  wire d2faf3;
  wire d2faf4;
  wire d2faf5;
  wire d2faf6;
  wire d2faf7;
  wire d2faf8;
  wire d2faf9;
  wire d2fafa;
  wire d2fafb;
  wire d2fafc;
  wire d2fafd;
  wire d2fafe;
  wire d2faff;
  wire d2fb00;
  wire d2fb01;
  wire d2fb02;
  wire d2fb03;
  wire d2fb04;
  wire d2fb05;
  wire d2fb06;
  wire d2fb07;
  wire d2fb08;
  wire d2fb09;
  wire d2fb0a;
  wire d2fb0b;
  wire d2fb0c;
  wire d2fb0d;
  wire d2fb0e;
  wire d2fb0f;
  wire d2fb10;
  wire d2fb11;
  wire d2fb12;
  wire d2fb13;
  wire d2fb14;
  wire d2fb15;
  wire d2fb16;
  wire d2fb17;
  wire d2fb18;
  wire d2fb19;
  wire d2fb1a;
  wire d2fb1b;
  wire d2fb1c;
  wire d2fb1d;
  wire d2fb1e;
  wire d2fb1f;
  wire d2fb20;
  wire d2fb21;
  wire d2fb22;
  wire d2fb23;
  wire d2fb24;
  wire d2fb25;
  wire d2fb26;
  wire d2fb27;
  wire d2fb28;
  wire d2fb29;
  wire d2fb2a;
  wire d2fb2b;
  wire d2fb2c;
  wire d2fb2d;
  wire d2fb2e;
  wire d2fb2f;
  wire d2fb30;
  wire d2fb31;
  wire d2fb32;
  wire d2fb33;
  wire d2fb34;
  wire d2fb35;
  wire d2fb36;
  wire d2fb37;
  wire d2fb38;
  wire d2fb39;
  wire d2fb3a;
  wire d2fb3b;
  wire d2fb3c;
  wire d2fb3d;
  wire d2fb3e;
  wire d2fb3f;
  wire d2fb40;
  wire d2fb41;
  wire d2fb42;
  wire d2fb43;
  wire d2fb44;
  wire d2fb45;
  wire d2fb46;
  wire d2fb47;
  wire d2fb48;
  wire d2fb49;
  wire d2fb4a;
  wire d2fb4b;
  wire d2fb4d;
  wire d2fb4e;
  wire d2fb4f;
  wire d2fb50;
  wire d2fb51;
  wire d2fb52;
  wire d2fb53;
  wire d2fb54;
  wire d2fb55;
  wire d2fb56;
  wire d2fb58;
  wire d2fb59;
  wire d2fb5a;
  wire d2fb5b;
  wire d2fb5c;
  wire d2fb5d;
  wire d2fb5e;
  wire d2fb5f;
  wire d2fb69;
  wire d2fb6a;
  wire d2fb6b;
  wire d2fb6c;
  wire d2fb6d;
  wire d2fb6e;
  wire d2fb6f;
  wire d2fb70;
  wire d2fb71;
  wire d2fb72;
  wire d2fb73;
  wire d2fb74;
  wire d2fb75;
  wire d2fb76;
  wire d2fb77;
  wire d2fb78;
  wire d2fb79;
  wire d2fb7a;
  wire d2fb7b;
  wire d2fb7c;
  wire d2fb7d;
  wire d2fb7e;
  wire d2fb7f;
  wire d2fb80;
  wire d2fb81;
  wire d2fb82;
  wire d2fb83;
  wire d2fb84;
  wire d2fb85;
  wire d2fb86;
  wire d2fb87;
  wire d2fb88;
  wire d2fb89;
  wire d2fb8a;
  wire d2fb8b;
  wire d2fb8c;
  wire d2fb8d;
  wire d2fb8e;
  wire d2fb8f;
  wire d2fb90;
  wire d2fb91;
  wire d2fb92;
  wire d2fb93;
  wire d2fb94;
  wire d2fb95;
  wire d2fb96;
  wire d2fb97;
  wire d2fb98;
  wire d2fb99;
  wire d2fb9a;
  wire d2fb9b;
  wire d2fb9c;
  wire d2fb9d;
  wire d2fb9e;
  wire d2fb9f;
  wire d2fba0;
  wire d2fba1;
  wire d2fba2;
  wire d2fba3;
  wire d2fba4;
  wire d2fba5;
  wire d2fba6;
  wire d2fba7;
  wire d2fba8;
  wire d2fba9;
  wire d2fbaa;
  wire d2fbab;
  wire d2fbac;
  wire d2fbad;
  wire d2fbae;
  wire d2fbaf;
  wire d2fbb0;
  wire d2fbb1;
  wire d2fbb2;
  wire d2fbb3;
  wire d2fbb4;
  wire d2fbb5;
  wire d2fbb6;
  wire d2fbb7;
  wire d2fbb8;
  wire d2fbb9;
  wire d2fbba;
  wire d2fbbb;
  wire d2fbbc;
  wire d2fbbd;
  wire d2fbbe;
  wire d2fbbf;
  wire d2fbc0;
  wire d2fbc1;
  wire d2fbc2;
  wire d2fbc3;
  wire d2fbc4;
  wire d2fbc5;
  wire d2fbc7;
  wire d2fbc8;
  wire d2fbc9;
  wire d2fbca;
  wire d2fbcb;
  wire d2fbcd;
  wire d2fbce;
  wire d2fbcf;
  wire d2fbd0;
  wire d2fbd1;
  wire d2fbd2;
  wire d2fbd3;
  wire d2fbd4;
  wire d2fbd5;
  wire d2fbd6;
  wire d2fbd7;
  wire d2fbd8;
  wire d2fbd9;
  wire d2fbda;
  wire d2fbdb;
  wire d2fbdc;
  wire d2fbdd;
  wire d2fbde;
  wire d2fbdf;
  wire d2fbe0;
  wire d2fbe1;
  wire d2fbe2;
  wire d2fbe3;
  wire d2fbe4;
  wire d2fbe5;
  wire d2fbe6;
  wire d2fbe7;
  wire d2fbe8;
  wire d2fbe9;
  wire d2fbea;
  wire d2fbeb;
  wire d2fbec;
  wire d2fbed;
  wire d2fbee;
  wire d2fbef;
  wire d2fbf0;
  wire d2fbf1;
  wire d2fbf2;
  wire d2fbf3;
  wire d2fbf4;
  wire d2fbf5;
  wire d2fbf6;
  wire d2fbf7;
  wire d2fbf8;
  wire d2fbf9;
  wire d2fbfa;
  wire d2fbfb;
  wire d2fbfc;
  wire d2fbfd;
  wire d2fbfe;
  wire d2fbff;
  wire d2fc00;
  wire d2fc01;
  wire d2fc03;
  wire d2fc04;
  wire d2fc05;
  wire d2fc06;
  wire d2fc07;
  wire d2fc08;
  wire d2fc09;
  wire d2fc0a;
  wire d2fc0b;
  wire d2fc0c;
  wire d2fc0d;
  wire d2fc0e;
  wire d2fc0f;
  wire d2fc10;
  wire d2fc11;
  wire d2fc12;
  wire d2fc13;
  wire d2fc14;
  wire d2fc15;
  wire d2fc16;
  wire d2fc17;
  wire d2fc18;
  wire d2fc19;
  wire d2fc1a;
  wire d2fc21;
  wire d2fc22;
  wire d2fc23;
  wire d2fc24;
  wire d2fc25;
  wire d2fc26;
  wire d2fc27;
  wire d2fc28;
  wire d2fc29;
  wire d2fc2a;
  wire d2fc2b;
  wire d2fc2c;
  wire d2fc2d;
  wire d2fc2e;
  wire d2fc2f;
  wire d2fc30;
  wire d2fc31;
  wire d2fc32;
  wire d2fc33;
  wire d2fc34;
  wire d2fc35;
  wire d2fc36;
  wire d2fc37;
  wire d2fc38;
  wire d2fc39;
  wire d2fc3a;
  wire d2fc3b;
  wire d2fc3c;
  wire d2fc3d;
  wire d2fc3e;
  wire d2fc3f;
  wire d2fc40;
  wire d2fc41;
  wire d2fc42;
  wire d2fc43;
  wire d2fc44;
  wire d2fc45;
  wire d2fc46;
  wire d2fc47;
  wire d2fc48;
  wire d2fc49;
  wire d2fc4a;
  wire d2fc4b;
  wire d2fc4c;
  wire d2fc4d;
  wire d2fc4e;
  wire d2fc4f;
  wire d2fc50;
  wire d2fc51;
  wire d2fc52;
  wire d2fc53;
  wire d2fc54;
  wire d2fc55;
  wire d2fc56;
  wire d2fc57;
  wire d2fc58;
  wire d2fc59;
  wire d2fc5a;
  wire d2fc5b;
  wire d2fc5c;
  wire d2fc5d;
  wire d2fc5e;
  wire d2fc5f;
  wire d2fc60;
  wire d2fc61;
  wire d2fc62;
  wire d2fc63;
  wire d2fc64;
  wire d2fc65;
  wire d2fc66;
  wire d2fc67;
  wire d2fc68;
  wire d2fc69;
  wire d2fc6a;
  wire d2fc6b;
  wire d2fc6c;
  wire d2fc6d;
  wire d2fc6e;
  wire d2fc6f;
  wire d2fc70;
  wire d2fc71;
  wire d2fc72;
  wire d2fc73;
  wire d2fc74;
  wire d2fc75;
  wire d2fc76;
  wire d2fc77;
  wire d2fc78;
  wire d2fc79;
  wire d2fc7a;
  wire d2fc7b;
  wire d2fc7c;
  wire d2fc7f;
  wire d2fc80;
  wire d2fc81;
  wire d2fc82;
  wire d2fc83;
  wire d2fc84;
  wire d2fc85;
  wire d2fc86;
  wire d2fc87;
  wire d2fc88;
  wire d2fc89;
  wire d2fc8a;
  wire d2fc8b;
  wire d2fc8c;
  wire d2fc8d;
  wire v845552;
  wire d2fc8e;
  wire d2fc8f;
  wire d2fcac;
  wire d2fcad;
  wire d2fcae;
  wire d2fcaf;
  wire d2fcb0;
  wire d2fcb1;
  wire d2fcb2;
  wire d2fcb3;
  wire d2fcb4;
  wire d2fcb5;
  wire d2fcb6;
  wire d2fcb7;
  wire d2fcb8;
  wire d2fcd8;
  wire d2fcd9;
  wire d2fce6;
  wire d2fce7;
  wire d2fce8;
  wire d2fce9;
  wire d2fcea;
  wire d2fceb;
  wire d2fcec;
  wire d2fcf3;
  wire d2fcf4;
  wire d2fcfb;
  wire d2fcfc;
  wire d2fcfd;
  wire d2fcfe;
  wire d2fcff;
  wire d2fd00;
  wire d2fd01;
  wire d2fd08;
  wire d2fd09;
  wire d2fd0a;
  wire d2fd0b;
  wire d2fd0c;
  wire d2fd0d;
  wire d2fd0e;
  wire d2fd0f;
  wire d2fd10;
  wire d2fd11;
  wire d2fd12;
  wire d2fd13;
  wire d2fd14;
  wire d2fd15;
  wire d2fd16;
  wire d2fd17;
  wire d2fd18;
  wire d2fd19;
  wire d2fd1a;
  wire d2fd1b;
  wire d2fd1c;
  wire d2fd1d;
  wire d2fd1e;
  wire d2fd1f;
  wire d2fd20;
  wire d2fd21;
  wire d2fd22;
  wire d2fd23;
  wire d2fd24;
  wire d2fd25;
  wire d2fd26;
  wire d2fd27;
  wire d2fd28;
  wire d2fd29;
  wire d2fd2a;
  wire d2fd2b;
  wire d2fd2c;
  wire d2fd2d;
  wire d2fd2e;
  wire d2fd2f;
  wire d2fd30;
  wire d2fd37;
  wire d2fd38;
  wire d2fd39;
  wire d2fd3a;
  wire d2fd3b;
  wire d2fd3c;
  wire d2fd3d;
  wire d2fd3e;
  wire d2fd3f;
  wire d2fd40;
  wire d2fd41;
  wire d2fd42;
  wire d2fd43;
  wire d2fd44;
  wire d2fd45;
  wire d2fd46;
  wire d2fd47;
  wire d2fd48;
  wire d2fd49;
  wire d2fd4a;
  wire d2fd4b;
  wire d2fd4c;
  wire d2fd4d;
  wire d2fd4e;
  wire d2fd4f;
  wire bf1f4d;
  wire bf1f4e;
  wire bf1f4f;
  wire bf1f50;
  wire bf1f51;
  wire bf1f52;
  wire bf1f53;
  wire bf1f54;
  wire bf1f55;
  wire bf1f56;
  wire bf1f57;
  wire bf1f58;
  wire bf1f59;
  wire bf1f5a;
  wire bf1f5b;
  wire bf1f5c;
  wire bf1f5d;
  wire bf1f5e;
  wire bf1f5f;
  wire bf1f60;
  wire bf1f61;
  wire bf1f62;
  wire bf1f63;
  wire bf1f64;
  wire bf1f65;
  wire bf1f66;
  wire bf1f67;
  wire bf1f68;
  wire bf1f69;
  wire bf1f6a;
  wire bf1f6b;
  wire bf1f6c;
  wire bf1f6d;
  wire bf1f6e;
  wire bf1f6f;
  wire bf1f70;
  wire bf1f71;
  wire bf1f72;
  wire bf1f73;
  wire bf1f74;
  wire bf1f75;
  wire bf1f76;
  wire bf1f77;
  wire bf1f78;
  wire bf1f79;
  wire bf1f7a;
  wire bf1f7b;
  wire bf1f7c;
  wire bf1f7d;
  wire bf1f7e;
  wire bf1f7f;
  wire bf1f80;
  wire bf1f81;
  wire bf1f82;
  wire bf1f83;
  wire bf1f84;
  wire bf1f85;
  wire bf1f86;
  wire bf1f87;
  wire bf1f88;
  wire bf1f89;
  wire bf1f8a;
  wire bf1f8b;
  wire bf1f8c;
  wire bf1f8d;
  wire bf1f8e;
  wire bf1f8f;
  wire bf1f90;
  wire bf1f91;
  wire bf1f92;
  wire bf1f93;
  wire bf1f94;
  wire bf1f95;
  wire bf1f96;
  wire bf1f97;
  wire bf1f98;
  wire bf1f99;
  wire bf1f9a;
  wire bf1f9b;
  wire bf1f9c;
  wire bf1f9d;
  wire bf1f9e;
  wire bf1f9f;
  wire bf1fa0;
  wire bf1fa1;
  wire bf1fa2;
  wire bf1fa3;
  wire bf1fa4;
  wire bf1fa5;
  wire bf1fa6;
  wire bf1fa7;
  wire bf1fa8;
  wire bf1fa9;
  wire bf1faa;
  wire bf1fab;
  wire v845555;
  wire v16a2664;
  wire v16a2665;
  wire v16a2666;
  wire v16a2667;
  wire v16a2668;
  wire v16a2669;
  wire v16a266a;
  wire v84554d;
  wire v16a266b;
  wire v845559;
  wire v16a266f;
  wire v16a2670;
  wire v16a2671;
  wire v16a2672;
  wire v16a2673;
  wire v16a2674;
  wire v16a2675;
  wire v16a2676;
  wire v16a2677;
  wire v16a2678;
  wire v16a2679;
  wire v16a267a;
  wire v16a267b;
  wire v16a1f93;
  wire v16a1f94;
  wire v16a1f95;
  wire v16a1f96;
  wire v16a1f97;
  wire v16a1f98;
  wire v16a1f99;
  wire v16a1f9a;
  wire v16a1f9b;
  wire v16a1f9c;
  wire v16a1f9d;
  wire v16a1f9e;
  wire v16a2058;
  wire v16a2059;
  wire v16a205a;
  wire v9109e4;
  wire v16a205b;
  wire v16a205c;
  wire v16a205d;
  wire v16a205e;
  wire v16a205f;
  wire v16a2060;
  wire v16a2061;
  wire v16a2062;
  wire v16a2063;
  wire v16a2064;
  wire v16a2065;
  wire v16a2066;
  wire v16a2067;
  wire v845582;
  wire v16a2068;
  wire v16a2069;
  wire v16a206a;
  wire v16a206b;
  wire v16a206c;
  wire v16a206d;
  wire v16a206e;
  wire v16a206f;
  wire v16a2070;
  wire v16a2071;
  wire v16a2072;
  wire v16a2073;
  wire v16a2074;
  wire v16a2075;
  wire v16a2076;
  wire v16a2077;
  wire v16a2078;
  wire v16a2079;
  wire v16a207a;
  wire v16a207b;
  wire v16a207c;
  wire v16a207d;
  wire v16a207e;
  wire v16a207f;
  wire v16a2080;
  wire v16a2081;
  wire v16a2082;
  wire v16a2083;
  wire v16a2084;
  wire v16a2085;
  wire v16a2086;
  wire v16a2087;
  wire v16a2088;
  wire v16a2089;
  wire v16a208a;
  wire v16a208b;
  wire v16a208c;
  wire v16a208d;
  wire v16a208e;
  wire v16a208f;
  wire v16a2090;
  wire v16a2091;
  wire v16a2092;
  wire v16a2093;
  wire v16a2094;
  wire v16a2095;
  wire v16a2096;
  wire v16a2097;
  wire v16a2098;
  wire v16a2099;
  wire v16a209a;
  wire v16a209b;
  wire v16a209c;
  wire v16a209d;
  wire v16a209e;
  wire v16a209f;
  wire v16a20a0;
  wire v16a20a1;
  wire v16a20a2;
  wire v16a20a3;
  wire v16a20a4;
  wire v16a20a5;
  wire v16a20a6;
  wire v845547;
  wire v16a2234;
  wire v16a2235;
  wire v16a2236;
  wire v16a2237;
  wire v16a2238;
  wire v16a2239;
  wire v16a223a;
  wire v16a223b;
  wire v16a223c;
  wire v16a223d;
  wire v16a223e;
  wire v16a223f;
  wire v16a2240;
  wire v16a2241;
  wire v16a2242;
  wire v16a2243;
  wire v16a2244;
  wire v16a2245;
  wire v16a2246;
  wire v16a2247;
  wire v16a2248;
  wire v16a2249;
  wire v16a224a;
  wire v16a224b;
  wire v16a224c;
  wire v16a224d;
  wire v16a224e;
  wire v16a224f;
  wire v16a1ab7;
  wire v16a1ab8;
  wire v16a1ab9;
  wire v16a1aba;
  wire v16a1abb;
  wire v16a1abc;
  wire v16a1abd;
  wire v16a1abe;
  wire v16a1abf;
  wire v16a1ac0;
  wire v16a1ac1;
  wire v16a1ac2;
  wire v16a1ac3;
  wire v16a1ac4;
  wire v16a1ac5;
  wire v16a1ac6;
  wire v16a1ac7;
  wire v16a1ac8;
  wire v16a1ac9;
  wire v16a1aca;
  wire v16a1acb;
  wire v16a1acc;
  wire v16a1acd;
  wire v16a1ace;
  wire v16a1acf;
  wire v16a1ad0;
  wire v16a1ad1;
  wire v16a1ad2;
  wire v16a1ad3;
  wire v16a1ad4;
  wire v16a1ad5;
  wire v16a1ad6;
  wire v16a1ad7;
  wire v16a1ad8;
  wire v16a1ad9;
  wire v16a1ada;
  wire v16a1adb;
  wire v16a1adc;
  wire v16a1add;
  wire v16a1ade;
  wire v16a1adf;
  wire v16a1ae0;
  wire v16a1ae1;
  wire v16a1ae2;
  wire v16a1ae3;
  wire v16a1ae4;
  wire v16a1ae5;
  wire v16a1ae6;
  wire v16a1ae7;
  wire v16a1ae8;
  wire v16a1ae9;
  wire v16a1aea;
  wire v16a1aeb;
  wire v16a1aec;
  wire v16a1aed;
  wire v16a1aee;
  wire v16a1aef;
  wire v16a1af0;
  wire v16a1af1;
  wire v16a1af2;
  wire v16a1af3;
  wire v16a1af4;
  wire v16a1af5;
  wire v16a1af6;
  wire v16a1af7;
  wire v16a1af8;
  wire v16a1af9;
  wire v16a1afa;
  wire v16a1afb;
  wire v16a1afc;
  wire v16a1afd;
  wire v16a1afe;
  wire v16a1aff;
  wire v16a1b00;
  wire v16a1b01;
  wire v16a1b02;
  wire v16a1b03;
  wire v16a1b62;
  wire v16a1b63;
  wire v16a1b64;
  wire v16a1b65;
  wire v16a1b66;
  wire v16a1b67;
  wire v16a1b68;
  wire v16a1b69;
  wire v16a1b6a;
  wire v16a1b6b;
  wire v16a1bb2;
  wire v16a1bb3;
  wire v16a1bb4;
  wire v16a1bb5;
  wire v16a1bb6;
  wire v16a1bb7;
  wire v16a1bb8;
  wire v16a1bb9;
  wire v16a1bba;
  wire v16a1bbb;
  wire v16a1bbc;
  wire v16a1bbd;
  wire v16a1bbe;
  wire v16a1bbf;
  wire v16a1bc0;
  wire v16a1bc1;
  wire v16a1bc2;
  wire v16a1bc3;
  wire v16a1bc4;
  wire v16a1bc5;
  wire v16a1bc6;
  wire v16a1bc7;
  wire v16a1bc8;
  wire v16a1bc9;
  wire v16a1bca;
  wire v16a1bcb;
  wire v16a1bcc;
  wire v16a1bcd;
  wire v16a1bce;
  wire v16a1bcf;
  wire v16a1bd0;
  wire v16a1bd1;
  wire v16a1bd2;
  wire v16a1bd3;
  wire v16a1bd4;
  wire v16a1bd5;
  wire v16a1bd6;
  wire v16a1bd7;
  wire v16a1bd8;
  wire v16a1bd9;
  wire v16a1bda;
  wire v16a1bdb;
  wire v16a1bdc;
  wire v16a1bdd;
  wire v16a1bde;
  wire v16a1bdf;
  wire v16a1be0;
  wire v16a1be1;
  wire v16a1be2;
  wire v16a1be3;
  wire v16a1be4;
  wire v16a1be5;
  wire v16a1be6;
  wire v16a1be7;
  wire v16a1be8;
  wire v16a1be9;
  wire v16a1bea;
  wire v16a1beb;
  wire v16a1bec;
  wire v16a1bed;
  wire v16a1bee;
  wire v16a1bef;
  wire v16a1bf0;
  wire v16a1bf1;
  wire v16a1bf2;
  wire v16a1bf3;
  wire v16a1bf4;
  wire v16a1bf5;
  wire v16a1bf6;
  wire v16a1bf7;
  wire v16a1bf8;
  wire v16a1bf9;
  wire v16a1bfa;
  wire v16a1bfb;
  wire v16a1bfc;
  wire v16a1bfd;
  wire v16a1bfe;
  wire v16a1bff;
  wire v16a1c00;
  wire v16a1c01;
  wire v16a1c02;
  wire v16a1c03;
  wire v16a1c04;
  wire v16a1c05;
  wire v16a1c95;
  wire v16a1c96;
  wire v16a1c97;
  wire v16a1c98;
  wire v16a1c99;
  wire v16a1c9a;
  wire v16a1c9b;
  wire v16a1c9c;
  wire v16a1c9d;
  wire v16a1c9e;
  wire v16a1c9f;
  wire v16a1ca0;
  wire v16a1ca1;
  wire v16a1ca2;
  wire v16a1ca3;
  wire v16a1ca4;
  wire v16a1ca5;
  wire v16a1ca6;
  wire v16a1ca7;
  wire v16a1ca8;
  wire v16a1cb9;
  wire v16a1cba;
  wire v16a1cbb;
  wire v16a1cbc;
  wire v16a1cbd;
  wire v16a1cbe;
  wire v16a1cbf;
  wire v16a1cc0;
  wire v16a1cc1;
  wire v16a1cc2;
  wire v16a1cc3;
  wire v16a1cc4;
  wire v16a1cc5;
  wire v16a1cc6;
  wire v16a1cc7;
  wire v16a1cc8;
  wire v16a1cc9;
  wire v16a1cca;
  wire v16a1ccb;
  wire v16a1ccc;
  wire v16a1ccd;
  wire v16a1cce;
  wire v16a1ccf;
  wire v16a1cd0;
  wire v16a1cd1;
  wire v16a1cd2;
  wire v16a1cd3;
  wire v16a1cd4;
  wire v16a1cd5;
  wire v16a1cd6;
  wire v16a1cd7;
  wire v16a1cd8;
  wire v16a1cd9;
  wire v16a1cda;
  wire v16a1cdb;
  wire v16a1cdc;
  wire v16a1cdd;
  wire v16a1cde;
  wire v16a1cdf;
  wire v16a1ce0;
  wire v16a1ce1;
  wire v16a1ce2;
  wire v16a1ce3;
  wire v16a1ce4;
  wire v16a1ce5;
  wire v16a1ce6;
  wire v16a1ce7;
  wire v16a1ce8;
  wire v16a1ce9;
  wire v16a1cea;
  wire v16a1ceb;
  wire v16a1cec;
  wire v16a1ced;
  wire v16a1cee;
  wire v16a1cef;
  wire v16a1cf0;
  wire v16a1cf1;
  wire v16a1cf2;
  wire v16a1cf3;
  wire v16a1cf4;
  wire v16a1cf5;
  wire v16a1cf6;
  wire v16a1cf7;
  wire v16a1cf8;
  wire v16a1cf9;
  wire v16a1cfa;
  wire v16a1cfb;
  wire v16a1cfc;
  wire v16a1cfd;
  wire v16a1cfe;
  wire v16a1cff;
  wire v16a1d00;
  wire v16a1d01;
  wire v16a1d02;
  wire v16a1d03;
  wire v16a1d04;
  wire v16a1d05;
  wire v16a1d0e;
  wire v16a1d0f;
  wire v16a1d10;
  wire v16a1d11;
  wire v16a1d12;
  wire v16a1d16;
  wire v16a1d17;
  wire v16a1d18;
  wire v16a1d19;
  wire v16a1d1a;
  wire v16a1d1b;
  wire v16a1d1e;
  wire v16a1d1f;
  wire v16a1d20;
  wire v16a1d21;
  wire v16a1d25;
  wire v16a1d26;
  wire v16a1d27;
  wire v16a1d28;
  wire v16a1d29;
  wire v16a1d2a;
  wire v16a1d2b;
  wire v16a1d2c;
  wire v16a1d2d;
  wire v16a1d2e;
  wire v16a1d2f;
  wire v16a1d30;
  wire v16a1d31;
  wire v16a1d32;
  wire v16a1d33;
  wire v16a1d34;
  wire v16a1d35;
  wire v16a1d36;
  wire v16a1d37;
  wire v16a1d39;
  wire v16a1d3a;
  wire v16a1d3b;
  wire v16a1d3c;
  wire v16a1d3d;
  wire v16a1d3e;
  wire v16a1d3f;
  wire v16a1d40;
  wire v16a1d41;
  wire v16a1d42;
  wire v16a1d43;
  wire v16a1d44;
  wire v16a1d45;
  wire v16a1d46;
  wire v16a1d47;
  wire v16a1d48;
  wire v16a1d49;
  wire v16a1d4a;
  wire v16a1d4b;
  wire v16a1d4c;
  wire v16a1d4d;
  wire v16a1d50;
  wire v16a1d51;
  wire v16a1d53;
  wire v16a1d54;
  wire v16a1d55;
  wire v16a1d56;
  wire v16a1d57;
  wire v16a1d58;
  wire v16a1d59;
  wire v16a1d5a;
  wire v16a1d5b;
  wire v16a1d5c;
  wire v16a1d5d;
  wire v16a1d5e;
  wire v16a1d5f;
  wire v16a1d60;
  wire v16a1d61;
  wire v16a1d62;
  wire v16a1d63;
  wire v16a1d64;
  wire v16a1d65;
  wire v16a1d66;
  wire v16a1d67;
  wire v16a1d68;
  wire v16a1d6a;
  wire v16a1d6b;
  wire v16a1d6c;
  wire v16a1d6d;
  wire v16a1d6e;
  wire v16a1d6f;
  wire v16a1d70;
  wire v16a1d73;
  wire v16a1d74;
  wire v16a1d76;
  wire v16a1d77;
  wire v16a1d78;
  wire v16a1d79;
  wire v16a1d7a;
  wire v16a1d7b;
  wire v16a1d7c;
  wire v16a1d7d;
  wire v16a1d7e;
  wire v16a1d7f;
  wire v16a1d80;
  wire v16a1d81;
  wire v16a1d82;
  wire v16a1d8c;
  wire v16a1d8d;
  wire v16a1d8e;
  wire v16a1d91;
  wire v16a1d92;
  wire v16a1d93;
  wire v16a1d94;
  wire v16a1d95;
  wire v16a1d97;
  wire v16a1d98;
  wire v16a1d99;
  wire v16a1d9a;
  wire v16a1d9b;
  wire v16a1d9c;
  wire v16a1d9d;
  wire v16a1d9e;
  wire v16a1d9f;
  wire v16a1da0;
  wire v16a1da1;
  wire v16a1da2;
  wire v16a1da3;
  wire v16a1da4;
  wire v16a1da5;
  wire v16a1da6;
  wire v16a1da7;
  wire v16a1da8;
  wire v16a1da9;
  wire v16a1daa;
  wire v16a1dab;
  wire v16a1dac;
  wire v16a1dad;
  wire v16a1dae;
  wire v16a1daf;
  wire v16a1db0;
  wire v16a1db1;
  wire v16a1db2;
  wire v16a1db3;
  wire v16a1db4;
  wire v16a1db5;
  wire v16a1db6;
  wire v16a1db7;
  wire v16a1db8;
  wire v16a1db9;
  wire v16a1dba;
  wire v16a1dbb;
  wire v16a1dbc;
  wire v16a1dbd;
  wire v16a1dbe;
  wire v16a1dbf;
  wire v16a1dc0;
  wire v16a1dc1;
  wire v16a1dd2;
  wire v16a1dd3;
  wire v16a1dd4;
  wire v16a1dd5;
  wire v16a1dd6;
  wire v16a1dd7;
  wire v16a1dd8;
  wire v16a1dd9;
  wire v16a1dda;
  wire v16a1deb;
  wire v16a1dec;
  wire v16a1ded;
  wire v16a1dfd;
  wire v16a1dfe;
  wire v16a1dff;
  wire v16a1e00;
  wire v16a1e01;
  wire v16a1e02;
  wire v16a1e03;
  wire v16a1e04;
  wire v16a1e05;
  wire v16a1e06;
  wire v16a1e07;
  wire v16a1e08;
  wire v16a1e09;
  wire v16a1e0a;
  wire v16a1e0b;
  wire v16a1e0c;
  wire v16a1e0d;
  wire v16a1e0e;
  wire v16a1e1f;
  wire v16a1e20;
  wire v16a1e21;
  wire v16a1e22;
  wire v16a1e23;
  wire v16a1e24;
  wire v16a1e25;
  wire v16a1e26;
  wire v16a1e27;
  wire v16a1e28;
  wire v16a1e29;
  wire v16a1e2a;
  wire v16a1e2b;
  wire v16a1e2c;
  wire v16a1e2d;
  wire v16a1e2e;
  wire v16a1e2f;
  wire v16a1e30;
  wire v16a1e49;
  wire v16a1e4a;
  wire v16a1e4b;
  wire v16a1e4c;
  wire v16a1e4d;
  wire v16a1e4e;
  wire v16a1e4f;
  wire v16a1e50;
  wire v16a1e51;
  wire v16a1e52;
  wire v16a1e53;
  wire v16a1e54;
  wire v16a1e55;
  wire v16a1e56;
  wire v16a1e57;
  wire v16a1e58;
  wire v16a1e59;
  wire v16a1e5a;
  wire v16a1e5b;
  wire v16a1e5c;
  wire v16a1e5d;
  wire v16a1e5e;
  wire v16a1e5f;
  wire v16a1e60;
  wire v16a1e61;
  wire v16a1e62;
  wire v16a1e63;
  wire v16a1e64;
  wire v16a1e65;
  wire v16a1e66;
  wire v16a1e67;
  wire v16a1e68;
  wire v16a1e69;
  wire v16a1e6a;
  wire v16a1e6b;
  wire v16a1e6c;
  wire v16a1e6d;
  wire v16a1e6e;
  wire v16a1e6f;
  wire v16a1e70;
  wire v16a1e71;
  wire v16a1e72;
  wire v16a1e73;
  wire v16a1e74;
  wire v16a1e75;
  wire v16a1e76;
  wire v16a1e77;
  wire v16a1e78;
  wire v16a1e79;
  wire v16a1e7a;
  wire v16a1e89;
  wire v16a1e8a;
  wire v16a1e8b;
  wire v16a1e8c;
  wire v16a1e8d;
  wire v16a1e8e;
  wire v16a1e8f;
  wire v16a1e90;
  wire v16a1e91;
  wire v16a1e92;
  wire v16a1e93;
  wire v16a1e94;
  wire v16a1e95;
  wire v16a1e96;
  wire v16a1e97;
  wire v16a1e98;
  wire v16a169c;
  wire v16a169d;
  wire v16a169e;
  wire v16a169f;
  wire v16a16a0;
  wire v16a16a1;
  wire v16a16a2;
  wire v16a16a3;
  wire v16a16a4;
  wire v16a16a5;
  wire v16a16a6;
  wire v16a16a7;
  wire v16a16a8;
  wire v16a16a9;
  wire v16a16aa;
  wire v16a16ab;
  wire v16a16ac;
  wire v16a16ad;
  wire v16a16ae;
  wire v16a16af;
  wire v16a16b0;
  wire v16a16b1;
  wire v16a16b2;
  wire v16a16b3;
  wire v16a16b4;
  wire v16a16b5;
  wire v16a16b6;
  wire v16a16b7;
  wire v16a183f;
  wire v16a1840;
  wire v16a1841;
  wire v16a1842;
  wire v16a1843;
  wire v16a1844;
  wire v16a1845;
  wire v16a1846;
  wire v16a1847;
  wire v16a1848;
  wire v16a1887;
  wire v16a1888;
  wire v16a1889;
  wire v16a188a;
  wire v16a188b;
  wire v16a188c;
  wire v16a188d;
  wire v16a188e;
  wire v16a188f;
  wire v16a1890;
  wire v16a18dd;
  wire v16a18de;
  wire v16a193d;
  wire v16a193e;
  wire v16a193f;
  wire v16a1940;
  wire v16a1941;
  wire v16a1942;
  wire v16a1943;
  wire v16a1944;
  wire v16a1945;
  wire v16a1946;
  wire v16a1947;
  wire v16a1948;
  wire v16a1949;
  wire v16a194a;
  wire v16a194b;
  wire v16a194c;
  wire v16a194d;
  wire v16a194e;
  wire v16a194f;
  wire v16a1950;
  wire v16a1951;
  wire v16a1952;
  wire v16a1953;
  wire v16a1954;
  wire v16a1955;
  wire v16a1956;
  wire v16a1957;
  wire v16a1958;
  wire v16a1959;
  wire v16a195a;
  wire v16a195b;
  wire v16a195c;
  wire v16a195d;
  wire v16a195e;
  wire v16a195f;
  wire v16a1960;
  wire v16a1961;
  wire v16a1962;
  wire v16a1963;
  wire v16a1964;
  wire v16a1965;
  wire v16a1966;
  wire v16a1967;
  wire v16a1968;
  wire v16a1969;
  wire v16a196a;
  wire v16a196b;
  wire v16a196c;
  wire v16a196d;
  wire v16a196e;
  wire v16a196f;
  wire v16a1970;
  wire v16a1971;
  wire v16a1972;
  wire v16a1973;
  wire v16a1974;
  wire v16a1975;
  wire v16a1976;
  wire v16a1977;
  wire v16a1978;
  wire v16a1979;
  wire v16a197a;
  wire v16a197b;
  wire v16a197c;
  wire v16a197d;
  wire v16a197e;
  wire v16a197f;
  wire v16a1980;
  wire v16a1981;
  wire v16a1982;
  wire v16a1983;
  wire v16a1984;
  wire v16a1985;
  wire v16a19a4;
  wire v16a19a5;
  wire v16a19a6;
  wire v16a19a7;
  wire v16a19a8;
  wire v16a19a9;
  wire v16a19aa;
  wire v16a19ab;
  wire v16a19ac;
  wire v16a19ad;
  wire v16a19ae;
  wire v16a19af;
  wire v16a19b0;
  wire v16a19b1;
  wire v16a19b2;
  wire v16a19b3;
  wire v16a19b4;
  wire v16a19b5;
  wire v16a19b6;
  wire v16a19b7;
  wire v16a19b8;
  wire v16a19b9;
  wire v16a19bf;
  wire v16a19c0;
  wire v16a19c1;
  wire v16a19c2;
  wire v16a19c3;
  wire v16a19c4;
  wire v16a19c5;
  wire v16a19c6;
  wire v16a19c7;
  wire v16a19c8;
  wire v16a19c9;
  wire v16a19ca;
  wire v16a19cb;
  wire v16a19cc;
  wire v16a19cd;
  wire v16a19ce;
  wire v16a19cf;
  wire v16a19d0;
  wire v16a19d1;
  wire v16a19d2;
  wire v16a19d3;
  wire v16a19d4;
  wire v16a19dd;
  wire v16a19de;
  wire v16a19df;
  wire v16a19e0;
  wire v16a19e1;
  wire v16a19e2;
  wire v16a19e3;
  wire v16a19e4;
  wire v16a19e5;
  wire v16a19e6;
  wire v16a1a20;
  wire v16a1a21;
  wire v16a1a22;
  wire v16a1a23;
  wire v16a1a24;
  wire v16a1a25;
  wire v16a1a26;
  wire v16a1a27;
  wire v16a1a28;
  wire v16a1a29;
  wire v16a1a2a;
  wire v16a1a2b;
  wire v16a1a2c;
  wire v16a1a2d;
  wire v16a1a2e;
  wire v16a1a2f;
  wire v16a1a30;
  wire v16a1a31;
  wire v16a1a75;
  wire v16a1a76;
  wire v16a1a77;
  wire v16a1a78;
  wire v16a1a79;
  wire v16a1a7a;
  wire v16a1a7b;
  wire v16a1a7c;
  wire v16a1a7d;
  wire v16a1a7e;
  wire v16a1a7f;
  wire v16a1a80;
  wire v16a1a81;
  wire v16a1a82;
  wire v16a1a83;
  wire v16a1a84;
  wire v16a1a85;
  wire v16a1a86;
  wire v16a1a87;
  wire v16a1a88;
  wire v16a1a89;
  wire v16a1a8a;
  wire v16a1a8b;
  wire v16a1a8c;
  wire v16a1a8d;
  wire v16a1a8e;
  wire v16a1a8f;
  wire v16a1a90;
  wire v16a1a91;
  wire v16a1a92;
  wire v16a1a93;
  wire v16a1a94;
  wire v16a1a95;
  wire v16a1a96;
  wire v16a1a97;
  wire v16a1a98;
  wire v16a1a99;
  wire v16a129c;
  wire v16a129d;
  wire v16a129e;
  wire v16a129f;
  wire v16a12be;
  wire v16a12bf;
  wire v16a12c0;
  wire v16a12c1;
  wire v16a12c2;
  wire v16a12c3;
  wire v16a12c4;
  wire v16a12c5;
  wire v16a12c6;
  wire v16a12c7;
  wire v16a12e4;
  wire v16a12e5;
  wire v16a12e6;
  wire v16a12e7;
  wire v16a12e8;
  wire v16a12e9;
  wire v16a12ea;
  wire v16a12eb;
  wire v16a12ec;
  wire v16a12ed;
  wire v16a12ee;
  wire v16a12ef;
  wire v16a12f0;
  wire v16a12f1;
  wire v16a12f2;
  wire v16a12f3;
  wire v16a12f4;
  wire v16a12f5;
  wire v16a12f6;
  wire v16a12f7;
  wire v16a12f8;
  wire v16a12f9;
  wire v16a131b;
  wire v16a131c;
  wire v16a131d;
  wire v16a131e;
  wire v16a131f;
  wire v16a1320;
  wire v16a1321;
  wire v16a1322;
  wire v16a1323;
  wire v16a1324;
  wire v16a1325;
  wire v16a1326;
  wire v16a1327;
  wire v16a1328;
  wire v16a1329;
  wire v16a132a;
  wire v16a132b;
  wire v16a132c;
  wire v16a132d;
  wire v16a132e;
  wire v16a132f;
  wire v16a1330;
  wire v16a1331;
  wire v16a1332;
  wire v16a1333;
  wire v16a1334;
  wire v16a1335;
  wire v16a1336;
  wire v16a1337;
  wire v16a1372;
  wire v16a1373;
  wire v16a1374;
  wire v16a1375;
  wire v16a1376;
  wire v16a1377;
  wire v16a1378;
  wire v16a1379;
  wire v16a137a;
  wire v16a137b;
  wire v16a137c;
  wire v16a137d;
  wire v16a137e;
  wire v16a137f;
  wire v16a1380;
  wire v16a1381;
  wire v16a1382;
  wire v16a1383;
  wire v16a1384;
  wire v16a1385;
  wire v16a1386;
  wire v16a1387;
  wire v16a1388;
  wire v16a1389;
  wire v16a138a;
  wire v16a138b;
  wire v16a138c;
  wire v16a138d;
  wire v16a138e;
  wire v16a138f;
  wire v16a1390;
  wire v16a1391;
  wire v16a1392;
  wire v16a1393;
  wire v16a1394;
  wire v16a1395;
  wire v16a1396;
  wire v16a1397;
  wire v16a1398;
  wire v16a1399;
  wire v16a139a;
  wire v16a139b;
  wire v16a139c;
  wire v16a139d;
  wire v16a139e;
  wire v16a139f;
  wire v16a13a7;
  wire v16a13a8;
  wire v16a13ba;
  wire v16a13c0;
  wire v16a13c1;
  wire v16a13c2;
  wire v16a13c3;
  wire v16a13c4;
  wire v16a13c5;
  wire v16a13c6;
  wire v16a13c7;
  wire v16a13c8;
  wire v16a13c9;
  wire v16a13ca;
  wire v16a13cb;
  wire v16a13cc;
  wire v16a13cd;
  wire v16a13ce;
  wire v16a13cf;
  wire v16a13d0;
  wire v16a13d1;
  wire v16a13d2;
  wire v16a13d3;
  wire v16a13d4;
  wire v16a13d5;
  wire v16a13d6;
  wire v16a13d7;
  wire v16a13d8;
  wire v16a13d9;
  wire v16a13da;
  wire v16a13db;
  wire v16a13dc;
  wire v16a13dd;
  wire v16a13de;
  wire v16a13df;
  wire v16a13e0;
  wire v16a13e1;
  wire v16a13e2;
  wire v16a13e3;
  wire v16a13e4;
  wire v16a13e5;
  wire v16a13e6;
  wire v16a13e7;
  wire v16a13e8;
  wire v16a13e9;
  wire v16a13ea;
  wire v16a13eb;
  wire v16a13ec;
  wire v16a13ed;
  wire v16a13ee;
  wire v16a13ef;
  wire v16a13f0;
  wire v16a13f1;
  wire v16a13f2;
  wire v16a13f3;
  wire v16a13f4;
  wire v16a13f5;
  wire v16a13f6;
  wire v16a13f7;
  wire v16a13f8;
  wire v16a13f9;
  wire v16a13fa;
  wire v16a13fb;
  wire v16a13fc;
  wire v16a13fd;
  wire v16a13fe;
  wire v16a13ff;
  wire v16a1400;
  wire v16a1401;
  wire v16a1402;
  wire v16a1403;
  wire v16a1404;
  wire v16a1405;
  wire v16a1406;
  wire v16a1407;
  wire v16a1408;
  wire v16a1409;
  wire v16a140a;
  wire v16a140b;
  wire v16a140c;
  wire v16a140d;
  wire v16a140e;
  wire v16a140f;
  wire v16a1410;
  wire v16a1411;
  wire v16a1412;
  wire v16a1413;
  wire v16a1414;
  wire v16a1415;
  wire v16a1416;
  wire v16a1417;
  wire v16a1418;
  wire v16a1419;
  wire v16a141a;
  wire v16a141b;
  wire v16a141c;
  wire v16a141d;
  wire v16a141e;
  wire v16a141f;
  wire v16a1420;
  wire v16a1421;
  wire v16a1422;
  wire v16a1423;
  wire v16a1424;
  wire v16a1425;
  wire v16a1426;
  wire v16a1427;
  wire v16a1428;
  wire v16a1429;
  wire v16a142a;
  wire v16a142b;
  wire v16a142c;
  wire v16a142d;
  wire v16a142e;
  wire v16a142f;
  wire v16a1430;
  wire v16a1431;
  wire v16a1432;
  wire v16a1433;
  wire v16a1434;
  wire v16a1435;
  wire v16a1436;
  wire v16a1437;
  wire v16a1438;
  wire v16a1439;
  wire v16a143a;
  wire v16a143b;
  wire v16a143c;
  wire v16a143d;
  wire v16a143e;
  wire v16a143f;
  wire v16a1440;
  wire v16a1441;
  wire v16a1442;
  wire v16a1443;
  wire v16a1444;
  wire v16a1445;
  wire v16a1446;
  wire v16a1447;
  wire v16a1448;
  wire v16a1449;
  wire v16a144a;
  wire v16a144b;
  wire v15167b6;
  wire v15167b7;
  wire v15167b8;
  wire v15167b9;
  wire v15167bd;
  wire v15167be;
  wire v15167bf;
  wire v15167c0;
  wire v15167c1;
  wire v15167c2;
  wire v15167c3;
  wire v15167c4;
  wire v15167e8;
  wire v15167e9;
  wire v15167ea;
  wire v15167eb;
  wire v9745f6;
  wire v15167ec;
  wire v15167ed;
  wire v15167ee;
  wire v15167ef;
  wire v15167f0;
  wire v15167f1;
  wire v15167f2;
  wire v15167f3;
  wire v15167f4;
  wire v15167f5;
  wire v15167f6;
  wire v15167f7;
  wire v15167f8;
  wire v15167f9;
  wire v15167fa;
  wire v15167fb;
  wire v15167fc;
  wire v15167fd;
  wire v15167fe;
  wire v15167ff;
  wire v1516800;
  wire v1516801;
  wire v1516802;
  wire v1516803;
  wire v1516804;
  wire v1516805;
  wire v1516806;
  wire v1516853;
  wire v1516854;
  wire v1516855;
  wire v15168a5;
  wire v15168a6;
  wire v15168a7;
  wire v15168a8;
  wire v15168a9;
  wire v15168aa;
  wire v15168ab;
  wire v15168ac;
  wire v15168ad;
  wire v15168ae;
  wire v15168af;
  wire v15168b0;
  wire v15168b1;
  wire v15168b2;
  wire v15168b3;
  wire v15168b4;
  wire v15168b5;
  wire v15168b6;
  wire v15168b7;
  wire v15168b8;
  wire v15168eb;
  wire v15168ec;
  wire v15168ed;
  wire v15168ee;
  wire v15168ef;
  wire v15168f0;
  wire v15168f1;
  wire v15168f2;
  wire v15168f3;
  wire v15168f4;
  wire v15168f5;
  wire v15168f6;
  wire v15168f7;
  wire v15168f8;
  wire v15168f9;
  wire v15168fa;
  wire v15168fb;
  wire v15168fc;
  wire v15168fd;
  wire v15168fe;
  wire v15168ff;
  wire v1516900;
  wire v1516957;
  wire v1516958;
  wire v1516959;
  wire v1516975;
  wire v1516979;
  wire v151697a;
  wire v151697b;
  wire v151697c;
  wire v151697d;
  wire v151697e;
  wire v151697f;
  wire v1516980;
  wire v1516981;
  wire v1516982;
  wire v1516988;
  wire v1516998;
  wire v1516999;
  wire v151699a;
  wire v151699b;
  wire v151699c;
  wire v151699d;
  wire v151699e;
  wire v151699f;
  wire v15169a0;
  wire v15161cb;
  wire v15161cc;
  wire v15161cd;
  wire v15161ce;
  wire v15161cf;
  wire v15161d0;
  wire v15161d1;
  wire v15161d2;
  wire v15161d3;
  wire v15161d4;
  wire v15161d5;
  wire v15161d6;
  wire v15161d7;
  wire v15161f9;
  wire v15161fa;
  wire v15161fb;
  wire v15161fc;
  wire v15161fd;
  wire v15161fe;
  wire v15161ff;
  wire v1516200;
  wire v1516201;
  wire v1516213;
  wire v1516214;
  wire v1516215;
  wire v1516216;
  wire v1516217;
  wire v1516218;
  wire v1516219;
  wire v151621a;
  wire v151621b;
  wire v151621c;
  wire v151621d;
  wire v151621e;
  wire v15160f9;
  wire v15160fa;
  wire v15160fb;
  wire v15160fc;
  wire v15160fd;
  wire v15160fe;
  wire v15160ff;
  wire v1516100;
  wire v1516101;
  wire v1516102;
  wire v1516103;
  wire v1516104;
  wire v1516105;
  wire v1516106;
  wire v1516107;
  wire v1515adf;
  wire v1515ae0;
  wire v1515ae1;
  wire v1515ae2;
  wire v1515ae3;
  wire v1515ae4;
  wire v1515ae5;
  wire v1515ae6;
  wire v1515ae7;
  wire v1515ae8;
  wire v1515ae9;
  wire v1515aea;
  wire v1515aeb;
  wire v1515aec;
  wire v1515aed;
  wire v1515aee;
  wire v1515aef;
  wire v1515bae;
  wire v1515baf;
  wire v1515bb0;
  wire v1515c7b;
  wire v1515c7c;
  wire v1515c7d;
  wire v1515c7e;
  wire v1515c7f;
  wire v1515c80;
  wire v1515c81;
  wire v1515c82;
  wire v1515c83;
  wire v1515c84;
  wire v1515c85;
  wire v1515c86;
  wire v1515c87;
  wire v1515c88;
  wire v15155e4;
  wire v15155e5;
  wire v15155e6;
  wire v15155e7;
  wire v15155e8;
  wire v15155e9;
  wire v15155ea;
  wire v15155eb;
  wire v15155ec;
  wire v15155ed;
  wire v15155ee;
  wire v15155ef;
  wire v15155f0;
  wire v15155f1;
  wire v15155f2;
  wire v15155f3;
  wire v15155f4;
  wire v15155f5;
  wire v15155f6;
  wire v15155f7;
  wire v15155f8;
  wire v15155f9;
  wire v15155fa;
  wire v15155fb;
  wire v15155fc;
  wire v15155fd;
  wire v15155fe;
  wire v15155ff;
  wire v1515600;
  wire v1515601;
  wire v1515602;
  wire v1515603;
  wire v1515604;
  wire v1515605;
  wire v1515606;
  wire v1515607;
  wire v1515608;
  wire v1515609;
  wire v151560a;
  wire v151560b;
  wire v151560c;
  wire v151560d;
  wire v151560e;
  wire v151560f;
  wire v1515610;
  wire v1515611;
  wire v1515612;
  wire v1515613;
  wire v1515614;
  wire v1515615;
  wire v1515616;
  wire v1515617;
  wire v1515618;
  wire v1515619;
  wire v151561a;
  wire v151561b;
  wire v151561c;
  wire v151561d;
  wire v151561e;
  wire v151561f;
  wire v1515620;
  wire v1515621;
  wire v1515622;
  wire v1515623;
  wire v1515624;
  wire v1515625;
  wire v1515626;
  wire v1515627;
  wire v1515628;
  wire v1515629;
  wire v151562a;
  wire v151562b;
  wire v151562c;
  wire v151562d;
  wire v151562e;
  wire v151562f;
  wire v1515630;
  wire v1515631;
  wire v1515632;
  wire v1515633;
  wire v1515634;
  wire v1515635;
  wire v1515636;
  wire v1515637;
  wire v1515638;
  wire v1515639;
  wire v151563a;
  wire v151563b;
  wire v151563c;
  wire v151563d;
  wire v151563e;
  wire v151563f;
  wire v1515640;
  wire v1515641;
  wire v1515642;
  wire v1515643;
  wire v1515644;
  wire v1515645;
  wire v1515646;
  wire v1515647;
  wire v1515648;
  wire v1515649;
  wire v151564a;
  wire v151564b;
  wire v151564c;
  wire v151564d;
  wire v151564e;
  wire v151564f;
  wire v1515650;
  wire v1515651;
  wire v1515652;
  wire v1515653;
  wire v1515654;
  wire v1515655;
  wire v1515656;
  wire v1515657;
  wire v1515658;
  wire v1515659;
  wire v151565a;
  wire v151565b;
  wire v1515667;
  wire v1515668;
  wire v1515669;
  wire v151566a;
  wire v151566b;
  wire v151566c;
  wire v151566d;
  wire v151566e;
  wire v151566f;
  wire v1515670;
  wire v1515671;
  wire v1515672;
  wire v1515673;
  wire v1515674;
  wire v1515675;
  wire v151567e;
  wire v151567f;
  wire v15156ad;
  wire v15156ae;
  wire v15156af;
  wire v15156b0;
  wire v15156b1;
  wire v15156b2;
  wire v15156b3;
  wire v15156b4;
  wire v15156b5;
  wire v15156b6;
  wire v15156b7;
  wire v15156b8;
  wire v15156b9;
  wire v15156ba;
  wire v15156bb;
  wire v15156bc;
  wire v15156bd;
  wire v15156be;
  wire v15156c6;
  wire v15156c7;
  wire v15156c8;
  wire v15156c9;
  wire v15156ca;
  wire v15156cb;
  wire v15156cc;
  wire v15156cd;
  wire v15156ce;
  wire v15156d5;
  wire v15156d6;
  wire v15156d7;
  wire v15156d8;
  wire v15156d9;
  wire v15156da;
  wire v15156db;
  wire v15156e3;
  wire v15156e4;
  wire v15156e5;
  wire v15156e6;
  wire v15156e7;
  wire v15156e8;
  wire v15156e9;
  wire v15156ea;
  wire v15156eb;
  wire v15156ec;
  wire v15156ed;
  wire v15156ee;
  wire v15156ef;
  wire v15156f0;
  wire v15156f1;
  wire v15156f2;
  wire v15156f3;
  wire v15156f4;
  wire v15156f5;
  wire v15156f6;
  wire v15156f7;
  wire v15156f8;
  wire v15156f9;
  wire v15156fa;
  wire v15156fb;
  wire v15156fc;
  wire v15156fd;
  wire v15156fe;
  wire v15156ff;
  wire v1515700;
  wire v1515701;
  wire v1515702;
  wire v1515703;
  wire v1515704;
  wire v1515705;
  wire v1515706;
  wire v1515707;
  wire v1515708;
  wire v1515709;
  wire v151570a;
  wire v151570b;
  wire v151570c;
  wire v151570d;
  wire v151570e;
  wire v151570f;
  wire v1515710;
  wire v1515711;
  wire v1515712;
  wire v1515713;
  wire v1515714;
  wire v1515715;
  wire v1515716;
  wire v1515717;
  wire v1515718;
  wire v1515719;
  wire v151571a;
  wire v151571b;
  wire v151571c;
  wire v151571d;
  wire v151571e;
  wire v151571f;
  wire v1515720;
  wire v1515721;
  wire v1515722;
  wire v1515723;
  wire v1515724;
  wire v1515725;
  wire v1515726;
  wire v1515727;
  wire v1515728;
  wire v1515729;
  wire v151572a;
  wire v151572b;
  wire v151572c;
  wire v151572d;
  wire v151572e;
  wire v151572f;
  wire v1515730;
  wire v1515731;
  wire v1515732;
  wire v1515733;
  wire v1515734;
  wire v1515735;
  wire v1515736;
  wire v1515737;
  wire v1515738;
  wire v1515739;
  wire v151573a;
  wire v151573b;
  wire v151573c;
  wire v151573d;
  wire v151573e;
  wire v151573f;
  wire v1515740;
  wire v1515741;
  wire v1515742;
  wire v1515743;
  wire v1515744;
  wire v1515745;
  wire v1515746;
  wire v1515747;
  wire v1515748;
  wire v1515749;
  wire v151574a;
  wire v151574b;
  wire v151574c;
  wire v151574d;
  wire v151574e;
  wire v151574f;
  wire v1515750;
  wire v1515751;
  wire v1515752;
  wire v1515753;
  wire v1515754;
  wire v1515755;
  wire v1515756;
  wire v1515757;
  wire v1515758;
  wire v1515759;
  wire v151575a;
  wire v151575b;
  wire v151575c;
  wire v151575d;
  wire v151575e;
  wire v151575f;
  wire v1515760;
  wire v1515761;
  wire v1515762;
  wire v1515763;
  wire v1515764;
  wire v1515765;
  wire v1515766;
  wire v1515767;
  wire v1515768;
  wire v1515769;
  wire v151576a;
  wire v151576b;
  wire v151576c;
  wire v151576d;
  wire v151576e;
  wire v151576f;
  wire v1515770;
  wire v1515771;
  wire v1515772;
  wire v1515773;
  wire v1515774;
  wire v1515775;
  wire v1515776;
  wire v1515777;
  wire v1515778;
  wire v1515779;
  wire v151577a;
  wire v151577b;
  wire v151577c;
  wire v151577d;
  wire v151577e;
  wire v151577f;
  wire v1515780;
  wire v1515781;
  wire v1515782;
  wire v1515783;
  wire v1515784;
  wire v1515785;
  wire v1515786;
  wire v1515787;
  wire v1515788;
  wire v1515789;
  wire v151578a;
  wire v151578b;
  wire v151578c;
  wire v151578d;
  wire v151578e;
  wire v151578f;
  wire v1515790;
  wire v1515791;
  wire v1515792;
  wire v1515793;
  wire v1515794;
  wire v1515795;
  wire v1515796;
  wire v1515797;
  wire v1515798;
  wire v1515799;
  wire v151579a;
  wire v151579b;
  wire v151579c;
  wire v151579d;
  wire v151579e;
  wire v151579f;
  wire v15157a0;
  wire v15157a1;
  wire v15157a2;
  wire v15157a3;
  wire v15157a4;
  wire v15157a5;
  wire v15157a6;
  wire v15157a7;
  wire v15157a8;
  wire v15157a9;
  wire v15157aa;
  wire v15157ab;
  wire v15157ac;
  wire v15157ad;
  wire v15157ae;
  wire v15157af;
  wire v15157b0;
  wire v15157b1;
  wire v15157b2;
  wire v15157b3;
  wire v15157b4;
  wire v15157b5;
  wire v15157b6;
  wire v15157b7;
  wire v15157b8;
  wire v15157b9;
  wire v15157ba;
  wire v15157bb;
  wire v15157bc;
  wire v15157bd;
  wire v15157be;
  wire v15157bf;
  wire v15157c0;
  wire v15157c1;
  wire v15157c2;
  wire v15157c3;
  wire v15157c4;
  wire v15157c5;
  wire v15157c6;
  wire v15157c7;
  wire v15157c8;
  wire v15157c9;
  wire v15157ca;
  wire v15157cb;
  wire v15157cc;
  wire v15157cd;
  wire v15157ce;
  wire v15157cf;
  wire v15157d0;
  wire v15157d1;
  wire v15157d2;
  wire v15157d3;
  wire v15157d4;
  wire v15157d5;
  wire v15157d6;
  wire v15157d7;
  wire v15157d8;
  wire v15157d9;
  wire v15157da;
  wire v15157db;
  wire v15157dc;
  wire v15157dd;
  wire v15157de;
  wire v15157df;
  wire v15157e0;
  wire v15157e1;
  wire v15157e2;
  wire v15157e3;
  wire v15157e4;
  wire v15157e5;
  wire v15157e6;
  wire v15157e7;
  wire v15157e8;
  wire v15157e9;
  wire v15157ea;
  wire v15157eb;
  wire v15157ec;
  wire v15157ed;
  wire v15157ee;
  wire v15157ef;
  wire v15157f0;
  wire v15157f1;
  wire v15157f2;
  wire v15157f3;
  wire v15157f4;
  wire v15157f5;
  wire v15157f6;
  wire v15157f7;
  wire v15157f8;
  wire v15157f9;
  wire v15157fa;
  wire v15157fb;
  wire v15157fc;
  wire v15157fd;
  wire v15157fe;
  wire v15157ff;
  wire v1515800;
  wire v1515801;
  wire v1515802;
  wire v1515803;
  wire v1515804;
  wire v1515805;
  wire v1515806;
  wire v1515807;
  wire v1515808;
  wire v1515809;
  wire v151580a;
  wire v151580b;
  wire v151580c;
  wire v151580d;
  wire v151580e;
  wire v151580f;
  wire v1515810;
  wire v1515811;
  wire v1515812;
  wire v1515813;
  wire v1515814;
  wire v1515815;
  wire v1515816;
  wire v1515817;
  wire v1515818;
  wire v1515819;
  wire v151581a;
  wire v151581b;
  wire v151581c;
  wire v151581d;
  wire v151581e;
  wire v151581f;
  wire v1515820;
  wire v1515821;
  wire v1515822;
  wire v1515823;
  wire v1515824;
  wire v1515825;
  wire v1515826;
  wire v1515827;
  wire v1515828;
  wire v1515829;
  wire v151582a;
  wire v151582b;
  wire v151582c;
  wire v151582d;
  wire v151582e;
  wire v151582f;
  wire v1515830;
  wire v1515831;
  wire v1515832;
  wire v1515833;
  wire v1515834;
  wire v1515835;
  wire v1515836;
  wire v1515837;
  wire v1515838;
  wire v1515839;
  wire v151583a;
  wire v151583b;
  wire v151583c;
  wire v151583d;
  wire v151583e;
  wire v151583f;
  wire v1515840;
  wire v1515841;
  wire v1515842;
  wire v1515843;
  wire v1515844;
  wire v1515845;
  wire v1515846;
  wire v1515847;
  wire v1515848;
  wire v1515849;
  wire v151584a;
  wire v151584b;
  wire v151584c;
  wire v151584d;
  wire v151584e;
  wire v151584f;
  wire v1515850;
  wire v1515851;
  wire v1515852;
  wire v1515853;
  wire v1515854;
  wire v1515855;
  wire v1515856;
  wire v1515857;
  wire v845578;
  wire v14eb679;
  wire v845566;
  wire v143fd77;
  wire v143fd78;
  wire v143fd79;
  wire v143fd7a;
  wire v143fd7b;
  wire v143fd7c;
  wire v143fd7d;
  wire v14838b7;
  wire v14838b8;
  wire v14838b9;
  wire v14838ba;
  wire v14838bb;
  wire v14838bc;
  wire v14838bd;
  wire v14838be;
  wire v14838bf;
  wire v134d1d9;
  wire v134d1da;
  wire v134d1db;
  wire v134d1dc;
  wire v134d1dd;
  wire v134d1de;
  wire v134d1df;
  wire v134d1e0;
  wire v134d1e1;
  wire v134d1e2;
  wire v134d1e3;
  wire v134d1e4;
  wire v134d1e5;
  wire v134d1e6;
  wire v134d1e7;
  wire v134d1e8;
  wire v134d1e9;
  wire v134d1ea;
  wire v134d1eb;
  wire v134d1ec;
  wire v134d1ed;
  wire v134d1ee;
  wire v134d1ef;
  wire v134d1f0;
  wire v134d1f1;
  wire v134d1f2;
  wire v134d1f3;
  wire v134d1f4;
  wire v134d1f5;
  wire v134d1f6;
  wire v134d1f7;
  wire v134d1f8;
  wire v134d1f9;
  wire v134d1fa;
  wire v134d1fb;
  wire v134d1fc;
  wire v134d1fd;
  wire v134d1fe;
  wire v134d1ff;
  wire v134d200;
  wire v134d201;
  wire v134d202;
  wire v134d203;
  wire v134d204;
  wire v134d205;
  wire v134d206;
  wire v134d207;
  wire v134d208;
  wire v134d209;
  wire v134d20a;
  wire v134d20b;
  wire v134d20c;
  wire v134d20d;
  wire v134d20e;
  wire v134d20f;
  wire v134d210;
  wire v134d211;
  wire v134d212;
  wire v134d213;
  wire v134d214;
  wire v134d215;
  wire v134d216;
  wire v134d217;
  wire v134d218;
  wire v134d219;
  wire v134d21a;
  wire v134d21b;
  wire v134d21c;
  wire v134d21d;
  wire v134d21e;
  wire v134d21f;
  wire v134d220;
  wire v134d221;
  wire v134d222;
  wire v134d223;
  wire v134d224;
  wire v134d225;
  wire v134d226;
  wire v134d227;
  wire v134d228;
  wire v134d229;
  wire v134d22a;
  wire v134d22b;
  wire v134d22c;
  wire v134d22d;
  wire v134d22e;
  wire v134d22f;
  wire v134d230;
  wire v134d231;
  wire v134d232;
  wire v134d233;
  wire v134d234;
  wire v134d235;
  wire v134d236;
  wire v134d237;
  wire v134d238;
  wire v134d239;
  wire v134d23a;
  wire v134d23b;
  wire v134d23c;
  wire v134d23d;
  wire v134d23e;
  wire v134d23f;
  wire v134d240;
  wire v134d241;
  wire v134d242;
  wire v134d243;
  wire v134d244;
  wire v134d245;
  wire v134d260;
  wire v134d261;
  wire v134d262;
  wire v134d263;
  wire v134d264;
  wire v134d265;
  wire v134d266;
  wire v134d267;
  wire v134d268;
  wire v134d269;
  wire v134d26a;
  wire v134d26b;
  wire v134d26c;
  wire v134d26d;
  wire v134d26e;
  wire v134d26f;
  wire v134d270;
  wire v134d271;
  wire v134d272;
  wire v134d273;
  wire v134d274;
  wire v134d275;
  wire v134d276;
  wire v134d277;
  wire v134d278;
  wire v134d279;
  wire v134d27a;
  wire v134d27b;
  wire v134d27c;
  wire v134d27d;
  wire v134d27e;
  wire v134d27f;
  wire v134d280;
  wire v134d281;
  wire v134d282;
  wire v134d283;
  wire v134d284;
  wire v134d285;
  wire v134d286;
  wire v134d287;
  wire v134d288;
  wire v134d289;
  wire v134d28a;
  wire v134d28b;
  wire v134d28c;
  wire v134d28d;
  wire v134d28e;
  wire v134d28f;
  wire v134d290;
  wire v134d291;
  wire v134d292;
  wire v134d293;
  wire v134d294;
  wire v134d295;
  wire v134d296;
  wire v134d308;
  wire v134d309;
  wire v134d30a;
  wire v134d30b;
  wire v134d30c;
  wire v134d30d;
  wire v134d30e;
  wire v134d30f;
  wire v134d310;
  wire v134d311;
  wire v134d312;
  wire v134d313;
  wire v134d314;
  wire v134d315;
  wire v134d316;
  wire v134d34f;
  wire v134d363;
  wire v134d364;
  wire v134d365;
  wire v134d366;
  wire v134d367;
  wire v134d368;
  wire v134d369;
  wire v134d36a;
  wire v134d36b;
  wire v134d36c;
  wire v134d36d;
  wire v134d36e;
  wire v134d36f;
  wire v134d370;
  wire v134d371;
  wire v134d372;
  wire v134d373;
  wire v134d374;
  wire v134d375;
  wire v134d376;
  wire v134d377;
  wire v134d378;
  wire v134d379;
  wire v134d37a;
  wire v134d37b;
  wire v134d37c;
  wire v134d37d;
  wire v134d37e;
  wire v134d37f;
  wire v134d380;
  wire v134d381;
  wire v134d382;
  wire v134d383;
  wire v134d384;
  wire v134d385;
  wire v134d386;
  wire v134d387;
  wire v134d388;
  wire v134d389;
  wire v134d38a;
  wire v134d38b;
  wire v134d38c;
  wire v134d38d;
  wire v134d38e;
  wire v134d38f;
  wire v134d390;
  wire v134d391;
  wire v134d392;
  wire v134d393;
  wire v134d394;
  wire v134d395;
  wire v134d396;
  wire v134d397;
  wire v134d398;
  wire v134d399;
  wire v134d39a;
  wire v134d39b;
  wire v134d39c;
  wire v134d3a9;
  wire v134d3aa;
  wire v134d3ab;
  wire v134d3ac;
  wire v134d3ad;
  wire v134d3ae;
  wire v134d3af;
  wire v134d3b0;
  wire v134d3b1;
  wire v134d3b2;
  wire v134d3b3;
  wire v134d3b4;
  wire v134d3b5;
  wire v134d3b6;
  wire v134d3b7;
  wire v134d3b8;
  wire v134d3b9;
  wire v134d3ba;
  wire v134d3bb;
  wire v134d3bc;
  wire v134d3bd;
  wire v134d3be;
  wire v134d3bf;
  wire v134d3c0;
  wire v134d3c1;
  wire v134d3c2;
  wire v134d3c3;
  wire v134d3c4;
  wire v134d3c5;
  wire v134d3c6;
  wire v134d3c7;
  wire v134d3c8;
  wire v134d3c9;
  wire v134d3ca;
  wire v134d3cb;
  wire v134d3cc;
  wire v134d3cd;
  wire v134d3ce;
  wire v134d3cf;
  wire v134d3d0;
  wire v134d3d1;
  wire v134d3d2;
  wire v134d3d3;
  wire v134d3d4;
  wire v134d3d5;
  wire v134d3d6;
  wire v134d3d7;
  wire v134d3d8;
  wire v134d3d9;
  wire v134d3da;
  wire v134d3db;
  wire v134d3dc;
  wire v134d3dd;
  wire v134d3de;
  wire v134d3df;
  wire v134d3e0;
  wire v134d3e1;
  wire v134d3e2;
  wire v134d3e3;
  wire v134d3e4;
  wire v134d3e5;
  wire v134d3e6;
  wire v134d3e7;
  wire v134d3e8;
  wire v134d3e9;
  wire v134d3fa;
  wire v134d3fb;
  wire v134d3fc;
  wire v134d425;
  wire v134d426;
  wire v134d427;
  wire v134d428;
  wire v134d429;
  wire v134d42a;
  wire v134d42b;
  wire v134d42c;
  wire v134d42d;
  wire v134d42e;
  wire v134d42f;
  wire v134d430;
  wire v134d431;
  wire v134d432;
  wire v134d433;
  wire v134d434;
  wire v134d43c;
  wire v134d43d;
  wire v134d43e;
  wire v134d43f;
  wire v134d440;
  wire v134d441;
  wire v134d442;
  wire v134d443;
  wire v134d444;
  wire v134d445;
  wire v134d446;
  wire v134d447;
  wire v134d448;
  wire v134d449;
  wire v134d44a;
  wire v134d44b;
  wire v134d44c;
  wire v134d44d;
  wire v134d44e;
  wire v134d44f;
  wire v134d450;
  wire v134d451;
  wire v134d452;
  wire v134d453;
  wire v134d454;
  wire v134d455;
  wire v134d456;
  wire v134d457;
  wire v134d458;
  wire v134d459;
  wire v134d45a;
  wire v134d45b;
  wire v134d45c;
  wire v134d45d;
  wire v134d45e;
  wire v134d45f;
  wire v134d460;
  wire v134d461;
  wire v134d462;
  wire v134d463;
  wire v134d464;
  wire v134d465;
  wire v134d466;
  wire v134d467;
  wire v134d468;
  wire v134d469;
  wire v134d46a;
  wire v134d46b;
  wire v134d46c;
  wire v134d46d;
  wire v134d495;
  wire v134d496;
  wire v134d497;
  wire v134d498;
  wire v134d499;
  wire v134d49a;
  wire v134d49b;
  wire v134d49c;
  wire v134d49f;
  wire v134d4a0;
  wire v134d4a1;
  wire v134d4a2;
  wire v134d4a3;
  wire v134d4a4;
  wire v134d4a5;
  wire v134d4a6;
  wire v134d4a7;
  wire v134d4a8;
  wire v134d4a9;
  wire v134d4aa;
  wire v134d4ab;
  wire v134d4ac;
  wire v134d4ad;
  wire v134d4ae;
  wire v134d4af;
  wire v134d4b0;
  wire v134d4b1;
  wire v134d4b2;
  wire v134d4b3;
  wire v134d4b4;
  wire v134d4b5;
  wire v134d4b6;
  wire v134d4b7;
  wire v134d4b8;
  wire v134d4b9;
  wire v134d4ba;
  wire v134d4bb;
  wire v134d4bc;
  wire v134d4c2;
  wire v134d4c3;
  wire v134d4c4;
  wire v134d4c5;
  wire v134d4c6;
  wire v134d4c7;
  wire v134d4c8;
  wire v134d4c9;
  wire v134d4ca;
  wire v134d4cb;
  wire v134d4cc;
  wire v134d4cd;
  wire v134d4ce;
  wire v134d4cf;
  wire v134d4d0;
  wire v134d4d1;
  wire v134d4d2;
  wire v134d4d3;
  wire v134d4d4;
  wire v134d4d5;
  wire v134d4d6;
  wire v134d4d7;
  wire v134d4d8;
  wire v134d4d9;
  wire v134d4da;
  wire v134d4db;
  wire v134d4dc;
  wire v134d4dd;
  wire v134d4de;
  wire v134d4df;
  wire v134d4e0;
  wire v134d4e1;
  wire v134d4e2;
  wire v134d4e3;
  wire v134d4e4;
  wire v134d4e5;
  wire v134d4e6;
  wire v134d4e7;
  wire v134d4e8;
  wire v134d4e9;
  wire v134d4ea;
  wire v134d4eb;
  wire v134d4ec;
  wire v134d4ed;
  wire v134d4ee;
  wire v134d4ef;
  wire v134d4f0;
  wire v134d4f1;
  wire v134d4f2;
  wire v134d4f3;
  wire v134d4f4;
  wire v134d4f5;
  wire v134d4f6;
  wire v134d4f7;
  wire v134d4f8;
  wire v134d4f9;
  wire v134d4fa;
  wire v134d4fb;
  wire v134d4fc;
  wire v134d4fd;
  wire v134d4fe;
  wire v134d4ff;
  wire v134d500;
  wire v134d501;
  wire v134d502;
  wire v134d503;
  wire v134d504;
  wire v134d505;
  wire v134d506;
  wire v134d507;
  wire v134d508;
  wire v134d509;
  wire v134d50a;
  wire v134d50b;
  wire v134d50c;
  wire v134d50d;
  wire v134d50e;
  wire v134d50f;
  wire v134d510;
  wire v134d511;
  wire v134d512;
  wire v134d513;
  wire v134d514;
  wire v134d515;
  wire v134d516;
  wire v134d517;
  wire v134d518;
  wire v134d519;
  wire v134d51a;
  wire v134d51b;
  wire v134d51c;
  wire v134d51d;
  wire v134d51e;
  wire v134d51f;
  wire v134d520;
  wire v134d521;
  wire v134d522;
  wire v134d523;
  wire v134d524;
  wire v134d525;
  wire v134d526;
  wire v134d527;
  wire v134d528;
  wire v134d529;
  wire v134d52a;
  wire v134d52b;
  wire v134d52c;
  wire v134d52d;
  wire v134d52e;
  wire v134d52f;
  wire v134d530;
  wire v134d531;
  wire v134d532;
  wire v134d533;
  wire v134d534;
  wire v134d535;
  wire v134d536;
  wire v134d537;
  wire v134d538;
  wire v134d539;
  wire v134d53a;
  wire v134d53b;
  wire v134d53c;
  wire v134d53d;
  wire v134d53e;
  wire v134d53f;
  wire v134d540;
  wire v134d541;
  wire v134cd44;
  wire v134cd45;
  wire v134cd55;
  wire v134cd56;
  wire v134cd57;
  wire v134cd58;
  wire v134cd59;
  wire v134cd5a;
  wire v134cd5b;
  wire v134cd5c;
  wire v134cd5d;
  wire v134cd5e;
  wire v134cd5f;
  wire v134cd60;
  wire v134cd61;
  wire v134cd62;
  wire v134cd63;
  wire v134cd64;
  wire v134cd65;
  wire v134cd66;
  wire v134cd67;
  wire v134cd68;
  wire v134cd69;
  wire v134cd6a;
  wire v134cd6b;
  wire v134cd6c;
  wire v134cd6d;
  wire v134cd6e;
  wire v134cd6f;
  wire v134cd70;
  wire v134cd71;
  wire v134cd72;
  wire v134cd73;
  wire v134cd74;
  wire v134cd75;
  wire v134cd76;
  wire v134cd77;
  wire v134cd78;
  wire v134cd79;
  wire v134cd7a;
  wire v134cd7b;
  wire v134cd7c;
  wire v134cd7d;
  wire v134cd7e;
  wire v134cd7f;
  wire v134cd80;
  wire v134cd81;
  wire v134cd82;
  wire v134cd83;
  wire v134cd84;
  wire v134cd85;
  wire v134cd86;
  wire v134cd87;
  wire v134cd88;
  wire v134cd89;
  wire v134cd8a;
  wire v134cd8b;
  wire v134cd8c;
  wire v134cd8d;
  wire v134cd8e;
  wire v134cd8f;
  wire v134cdc2;
  wire v134cdc3;
  wire v134cdc4;
  wire v134cdc5;
  wire v134cdc6;
  wire v134cdc7;
  wire v134cdc8;
  wire v134cdc9;
  wire v134cdca;
  wire v134cdcb;
  wire v134cdcc;
  wire v134cdcd;
  wire v134cdce;
  wire v134cdcf;
  wire v134ce33;
  wire v134ce34;
  wire v134ce35;
  wire v134ce36;
  wire v134ce37;
  wire v134ce38;
  wire v134ce39;
  wire v134ce3a;
  wire v134ce3b;
  wire v134ce3c;
  wire v134ce3d;
  wire v134ce3e;
  wire v134ce3f;
  wire v134ce40;
  wire v134ce41;
  wire v134ce42;
  wire v134ce43;
  wire v134ce44;
  wire v134ce45;
  wire v134ce46;
  wire v134ce47;
  wire v134ce48;
  wire v134ce52;
  wire v134ce53;
  wire v134ce54;
  wire v134ce55;
  wire v134ce56;
  wire v134ce57;
  wire v134ce58;
  wire v134ce59;
  wire v134ce5a;
  wire v134ce5b;
  wire v134ce5c;
  wire v134ce5d;
  wire v134ce5e;
  wire v134ce5f;
  wire v134ce60;
  wire v134ce61;
  wire v134ce62;
  wire v134ce63;
  wire v134ce64;
  wire v134ce65;
  wire v134ce66;
  wire v134ce67;
  wire v134ce68;
  wire v134ce69;
  wire v134ce6a;
  wire v134ce6b;
  wire v134ce6c;
  wire v134ce6d;
  wire v134ce6e;
  wire v134ce6f;
  wire v134ce70;
  wire v134ce71;
  wire v134ce72;
  wire v134ce73;
  wire v134ce74;
  wire v134ce75;
  wire v134ce76;
  wire v134ce77;
  wire v134ce78;
  wire v134ce79;
  wire v134ce7a;
  wire v134ce7b;
  wire v134ce7c;
  wire v134ce7d;
  wire v134ce7e;
  wire v134ce7f;
  wire v134ce80;
  wire v134ce81;
  wire v134ce82;
  wire v134ce83;
  wire v134ce84;
  wire v134ce85;
  wire v134ce86;
  wire v134ce87;
  wire v134ce88;
  wire v134ce89;
  wire v134ce8a;
  wire v134ce8b;
  wire v134ce8c;
  wire v134ce8d;
  wire v134ce8e;
  wire v134ce8f;
  wire v134ce90;
  wire v134ce91;
  wire v134ce92;
  wire v134ce93;
  wire v134ce94;
  wire v134ce95;
  wire v134ce96;
  wire v134ce97;
  wire v134ce98;
  wire v134ce99;
  wire v134ce9a;
  wire v134ce9b;
  wire v134ce9c;
  wire v134ce9d;
  wire v134ce9e;
  wire v134ce9f;
  wire v134cea0;
  wire v134cea1;
  wire v134cea2;
  wire v134cea3;
  wire v134cea4;
  wire v134cea5;
  wire v134cea6;
  wire v134cea7;
  wire v134cea8;
  wire v134cea9;
  wire v134ceb8;
  wire v134ceb9;
  wire v134ceba;
  wire v134cebb;
  wire v134cebc;
  wire v134cebd;
  wire v134cebe;
  wire v134cebf;
  wire v134cec0;
  wire v134cec1;
  wire v134cec2;
  wire v134cec3;
  wire v134cec4;
  wire v134cec5;
  wire v134cec6;
  wire v134cec7;
  wire v134cec8;
  wire v134cec9;
  wire v134ceca;
  wire v134cecb;
  wire v134cecc;
  wire v134cecd;
  wire v134cece;
  wire v134cecf;
  wire v134ced0;
  wire v134ced8;
  wire v134ced9;
  wire v134ceda;
  wire v134cedb;
  wire v134cedc;
  wire v134cedd;
  wire v134cede;
  wire v134cedf;
  wire v134cee0;
  wire v134cee1;
  wire v134cee2;
  wire v134cee3;
  wire v134cee4;
  wire v134cee5;
  wire v134cee6;
  wire v134cee7;
  wire v134cf3f;
  wire v134cf40;
  wire v134cf41;
  wire v134cf42;
  wire v134cf6a;
  wire v134cf6b;
  wire v134cf6c;
  wire v134cf6d;
  wire v134cf6e;
  wire v134cf6f;
  wire v134cf70;
  wire v138a2f7;
  wire v138a2f8;
  wire v138a2f9;
  wire v138a2fa;
  wire v138a2fb;
  wire v138a2fc;
  wire v138a2fd;
  wire v138a2fe;
  wire v138a2ff;
  wire v138a300;
  wire v138a301;
  wire v138a302;
  wire v138a303;
  wire v138a304;
  wire v138a305;
  wire v138a306;
  wire v138a307;
  wire v138a308;
  wire v138a309;
  wire v138a30a;
  wire v138a30b;
  wire v138a30c;
  wire v138a30d;
  wire v138a30e;
  wire v138a30f;
  wire v138a310;
  wire v138a311;
  wire v138a312;
  wire v138a313;
  wire v138a314;
  wire v138a315;
  wire v138a316;
  wire v138a317;
  wire v138a318;
  wire v138a319;
  wire v138a31a;
  wire v138a31b;
  wire v138a31c;
  wire v138a31d;
  wire v138a31e;
  wire v138a31f;
  wire v138a320;
  wire v845562;
  wire v138a321;
  wire v138a322;
  wire v138a323;
  wire v138a324;
  wire v138a325;
  wire v1180b7b;
  wire v138a326;
  wire v138a327;
  wire v138a328;
  wire v138a329;
  wire v138a32a;
  wire v138a32b;
  wire v138a32c;
  wire v138a32d;
  wire v138a32e;
  wire v138a32f;
  wire v138a330;
  wire v138a331;
  wire v138a332;
  wire v138a333;
  wire v138a334;
  wire v138a335;
  wire v138a336;
  wire v138a337;
  wire v138a338;
  wire v138a339;
  wire v138a33a;
  wire v138a33b;
  wire v138a33c;
  wire v138a33d;
  wire v138a33e;
  wire v138a33f;
  wire v138a340;
  wire v138a341;
  wire v138a342;
  wire v138a343;
  wire v138a344;
  wire v138a345;
  wire v138a346;
  wire v138a347;
  wire v138a348;
  wire v138a349;
  wire v138a34a;
  wire v138a34b;
  wire v138a34c;
  wire v138a34d;
  wire v138a34e;
  wire v138a34f;
  wire v138a350;
  wire v138a351;
  wire v138a352;
  wire v138a353;
  wire v138a354;
  wire v138a355;
  wire v138a356;
  wire v138a357;
  wire v138a358;
  wire v138a359;
  wire v138a35a;
  wire v138a35b;
  wire v138a35c;
  wire v138a35d;
  wire v138a35e;
  wire v138a35f;
  wire v138a360;
  wire v138a361;
  wire v138a362;
  wire v138a363;
  wire v138a364;
  wire v138a365;
  wire v138a366;
  wire v138a38e;
  wire v138a38f;
  wire v138a390;
  wire v138a391;
  wire v138a392;
  wire v138a393;
  wire v138a394;
  wire v138a395;
  wire v138a396;
  wire v138a397;
  wire v138a398;
  wire v138a399;
  wire v138a39a;
  wire v138a39b;
  wire v138a39c;
  wire v138a39d;
  wire v138a39e;
  wire v138a39f;
  wire v138a3a0;
  wire v138a3a1;
  wire v138a3a2;
  wire v138a3a3;
  wire v138a3a4;
  wire v138a3a5;
  wire v138a3a6;
  wire v138a3a7;
  wire v138a3a8;
  wire v138a3a9;
  wire v138a3aa;
  wire v138a3ab;
  wire v138a3ac;
  wire v138a3ad;
  wire v138a3ae;
  wire v138a3bf;
  wire v138a3c0;
  wire v138a3c1;
  wire v138a3c2;
  wire v138a3c3;
  wire v138a3c4;
  wire v138a3c5;
  wire v138a3c6;
  wire v138a3c7;
  wire v138a3c8;
  wire v138a3c9;
  wire v138a3ca;
  wire v138a3cb;
  wire v138a3cc;
  wire v138a3cd;
  wire v138a3ce;
  wire v138a3cf;
  wire v138a3d0;
  wire v138a3d1;
  wire v138a3d2;
  wire v138a3d3;
  wire v138a3d4;
  wire v138a3d5;
  wire v138a3d6;
  wire v138a3d7;
  wire v138a3d8;
  wire v138a3d9;
  wire v138a3da;
  wire v138a3db;
  wire v138a3dc;
  wire v138a3dd;
  wire v138a3de;
  wire v138a3df;
  wire v138a3e0;
  wire v138a3e1;
  wire v138a3e2;
  wire v138a3e3;
  wire v138a3e4;
  wire v138a3e5;
  wire v138a3e6;
  wire v138a3e7;
  wire v138a3e8;
  wire v138a3e9;
  wire v138a3ea;
  wire v138a3eb;
  wire v138a3ec;
  wire v138a3ed;
  wire v138a3ee;
  wire v138a3ef;
  wire v138a3f0;
  wire v138a3f1;
  wire v138a3f2;
  wire v138a3f3;
  wire v138a3f4;
  wire v138a3f5;
  wire v138a3f6;
  wire v138a3f7;
  wire v138a3f8;
  wire v138a3f9;
  wire v138a3fa;
  wire v138a3fb;
  wire v138a3fc;
  wire v84557c;
  wire v138a402;
  wire v138a403;
  wire v138a404;
  wire v138a405;
  wire v138a406;
  wire v138a407;
  wire v138a434;
  wire v138a435;
  wire v138a436;
  wire v138a437;
  wire v138a438;
  wire v138a439;
  wire v138a43a;
  wire v138a43b;
  wire v138a43c;
  wire v138a43d;
  wire v138a43e;
  wire v138a43f;
  wire v138a440;
  wire v138a441;
  wire v138a442;
  wire v138a443;
  wire v138a444;
  wire v138a445;
  wire v138a446;
  wire v138a447;
  wire v138a448;
  wire v138a449;
  wire v138a44a;
  wire v138a44b;
  wire v138a44c;
  wire v138a44d;
  wire v138a44e;
  wire v138a44f;
  wire v138a450;
  wire v138a451;
  wire v138a452;
  wire v138a453;
  wire v138a454;
  wire v138a455;
  wire v138a456;
  wire v138a457;
  wire v138a458;
  wire v138a459;
  wire v138a45a;
  wire v138a45b;
  wire v138a45c;
  wire v138a45d;
  wire v138a45e;
  wire v138a45f;
  wire v138a460;
  wire v138a461;
  wire v138a462;
  wire v138a463;
  wire v138a464;
  wire v138a475;
  wire v138a476;
  wire v138a477;
  wire v138a478;
  wire v138a479;
  wire v138a47a;
  wire v138a47b;
  wire v138a47c;
  wire v138a47d;
  wire v138a47e;
  wire v138a47f;
  wire v138a480;
  wire v138a481;
  wire v138a482;
  wire v138a483;
  wire v138a484;
  wire v138a485;
  wire v138a486;
  wire v138a487;
  wire v138a48d;
  wire v138a48e;
  wire v138a49f;
  wire v138a4a0;
  wire v138a4a1;
  wire v138a4a2;
  wire v1389d58;
  wire v1389d59;
  wire v1389d5a;
  wire v1389d5b;
  wire v1389d5c;
  wire v1389d71;
  wire v1389d72;
  wire v1389d73;
  wire v1389d74;
  wire v1389d75;
  wire v1389d76;
  wire v1389d77;
  wire v1389d78;
  wire v1389ddf;
  wire v1389de0;
  wire v1389de1;
  wire v1389de4;
  wire v1389de5;
  wire v1389de6;
  wire v1389de7;
  wire v1389df9;
  wire v1389dfa;
  wire v1389dfb;
  wire v1389e25;
  wire v1389e26;
  wire v1389e27;
  wire v1389e2a;
  wire v1389e2b;
  wire v1389e2c;
  wire v1389e2d;
  wire v1389e31;
  wire v1389e32;
  wire v1389e33;
  wire v1389e36;
  wire v1389e37;
  wire v1389efc;
  wire v1389efd;
  wire v1389efe;
  wire v1389f82;
  wire v1389f83;
  wire v1389f84;
  wire v1389f85;
  wire v1389f86;
  wire v1389f87;
  wire v1389f8b;
  wire v1389f8c;
  wire v1389f8d;
  wire v1389f8e;
  wire v1389f8f;
  wire v1389f90;
  wire v1389f91;
  wire v1389f92;
  wire v1389f93;
  wire v1389f94;
  wire v1389f97;
  wire v1389f98;
  wire v1389fb3;
  wire v1389fb4;
  wire v1389fb8;
  wire v1389fb9;
  wire v1389fba;
  wire v1389fbb;
  wire v1389fbc;
  wire v1389fbd;
  wire v1389fbe;
  wire v1389fbf;
  wire v1389fc0;
  wire v1389fc3;
  wire v1389fc4;
  wire v1389fca;
  wire v1389fcb;
  wire v1389fcc;
  wire v1389fcd;
  wire v1389fce;
  wire v1389fdb;
  wire v1389fdc;
  wire v1389fdd;
  wire v1389fe7;
  wire v1389fe8;
  wire v1389fe9;
  wire v1389ff2;
  wire v1389ff5;
  wire v1389ffb;
  wire v1389ffc;
  wire v1389ffd;
  wire v1389ffe;
  wire v1389fff;
  wire v138a000;
  wire v138a001;
  wire v138a002;
  wire v138a006;
  wire v138a007;
  wire v138a008;
  wire v138a010;
  wire v138a011;
  wire v138a02b;
  wire v138a02c;
  wire v138a02d;
  wire v138a02e;
  wire v138a032;
  wire v138a033;
  wire v138a034;
  wire v138a037;
  wire v138a038;
  wire v138a039;
  wire v138a03a;
  wire v138a059;
  wire v138a05a;
  wire v138a05b;
  wire v138a066;
  wire v138a067;
  wire v138a068;
  wire v138a069;
  wire v138a06a;
  wire v138a074;
  wire v138a075;
  wire v138a076;
  wire v138a07e;
  wire v138a07f;
  wire v138a090;
  wire v138a091;
  wire v138a092;
  wire v138a093;
  wire v138a0c6;
  wire v138a0c7;
  wire v1389538;
  wire v1389539;
  wire v138953a;
  wire v138953b;
  wire v138953c;
  wire v138959f;
  wire v13895a0;
  wire v13895a1;
  wire v13895a2;
  wire v13895a3;
  wire v13895a4;
  wire v13895a5;
  wire v13895a6;
  wire v13897dd;
  wire v13897de;
  wire v13897df;
  wire v13897e0;
  wire v13897ef;
  wire v13897f0;
  wire v13897f1;
  wire v1389808;
  wire v1389809;
  wire v138980a;
  wire v138980d;
  wire v138980e;
  wire v138980f;
  wire v1389810;
  wire v1389814;
  wire v1389815;
  wire v1389816;
  wire v1389817;
  wire v1389818;
  wire v1389819;
  wire v138981c;
  wire v138981d;
  wire v1389168;
  wire v1389169;
  wire v138916a;
  wire v13891a1;
  wire v13891a2;
  wire v13891a3;
  wire v13891a4;
  wire v13891a5;
  wire v13891a6;
  wire v13891a7;
  wire v13891a8;
  wire v138932c;
  wire v138932d;
  wire v138936c;
  wire v138936d;
  wire v138936e;
  wire v138936f;
  wire v1389370;
  wire v1389371;
  wire v1389372;
  wire v1389373;
  wire v1389374;
  wire v138937d;
  wire v138937e;
  wire v138937f;
  wire v1389380;
  wire v1389389;
  wire v138938a;
  wire v138938b;
  wire v138938c;
  wire v138938d;
  wire v138938e;
  wire v138938f;
  wire v1389390;
  wire v1389391;
  wire v1389392;
  wire v1389393;
  wire v1389394;
  wire v13893b5;
  wire v13893b6;
  wire v13893b7;
  wire v1389411;
  wire v1389430;
  wire v1389444;
  wire v1389445;
  wire v1389446;
  wire v1389447;
  wire v1389448;
  wire v1389449;
  wire v138944a;
  wire v138944b;
  wire v138944c;
  wire v138944d;
  wire v138944e;
  wire v138944f;
  wire v1389450;
  wire v1389451;
  wire v1389458;
  wire v1389459;
  wire v138945a;
  wire v138945b;
  wire v138945c;
  wire v138945d;
  wire v138945e;
  wire v138945f;
  wire v1389460;
  wire v1389461;
  wire v1389462;
  wire v1389463;
  wire v1389464;
  wire v1389465;
  wire v1389466;
  wire v1389498;
  wire v1389499;
  wire v138949a;
  wire v1388ce7;
  wire v1388ce8;
  wire v1388ce9;
  wire v140582a;
  wire v85e755;
  wire v1405838;
  wire v1405839;
  wire v140583a;
  wire v140583b;
  wire v140583c;
  wire v140583d;
  wire v85e70d;
  wire v140583e;
  wire v140583f;
  wire v1405840;
  wire v1405841;
  wire v1405842;
  wire v1405843;
  wire v1405844;
  wire v1405845;
  wire v1405846;
  wire v1405847;
  wire v1405848;
  wire v1405849;
  wire v140584a;
  wire v140584b;
  wire v140584c;
  wire v140584d;
  wire v140584e;
  wire v140584f;
  wire v1405850;
  wire v1405851;
  wire v1405852;
  wire v1405853;
  wire v1405854;
  wire v1405855;
  wire v1405856;
  wire v1405857;
  wire v1405858;
  wire v1405859;
  wire v140585a;
  wire v140585b;
  wire v140585c;
  wire v140585d;
  wire v140585e;
  wire v146b550;
  wire v140585f;
  wire v1405860;
  wire v1405861;
  wire v1405862;
  wire v1405863;
  wire v1405864;
  wire v1405865;
  wire v1405866;
  wire v1405867;
  wire v1405868;
  wire v1405869;
  wire v140586a;
  wire v140586b;
  wire v140586c;
  wire v140586d;
  wire v140586e;
  wire v140586f;
  wire v1405870;
  wire v1405871;
  wire v1405872;
  wire v1405873;
  wire v1405874;
  wire v1405875;
  wire v1405876;
  wire v1405877;
  wire v1405878;
  wire v1405879;
  wire v140587a;
  wire v140587b;
  wire v140587c;
  wire v140587d;
  wire v140587e;
  wire v140587f;
  wire v1405880;
  wire v1405881;
  wire v1405882;
  wire v1405883;
  wire v1405884;
  wire v1405885;
  wire v1405886;
  wire v1405887;
  wire v1405888;
  wire v1405889;
  wire v140588a;
  wire v140588b;
  wire v140588c;
  wire v140588d;
  wire v140588e;
  wire v140588f;
  wire v1405890;
  wire v1405891;
  wire v1405892;
  wire v1405893;
  wire v1405894;
  wire v1405895;
  wire v1405896;
  wire v1405897;
  wire v1405898;
  wire v1405899;
  wire v140589a;
  wire v140589b;
  wire v140589c;
  wire v140589d;
  wire v140589e;
  wire v140589f;
  wire v14058a0;
  wire v14058a1;
  wire v14058a2;
  wire v14058a3;
  wire v14058a4;
  wire v14058a5;
  wire v14058a6;
  wire v14058a7;
  wire v14058a8;
  wire v14058a9;
  wire v14058aa;
  wire v14058ab;
  wire v14058ac;
  wire v14058ad;
  wire v14058ae;
  wire v14058af;
  wire v14058b0;
  wire v14058b1;
  wire v14058b2;
  wire v14058b3;
  wire v14058b4;
  wire v14058b5;
  wire v14058b6;
  wire v14058b7;
  wire v14058b8;
  wire v14058b9;
  wire v14058ba;
  wire v14058bb;
  wire v14058bc;
  wire v14058bd;
  wire v14058be;
  wire v14058bf;
  wire v14058c0;
  wire v14058c1;
  wire v14058c2;
  wire v14058c3;
  wire v14058c4;
  wire v14058c5;
  wire v14058c6;
  wire v14058c7;
  wire v14058c8;
  wire v14058c9;
  wire v14058ca;
  wire v14058cb;
  wire v14058cc;
  wire v14058cd;
  wire v14058ce;
  wire v14058cf;
  wire v14058d0;
  wire v14058d1;
  wire v14058d2;
  wire v14058d3;
  wire v14058d4;
  wire v14058d5;
  wire v14058d6;
  wire v14058d7;
  wire v14058d8;
  wire v14058d9;
  wire v14058da;
  wire v14058db;
  wire v14058dc;
  wire v14058dd;
  wire v14058de;
  wire v14058df;
  wire v14058e0;
  wire v14058e1;
  wire v14058e2;
  wire v14058e3;
  wire v14058e4;
  wire v14058e5;
  wire v14058e6;
  wire v14058e7;
  wire v14058e8;
  wire v14058e9;
  wire v14058ea;
  wire v14058eb;
  wire v14058ec;
  wire v14058ed;
  wire v14058ee;
  wire v14058ef;
  wire v14058f0;
  wire v14058f1;
  wire v14058f2;
  wire v14058f3;
  wire v14058f4;
  wire v14058f5;
  wire v14058f6;
  wire v14058f7;
  wire v14058f8;
  wire v14058f9;
  wire v14058fa;
  wire v14058fb;
  wire v14058fc;
  wire v14058fd;
  wire v14058fe;
  wire v14058ff;
  wire v1405900;
  wire v1405901;
  wire v1405902;
  wire v1405903;
  wire v1405904;
  wire v1405905;
  wire v1405906;
  wire v1405907;
  wire v1405908;
  wire v1405909;
  wire v140590a;
  wire v140590b;
  wire v140590c;
  wire v140590d;
  wire v140590e;
  wire v140590f;
  wire v1405910;
  wire v1405911;
  wire v1405912;
  wire v1405913;
  wire v1405914;
  wire v1405915;
  wire v1405916;
  wire v1405917;
  wire v1405918;
  wire v1405919;
  wire v140591a;
  wire v140591b;
  wire v140591c;
  wire v140591d;
  wire v140591e;
  wire v140591f;
  wire v1405920;
  wire v1405921;
  wire v1405922;
  wire v1405923;
  wire v1405924;
  wire v1405925;
  wire v1405926;
  wire v1405927;
  wire v1405928;
  wire v1405929;
  wire v140592a;
  wire v140592b;
  wire v140592c;
  wire v140592d;
  wire v140592e;
  wire v140592f;
  wire v1405930;
  wire v1405931;
  wire v1405932;
  wire v1405933;
  wire v1405934;
  wire v1405935;
  wire v1405936;
  wire v1405937;
  wire v1405938;
  wire v1405939;
  wire v140593a;
  wire v140593b;
  wire v140593c;
  wire v140593d;
  wire v140593e;
  wire v140593f;
  wire v1405940;
  wire v1405941;
  wire v1405942;
  wire v85e75b;
  wire v1405a7d;
  wire v1405a7e;
  wire v1405a7f;
  wire v1405a80;
  wire v1405a84;
  wire v85e750;
  wire v1405a85;
  wire v1405a86;
  wire v1405a87;
  wire v1405a88;
  wire v1405a89;
  wire v1405a8a;
  wire v1405a8b;
  wire v1405a8c;
  wire v1405a8d;
  wire v1405a8e;
  wire v1405a8f;
  wire v1405a90;
  wire v1405a91;
  wire v1405a92;
  wire v1405a93;
  wire v1405a94;
  wire v1405a95;
  wire v1405a96;
  wire v1405a97;
  wire v1405a98;
  wire v1405a99;
  wire v1405a9a;
  wire v1405a9b;
  wire v1405a9c;
  wire v1405a9d;
  wire v1405a9e;
  wire v1405a9f;
  wire v1405aa0;
  wire v1405aa1;
  wire v1405aa2;
  wire v1405aa3;
  wire v1405aa4;
  wire v1405aa5;
  wire v1405aa6;
  wire v1405aa7;
  wire v1405aa8;
  wire v1405aa9;
  wire v1405aaa;
  wire v1405aab;
  wire v1405aac;
  wire v1405aad;
  wire v1405aae;
  wire v1405aaf;
  wire v1405ab0;
  wire v1405ab1;
  wire v1405ab2;
  wire v1405ab3;
  wire v1405ab4;
  wire v1405ab5;
  wire v1405ab6;
  wire v1405ab7;
  wire v1405ab8;
  wire v1405ab9;
  wire v1405aba;
  wire v1405abb;
  wire v1405abc;
  wire v1405abd;
  wire v1405abe;
  wire v1405abf;
  wire v1405ac0;
  wire v1405ac1;
  wire v1405ac2;
  wire v1405ac3;
  wire v1405ac4;
  wire v1405ac5;
  wire v1405ac6;
  wire v1405ac7;
  wire v1405ac8;
  wire v1405ac9;
  wire v1405aca;
  wire v1405acb;
  wire v1405acc;
  wire v1405acd;
  wire v1405ace;
  wire v1405acf;
  wire v1405ad0;
  wire v1405ad1;
  wire v1405ad2;
  wire v1405ad3;
  wire v1405ad4;
  wire v1405ad5;
  wire v1405ad6;
  wire v1405ad7;
  wire v1405ad8;
  wire v1405ad9;
  wire v1405ada;
  wire v1405adb;
  wire v1405adc;
  wire v1405add;
  wire v1405ade;
  wire v1405adf;
  wire v1405ae0;
  wire v1405ae1;
  wire v1405ae2;
  wire v1405ae3;
  wire v1405ae4;
  wire v1405ae5;
  wire v1405ae6;
  wire v1405ae7;
  wire v1405ae8;
  wire v1405ae9;
  wire v1405aea;
  wire v1405aeb;
  wire v1405aec;
  wire v1405aed;
  wire v1405aee;
  wire v1405aef;
  wire v1405af0;
  wire v1405af1;
  wire v1405af2;
  wire v1405af3;
  wire v1405af4;
  wire v1405af5;
  wire v1405af6;
  wire v1405af7;
  wire v1405af8;
  wire v1405af9;
  wire v1405afa;
  wire v1405afb;
  wire v1405afc;
  wire v1405afd;
  wire v1405afe;
  wire v1405aff;
  wire v1405b00;
  wire v1405b01;
  wire v1405b02;
  wire v1405b03;
  wire v1405b04;
  wire v1405b05;
  wire v1405b06;
  wire v1405b07;
  wire v1405b08;
  wire v1405b09;
  wire v1405b0a;
  wire v1405b0b;
  wire v1405b0c;
  wire v1405b0d;
  wire v1405b0e;
  wire v1405b0f;
  wire v1405b10;
  wire v1405b11;
  wire v1405b12;
  wire v1405b13;
  wire v1405b14;
  wire v1405b15;
  wire v1405b16;
  wire v1405b17;
  wire v1405b18;
  wire v1405b19;
  wire v1405b1a;
  wire v1405b1b;
  wire v1405b1c;
  wire v1405b1d;
  wire v1405b1e;
  wire v1405b1f;
  wire v1405b20;
  wire v1405b21;
  wire v1405b22;
  wire v1405b23;
  wire v1405b24;
  wire v1405b25;
  wire v1405b26;
  wire v1405b27;
  wire v1405b28;
  wire v1405b29;
  wire v1405b2a;
  wire v1405b2b;
  wire v1405b2c;
  wire v1405b2d;
  wire v1405b2e;
  wire v1405b2f;
  wire v1405b30;
  wire v1405b31;
  wire v1405b32;
  wire v1405b33;
  wire v1405b34;
  wire v1405b35;
  wire v1405b36;
  wire v1405b37;
  wire v1405b38;
  wire v1405b39;
  wire v1405b3a;
  wire v1405b3b;
  wire v1405b3c;
  wire v1405b3d;
  wire v1405b3e;
  wire v1405b3f;
  wire v1405b40;
  wire v1405b41;
  wire v1405b42;
  wire v1405b43;
  wire v1405b44;
  wire v1405b45;
  wire v1405b46;
  wire v1405b47;
  wire v1405b48;
  wire v1405b49;
  wire v1405b4a;
  wire v1405b4b;
  wire v1405b4c;
  wire v1405b4d;
  wire v1405b4e;
  wire v1405b4f;
  wire v1405b50;
  wire v1405b51;
  wire v1405b52;
  wire v1405b53;
  wire v1405b54;
  wire v1405b55;
  wire v1405b56;
  wire v1405b57;
  wire v1405b58;
  wire v1405b59;
  wire v1405b5a;
  wire v1405b5b;
  wire v1405b5c;
  wire v1405b5d;
  wire v1405b5e;
  wire v1405b5f;
  wire v1405b60;
  wire v1405b61;
  wire v1405b62;
  wire v1405b63;
  wire v1405b64;
  wire v1405b65;
  wire v1405b66;
  wire v1405b67;
  wire v1405b68;
  wire v1405b69;
  wire v12afda1;
  wire v12afda2;
  wire v12afda3;
  wire v12afda4;
  wire v12afda5;
  wire v12afda6;
  wire v12afda7;
  wire v12afda8;
  wire v12afda9;
  wire v12afdaa;
  wire v12afdab;
  wire v12afdac;
  wire v12afdad;
  wire v12afdae;
  wire v12afdaf;
  wire v12afdb0;
  wire v12afdb1;
  wire v12afdb2;
  wire v12afdb3;
  wire v12afdb4;
  wire v12afdb5;
  wire v12afe3b;
  wire v12afe3c;
  wire v12afe3d;
  wire v12afe3e;
  wire v12afe3f;
  wire v12afe40;
  wire v12afe44;
  wire v12afe45;
  wire v12afe46;
  wire v12afe47;
  wire v12afe4d;
  wire v12afe4e;
  wire v12afe4f;
  wire v12afe50;
  wire v12afe51;
  wire v12afe52;
  wire v12afe53;
  wire v12afe54;
  wire v12afe55;
  wire v12afe56;
  wire v12afe57;
  wire v12afe58;
  wire v12afe59;
  wire v12afe5a;
  wire v12afe5b;
  wire v12afe5c;
  wire v12afe5d;
  wire v12afe5e;
  wire v12afe5f;
  wire v12afe60;
  wire v12afe61;
  wire v12afe62;
  wire v12afe63;
  wire v12afe64;
  wire v12afe65;
  wire v12afe66;
  wire v12afe67;
  wire v12afe68;
  wire v12afe6f;
  wire v12afe70;
  wire v12afe71;
  wire v12afe72;
  wire v12afe73;
  wire v12afe74;
  wire v12afe75;
  wire v12afe76;
  wire v12afe77;
  wire v12af73c;
  wire v12af73d;
  wire v12af73e;
  wire v12af73f;
  wire v12af7e1;
  wire v12af7e2;
  wire v12af7f4;
  wire v12af7f5;
  wire v12af7f6;
  wire v12af7f7;
  wire v12af983;
  wire v12af984;
  wire v12af985;
  wire v12af986;
  wire v12af987;
  wire v12af988;
  wire v12af989;
  wire v12af98a;
  wire v12af98b;
  wire v12af98c;
  wire v12af98d;
  wire v12af98e;
  wire v12af98f;
  wire v12af9b1;
  wire v12af9b2;
  wire v12af9b3;
  wire v12af9b4;
  wire v12af9b5;
  wire v12af9b6;
  wire v12af9b7;
  wire v12af9b8;
  wire v12af9b9;
  wire v12af9bc;
  wire v12af9bd;
  wire v12af9be;
  wire v12af9bf;
  wire v12af9c0;
  wire v12af9c1;
  wire v12af9c2;
  wire v12af9c3;
  wire v12af9ce;
  wire v12af9cf;
  wire v12af9d0;
  wire v12af9d1;
  wire v12af9d2;
  wire v12af9d3;
  wire v12af9d4;
  wire v12af9d5;
  wire v12af9d6;
  wire v12af9d7;
  wire v12af9d8;
  wire v12af9d9;
  wire v12af9da;
  wire v12afa0a;
  wire v12afa0b;
  wire v12afa0c;
  wire v12afa0d;
  wire v12afa0e;
  wire v12afa0f;
  wire v12afa10;
  wire v12afa11;
  wire v12afa32;
  wire v12afa33;
  wire v12afa34;
  wire v12afa35;
  wire v12af3a4;
  wire v12af3a5;
  wire v12af3a6;
  wire v12af3a7;
  wire v12af3a8;
  wire v12af3a9;
  wire v12af3aa;
  wire v12af3ab;
  wire v12af3ac;
  wire v12af3ad;
  wire v12af3ae;
  wire v12af58d;
  wire v12af58e;
  wire v12af58f;
  wire v12af590;
  wire v12af5a2;
  wire v12af5a3;
  wire v12af5a4;
  wire v12af5a5;
  wire v12af5a6;
  wire v12af5a7;
  wire v12af5a8;
  wire v12af5a9;
  wire v12af5aa;
  wire v12af5ab;
  wire v12af5ac;
  wire v12af5ad;
  wire v12af5ae;
  wire v12af5af;
  wire v12af5b0;
  wire v12af5c4;
  wire v12aef09;
  wire v12aef0a;
  wire v12aef0b;
  wire v12af1b9;
  wire v12af1ba;
  wire v12af1bb;
  wire v12af1bc;
  wire v12af1bd;
  wire v12af1be;
  wire v12af1bf;
  wire v12af1c0;
  wire v12af1c1;
  wire v12af1c2;
  wire v12af1c3;
  wire v12af1c4;
  wire v12af21b;
  wire v12af21c;
  wire v12af21d;
  wire v12af21e;
  wire v12af21f;
  wire v12af220;
  wire v12af221;
  wire v12af222;
  wire v12af223;
  wire v12af224;
  wire v12af225;
  wire v12af226;
  wire v12af227;
  wire v12af228;
  wire v12af229;
  wire v12af22a;
  wire v12af22b;
  wire v12af22c;
  wire v12aead3;
  wire v12aead4;
  wire v12aead5;
  wire v12aead6;
  wire v12aead7;
  wire v12aeb18;
  wire v12aeb19;
  wire v12aeb1a;
  wire v12aeb1b;
  wire v12aeb1c;
  wire v12aeb1d;
  wire v12aeb1e;
  wire v12aeb1f;
  wire v12aeb22;
  wire v12aeb23;
  wire v12aeb40;
  wire v12aeb70;
  wire v12aeb71;
  wire v12aeb72;
  wire v12aeb73;
  wire v12aeb74;
  wire v12aeb75;
  wire v12aeb76;
  wire v12aeb77;
  wire v12aeb78;
  wire v12aeb7b;
  wire v12aeb7c;
  wire v12aeb82;
  wire v12aeb83;
  wire v12aeb84;
  wire v12aeb85;
  wire v12aec08;
  wire v12aec09;
  wire v12aec0a;
  wire v12aec0b;
  wire v12aec16;
  wire v12aec47;
  wire v12aec48;
  wire v12aec49;
  wire v12aec4a;
  wire v12aec4d;
  wire v12aec4e;
  wire v12aec4f;
  wire v12aecda;
  wire v12aecdb;
  wire v12aecdc;
  wire v12aed9e;
  wire v12aed9f;
  wire v12aedde;
  wire v12aee5c;
  wire v12aee5d;
  wire v12aee5e;
  wire v12aee5f;
  wire v12ae6da;
  wire v12ae6db;
  wire v12ae6fe;
  wire v12ae76a;
  wire v12ae76b;
  wire v12ae76c;
  wire v12ae83c;
  wire v12ae83d;
  wire v12ae83e;
  wire v12adf5d;
  wire v12adf5e;
  wire v12adf5f;
  wire v12adf60;
  wire v12adf61;
  wire v12adf62;
  wire v12adf63;
  wire v12adf64;
  wire v12adf65;
  wire v12adf66;
  wire v12adf67;
  wire v12ae1ef;
  wire v12ae1f0;
  wire v12ae1f1;
  wire v12ae1f2;
  wire v12ae1f3;
  wire v12ae1f4;
  wire v12ae1f5;
  wire v12ae1f6;
  wire v12ae1f7;
  wire v12ae1f8;
  wire v12ae1f9;
  wire v12ae1fa;
  wire v12ae1fb;
  wire v12ae1fc;
  wire v12ae1fd;
  wire v12ae1fe;
  wire v12ae1ff;
  wire v12ae200;
  wire v12ae201;
  wire v12ae209;
  wire v12adbea;
  wire v12adbeb;
  wire v12adbec;
  wire v12add46;
  wire v12add47;
  wire v12add48;
  wire v12add49;
  wire v12add4a;
  wire v12add4b;
  wire v12add4c;
  wire v12ad8e3;
  wire v12ad8e4;
  wire v12ad8e5;
  wire v12ad8e6;
  wire v12ad8e7;
  wire v12ad8e8;
  wire v12ad8e9;
  wire v12ad8ea;
  wire v12ad8eb;
  wire v12ad8ec;
  wire v12ad8ed;
  wire v12ad951;
  wire v12ad952;
  wire v12ad953;
  wire v12ad31a;
  wire v12ad31b;
  wire v12ad31c;
  wire v12ad31d;
  wire v12ad31e;
  wire v12ad31f;
  wire v12ad320;
  wire v12ad321;
  wire v12ad322;
  wire v12ad323;
  wire v12ad324;
  wire v12ad325;
  wire v12ad326;
  wire v12ad327;
  wire v12ad328;
  wire v12ad329;
  wire v12ad32a;
  wire v12ad32b;
  wire v12ad32c;
  wire v12ad32d;
  wire v12ad4be;
  wire v12ad4bf;
  wire v12ad4c0;
  wire v12ad4c1;
  wire v12ad4c2;
  wire v12ad4c3;
  wire v12ad4c4;
  wire v12ad4c5;
  wire v12ad4c6;
  wire v12ad4c7;
  wire v12ad4c8;
  wire v12ad4c9;
  wire v12ad4ca;
  wire v12ad4cc;
  wire v12ad4cd;
  wire v12ad4ce;
  wire v12ad4d0;
  wire v12ad4d1;
  wire v12ad4d2;
  wire v12ad4d3;
  wire v12ad4d4;
  wire v12ad4d5;
  wire v12ad4d6;
  wire v12ad4d7;
  wire v12ad4d8;
  wire v12ad4d9;
  wire v12ad4da;
  wire v12ad4db;
  wire v12ad4dc;
  wire v12ad4dd;
  wire v12ad4de;
  wire v12ad4df;
  wire v12ad4e0;
  wire v12ad4e1;
  wire v12ad4e2;
  wire v12ad4e3;
  wire v12ad4e4;
  wire v12ad4e5;
  wire v12ad4e6;
  wire v12ad4e7;
  wire v12ad4e8;
  wire v12ad4e9;
  wire v12ad4ea;
  wire v12ad4eb;
  wire v12ad4ec;
  wire v12ad4ed;
  wire v12ad4ee;
  wire v12ad4ef;
  wire v12ad4f0;
  wire v12ad4f1;
  wire v12ad4f2;
  wire v12ad4f3;
  wire v12ad4f4;
  wire v12ad4f5;
  wire v12ad4f6;
  wire v12ad4f7;
  wire v12ad4f8;
  wire v12ad4f9;
  wire v12ad4fa;
  wire v12ad4fb;
  wire v12ad4fc;
  wire v12ad4fd;
  wire v12ad4fe;
  wire v12ad4ff;
  wire v12ad500;
  wire v12ad501;
  wire v12ad502;
  wire v12ad503;
  wire v12ad504;
  wire v12ad505;
  wire v12ad506;
  wire v12ad507;
  wire v12ad508;
  wire v12ad509;
  wire v12ad50a;
  wire v12ad50b;
  wire v12ad50c;
  wire v12ad50d;
  wire v12ad50e;
  wire v12ad50f;
  wire v12ad510;
  wire v12ad511;
  wire v12ad512;
  wire v12ad513;
  wire v12ad514;
  wire v12ad515;
  wire v12ad516;
  wire v12ad517;
  wire v12ad518;
  wire v12ad519;
  wire v12ad51a;
  wire v12ad51b;
  wire v12ad51c;
  wire v12ad51d;
  wire v12ad51e;
  wire v12ad51f;
  wire v12ad520;
  wire v12ad521;
  wire v12ad522;
  wire v12ad523;
  wire v12ad524;
  wire v12ad525;
  wire v12ad526;
  wire v12ad527;
  wire v12ad528;
  wire v12ad529;
  wire v12ad52a;
  wire v12ad52b;
  wire v12ad52c;
  wire v12ad52d;
  wire v12ad52e;
  wire v12ad52f;
  wire v12ad530;
  wire v12ad531;
  wire v12ad532;
  wire v12ad533;
  wire v12ad534;
  wire v12ad535;
  wire v12ad536;
  wire v12ad537;
  wire v12ad538;
  wire v12ad539;
  wire v12ad53a;
  wire v12ad53b;
  wire v12ad53c;
  wire v12ad53d;
  wire v12ad53e;
  wire v12ad53f;
  wire v12ad540;
  wire v12ad541;
  wire v12ad542;
  wire v12ad543;
  wire v12ad544;
  wire v12ad545;
  wire v12ad546;
  wire v12ad547;
  wire v12ad548;
  wire v12ad549;
  wire v12ad54a;
  wire v12ad54b;
  wire v12ad54c;
  wire v12ad54d;
  wire v12ad54e;
  wire v12ad54f;
  wire v12ad550;
  wire v12ad551;
  wire v12ad552;
  wire v12ad553;
  wire v12ad554;
  wire v12ad555;
  wire v12ad556;
  wire v12ad557;
  wire v12ad558;
  wire v12ad559;
  wire v12ad55a;
  wire v12ad55b;
  wire v12ad55c;
  wire v12ad55d;
  wire v12ad55e;
  wire v12ad55f;
  wire v12ad560;
  wire v12ad561;
  wire v12ad562;
  wire v12ad563;
  wire v12ad564;
  wire v12ad565;
  wire v12ad566;
  wire v12ad567;
  wire v12ad568;
  wire v12ad569;
  wire v12ad56a;
  wire v12ad56b;
  wire v12ad56c;
  wire v12ad56d;
  wire v12ad56e;
  wire v12ad56f;
  wire v12ad570;
  wire v12ad571;
  wire v12ad572;
  wire v12ad573;
  wire v12ad574;
  wire v12ad575;
  wire v12ad576;
  wire v12ad577;
  wire v12ad578;
  wire v12ad579;
  wire v12ad57a;
  wire v12ad57b;
  wire v12ad57c;
  wire v12ad57d;
  wire v12ad57e;
  wire v12ad57f;
  wire v12ad580;
  wire v12ad581;
  wire v12ad582;
  wire v12ad583;
  wire v12ad584;
  wire v12ad585;
  wire v12ad586;
  wire v12ad587;
  wire v12ad588;
  wire v12ad589;
  wire v12ad58a;
  wire v12ad58b;
  wire v12ad58c;
  wire v12ad58d;
  wire v12ad58e;
  wire v12ad58f;
  wire v12ad590;
  wire v12ad591;
  wire v12ad592;
  wire v12ad593;
  wire v12ad594;
  wire v12ad595;
  wire v12ad596;
  wire v12ad597;
  wire v12ad598;
  wire v12ad599;
  wire v12ad59a;
  wire v12ad59c;
  wire v12ad59d;
  wire v12ad59e;
  wire v12ad59f;
  wire v12ad5a0;
  wire v12ad5a1;
  wire v12ad5a2;
  wire v12ad5a3;
  wire v12ad5a4;
  wire v12ad5a5;
  wire v12ad5a6;
  wire v12ad5a7;
  wire v12ad5a8;
  wire v12ad5a9;
  wire v12ad5aa;
  wire v12ad5ab;
  wire v12ad5ac;
  wire v12ad5ad;
  wire v12ad5ae;
  wire v12ad5af;
  wire v12ad5b0;
  wire v12ad5b1;
  wire v12ad5b2;
  wire v12ad5b3;
  wire v12ad5b4;
  wire v12ad5b5;
  wire v12ad5b6;
  wire v12ad5b7;
  wire v12ad5b8;
  wire v12ad5b9;
  wire v12ad5ba;
  wire v12ad5bb;
  wire v12ad5bc;
  wire v12ad5bd;
  wire v12ad5be;
  wire v12ad5bf;
  wire v12ad5c0;
  wire v12ad5c1;
  wire v12ad5c2;
  wire v12ad5c3;
  wire v12ad5c4;
  wire v12ad5c5;
  wire v12ad5c6;
  wire v12ad5c7;
  wire v12ad5c8;
  wire v12ad5c9;
  wire v12ad5ca;
  wire v12ad5cb;
  wire v12ad5cc;
  wire v12ad5cd;
  wire v12ad5ce;
  wire v12ad5cf;
  wire v12ad5d0;
  wire v12ad5d1;
  wire v12ad5d2;
  wire v12ad5d3;
  wire v12ad5d4;
  wire v12ad5d5;
  wire v12ad5d6;
  wire v12ad5d7;
  wire v12ad5d8;
  wire v12ad5d9;
  wire v12ad5da;
  wire v12ad5db;
  wire v12ad5dc;
  wire v12ad5dd;
  wire v12ad5de;
  wire v12ad5df;
  wire v12ad5e0;
  wire v12ad5e1;
  wire v12ad5e2;
  wire v12ad5e3;
  wire v12ad5e4;
  wire v12ad5e5;
  wire v12ad5e6;
  wire v12ad5e7;
  wire v12ad5e8;
  wire v12ad5e9;
  wire v12ad5ea;
  wire v12ad5eb;
  wire v12ad5ec;
  wire v12ad5ed;
  wire v12ad5ee;
  wire v12ad5ef;
  wire v12ad5f0;
  wire v12ad5f1;
  wire v12ad5f2;
  wire v12ad5f3;
  wire v12ad5f4;
  wire v12ad5f5;
  wire v12ad5f6;
  wire v12ad5f7;
  wire v12ad5f8;
  wire v12ad5f9;
  wire v12ad5fa;
  wire v12ad5fb;
  wire v12ad5fc;
  wire v12ad5fd;
  wire v12ad5fe;
  wire v12ad600;
  wire v12ad601;
  wire v12ad602;
  wire v12ad609;
  wire v12ad60b;
  wire v12ad60c;
  wire v12ad60d;
  wire v12ad60e;
  wire v12ad60f;
  wire v12ad610;
  wire v12ad611;
  wire v12ad612;
  wire v12ad613;
  wire v12ad614;
  wire v12ad615;
  wire v12ad616;
  wire v12ad617;
  wire v12ad618;
  wire v12ad619;
  wire v12ad61a;
  wire v12ad61b;
  wire v12ad61c;
  wire v12ad61d;
  wire v12ad61e;
  wire v12ad61f;
  wire v12ad620;
  wire v12ad621;
  wire v12ad622;
  wire v12ad623;
  wire v12ad624;
  wire v12ad625;
  wire v12ad626;
  wire v12ad627;
  wire v12ad62e;
  wire v12ad62f;
  wire v12ad630;
  wire v12ad631;
  wire v12ad632;
  wire v12ad633;
  wire v12ad634;
  wire v12ad635;
  wire v12ad643;
  wire v12ad644;
  wire v12ad645;
  wire v12ad65a;
  wire v12ad65b;
  wire v12ad65c;
  wire v12ad65d;
  wire v12ad65e;
  wire v12ad65f;
  wire v12ad660;
  wire v12ad661;
  wire v12ad662;
  wire v12ad663;
  wire v12ad664;
  wire v12ad665;
  wire v12ad666;
  wire v12ad667;
  wire v12ad668;
  wire v12ad669;
  wire v12ad66a;
  wire v12ad66b;
  wire v12ad66c;
  wire v12ad66d;
  wire v12ad66e;
  wire v12ad66f;
  wire v12ad670;
  wire v12ad671;
  wire v12ad672;
  wire v12ad673;
  wire v12ad674;
  wire v12ad675;
  wire v12ad676;
  wire v12ad677;
  wire v12ad678;
  wire v12ad679;
  wire v12ad67a;
  wire v12ad67b;
  wire v12ad67c;
  wire v12ad67d;
  wire v12ad67e;
  wire v12ad67f;
  wire v12ad680;
  wire v12ad681;
  wire v12acfb2;
  wire v12acfb3;
  wire v12acfb4;
  wire v12acfb5;
  wire v12acfb6;
  wire v12acfb7;
  wire v12acfb8;
  wire v12acfb9;
  wire v12acfba;
  wire v12acfbb;
  wire v12acfbc;
  wire v12acfbd;
  wire v12acfbe;
  wire v12acfbf;
  wire v12acfc0;
  wire v12acfc1;
  wire v12acfc2;
  wire v12acfc3;
  wire v12acfc4;
  wire v12acfc5;
  wire v12acfc6;
  wire v12acfc7;
  wire v12acfc8;
  wire v12acfc9;
  wire v12acfca;
  wire v12acfcb;
  wire v12acfcc;
  wire v12acfcd;
  wire v12acfce;
  wire v12acfcf;
  wire v12acfd0;
  wire v12acfd1;
  wire v12acfd2;
  wire v12acfd3;
  wire v12acfd4;
  wire v12acfd5;
  wire v12acfd6;
  wire v12acfd7;
  wire v12acfd8;
  wire v12acfd9;
  wire v12acfda;
  wire v12acfdb;
  wire v12acfdc;
  wire v12acfdd;
  wire v12acfde;
  wire v12acfdf;
  wire v12acfe0;
  wire v12acfe1;
  wire v12acfe2;
  wire v12acfe3;
  wire v12acfe4;
  wire v12acfe5;
  wire v12acfe6;
  wire v12acfe7;
  wire v12acfe8;
  wire v12acfe9;
  wire v12acfea;
  wire v12acfeb;
  wire v12acfec;
  wire v12acfed;
  wire v12acfee;
  wire v12acfef;
  wire v12acff0;
  wire v12acff1;
  wire v12acff2;
  wire v12acff3;
  wire v12acff4;
  wire v12acff5;
  wire v12acff6;
  wire v12acff7;
  wire v12acff8;
  wire v12acff9;
  wire v12acffa;
  wire v12acffb;
  wire v12acffc;
  wire v12acffd;
  wire v12acffe;
  wire v12acfff;
  wire v12ad000;
  wire v12ad001;
  wire v12ad002;
  wire v12ad003;
  wire v12ad004;
  wire v12ad005;
  wire v12ad006;
  wire v12ad007;
  wire v12ad008;
  wire v12ad009;
  wire v12ad00a;
  wire v12ad00b;
  wire v12ad00c;
  wire v12ad00d;
  wire v12ad00e;
  wire v12ad00f;
  wire v12ad010;
  wire v12ad011;
  wire v12ad012;
  wire v12ad013;
  wire v12ad014;
  wire v12ad015;
  wire v12ad016;
  wire v12ad017;
  wire v12ad018;
  wire v12ad019;
  wire v12ad01a;
  wire v12ad01b;
  wire v12ad01c;
  wire v12ad01d;
  wire v12ad01e;
  wire v12ad01f;
  wire v12ad020;
  wire v12ad021;
  wire v12ad022;
  wire v12ad023;
  wire v12ad024;
  wire v12ad025;
  wire v12ad026;
  wire v12ad027;
  wire v12ad028;
  wire v12ad029;
  wire v12ad02a;
  wire v12ad02b;
  wire v12ad02c;
  wire v12ad02d;
  wire v12ad02e;
  wire v12ad02f;
  wire v12ad030;
  wire v12ad031;
  wire v12ad032;
  wire v12ad033;
  wire v12ad034;
  wire v12ad035;
  wire v12ad036;
  wire v12ad039;
  wire v12ad03a;
  wire v12ad03b;
  wire v12ad03c;
  wire v12ad03d;
  wire v12ad0b0;
  wire v12ad0b1;
  wire v12ad0b2;
  wire v12ad0b3;
  wire v12ad0b4;
  wire v12ad0b5;
  wire v12ad0b6;
  wire v12ad0b7;
  wire v12ad0b8;
  wire v12ad0b9;
  wire v12ad0ba;
  wire v12ad0bb;
  wire v12ad0bc;
  wire v12ad0bd;
  wire v12ad0ca;
  wire v12ad0cb;
  wire v12ad0cc;
  wire v12ad13c;
  wire v12ad13d;
  wire v12ad13e;
  wire v12ad13f;
  wire v12ad140;
  wire v12ad1b0;
  wire v12ad1b1;
  wire v12ad1b3;
  wire v12ad1fc;
  wire v12ad1fd;
  wire v12ad1fe;
  wire v12ad1ff;
  wire v12ad22c;
  wire v12ad22d;
  wire v12ad22e;
  wire v12ad279;
  wire v12ad27a;
  wire v12ad27b;
  wire v12ad27c;
  wire v12acd05;
  wire v12acd06;
  wire v12acd07;
  wire v131be8a;
  wire v131be8b;
  wire v131be8c;
  wire v131be8d;
  wire v131be8e;
  wire v131be8f;
  wire v131be90;
  wire v1284c8d;
  wire v1284c8e;
  wire v1284c8f;
  wire v1284c90;
  wire v1284c91;
  wire v1284c92;
  wire v1284c93;
  wire v1284c94;
  wire v1284c95;
  wire v1284c96;
  wire v1284c97;
  wire v1284c98;
  wire v1284c99;
  wire v1284c9a;
  wire v1284c9b;
  wire v1284c9c;
  wire v1284c9d;
  wire v1284c9e;
  wire v1284c9f;
  wire v1284ca0;
  wire v1284ca1;
  wire v1284ca2;
  wire v1284ca3;
  wire v1284ca4;
  wire v1284ca5;
  wire v1284ca6;
  wire v1284ca7;
  wire v1284ca8;
  wire v1284ca9;
  wire v1284caa;
  wire v1284cab;
  wire v1284cac;
  wire v1284cad;
  wire v1284cae;
  wire v1284caf;
  wire v1284cb0;
  wire v1284cb1;
  wire v1284cb2;
  wire v1284cb3;
  wire v1284cb4;
  wire v1284cb5;
  wire v1284cb6;
  wire v1284cb7;
  wire v1284cb8;
  wire v1284cb9;
  wire v1284cba;
  wire v1284cbb;
  wire v1284cbc;
  wire v1284cbd;
  wire v1284cbe;
  wire v1284cbf;
  wire v1284cc0;
  wire v1284cc1;
  wire v1284cc2;
  wire v1284cc3;
  wire v1284cc4;
  wire v1284cc5;
  wire v1284cc6;
  wire v1284cc7;
  wire v1284cc8;
  wire v1284cc9;
  wire v1284cca;
  wire v1284ccb;
  wire v1284ccc;
  wire v1284ccd;
  wire v1284cce;
  wire v1284ccf;
  wire v1284cd0;
  wire v1284cd1;
  wire v1284cd2;
  wire v1284cd3;
  wire v1284cd4;
  wire v1284cd5;
  wire v1284cd6;
  wire v1284cd7;
  wire v1284cd8;
  wire v1284cd9;
  wire v1284cda;
  wire v1284cdb;
  wire v1284cdc;
  wire v1284cdd;
  wire v1284cde;
  wire v1284cdf;
  wire v1284ce0;
  wire v1284ce1;
  wire v1284ce2;
  wire v1284ce3;
  wire v1284ce5;
  wire v1284ce6;
  wire v1284ce7;
  wire v1284ce8;
  wire v1284ce9;
  wire v1284cea;
  wire v1284ceb;
  wire v1284cec;
  wire v1284ced;
  wire v1284cee;
  wire v1284cef;
  wire v1284cf0;
  wire v1284cf2;
  wire v1284cf3;
  wire v1284cf4;
  wire v1284cf5;
  wire v1284cf6;
  wire v1284cf7;
  wire v1284cf8;
  wire v1284cf9;
  wire v1284cfa;
  wire v1284cfb;
  wire v1284cfc;
  wire v1284cfd;
  wire v1284cfe;
  wire v1284cff;
  wire v1284d00;
  wire v1284d01;
  wire v1284d02;
  wire v1284d03;
  wire v1284d04;
  wire v1284d05;
  wire v1284d06;
  wire v1284d07;
  wire v1284d08;
  wire v1284d09;
  wire v1284d0a;
  wire v1284d0b;
  wire v1284d0c;
  wire v1284d0d;
  wire v1284d0e;
  wire v1284d0f;
  wire v1284d10;
  wire v1284d11;
  wire v1284d12;
  wire v1284d13;
  wire v1284d14;
  wire v1284d15;
  wire v1284d16;
  wire v1284d17;
  wire v1284d18;
  wire v1284d19;
  wire v1284d1a;
  wire v1284d1b;
  wire v1284d1c;
  wire v1284d1d;
  wire v1284d1e;
  wire v1284d1f;
  wire v1284d20;
  wire v1284d21;
  wire v1284d22;
  wire v1284d23;
  wire v1284d24;
  wire v1284d25;
  wire v1284d26;
  wire v1284d27;
  wire v1284d28;
  wire v1284d29;
  wire v1284d2a;
  wire v1284d2c;
  wire v1284d2d;
  wire v1284d2e;
  wire v1284d2f;
  wire v1284d30;
  wire v1284d31;
  wire v1284d32;
  wire v1284d33;
  wire v1284d34;
  wire v1284d35;
  wire v1284d36;
  wire v1284d37;
  wire v1284d39;
  wire v1284d3a;
  wire v1284d3b;
  wire v1284d3c;
  wire v1284d3d;
  wire v1284d3e;
  wire v1284d3f;
  wire v1284d40;
  wire v1284d41;
  wire v1284d42;
  wire v1284d43;
  wire v1284d44;
  wire v1284d45;
  wire v1284d46;
  wire v1284d47;
  wire v1284d48;
  wire v1284d49;
  wire v1284d4a;
  wire v1284d4b;
  wire v1284d4c;
  wire v1284d4d;
  wire v1284d4e;
  wire v1284d4f;
  wire v1284d50;
  wire v1284d51;
  wire v1284d52;
  wire v1284d53;
  wire v1284d54;
  wire v1284d55;
  wire v1284d56;
  wire v1284d57;
  wire v1284d58;
  wire v1284d59;
  wire v1284d5a;
  wire v1284d5b;
  wire v1284d5c;
  wire v1284d5d;
  wire v1284d5e;
  wire v1284d5f;
  wire v1284d60;
  wire v1284d61;
  wire v1284d62;
  wire v1284d63;
  wire v1284d64;
  wire v1284d65;
  wire v1284d66;
  wire v1284d67;
  wire v1284d68;
  wire v8b6f6a;
  wire v1284d69;
  wire v11e593a;
  wire v11e593b;
  wire v11e593c;
  wire v11e593d;
  wire v11e593e;
  wire v11e593f;
  wire v11e5940;
  wire v11e5941;
  wire v11e5942;
  wire v11e5943;
  wire v11e5944;
  wire v11e5945;
  wire v11e5946;
  wire v11e5947;
  wire v11e5948;
  wire v11e5949;
  wire v11e594a;
  wire v11e594b;
  wire v11e594c;
  wire v11e594d;
  wire v11e594e;
  wire v11e594f;
  wire v11e5950;
  wire v11e5951;
  wire v11e5952;
  wire v11e5953;
  wire v11e5954;
  wire v11e5955;
  wire v11e5956;
  wire v11e5957;
  wire v11e5958;
  wire v11e5959;
  wire v11e595a;
  wire v11e595b;
  wire v11e595c;
  wire v11e595d;
  wire v11e595e;
  wire v11e595f;
  wire v11e5960;
  wire v11e5961;
  wire v11e5962;
  wire v11e5963;
  wire v11e5964;
  wire v11e5965;
  wire v11e5966;
  wire v11e5967;
  wire v11e5968;
  wire v11e5969;
  wire v11e596a;
  wire v11e596b;
  wire v11e596c;
  wire v11e596d;
  wire v11e596e;
  wire v11e596f;
  wire v11e5970;
  wire v11e5971;
  wire v11e5972;
  wire v11e5973;
  wire v11e5974;
  wire v11e5975;
  wire v11e5976;
  wire v11e5977;
  wire v11e5978;
  wire v11e5979;
  wire v11e597a;
  wire v11e597b;
  wire v11e597c;
  wire v11e597d;
  wire v11e597e;
  wire v11e597f;
  wire v11e5980;
  wire v11e5981;
  wire v11e5982;
  wire v11e5983;
  wire v1216a5a;
  wire v1216a5b;
  wire v1216a5c;
  wire v1216a5d;
  wire v1216a5e;
  wire v1216a5f;
  wire v1216a60;
  wire v1216a61;
  wire v1216a62;
  wire v1216a63;
  wire v1216a64;
  wire v1216a65;
  wire v1216a66;
  wire v1216a67;
  wire v1216a68;
  wire v1216a69;
  wire v1216a6a;
  wire v1216a6b;
  wire v1216a6c;
  wire v1216a6d;
  wire v1216a6e;
  wire v1216a6f;
  wire v1216a70;
  wire v1216a71;
  wire v1216a72;
  wire v1216a73;
  wire v1216a74;
  wire v1216a75;
  wire v1216a76;
  wire v1216a77;
  wire v1216a78;
  wire v1216a79;
  wire v1216a7a;
  wire v1216a7b;
  wire v1216a7c;
  wire v1216a7d;
  wire v1216a7e;
  wire v1216a7f;
  wire v1216a80;
  wire v1216a81;
  wire v1216a82;
  wire v1216a83;
  wire v1216a84;
  wire v118e18f;
  wire v1216a85;
  wire v1216a86;
  wire v1216a87;
  wire v1216a88;
  wire v1216a89;
  wire v1216a8a;
  wire v1216a8b;
  wire v1216a8c;
  wire v1216a8d;
  wire v1216a8e;
  wire v1216a8f;
  wire v1216a90;
  wire v1216a91;
  wire v1216a92;
  wire v1216a93;
  wire v1216a94;
  wire v1216a95;
  wire v1216a96;
  wire v1216a97;
  wire v1216a98;
  wire v1216a99;
  wire v1216a9a;
  wire v1216a9b;
  wire v1216a9c;
  wire v1216a9d;
  wire v1216a9e;
  wire v1216a9f;
  wire v1216aa0;
  wire v1216aa1;
  wire v1216aa2;
  wire v1216aa3;
  wire v1216aa4;
  wire v1216aa5;
  wire v1216aa6;
  wire v1216aa7;
  wire v1216aa8;
  wire v1216aa9;
  wire v1216aac;
  wire v1216aad;
  wire v1216aae;
  wire v1216aaf;
  wire v1216ab0;
  wire v1216ab1;
  wire v1216ab2;
  wire v1216ab3;
  wire v1216ab8;
  wire v1216ab9;
  wire v1216aba;
  wire v1216abb;
  wire v1216abc;
  wire v1216abd;
  wire v1216abe;
  wire v1216ac3;
  wire v1216ac7;
  wire v1216acc;
  wire v1216acd;
  wire v1216ace;
  wire v1216acf;
  wire v1216ad0;
  wire v1216ad1;
  wire v1216ad2;
  wire v1216ad3;
  wire v1216ad4;
  wire v1216ad5;
  wire v1216ad6;
  wire v1216ada;
  wire v1216adb;
  wire v1216adc;
  wire v1216add;
  wire v1216ade;
  wire v1216adf;
  wire v1216ae3;
  wire v1216ae4;
  wire v1216ae5;
  wire v1216ae6;
  wire v1216aea;
  wire v1216aeb;
  wire v1216aec;
  wire v1216aed;
  wire v1216aee;
  wire v1216aef;
  wire v1216af3;
  wire v1216af4;
  wire v1216af5;
  wire v1216af6;
  wire v1216af7;
  wire v1216af8;
  wire v1216af9;
  wire v1216afa;
  wire v1216afb;
  wire v1216afc;
  wire v1216afd;
  wire v1216afe;
  wire v1216aff;
  wire v1216b00;
  wire v1216b01;
  wire v1216b02;
  wire v1216b03;
  wire v1216b04;
  wire v1216b05;
  wire v1216b06;
  wire v1216b07;
  wire v1216b08;
  wire v1216b0d;
  wire v1216b0e;
  wire v1216b0f;
  wire v1216b10;
  wire v1216b11;
  wire v1216b12;
  wire v1216b13;
  wire v1216b14;
  wire v1216b15;
  wire v1216b16;
  wire v1216b17;
  wire v12164c0;
  wire v12164c1;
  wire v12164c2;
  wire v12164c3;
  wire v12164c4;
  wire v12164c5;
  wire v12164c6;
  wire v12164c7;
  wire v12164c8;
  wire v12164c9;
  wire v12164ca;
  wire v12164cd;
  wire v12164ce;
  wire v12164cf;
  wire v12164d0;
  wire v12164d1;
  wire v12164d2;
  wire v12164d3;
  wire v12164d4;
  wire v12164d5;
  wire v12164d6;
  wire v12164d7;
  wire v12164d8;
  wire v12164d9;
  wire v12164da;
  wire v12164db;
  wire v12164dc;
  wire v12164dd;
  wire v12164de;
  wire v12164df;
  wire v12164e0;
  wire v12164e1;
  wire v12164e2;
  wire v12164e3;
  wire v12164e4;
  wire v12164e5;
  wire v12164e6;
  wire v12164e7;
  wire v1216518;
  wire v1216519;
  wire v121651a;
  wire v121651b;
  wire v121651c;
  wire v121651d;
  wire v121651e;
  wire v121651f;
  wire v1216520;
  wire v1216521;
  wire v1216522;
  wire v1216523;
  wire v1216524;
  wire v1216525;
  wire v1216526;
  wire v1216527;
  wire v1216528;
  wire v1216529;
  wire v121652a;
  wire v121652b;
  wire v121652c;
  wire v121652d;
  wire v121652e;
  wire v121652f;
  wire v1216530;
  wire v1216531;
  wire v1216532;
  wire v1216533;
  wire v1216534;
  wire v1216535;
  wire v1216536;
  wire v1216537;
  wire v1216538;
  wire v1216539;
  wire v121653a;
  wire v121653b;
  wire v121653c;
  wire v121653d;
  wire v121653e;
  wire v121653f;
  wire v1216540;
  wire v1216541;
  wire v1216542;
  wire v1216543;
  wire v1216544;
  wire v1216545;
  wire v1216546;
  wire v1216547;
  wire v1216548;
  wire v1216549;
  wire v121654a;
  wire v121654b;
  wire v121654c;
  wire v121654d;
  wire v121654e;
  wire v121654f;
  wire v1216550;
  wire v1216551;
  wire v1216552;
  wire v1216553;
  wire v1216554;
  wire v1216555;
  wire v1216556;
  wire v1216557;
  wire v1216558;
  wire v1216559;
  wire v121655a;
  wire v121655b;
  wire v121655c;
  wire v121655d;
  wire v121655e;
  wire v121655f;
  wire v1216560;
  wire v1216561;
  wire v1216562;
  wire v1216563;
  wire v1216564;
  wire v1216565;
  wire v1216566;
  wire v1216567;
  wire v1216568;
  wire v1216569;
  wire v121656a;
  wire v121656b;
  wire v121656c;
  wire v121656d;
  wire v121656e;
  wire v121656f;
  wire v1216570;
  wire v1216571;
  wire v1216572;
  wire v1216573;
  wire v1216574;
  wire v1216575;
  wire v1216576;
  wire v1216577;
  wire v1216578;
  wire v1216579;
  wire v121657a;
  wire v121657b;
  wire v121657c;
  wire v121657d;
  wire v121657e;
  wire v121657f;
  wire v1216580;
  wire v1216581;
  wire v1216582;
  wire v1216583;
  wire v1216584;
  wire v1216585;
  wire v1216586;
  wire v1216587;
  wire v1216588;
  wire v1216589;
  wire v121658a;
  wire v121658b;
  wire v121658c;
  wire v121658d;
  wire v121658e;
  wire v121658f;
  wire v1216590;
  wire v1216591;
  wire v1216592;
  wire v1216593;
  wire v1216594;
  wire v1216595;
  wire v1216596;
  wire v1216597;
  wire v1216598;
  wire v1216599;
  wire v121659a;
  wire v121659b;
  wire v121659c;
  wire v121659d;
  wire v121659e;
  wire v121659f;
  wire v12165a0;
  wire v12165a1;
  wire v12165a2;
  wire v12165a3;
  wire v12165a4;
  wire v12165a5;
  wire v12165a6;
  wire v12165a7;
  wire v12165a8;
  wire v12165a9;
  wire v12165aa;
  wire v12165ab;
  wire v12165ac;
  wire v12165ad;
  wire v12165ae;
  wire v12165af;
  wire v12165b0;
  wire v12165b1;
  wire v12165b2;
  wire v12165b3;
  wire v12165b4;
  wire v12166c1;
  wire v12166c2;
  wire v12166c3;
  wire v12166c4;
  wire v12166c5;
  wire v12166c6;
  wire v12166c7;
  wire v12166c8;
  wire v12166c9;
  wire v12166ca;
  wire v12166cb;
  wire v12166cc;
  wire v12166cd;
  wire v12166ce;
  wire v12166cf;
  wire v12166d0;
  wire v12166d1;
  wire v12166d2;
  wire v12166d3;
  wire v12166d4;
  wire v12166d5;
  wire v12166d6;
  wire v12166d7;
  wire v12166d8;
  wire v12166d9;
  wire v12166da;
  wire v12166db;
  wire v12166dc;
  wire v12166dd;
  wire v12166de;
  wire v12166df;
  wire v12166e0;
  wire v12166e1;
  wire v12166e2;
  wire v12166e3;
  wire v12166e4;
  wire v12166e5;
  wire v12166e6;
  wire v12166e7;
  wire v12166e8;
  wire v12166e9;
  wire v12166ea;
  wire v12166eb;
  wire v12166ec;
  wire v12166ed;
  wire v12166ee;
  wire v12166ef;
  wire v12166f0;
  wire v12166f1;
  wire v12166f2;
  wire v12166f3;
  wire v12166f4;
  wire v12166f5;
  wire v12166f6;
  wire v12166f7;
  wire v12166f8;
  wire v12166f9;
  wire v12166fa;
  wire v12166fb;
  wire v12166fc;
  wire v12166fd;
  wire v12166fe;
  wire v12166ff;
  wire v1216700;
  wire v1216701;
  wire v1216702;
  wire v1216703;
  wire v1216704;
  wire v1216705;
  wire v1216706;
  wire v1216707;
  wire v1216708;
  wire v1216709;
  wire v121670a;
  wire v121670b;
  wire v121670c;
  wire v121670d;
  wire v121670e;
  wire v121670f;
  wire v1216710;
  wire v1216711;
  wire v1216712;
  wire v1216713;
  wire v1216714;
  wire v1216715;
  wire v1216716;
  wire v1216717;
  wire v1216718;
  wire v1216719;
  wire v121671a;
  wire v121678b;
  wire v121678c;
  wire v121678d;
  wire v121678e;
  wire v121678f;
  wire v1216790;
  wire v1216791;
  wire v1216792;
  wire v1216793;
  wire v1216794;
  wire v1216795;
  wire v1216796;
  wire v1216799;
  wire v121679a;
  wire v121679b;
  wire v121679c;
  wire v121679d;
  wire v121679e;
  wire v121679f;
  wire v12167a0;
  wire v12167a1;
  wire v12167a2;
  wire v12167a3;
  wire v12167a4;
  wire v12167a5;
  wire v12167a6;
  wire v12167a7;
  wire v12167a8;
  wire v12167a9;
  wire v12167aa;
  wire v12167ab;
  wire v12167ac;
  wire v12167af;
  wire v1215fb2;
  wire v1215fb3;
  wire v1215fb4;
  wire v1215fb5;
  wire v1215fb6;
  wire v1215fb7;
  wire v1215fb8;
  wire v1215fb9;
  wire v1215fba;
  wire v1215fbb;
  wire v1215fbc;
  wire v1215fbd;
  wire v1215fbe;
  wire v1215fbf;
  wire v1215fc0;
  wire v1215fc1;
  wire v1215fe2;
  wire v1215fe3;
  wire v1215fe4;
  wire v1215fe5;
  wire v1215fe6;
  wire v1215fe7;
  wire v1215fe8;
  wire v1215fe9;
  wire v1215fea;
  wire v1215feb;
  wire v1215fec;
  wire v1215fed;
  wire v1215fee;
  wire v1215fef;
  wire v1215ff0;
  wire v1215ff1;
  wire v1215ff2;
  wire v1215ff3;
  wire v1215ff4;
  wire v1215ff5;
  wire v1215ff6;
  wire v1215ff7;
  wire v1215ff8;
  wire v1215ff9;
  wire v1215ffa;
  wire v1215ffb;
  wire v1215ffc;
  wire v1215ffd;
  wire v1215ffe;
  wire v1215fff;
  wire v1216000;
  wire v1216001;
  wire v1216002;
  wire v1216003;
  wire v1216004;
  wire v1216005;
  wire v1216006;
  wire v1216007;
  wire v1216008;
  wire v1216009;
  wire v121600a;
  wire v121600b;
  wire v121600c;
  wire v121600d;
  wire v121600e;
  wire v121600f;
  wire v1216010;
  wire v1216011;
  wire v1216012;
  wire v1216013;
  wire v1216014;
  wire v1216015;
  wire v1216016;
  wire v1216017;
  wire v1216018;
  wire v1216019;
  wire v121601a;
  wire v121601b;
  wire v121601c;
  wire v121601d;
  wire v121601e;
  wire v121601f;
  wire v1216020;
  wire v1216021;
  wire v1216022;
  wire v1216023;
  wire v1216024;
  wire v1216025;
  wire v1216026;
  wire v1216027;
  wire v1216028;
  wire v1216029;
  wire v121602a;
  wire v121602b;
  wire v121602c;
  wire v121602d;
  wire v121602e;
  wire v121602f;
  wire v1216030;
  wire v1216031;
  wire v1216032;
  wire v1216033;
  wire v1216034;
  wire v1216035;
  wire v1216036;
  wire v1216037;
  wire v1216038;
  wire v1216039;
  wire v121603a;
  wire v121603b;
  wire v121603c;
  wire v121603d;
  wire v121603e;
  wire v121603f;
  wire v1216040;
  wire v1216041;
  wire v1216042;
  wire v1216043;
  wire v1216044;
  wire v1216045;
  wire v1216046;
  wire v1216047;
  wire v1216048;
  wire v1216049;
  wire v121604a;
  wire v121604b;
  wire v121604c;
  wire v121604d;
  wire v121604e;
  wire v121604f;
  wire v1216050;
  wire v1216051;
  wire v1216052;
  wire v1216053;
  wire v1216054;
  wire v1216055;
  wire v1216056;
  wire v1216057;
  wire v1216058;
  wire v1216059;
  wire v121605a;
  wire v121605b;
  wire v121605c;
  wire v121605d;
  wire v121605e;
  wire v121605f;
  wire v1216060;
  wire v1216061;
  wire v1216062;
  wire v1216063;
  wire v1216064;
  wire v1216065;
  wire v1216066;
  wire v1216067;
  wire v1216068;
  wire v1216069;
  wire v121606a;
  wire v121606b;
  wire v121606c;
  wire v121606d;
  wire v121606e;
  wire v121606f;
  wire v1216070;
  wire v1216071;
  wire v1216072;
  wire v1216073;
  wire v1216074;
  wire v1216075;
  wire v1216076;
  wire v1216077;
  wire v1216078;
  wire v1216079;
  wire v121607a;
  wire v121607b;
  wire v121607c;
  wire v121607d;
  wire v121607e;
  wire v121607f;
  wire v1216080;
  wire v1216081;
  wire v1216082;
  wire v1216083;
  wire v1216084;
  wire v1216085;
  wire v1216086;
  wire v1216087;
  wire v1216088;
  wire v1216089;
  wire v121608a;
  wire v121608b;
  wire v121608c;
  wire v121608d;
  wire v121608e;
  wire v121608f;
  wire v1216090;
  wire v1216091;
  wire v1216092;
  wire v1216093;
  wire v1216094;
  wire v1216095;
  wire v1216096;
  wire v1216097;
  wire v1216098;
  wire v1216099;
  wire v121609a;
  wire v121609b;
  wire v121609c;
  wire v121609d;
  wire v121609e;
  wire v121609f;
  wire v12160a0;
  wire v12160a1;
  wire v12160a2;
  wire v12160a3;
  wire v12160a4;
  wire v12160a5;
  wire v12160a6;
  wire v12160a7;
  wire v12160a8;
  wire v12160a9;
  wire v12160aa;
  wire v12160ab;
  wire v12160ac;
  wire v12160ad;
  wire v12160ae;
  wire v12160af;
  wire v12160b0;
  wire v12160b1;
  wire v12160b2;
  wire v12160b3;
  wire v12160b4;
  wire v12160b5;
  wire v12160b6;
  wire v12160b7;
  wire v12160b8;
  wire v12160b9;
  wire v12160ba;
  wire v12160bb;
  wire v12160bc;
  wire v12160bd;
  wire v12160be;
  wire v12160bf;
  wire v12160c0;
  wire v12160c1;
  wire v12160c2;
  wire v12160c3;
  wire v12160c4;
  wire v12160c5;
  wire v12160c6;
  wire v12160c7;
  wire v12160c8;
  wire v12160c9;
  wire v12160ca;
  wire v12160cb;
  wire v12160cc;
  wire v12160cd;
  wire v12160ce;
  wire v12160cf;
  wire v12160d0;
  wire v12160d1;
  wire v12160d2;
  wire v12160d3;
  wire v12160d4;
  wire v12160d5;
  wire v12160d6;
  wire v12160d7;
  wire v12160d8;
  wire v12160d9;
  wire v12160da;
  wire v12160db;
  wire v12160dc;
  wire v12160dd;
  wire v12160de;
  wire v12160df;
  wire v12160e0;
  wire v12160e1;
  wire v12160e2;
  wire v12160e3;
  wire v12160e4;
  wire v12160e5;
  wire v12160e6;
  wire v12160e7;
  wire v12160e8;
  wire v12160e9;
  wire v12160ea;
  wire v12160eb;
  wire v12160ec;
  wire v12160ed;
  wire v12160ee;
  wire v12160ef;
  wire v12160f0;
  wire v12160f1;
  wire v12160f2;
  wire v12160f3;
  wire v12160f4;
  wire v12160f5;
  wire v12160f6;
  wire v12160f7;
  wire v12160f8;
  wire v12160f9;
  wire v12160fa;
  wire v12160fb;
  wire v12160fc;
  wire v12160fd;
  wire v12160fe;
  wire v12160ff;
  wire v1216100;
  wire v1216101;
  wire v1216102;
  wire v1216103;
  wire v1216104;
  wire v1216105;
  wire v1216106;
  wire v1216107;
  wire v1216108;
  wire v1216109;
  wire v121610a;
  wire v121610b;
  wire v121610c;
  wire v121610d;
  wire v121610e;
  wire v121610f;
  wire v1216110;
  wire v1216111;
  wire v1216112;
  wire v1216113;
  wire v1216114;
  wire v1216115;
  wire v1216116;
  wire v1216117;
  wire v1216118;
  wire v1216119;
  wire v121611a;
  wire v121611b;
  wire v121611c;
  wire v121611d;
  wire v121611e;
  wire v121611f;
  wire v1216120;
  wire v1216121;
  wire v1216122;
  wire v1216123;
  wire v1216124;
  wire v1216125;
  wire v1216126;
  wire v1216127;
  wire v1216128;
  wire v1216129;
  wire v121612a;
  wire v121612b;
  wire v121612c;
  wire v121612d;
  wire v121612e;
  wire v121612f;
  wire v1216130;
  wire v1216131;
  wire v1216132;
  wire v1216133;
  wire v1216134;
  wire v1216135;
  wire v1216136;
  wire v1216137;
  wire v1216138;
  wire v1216139;
  wire v121613a;
  wire v121613b;
  wire v121613c;
  wire v121613d;
  wire v121613e;
  wire v121613f;
  wire v1216140;
  wire v1216141;
  wire v1216142;
  wire v1216143;
  wire v1216144;
  wire v1216145;
  wire v1216146;
  wire v1216147;
  wire v1216148;
  wire v1216149;
  wire v121614a;
  wire v121614b;
  wire v121614c;
  wire v121614d;
  wire v121614e;
  wire v121614f;
  wire v1216150;
  wire v1216151;
  wire v1216152;
  wire v1216153;
  wire v1216154;
  wire v1216155;
  wire v1216156;
  wire v1216157;
  wire v1216158;
  wire v1216159;
  wire v121615a;
  wire v121615b;
  wire v121615c;
  wire v121615d;
  wire v121615e;
  wire v121615f;
  wire v1216160;
  wire v1216161;
  wire v1216162;
  wire v1216163;
  wire v1216164;
  wire v1216165;
  wire v1216166;
  wire v1216167;
  wire v1216168;
  wire v1216169;
  wire v121616a;
  wire v121616b;
  wire v121616c;
  wire v121616d;
  wire v121616e;
  wire v121616f;
  wire v1216170;
  wire v1216171;
  wire v1216172;
  wire v1216173;
  wire v1216174;
  wire v1216175;
  wire v1216176;
  wire v1216177;
  wire v1216178;
  wire v1216179;
  wire v121617a;
  wire v121617b;
  wire v121617c;
  wire v121617d;
  wire v121617e;
  wire v121617f;
  wire v1216180;
  wire v1216181;
  wire v1216182;
  wire v1216183;
  wire v1216184;
  wire v1216185;
  wire v1216186;
  wire v1216187;
  wire v1216188;
  wire v1216189;
  wire v121618a;
  wire v121618b;
  wire v121618c;
  wire v121618d;
  wire v121618e;
  wire v121618f;
  wire v1216190;
  wire v1216191;
  wire v1216192;
  wire v1216193;
  wire v1216194;
  wire v1216195;
  wire v1216196;
  wire v1216197;
  wire v1216198;
  wire v1216199;
  wire v121619a;
  wire v121619b;
  wire v121619c;
  wire v121619d;
  wire v121619e;
  wire v121619f;
  wire v12161a0;
  wire v12161a1;
  wire v12161a2;
  wire v12161a3;
  wire v12161a4;
  wire v12161a5;
  wire v12161a6;
  wire v12161a7;
  wire v12161a8;
  wire v12161a9;
  wire v12161aa;
  wire v12161ab;
  wire v12161ac;
  wire v12161ad;
  wire v12161ae;
  wire v12161af;
  wire v12161b0;
  wire v12161b1;
  wire v12161b2;
  wire v12161b3;
  wire v12161b4;
  wire v12161b5;
  wire v12161cc;
  wire v12161cd;
  wire v12161ce;
  wire v12161cf;
  wire v12161d0;
  wire v12161d1;
  wire v12161d2;
  wire v12161d3;
  wire v12161d4;
  wire v12161d5;
  wire v12161d6;
  wire v12161d7;
  wire v12161d8;
  wire v12161d9;
  wire v12161da;
  wire v12161db;
  wire v12161dc;
  wire v12161dd;
  wire v12161ec;
  wire v12161ed;
  wire v12161ee;
  wire v12161ef;
  wire v12161f0;
  wire v12161f1;
  wire v12161f2;
  wire v12161f3;
  wire v12161f4;
  wire v12161f5;
  wire v12161f6;
  wire v12161f7;
  wire v12161f8;
  wire v12161f9;
  wire v12161fa;
  wire v12161fb;
  wire v12161fc;
  wire v12161fd;
  wire v12161fe;
  wire v12161ff;
  wire v1216200;
  wire v1216201;
  wire v1216202;
  wire v1216203;
  wire v1216204;
  wire v1216205;
  wire v1216206;
  wire v1216207;
  wire v1216208;
  wire v1216209;
  wire v121620a;
  wire v121620b;
  wire v121620c;
  wire v121620d;
  wire v121620e;
  wire v121620f;
  wire v1216210;
  wire v1216211;
  wire v1216212;
  wire v1216213;
  wire v1216214;
  wire v1216215;
  wire v1216216;
  wire v1216217;
  wire v1216218;
  wire v1216219;
  wire v121621a;
  wire v121621b;
  wire v121621c;
  wire v121621d;
  wire v121621e;
  wire v121621f;
  wire v1216220;
  wire v1216221;
  wire v1216222;
  wire v1216223;
  wire v1216224;
  wire v1216225;
  wire v1216226;
  wire v1216227;
  wire v1216228;
  wire v1216229;
  wire v121622a;
  wire v121622b;
  wire v121622c;
  wire v121622d;
  wire v121622e;
  wire v121622f;
  wire v1216230;
  wire v1216231;
  wire v1216232;
  wire v1216233;
  wire v1216234;
  wire v1216235;
  wire v1216236;
  wire v1216237;
  wire v1216238;
  wire v1216239;
  wire v121623a;
  wire v121623b;
  wire v121623c;
  wire v121623d;
  wire v121623e;
  wire v121623f;
  wire v1216240;
  wire v1216241;
  wire v1216242;
  wire v1216243;
  wire v1216244;
  wire v1216245;
  wire v1216246;
  wire v1216247;
  wire v1216248;
  wire v1216249;
  wire v121624a;
  wire v121624b;
  wire v121624c;
  wire v121624d;
  wire v121624e;
  wire v121624f;
  wire v1216250;
  wire v1216251;
  wire v1216252;
  wire v1216253;
  wire v1216254;
  wire v1216255;
  wire v1216256;
  wire v1216257;
  wire v1216258;
  wire v1216259;
  wire v121625a;
  wire v121625b;
  wire v121625c;
  wire v121625d;
  wire v121625e;
  wire v121625f;
  wire v1216260;
  wire v1216261;
  wire v1216262;
  wire v1216263;
  wire v1216264;
  wire v1216265;
  wire v1216266;
  wire v1216267;
  wire v1216268;
  wire v1216269;
  wire v121626a;
  wire v121626b;
  wire v121626c;
  wire v121626d;
  wire v121626e;
  wire v121626f;
  wire v1216270;
  wire v1216271;
  wire v1216272;
  wire v1216273;
  wire v1216274;
  wire v1216275;
  wire v1216276;
  wire v1216277;
  wire v1216278;
  wire v1216279;
  wire v121627a;
  wire v121627b;
  wire v121627c;
  wire v121627d;
  wire v121627e;
  wire v121627f;
  wire v1216280;
  wire v1216281;
  wire v1216282;
  wire v1216283;
  wire v1216284;
  wire v1216285;
  wire v1216286;
  wire v1216287;
  wire v1216288;
  wire v1216289;
  wire v121628a;
  wire v121628b;
  wire v121628c;
  wire v121628d;
  wire v121628e;
  wire v121628f;
  wire v1216290;
  wire v1216291;
  wire v1216292;
  wire v1216293;
  wire v1216294;
  wire v1216295;
  wire v1216296;
  wire v1216297;
  wire v1216298;
  wire v1216299;
  wire v121629a;
  wire v121629b;
  wire v121629c;
  wire v121629d;
  wire v121629e;
  wire v121629f;
  wire v12162a0;
  wire v12162a1;
  wire v12162b2;
  wire v12162b3;
  wire v12162b4;
  wire v12162b5;
  wire v12162b6;
  wire v12162b7;
  wire v12162b8;
  wire v12162b9;
  wire v12162ba;
  wire v12162bb;
  wire v12162bc;
  wire v12162bd;
  wire v12162be;
  wire v12162bf;
  wire v12162c0;
  wire v12162c1;
  wire v12162c2;
  wire v12162c3;
  wire v12162c4;
  wire v12162c5;
  wire v12162c6;
  wire v12162c7;
  wire v12162c8;
  wire v12162c9;
  wire v12162ca;
  wire v12162cb;
  wire v12162cc;
  wire v12162cd;
  wire v12162ce;
  wire v12162cf;
  wire v12162d0;
  wire v12162d1;
  wire v12162d2;
  wire v12162d3;
  wire v12162d4;
  wire v12162d5;
  wire v12162d6;
  wire v12162d7;
  wire v12162d8;
  wire v12162d9;
  wire v12162da;
  wire v12162db;
  wire v12162dc;
  wire v12162dd;
  wire v12162de;
  wire v12162df;
  wire v12162e0;
  wire v12162e1;
  wire v12162e2;
  wire v12162e3;
  wire v12162e4;
  wire v12162e8;
  wire v12162e9;
  wire v12162ea;
  wire v12162eb;
  wire v12162ec;
  wire v12162ed;
  wire v12162ee;
  wire v12162ef;
  wire v12162f0;
  wire v12162f1;
  wire v12162f2;
  wire v12162f3;
  wire v12162f4;
  wire v12162f5;
  wire v12162f6;
  wire v12162f7;
  wire v12162f8;
  wire v12162f9;
  wire v12162fa;
  wire v12162fb;
  wire v12162fc;
  wire v12162fd;
  wire v12162fe;
  wire v12162ff;
  wire v1216300;
  wire v1216301;
  wire v1216302;
  wire v1216303;
  wire v1216304;
  wire v1216307;
  wire v1216308;
  wire v121630c;
  wire v121630d;
  wire v121630e;
  wire v121630f;
  wire v1216312;
  wire v1216313;
  wire v1216314;
  wire v1216318;
  wire v1216319;
  wire v121631a;
  wire v121631b;
  wire v121631c;
  wire v121631d;
  wire v121631e;
  wire v121631f;
  wire v1216320;
  wire v1216321;
  wire v1216322;
  wire v1216323;
  wire v1216326;
  wire v1216327;
  wire v121632b;
  wire v121632c;
  wire v121632f;
  wire v1216330;
  wire v1216399;
  wire v121639a;
  wire v121639e;
  wire v121639f;
  wire v12163a0;
  wire v12163a1;
  wire v12163a2;
  wire v12163a3;
  wire v12163a4;
  wire v12163a5;
  wire v12163a6;
  wire v12163a7;
  wire v12163a8;
  wire v12163a9;
  wire v12163aa;
  wire v12163ab;
  wire v12163ac;
  wire v12163ad;
  wire v1215bb4;
  wire v1215bb5;
  wire v1215bb6;
  wire v1215bb7;
  wire v1215bb8;
  wire v1215bbb;
  wire v1215bbf;
  wire v1215bc0;
  wire v1215bc1;
  wire v1215bc2;
  wire v1215bc3;
  wire v1215bc4;
  wire v1215bc5;
  wire v1215bc6;
  wire v1215bca;
  wire v1215bcb;
  wire v1215bcc;
  wire v1215bcd;
  wire v1215bd3;
  wire v1215bd4;
  wire v1215bd5;
  wire v1215bd7;
  wire v1215bd8;
  wire v1215bd9;
  wire v1215bda;
  wire v1215bdb;
  wire v1215bdc;
  wire v1215bdd;
  wire v1215bde;
  wire v1215bdf;
  wire v1215be0;
  wire v1215be1;
  wire v1215be2;
  wire v1215be3;
  wire v1215be4;
  wire v1215be5;
  wire v1215be6;
  wire v1215be7;
  wire v1215be8;
  wire v1215be9;
  wire v1215bea;
  wire v1215beb;
  wire v1215bec;
  wire v1215bed;
  wire v1215bef;
  wire v1215bf0;
  wire v1215bf1;
  wire v1215bf2;
  wire v1215bf3;
  wire v1215bf4;
  wire v1215bf5;
  wire v1215bf6;
  wire v1215bf7;
  wire v1215bf8;
  wire v1215bf9;
  wire v1215bfa;
  wire v1215bfb;
  wire v1215bfc;
  wire v1215bfd;
  wire v1215bfe;
  wire v1215bff;
  wire v1215c00;
  wire v1215c01;
  wire v1215c02;
  wire v1215c03;
  wire v1215c04;
  wire v1215c05;
  wire v1215c06;
  wire v1215c07;
  wire v1215c08;
  wire v1215c09;
  wire v1215c0a;
  wire v1215c0b;
  wire v1215c0c;
  wire v1215c0d;
  wire v1215c0e;
  wire v1215c0f;
  wire v1215c10;
  wire v1215c11;
  wire v1215c12;
  wire v1215c13;
  wire v1215c14;
  wire v1215c15;
  wire v1215c16;
  wire v1215c17;
  wire v1215c18;
  wire v1215c19;
  wire v1215c1a;
  wire v1215c1b;
  wire v1215c1c;
  wire v1215c1d;
  wire v1215c1e;
  wire v1215c1f;
  wire v1215c20;
  wire v1215c21;
  wire v1215c22;
  wire v1215c23;
  wire v1215c24;
  wire v1215c25;
  wire v1215c26;
  wire v1215c27;
  wire v1215c28;
  wire v1215c29;
  wire v1215c2a;
  wire v1215c2b;
  wire v1215c2c;
  wire v1215c2d;
  wire v1215c2e;
  wire v1215c2f;
  wire v1215c30;
  wire v1215c31;
  wire v1215c32;
  wire v1215c33;
  wire v1215c34;
  wire v1215c35;
  wire v1215c36;
  wire v1215c37;
  wire v1215c38;
  wire v1215c39;
  wire v1215c3c;
  wire v1215c3d;
  wire v1215c3e;
  wire v1215c3f;
  wire v1215c40;
  wire v1215c41;
  wire v1215c42;
  wire v1215c43;
  wire v1215c44;
  wire v1215c45;
  wire v1215c46;
  wire v1215c47;
  wire v1215c48;
  wire v1215c49;
  wire v1215c4a;
  wire v1215c4b;
  wire v1215c4c;
  wire v1215c4d;
  wire v1215c4e;
  wire v1215c4f;
  wire v1215c50;
  wire v1215c51;
  wire v1215c52;
  wire v1215c54;
  wire v1215c55;
  wire v1215c56;
  wire v1215c57;
  wire v1215c58;
  wire v1215c59;
  wire v1215c5a;
  wire v1215c5b;
  wire v1215c5c;
  wire v1215c5d;
  wire v1215c5e;
  wire v1215c5f;
  wire v1215c60;
  wire v1215c61;
  wire v1215c62;
  wire v1215c63;
  wire v1215c64;
  wire v1215c65;
  wire v1215c66;
  wire v1215c67;
  wire v1215c68;
  wire v1215c69;
  wire v1215c6a;
  wire v1215c6b;
  wire v1215c6c;
  wire v1215c6f;
  wire v1215c70;
  wire v1215c71;
  wire v1215c72;
  wire v1215c73;
  wire v1215c74;
  wire v1215c75;
  wire v1215c76;
  wire v1215c77;
  wire v1215c78;
  wire v1215c79;
  wire v1215c7a;
  wire v1215c7b;
  wire v1215c7c;
  wire v1215c7d;
  wire v1215c7e;
  wire v1215c7f;
  wire v1215c80;
  wire v1215c81;
  wire v1215c82;
  wire v1215c83;
  wire v1215c84;
  wire v1215c85;
  wire v1215c87;
  wire v1215c88;
  wire v1215c89;
  wire v1215c8a;
  wire v1215c8b;
  wire v1215c8c;
  wire v1215c8d;
  wire v1215c8e;
  wire v1215c8f;
  wire v1215c90;
  wire v1215c91;
  wire v1215c92;
  wire v1215c93;
  wire v1215c94;
  wire v1215c95;
  wire v1215c96;
  wire v1215c97;
  wire v1215c98;
  wire v1215c99;
  wire v1215c9a;
  wire v1215c9b;
  wire v1215c9c;
  wire v1215c9d;
  wire v1215c9e;
  wire v1215c9f;
  wire v1215ca0;
  wire v1215ca1;
  wire v1215ca2;
  wire v1215ca3;
  wire v1215ca4;
  wire v1215ca5;
  wire v1215ca6;
  wire v1215ca7;
  wire v1215ca8;
  wire v1215ca9;
  wire v1215caa;
  wire v1215cab;
  wire v1215cac;
  wire v1215cad;
  wire v1215cae;
  wire v1215caf;
  wire v1215cb0;
  wire v1215cb1;
  wire v1215cb2;
  wire v1215cb3;
  wire v1215cb4;
  wire v1215cb5;
  wire v1215cb6;
  wire v1215cb7;
  wire v1215cb8;
  wire v1215cb9;
  wire v1215cba;
  wire v1215cbb;
  wire v1215cbc;
  wire v1215cbd;
  wire v1215cbe;
  wire v1215cbf;
  wire v1215cc0;
  wire v1215cc1;
  wire v1215cc2;
  wire v1215cc3;
  wire v1215cc4;
  wire v1215cc5;
  wire v1215cc6;
  wire v1215cc7;
  wire v1215cc8;
  wire v1215cc9;
  wire v1215cca;
  wire v1215ccd;
  wire v1215cce;
  wire v1215ccf;
  wire v1215cd0;
  wire v1215cd1;
  wire v1215cd2;
  wire v1215cd3;
  wire v1215cd4;
  wire v1215cd5;
  wire v1215cd6;
  wire v1215cd7;
  wire v1215cd8;
  wire v1215cd9;
  wire v1215cda;
  wire v1215cdb;
  wire v1215cdc;
  wire v1215cdd;
  wire v1215cde;
  wire v1215cdf;
  wire v1215ce0;
  wire v1215ce2;
  wire v1215ce3;
  wire v1215ce4;
  wire v1215ce5;
  wire v1215ce6;
  wire v1215ce7;
  wire v1215ce8;
  wire v1215ce9;
  wire v1215cea;
  wire v1215ceb;
  wire v1215cec;
  wire v1215ced;
  wire v1215cee;
  wire v1215cef;
  wire v1215cf0;
  wire v1215cf1;
  wire v1215cf2;
  wire v1215cf3;
  wire v1215cf4;
  wire v1215cf5;
  wire v1215cf6;
  wire v1215cf7;
  wire v1215cf8;
  wire v1215cf9;
  wire v1215cfa;
  wire v1215cfb;
  wire v1215cfc;
  wire v1215cff;
  wire v1215d00;
  wire v1215d01;
  wire v1215d02;
  wire v1215d03;
  wire v1215d04;
  wire v1215d05;
  wire v1215d06;
  wire v1215d07;
  wire v1215d08;
  wire v1215d09;
  wire v1215d0a;
  wire v1215d0b;
  wire v1215d0c;
  wire v1215d0d;
  wire v1215d27;
  wire v1215d28;
  wire v1215d29;
  wire v1215d2a;
  wire v1215d2b;
  wire v1215d2c;
  wire v1215d2e;
  wire v1215d2f;
  wire v1215d30;
  wire v1215d31;
  wire v1215d32;
  wire v1215d33;
  wire v1215d34;
  wire v1215d35;
  wire v1215d36;
  wire v1215d37;
  wire v1215d38;
  wire v1215d39;
  wire v1215d3a;
  wire v1215d3b;
  wire v1215d3c;
  wire v1215d3d;
  wire v1215d3e;
  wire v1215d41;
  wire v1215d42;
  wire v1215d43;
  wire v1215d44;
  wire v1215d45;
  wire v1215d46;
  wire v1215d47;
  wire v1215d63;
  wire v1215d64;
  wire v1215d65;
  wire v1215d66;
  wire v1215d67;
  wire v1215d68;
  wire v1215d69;
  wire v1215d6b;
  wire v1215d6c;
  wire v1215d6d;
  wire v1215d6e;
  wire v1215d6f;
  wire v1215d70;
  wire v1215d71;
  wire v1215d72;
  wire v1215d73;
  wire v1215d74;
  wire v1215d75;
  wire v1215d76;
  wire v1215d77;
  wire v1215d78;
  wire v1215d79;
  wire v1215d7a;
  wire v1215d7b;
  wire v1215d7c;
  wire v1215d7d;
  wire v1215d80;
  wire v1215d81;
  wire v1215d82;
  wire v1215d83;
  wire v1215d84;
  wire v1215d85;
  wire v1215d86;
  wire v1215d88;
  wire v1215d89;
  wire v1215d8a;
  wire v1215d8b;
  wire v1215d8e;
  wire v1215d8f;
  wire v1215d95;
  wire v1215d97;
  wire v1215d98;
  wire v1215d99;
  wire v1215d9a;
  wire v1215d9b;
  wire v1215d9c;
  wire v1215d9d;
  wire v1215da0;
  wire v1215da1;
  wire v1215da2;
  wire v1215da4;
  wire v1215da5;
  wire v1215da8;
  wire v1215da9;
  wire v1215dac;
  wire v1215dad;
  wire v1215dae;
  wire v1215daf;
  wire v1215db0;
  wire v1215dc1;
  wire v1215dc2;
  wire v1215dda;
  wire v1215ddb;
  wire v1215ddc;
  wire v1215ddd;
  wire v1215dde;
  wire v1215ddf;
  wire v1215b76;
  wire v1215b77;
  wire v1215b78;
  wire v1215b79;
  wire v1215b7a;
  wire v1215b7b;
  wire v1215b7c;
  wire v1215b7d;
  wire v1215b7e;
  wire v1215b7f;
  wire v1215b80;
  wire v1215b81;
  wire v1215b82;
  wire v1215b83;
  wire v1215b84;
  wire v1215b85;
  wire v1215b86;
  wire v1215b87;
  wire v1215b88;
  wire v1215b89;
  wire v1215b8a;
  wire v1215b8b;
  wire v1215b8c;
  wire v1215b8d;
  wire v1215b8e;
  wire v1215b8f;
  wire v1215b90;
  wire v1215b91;
  wire v1215b92;
  wire v1215b93;
  wire v1215b94;
  wire v1215b95;
  wire v1215b96;
  wire v1215b97;
  wire v1215b98;
  wire v1215b99;
  wire v1215b9a;
  wire v1215b9b;
  wire v1215b9c;
  wire v1215b9d;
  wire v1215b9e;
  wire v1215b9f;
  wire v1215ba0;
  wire v1215ba1;
  wire v1215ba2;
  wire v1215ba3;
  wire v1215ba4;
  wire v1215ba5;
  wire v1215ba6;
  wire v1215ba7;
  wire v1215ba8;
  wire v1215ba9;
  wire v1215baa;
  wire v1215bab;
  wire v1215bac;
  wire v1215bad;
  wire v1215bae;
  wire v1215baf;
  wire v1215bb0;
  wire v12153b4;
  wire v12153b5;
  wire v12153b6;
  wire v12153b7;
  wire v12153b8;
  wire v12153b9;
  wire v12153ba;
  wire v12153bb;
  wire v12153bc;
  wire v12153bd;
  wire v12153be;
  wire v12153bf;
  wire v12153c0;
  wire v12153c1;
  wire v12153c2;
  wire v12153c3;
  wire v12153c4;
  wire v12153cd;
  wire v12153ce;
  wire v12153cf;
  wire v12153d0;
  wire v12153d1;
  wire v12153d2;
  wire v12153d3;
  wire v12153d4;
  wire v12153d5;
  wire v12153d6;
  wire v12153d7;
  wire v12153d8;
  wire v12153d9;
  wire v12153da;
  wire v12153db;
  wire v12153dc;
  wire v12153dd;
  wire v12153de;
  wire v12153df;
  wire v12153e0;
  wire v12153e1;
  wire v12153e2;
  wire v12153e3;
  wire v12153e4;
  wire v12153e5;
  wire v12153e6;
  wire v12153e7;
  wire v12153e8;
  wire v12153e9;
  wire v12153ea;
  wire v12153eb;
  wire v12153ec;
  wire v12153ed;
  wire v12153ee;
  wire v12153ef;
  wire v12153f0;
  wire v12153f1;
  wire v12153f2;
  wire v12153f3;
  wire v12153f4;
  wire v12153f5;
  wire v12153f6;
  wire v12153f7;
  wire v12153f8;
  wire v12153f9;
  wire v12153fa;
  wire v12153fb;
  wire v12153fc;
  wire v12153fd;
  wire v12153fe;
  wire v1215407;
  wire v1215408;
  wire v1215409;
  wire v121540a;
  wire v121540b;
  wire v121540c;
  wire v121540d;
  wire v121540e;
  wire v121540f;
  wire v1215410;
  wire v1215411;
  wire v1215412;
  wire v1215413;
  wire v1215414;
  wire v1215415;
  wire v1215416;
  wire v1215417;
  wire v1215418;
  wire v1215419;
  wire v121541a;
  wire v121541b;
  wire v1215435;
  wire v1215436;
  wire v1215437;
  wire v1215438;
  wire v1215439;
  wire v121543a;
  wire v121543b;
  wire v121543c;
  wire v121543d;
  wire v121543e;
  wire v121543f;
  wire v1215440;
  wire v1215441;
  wire v1215442;
  wire v1215443;
  wire v1215444;
  wire v1215445;
  wire v1215446;
  wire v1215447;
  wire v1215448;
  wire v1215449;
  wire v121544a;
  wire v121544b;
  wire v121544c;
  wire v121544d;
  wire v121544e;
  wire v121544f;
  wire v1215450;
  wire v1215451;
  wire v1215452;
  wire v1215453;
  wire v1215454;
  wire v1215455;
  wire v1215456;
  wire v1215457;
  wire v1215458;
  wire v1215459;
  wire v121545a;
  wire v121545b;
  wire v121545c;
  wire v121545d;
  wire v121545e;
  wire v121545f;
  wire v1215460;
  wire v1215461;
  wire v1215462;
  wire v1215463;
  wire v1215464;
  wire v1215465;
  wire v1215466;
  wire v1215467;
  wire v1215468;
  wire v1215469;
  wire v121546a;
  wire v121546b;
  wire v121546c;
  wire v121546d;
  wire v121546e;
  wire v121546f;
  wire v1215470;
  wire v1215471;
  wire v1215472;
  wire v1215473;
  wire v1215474;
  wire v1215475;
  wire v1215476;
  wire v1215707;
  wire v1215708;
  wire v1215709;
  wire v121570a;
  wire v121570b;
  wire v121570c;
  wire v121570d;
  wire v121570e;
  wire v121570f;
  wire v1215710;
  wire v1215711;
  wire v1215712;
  wire v1215713;
  wire v1215714;
  wire v1215715;
  wire v1215716;
  wire v1215717;
  wire v1215718;
  wire v1215719;
  wire v121571a;
  wire v121571b;
  wire v121571c;
  wire v121571d;
  wire v121571e;
  wire v121571f;
  wire v1215720;
  wire v1215721;
  wire v1215722;
  wire v1215723;
  wire v1215724;
  wire v1215725;
  wire v1215726;
  wire v1215727;
  wire v1215728;
  wire v1215729;
  wire v121572a;
  wire v121572b;
  wire v121572c;
  wire v121572d;
  wire v121572e;
  wire v121572f;
  wire v1215730;
  wire v1215731;
  wire v1215732;
  wire v1215733;
  wire v1215734;
  wire v1215735;
  wire v1215736;
  wire v1215737;
  wire v1215738;
  wire v1215739;
  wire v121573a;
  wire v121573b;
  wire v121573c;
  wire v121573d;
  wire v121573e;
  wire v121573f;
  wire v1215740;
  wire v1215741;
  wire v1215742;
  wire v1215743;
  wire v1215744;
  wire v1215745;
  wire v1215746;
  wire v1215747;
  wire v1215748;
  wire v1215749;
  wire v121574a;
  wire v121574b;
  wire v121574c;
  wire v121574d;
  wire v121574e;
  wire v121574f;
  wire v1215750;
  wire v1215751;
  wire v1215752;
  wire v1215753;
  wire v1215754;
  wire v1215755;
  wire v1215756;
  wire v1215757;
  wire v1215758;
  wire v1215759;
  wire v121575a;
  wire v121575b;
  wire v121575c;
  wire v121575d;
  wire v121575e;
  wire v121575f;
  wire v1215760;
  wire v1215761;
  wire v1215762;
  wire v1215763;
  wire v1215764;
  wire v1215765;
  wire v1215766;
  wire v1215767;
  wire v1215768;
  wire v1215769;
  wire v121576a;
  wire v121576b;
  wire v121576c;
  wire v121576d;
  wire v121576e;
  wire v121576f;
  wire v1215770;
  wire v1215771;
  wire v1215772;
  wire v1215773;
  wire v1215774;
  wire v1215775;
  wire v1215776;
  wire v1215777;
  wire v1215778;
  wire v1215779;
  wire v121577a;
  wire v121577b;
  wire v121577c;
  wire v121577d;
  wire v121577e;
  wire v121577f;
  wire v1215780;
  wire v1215781;
  wire v1215782;
  wire v1215783;
  wire v1215784;
  wire v1215785;
  wire v1215786;
  wire v1215787;
  wire v1215788;
  wire v1215789;
  wire v121578a;
  wire v121578b;
  wire v121578c;
  wire v121578d;
  wire v121578e;
  wire v121578f;
  wire v1215790;
  wire v1215791;
  wire v1215792;
  wire v1215793;
  wire v1215794;
  wire v1215795;
  wire v1215796;
  wire v1215797;
  wire v1215798;
  wire v1215799;
  wire v121579a;
  wire v121579b;
  wire v121579c;
  wire v121579d;
  wire v121579e;
  wire v121579f;
  wire v12157a0;
  wire v12157a1;
  wire v12157a2;
  wire v12157a3;
  wire v12157a4;
  wire v12157a5;
  wire v12157a6;
  wire v12157a7;
  wire v12157a8;
  wire v12157a9;
  wire v12157aa;
  wire v12157ab;
  wire v12157ac;
  wire v12157ad;
  wire v12157ae;
  wire v12157af;
  wire v12157b0;
  wire v12157b1;
  wire v1214fb4;
  wire v1214fb5;
  wire v1214fb6;
  wire v1214fb7;
  wire v1214fb8;
  wire v1214fb9;
  wire v1214fba;
  wire v1214fbb;
  wire v1214fbc;
  wire v1214fbd;
  wire v1214fbe;
  wire v1214fbf;
  wire v1214fc0;
  wire v1214fc1;
  wire v1214fc2;
  wire v1214fc3;
  wire v1214fc4;
  wire v1214fc5;
  wire v1214fc6;
  wire v1214fc7;
  wire v1214fc8;
  wire v1214fc9;
  wire v1214fca;
  wire v1214fe1;
  wire v1214fe2;
  wire v1214fe3;
  wire v1214fe4;
  wire v1214fe5;
  wire v1214fe6;
  wire v1214fea;
  wire v1214feb;
  wire v1214fec;
  wire v1214fed;
  wire v1214fee;
  wire v1214fef;
  wire v1214ff0;
  wire v1214ff1;
  wire v1214ff5;
  wire v1214ff6;
  wire v1214ff7;
  wire v1214ff8;
  wire v1214ff9;
  wire v1214ffa;
  wire v1214ffe;
  wire v1214fff;
  wire v1215000;
  wire v1215001;
  wire v121500e;
  wire v121500f;
  wire v1215010;
  wire v1215011;
  wire v1215012;
  wire v1215013;
  wire v1215014;
  wire v1215015;
  wire v1215016;
  wire v1215017;
  wire v1215018;
  wire v1215019;
  wire v121501a;
  wire v121501b;
  wire v121501c;
  wire v121501d;
  wire v121501e;
  wire v121501f;
  wire v1215020;
  wire v1215021;
  wire v1215022;
  wire v1215023;
  wire v1215024;
  wire v1215025;
  wire v1215026;
  wire v1215027;
  wire v1215028;
  wire v1215029;
  wire v121502a;
  wire v121502b;
  wire v121502c;
  wire v121502d;
  wire v121502e;
  wire v121502f;
  wire v1215030;
  wire v1215031;
  wire v1215032;
  wire v1215033;
  wire v1215034;
  wire v1215035;
  wire v1215036;
  wire v1215037;
  wire v1215038;
  wire v1215039;
  wire v121503a;
  wire v121503b;
  wire v121503c;
  wire v121503d;
  wire v121503e;
  wire v121503f;
  wire v1215040;
  wire v1215041;
  wire v1215042;
  wire v1215043;
  wire v1215044;
  wire v1215045;
  wire v1215046;
  wire v1215047;
  wire v1215048;
  wire v1215049;
  wire v121504a;
  wire v121504b;
  wire v121504c;
  wire v121504d;
  wire v121504e;
  wire v121504f;
  wire v1215050;
  wire v1215051;
  wire v1215052;
  wire v1215053;
  wire v1215054;
  wire v1215055;
  wire v1215056;
  wire v1215057;
  wire v1215058;
  wire v1215059;
  wire v121505a;
  wire v121505b;
  wire v121505c;
  wire v121505d;
  wire v121505e;
  wire v121505f;
  wire v1215060;
  wire v1215061;
  wire v1215062;
  wire v1215063;
  wire v1215064;
  wire v1215065;
  wire v1215066;
  wire v1215067;
  wire v1215068;
  wire v1215069;
  wire v121506a;
  wire v121506b;
  wire v121506c;
  wire v121506d;
  wire v121506e;
  wire v121506f;
  wire v1215070;
  wire v1215071;
  wire v1215072;
  wire v1215073;
  wire v1215074;
  wire v1215075;
  wire v1215076;
  wire v1215077;
  wire v1215078;
  wire v1215079;
  wire v121507a;
  wire v121507b;
  wire v121507c;
  wire v121507d;
  wire v121507e;
  wire v121507f;
  wire v1215080;
  wire v1215081;
  wire v1215082;
  wire v1215083;
  wire v1215084;
  wire v1215085;
  wire v1215086;
  wire v1215087;
  wire v1215088;
  wire v1215089;
  wire v121508a;
  wire v121508b;
  wire v121508c;
  wire v121508d;
  wire v1215091;
  wire v1215092;
  wire v1215093;
  wire v1215094;
  wire v1215095;
  wire v1215096;
  wire v1215097;
  wire v1215098;
  wire v1215099;
  wire v121509a;
  wire v121509b;
  wire v121509c;
  wire v121509d;
  wire v121509e;
  wire v121509f;
  wire v12150a0;
  wire v12150a1;
  wire v12150a2;
  wire v12150a3;
  wire v12150a4;
  wire v12150a5;
  wire v12150a6;
  wire v12150a7;
  wire v12150a8;
  wire v12150a9;
  wire v12150aa;
  wire v12150ab;
  wire v12150ac;
  wire v12150ad;
  wire v12150ae;
  wire v12150af;
  wire v12150b0;
  wire v12150b1;
  wire v12150b2;
  wire v12150b3;
  wire v12150b4;
  wire v12150b5;
  wire v12150b6;
  wire v12150b7;
  wire v12150b8;
  wire v12150b9;
  wire v12150ba;
  wire v12150bb;
  wire v12150bc;
  wire v12150bd;
  wire v12150be;
  wire v12150bf;
  wire v12150c0;
  wire v12150c1;
  wire v12150c2;
  wire v12150c3;
  wire v12150c4;
  wire v12150c5;
  wire v12150c6;
  wire v12150c7;
  wire v12150c8;
  wire v12150c9;
  wire v12150ca;
  wire v12150cb;
  wire v12150cc;
  wire v12150cd;
  wire v12150ce;
  wire v12150cf;
  wire v12150d0;
  wire v12150d1;
  wire v12150d2;
  wire v12150d3;
  wire v12150d4;
  wire v12150dd;
  wire v12150de;
  wire v12150df;
  wire v12150e0;
  wire v12150e1;
  wire v12150e2;
  wire v12150e3;
  wire v12150ec;
  wire v12150ed;
  wire v12150ee;
  wire v12150ef;
  wire v12150f0;
  wire v12150f1;
  wire v12150f2;
  wire v12150f3;
  wire v12150f4;
  wire v12150f5;
  wire v12150f6;
  wire v12150f7;
  wire v12150f8;
  wire v12150f9;
  wire v12150fa;
  wire v12150fb;
  wire v12150fc;
  wire v1215108;
  wire v1215109;
  wire v121510a;
  wire v121510b;
  wire v121510c;
  wire v121510d;
  wire v121510e;
  wire v121510f;
  wire v1215110;
  wire v1215111;
  wire v1215112;
  wire v12152e4;
  wire v12152e5;
  wire v12152e6;
  wire v12152e7;
  wire v12152e8;
  wire v12152e9;
  wire v12152ea;
  wire v12152eb;
  wire v12152ec;
  wire v12152ed;
  wire v12152ee;
  wire v12152ef;
  wire v12152f0;
  wire v12152f1;
  wire v12152f2;
  wire v12152f3;
  wire v12152f4;
  wire v12152f5;
  wire v12152f6;
  wire v12152f7;
  wire v12152f8;
  wire v12152f9;
  wire v12152fa;
  wire v12152fb;
  wire v12152fc;
  wire v12152fd;
  wire v12152fe;
  wire v12152ff;
  wire v1215300;
  wire v1215301;
  wire v1215302;
  wire v1215313;
  wire v1215314;
  wire v1215315;
  wire v1215316;
  wire v1215317;
  wire v1215318;
  wire v1215319;
  wire v121531a;
  wire v121531b;
  wire v121531c;
  wire v121531d;
  wire v121531e;
  wire v121531f;
  wire v1215320;
  wire v1215321;
  wire v1215322;
  wire v1215323;
  wire v1215324;
  wire v1215325;
  wire v1215326;
  wire v1215327;
  wire v1215328;
  wire v1215329;
  wire v121532a;
  wire v121532b;
  wire v121532c;
  wire v121532d;
  wire v121532e;
  wire v121532f;
  wire v1215330;
  wire v1215331;
  wire v1215332;
  wire v1215333;
  wire v1215334;
  wire v1215335;
  wire v1215336;
  wire v1215337;
  wire v1215338;
  wire v1215339;
  wire v121533a;
  wire v121533b;
  wire v121533c;
  wire v121533d;
  wire v121533e;
  wire v121533f;
  wire v1215340;
  wire v1215341;
  wire v1215342;
  wire v1215343;
  wire v1215344;
  wire v1215345;
  wire v1215346;
  wire v1215347;
  wire v1215348;
  wire v1215349;
  wire v121534a;
  wire v121534b;
  wire v121534c;
  wire v121534d;
  wire v121534e;
  wire v121534f;
  wire v1215350;
  wire v1215351;
  wire v1215352;
  wire v1215353;
  wire v1215354;
  wire v1215355;
  wire v1215356;
  wire v1215357;
  wire v1215358;
  wire v1215359;
  wire v121535a;
  wire v121535b;
  wire v121535c;
  wire v121535d;
  wire v121535e;
  wire v121535f;
  wire v1215360;
  wire v1215361;
  wire v1215362;
  wire v1215363;
  wire v1215364;
  wire v1215365;
  wire v1215366;
  wire v1215367;
  wire v1215368;
  wire v1215369;
  wire v121536a;
  wire v121536b;
  wire v121536c;
  wire v121536d;
  wire v121536e;
  wire v121536f;
  wire v1215370;
  wire v1215371;
  wire v1215372;
  wire v1215373;
  wire v1215374;
  wire v1215375;
  wire v1215376;
  wire v1215377;
  wire v1215378;
  wire v1215379;
  wire v121537a;
  wire v121537b;
  wire v121537c;
  wire v121537d;
  wire v121537e;
  wire v121537f;
  wire v1215380;
  wire v1215381;
  wire v1215382;
  wire v1215383;
  wire v1215384;
  wire v1215385;
  wire v1215386;
  wire v1215387;
  wire v1215388;
  wire v1215389;
  wire v121538a;
  wire v121538b;
  wire v121538c;
  wire v121538d;
  wire v121538e;
  wire v121538f;
  wire v1215390;
  wire v1215391;
  wire v1215392;
  wire v1215394;
  wire v1215395;
  wire v1215396;
  wire v1215398;
  wire v1215399;
  wire v121539a;
  wire v121539b;
  wire v121539c;
  wire v121539d;
  wire v121539e;
  wire v121539f;
  wire v12153a0;
  wire v12153a1;
  wire v12153a2;
  wire v12153a3;
  wire v12153a4;
  wire v12153a5;
  wire v12153a6;
  wire v12153a7;
  wire v12153a8;
  wire v12153a9;
  wire v12153aa;
  wire v12153ab;
  wire v12153ac;
  wire v12153ad;
  wire v12153ae;
  wire v12153af;
  wire v12153b0;
  wire v12153b1;
  wire v1214bb5;
  wire v1214bb6;
  wire v1214bb7;
  wire v1214bb8;
  wire v1214bb9;
  wire v1214bba;
  wire v1214bbb;
  wire v1214bbc;
  wire v1214bbd;
  wire v1214bbe;
  wire v1214bbf;
  wire v1214bc0;
  wire v1214bc1;
  wire v1214bc2;
  wire v1214bc3;
  wire v1214bc4;
  wire v1214bc5;
  wire v1214bc6;
  wire v1214bc7;
  wire v1214bc8;
  wire v1214bc9;
  wire v1214bca;
  wire v1214bcb;
  wire v1214bcc;
  wire v1214bcd;
  wire v1214bce;
  wire v1214bcf;
  wire v1214bd0;
  wire v1214bd1;
  wire v1214bd2;
  wire v1214bd3;
  wire v1214bd4;
  wire v1214bd5;
  wire v1214bd6;
  wire v1214bd7;
  wire v1214bd8;
  wire v1214bd9;
  wire v1214bda;
  wire v1214bdb;
  wire v1214bdc;
  wire v1214bf0;
  wire v1214bf1;
  wire v1214bf2;
  wire v1214bf3;
  wire v1214bf4;
  wire v1214bf5;
  wire v1214bf6;
  wire v1214bf7;
  wire v1214bf8;
  wire v1214bf9;
  wire v1214bfa;
  wire v1214bfb;
  wire v1214bfc;
  wire v1214bfd;
  wire v1214bfe;
  wire v1214bff;
  wire v1214c00;
  wire v1214c01;
  wire v1214c02;
  wire v1214c03;
  wire v1214c04;
  wire v1214c05;
  wire v1214c06;
  wire v1214c07;
  wire v1214c08;
  wire v1214c09;
  wire v1214c0a;
  wire v1214c0b;
  wire v1214c0c;
  wire v1214c0d;
  wire v1214c0e;
  wire v1214c0f;
  wire v1214c10;
  wire v1214c11;
  wire v1214c12;
  wire v1214c13;
  wire v1214c14;
  wire v1214c15;
  wire v1214c16;
  wire v1214c17;
  wire v1214c18;
  wire v1214c19;
  wire v1214c1a;
  wire v1214c1b;
  wire v1214c1c;
  wire v1214c1d;
  wire v1214c1e;
  wire v1214c1f;
  wire v1214c20;
  wire v1214c21;
  wire v1214c22;
  wire v1214c23;
  wire v1214c24;
  wire v1214c25;
  wire v1214c26;
  wire v1214c27;
  wire v1214c28;
  wire v1214c29;
  wire v1214c2a;
  wire v1214c2b;
  wire v1214c2c;
  wire v1214c2d;
  wire v1214c2e;
  wire v1214c2f;
  wire v1214c30;
  wire v1214c31;
  wire v1214c32;
  wire v1214c33;
  wire v1214c34;
  wire v1214c35;
  wire v1214c36;
  wire v1214c37;
  wire v1214c38;
  wire v1214c39;
  wire v1214c3a;
  wire v1214c3b;
  wire v1214c3c;
  wire v1214c3d;
  wire v1214c3e;
  wire v1214c3f;
  wire v1214c40;
  wire v1214c41;
  wire v1214c42;
  wire v1214c43;
  wire v1214c44;
  wire v1214c45;
  wire v1214c46;
  wire v1214c47;
  wire v1214c48;
  wire v1214c49;
  wire v1214c4a;
  wire v1214c4b;
  wire v1214c4c;
  wire v1214c4d;
  wire v1214c4e;
  wire v1214c4f;
  wire v1214c50;
  wire v1214c51;
  wire v1214c52;
  wire v1214c53;
  wire v1214c54;
  wire v1214c55;
  wire v1214c56;
  wire v1214c57;
  wire v1214c58;
  wire v1214c59;
  wire v1214c5a;
  wire v1214c5b;
  wire v1214c5c;
  wire v1214c5d;
  wire v1214c5e;
  wire v1214c5f;
  wire v1214c60;
  wire v1214c61;
  wire v1214c62;
  wire v1214c63;
  wire v1214c64;
  wire v1214c65;
  wire v1214c66;
  wire v1214c67;
  wire v1214c68;
  wire v1214c69;
  wire v1214c6a;
  wire v1214c6b;
  wire v1214c6c;
  wire v1214c6d;
  wire v1214c6e;
  wire v1214c6f;
  wire v1214c70;
  wire v1214c71;
  wire v1214c72;
  wire v1214c73;
  wire v1214c74;
  wire v1214c75;
  wire v1214c76;
  wire v1214c77;
  wire v1214c78;
  wire v1214c79;
  wire v1214c7a;
  wire v1214c7b;
  wire v1214c7c;
  wire v1214c7d;
  wire v1214c7e;
  wire v1214c7f;
  wire v1214c80;
  wire v1214c81;
  wire v1214c82;
  wire v1214c83;
  wire v1214c84;
  wire v1214c85;
  wire v1214c86;
  wire v1214c87;
  wire v1214c88;
  wire v1214c89;
  wire v1214c8a;
  wire v1214c8b;
  wire v1214c8c;
  wire v1214c8d;
  wire v1214c8e;
  wire v1214c8f;
  wire v1214c90;
  wire v1214c91;
  wire v1214c92;
  wire v1214c93;
  wire v1214c94;
  wire v1214c95;
  wire v1214c96;
  wire v1214c97;
  wire v1214c98;
  wire v1214c99;
  wire v1214c9a;
  wire v1214c9b;
  wire v1214c9c;
  wire v1214c9d;
  wire v1214c9e;
  wire v1214c9f;
  wire v1214ca0;
  wire v1214ca1;
  wire v1214ca2;
  wire v1214cb9;
  wire v1214cba;
  wire v1214cbb;
  wire v1214cbc;
  wire v1214cbd;
  wire v1214cbe;
  wire v1214cbf;
  wire v1214cc0;
  wire v1214cc1;
  wire v1214cc2;
  wire v1214cc3;
  wire v1214cc4;
  wire v1214cc5;
  wire v1214cc6;
  wire v1214cc7;
  wire v1214cc8;
  wire v1214cc9;
  wire v1214cca;
  wire v1214ccb;
  wire v1214ccc;
  wire v1214ccd;
  wire v1214cce;
  wire v1214ccf;
  wire v1214cd0;
  wire v1214cd1;
  wire v1214cd2;
  wire v1214cd3;
  wire v1214cd4;
  wire v1214cd5;
  wire v1214cd6;
  wire v1214cd7;
  wire v1214cd8;
  wire v1214cd9;
  wire v1214cda;
  wire v1214cdb;
  wire v1214cdc;
  wire v1214cdd;
  wire v1214cde;
  wire v1214cdf;
  wire v1214ce0;
  wire v1214ce1;
  wire v1214ce2;
  wire v1214ce3;
  wire v1214ce4;
  wire v1214ce5;
  wire v1214ce6;
  wire v1214ce7;
  wire v1214ce8;
  wire v1214ce9;
  wire v1214cea;
  wire v1214ceb;
  wire v1214cec;
  wire v1214ced;
  wire v1214cee;
  wire v1214cef;
  wire v1214cf0;
  wire v1214cf1;
  wire v1214cf2;
  wire v1214cf3;
  wire v1214cf4;
  wire v1214cf5;
  wire v1214cf6;
  wire v1214cf7;
  wire v1214cf8;
  wire v1214cf9;
  wire v1214cfa;
  wire v1214cfb;
  wire v1214cfc;
  wire v1214cfd;
  wire v1214cfe;
  wire v1214cff;
  wire v1214d00;
  wire v1214d01;
  wire v1214d02;
  wire v1214d03;
  wire v1214d04;
  wire v1214d05;
  wire v1214d06;
  wire v1214d07;
  wire v1214d08;
  wire v1214d09;
  wire v1214d0a;
  wire v1214d0b;
  wire v1214d0c;
  wire v1214d0d;
  wire v1214d0e;
  wire v1214d0f;
  wire v1214d10;
  wire v1214d11;
  wire v1214d12;
  wire v1214d13;
  wire v1214d14;
  wire v1214d15;
  wire v1214d16;
  wire v1214d17;
  wire v1214d18;
  wire v1214d19;
  wire v1214d1a;
  wire v1214d1b;
  wire v1214d1c;
  wire v1214d1d;
  wire v1214d1e;
  wire v1214d1f;
  wire v1214d20;
  wire v1214d21;
  wire v1214d22;
  wire v1214d23;
  wire v1214d24;
  wire v1214d25;
  wire v1214d26;
  wire v1214d27;
  wire v1214d28;
  wire v1214d29;
  wire v1214d2a;
  wire v1214d2b;
  wire v1214d2c;
  wire v1214d2d;
  wire v1214d2e;
  wire v1214d2f;
  wire v1214d30;
  wire v1214d31;
  wire v1214d32;
  wire v1214d33;
  wire v1214d34;
  wire v1214d35;
  wire v1214d36;
  wire v1214d37;
  wire v1214d38;
  wire v1214d39;
  wire v1214d3a;
  wire v1214d3b;
  wire v1214d3c;
  wire v1214d3d;
  wire v1214d3e;
  wire v1214d3f;
  wire v1214d40;
  wire v1214d41;
  wire v1214d42;
  wire v1214d43;
  wire v1214d44;
  wire v1214d45;
  wire v1214d46;
  wire v1214d47;
  wire v1214d48;
  wire v1214d49;
  wire v1214d4a;
  wire v1214d4b;
  wire v1214d4c;
  wire v1214d4d;
  wire v1214d4e;
  wire v1214d4f;
  wire v1214d50;
  wire v1214d51;
  wire v1214d52;
  wire v1214d53;
  wire v1214d54;
  wire v1214d55;
  wire v1214d56;
  wire v1214d57;
  wire v1214d58;
  wire v1214d59;
  wire v1214d5a;
  wire v1214d5b;
  wire v1214d5c;
  wire v1214d5d;
  wire v1214d5e;
  wire v1214d5f;
  wire v1214d60;
  wire v1214d61;
  wire v1214d62;
  wire v1214d63;
  wire v1214d64;
  wire v1214d65;
  wire v1214d66;
  wire v1214d67;
  wire v1214d68;
  wire v1214d69;
  wire v1214d6a;
  wire v1214d6b;
  wire v1214d6c;
  wire v1214d6d;
  wire v1214d6e;
  wire v1214d6f;
  wire v1214d70;
  wire v1214d71;
  wire v1214d72;
  wire v1214d73;
  wire v1214d74;
  wire v1214d75;
  wire v1214d76;
  wire v1214d77;
  wire v1214d78;
  wire v1214d79;
  wire v1214d7a;
  wire v1214d7b;
  wire v1214d7c;
  wire v1214d7d;
  wire v1214d7e;
  wire v1214d7f;
  wire v1214d80;
  wire v1214d81;
  wire v1214d82;
  wire v1214d83;
  wire v1214d84;
  wire v1214d85;
  wire v1214d86;
  wire v1214d87;
  wire v1214d88;
  wire v1214d89;
  wire v1214d8a;
  wire v1214d8b;
  wire v1214d9c;
  wire v1214d9d;
  wire v1214d9e;
  wire v1214d9f;
  wire v1214da0;
  wire v1214da1;
  wire v1214da2;
  wire v1214da3;
  wire v1214da4;
  wire v1214da5;
  wire v1214da6;
  wire v1214da7;
  wire v1214da8;
  wire v1214da9;
  wire v1214daa;
  wire v1214dab;
  wire v1214dac;
  wire v1214dad;
  wire v1214dae;
  wire v1214daf;
  wire v1214db0;
  wire v1214db1;
  wire v1214db2;
  wire v1214db3;
  wire v1214db4;
  wire v1214db5;
  wire v1214db6;
  wire v1214db7;
  wire v1214db8;
  wire v1214db9;
  wire v1214dba;
  wire v1214dbb;
  wire v1214dbc;
  wire v1214dbd;
  wire v1214dbe;
  wire v1214dbf;
  wire v1214dc0;
  wire v1214dc1;
  wire v1214dc2;
  wire v1214dc3;
  wire v1214dc4;
  wire v1214dc5;
  wire v1214dc6;
  wire v1214dc7;
  wire v1214dc8;
  wire v1214dc9;
  wire v1214dca;
  wire v1214dcb;
  wire v1214dcc;
  wire v1214dcd;
  wire v1214dce;
  wire v1214dcf;
  wire v1214dd0;
  wire v1214dd1;
  wire v1214dd2;
  wire v1214dd3;
  wire v1214dd4;
  wire v1214dd5;
  wire v1214dd6;
  wire v1214dd7;
  wire v1214dd8;
  wire v1214dd9;
  wire v1214dda;
  wire v1214ddb;
  wire v1214ddc;
  wire v1214ddd;
  wire v1214dde;
  wire v1214ddf;
  wire v1214de0;
  wire v1214de1;
  wire v1214de2;
  wire v1214de3;
  wire v1214dea;
  wire v1214df1;
  wire v1214df2;
  wire v1214df3;
  wire v1214df4;
  wire v1214df5;
  wire v1214df6;
  wire v1214df7;
  wire v1214e0b;
  wire v1214e0c;
  wire v1214e0d;
  wire v1214e0e;
  wire v1214e0f;
  wire v1214e10;
  wire v1214e1a;
  wire v1214e40;
  wire v1214e41;
  wire v1214e42;
  wire v1214e50;
  wire v1214e57;
  wire v1214e58;
  wire v1214e59;
  wire v1214e5a;
  wire v1214e5b;
  wire v1214e62;
  wire v1214e63;
  wire v1214e64;
  wire v1214e65;
  wire v1214e66;
  wire v1214e67;
  wire v1214e6e;
  wire v1214e6f;
  wire v1214e70;
  wire v1214e71;
  wire v1214e72;
  wire v1214e73;
  wire v1214e74;
  wire v1214e7b;
  wire v1214e7c;
  wire v1214e7d;
  wire v1214e7e;
  wire v1214e7f;
  wire v1214e80;
  wire v1214e81;
  wire v1214e82;
  wire v1214eb2;
  wire v1214eb3;
  wire v1214eb4;
  wire v1214eb5;
  wire v1214eb6;
  wire v1214eb7;
  wire v1214eb8;
  wire v1214eb9;
  wire v1214eba;
  wire v1214ebb;
  wire v1214ebc;
  wire v1214ebd;
  wire v1214ec0;
  wire v1214ec1;
  wire v1214ec2;
  wire v1214ec3;
  wire v1214ec4;
  wire v1214ec5;
  wire v1214ec6;
  wire v1214ec7;
  wire v1214ec8;
  wire v1214ec9;
  wire v1214eca;
  wire v1214ecb;
  wire v1214ecc;
  wire v1214ecd;
  wire v1214ece;
  wire v1214ecf;
  wire v1214ed0;
  wire v1214ed1;
  wire v1214ed2;
  wire v1214ed3;
  wire v1214ed4;
  wire v1214ed5;
  wire v1214ed6;
  wire v1214ed7;
  wire v1214ed8;
  wire v1214ed9;
  wire v1214eda;
  wire v1214edb;
  wire v1214edc;
  wire v1214edd;
  wire v1214ede;
  wire v1214edf;
  wire v1214ee0;
  wire v1214ee1;
  wire v1214ee2;
  wire v1214ee3;
  wire v1214ee4;
  wire v1214ee5;
  wire v1214ee6;
  wire v1214ee7;
  wire v1214ee8;
  wire v1214ee9;
  wire v1214eea;
  wire v1214eeb;
  wire v1214eec;
  wire v1214eed;
  wire v1214eee;
  wire v1214eef;
  wire v1214ef0;
  wire v1214ef1;
  wire v1214ef2;
  wire v1214ef3;
  wire v1214ef4;
  wire v1214ef5;
  wire v1214ef6;
  wire v1214ef7;
  wire v1214ef8;
  wire v1214ef9;
  wire v1214efa;
  wire v1214efb;
  wire v1214efc;
  wire v1214efd;
  wire v1214efe;
  wire v1214eff;
  wire v1214f00;
  wire v1214f01;
  wire v1214f02;
  wire v1214f03;
  wire v1214f04;
  wire v1214f05;
  wire v1214f06;
  wire v1214f07;
  wire v1214f08;
  wire v1214f09;
  wire v1214f0a;
  wire v1214f0b;
  wire v1214f0c;
  wire v1214f0d;
  wire v1214f0e;
  wire v1214f0f;
  wire v1214f10;
  wire v1214f11;
  wire v1214f12;
  wire v1214f13;
  wire v1214f14;
  wire v1214f15;
  wire v1214f16;
  wire v1214f17;
  wire v1214f18;
  wire v1214f19;
  wire v1214f1a;
  wire v1214f1b;
  wire v1214f38;
  wire v1214f39;
  wire v1214f3a;
  wire v1214f3b;
  wire v1214f3c;
  wire v1214f3d;
  wire v1214f4e;
  wire v1214f4f;
  wire v1214f50;
  wire v1214f51;
  wire v1214f53;
  wire v1214f54;
  wire v1214f55;
  wire v1214f56;
  wire v1214f57;
  wire v1214f58;
  wire v1214f59;
  wire v1214f5a;
  wire v1214f5b;
  wire v1214f5c;
  wire v1214f5d;
  wire v1214f5e;
  wire v1214f5f;
  wire v1214f60;
  wire v1214f61;
  wire v1214f62;
  wire v1214f63;
  wire v1214f64;
  wire v1214f65;
  wire v1214f66;
  wire v1214f67;
  wire v1214f68;
  wire v1214f69;
  wire v1214f6a;
  wire v1214f6b;
  wire v1214f6e;
  wire v1214f6f;
  wire v1214f70;
  wire v1214f71;
  wire v1214f7d;
  wire v1214f7e;
  wire v12147e5;
  wire v12147e6;
  wire v12147e7;
  wire v12147e8;
  wire v12147e9;
  wire v12147ea;
  wire v12147ed;
  wire v12147ee;
  wire v12147ef;
  wire v12147f0;
  wire v12147f1;
  wire v12147fd;
  wire v12147fe;
  wire v12147ff;
  wire v1214800;
  wire v1214815;
  wire v1214816;
  wire v1214817;
  wire v1214818;
  wire v1214819;
  wire v121481a;
  wire v121481b;
  wire v121482c;
  wire v121482d;
  wire v121482e;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hbusreq2_p;
  input hbusreq2;
  reg hlock2_p;
  input hlock2;
  reg hbusreq3_p;
  input hbusreq3;
  reg hlock3_p;
  input hlock3;
  reg hbusreq4_p;
  input hbusreq4;
  reg hlock4_p;
  input hlock4;
  reg hbusreq5_p;
  input hbusreq5;
  reg hlock5_p;
  input hlock5;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmaster1_p;
  output hmaster1;
  reg hmaster2_p;
  output hmaster2;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg hgrant2_p;
  output hgrant2;
  reg hgrant3_p;
  output hgrant3;
  reg hgrant4_p;
  output hgrant4;
  reg hgrant5_p;
  output hgrant5;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg stateG10_2_p;
  output stateG10_2;
  reg stateG10_3_p;
  output stateG10_3;
  reg stateG10_4_p;
  output stateG10_4;
  reg stateG10_5_p;
  output stateG10_5;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;
  reg jx2_p;
  output jx2;

assign v1445f9b = hbusreq1_p & v14463b7 | !hbusreq1_p & v14463bb;
assign v12ad681 = hbusreq5_p & v12ad51d | !hbusreq5_p & !v12ad680;
assign v134d50f = hmaster2_p & v134d50d | !hmaster2_p & v134d50e;
assign v1214dc4 = hbusreq2 & v1214dba | !hbusreq2 & v1214dc3;
assign v144649f = hgrant5_p & v845542 | !hgrant5_p & v144649e;
assign v13891a4 = hmaster0_p & v13891a3 | !hmaster0_p & v845542;
assign v12163a8 = hbusreq0 & v12163a6 | !hbusreq0 & v12163a7;
assign v134cdc2 = hmaster0_p & v134cd71 | !hmaster0_p & v845542;
assign v1214d32 = decide_p & v1214c27 | !decide_p & v1214d31;
assign v12ad549 = hmaster2_p & v12ad519 | !hmaster2_p & !v12ad51c;
assign v1446425 = hbusreq1 & v1446421 | !hbusreq1 & v1446424;
assign v1445e01 = hbusreq0 & v1445dff | !hbusreq0 & v1445e00;
assign v1552d5c = hgrant5_p & v1552d5b | !hgrant5_p & v1553391;
assign v1668c28 = hmaster2_p & v845542 | !hmaster2_p & !a66275;
assign v1445e97 = hbusreq0_p & v144639c | !hbusreq0_p & v1445e56;
assign v14465cf = hlock1 & v14465ce | !hlock1 & v14465cb;
assign v151574b = hgrant5_p & v151573d | !hgrant5_p & v151574a;
assign a658ed = hbusreq2_p & a658e7 | !hbusreq2_p & a658eb;
assign v12163a3 = hbusreq5_p & v12163a2 | !hbusreq5_p & v1216acf;
assign v1214ce6 = hmaster0_p & v1214c2e | !hmaster0_p & v1214c2c;
assign a6548f = hmaster0_p & a658e8 | !hmaster0_p & a658f1;
assign v138a3a5 = hbusreq2_p & v138a3a2 | !hbusreq2_p & v138a3a4;
assign a653e0 = hgrant1_p & a653c7 | !hgrant1_p & !a653df;
assign v1446655 = hbusreq5_p & v1446654 | !hbusreq5_p & v1446636;
assign d30154 = hbusreq5_p & d30153 | !hbusreq5_p & d30152;
assign d30827 = hgrant5_p & d306d0 | !hgrant5_p & d307dc;
assign v140585b = hmaster1_p & v140585a | !hmaster1_p & v140584d;
assign v16a1d6c = hbusreq0 & v16a207a | !hbusreq0 & v16a1d6b;
assign d2fb73 = hlock5_p & d2fb71 | !hlock5_p & d2fb72;
assign v15155e7 = hlock0_p & v1668c2d | !hlock0_p & v15155e6;
assign v1216218 = hgrant1_p & v845542 | !hgrant1_p & v1216217;
assign f2f35e = hmaster2_p & f2f295 | !hmaster2_p & v845542;
assign d80765 = decide_p & d80752 | !decide_p & d80764;
assign v121617a = hgrant5_p & v121600e | !hgrant5_p & v1216179;
assign v1446648 = hbusreq5_p & v1446647 | !hbusreq5_p & v1446643;
assign v1515773 = hgrant4_p & v151576f | !hgrant4_p & v1515772;
assign d2f9a1 = hbusreq1_p & d2fec0 | !hbusreq1_p & d2f9a0;
assign v134d3da = hgrant0_p & v845542 | !hgrant0_p & v134d3d9;
assign a65b32 = hgrant3_p & a65b28 | !hgrant3_p & a65b31;
assign d807bb = decide_p & d80751 | !decide_p & d807ba;
assign v134d4ba = decide_p & v134d3fa | !decide_p & v134d4b9;
assign v1216295 = hgrant2_p & v1216289 | !hgrant2_p & !v1216294;
assign v1445789 = hmaster2_p & v1445de5 | !hmaster2_p & v1445ec0;
assign v12152f4 = hbusreq2 & v12152f0 | !hbusreq2 & v12152f3;
assign d2f9a8 = hbusreq0 & d2f9a3 | !hbusreq0 & d2f9a7;
assign v1445871 = hbusreq1 & v144586d | !hbusreq1 & v1445870;
assign v10d40a5 = hmaster0_p & v10d3ffd | !hmaster0_p & v10d3ff1;
assign v1405b18 = hgrant0_p & v1405abf | !hgrant0_p & !v1405a87;
assign v16a1e08 = hgrant2_p & v845542 | !hgrant2_p & !v16a1e06;
assign v15156e5 = hmaster0_p & v15156e4 | !hmaster0_p & !v15156b0;
assign v12af3a4 = hbusreq1_p & v12afda1 | !hbusreq1_p & v12afda3;
assign v16a1aba = decide_p & v16a1f9e | !decide_p & v16a1ab9;
assign v1215779 = hbusreq5_p & v1215777 | !hbusreq5_p & !v1215778;
assign d80779 = hlock4_p & d80733 | !hlock4_p & !v845542;
assign v1445b14 = hlock2 & v1445af2 | !hlock2 & v1445b12;
assign v121655d = hlock4_p & v121655c | !hlock4_p & !v845542;
assign v1515604 = decide_p & v1515603 | !decide_p & v845576;
assign d2fb4a = hgrant3_p & d2f9d9 | !hgrant3_p & !d2fb49;
assign v1284d0b = hgrant4_p & v140587c | !hgrant4_p & v1284d0a;
assign v12161fe = hgrant2_p & v12161f9 | !hgrant2_p & v12161fd;
assign v134d21f = hmaster2_p & v134d1e8 | !hmaster2_p & v134d1f5;
assign d30655 = hgrant1_p & d30654 | !hgrant1_p & v845542;
assign v1446711 = hlock3 & v1446702 | !hlock3 & v1446710;
assign v12153f1 = hlock2_p & v12153ed | !hlock2_p & v12153f0;
assign d2f9cb = hmaster0_p & d2f9ca | !hmaster0_p & d2f994;
assign v144599a = hgrant4_p & v14458d2 | !hgrant4_p & v144639c;
assign v10d4032 = hgrant1_p & v10d402c | !hgrant1_p & !v10d4031;
assign a6627d = hbusreq5_p & a6627a | !hbusreq5_p & a6627c;
assign v16a1e68 = hmaster0_p & v16a1e63 | !hmaster0_p & v16a1e5f;
assign v1445522 = hbusreq2_p & v1445521 | !hbusreq2_p & v1445bdb;
assign d2fcaf = hbusreq1_p & d2fcae | !hbusreq1_p & !v845542;
assign v1214edb = hgrant5_p & v1214ed9 | !hgrant5_p & v1214eda;
assign v121606d = hmaster1_p & v121606c | !hmaster1_p & v121605d;
assign v1445ea3 = hlock1 & v1445e8d | !hlock1 & v1445ea2;
assign v155343e = hmaster2_p & v155343d | !hmaster2_p & v845542;
assign v16a1d16 = stateA1_p & v84557e | !stateA1_p & !v845582;
assign v1216556 = hlock0_p & v1216a61 | !hlock0_p & v845547;
assign v1214d10 = hgrant2_p & v1214d0a | !hgrant2_p & v1214d0f;
assign v12153e1 = hlock0_p & v12153d0 | !hlock0_p & v845547;
assign bf1f83 = hmaster2_p & bf1f80 | !hmaster2_p & bf1f82;
assign v1216040 = hmaster2_p & v121603d | !hmaster2_p & v121603f;
assign v1668c9b = hbusreq5_p & v1668c99 | !hbusreq5_p & v1668c9a;
assign d807a4 = decide_p & d80787 | !decide_p & d807a3;
assign d2fb05 = hmaster2_p & d306b0 | !hmaster2_p & d2fb04;
assign d2f98a = hbusreq1 & d2feb4 | !hbusreq1 & d2f989;
assign v1445785 = hmaster1_p & v1445784 | !hmaster1_p & v1445e1b;
assign v12152fc = hmaster1_p & v12152fb | !hmaster1_p & v1214fbf;
assign v134cdcc = decide_p & v134d3ce | !decide_p & v134cd8c;
assign d2fd29 = hbusreq2 & d2fd28 | !hbusreq2 & d302f3;
assign v10d4096 = hbusreq2_p & v10d408e | !hbusreq2_p & v10d4095;
assign v138a33d = hgrant4_p & v138a33c | !hgrant4_p & a658e0;
assign v1216ab2 = hlock5_p & v1216aae | !hlock5_p & !v1216ab1;
assign d300f4 = hgrant5_p & d300e4 | !hgrant5_p & d300f3;
assign bf1f8d = hgrant0_p & a6537d | !hgrant0_p & d2fc50;
assign v134ce3f = hgrant4_p & v134ce3e | !hgrant4_p & v845542;
assign v144600b = hready_p & v144639b | !hready_p & v144600a;
assign v1216118 = hmaster2_p & v1216100 | !hmaster2_p & v845542;
assign v134d239 = hbusreq3 & v134d21e | !hbusreq3 & v134d238;
assign v1214c6b = hlock4_p & v1214c6a | !hlock4_p & v845547;
assign v1445355 = hmaster0_p & v1445902 | !hmaster0_p & v1445a6b;
assign v140593d = decide_p & v1405918 | !decide_p & v1405902;
assign v1214dcf = hmaster0_p & v1216a68 | !hmaster0_p & v845542;
assign v1216299 = hgrant5_p & v121602d | !hgrant5_p & v1216132;
assign a6564b = hbusreq1_p & a653df | !hbusreq1_p & a6564a;
assign v121539c = hlock1_p & v121539a | !hlock1_p & v121539b;
assign v1284ced = hgrant5_p & v1284cca | !hgrant5_p & !v1284cec;
assign f2f416 = hmaster0_p & f2f2a4 | !hmaster0_p & f2f296;
assign v1445b48 = hmaster1_p & v1445b47 | !hmaster1_p & v1445a61;
assign v1214ff5 = hgrant4_p & v845542 | !hgrant4_p & v1215bac;
assign v1405aa9 = hbusreq5_p & v1405aa8 | !hbusreq5_p & v1405aa6;
assign v16a1dae = decide_p & v16a1dad | !decide_p & !v16a2065;
assign stateG3_0 = !v134cf70;
assign v1215d79 = hmaster0_p & v1215d75 | !hmaster0_p & v1215d78;
assign d307c0 = hmaster2_p & d307bf | !hmaster2_p & d30655;
assign v16a2237 = busreq_p & v16a2236 | !busreq_p & v845542;
assign v1446257 = hmaster1_p & v144621d | !hmaster1_p & v1446250;
assign v12ad5b3 = hgrant5_p & v12ad4f3 | !hgrant5_p & v12ad5b1;
assign v151577d = hlock0_p & a6588d | !hlock0_p & !v151577c;
assign v1215ba1 = hmaster0_p & v1215b9f | !hmaster0_p & v1215ba0;
assign v12161b5 = hbusreq5 & v121618b | !hbusreq5 & v12161b4;
assign v12aef0a = hready_p & v12af5c4 | !hready_p & v12aef09;
assign v134d4b3 = hlock2 & v134d4b0 | !hlock2 & v134d4b2;
assign v1515706 = hmaster1_p & v15156fb | !hmaster1_p & !v15156da;
assign v144662d = hbusreq5_p & v144662c | !hbusreq5_p & v1446611;
assign d3072e = hmaster2_p & d3071b | !hmaster2_p & v84554e;
assign v1446279 = hbusreq5_p & v1446411 | !hbusreq5_p & v1446278;
assign v134cd72 = hmaster0_p & v845542 | !hmaster0_p & v134cd71;
assign v1405b21 = hbusreq5_p & v1405b1d | !hbusreq5_p & v1405b20;
assign v1445b6a = hmaster1_p & v1446323 | !hmaster1_p & v1445b5f;
assign v134d386 = hgrant1_p & v845542 | !hgrant1_p & v134d385;
assign v1215bef = hbusreq1 & v121601c | !hbusreq1 & !v845542;
assign v144645f = hready_p & v144639b | !hready_p & v144645e;
assign v16a1442 = hmaster1_p & v16a1441 | !hmaster1_p & v16a209c;
assign v121538c = hmaster1_p & v121538b | !hmaster1_p & v1215388;
assign v1389df9 = hmaster0_p & v1389de7 | !hmaster0_p & v1389de1;
assign d2fc3a = hbusreq0 & d2fc36 | !hbusreq0 & d2fc39;
assign d80797 = hgrant0_p & d80796 | !hgrant0_p & !v845542;
assign v1214d9d = hmaster1_p & v1214d9c | !hmaster1_p & v1215388;
assign v12ad58c = hmaster1_p & v12ad531 | !hmaster1_p & v12ad54f;
assign v1405853 = stateG3_2_p & v845542 | !stateG3_2_p & v845584;
assign v12163ad = hbusreq2_p & v12163ac | !hbusreq2_p & v12163ab;
assign v12ad4c9 = hbusreq3_p & v12adbec | !hbusreq3_p & v12ad4c8;
assign v1668d8b = hmaster0_p & v1668d61 | !hmaster0_p & v1668d8a;
assign v1214c9d = hlock2_p & v1214c81 | !hlock2_p & v1214c9c;
assign v1668db3 = hgrant5_p & v1668da6 | !hgrant5_p & v1668d29;
assign v1216399 = hbusreq3 & v1216330 | !hbusreq3 & v845542;
assign v14457c5 = hbusreq2_p & v14457c3 | !hbusreq2_p & v14457c4;
assign d30246 = hbusreq5_p & d30244 | !hbusreq5_p & d30245;
assign v12ad601 = hbusreq5_p & v12ad5fe | !hbusreq5_p & !v12ad600;
assign d3012e = hbusreq2 & d30122 | !hbusreq2 & d3012d;
assign v1215b86 = hbusreq4_p & v1215b85 | !hbusreq4_p & v845542;
assign v144545c = hlock3 & v1445446 | !hlock3 & v144545a;
assign d2fc35 = hmaster2_p & d2fb78 | !hmaster2_p & d30690;
assign f2f3d5 = hgrant5_p & f2f2a8 | !hgrant5_p & !f2f3a4;
assign v1446722 = hbusreq5 & v144671e | !hbusreq5 & v1446721;
assign v1446600 = hgrant4_p & v1446423 | !hgrant4_p & v144639c;
assign d30706 = hmaster0_p & d306ff | !hmaster0_p & d30705;
assign v1214ca0 = hbusreq2_p & v1214c9e | !hbusreq2_p & v1214c9f;
assign v140588d = hmastlock_p & v146b550 | !hmastlock_p & v845542;
assign d300ba = hgrant0_p & a6537d | !hgrant0_p & d300b9;
assign a6549b = hmaster1_p & a658f1 | !hmaster1_p & a65476;
assign v1216a5b = hburst0_p & v134d1d9 | !hburst0_p & v845542;
assign v12ad27b = hgrant3_p & v12ad1ff | !hgrant3_p & v12ad27a;
assign v12161d8 = hbusreq1_p & v12161d7 | !hbusreq1_p & !v845542;
assign f2f38c = hbusreq1_p & f2f38b | !hbusreq1_p & v845542;
assign bf1fab = hbusreq3_p & bf1f8a | !hbusreq3_p & !bf1faa;
assign v1668d1e = hmaster0_p & v1668d1b | !hmaster0_p & v1668d1d;
assign v1284cc8 = hmaster2_p & v1284cc7 | !hmaster2_p & v14463b1;
assign v10d42b6 = hgrant2_p & v10d408a | !hgrant2_p & v10d42b5;
assign v1553232 = hlock0_p & v1553138 | !hlock0_p & v845542;
assign d30197 = hbusreq3 & d30192 | !hbusreq3 & d308f7;
assign v1405888 = hlock1_p & v140583d | !hlock1_p & v140583c;
assign v16a1388 = hbusreq2_p & v16a1a99 | !hbusreq2_p & v16a1387;
assign a656b8 = hgrant3_p & a654cb | !hgrant3_p & a656b6;
assign a662ca = hgrant1_p & v845542 | !hgrant1_p & !a662c7;
assign a662a4 = decide_p & a6627f | !decide_p & a662a2;
assign v1215729 = hgrant4_p & v845542 | !hgrant4_p & v1215728;
assign d2fbed = hgrant1_p & d2fbe8 | !hgrant1_p & d2fbec;
assign v138a3f0 = hbusreq2_p & v138a3e2 | !hbusreq2_p & v138a3ef;
assign v1214c0a = hbusreq2_p & v1214c09 | !hbusreq2_p & v1214c08;
assign v140583f = locked_p & v140583e | !locked_p & v14463b1;
assign v151573f = hbusreq1 & a653c8 | !hbusreq1 & !v151563e;
assign v144617e = hgrant2_p & v144617d | !hgrant2_p & v144616e;
assign v10d401f = hbusreq1_p & v10d3fdb | !hbusreq1_p & !v10d3fd8;
assign v1446133 = hlock3 & v1446127 | !hlock3 & v1446132;
assign v1284ce2 = hmaster2_p & v1284cc7 | !hmaster2_p & v1405844;
assign v14463c4 = hmaster2_p & v144639c | !hmaster2_p & v14463a2;
assign v16a206d = hgrant1_p & v84554d | !hgrant1_p & v16a206c;
assign v1445872 = hbusreq1_p & v144639c | !hbusreq1_p & v1445871;
assign v15161d5 = hbusreq2_p & v15161d4 | !hbusreq2_p & !v845542;
assign v144587e = hgrant5_p & v144587b | !hgrant5_p & !v144587d;
assign busreq = v16a144b;
assign v138a038 = hbusreq5 & v1389ff5 | !hbusreq5 & v138a037;
assign d2fe8a = hbusreq4_p & d2fe89 | !hbusreq4_p & v845542;
assign v1284cac = hlock2_p & v1284ca8 | !hlock2_p & v1284cab;
assign v1515643 = hbusreq2 & v1515642 | !hbusreq2 & !v845542;
assign v12150b3 = hready_p & v1215022 | !hready_p & v12150b2;
assign v1216110 = hbusreq1_p & v121610f | !hbusreq1_p & v845542;
assign v1445851 = hlock2 & v14457f6 | !hlock2 & v1445850;
assign v138a39f = hbusreq2_p & v138a39c | !hbusreq2_p & v138a39e;
assign v1215747 = hgrant1_p & v1215746 | !hgrant1_p & v121573b;
assign v121614b = hgrant0_p & v121614a | !hgrant0_p & v845542;
assign v1215bea = hmaster2_p & v1216021 | !hmaster2_p & v1216024;
assign v10d427f = hmastlock_p & v10d427e | !hmastlock_p & v10d3fd3;
assign v1284cd9 = hlock0_p & v1284c8f | !hlock0_p & !v14058aa;
assign v1668d2a = hgrant5_p & v1668d15 | !hgrant5_p & v1668d29;
assign v1405ab6 = hmaster1_p & v1405ab5 | !hmaster1_p & v1405aae;
assign a65b26 = hmaster1_p & v845542 | !hmaster1_p & a65b25;
assign v1445e9a = hbusreq4_p & v1445e99 | !hbusreq4_p & v144660d;
assign v134d263 = hlock2_p & v134d261 | !hlock2_p & v134d262;
assign v1446413 = hmaster2_p & v1446406 | !hmaster2_p & v1446412;
assign d30209 = hbusreq1_p & d30208 | !hbusreq1_p & d30207;
assign v12160f6 = hlock1_p & v12160f1 | !hlock1_p & v12160f5;
assign v1389f8b = hmaster2_p & v15168ad | !hmaster2_p & v845542;
assign v12ad5e5 = hbusreq0 & v12ad5e4 | !hbusreq0 & v845542;
assign v1216277 = hbusreq2_p & v1216274 | !hbusreq2_p & v1216276;
assign v1215362 = hmaster1_p & v1215361 | !hmaster1_p & v845542;
assign v16a1e4e = hgrant2_p & v16a1d32 | !hgrant2_p & v16a1e4d;
assign d30875 = hmaster0_p & d30874 | !hmaster0_p & d3086e;
assign v1214d3c = hmaster1_p & v1214d3b | !hmaster1_p & v1215388;
assign f2e4f2 = hbusreq2_p & f2f52e | !hbusreq2_p & f2ed94;
assign v15157cd = hgrant5_p & v845570 | !hgrant5_p & v15157cc;
assign d3027c = hlock5_p & d3027a | !hlock5_p & !d3027b;
assign v155314d = hmaster2_p & v1553148 | !hmaster2_p & v155314c;
assign v1215061 = hmaster2_p & v121545f | !hmaster2_p & !v1215060;
assign v12ad50e = stateG2_p & v845542 | !stateG2_p & !v9a051b;
assign v1445896 = hbusreq0 & v1445894 | !hbusreq0 & v1445895;
assign v1214d5f = hmaster0_p & v1214d5e | !hmaster0_p & v1214d4a;
assign v1215c48 = hgrant2_p & v1215c39 | !hgrant2_p & !v1215c47;
assign v151565b = hbusreq5_p & v1515659 | !hbusreq5_p & !v151565a;
assign v1216570 = hgrant1_p & v845542 | !hgrant1_p & v121656f;
assign v1445beb = hmaster0_p & v144643d | !hmaster0_p & v144639c;
assign d300f9 = hlock1_p & d300f7 | !hlock1_p & d300f8;
assign d2fd2b = hlock2_p & v845542 | !hlock2_p & d2fd2a;
assign v1405a9d = hbusreq2_p & v1405a9a | !hbusreq2_p & v1405a9c;
assign v138a449 = decide_p & v138a448 | !decide_p & v845542;
assign v144645b = hlock5 & v1446455 | !hlock5 & v144645a;
assign v12162c5 = hgrant2_p & v12162c3 | !hgrant2_p & v12162c4;
assign v1216024 = hlock0_p & v845547 | !hlock0_p & v1216023;
assign v1446447 = hbusreq0 & v1446446 | !hbusreq0 & v144643e;
assign v12ad505 = hbusreq2_p & v12ad500 | !hbusreq2_p & v12ad504;
assign d306a3 = hgrant0_p & v84554a | !hgrant0_p & v845548;
assign v134d23f = hlock2_p & v134d23d | !hlock2_p & v134d23e;
assign v16a1ab9 = hbusreq5 & v16a1ab8 | !hbusreq5 & v16a2064;
assign v1446343 = hgrant2_p & v14462e9 | !hgrant2_p & v1446342;
assign d307ec = hbusreq1_p & d307eb | !hbusreq1_p & v845542;
assign f2f331 = hmaster1_p & f2f2cc | !hmaster1_p & !f2f330;
assign v1668dbd = hgrant5_p & v845570 | !hgrant5_p & v1668d3d;
assign v134d4e3 = hbusreq2_p & v134d4de | !hbusreq2_p & v134d4e2;
assign v1668d60 = hbusreq5_p & v1668d5c | !hbusreq5_p & !v1668d5f;
assign v1214c81 = hmaster1_p & v1214c80 | !hmaster1_p & v845542;
assign a653e9 = hgrant2_p & a6535d | !hgrant2_p & a653e8;
assign v16693af = hbusreq3 & v16693a9 | !hbusreq3 & v16693ae;
assign v1405927 = hbusreq0_p & v140588e | !hbusreq0_p & v1405926;
assign v16a12e5 = hready_p & v845555 | !hready_p & !v16a12e4;
assign v12150d3 = hmaster1_p & v12153ee | !hmaster1_p & v12150d1;
assign v12153f8 = hbusreq2 & v12153f2 | !hbusreq2 & v12153f7;
assign v1214cea = hgrant0_p & v1214ce9 | !hgrant0_p & !v845542;
assign v10d4264 = stateG3_2_p & v845542 | !stateG3_2_p & !v88d3e4;
assign v14465e8 = hlock1 & v144641d | !hlock1 & v14465e7;
assign v16a2089 = hgrant4_p & v845559 | !hgrant4_p & !v845542;
assign v16a12c6 = hbusreq3 & v16a12c2 | !hbusreq3 & v16a12c5;
assign bf1fa0 = hgrant1_p & f2f227 | !hgrant1_p & bf1f9f;
assign v10d42cc = hbusreq5_p & v10d4273 | !hbusreq5_p & !v10d42cb;
assign v1445918 = hbusreq5_p & v14458e6 | !hbusreq5_p & v1445917;
assign v138a30c = hbusreq3 & v138a307 | !hbusreq3 & v138a30b;
assign f2f2d9 = hmaster2_p & f2f2d3 | !hmaster2_p & !f2f2d8;
assign v16a1cf7 = hbusreq5_p & v16a1be0 | !hbusreq5_p & v16a1cf6;
assign d30101 = hgrant5_p & d2fea1 | !hgrant5_p & d300ff;
assign v12160b8 = hbusreq2 & v12160b2 | !hbusreq2 & v12160b7;
assign v138a05b = hgrant3_p & v1389fce | !hgrant3_p & v138a05a;
assign f2f437 = hgrant5_p & f2f385 | !hgrant5_p & !f2f436;
assign v1284d65 = hgrant3_p & v1284d41 | !hgrant3_p & v1284d64;
assign v1445895 = hmaster2_p & v1445891 | !hmaster2_p & v14463bb;
assign f2f451 = hgrant5_p & v84554c | !hgrant5_p & f2f436;
assign v144614f = hlock2 & v1446125 | !hlock2 & v144614d;
assign v16a1aff = hmaster1_p & v16a1afe | !hmaster1_p & v16a2672;
assign v1445bdc = hbusreq2_p & v1445bd7 | !hbusreq2_p & v1445bdb;
assign v1214d0f = hmaster1_p & v1214d0e | !hmaster1_p & v1214d04;
assign a65446 = hmaster1_p & a65445 | !hmaster1_p & a65439;
assign v12ad514 = hbusreq0_p & v12ad513 | !hbusreq0_p & !v845542;
assign v144634d = hlock3 & v144632f | !hlock3 & v144634c;
assign v134d4db = hgrant5_p & v845542 | !hgrant5_p & v134d4da;
assign d30138 = hmaster2_p & d30124 | !hmaster2_p & d2fe80;
assign bf1f66 = hgrant4_p & v845570 | !hgrant4_p & a65382;
assign v14459b5 = hbusreq0_p & v14459b4 | !hbusreq0_p & v14465bb;
assign f2f3f9 = hmaster0_p & f2f2e8 | !hmaster0_p & f2f2cc;
assign v1214c1e = hbusreq2_p & v1214c1d | !hbusreq2_p & v1214c1c;
assign v1445b86 = hlock3 & v144632f | !hlock3 & v1445b85;
assign v15161fb = hlock2_p & v15161fa | !hlock2_p & !v845542;
assign v14454a4 = hlock5 & v144546f | !hlock5 & v144549f;
assign v16695c7 = hbusreq3_p & v16695c6 | !hbusreq3_p & !v1668c39;
assign v14058bd = hmaster1_p & v14058bc | !hmaster1_p & v14058b1;
assign v144611a = hmaster0_p & v1446079 | !hmaster0_p & v1445fe3;
assign v1215766 = hlock0_p & v1215b90 | !hlock0_p & !v845542;
assign v1668dad = hmaster1_p & v1668dac | !hmaster1_p & v845542;
assign v1215025 = hbusreq4 & v845542 | !hbusreq4 & v845547;
assign v1445fe7 = hbusreq1_p & v1446444 | !hbusreq1_p & v1446406;
assign d300d8 = hlock4_p & d307ac | !hlock4_p & !v845542;
assign f2f35a = hgrant5_p & f2f293 | !hgrant5_p & !f2f359;
assign v1446437 = hmaster1_p & v1446405 | !hmaster1_p & v1446436;
assign v14458b0 = hmaster1_p & v144639c | !hmaster1_p & v14458af;
assign v1515aee = hbusreq2 & v1515ae3 | !hbusreq2 & v1515aed;
assign v1445d93 = hbusreq5_p & v1445d8e | !hbusreq5_p & v1445d92;
assign v134d1e5 = hburst1_p & v134d1e4 | !hburst1_p & v845584;
assign d307be = hbusreq1_p & d307bd | !hbusreq1_p & v845542;
assign v134cebc = hlock3 & v134d270 | !hlock3 & v134cebb;
assign d30869 = hmaster2_p & d30867 | !hmaster2_p & d30868;
assign v12aec4e = hlock3_p & v12aec16 | !hlock3_p & v12aec4d;
assign v16a1e0c = hgrant2_p & v845542 | !hgrant2_p & v16a1e0a;
assign v1216538 = hgrant1_p & v1216522 | !hgrant1_p & v1216537;
assign a6538e = hbusreq5_p & a6538b | !hbusreq5_p & a6538d;
assign a6628c = hgrant5_p & v845542 | !hgrant5_p & a6628b;
assign a653cb = hlock0_p & a6585c | !hlock0_p & a653c9;
assign f2f350 = hbusreq1_p & f2f34f | !hbusreq1_p & v845542;
assign v1668d23 = hbusreq1_p & v1668d21 | !hbusreq1_p & v1668d22;
assign v1405b09 = hmaster0_p & v1405b01 | !hmaster0_p & !v1405b08;
assign d30954 = hmaster2_p & v845542 | !hmaster2_p & !d30952;
assign v16a1415 = hbusreq2 & v16a1414 | !hbusreq2 & v16a2060;
assign d300e4 = hmaster2_p & d300d8 | !hmaster2_p & d2fe9d;
assign v134d206 = hlock0_p & v134d1e8 | !hlock0_p & v845542;
assign v16a1d81 = hbusreq5 & v16a1d76 | !hbusreq5 & v16a1d80;
assign v16a20a4 = hbusreq2 & v16a20a2 | !hbusreq2 & !v16a20a3;
assign v144674c = hmaster1_p & v144674b | !hmaster1_p & v1446436;
assign v16a1beb = hgrant2_p & v845542 | !hgrant2_p & v16a1be9;
assign v1215d3e = hmaster1_p & v1215d3d | !hmaster1_p & v1215d2b;
assign v144602c = hbusreq2_p & v1446019 | !hbusreq2_p & v144602b;
assign v14458b9 = stateG10_5_p & v144588a | !stateG10_5_p & !v14458b8;
assign v1216119 = hgrant5_p & v1216117 | !hgrant5_p & v1216118;
assign v134d376 = hgrant5_p & v134d36a | !hgrant5_p & v134d375;
assign v1445e21 = hbusreq2 & v1445e1a | !hbusreq2 & v1445e20;
assign v1516219 = decide_p & v15167ee | !decide_p & !v845576;
assign v134cd65 = hbusreq1 & v134cd63 | !hbusreq1 & v134cd64;
assign v16a1d93 = hmaster1_p & v16a1d92 | !hmaster1_p & !v16a2672;
assign v12157a4 = hbusreq0 & v12157a2 | !hbusreq0 & v12157a3;
assign v1446192 = hlock2 & v144618c | !hlock2 & v1446191;
assign v1214d87 = hgrant2_p & v1214c9d | !hgrant2_p & v1214d82;
assign v11e5955 = hgrant1_p & v845542 | !hgrant1_p & !v11e5954;
assign a65854 = hburst1_p & v1553931 | !hburst1_p & a65853;
assign v134d4cc = hgrant1_p & v134d4cb | !hgrant1_p & v845542;
assign v15156be = hmaster1_p & v15156bd | !hmaster1_p & v151566b;
assign v12ad55f = hmaster1_p & v12ad544 | !hmaster1_p & v12ad54f;
assign a653dd = hgrant0_p & a653dc | !hgrant0_p & v845570;
assign v1215ca2 = hlock1_p & v1215ca1 | !hlock1_p & !v845542;
assign v143fd77 = hready_p & v845542 | !hready_p & v845566;
assign v121629d = hmaster1_p & v12161a1 | !hmaster1_p & v121629c;
assign v11e5975 = hgrant0_p & v845542 | !hgrant0_p & !v11e5974;
assign v1445369 = hbusreq2_p & v1445363 | !hbusreq2_p & v1445368;
assign v1214c4a = hgrant0_p & v845542 | !hgrant0_p & !v1214c49;
assign v12ad61c = hbusreq5_p & v12ad61a | !hbusreq5_p & !v12ad61b;
assign d308ce = hbusreq2 & d308ca | !hbusreq2 & d308cd;
assign v12165ae = hbusreq5_p & v12165ad | !hbusreq5_p & v845542;
assign d3028b = hgrant2_p & d3028a | !hgrant2_p & d30284;
assign v1445780 = hbusreq2_p & v144577a | !hbusreq2_p & v144577f;
assign v14463f4 = hbusreq5_p & v14463f3 | !hbusreq5_p & v14463c5;
assign v1215ffb = hmaster2_p & v1215ffa | !hmaster2_p & v845542;
assign v12157a1 = hgrant2_p & v121570b | !hgrant2_p & v12157a0;
assign v14058e4 = decide_p & v14058bf | !decide_p & v14058e3;
assign v1553099 = hmaster0_p & v1553098 | !hmaster0_p & v155305e;
assign v134d26e = hmaster1_p & v134d20a | !hmaster1_p & v134d23c;
assign v12afdb5 = hmaster1_p & v845542 | !hmaster1_p & v12afdb4;
assign v1446084 = hgrant2_p & v144607b | !hgrant2_p & v1446083;
assign v14460b2 = hgrant5_p & v14460af | !hgrant5_p & v14460b1;
assign d30291 = hlock5_p & d30290 | !hlock5_p & d30277;
assign v1446203 = decide_p & v1446117 | !decide_p & v1446202;
assign a6567b = hgrant2_p & a6561c | !hgrant2_p & a6567a;
assign v121508a = hgrant0_p & v121545e | !hgrant0_p & !v845559;
assign v1515737 = hmaster2_p & v151572a | !hmaster2_p & v845542;
assign v1215fe7 = hbusreq3_p & v121678f | !hbusreq3_p & v1215fe6;
assign v12ad591 = hbusreq3 & v12ad587 | !hbusreq3 & v12ad590;
assign v1284d3a = hbusreq4_p & v140588d | !hbusreq4_p & v1284d39;
assign v1216263 = hmaster0_p & v121625e | !hmaster0_p & v1216262;
assign v1445832 = hmaster1_p & v144580a | !hmaster1_p & v1445ef0;
assign v12ad540 = hmaster1_p & v12ad52d | !hmaster1_p & !v12ad525;
assign v121482c = jx2_p & v121481b | !jx2_p & v1215ddc;
assign v14466d9 = hmaster1_p & v14466d8 | !hmaster1_p & v14463ef;
assign v16a223f = hgrant5_p & v16a2234 | !hgrant5_p & v16a223e;
assign d30786 = hgrant4_p & d30783 | !hgrant4_p & d30785;
assign v11e597d = hmaster1_p & v11e597c | !hmaster1_p & !v11e595c;
assign d2fc7a = hbusreq2 & d2fc78 | !hbusreq2 & d2fc79;
assign v138a301 = hmaster0_p & v138a2fe | !hmaster0_p & v138a300;
assign v1552d92 = hmaster0_p & v845542 | !hmaster0_p & v1552d91;
assign v1389819 = hgrant2_p & v845542 | !hgrant2_p & !v1389818;
assign v1445e27 = hlock0 & v1445e26 | !hlock0 & v1445e25;
assign v144643f = hbusreq0 & v144643c | !hbusreq0 & v144643e;
assign v16a1d1a = hmaster2_p & v16a1d19 | !hmaster2_p & v845542;
assign v16a1b00 = hbusreq2 & v16a1afc | !hbusreq2 & v16a1aff;
assign v1445ec4 = hmaster0_p & v1446404 | !hmaster0_p & v1445ec3;
assign d301c6 = hmaster2_p & v845542 | !hmaster2_p & d301c5;
assign v134ce8a = hbusreq1 & v134d1ec | !hbusreq1 & v134ce89;
assign d30644 = hmastlock_p & v1553934 | !hmastlock_p & !v845542;
assign v14466d8 = hmaster0_p & v14463f6 | !hmaster0_p & v144639c;
assign v1389445 = hgrant1_p & v1389444 | !hgrant1_p & v15168ad;
assign v121545d = hlock3_p & v1215442 | !hlock3_p & v121545c;
assign v1668d33 = hbusreq5_p & v1668d31 | !hbusreq5_p & v1668d32;
assign d30161 = hbusreq2 & d3015d | !hbusreq2 & d30160;
assign f2f2cb = hbusreq1_p & f2f2ca | !hbusreq1_p & v845542;
assign v1445e74 = hgrant1_p & v1445df2 | !hgrant1_p & v1445e73;
assign v15157a8 = hbusreq1_p & v15157a7 | !hbusreq1_p & !v845542;
assign v1515710 = hbusreq1 & v1515609 | !hbusreq1 & v845570;
assign v1445bd5 = hmaster0_p & v1445bd4 | !hmaster0_p & v1446611;
assign v1214bcc = hlock5_p & v1214bca | !hlock5_p & v1214bcb;
assign v16a1981 = hgrant2_p & v845542 | !hgrant2_p & !v16a1980;
assign d2fad6 = hmaster1_p & d2fad5 | !hmaster1_p & !d2f97d;
assign v14466f3 = hmaster1_p & v14466f2 | !hmaster1_p & v1446436;
assign d30729 = hbusreq1_p & d30728 | !hbusreq1_p & v845542;
assign v1215722 = hmaster2_p & v1215717 | !hmaster2_p & v1215721;
assign v1216a84 = hlock3_p & v1216a7e | !hlock3_p & v1216a83;
assign v14458e1 = hbusreq0_p & v1446407 | !hbusreq0_p & v1446406;
assign v134d52b = decide_p & v134d3fa | !decide_p & v134d52a;
assign v12ad32c = hbusreq2_p & v12ae201 | !hbusreq2_p & v12ad32b;
assign v121657a = hmaster0_p & v845542 | !hmaster0_p & v1216a7a;
assign v1668d52 = hbusreq1 & a65861 | !hbusreq1 & v845542;
assign v14466aa = hmaster1_p & v14465b8 | !hmaster1_p & v14466a9;
assign v134d3af = hmaster1_p & v134d3ae | !hmaster1_p & v845542;
assign v14458de = hbusreq0_p & v14458dd | !hbusreq0_p & v1446406;
assign v1445f64 = hmaster1_p & v1445f63 | !hmaster1_p & v14466a9;
assign d30162 = hbusreq5 & d3012e | !hbusreq5 & d30161;
assign v14460cd = hbusreq0 & v14460cc | !hbusreq0 & v1446053;
assign v16a1dad = hbusreq5 & v16a1dac | !hbusreq5 & v16a1ad4;
assign v14466de = hbusreq2_p & v14466d9 | !hbusreq2_p & v14466dd;
assign v1445443 = hmaster0_p & v144621c | !hmaster0_p & v144639c;
assign v12afda2 = hmaster2_p & v845542 | !hmaster2_p & !v12afda1;
assign v134ce3b = hbusreq0 & v134ce3a | !hbusreq0 & v134d379;
assign v1668da1 = hbusreq0 & v1668d9c | !hbusreq0 & v1668da0;
assign v140587f = hmaster0_p & v140587d | !hmaster0_p & v140587e;
assign v1214ce1 = hmaster0_p & v1214cc1 | !hmaster0_p & v1214ce0;
assign v16a1f99 = hbusreq2 & v16a1f97 | !hbusreq2 & v16a1f98;
assign v12153eb = hbusreq0 & v12153e5 | !hbusreq0 & v12153ea;
assign a65619 = hgrant2_p & a65614 | !hgrant2_p & a65616;
assign v10d4026 = hgrant5_p & v10d3fdc | !hgrant5_p & v10d4025;
assign v134d1ea = hmastlock_p & v134d1e9 | !hmastlock_p & v845542;
assign v1552d6c = decide_p & v1553216 | !decide_p & v1552d6b;
assign v12167a6 = hmaster0_p & v1668c1f | !hmaster0_p & v12165a9;
assign v144621b = hbusreq0 & v14463c4 | !hbusreq0 & v144639c;
assign v1445f54 = hmaster0_p & v1446448 | !hmaster0_p & v1446657;
assign a65652 = hmaster0_p & a65640 | !hmaster0_p & a65650;
assign v12152fb = hmaster0_p & v1214fc4 | !hmaster0_p & v1214fb6;
assign v1215320 = hmaster0_p & v121505b | !hmaster0_p & v1215030;
assign v1215d63 = hmaster2_p & v12164cf | !hmaster2_p & v845542;
assign v14459da = hgrant4_p & v14459d6 | !hgrant4_p & v14459d9;
assign v1214dac = hmaster0_p & v1214c3c | !hmaster0_p & v1214d08;
assign v1215bd5 = hlock3_p & v121639a | !hlock3_p & !v1215bd4;
assign v1214dae = hmaster1_p & v1214d0d | !hmaster1_p & v1214d04;
assign v151580b = hgrant3_p & v151570e | !hgrant3_p & !v151580a;
assign v144647a = hmaster2_p & v845542 | !hmaster2_p & v1446479;
assign d300ce = hmaster2_p & d300cd | !hmaster2_p & d300c4;
assign v1216ae6 = hbusreq5_p & v1216ae5 | !hbusreq5_p & v845542;
assign v1553439 = hgrant0_p & v845542 | !hgrant0_p & v1553438;
assign v1553052 = hmaster2_p & v845542 | !hmaster2_p & v1553051;
assign f2e4f9 = hready_p & f2e4f4 | !hready_p & f2e4f8;
assign v1215316 = hmaster1_p & v1215315 | !hmaster1_p & v1215016;
assign v1445841 = hbusreq3 & v144583f | !hbusreq3 & v1445840;
assign v138a30d = hbusreq5 & v138a30c | !hbusreq5 & v845542;
assign v15167c3 = hbusreq2_p & v15167c2 | !hbusreq2_p & v845542;
assign d306ad = hbusreq5_p & d30653 | !hbusreq5_p & !d306ac;
assign v12afe45 = hgrant4_p & v845542 | !hgrant4_p & !v12afe44;
assign v1405933 = hbusreq2_p & v1405922 | !hbusreq2_p & v1405932;
assign v1214db9 = hgrant2_p & v1214dad | !hgrant2_p & v1214db8;
assign v138938c = hlock5_p & v138938b | !hlock5_p & v845542;
assign v134d4ea = hgrant1_p & v134d4e9 | !hgrant1_p & v845542;
assign v1445ad3 = hbusreq2_p & v1445acf | !hbusreq2_p & v1445ad2;
assign v1445be1 = decide_p & v1446224 | !decide_p & v1446275;
assign v14465c7 = hbusreq1_p & v144639c | !hbusreq1_p & v14465c6;
assign f2f297 = hmaster0_p & f2f296 | !hmaster0_p & f2f293;
assign v121632c = hlock2_p & v121632b | !hlock2_p & v121631d;
assign a662c5 = decide_p & a662c3 | !decide_p & v845542;
assign v1215335 = hgrant2_p & v1215329 | !hgrant2_p & v1215334;
assign a6567d = hgrant2_p & a6540a | !hgrant2_p & a65663;
assign v12166f2 = hmaster2_p & v12164cf | !hmaster2_p & !v12166ce;
assign d307f8 = hmaster0_p & d306fd | !hmaster0_p & d307f7;
assign v1668c44 = hmaster0_p & v1668c43 | !hmaster0_p & v1668c3f;
assign v15530a5 = hbusreq5 & v15530a3 | !hbusreq5 & v15530a4;
assign v14461dd = hlock3 & v144617b | !hlock3 & v14461db;
assign hgrant1 = !f2e506;
assign v144600f = hgrant5_p & v144600e | !hgrant5_p & v144647a;
assign v1215386 = hmaster2_p & v1215385 | !hmaster2_p & v845542;
assign a65665 = hgrant2_p & a65614 | !hgrant2_p & a65663;
assign v14458fb = hbusreq0 & v14458f9 | !hbusreq0 & v14458fa;
assign v12ad5ef = hgrant2_p & v12ad5e7 | !hgrant2_p & v12ad5ee;
assign d3060e = hmaster1_p & d3060d | !hmaster1_p & d30608;
assign v134cd79 = hlock3 & v134d3b5 | !hlock3 & v134cd78;
assign v14457d0 = hbusreq3 & v14457c2 | !hbusreq3 & v14457cf;
assign v134d441 = hmaster0_p & v845542 | !hmaster0_p & v134d440;
assign v14058b8 = hgrant5_p & v140584f | !hgrant5_p & v14058b7;
assign a65ada = hmaster1_p & a662cb | !hmaster1_p & a65ad7;
assign v16a2078 = hgrant5_p & v845542 | !hgrant5_p & v16a2077;
assign d306f4 = hbusreq1 & d306f3 | !hbusreq1 & !v845542;
assign v1515627 = locked_p & v1515626 | !locked_p & v845542;
assign d2fbd9 = hlock5_p & d2fbd7 | !hlock5_p & d2fbd8;
assign d30892 = hmaster2_p & d3088f | !hmaster2_p & d30891;
assign v15157a3 = hgrant5_p & v845542 | !hgrant5_p & !v15157a1;
assign d3067a = hbusreq5_p & v845542 | !hbusreq5_p & d30656;
assign a646da = hbusreq2_p & a65aff | !hbusreq2_p & a65b26;
assign v14058da = hgrant2_p & v1405884 | !hgrant2_p & v14058d9;
assign v134d4d6 = hlock0_p & v134d1dd | !hlock0_p & v134d4d5;
assign d30621 = hbusreq2_p & d30620 | !hbusreq2_p & d3061f;
assign v1215d0b = hbusreq3 & v1215d0a | !hbusreq3 & v845542;
assign v134d3d7 = decide_p & v134d3cf | !decide_p & v134d3d6;
assign f2f33b = hmaster1_p & f2f2e3 | !hmaster1_p & !f2f330;
assign v1214fc0 = hmaster1_p & v1214fb6 | !hmaster1_p & v1214fbf;
assign v1405b1e = hgrant1_p & v1405abf | !hgrant1_p & v1405b19;
assign v1214eb3 = hbusreq3 & v1214e7e | !hbusreq3 & v1214eb2;
assign v10d429b = hbusreq5_p & v10d4297 | !hbusreq5_p & !v10d429a;
assign v1216b07 = hbusreq2_p & v1216b06 | !hbusreq2_p & v1216afd;
assign v134d498 = hbusreq0 & v134d396 | !hbusreq0 & v134d388;
assign d2fea6 = hmaster1_p & d2fea5 | !hmaster1_p & !d2fea2;
assign v1215349 = hbusreq0 & v1215348 | !hbusreq0 & v845542;
assign f2f41c = hmaster1_p & f2f41b | !hmaster1_p & f2f39d;
assign v15155fa = hmaster2_p & v845570 | !hmaster2_p & !v15155f9;
assign v1553422 = hbusreq3 & v1553420 | !hbusreq3 & v1553421;
assign v12153d1 = hbusreq4 & v1216ab0 | !hbusreq4 & v845542;
assign v138a3e6 = hgrant5_p & v845570 | !hgrant5_p & !v1515833;
assign v12afe52 = hbusreq5_p & v12afe51 | !hbusreq5_p & v12afe47;
assign d3074d = hlock2_p & d3074c | !hlock2_p & d30748;
assign v1445a44 = hmaster0_p & v14459a3 | !hmaster0_p & v1445a43;
assign a65476 = hmaster0_p & a65471 | !hmaster0_p & !a65475;
assign v144622b = hmaster2_p & v14463b1 | !hmaster2_p & !v14463db;
assign v12162ec = hlock1_p & v12162eb | !hlock1_p & v845547;
assign v10d402a = hlock1_p & v10d3fd9 | !hlock1_p & v10d3fef;
assign d2fb91 = hlock2_p & d2fb8e | !hlock2_p & d2fb90;
assign a6591e = hmaster1_p & a658f2 | !hmaster1_p & !a65916;
assign v12ad619 = hgrant2_p & v12ad597 | !hgrant2_p & v12ad618;
assign v1515817 = hbusreq3 & v1515811 | !hbusreq3 & !v1515816;
assign v16693a6 = hbusreq4_p & a66275 | !hbusreq4_p & v84556a;
assign v1215c4c = hmaster1_p & v1215c4b | !hmaster1_p & v845542;
assign v134d46b = hgrant3_p & v134d468 | !hgrant3_p & v134d46a;
assign v16a1953 = hbusreq4_p & v16a1952 | !hbusreq4_p & v845542;
assign v1446155 = hmaster1_p & v1446139 | !hmaster1_p & v1445ffc;
assign v1215c9b = hgrant5_p & v1215c92 | !hgrant5_p & v1215c9a;
assign f2f4a7 = hbusreq1 & a66275 | !hbusreq1 & !v16693aa;
assign v121604f = hbusreq5_p & v121604e | !hbusreq5_p & v16a2243;
assign a658ce = hbusreq1_p & a658bf | !hbusreq1_p & !a658cc;
assign v121546b = hbusreq0_p & v12160f2 | !hbusreq0_p & v1215465;
assign v15532c5 = hgrant1_p & v845542 | !hgrant1_p & v15532c4;
assign v1214dc9 = hgrant3_p & v1214d73 | !hgrant3_p & v1214dc8;
assign v1445a49 = hbusreq1 & v14459b1 | !hbusreq1 & v1445a48;
assign v14459ff = hmaster2_p & v14459db | !hmaster2_p & v14459fc;
assign d2fe91 = hbusreq2_p & d2fe8d | !hbusreq2_p & d2fe90;
assign v1446703 = hmaster0_p & v1446657 | !hmaster0_p & v1446404;
assign v1668c9f = hmaster2_p & a658ca | !hmaster2_p & !v1668c77;
assign v1216103 = hgrant5_p & v121601e | !hgrant5_p & !v1216101;
assign d302d8 = hbusreq5_p & d305fe | !hbusreq5_p & d30691;
assign v1668cf6 = hbusreq2 & v1668cec | !hbusreq2 & v1668cf5;
assign v134d3c7 = hbusreq2_p & v134d263 | !hbusreq2_p & v134d3c6;
assign v12af22a = hgrant2_p & v12af73f | !hgrant2_p & v12af229;
assign d301cc = hlock2_p & d301c2 | !hlock2_p & !d301cb;
assign v1284d45 = hmaster0_p & v1284ce3 | !hmaster0_p & v1284cc9;
assign v16a1c9b = hgrant5_p & v845568 | !hgrant5_p & v16a1c9a;
assign v1552f75 = hlock2 & v155341e | !hlock2 & v1552f6b;
assign d30686 = hbusreq5 & d30685 | !hbusreq5 & !v845542;
assign d2fc4c = hbusreq4_p & d2fbd0 | !hbusreq4_p & d2fc4b;
assign v144539e = hbusreq2_p & v1445392 | !hbusreq2_p & v144539d;
assign a65925 = hmaster1_p & a6590b | !hmaster1_p & !a65916;
assign v1284cdf = hmaster0_p & v1284cd4 | !hmaster0_p & !v1284cde;
assign v138a454 = hmaster1_p & v138a453 | !hmaster1_p & v138a341;
assign v1515789 = hburst1_p & v1553931 | !hburst1_p & v1515788;
assign v1446057 = hbusreq1_p & v1446056 | !hbusreq1_p & v1446427;
assign v134d30a = hgrant1_p & v134d1dd | !hgrant1_p & v845542;
assign v140586e = hmaster2_p & v140586c | !hmaster2_p & v140586d;
assign v1515674 = hburst0 & v151566f | !hburst0 & v1515673;
assign v1389e33 = hgrant2_p & v845542 | !hgrant2_p & !v1389e32;
assign v10d42c4 = hlock0_p & v10d4267 | !hlock0_p & v10d42c3;
assign v12162d3 = hmaster1_p & v12162c9 | !hmaster1_p & !v121624b;
assign v1445510 = hlock3 & v1445501 | !hlock3 & v144550f;
assign v1515c7d = hmastlock_p & v1515c7c | !hmastlock_p & v845542;
assign v1445dcb = hmaster2_p & v1445db5 | !hmaster2_p & v1445d85;
assign d2fcfd = hbusreq5_p & d2fcfc | !hbusreq5_p & d2fcb1;
assign v1553229 = hmaster2_p & v845542 | !hmaster2_p & v1553228;
assign v1446678 = hmaster2_p & v144639c | !hmaster2_p & v1446677;
assign v14465f9 = hgrant0_p & v14465f7 | !hgrant0_p & !v14465f8;
assign v1389fbd = hlock5_p & v1389fbc | !hlock5_p & v845542;
assign v14461b0 = hmaster1_p & v1446166 | !hmaster1_p & v1445ffc;
assign v144610d = hmaster1_p & v1445fa9 | !hmaster1_p & v1445fbd;
assign v16a1da9 = hmaster1_p & v16a1ad0 | !hmaster1_p & !v16a2672;
assign v1405b04 = hgrant0_p & v1405a88 | !hgrant0_p & !v1405a92;
assign v12ad57a = hlock2_p & v12ad578 | !hlock2_p & v12ad579;
assign d307b2 = hgrant0_p & d307b1 | !hgrant0_p & d306d4;
assign f2eda1 = hready_p & f2eda0 | !hready_p & f2ed9c;
assign v14459dd = hlock1 & v14459cb | !hlock1 & v14459c2;
assign f2f336 = hbusreq2_p & f2f334 | !hbusreq2_p & f2f335;
assign v14458f2 = hbusreq4 & v14458f1 | !hbusreq4 & v14458dc;
assign v1446744 = hlock2 & v144673f | !hlock2 & v1446743;
assign v1214fbd = hgrant5_p & v845542 | !hgrant5_p & v1214fbc;
assign d308d2 = hgrant3_p & d3087c | !hgrant3_p & !d308d1;
assign v134d458 = hbusreq3 & v134d456 | !hbusreq3 & v134d457;
assign d30108 = hmaster2_p & d30662 | !hmaster2_p & d30107;
assign v16a1d9e = hbusreq5 & v16a1d97 | !hbusreq5 & v16a1d9d;
assign v144580f = hmaster1_p & v144580e | !hmaster1_p & v1445e07;
assign v10d4050 = hmaster1_p & v10d4028 | !hmaster1_p & !v10d404f;
assign v13895a1 = hbusreq5_p & v13895a0 | !hbusreq5_p & v845542;
assign v1216048 = hready & v1216047 | !hready & !v845542;
assign a65b2e = hbusreq2_p & a65b29 | !hbusreq2_p & a65b2c;
assign v1445ae8 = hmaster1_p & v1445ae7 | !hmaster1_p & v14458fd;
assign f2e4ca = hmaster0_p & f2f21d | !hmaster0_p & v845542;
assign v15168a8 = hbusreq2_p & v15168a7 | !hbusreq2_p & v845542;
assign d302e3 = hbusreq5_p & d302e2 | !hbusreq5_p & d30663;
assign d2faf8 = hgrant5_p & d2faf2 | !hgrant5_p & d2faf7;
assign v12acfde = hmaster1_p & v12acfbc | !hmaster1_p & v12ad54f;
assign v12aeb73 = hmaster1_p & v845542 | !hmaster1_p & v12aeb72;
assign v1216b12 = hbusreq2_p & v1216b11 | !hbusreq2_p & v1216b10;
assign v1405b30 = hgrant2_p & v1405b11 | !hgrant2_p & v1405b2f;
assign v1214bc6 = hlock2_p & v1214bc3 | !hlock2_p & v1214bc5;
assign v12157aa = hready & v845542 | !hready & v12157a9;
assign v12153b8 = hmaster2_p & v12153b4 | !hmaster2_p & v12153b7;
assign a658e8 = hmaster2_p & a658b0 | !hmaster2_p & !a658c7;
assign v1214bfe = hmaster0_p & v12153ab | !hmaster0_p & v12153b1;
assign v16a1dfe = hbusreq3 & v16a1d2f | !hbusreq3 & v16a1dfd;
assign v1446122 = hmaster1_p & v1446121 | !hmaster1_p & v1445fef;
assign v138a34c = hmaster0_p & v138a32d | !hmaster0_p & v138a34b;
assign d30127 = hmaster1_p & d30126 | !hmaster1_p & d2fe97;
assign v1215cc1 = hgrant1_p & v1215cb9 | !hgrant1_p & v121615d;
assign v10d3ff9 = hlock0_p & v10d3fd8 | !hlock0_p & v10d3ff8;
assign v121576d = hgrant5_p & v1215ba0 | !hgrant5_p & v121576b;
assign v16a1cfc = hgrant2_p & v845542 | !hgrant2_p & v16a1cf9;
assign a653c7 = hbusreq1_p & a653c2 | !hbusreq1_p & a653c6;
assign bf1f57 = hready_p & bf1f51 | !hready_p & bf1f56;
assign v14466c7 = hready_p & v14465a9 | !hready_p & v14466c6;
assign v1214cf6 = hmaster2_p & v1214cbc | !hmaster2_p & v1214cf5;
assign v12adf65 = hmaster1_p & v845542 | !hmaster1_p & v12adf64;
assign d3089a = hmaster2_p & d30891 | !hmaster2_p & d306aa;
assign v1552d91 = hmaster2_p & v845542 | !hmaster2_p & v1552d7c;
assign v14461e5 = hmaster1_p & v144616d | !hmaster1_p & v14460cf;
assign v10d42b1 = hgrant4_p & v10d3fd4 | !hgrant4_p & v10d42b0;
assign v10d3fe9 = hmaster0_p & v10d3fe4 | !hmaster0_p & v10d3fe8;
assign v84557a = hgrant4_p & v845542 | !hgrant4_p & !v845542;
assign v138a3f9 = hmaster1_p & v138a3f8 | !hmaster1_p & v845542;
assign v134cf6e = jx2_p & v134cf42 | !jx2_p & v134cf6d;
assign v121508b = hbusreq4_p & v121508a | !hbusreq4_p & v1216714;
assign v16a1a79 = hmaster2_p & v16a1a78 | !hmaster2_p & v16a206f;
assign v1216596 = hgrant1_p & v1216595 | !hgrant1_p & v1216a93;
assign v1553222 = hgrant1_p & v845542 | !hgrant1_p & v1553221;
assign v1215c23 = hbusreq0 & v1215c18 | !hbusreq0 & v1215c22;
assign v1446145 = hbusreq2_p & v1446141 | !hbusreq2_p & v1446144;
assign a65429 = hgrant5_p & a6541f | !hgrant5_p & a653b9;
assign v1445f49 = hmaster0_p & v1445db8 | !hmaster0_p & v1445da9;
assign v1405b4d = hbusreq1_p & v1405ad5 | !hbusreq1_p & v1405b4c;
assign v12162c0 = hmaster1_p & v12162bf | !hmaster1_p & v1216224;
assign v14463fb = hbusreq2_p & v14463f0 | !hbusreq2_p & v14463fa;
assign v1445dd1 = hmaster0_p & v1445dd0 | !hmaster0_p & v1445da3;
assign v144583c = hbusreq2_p & v1445830 | !hbusreq2_p & v144583b;
assign v1515830 = decide_p & v151582f | !decide_p & v845542;
assign v1284d23 = hgrant5_p & v1284cbc | !hgrant5_p & v1284d22;
assign v121501a = hmaster0_p & v12153b5 | !hmaster0_p & v1215019;
assign a654cb = hready_p & a65464 | !hready_p & a654c9;
assign v1445a73 = hbusreq3 & v1445a71 | !hbusreq3 & v1445a72;
assign v1214fca = hbusreq5 & v121578b | !hbusreq5 & v1214fc9;
assign v12acfc4 = hbusreq0 & v12acfc3 | !hbusreq0 & !v12af7f7;
assign v10d4292 = hgrant0_p & v10d3fe0 | !hgrant0_p & v10d4291;
assign v1284cc1 = hready_p & v1284c97 | !hready_p & !v1284cc0;
assign v1515744 = hbusreq4 & v151560d | !hbusreq4 & v845570;
assign d308a4 = hbusreq5_p & d307df | !hbusreq5_p & d308a3;
assign v16a169e = hbusreq0 & v16a1e92 | !hbusreq0 & v16a169d;
assign v1668cdc = hburst0 & v156645f | !hburst0 & v1668cdb;
assign v15161cb = hmaster0_p & v845570 | !hmaster0_p & v1668c17;
assign d306fc = hlock1_p & v845580 | !hlock1_p & v845542;
assign v1405aa4 = hlock1_p & v1405a87 | !hlock1_p & !v845542;
assign v1445b56 = hmaster2_p & v144665b | !hmaster2_p & v14465d2;
assign v1216144 = hbusreq0_p & v1216523 | !hbusreq0_p & v121611e;
assign d306c5 = hready_p & d306c4 | !hready_p & d306a1;
assign v1668d13 = decide_p & v1668d12 | !decide_p & !v845542;
assign d3020f = hbusreq5_p & d3020e | !hbusreq5_p & d3020d;
assign v16a1ac1 = hmaster1_p & v16a1ac0 | !hmaster1_p & !v16a2672;
assign v1445519 = hbusreq2_p & v1445518 | !hbusreq2_p & v1445bdb;
assign d2fd0e = hbusreq5 & d2fcf4 | !hbusreq5 & d2fd0d;
assign d30711 = hbusreq3 & d3070b | !hbusreq3 & !d30710;
assign v12ad5bf = hlock0_p & v1515745 | !hlock0_p & v845542;
assign d2fc73 = hbusreq5_p & d2fc0e | !hbusreq5_p & d2fc63;
assign v1668c18 = hbusreq5_p & v1668c17 | !hbusreq5_p & v845570;
assign v10d400f = hmaster0_p & v10d400a | !hmaster0_p & v10d400e;
assign v16a1cd0 = hbusreq5_p & v16a1afd | !hbusreq5_p & v16a1ccf;
assign v16a1e89 = decide_p & v16a1e7a | !decide_p & !v16a1e03;
assign f2ec20 = hbusreq1 & v16693a6 | !hbusreq1 & !v16693ab;
assign v1216095 = hlock5_p & v121607e | !hlock5_p & v1216094;
assign v1553146 = hbusreq5_p & v1553145 | !hbusreq5_p & v1553144;
assign v1216006 = hbusreq0_p & v1216a5a | !hbusreq0_p & v845570;
assign v1446730 = hmaster1_p & v144672f | !hmaster1_p & v1446436;
assign d2faf1 = hbusreq0 & d2fae5 | !hbusreq0 & d2faf0;
assign v134d540 = hgrant3_p & v134d53c | !hgrant3_p & v134d53f;
assign d2f9d7 = hbusreq5 & d2f9bd | !hbusreq5 & d2f9d6;
assign d301f5 = hmaster2_p & d301f4 | !hmaster2_p & d301ec;
assign v1389d5a = hbusreq5_p & v1389d59 | !hbusreq5_p & !v845542;
assign v845570 = locked_p & v845542 | !locked_p & !v845542;
assign v134cd6b = hmaster0_p & v134cd5e | !hmaster0_p & v134cd6a;
assign v138a35e = hmaster1_p & v138a34b | !hmaster1_p & v138a341;
assign v16a1379 = hmaster1_p & v16a1333 | !hmaster1_p & v16a1f96;
assign v1405875 = hbusreq2_p & v1405874 | !hbusreq2_p & v1405873;
assign v16a1372 = hbusreq2 & v16a1335 | !hbusreq2 & v16a1337;
assign v156645f = stateG3_2_p & v845542 | !stateG3_2_p & !v906a5a;
assign d8077f = hgrant4_p & v845542 | !hgrant4_p & !d8077e;
assign f2ec27 = hready_p & v845542 | !hready_p & f2ec26;
assign v1216318 = hmaster2_p & v1216aea | !hmaster2_p & v12162ed;
assign d2fd4d = jx2_p & d2fd4c | !jx2_p & d302f7;
assign f2e276 = hbusreq1_p & f2e275 | !hbusreq1_p & !v845542;
assign v1445eb2 = hmaster1_p & v1445eb1 | !hmaster1_p & v1445e07;
assign v14461ba = hgrant2_p & v14461b8 | !hgrant2_p & v14461b9;
assign v1284d26 = hgrant2_p & v1284d08 | !hgrant2_p & v1284d25;
assign v1216168 = hbusreq1_p & v1216167 | !hbusreq1_p & v845542;
assign v14461cd = hbusreq2_p & v14461c4 | !hbusreq2_p & v14461cc;
assign v1389d73 = hbusreq5_p & v1389d72 | !hbusreq5_p & v845542;
assign a658f2 = hmaster0_p & a658b7 | !hmaster0_p & a658f1;
assign a65ae9 = hbusreq5_p & a662cd | !hbusreq5_p & a65ae8;
assign v1214cc5 = locked_p & v1214cc4 | !locked_p & v845542;
assign f2e4d6 = hgrant3_p & f2e4cd | !hgrant3_p & f2e4d5;
assign v12acfbc = hmaster0_p & v12ad528 | !hmaster0_p & v12ad52d;
assign v1214f01 = hgrant5_p & v845542 | !hgrant5_p & v1214ecf;
assign v12afe70 = hmaster0_p & v12afe47 | !hmaster0_p & v12afe6f;
assign v1446315 = hgrant2_p & v1446309 | !hgrant2_p & v1446314;
assign v16a1410 = hbusreq2_p & v16a140f | !hbusreq2_p & v16a205b;
assign d30133 = hgrant5_p & d2fe80 | !hgrant5_p & d300ce;
assign v1445a9b = hmaster0_p & v1445a9a | !hmaster0_p & v1445a31;
assign d30637 = hbusreq2_p & d30636 | !hbusreq2_p & d30635;
assign v1215cfc = hgrant2_p & v1215c85 | !hgrant2_p & v1215cfb;
assign v1552fcb = hmaster0_p & v1552f6f | !hmaster0_p & v845542;
assign v1284ca7 = hmaster0_p & v1284ca2 | !hmaster0_p & v1284ca6;
assign v151563d = hbusreq2 & v151563c | !hbusreq2 & v845542;
assign v16a1e8b = hgrant0_p & v845542 | !hgrant0_p & v16a1e5b;
assign v138a3d2 = hmaster2_p & v845542 | !hmaster2_p & v1515757;
assign v144585c = hgrant2_p & v144583a | !hgrant2_p & v1445858;
assign v1668cc2 = hburst1 & v156645f | !hburst1 & v1668cc1;
assign v144537c = hmaster1_p & v1445b36 | !hmaster1_p & v144591b;
assign v1515849 = hmaster0_p & v1515848 | !hmaster0_p & v15157e4;
assign d3063c = hbusreq2 & d30637 | !hbusreq2 & d3063b;
assign f2f234 = hgrant1_p & f2f233 | !hgrant1_p & !v845542;
assign v1446065 = hmaster2_p & v1446062 | !hmaster2_p & v1446064;
assign v144640b = hlock4 & v1446407 | !hlock4 & v1446406;
assign v1515851 = decide_p & v151582f | !decide_p & !v845576;
assign v12166d4 = hgrant5_p & v845542 | !hgrant5_p & v12166d3;
assign d2feb8 = hbusreq1 & d2feb4 | !hbusreq1 & d2feb7;
assign d3084a = hbusreq1_p & d306fc | !hbusreq1_p & v845542;
assign v1215047 = hgrant1_p & v121546d | !hgrant1_p & v1215046;
assign v1446095 = hgrant2_p & v144608c | !hgrant2_p & v1446094;
assign v1446070 = hgrant5_p & v1445fdc | !hgrant5_p & v144606f;
assign v1215c0f = hgrant5_p & v1215c07 | !hgrant5_p & v1215c0e;
assign v1445848 = hmaster1_p & v14457e4 | !hmaster1_p & v1445f09;
assign v134d3ca = hbusreq2 & v134d3c5 | !hbusreq2 & v134d3c9;
assign v12166cc = hmastlock_p & v12166cb | !hmastlock_p & v845542;
assign v1284d1f = hmaster0_p & v1284d17 | !hmaster0_p & v1284d1e;
assign d30221 = hmaster2_p & d301d1 | !hmaster2_p & d301f4;
assign v10d40be = hbusreq4_p & v10d401c | !hbusreq4_p & v10d40bd;
assign v155305f = hmaster0_p & v1553054 | !hmaster0_p & v155305e;
assign v16a188f = hbusreq3 & v16a188b | !hbusreq3 & v16a188e;
assign v1216b01 = hmaster2_p & v845542 | !hmaster2_p & v1216acd;
assign v12ad58d = hlock2_p & v12ad58b | !hlock2_p & v12ad58c;
assign v10d4099 = hgrant3_p & v10d4013 | !hgrant3_p & v10d4098;
assign v12166e0 = hgrant5_p & v845542 | !hgrant5_p & v12166df;
assign v1445f6e = hlock2 & v144673f | !hlock2 & v1445f6c;
assign v16a1385 = hbusreq2_p & v16a1a95 | !hbusreq2_p & v16a1384;
assign v14838bd = decide_p & v14838b7 | !decide_p & v14838bc;
assign v16a1c97 = hbusreq1 & v16a223c | !hbusreq1 & v845542;
assign v1405af6 = hmaster2_p & v1405ad6 | !hmaster2_p & v1405a87;
assign a6587a = hmaster1_p & a65879 | !hmaster1_p & a6586e;
assign v1215d6b = hmaster2_p & v12166c5 | !hmaster2_p & v845542;
assign v1389808 = hgrant5_p & a6587e | !hgrant5_p & !v845542;
assign a6549a = hmaster1_p & a65499 | !hmaster1_p & a65476;
assign v134ce87 = hbusreq2_p & v134ce86 | !hbusreq2_p & v134d23e;
assign v1446224 = hmaster1_p & v144639c | !hmaster1_p & v1446223;
assign v121510b = hbusreq5 & v12150e3 | !hbusreq5 & v121510a;
assign v1552d84 = hbusreq4_p & v1553138 | !hbusreq4_p & v1552d7c;
assign v1284c8f = locked_p & v1284c8e | !locked_p & !v14463b1;
assign v1445760 = hlock2 & v1445759 | !hlock2 & v144575f;
assign v12ad52c = hmaster2_p & v12ad514 | !hmaster2_p & v12ad519;
assign v12ae1f2 = hmaster2_p & v12afe46 | !hmaster2_p & v12ae1f1;
assign v1215017 = hmaster1_p & v1214fed | !hmaster1_p & v1215016;
assign v1215b92 = hbusreq4_p & v1215b91 | !hbusreq4_p & v845542;
assign v14457a3 = hmaster0_p & v144579d | !hmaster0_p & v1445e0c;
assign v1445f00 = hbusreq2 & v1445efb | !hbusreq2 & v1445eff;
assign v1668c2f = hbusreq5_p & v1668c2e | !hbusreq5_p & v845568;
assign v1389fce = hready_p & v845542 | !hready_p & v1389fcd;
assign v1216191 = hlock5_p & v1216190 | !hlock5_p & v121611a;
assign d2fecb = hlock2_p & d2fec7 | !hlock2_p & d2feca;
assign v144547d = hbusreq0 & v1446678 | !hbusreq0 & v144639c;
assign v1215c60 = hbusreq5_p & v1215c5e | !hbusreq5_p & v1215c5f;
assign f2f3b6 = hbusreq2_p & f2f3af | !hbusreq2_p & !f2f3b5;
assign a67ea5 = hburst0_p & v845542 | !hburst0_p & v893df7;
assign v138a486 = hbusreq2_p & v138a482 | !hbusreq2_p & !v138a485;
assign v845550 = hbusreq2_p & v845542 | !hbusreq2_p & !v845542;
assign v1668c2e = hmaster2_p & v845542 | !hmaster2_p & v1668c2d;
assign v14453e1 = hmaster0_p & v144639c | !hmaster0_p & v14463c5;
assign v1214c43 = hmaster1_p & v1214c42 | !hmaster1_p & v1215357;
assign v144584e = hlock2 & v1445847 | !hlock2 & v144584d;
assign d3064a = hgrant1_p & f2f227 | !hgrant1_p & d30649;
assign f2f22e = hlock1_p & f2f22d | !hlock1_p & !v845542;
assign v16a16a7 = hgrant5_p & v845542 | !hgrant5_p & !v16a1e98;
assign d30214 = hgrant5_p & d301c9 | !hgrant5_p & d30212;
assign a65368 = hburst0 & a65366 | !hburst0 & a65367;
assign v1515756 = hbusreq1_p & v151572c | !hbusreq1_p & v1515755;
assign d308a9 = hmaster2_p & d308a6 | !hmaster2_p & d308a8;
assign v1216aa1 = decide_p & v1216a84 | !decide_p & v1216aa0;
assign v15168ad = hmastlock_p & v15168ac | !hmastlock_p & v845542;
assign v14465ee = hgrant0_p & v144641b | !hgrant0_p & v14463e1;
assign v11ac67b = hready_p & v84554c | !hready_p & v11ac67a;
assign v1216533 = hbusreq5_p & v1216532 | !hbusreq5_p & v845542;
assign v15156f5 = hmaster0_p & v15156f4 | !hmaster0_p & v1515675;
assign v144627a = hbusreq0 & v1446279 | !hbusreq0 & v1446265;
assign v1445ff1 = hmaster0_p & v144639c | !hmaster0_p & v1445fe1;
assign v1405acb = hmaster0_p & v1405abc | !hmaster0_p & v1405aca;
assign v1445b35 = hgrant2_p & v1445b32 | !hgrant2_p & v1445b34;
assign v1553933 = stateG3_2_p & v845542 | !stateG3_2_p & v1553932;
assign v1552d65 = hlock2 & v1552d62 | !hlock2 & v1552d64;
assign v1515728 = hgrant0_p & a6537d | !hgrant0_p & v1515720;
assign d3083e = hgrant2_p & d307f9 | !hgrant2_p & !d3083d;
assign v1553517 = hready_p & v1553427 | !hready_p & v1553516;
assign v121625f = hmaster1_p & v121625e | !hmaster1_p & !v121624b;
assign v138a090 = decide_p & v138a074 | !decide_p & v138a406;
assign v1215ba6 = hbusreq2_p & v1215ba2 | !hbusreq2_p & v1215ba5;
assign v12afe59 = hlock0_p & d305de | !hlock0_p & v845542;
assign v134ce85 = hmaster1_p & v134ce84 | !hmaster1_p & v134d23c;
assign v134d20e = hbusreq2_p & v134d20d | !hbusreq2_p & v134d20c;
assign v144553c = hgrant3_p & v14454a8 | !hgrant3_p & v144553b;
assign a6629a = hmaster2_p & a66299 | !hmaster2_p & a66286;
assign v16695a5 = hready_p & v166959d | !hready_p & !v16695a4;
assign v14460ab = hbusreq2 & v1446097 | !hbusreq2 & v14460aa;
assign v12165a1 = hgrant1_p & v1216a98 | !hgrant1_p & v12165a0;
assign v1284ccb = hlock1_p & v1284c8f | !hlock1_p & !v1405854;
assign v12afe4f = hgrant1_p & v845542 | !hgrant1_p & v12afe4e;
assign v16a1323 = hlock0_p & v16a1320 | !hlock0_p & v16a1322;
assign d308e7 = hmaster1_p & v845542 | !hmaster1_p & d308e6;
assign v16a1ccb = hmaster2_p & v16a1cca | !hmaster2_p & v845542;
assign v1215c37 = hgrant2_p & v1215bed | !hgrant2_p & v1215c36;
assign v1552d54 = hmaster1_p & v1552d53 | !hmaster1_p & v845542;
assign v11e5961 = hgrant1_p & v11e593a | !hgrant1_p & !v845542;
assign f2f327 = hmaster1_p & f2f2e3 | !hmaster1_p & f2f2db;
assign v1445431 = hlock3 & v144541f | !hlock3 & v1445430;
assign v15167b7 = hmaster1_p & v15167b6 | !hmaster1_p & v845542;
assign v134d217 = hbusreq0 & v134d216 | !hbusreq0 & v134d1e8;
assign v12ad564 = hmaster2_p & v12ad514 | !hmaster2_p & !a658d4;
assign v1445bf1 = hgrant2_p & v1445bec | !hgrant2_p & v1445bf0;
assign v12af9ce = hbusreq5_p & v12afe51 | !hbusreq5_p & v12af9c2;
assign v1214fc7 = hgrant2_p & v1215786 | !hgrant2_p & v1214fc6;
assign v1215730 = hbusreq0 & v1215725 | !hbusreq0 & v121572f;
assign a658e1 = hbusreq4_p & a658e0 | !hbusreq4_p & !v845542;
assign a65494 = hmaster1_p & a65493 | !hmaster1_p & a65476;
assign v138945b = hready_p & v845542 | !hready_p & v138945a;
assign v1405941 = jx2_p & v85e755 | !jx2_p & v1405940;
assign v1405ae4 = hbusreq5_p & v1405ae0 | !hbusreq5_p & v1405ae3;
assign v138a2fc = hmaster2_p & v845542 | !hmaster2_p & v151560e;
assign v1216575 = hmaster0_p & v121654f | !hmaster0_p & v1216574;
assign v144540a = hbusreq2_p & v1445409 | !hbusreq2_p & v1445bc8;
assign v1668ddb = hgrant5_p & v845542 | !hgrant5_p & !v1668d9d;
assign a656ca = hgrant5_p & v845542 | !hgrant5_p & a656c9;
assign v16a1d8e = hgrant2_p & v16a2058 | !hgrant2_p & v16a1d8d;
assign v1215bfe = hgrant5_p & v1215bfc | !hgrant5_p & v1215bfd;
assign v1445779 = hmaster0_p & v1445778 | !hmaster0_p & v1445de7;
assign v12165a8 = hmaster2_p & v845570 | !hmaster2_p & !v1216594;
assign v1445ad8 = hmaster1_p & v1445ac4 | !hmaster1_p & v14458c1;
assign v16a1bbb = hgrant4_p & v845559 | !hgrant4_p & v16a1bba;
assign v12ad8e9 = hmaster2_p & d30690 | !hmaster2_p & v12ad8e8;
assign v1215cb6 = hgrant5_p & v845542 | !hgrant5_p & !v1215cb5;
assign v121608a = hbusreq2_p & v1216089 | !hbusreq2_p & v1216088;
assign v16a141d = hready_p & v16a1409 | !hready_p & v16a141c;
assign v1215347 = hlock0_p & v1216a61 | !hlock0_p & v1215346;
assign v16a13df = hmaster0_p & v16a13db | !hmaster0_p & v16a13de;
assign v16a1cda = hbusreq2 & v16a1cd7 | !hbusreq2 & v16a1cd9;
assign v1552f5d = hbusreq0_p & v1553217 | !hbusreq0_p & v1552f53;
assign v15168b4 = hlock2_p & v15168b3 | !hlock2_p & v845542;
assign v14461fc = hlock2 & v144617b | !hlock2 & v14461fb;
assign v1446626 = hgrant0_p & v1446625 | !hgrant0_p & !v144661b;
assign v121574e = hgrant5_p & v1215740 | !hgrant5_p & v121574c;
assign a66286 = hgrant1_p & v845542 | !hgrant1_p & !a66285;
assign v1214d50 = hbusreq5_p & v1214bb7 | !hbusreq5_p & v1214d4f;
assign v16a19d4 = hmaster1_p & v16a19d3 | !hmaster1_p & v16a2672;
assign d3069d = hmaster0_p & d3069b | !hmaster0_p & d3069c;
assign v1552f57 = hbusreq1_p & v1553217 | !hbusreq1_p & v1552f56;
assign v14460f2 = hbusreq2_p & v14460f0 | !hbusreq2_p & v14460f1;
assign v1445b1c = hlock2 & v1445af2 | !hlock2 & v1445b1a;
assign v16a1be1 = hgrant5_p & v845542 | !hgrant5_p & !v16a1bcc;
assign f2f53b = hmaster1_p & f2f53a | !hmaster1_p & f2f52c;
assign a656c3 = decide_p & a656c2 | !decide_p & a662a2;
assign v12af9bf = hgrant4_p & d3068f | !hgrant4_p & !v12af9be;
assign v1445775 = hmaster2_p & v1445de5 | !hmaster2_p & v1445e70;
assign v12ae1f6 = hlock0_p & v1515ae5 | !hlock0_p & v845542;
assign v16a19ae = hgrant2_p & v16a2058 | !hgrant2_p & v16a19ad;
assign v1214e50 = hbusreq2 & v1214e42 | !hbusreq2 & v845542;
assign v1446476 = locked_p & v1446475 | !locked_p & v845542;
assign v1215c95 = hmaster2_p & v1215c87 | !hmaster2_p & v1215c94;
assign v16a1d7b = hmaster0_p & v16a1d78 | !hmaster0_p & v16a1d7a;
assign v845580 = stateA1_p & v845542 | !stateA1_p & !v845542;
assign v12160ea = hlock2_p & v12160e9 | !hlock2_p & !v1216028;
assign d30919 = hmaster1_p & d3090e | !hmaster1_p & d30918;
assign v1215fc0 = hbusreq2_p & v1215fbf | !hbusreq2_p & v1215fb9;
assign v14058c1 = hgrant4_p & v140583d | !hgrant4_p & v14058c0;
assign d2fe7a = hlock4_p & d306c8 | !hlock4_p & v845570;
assign v14466cb = decide_p & v14466ca | !decide_p & v144639b;
assign v14458c1 = hmaster0_p & v14458c0 | !hmaster0_p & v144589e;
assign v1445a80 = hbusreq0 & v1445a79 | !hbusreq0 & v1445a7f;
assign f2f3a3 = hbusreq5_p & f2f3a0 | !hbusreq5_p & f2f3a2;
assign v10d4079 = hgrant1_p & v10d3fe7 | !hgrant1_p & v10d4078;
assign v138a32d = hbusreq5_p & v138a32c | !hbusreq5_p & !v845542;
assign v144607b = hmaster1_p & v144607a | !hmaster1_p & v1445fde;
assign v15157c6 = hgrant4_p & v15157bb | !hgrant4_p & a65382;
assign v1216260 = hgrant2_p & v1216234 | !hgrant2_p & v121625f;
assign d807ae = hmaster2_p & d80760 | !hmaster2_p & !d8078a;
assign v134d4e8 = hbusreq1 & v134d4e6 | !hbusreq1 & v134d4e7;
assign v1215c09 = hlock1_p & v1215c08 | !hlock1_p & v845547;
assign v1216032 = hlock3_p & v121601b | !hlock3_p & !v1216031;
assign v1446042 = hgrant5_p & v1446040 | !hgrant5_p & v1446041;
assign a662c2 = hmaster0_p & v845542 | !hmaster0_p & !a662c1;
assign v121619c = hmaster0_p & v1216198 | !hmaster0_p & v121619b;
assign v121534a = hbusreq0_p & v1216a5a | !hbusreq0_p & v845542;
assign v16a132d = hgrant5_p & v845542 | !hgrant5_p & v16a132c;
assign v1215c73 = hmaster1_p & v1215c72 | !hmaster1_p & v1215c6a;
assign v1216afe = hlock2_p & v1216af9 | !hlock2_p & v1216afd;
assign v15157f3 = hgrant5_p & v845542 | !hgrant5_p & !v1515775;
assign v1445b92 = hbusreq2_p & v1445b8f | !hbusreq2_p & v1445b91;
assign v1668cd4 = hmaster2_p & v1668cd0 | !hmaster2_p & !v1668cd3;
assign v144667e = hbusreq0 & v144667d | !hbusreq0 & v1446638;
assign v1668c3f = hbusreq1_p & v845570 | !hbusreq1_p & v845542;
assign v134d4d7 = hgrant0_p & v134d4d6 | !hgrant0_p & v845542;
assign v12162f5 = hmaster1_p & v12162ea | !hmaster1_p & v12162f4;
assign v12ad5ed = hmaster0_p & v12ad5b5 | !hmaster0_p & v12ad5ec;
assign v12160b4 = hmaster1_p & v12160b3 | !hmaster1_p & v121605d;
assign v1216083 = hmaster1_p & v121604c | !hmaster1_p & v1216082;
assign f2f3e0 = hbusreq2 & f2f3dc | !hbusreq2 & f2f3df;
assign v14457ac = hlock3 & v1445786 | !hlock3 & v14457ab;
assign v144616f = hgrant2_p & v144616c | !hgrant2_p & v144616e;
assign v12162b9 = hmaster1_p & v12161fb | !hmaster1_p & v12161f4;
assign v16a1cfd = hbusreq2_p & v16a1beb | !hbusreq2_p & v16a1cfc;
assign v1214fe2 = hmaster1_p & v1214fe1 | !hmaster1_p & v12153bf;
assign v1214ed2 = hbusreq5_p & v1214ed0 | !hbusreq5_p & v1214ed1;
assign v1214d35 = hmaster0_p & v845547 | !hmaster0_p & v1215365;
assign v1552f67 = hbusreq0 & v1552f66 | !hbusreq0 & v15533a7;
assign v1445fc3 = hlock2 & v1445fc0 | !hlock2 & v1445fc2;
assign a6470f = hbusreq2 & a6470e | !hbusreq2 & a65b2e;
assign v1389465 = hbusreq5 & v138945d | !hbusreq5 & v1389464;
assign v12162e0 = decide_p & v12160ce | !decide_p & v12162df;
assign v1215bad = hbusreq4 & v1216a8d | !hbusreq4 & v845542;
assign f2f2a4 = hmaster2_p & f2f293 | !hmaster2_p & f2f29a;
assign a6543c = hgrant2_p & a6535d | !hgrant2_p & a6543a;
assign v1284cb1 = hmaster0_p & v1284ca9 | !hmaster0_p & v1284c98;
assign v12ad56f = hmaster1_p & v12ad56e | !hmaster1_p & !v12ad525;
assign v1216138 = hbusreq4_p & v121652c | !hbusreq4_p & v1216122;
assign v16a1333 = hmaster0_p & v16a132e | !hmaster0_p & v16a1329;
assign v1553446 = hready_p & v1553444 | !hready_p & v1553445;
assign v16a19a9 = hgrant4_p & v16a19a5 | !hgrant4_p & v16a19a8;
assign v16a13c1 = hlock2_p & v16a13ba | !hlock2_p & !v16a13c0;
assign v12acfca = hmaster1_p & v12acfc9 | !hmaster1_p & !v12ad525;
assign v1668cde = hbusreq1 & v1668cbd | !hbusreq1 & !v1668cdd;
assign v1216a7a = hbusreq5_p & v1216a79 | !hbusreq5_p & v845542;
assign v12afdac = hlock0_p & d305f0 | !hlock0_p & v845542;
assign v121504d = hgrant0_p & v121504c | !hgrant0_p & v845542;
assign v1284cb8 = hlock3_p & v1284cb0 | !hlock3_p & v1284cb7;
assign f2f377 = hbusreq5_p & f2f371 | !hbusreq5_p & !f2f376;
assign d30763 = hbusreq2_p & d30762 | !hbusreq2_p & d3075e;
assign a6566d = hbusreq5_p & a65422 | !hbusreq5_p & !a6566c;
assign v15168ab = hburst1 & v15168a9 | !hburst1 & v15168aa;
assign v138a32c = hmaster2_p & v138a32b | !hmaster2_p & !a658b5;
assign v1445fcd = hmaster2_p & v1445fcc | !hmaster2_p & v1446412;
assign v1215055 = hmaster1_p & v1215030 | !hmaster1_p & v1215054;
assign v1445d8b = stateG10_5_p & v1445d8a | !stateG10_5_p & !v1445d89;
assign v1214c33 = hmaster2_p & v1214c30 | !hmaster2_p & v1214c31;
assign v1215718 = hbusreq1 & v1215b7d | !hbusreq1 & v845542;
assign v14460e4 = hmaster0_p & v144601a | !hmaster0_p & v845542;
assign d3061f = hmaster1_p & d3061e | !hmaster1_p & d30608;
assign v12160a3 = hmaster1_p & v121605f | !hmaster1_p & v121605d;
assign v121678c = hbusreq5 & v1216713 | !hbusreq5 & v121678b;
assign v12162be = hmaster1_p & v12162bd | !hmaster1_p & v12160e0;
assign v12af3ab = hmaster0_p & v845542 | !hmaster0_p & v12af3aa;
assign v1445a3c = hgrant5_p & v14458ff | !hgrant5_p & v1445a3b;
assign f2f3e3 = decide_p & f2f340 | !decide_p & f2f23c;
assign v1389f93 = hmaster0_p & v1389f92 | !hmaster0_p & v845542;
assign v138a3c2 = hready_p & v138a320 | !hready_p & !v138a3c1;
assign v1445ddf = hlock5 & v1445dca | !hlock5 & v1445dde;
assign v1215371 = hmaster0_p & v1215370 | !hmaster0_p & v845542;
assign v138a35d = hbusreq2_p & v138a35a | !hbusreq2_p & v138a35c;
assign v121533d = hbusreq2_p & v121533a | !hbusreq2_p & v121533c;
assign v1445ef4 = hmaster1_p & v1445ebb | !hmaster1_p & v1445ef0;
assign v1214c79 = hgrant5_p & v845547 | !hgrant5_p & v1214c77;
assign d2fad5 = hmaster0_p & d2f974 | !hmaster0_p & d2f970;
assign v16a16b2 = decide_p & v16a1e7a | !decide_p & !v16a1e56;
assign v138a320 = decide_p & v138a31f | !decide_p & v845542;
assign v134d281 = hmaster2_p & v134d1dd | !hmaster2_p & v845542;
assign v1214f69 = hbusreq2_p & v1214f68 | !hbusreq2_p & v845542;
assign v16a2242 = hgrant2_p & v16a2058 | !hgrant2_p & v16a2241;
assign d308da = hlock1_p & d308d9 | !hlock1_p & v845542;
assign v1668d68 = stateG3_2_p & v88d3e4 | !stateG3_2_p & v1668d67;
assign a658f9 = hbusreq2 & a658ed | !hbusreq2 & a658f6;
assign d308ab = hbusreq5_p & d307f1 | !hbusreq5_p & d308aa;
assign v16a1b01 = hmaster0_p & v16a1afd | !hmaster0_p & v16a1afb;
assign v16a1d20 = hmaster1_p & v16a1d1f | !hmaster1_p & v16a2672;
assign f2f37c = hbusreq1 & v1668d7b | !hbusreq1 & v845542;
assign d807bd = decide_p & d80751 | !decide_p & d807b2;
assign v1445e57 = hbusreq4_p & v1445e56 | !hbusreq4_p & v14465bb;
assign v1515701 = hmaster1_p & v15156f2 | !hmaster1_p & !v15156da;
assign v1515813 = hmaster1_p & v1515812 | !hmaster1_p & v845542;
assign v1668cca = stateG3_2_p & v845542 | !stateG3_2_p & !v92fc87;
assign d3095b = hmaster1_p & d3090c | !hmaster1_p & d3095a;
assign v16a1a92 = hbusreq0_p & v16a2668 | !hbusreq0_p & v845542;
assign f2f226 = hlock1_p & v845570 | !hlock1_p & !v845542;
assign v12ad4e5 = hbusreq0_p & v1515630 | !hbusreq0_p & v845542;
assign d301ff = hmaster2_p & d301fe | !hmaster2_p & d301f9;
assign v12153ec = hmaster0_p & v12153e0 | !hmaster0_p & v12153eb;
assign d30283 = hmaster0_p & d30279 | !hmaster0_p & d30282;
assign v1214d1f = hmaster1_p & v1214cef | !hmaster1_p & !v1214d1e;
assign d3095a = hmaster0_p & d30956 | !hmaster0_p & d30959;
assign v16a1426 = hbusreq2_p & v16a13d4 | !hbusreq2_p & !v16a1ad1;
assign v138a348 = hmaster2_p & v138a32b | !hmaster2_p & v138a32f;
assign v1552d8b = hgrant1_p & v845542 | !hgrant1_p & v1552d8a;
assign v16a1dd7 = hmaster1_p & v845568 | !hmaster1_p & !v16a1f96;
assign v10d3fd3 = stateA1_p & v84557e | !stateA1_p & !v845542;
assign v1215c5d = hgrant5_p & v16a2243 | !hgrant5_p & v1215c0e;
assign v10d4017 = hmaster1_p & v10d4016 | !hmaster1_p & v10d3ffb;
assign v138a341 = hmaster0_p & v138a33a | !hmaster0_p & !v138a340;
assign v12acff3 = hmaster0_p & v12ad5ec | !hmaster0_p & v12ad5b5;
assign v12ad589 = hmaster1_p & v12ad574 | !hmaster1_p & v12ad54f;
assign v12aeb78 = hmaster1_p & v845542 | !hmaster1_p & v12aeb77;
assign a653b5 = hmaster2_p & a653b4 | !hmaster2_p & a653a3;
assign a6566b = hbusreq0 & a65667 | !hbusreq0 & a6566a;
assign d301fb = hgrant5_p & d301bd | !hgrant5_p & d301fa;
assign v1668d92 = hbusreq5_p & v1668d90 | !hbusreq5_p & !v1668d91;
assign d807b7 = hmaster1_p & d807b6 | !hmaster1_p & v845542;
assign v1389fbf = hmaster0_p & v1389fbe | !hmaster0_p & v845542;
assign v151571f = hmastlock_p & v151571e | !hmastlock_p & v10d3fd3;
assign d2fbdb = hbusreq0 & d2fbda | !hbusreq0 & v845542;
assign v1215ced = hmaster2_p & v1216014 | !hmaster2_p & v845542;
assign v1668d7e = hgrant5_p & v1668d1d | !hgrant5_p & v1668d7d;
assign d2fe83 = hlock4_p & d306d4 | !hlock4_p & v845570;
assign v121544f = hlock2_p & v121544d | !hlock2_p & v121544e;
assign v1668d01 = hmaster0_p & v1668d00 | !hmaster0_p & !v1668ce5;
assign d2fb3e = hbusreq2_p & d2fefb | !hbusreq2_p & d2fb3d;
assign v1214d8a = hbusreq2 & v1214d86 | !hbusreq2 & v1214d89;
assign v1515633 = hmaster1_p & v1515632 | !hmaster1_p & v845570;
assign v1215c7a = hbusreq3 & v1215c79 | !hbusreq3 & v845542;
assign d307d3 = hbusreq4_p & d307d2 | !hbusreq4_p & d307d1;
assign v14458a8 = hmaster1_p & v14458a7 | !hmaster1_p & v144589f;
assign a65682 = decide_p & a65681 | !decide_p & a662a2;
assign f2f32f = hbusreq5_p & f2f32d | !hbusreq5_p & f2f32e;
assign v10d3fe2 = hmaster2_p & v10d3fdb | !hmaster2_p & v10d3fe1;
assign f2f406 = hbusreq2_p & f2f404 | !hbusreq2_p & f2f405;
assign d30958 = hmaster2_p & a66278 | !hmaster2_p & !d30957;
assign v16a1d2b = hlock3_p & v16a1d12 | !hlock3_p & v16a1d2a;
assign d80792 = hbusreq4_p & d80733 | !hbusreq4_p & !d8078a;
assign v1668db0 = hbusreq2 & v1668da5 | !hbusreq2 & v1668daf;
assign v1552fd4 = hready_p & v1553427 | !hready_p & v1552fd3;
assign v1216211 = hbusreq1_p & v1216210 | !hbusreq1_p & v845542;
assign v12ad65c = hmaster1_p & v12ad635 | !hmaster1_p & v12ad65b;
assign v1216200 = decide_p & v12161b5 | !decide_p & v12161ff;
assign v1515798 = hgrant5_p & v845542 | !hgrant5_p & !v1515796;
assign v16a1d29 = hbusreq3 & v16a1d28 | !hbusreq3 & !v16a1f9c;
assign v1445f4f = hlock2 & v1445f40 | !hlock2 & v1445f4d;
assign v1215062 = hmaster0_p & v1215463 | !hmaster0_p & v1215061;
assign v12162de = hbusreq3 & v12162d6 | !hbusreq3 & v12162dd;
assign v12161ef = hbusreq1 & v12165a0 | !hbusreq1 & v845542;
assign v1445412 = hgrant1_p & v14465ae | !hgrant1_p & v144639c;
assign v1445f6a = hmaster1_p & v1445f69 | !hmaster1_p & v14466a9;
assign v12ad570 = hbusreq2_p & v12ad56d | !hbusreq2_p & v12ad56f;
assign v14459f1 = hbusreq0 & v14459e3 | !hbusreq0 & v14459f0;
assign v1553154 = hbusreq2_p & v1553153 | !hbusreq2_p & v1553152;
assign v14453ad = hlock2 & v14453a9 | !hlock2 & v14453ac;
assign d2fc0c = hmaster2_p & d2fc03 | !hmaster2_p & d2fb4d;
assign v14462f0 = hmaster2_p & v1446645 | !hmaster2_p & v14465e1;
assign v1515799 = hbusreq5_p & v1515797 | !hbusreq5_p & !v1515798;
assign v14458e7 = hlock1 & v14458e2 | !hlock1 & v14458db;
assign v1445da5 = hmaster1_p & v144639c | !hmaster1_p & v1445da4;
assign v12147ed = hmaster0_p & v1215d80 | !hmaster0_p & v1215d6c;
assign d30298 = hgrant2_p & d3028a | !hgrant2_p & d30294;
assign v1214c72 = hbusreq5_p & v1214c70 | !hbusreq5_p & v1214c71;
assign v14461eb = hlock2 & v144617b | !hlock2 & v14461ea;
assign v1446563 = hmaster1_p & v1446466 | !hmaster1_p & v1446562;
assign v1445b24 = hlock2 & v1445b21 | !hlock2 & v1445b23;
assign v1215c10 = hgrant5_p & v1215be7 | !hgrant5_p & v1215c0e;
assign v1405af3 = hmaster2_p & v1405a86 | !hmaster2_p & d3070c;
assign v1284d01 = hmaster0_p & v1405856 | !hmaster0_p & v1284d00;
assign f2ed92 = hmaster0_p & f2f236 | !hmaster0_p & f2f22b;
assign d80736 = hmaster1_p & d80735 | !hmaster1_p & v845542;
assign v16a129d = hmaster0_p & v16a1a97 | !hmaster0_p & v16a1a94;
assign v16a1cc4 = hbusreq2 & v16a1cc1 | !hbusreq2 & v16a1cc3;
assign v121610f = hlock1_p & v121610c | !hlock1_p & v121610e;
assign v1668dd0 = hbusreq5_p & v1668dce | !hbusreq5_p & !v1668dcf;
assign v1215d73 = hmaster2_p & v12166c5 | !hmaster2_p & v12166d2;
assign v1515642 = hlock2_p & v1515641 | !hlock2_p & v845542;
assign v1214d21 = hmaster1_p & v1214d0e | !hmaster1_p & !v1214d1e;
assign v10d4087 = hbusreq2_p & v10d407e | !hbusreq2_p & v10d4086;
assign v14462f1 = stateG10_5_p & v14465e2 | !stateG10_5_p & v14462f0;
assign d30202 = hbusreq0 & d301f7 | !hbusreq0 & d30201;
assign v1216ad1 = hbusreq5_p & v1216ad0 | !hbusreq5_p & v845542;
assign v1216a70 = hbusreq5_p & v1216a6f | !hbusreq5_p & v845542;
assign d2fe9b = hmaster2_p & d2fe9a | !hmaster2_p & !v84555a;
assign v10d4082 = hmaster2_p & v10d405f | !hmaster2_p & v10d406d;
assign v1215fbe = hmaster1_p & v1215fbd | !hmaster1_p & v12166ef;
assign v1214d25 = hbusreq2_p & v1214d24 | !hbusreq2_p & v1214d22;
assign v134d4a2 = hmaster1_p & v134d4a1 | !hmaster1_p & v845542;
assign f2f424 = hmaster2_p & f2f422 | !hmaster2_p & f2f423;
assign v1216560 = hgrant4_p & v845542 | !hgrant4_p & v1216a67;
assign v1216af4 = hmaster2_p & v1216adf | !hmaster2_p & !v1216af3;
assign v155323a = hgrant2_p & v155321f | !hgrant2_p & v1553239;
assign v1668c51 = hbusreq3 & v1668c4c | !hbusreq3 & v1668c50;
assign v134d4f6 = hbusreq5_p & v134d4f3 | !hbusreq5_p & v134d4f5;
assign f2f3eb = hmaster0_p & f2f3b2 | !hmaster0_p & v84554c;
assign d307c7 = hbusreq4_p & d307c5 | !hbusreq4_p & d307c6;
assign v1553152 = hmaster1_p & v1553151 | !hmaster1_p & v155314e;
assign v1445ded = hlock1 & v1445dec | !hlock1 & v1445dea;
assign v14465be = hbusreq4 & v14465bc | !hbusreq4 & v14465bd;
assign v12ad025 = hbusreq5_p & v12ad61a | !hbusreq5_p & !v12ad024;
assign d300c8 = hlock5_p & d300c6 | !hlock5_p & !d300c7;
assign v144590c = hbusreq2_p & v14458fe | !hbusreq2_p & v144590b;
assign v1445a98 = hbusreq0 & v1445a97 | !hbusreq0 & v14459f0;
assign v12150b4 = hgrant3_p & v1215476 | !hgrant3_p & v12150b3;
assign v12161ac = hbusreq5_p & v12161aa | !hbusreq5_p & v12161ab;
assign v1405b69 = jx0_p & v1405942 | !jx0_p & !v1405b68;
assign v1214c02 = hlock2_p & v1214bff | !hlock2_p & v1214c01;
assign v1284d58 = hgrant2_p & v1284d56 | !hgrant2_p & v1284d57;
assign v1445820 = hmaster1_p & v14457dd | !hmaster1_p & v1445e28;
assign v1214eec = hmaster0_p & v1214ee4 | !hmaster0_p & v1214eeb;
assign v121615c = hbusreq1 & v121615b | !hbusreq1 & v845542;
assign v16a13eb = hgrant5_p & v845542 | !hgrant5_p & !v16a2070;
assign v134cee5 = hbusreq5 & v134cee3 | !hbusreq5 & v134cee4;
assign d80793 = hgrant4_p & d80792 | !hgrant4_p & !v845542;
assign d2fe7d = hbusreq4_p & d2fe7c | !hbusreq4_p & v845542;
assign d301d1 = hgrant1_p & d301d0 | !hgrant1_p & d30786;
assign v16a1e61 = hbusreq2_p & v16a1da2 | !hbusreq2_p & v16a1e60;
assign v144634e = hbusreq3 & v1446338 | !hbusreq3 & v144634d;
assign v1668c8d = hgrant2_p & v1668c8b | !hgrant2_p & v1668c8c;
assign v1214dbf = hmaster1_p & v1214dbe | !hmaster1_p & !v1214d1e;
assign v144549f = hbusreq3 & v144549c | !hbusreq3 & v144549e;
assign v1405902 = hgrant2_p & v14058e6 | !hgrant2_p & v1405901;
assign v1445e32 = hbusreq3 & v1445e30 | !hbusreq3 & v1445e31;
assign v16a19d1 = hbusreq1_p & v16a183f | !hbusreq1_p & v16a19d0;
assign v1516959 = hgrant3_p & v15168b8 | !hgrant3_p & !v1516958;
assign v10d4067 = hgrant4_p & v10d3fe0 | !hgrant4_p & v10d4066;
assign a65498 = hbusreq2_p & a65494 | !hbusreq2_p & a65496;
assign v1214f14 = hbusreq5_p & v1214f13 | !hbusreq5_p & v1216547;
assign v10d408a = hmaster1_p & v10d4089 | !hmaster1_p & !v10d3fe9;
assign v14457d7 = hlock0 & v14457d6 | !hlock0 & v1445eb3;
assign v16a19e2 = hbusreq2_p & v16a1844 | !hbusreq2_p & v16a19e1;
assign v1284d60 = hmaster1_p & v1284d23 | !hmaster1_p & !v1284d1f;
assign v15160ff = hbusreq4_p & v15160fe | !hbusreq4_p & !v845542;
assign d2febb = hmaster2_p & d2feb4 | !hmaster2_p & d2feba;
assign v11e593e = hlock3_p & v11e593d | !hlock3_p & bf1f4f;
assign v12ad027 = hgrant5_p & v12ad60f | !hgrant5_p & !v12ad00b;
assign v1215b77 = hready & v845542 | !hready & v1216013;
assign v1445a36 = hmaster2_p & v14458d2 | !hmaster2_p & v144660b;
assign v12153e8 = hlock4_p & v12153e6 | !hlock4_p & !v12153e7;
assign v15534f3 = hbusreq2_p & v15534dd | !hbusreq2_p & v15534f2;
assign v1214bd7 = hbusreq2_p & v1214bd6 | !hbusreq2_p & v1214bd5;
assign v16a195a = hbusreq0 & v16a1957 | !hbusreq0 & v16a1959;
assign v1668c21 = hmaster2_p & v845542 | !hmaster2_p & v845570;
assign v1516803 = hbusreq2_p & v1516802 | !hbusreq2_p & !v845542;
assign d305e1 = hbusreq5_p & d305e0 | !hbusreq5_p & v845542;
assign v121503e = hgrant1_p & v1215466 | !hgrant1_p & v1215038;
assign v12165a4 = hbusreq5_p & v12165a3 | !hbusreq5_p & v845542;
assign v1214cd7 = hbusreq0 & v1214cd6 | !hbusreq0 & v845542;
assign v14058de = hmaster2_p & v14058c2 | !hmaster2_p & v1405844;
assign v1446283 = hmaster1_p & v1446282 | !hmaster1_p & v144627e;
assign d3013d = hgrant5_p & v84555a | !hgrant5_p & d300ea;
assign v1216188 = hgrant2_p & v1216187 | !hgrant2_p & v1216170;
assign v1215377 = locked_p & v1215376 | !locked_p & !v845542;
assign v121621f = hbusreq1_p & v121621e | !hbusreq1_p & v845542;
assign v12165b4 = decide_p & v1216583 | !decide_p & v12165b3;
assign v1445e1e = hmaster1_p & v1445e1d | !hmaster1_p & v1445e1b;
assign v12153db = hlock1_p & v12153da | !hlock1_p & v1215b97;
assign d2fb34 = hbusreq1_p & d2feb9 | !hbusreq1_p & d30660;
assign d30822 = hgrant5_p & v84554e | !hgrant5_p & d307b8;
assign v1446642 = hmaster2_p & v144639c | !hmaster2_p & v14465d8;
assign v1215d41 = hgrant5_p & v845570 | !hgrant5_p & v12165ac;
assign v12162ca = hmaster1_p & v12162c9 | !hmaster1_p & v1216224;
assign a65362 = hbusreq1_p & a6535e | !hbusreq1_p & a65361;
assign v1214c3a = hmaster1_p & v1214c2f | !hmaster1_p & v1214c39;
assign v14459ad = hready & v144639e | !hready & v14459a7;
assign v12ad672 = hbusreq0_p & v12ad671 | !hbusreq0_p & v845542;
assign a658a3 = stateG3_2_p & v845542 | !stateG3_2_p & !v9a051b;
assign v1216792 = hmaster0_p & v12165a9 | !hmaster0_p & v1668c1f;
assign v1445e8e = hlock1 & v1445e8d | !hlock1 & v1445e8b;
assign v10d4070 = hbusreq5_p & v10d406b | !hbusreq5_p & !v10d406f;
assign v144624b = stateG10_5_p & v144622b | !stateG10_5_p & !v144624a;
assign d306a1 = decide_p & d306a0 | !decide_p & v845570;
assign v1445411 = hmaster1_p & v14465aa | !hmaster1_p & v144626a;
assign v16a1dd6 = hmaster1_p & v9337f3 | !hmaster1_p & !v16a1f96;
assign d308bb = hbusreq5_p & d30839 | !hbusreq5_p & d308ba;
assign v151564e = hmaster2_p & v151564d | !hmaster2_p & a658b5;
assign v12ad631 = hmaster0_p & v12ad5e5 | !hmaster0_p & v12ad4f4;
assign d3026d = hbusreq5_p & d3026c | !hbusreq5_p & !d3026b;
assign v114a22f = hready_p & v845542 | !hready_p & !v845568;
assign d2f9ba = hmaster1_p & d2f9b9 | !hmaster1_p & d2f995;
assign v1668c82 = hgrant2_p & v1668c7e | !hgrant2_p & v1668c81;
assign v138a358 = hbusreq2 & v138a347 | !hbusreq2 & v138a357;
assign v16a2073 = hready & v16a2072 | !hready & !v845542;
assign v134ce6c = hlock5 & v134ce5d | !hlock5 & v134ce6b;
assign v1405aab = hbusreq4_p & v1405aaa | !hbusreq4_p & v1405a87;
assign v16a1395 = hbusreq2_p & v16a12c3 | !hbusreq2_p & v16a1394;
assign v15530a2 = hbusreq3 & v15530a0 | !hbusreq3 & v15530a1;
assign v138a391 = hmaster1_p & v845542 | !hmaster1_p & !v138a390;
assign f2e4dd = hgrant2_p & v845542 | !hgrant2_p & f2e4dc;
assign v14454f1 = hmaster1_p & v14454f0 | !hmaster1_p & v14462ff;
assign v15156ad = hbusreq1_p & v1668cd3 | !hbusreq1_p & v1668ce3;
assign v144616a = hbusreq2_p & v1446165 | !hbusreq2_p & v1446169;
assign v12153ab = hmaster2_p & v1215392 | !hmaster2_p & v845547;
assign d3024a = hgrant5_p & v845542 | !hgrant5_p & d301ff;
assign v12ad02f = hgrant2_p & v12acff7 | !hgrant2_p & v12ad02e;
assign v1405b59 = hbusreq2_p & v1405b56 | !hbusreq2_p & v1405b58;
assign v1515818 = decide_p & v1515817 | !decide_p & v845542;
assign v1405ac8 = hmaster0_p & v1405ac3 | !hmaster0_p & v1405ac7;
assign v1215773 = hmaster2_p & v12160ec | !hmaster2_p & !v1215734;
assign bf1f9c = hgrant0_p & v845570 | !hgrant0_p & d2fc50;
assign v151566c = hmaster1_p & v1515650 | !hmaster1_p & v151566b;
assign v1445fd2 = hbusreq0 & v1445fce | !hbusreq0 & v1445fd1;
assign v1445dfb = hbusreq4_p & v1446421 | !hbusreq4_p & v1446429;
assign v87abb5 = stateG3_0_p & v845542 | !stateG3_0_p & a81304;
assign v1216582 = hbusreq2 & v1216579 | !hbusreq2 & v1216581;
assign v12164d5 = hbusreq5_p & v12164d4 | !hbusreq5_p & v16a2243;
assign d301bb = hmaster2_p & d306c8 | !hmaster2_p & v845542;
assign v1216a64 = hburst1_p & v134d1d9 | !hburst1_p & v1216a63;
assign d3082c = hgrant5_p & v84554e | !hgrant5_p & d307ee;
assign v144628a = hlock3 & v1446275 | !hlock3 & v1446289;
assign d2fb1e = hbusreq5_p & d30157 | !hbusreq5_p & d2fb1d;
assign d2fc57 = hmaster2_p & d2fc4f | !hmaster2_p & d2fc56;
assign v1446616 = hgrant5_p & v144642c | !hgrant5_p & v1446615;
assign a65b3f = jx2_p & a65b38 | !jx2_p & a65b3d;
assign v1214c8c = hlock5_p & v1214c8a | !hlock5_p & v1214c8b;
assign v121628f = hbusreq2_p & v121628d | !hbusreq2_p & v121628e;
assign v1668d83 = hgrant1_p & v1668d65 | !hgrant1_p & v1668d82;
assign v16a1973 = hmaster2_p & v16a208a | !hmaster2_p & v16a1970;
assign v1405a8e = hmaster2_p & v1405a87 | !hmaster2_p & !v1405a8c;
assign v10d4013 = hready_p & v10d4002 | !hready_p & !v10d4012;
assign v1284d32 = hmaster0_p & v1284cad | !hmaster0_p & v1284c98;
assign v144649b = hgrant0_p & v144649a | !hgrant0_p & v845542;
assign v134d3e0 = hgrant5_p & v845542 | !hgrant5_p & v134d3df;
assign d307c4 = hbusreq4 & v845542 | !hbusreq4 & !d3070c;
assign v1445852 = hbusreq2 & v144584e | !hbusreq2 & v1445851;
assign v144644d = hmaster0_p & v1446417 | !hmaster0_p & v144642d;
assign v12153a8 = hbusreq0 & v12153a7 | !hbusreq0 & v845542;
assign v1445e48 = hmaster2_p & v1446493 | !hmaster2_p & v1445e47;
assign v1446264 = hmaster2_p & v1446407 | !hmaster2_p & v1446415;
assign f2f3fa = hmaster1_p & f2f3f9 | !hmaster1_p & f2f2db;
assign v151575d = hbusreq5_p & v1515759 | !hbusreq5_p & !v151575c;
assign a65b19 = hbusreq2_p & a65b0d | !hbusreq2_p & a65b18;
assign f2f21c = hbusreq1_p & f2f21b | !hbusreq1_p & !v845542;
assign d306a8 = hgrant5_p & v845542 | !hgrant5_p & !d306a7;
assign v1668c61 = hmaster0_p & v1668c5f | !hmaster0_p & v1668c60;
assign v15156b6 = stateA1_p & v146af2e | !stateA1_p & !v110b6cc;
assign d8075c = hmastlock_p & d8075b | !hmastlock_p & !v845542;
assign d300f2 = hgrant1_p & d300e8 | !hgrant1_p & d300c3;
assign v140584c = hmaster2_p & v1405849 | !hmaster2_p & v140584b;
assign v1214ee2 = hlock5_p & v1214ee0 | !hlock5_p & v1214ee1;
assign hgrant5 = !v1388ce9;
assign a65475 = hbusreq0 & a658d8 | !hbusreq0 & a65474;
assign v1215443 = hmaster0_p & v12153ee | !hmaster0_p & v12153d4;
assign v10d4305 = jx0_p & v10d40de | !jx0_p & v10d4304;
assign a65921 = hmaster1_p & a658fb | !hmaster1_p & !a65916;
assign v1214efb = hmaster1_p & v1214eef | !hmaster1_p & v1214efa;
assign v1214c96 = hbusreq0 & v1214c95 | !hbusreq0 & v845542;
assign d3081f = hgrant5_p & d3081e | !hgrant5_p & d307a8;
assign v144631b = hbusreq0 & v144631a | !hbusreq0 & v14462e7;
assign d2f99b = hmaster2_p & d2f99a | !hmaster2_p & d3068e;
assign d306b5 = hbusreq0 & d306b3 | !hbusreq0 & d306b4;
assign a66280 = decide_p & a6627f | !decide_p & v845542;
assign v1445ed7 = hmaster1_p & v1445ed6 | !hmaster1_p & v1445e1b;
assign v12acfec = hbusreq2 & v12acfe6 | !hbusreq2 & v12acfeb;
assign v1214dd4 = hmaster0_p & v1216a74 | !hmaster0_p & v845542;
assign v16a1bb4 = stateA1_p & v845542 | !stateA1_p & !v16a1af5;
assign v1214bdc = hbusreq2_p & v1214bdb | !hbusreq2_p & v1214bda;
assign v1446304 = hlock0 & v1446303 | !hlock0 & v1446302;
assign v151567e = hmaster2_p & v1515675 | !hmaster2_p & !v1668cbd;
assign v155309a = hmaster1_p & v1553385 | !hmaster1_p & v1553099;
assign a662cf = hbusreq1_p & a66298 | !hbusreq1_p & a66289;
assign v1215763 = hbusreq5_p & v1215761 | !hbusreq5_p & v1215762;
assign v12ad519 = hlock0_p & v1515654 | !hlock0_p & v12ad518;
assign v1216a6c = hbusreq5_p & v1216a6b | !hbusreq5_p & v845542;
assign v16a2094 = hbusreq0 & v16a207a | !hbusreq0 & v16a2093;
assign v134d36e = hready & v134d36d | !hready & v134d273;
assign v140582a = jx2_p & v85e75f | !jx2_p & v85e749;
assign v134cece = decide_p & v134cec0 | !decide_p & v134cecd;
assign v1215467 = hbusreq1_p & v1215bac | !hbusreq1_p & v1215466;
assign v12161a8 = hlock2_p & v1216183 | !hlock2_p & v12161a7;
assign v144554f = hmaster1_p & v1446310 | !hmaster1_p & v1445544;
assign v15157ae = hgrant1_p & v15157a8 | !hgrant1_p & v151579a;
assign v1214bfa = hmaster1_p & v1214bf9 | !hmaster1_p & v12153a9;
assign ab83a0 = stateG3_2_p & v88d3e4 | !stateG3_2_p & v92fc87;
assign d306be = hbusreq5_p & v845542 | !hbusreq5_p & !d306b2;
assign v144541d = hmaster1_p & v1445414 | !hmaster1_p & v1446329;
assign v1215d03 = hbusreq0 & v1215d00 | !hbusreq0 & v1215d02;
assign v16a12f7 = hbusreq2 & v16a12f5 | !hbusreq2 & !v16a12f6;
assign v134cd83 = hgrant2_p & v134cd73 | !hgrant2_p & v134cd81;
assign d30671 = hbusreq2_p & d3066f | !hbusreq2_p & d30670;
assign v1445ade = hbusreq2 & v1445adc | !hbusreq2 & v1445add;
assign v140589e = hgrant5_p & v1405897 | !hgrant5_p & v140589d;
assign v1446038 = decide_p & v144602c | !decide_p & v1446564;
assign v1445a65 = hmaster1_p & v1445a64 | !hmaster1_p & v144590e;
assign d2fb29 = hbusreq0 & d2fb26 | !hbusreq0 & d2fb28;
assign d2fadb = hbusreq1_p & d300bd | !hbusreq1_p & d2fada;
assign v138a477 = hready_p & v138a449 | !hready_p & !v138a476;
assign v12166c5 = hgrant1_p & v12164cf | !hgrant1_p & v12166c4;
assign v1446044 = hmaster2_p & v1446043 | !hmaster2_p & v1446412;
assign v1668dc1 = hmaster0_p & v1668db9 | !hmaster0_p & v1668dc0;
assign v16a19ce = hready_p & v16a1985 | !hready_p & v16a19cd;
assign v121535b = hmaster1_p & v121535a | !hmaster1_p & v1215357;
assign d30613 = hbusreq5_p & d30612 | !hbusreq5_p & v845542;
assign v16a194e = hgrant5_p & v845542 | !hgrant5_p & v16a194d;
assign v1216a8c = locked_p & v1216a8b | !locked_p & !v845542;
assign v151584b = hlock2_p & v151584a | !hlock2_p & v1515802;
assign v151561c = locked_p & v151561b | !locked_p & !v845542;
assign v12ad014 = hgrant5_p & v12ad644 | !hgrant5_p & v12ad013;
assign d30118 = hbusreq5_p & d30117 | !hbusreq5_p & !d30116;
assign v14466ae = hbusreq0 & v14466ad | !hbusreq0 & v1446648;
assign v16a1ca4 = hmaster0_p & v16a1c9f | !hmaster0_p & v16a1c9b;
assign f2f3f0 = hmaster1_p & f2f3ef | !hmaster1_p & f2f2db;
assign v16a13c3 = hbusreq2 & v16a13c2 | !hbusreq2 & v16a1da5;
assign v12ad610 = hgrant5_p & v12ad60f | !hgrant5_p & !v12ad5cc;
assign f2f4b4 = hmaster2_p & v845542 | !hmaster2_p & !f2f4b3;
assign d80742 = hlock4_p & d80732 | !hlock4_p & !v845542;
assign f2f380 = hgrant5_p & f2f2a1 | !hgrant5_p & !f2f37f;
assign v1284d2a = hgrant3_p & v1284cc1 | !hgrant3_p & v1284d29;
assign d307cf = hlock0_p & v845542 | !hlock0_p & d307ce;
assign v11e595b = hgrant5_p & v845542 | !hgrant5_p & v11e595a;
assign v15156c8 = hmaster2_p & v1515675 | !hmaster2_p & v15156c7;
assign v134d518 = hbusreq0 & v134d516 | !hbusreq0 & v134d517;
assign v12ad5a6 = hgrant0_p & a6537d | !hgrant0_p & !v12ad5a5;
assign v1515ae5 = hbusreq4 & d305de | !hbusreq4 & d30645;
assign d2fbd6 = hmaster2_p & d2fbd2 | !hmaster2_p & d2fbd5;
assign v1446558 = hgrant1_p & v1446398 | !hgrant1_p & v845542;
assign v1445a1d = hgrant1_p & v14458f6 | !hgrant1_p & v1445a17;
assign v1445fae = hmaster0_p & v1445f8f | !hmaster0_p & v1445f99;
assign v12160ee = hlock0_p & v1215fe8 | !hlock0_p & !v121601c;
assign v1515715 = hbusreq4_p & v1515713 | !hbusreq4_p & v1515714;
assign a653f5 = hmaster2_p & a65372 | !hmaster2_p & a653b4;
assign v1215bc3 = hmaster1_p & v121639f | !hmaster1_p & v1215bc2;
assign d2fed3 = hbusreq2_p & d2fed2 | !hbusreq2_p & d2feca;
assign v16a209c = hbusreq0 & v16a209a | !hbusreq0 & v16a209b;
assign v144586a = hgrant3_p & v14457d5 | !hgrant3_p & v1445869;
assign v144548d = hlock3 & v144546f | !hlock3 & v144548c;
assign v10d4041 = hbusreq4_p & v10d4022 | !hbusreq4_p & v10d402f;
assign a6563b = hgrant1_p & a6539b | !hgrant1_p & !a6562d;
assign v1215fbd = hmaster0_p & v12166f7 | !hmaster0_p & v1216702;
assign v14465c9 = hgrant4_p & v144640a | !hgrant4_p & v14465c8;
assign v1445378 = hbusreq3 & v1445376 | !hbusreq3 & v1445377;
assign v1445aa3 = hbusreq2_p & v1445a9d | !hbusreq2_p & v1445aa2;
assign v151578c = stateA1_p & v1515670 | !stateA1_p & v151578b;
assign v121670f = hmaster1_p & v1216702 | !hmaster1_p & v12166ef;
assign v138a315 = hmaster1_p & v138a310 | !hmaster1_p & v138a314;
assign v15168f7 = hlock1_p & v15168f5 | !hlock1_p & !v15168f6;
assign f2f4ae = hburst1 & a658a5 | !hburst1 & f2f4ad;
assign d80749 = hmaster0_p & d8073b | !hmaster0_p & d80748;
assign v1215c19 = hbusreq1_p & v1216537 | !hbusreq1_p & v121612e;
assign f2f4ba = hbusreq2_p & f2f4ac | !hbusreq2_p & f2f4b9;
assign v1446335 = hgrant2_p & v1446334 | !hgrant2_p & v1446324;
assign v1214db0 = hbusreq2_p & v1214dab | !hbusreq2_p & v1214daf;
assign v1445bb5 = hmaster0_p & v1446636 | !hmaster0_p & v1446404;
assign d80769 = hlock2_p & d80768 | !hlock2_p & v845542;
assign v1215392 = hlock0_p & v1215391 | !hlock0_p & !v845542;
assign v15530ad = hlock3 & v155321a | !hlock3 & v15530ac;
assign v1445e6a = hbusreq1 & v1445e66 | !hbusreq1 & v1445e69;
assign v12161a1 = hbusreq0 & v121619f | !hbusreq0 & v12161a0;
assign v1445b6b = hgrant2_p & v1445b69 | !hgrant2_p & v1445b6a;
assign d2fb48 = decide_p & d2fb47 | !decide_p & v845570;
assign f2ed9d = hready_p & f2ed9b | !hready_p & f2ed9c;
assign v1215ca9 = hlock5_p & v1215ca7 | !hlock5_p & !v1215ca8;
assign v1446408 = hready & v1446406 | !hready & v1446407;
assign v1215bdc = hmaster0_p & v1215bda | !hmaster0_p & v1215bdb;
assign v10d429f = hmaster2_p & v10d429e | !hmaster2_p & v10d4079;
assign d2fb5f = decide_p & d2fb5e | !decide_p & v845570;
assign v1445807 = hgrant2_p & v1445804 | !hgrant2_p & v1445806;
assign v1445ebf = hlock1 & v1446606 | !hlock1 & v1445e57;
assign v16a1cec = hmaster2_p & v16a1ceb | !hmaster2_p & v16a206f;
assign v1445529 = hbusreq3 & v1445527 | !hbusreq3 & v1445528;
assign v12164db = hbusreq5_p & v12164da | !hbusreq5_p & v845542;
assign v16a1401 = hbusreq2_p & v16a1400 | !hbusreq2_p & v16a1d54;
assign a653ef = hmaster2_p & a653a9 | !hmaster2_p & !a653aa;
assign d2fb81 = hlock2_p & d2fb7c | !hlock2_p & d2fb80;
assign d2fd14 = hlock2_p & v845542 | !hlock2_p & !d2fd13;
assign v16a19c9 = hgrant2_p & v16a1f9b | !hgrant2_p & v16a19c8;
assign v1216258 = hgrant2_p & v1216229 | !hgrant2_p & v1216257;
assign v1553105 = decide_p & v155342e | !decide_p & v1553104;
assign v144639f = hlock4 & v144639c | !hlock4 & v144639e;
assign a66294 = hmastlock_p & a66293 | !hmastlock_p & v845542;
assign v15156ee = hbusreq2 & v15156ed | !hbusreq2 & v15167ed;
assign v12ad500 = hmaster1_p & v12ad4f5 | !hmaster1_p & v12ad4ff;
assign v14463e5 = hbusreq0_p & v14463b1 | !hbusreq0_p & !v14463d8;
assign v12152ea = hmaster1_p & v12152e9 | !hmaster1_p & v1215770;
assign a654be = hmaster1_p & a658f1 | !hmaster1_p & !a654b0;
assign v1446429 = hlock0_p & v1446403 | !hlock0_p & v1446428;
assign v1214d2c = hmaster1_p & v1214d2b | !hmaster1_p & !v1214d1e;
assign v16a1c05 = decide_p & v16a1bed | !decide_p & v16a1c04;
assign a64716 = jx2_p & a64715 | !jx2_p & a65b3d;
assign v10d4039 = hbusreq1_p & v10d3fe0 | !hbusreq1_p & v10d3fdf;
assign v1216700 = hmaster2_p & v12166c5 | !hmaster2_p & v845570;
assign v16a142f = hbusreq2 & v16a142e | !hbusreq2 & !v16a1aed;
assign v16a1449 = jx2_p & v16a1435 | !jx2_p & v16a1448;
assign v134cea5 = hbusreq2 & v134cea4 | !hbusreq2 & v134d240;
assign d3086f = hmaster0_p & d30866 | !hmaster0_p & d3086e;
assign v1445bda = hmaster1_p & v1446643 | !hmaster1_p & v1445bd5;
assign v16a1ae7 = hbusreq5_p & v16a209a | !hbusreq5_p & v16a1ae6;
assign v13897f0 = hmaster1_p & v1389de1 | !hmaster1_p & v13897ef;
assign v16a1a2e = hbusreq3 & v16a1a28 | !hbusreq3 & v16a1a2d;
assign v134d42e = hmaster2_p & v134d427 | !hmaster2_p & v134d42d;
assign a656a2 = hmaster1_p & a6548f | !hmaster1_p & !a65916;
assign v12afa0b = hbusreq0 & v12af9c3 | !hbusreq0 & v12afa0a;
assign v14460a2 = hbusreq1_p & v1446677 | !hbusreq1_p & v14465bb;
assign v144604e = hbusreq1_p & v14465ce | !hbusreq1_p & v14465d7;
assign v1446660 = hgrant5_p & v1446445 | !hgrant5_p & v144665f;
assign v134cd61 = hgrant0_p & v134cd60 | !hgrant0_p & v845542;
assign v16a137f = hbusreq5 & v16a1373 | !hbusreq5 & v16a137e;
assign v10d4286 = stateA1_p & v845542 | !stateA1_p & v10d4264;
assign d2fc6f = hgrant2_p & d2fc28 | !hgrant2_p & d2fc6e;
assign v12162fe = hmaster2_p & v845547 | !hmaster2_p & v12162fc;
assign f2f29d = hbusreq1 & v1668d1c | !hbusreq1 & v845542;
assign v12ad035 = hbusreq5 & v12ad020 | !hbusreq5 & v12ad034;
assign v14463d3 = hbusreq2 & v14463cc | !hbusreq2 & v14463d2;
assign a65646 = hmaster2_p & a662ac | !hmaster2_p & a65645;
assign v12acfda = hbusreq0 & v12acfd9 | !hbusreq0 & !v12af73f;
assign v1552f61 = hgrant4_p & v845542 | !hgrant4_p & v1552f60;
assign v1445db2 = hmaster0_p & v144639c | !hmaster0_p & v1445da9;
assign v16a1940 = hgrant4_p & v845559 | !hgrant4_p & v16a193f;
assign v1445ec6 = hmaster2_p & v144639c | !hmaster2_p & v1445e10;
assign v1214c36 = hbusreq4_p & d2fbe5 | !hbusreq4_p & v1214c30;
assign v12167a4 = hmaster1_p & v12167a3 | !hmaster1_p & v12165a5;
assign f2ed93 = hmaster1_p & f2f22b | !hmaster1_p & f2ed92;
assign f2f2d4 = hbusreq1 & a658d6 | !hbusreq1 & v845542;
assign v1552f82 = hbusreq2_p & v1552f80 | !hbusreq2_p & v1552f81;
assign v11e595c = hmaster0_p & v11e5951 | !hmaster0_p & !v11e595b;
assign v1214d82 = hmaster1_p & v1214d81 | !hmaster1_p & v1214c92;
assign v16a2247 = hmaster0_p & v16a2240 | !hmaster0_p & v16a2246;
assign f2f52d = hmaster1_p & f2f229 | !hmaster1_p & f2f52c;
assign v12160d5 = hmaster2_p & v12160d1 | !hmaster2_p & f2f2a8;
assign v1284d39 = hlock0_p & v140588d | !hlock0_p & v1284d37;
assign v1553380 = hmaster1_p & v155337f | !hmaster1_p & v845542;
assign v14457f4 = hmaster1_p & v1445eb8 | !hmaster1_p & v1445ed3;
assign v16a1d55 = hgrant2_p & v845542 | !hgrant2_p & !v16a1d53;
assign d30243 = hgrant5_p & d30242 | !hgrant5_p & !d301ed;
assign d2fb95 = hlock2_p & d2fb94 | !hlock2_p & d2fb90;
assign v1446013 = hbusreq1_p & v1446484 | !hbusreq1_p & v144649c;
assign v12af21b = hbusreq1_p & v12afe4e | !hbusreq1_p & v12af9bf;
assign v1553092 = hbusreq2 & v1553090 | !hbusreq2 & v1553091;
assign v1405ad2 = hlock2_p & v1405ad1 | !hlock2_p & v1405a9a;
assign v14458ed = hmaster2_p & v14458e2 | !hmaster2_p & v14458eb;
assign v14460c1 = hlock2 & v14460bc | !hlock2 & v14460c0;
assign v1284cb4 = hlock2_p & v1284cb2 | !hlock2_p & v1284cb3;
assign v1445540 = decide_p & v144553f | !decide_p & v1446275;
assign v121533b = hmaster1_p & v12150aa | !hmaster1_p & !v12150a6;
assign d3019d = hbusreq5_p & d3019c | !hbusreq5_p & d30913;
assign v16a1d5f = hbusreq0 & v16a209a | !hbusreq0 & v16a1d5e;
assign v1214fb7 = hgrant0_p & v1215766 | !hgrant0_p & v845542;
assign v1445371 = hmaster1_p & v1445370 | !hmaster1_p & v14458fd;
assign v12af984 = hbusreq4_p & v12afda3 | !hbusreq4_p & v12af983;
assign v134d3fa = hlock3_p & v134d240 | !hlock3_p & v134d270;
assign v1445d99 = hbusreq4_p & v14463b5 | !hbusreq4_p & v14463bb;
assign v138a06a = hmaster1_p & v845542 | !hmaster1_p & !v138a069;
assign v134cec6 = hbusreq3 & v134cec4 | !hbusreq3 & v134cec5;
assign v14058b0 = hgrant5_p & v140584c | !hgrant5_p & v14058af;
assign d308d9 = hbusreq1 & v845542 | !hbusreq1 & d30740;
assign d30807 = hgrant2_p & d307f9 | !hgrant2_p & !d30806;
assign v1216540 = hbusreq1_p & v121653f | !hbusreq1_p & v845547;
assign v1445b38 = hmaster1_p & v1445a43 | !hmaster1_p & v1445a32;
assign v1214ef1 = hgrant5_p & v1214ef0 | !hgrant5_p & v1216547;
assign v134d538 = hbusreq3 & v134d536 | !hbusreq3 & v134d537;
assign v1515845 = hgrant5_p & v845570 | !hgrant5_p & v1515837;
assign f2f4c4 = hready_p & v845542 | !hready_p & f2f4c3;
assign v84555a = hlock4_p & v845542 | !hlock4_p & !v845542;
assign d2fb79 = hmaster2_p & d2fb78 | !hmaster2_p & v845542;
assign d3015e = hgrant2_p & d3012a | !hgrant2_p & d3014f;
assign v1445ab6 = hmaster1_p & v14458a6 | !hmaster1_p & v144589f;
assign v1446187 = hmaster0_p & v1445fea | !hmaster0_p & v1446079;
assign v1215b7f = hmaster0_p & v1215b7c | !hmaster0_p & v1215b7e;
assign v1215d0d = hlock3_p & v1215c7b | !hlock3_p & v1215d0c;
assign v134ce98 = hmaster2_p & v134ce8c | !hmaster2_p & v134d1fc;
assign v16a13ff = hmaster1_p & v16a13fe | !hmaster1_p & v16a1d6d;
assign a65867 = hmaster2_p & a65863 | !hmaster2_p & a65864;
assign v134d267 = hlock2_p & v134d266 | !hlock2_p & v134d244;
assign v84556a = hmastlock_p & v845542 | !hmastlock_p & !v845542;
assign d2fef4 = hbusreq2_p & d2fef3 | !hbusreq2_p & d2feef;
assign d30855 = hbusreq1_p & d30704 | !hbusreq1_p & !v845542;
assign f2f2c8 = hbusreq1 & a658ad | !hbusreq1 & v845542;
assign v16a1433 = hready_p & v16a1431 | !hready_p & v16a1432;
assign v1214d08 = hbusreq0 & v1214d07 | !hbusreq0 & v16a2243;
assign v16a1d43 = hbusreq0 & v16a1d3b | !hbusreq0 & v16a1d42;
assign d2fc44 = hbusreq2_p & d2fbbf | !hbusreq2_p & d2fc42;
assign v1445fa5 = hbusreq2_p & v1445f9f | !hbusreq2_p & v1445fa4;
assign v14458ae = hlock2 & v14458a9 | !hlock2 & v14458ad;
assign v12153a5 = hlock4_p & v12153a4 | !hlock4_p & v1215364;
assign v1553235 = hgrant1_p & v845542 | !hgrant1_p & v1553234;
assign v14457c2 = hlock3 & v14457b9 | !hlock3 & v14457c1;
assign d30151 = hgrant5_p & d2fe80 | !hgrant5_p & d30114;
assign v1445ee8 = hmaster1_p & v14465aa | !hmaster1_p & v1445e28;
assign v1516982 = hbusreq2 & v151697c | !hbusreq2 & v1516981;
assign d2fc8c = hbusreq2 & d2fc8b | !hbusreq2 & v845542;
assign d2fecf = hmaster2_p & d2feb2 | !hmaster2_p & d2fece;
assign v16a20a0 = hbusreq5 & v16a2099 | !hbusreq5 & v16a209f;
assign v1216140 = hbusreq1 & v121613f | !hbusreq1 & v845542;
assign v12ad598 = hbusreq1 & v12ad4ca | !hbusreq1 & v12ad4e4;
assign d3071f = hmaster2_p & d3071d | !hmaster2_p & v84554e;
assign v16a1e90 = hmaster2_p & v16a1e8f | !hmaster2_p & v16a206f;
assign v1446141 = hmaster1_p & v1446118 | !hmaster1_p & v1445ffc;
assign v1445ad9 = hbusreq2_p & v1445ad7 | !hbusreq2_p & v1445ad8;
assign v12af9b2 = hbusreq5_p & v12afdb1 | !hbusreq5_p & v12af98a;
assign d300e9 = hgrant1_p & d300e8 | !hgrant1_p & d300dd;
assign f2f3c9 = hgrant5_p & v84554c | !hgrant5_p & f2f37f;
assign v121616a = hmaster2_p & v1216161 | !hmaster2_p & v1216169;
assign v1214d48 = hmaster2_p & v1214d47 | !hmaster2_p & v845542;
assign v134ce34 = hlock0_p & v134d370 | !hlock0_p & v134ce33;
assign v12ad0b7 = hgrant1_p & v12ad0b6 | !hgrant1_p & v12afdab;
assign v15534d1 = hmaster2_p & v15534d0 | !hmaster2_p & v15533a2;
assign v144544d = hbusreq2_p & v144544c | !hbusreq2_p & v1445bb3;
assign v1446401 = hlock5 & v14463d1 | !hlock5 & v1446400;
assign v16a1bdf = hbusreq2 & v16a1bdd | !hbusreq2 & !v16a1bde;
assign v1216149 = hbusreq0_p & v845547 | !hbusreq0_p & v121611d;
assign v1405b3d = hmaster0_p & v1405a96 | !hmaster0_p & v1405a89;
assign d2fc28 = hmaster1_p & d2fc23 | !hmaster1_p & d2fc27;
assign d2feef = hmaster1_p & d2fed8 | !hmaster1_p & d2fee5;
assign v14460ee = hlock2 & v14460ea | !hlock2 & v14460ed;
assign v10d40b7 = hgrant2_p & v10d40b4 | !hgrant2_p & v10d40b6;
assign v1214c1d = hlock2_p & v1214c1b | !hlock2_p & v1214c1c;
assign v140591c = hmaster1_p & v140591b | !hmaster1_p & v140584d;
assign f2f40c = hmaster1_p & f2f3fb | !hmaster1_p & !f2f330;
assign v1216154 = hlock1_p & v121614d | !hlock1_p & v1216153;
assign d30777 = hbusreq2_p & d30776 | !hbusreq2_p & d30772;
assign d30220 = hmaster2_p & d306c8 | !hmaster2_p & d306d4;
assign v14453b2 = hmaster1_p & v1445361 | !hmaster1_p & v1445a9b;
assign v155298e = jx2_p & v1552963 | !jx2_p & v155298d;
assign v12af1c0 = hmaster0_p & v12af73f | !hmaster0_p & v12af1bf;
assign d2fc17 = hbusreq2_p & d2fc16 | !hbusreq2_p & d2fc14;
assign v90d5cd = hmaster0_p & b09421 | !hmaster0_p & !v84555c;
assign v10d40c1 = hgrant1_p & v10d4019 | !hgrant1_p & v10d40c0;
assign v16a1bfb = hgrant5_p & v845542 | !hgrant5_p & !v16a1bf0;
assign v10d426f = hbusreq5_p & v10d426d | !hbusreq5_p & !v10d426e;
assign v1445547 = hmaster1_p & v144632c | !hmaster1_p & v1445544;
assign v14463c7 = hbusreq5_p & v144639c | !hbusreq5_p & v14463c5;
assign v1216714 = hgrant0_p & v845547 | !hgrant0_p & v845542;
assign v14462f9 = hgrant5_p & v1446433 | !hgrant5_p & v144662b;
assign v1445ac5 = hmaster1_p & v1445ac4 | !hmaster1_p & v144589f;
assign d308b8 = hgrant5_p & d30654 | !hgrant5_p & d3088b;
assign d3075a = hlock2_p & d30759 | !hlock2_p & d30756;
assign v15533b4 = hbusreq0 & v15533b3 | !hbusreq0 & v15533a8;
assign v1445757 = hmaster1_p & v1445f27 | !hmaster1_p & v1445dd1;
assign d2ff08 = hbusreq2_p & d2ff07 | !hbusreq2_p & d2ff03;
assign v1446493 = hgrant1_p & v845542 | !hgrant1_p & v144648d;
assign v1215da1 = hgrant2_p & v1215d7d | !hgrant2_p & v1215da0;
assign v16a1375 = hgrant2_p & v16a205f | !hgrant2_p & v16a1374;
assign v1445998 = hgrant0_p & v144639c | !hgrant0_p & v1445997;
assign v1668d9d = hmaster2_p & v1668d2f | !hmaster2_p & v1668d5d;
assign v1215472 = hmaster0_p & v1215462 | !hmaster0_p & v1215471;
assign d2feec = hbusreq2_p & d2feeb | !hbusreq2_p & d2fee7;
assign v1215369 = hbusreq5_p & v1215367 | !hbusreq5_p & v1215368;
assign v1445e19 = hbusreq2_p & v1445e08 | !hbusreq2_p & v1445e18;
assign v1215c64 = hgrant5_p & v16a2243 | !hgrant5_p & v1215c20;
assign v1216091 = hlock1_p & v1216090 | !hlock1_p & !v84554d;
assign v12ad5a3 = locked_p & v151571b | !locked_p & v12ad5a2;
assign v15167f4 = hlock2_p & v15167f3 | !hlock2_p & !v845542;
assign v15155f3 = hmaster1_p & v15155f2 | !hmaster1_p & v845570;
assign v16a13f4 = hbusreq0 & v16a13f2 | !hbusreq0 & v16a13f3;
assign v1215325 = hmaster1_p & v121505b | !hmaster1_p & v1215054;
assign v151579c = hmaster2_p & v1515793 | !hmaster2_p & v151579b;
assign v14465b4 = hmaster2_p & v14465b0 | !hmaster2_p & v14465b3;
assign v1445b12 = hbusreq2_p & v1445b0e | !hbusreq2_p & v1445b11;
assign v1389538 = hmaster2_p & v16693a6 | !hmaster2_p & !v845542;
assign v1445f08 = hlock0 & v1445f07 | !hlock0 & v1445f06;
assign v1215c59 = hbusreq0 & v1215c57 | !hbusreq0 & v1215c58;
assign v1445abe = hmaster1_p & v14458a2 | !hmaster1_p & v14458af;
assign v1446167 = hmaster1_p & v1446166 | !hmaster1_p & v1445fde;
assign v1445b31 = hmaster0_p & v1445902 | !hmaster0_p & v14458d3;
assign v14453a2 = hlock3 & v1445354 | !hlock3 & v14453a0;
assign v1215daf = hready_p & v1215d47 | !hready_p & v1215dae;
assign v1668d59 = hbusreq1_p & v1668d3b | !hbusreq1_p & v1668d58;
assign v16a1be4 = hbusreq0 & v16a209a | !hbusreq0 & v16a1be3;
assign v1214cbc = hgrant1_p & d2fbe5 | !hgrant1_p & v1214cbb;
assign v1445b81 = hgrant2_p & v1445b6e | !hgrant2_p & v1445b80;
assign v138a067 = hlock5_p & v138a066 | !hlock5_p & !v845542;
assign v1446159 = hbusreq2 & v1446157 | !hbusreq2 & v1446158;
assign v14463a0 = hbusreq4 & v144639e | !hbusreq4 & v144639f;
assign v144615d = hlock5 & v1446125 | !hlock5 & v144615b;
assign v1214c0e = hlock2_p & v1214c0c | !hlock2_p & v1214c0d;
assign v1214cfc = hbusreq5_p & v1214cf7 | !hbusreq5_p & !v1214cfb;
assign v1215355 = hmaster2_p & v1215354 | !hmaster2_p & v845542;
assign v1446483 = hgrant0_p & v1446482 | !hgrant0_p & v845542;
assign v12166e1 = hbusreq5_p & v12166e0 | !hbusreq5_p & v845542;
assign v1515618 = stateA1_p & v845542 | !stateA1_p & !a65364;
assign v140589d = hmaster2_p & v14463b1 | !hmaster2_p & v140589c;
assign v14461e9 = hgrant2_p & v14461bd | !hgrant2_p & v14461e5;
assign v1215cb7 = hbusreq5_p & v1215cb3 | !hbusreq5_p & !v1215cb6;
assign v1515610 = hmaster2_p & v151560d | !hmaster2_p & v151560e;
assign d30117 = hlock5_p & d30115 | !hlock5_p & !d30116;
assign v1445470 = hlock2 & v144546f | !hlock2 & v144546e;
assign v144632b = hgrant2_p & v1446328 | !hgrant2_p & v144632a;
assign v12ad553 = hmaster1_p & v12ad52e | !hmaster1_p & v12ad54f;
assign v1445393 = hmaster1_p & v1445364 | !hmaster1_p & v144591b;
assign v138a059 = decide_p & v1389fcc | !decide_p & v138a406;
assign v12ad8ea = hbusreq5_p & v12add49 | !hbusreq5_p & v12ad8e9;
assign v10d42a2 = hmaster1_p & v10d428d | !hmaster1_p & !v10d42a1;
assign a658b6 = hbusreq4_p & a658b5 | !hbusreq4_p & v845542;
assign v1515c84 = hlock2_p & v1515c83 | !hlock2_p & v845542;
assign v144581c = hbusreq3 & v144581a | !hbusreq3 & v144581b;
assign v1446464 = hgrant1_p & v845542 | !hgrant1_p & v1446463;
assign v1405b37 = hmaster0_p & v1405af3 | !hmaster0_p & v1405a96;
assign d2fc63 = hgrant5_p & v84554a | !hgrant5_p & d2fc62;
assign v1214ec9 = hgrant5_p & v845547 | !hgrant5_p & v121652f;
assign v12ad4d6 = hmaster2_p & v12ad4d0 | !hmaster2_p & v12ad4d5;
assign v1445f8a = stateG10_5_p & v1445f89 | !stateG10_5_p & !v1445f88;
assign v144625a = hlock2 & v1446224 | !hlock2 & v1446258;
assign v121604a = hbusreq1 & v1216aad | !hbusreq1 & v845542;
assign v12ad626 = hbusreq5 & v12ad5fd | !hbusreq5 & v12ad625;
assign v1553508 = hlock5 & v15534f8 | !hlock5 & v1553507;
assign v1445e3d = hmaster2_p & v1445e38 | !hmaster2_p & v845542;
assign v12afa33 = hready_p & v12afa11 | !hready_p & v12afa32;
assign v1553389 = locked_p & v1553388 | !locked_p & v845542;
assign v16a1e73 = hbusreq2 & v16a1e70 | !hbusreq2 & v16a1e72;
assign v121502b = hgrant0_p & v12160f2 | !hgrant0_p & !v845542;
assign d2fe8e = hmaster2_p & d2fe7b | !hmaster2_p & d2fe84;
assign v1516215 = hgrant3_p & v15169a0 | !hgrant3_p & !v1516214;
assign v12157af = hbusreq4_p & v12157ae | !hbusreq4_p & v845542;
assign v1445818 = hlock2 & v14457f6 | !hlock2 & v1445817;
assign v16a13cb = hbusreq2 & v16a13ca | !hbusreq2 & !v16a205c;
assign v16a131b = hbusreq0_p & v845547 | !hbusreq0_p & v845542;
assign f2f432 = hgrant5_p & f2f385 | !hgrant5_p & !f2f431;
assign v15155fd = hbusreq0 & v1668da6 | !hbusreq0 & v845542;
assign v16a1cbb = hmaster1_p & v16a1c9b | !hmaster1_p & v16a1f96;
assign v1446112 = hlock3 & v1446109 | !hlock3 & v1446111;
assign v134d434 = hgrant2_p & v134d364 | !hgrant2_p & v134d433;
assign v1214c58 = hbusreq1 & v1215347 | !hbusreq1 & v121535e;
assign d3073f = hburst0 & d3073c | !hburst0 & d3073e;
assign v16a1bd9 = hgrant5_p & v845542 | !hgrant5_p & v16a1bcb;
assign v1215feb = hbusreq1 & v1216a61 | !hbusreq1 & v845542;
assign f2f44d = hbusreq5_p & f2f3c4 | !hbusreq5_p & !f2f44c;
assign v1284cf4 = hgrant4_p & v1284cf3 | !hgrant4_p & !v1405849;
assign v1214cdc = hbusreq0 & v1214cdb | !hbusreq0 & v845542;
assign v1446468 = stateG3_2_p & v845542 | !stateG3_2_p & !v845584;
assign a65370 = hbusreq4_p & a6536e | !hbusreq4_p & v845542;
assign v1405923 = hmaster0_p & v1405859 | !hmaster0_p & v14058b4;
assign d2f985 = hbusreq2_p & v84555a | !hbusreq2_p & d2f984;
assign a65405 = hmaster1_p & a65403 | !hmaster1_p & a653e7;
assign d306d4 = locked_p & v845542 | !locked_p & a65861;
assign a6537d = hlock0_p & v845570 | !hlock0_p & !v845542;
assign v134d453 = hbusreq2_p & v134d451 | !hbusreq2_p & v134d452;
assign v1446256 = hbusreq2_p & v1446254 | !hbusreq2_p & v1446255;
assign v1668cba = stateA1_p & v845542 | !stateA1_p & !a658a8;
assign v1215cce = hgrant5_p & v845542 | !hgrant5_p & !v1215c87;
assign v1445384 = hmaster1_p & v1445b40 | !hmaster1_p & v1445a82;
assign v1445fc0 = hbusreq2_p & v1445fbe | !hbusreq2_p & v1445fbf;
assign d2f991 = hlock4_p & v845542 | !hlock4_p & !d30957;
assign d2fba2 = hmaster1_p & d2fb86 | !hmaster1_p & d2fb9d;
assign v1214cee = hgrant5_p & v1214c2d | !hgrant5_p & v1214ced;
assign v121630d = hmaster0_p & v12162e8 | !hmaster0_p & v121630c;
assign d30793 = hgrant1_p & v845542 | !hgrant1_p & d30792;
assign d2fba9 = hbusreq2_p & d2fba8 | !hbusreq2_p & d2fba7;
assign d2faee = hmaster2_p & d2fae9 | !hmaster2_p & d2faed;
assign v1445923 = hbusreq2 & v1445921 | !hbusreq2 & v1445922;
assign v14461ef = hmaster1_p & v1446189 | !hmaster1_p & v14460cf;
assign d2fd2a = hmaster1_p & d2fd24 | !hmaster1_p & !d30293;
assign v1214bd8 = hbusreq2 & v1214bd3 | !hbusreq2 & v1214bd7;
assign v16a196e = hbusreq4_p & v845572 | !hbusreq4_p & v845542;
assign v10d40da = hbusreq2_p & v10d40d5 | !hbusreq2_p & v10d40d9;
assign d306d6 = hlock1_p & d306d5 | !hlock1_p & v845570;
assign v151576d = hbusreq0_p & v1668d25 | !hbusreq0_p & !v1515745;
assign f2e4cf = hbusreq0 & f2f51a | !hbusreq0 & f2f236;
assign d2fb14 = hgrant2_p & d3012a | !hgrant2_p & d2fad3;
assign v121481a = hgrant3_p & v1214f7e | !hgrant3_p & v1214819;
assign v1215dc1 = decide_p & v845542 | !decide_p & v12164e7;
assign v134cd5a = hgrant1_p & v134cd59 | !hgrant1_p & v845542;
assign v138a3d6 = hlock5_p & v138a3d3 | !hlock5_p & !v138a3d5;
assign v1446300 = hmaster1_p & v14465b7 | !hmaster1_p & v14462ff;
assign v16a1ad5 = hbusreq5 & v16a1ac8 | !hbusreq5 & !v16a1ad4;
assign v14453b7 = hmaster1_p & v1445a5a | !hmaster1_p & v1445a9b;
assign v1215754 = hbusreq0 & v121574a | !hbusreq0 & v1215753;
assign v1215c96 = hgrant5_p & v1215c92 | !hgrant5_p & v1215c95;
assign v134d3b3 = hmaster0_p & v134d379 | !hmaster0_p & v134d38b;
assign v1669596 = hmaster1_p & v1669595 | !hmaster1_p & v845570;
assign v1446605 = hgrant5_p & v14465ea | !hgrant5_p & v1446604;
assign v134d39b = hmaster1_p & v134d369 | !hmaster1_p & v134d39a;
assign v1446693 = hbusreq5_p & v144668e | !hbusreq5_p & v14465dd;
assign v1445b50 = hmaster1_p & v1445a3e | !hmaster1_p & v1445a61;
assign d807b0 = hmaster1_p & d807af | !hmaster1_p & !v845542;
assign v16a1969 = hmaster1_p & v16a1962 | !hmaster1_p & v16a1968;
assign v16a1e1f = hgrant0_p & v845547 | !hgrant0_p & !v16a1bc6;
assign v12164cf = hready & v845570 | !hready & !v845542;
assign v134d1db = stateG2_p & v845542 | !stateG2_p & v134d1da;
assign v16a1e96 = hbusreq1_p & v16a207f | !hbusreq1_p & v16a1e95;
assign v1445bbd = hready_p & v1445bac | !hready_p & v1445bbc;
assign v1405865 = hmaster2_p & v14463b1 | !hmaster2_p & v1405863;
assign f2f28b = hmaster1_p & f2f284 | !hmaster1_p & f2f28a;
assign v1445b57 = stateG10_5_p & v14465d3 | !stateG10_5_p & v1445b56;
assign v1215070 = hgrant2_p & v1215059 | !hgrant2_p & v121506f;
assign v1284ca2 = hbusreq5_p & v1284c9d | !hbusreq5_p & v1284ca1;
assign v121531d = decide_p & v1215302 | !decide_p & v121531c;
assign v16a1a26 = hmaster1_p & v16a19e0 | !hmaster1_p & !v16a1f96;
assign v14453f0 = hlock5 & v14453e4 | !hlock5 & v14453ee;
assign v1215ddc = hgrant3_p & v1215dc2 | !hgrant3_p & v1215ddb;
assign v1215112 = hready_p & v12150c0 | !hready_p & !v1215111;
assign d306da = hbusreq4_p & v845542 | !hbusreq4_p & d306d4;
assign v1668d76 = hbusreq0_p & v1668d24 | !hbusreq0_p & v1668d47;
assign v1405afc = hgrant1_p & v1405a88 | !hgrant1_p & !v1405a8c;
assign v14460d4 = hbusreq2_p & v14460d1 | !hbusreq2_p & v14460d3;
assign d2fd38 = hgrant3_p & d2fd1a | !hgrant3_p & d2fd37;
assign v151572e = hmaster2_p & v151572a | !hmaster2_p & v151572d;
assign v10d3ff2 = hmaster0_p & v10d3ff0 | !hmaster0_p & v10d3ff1;
assign v16a1a97 = hbusreq0 & v16a1a96 | !hbusreq0 & v845542;
assign v134d291 = hgrant1_p & v845542 | !hgrant1_p & v134d290;
assign d2fc84 = hmaster1_p & d2fc83 | !hmaster1_p & v845570;
assign v134d53b = decide_p & v134d3ce | !decide_p & v134d53a;
assign v16a1320 = hready & v16a131f | !hready & v845542;
assign v1216aec = hlock0_p & v1216ab9 | !hlock0_p & v845547;
assign v1668cfe = hmaster1_p & v1668cbf | !hmaster1_p & !v1668cfd;
assign v134d508 = hlock1 & v134d507 | !hlock1 & v134d503;
assign v12acfd3 = hmaster1_p & v12acfc4 | !hmaster1_p & !v12acfb9;
assign v16a1d31 = hmaster1_p & v16a2234 | !hmaster1_p & v16a1f96;
assign v1668d82 = hgrant4_p & v1668d70 | !hgrant4_p & a65382;
assign v14459f4 = hbusreq1_p & v144639c | !hbusreq1_p & v14459f3;
assign d2fb24 = hbusreq0 & d2fb21 | !hbusreq0 & d2fb23;
assign v1214f5b = hgrant2_p & v845542 | !hgrant2_p & v1214f5a;
assign v1516103 = hlock2_p & v1516102 | !hlock2_p & v845542;
assign v138980a = hbusreq5_p & v1389809 | !hbusreq5_p & !v845542;
assign v1515782 = hgrant5_p & v1515615 | !hgrant5_p & v1515781;
assign v1216adc = hready & v1446394 | !hready & !v1668cba;
assign v10d3fea = hmaster1_p & v10d3fdd | !hmaster1_p & v10d3fe9;
assign a65454 = hbusreq5 & a65412 | !hbusreq5 & a65452;
assign v1445e81 = hmaster2_p & v1445e80 | !hmaster2_p & v1445e7c;
assign v1445e70 = hbusreq1 & v1445e55 | !hbusreq1 & v1445e6f;
assign v14466ed = hbusreq3 & v14466eb | !hbusreq3 & v14466ec;
assign v12af5ac = hgrant5_p & v845542 | !hgrant5_p & v12af5ab;
assign v1445aaf = hgrant3_p & v144592a | !hgrant3_p & v1445aae;
assign v16695ca = jx0_p & v1668e10 | !jx0_p & v16695c9;
assign v16a1960 = hgrant5_p & v845542 | !hgrant5_p & !v16a1942;
assign v1446170 = hbusreq2_p & v1446165 | !hbusreq2_p & v144616f;
assign v134d1fa = hlock5_p & v134d1f3 | !hlock5_p & v134d1f9;
assign v16a1334 = hmaster1_p & v16a1333 | !hmaster1_p & !v16a2672;
assign v14459b1 = hlock0_p & v14459af | !hlock0_p & v14459b0;
assign bf1f73 = hbusreq2_p & bf1f71 | !hbusreq2_p & !bf1f72;
assign v1445f14 = hbusreq2_p & v1445f0b | !hbusreq2_p & v1445f13;
assign v121577c = hgrant5_p & v1215ba3 | !hgrant5_p & !v121577a;
assign v16a1d77 = hgrant5_p & v845542 | !hgrant5_p & !v16a1d6a;
assign d2fedf = hbusreq2_p & d2fede | !hbusreq2_p & d2fed9;
assign d30811 = hgrant2_p & d30810 | !hgrant2_p & d307f5;
assign v12ad535 = hmaster2_p & v12ad514 | !hmaster2_p & a658ca;
assign v14458ef = hbusreq0 & v14458ea | !hbusreq0 & v14458ee;
assign v155313a = hmaster0_p & v1553139 | !hmaster0_p & v845542;
assign v12150a9 = hmaster2_p & v121508d | !hmaster2_p & v121509b;
assign v12acfb6 = hmaster2_p & v12acfb5 | !hmaster2_p & !v12af985;
assign v1284d5c = hmaster1_p & v1284d5b | !hmaster1_p & !v1445bb7;
assign v14463db = hbusreq1_p & v144639c | !hbusreq1_p & v14463da;
assign v1405a89 = hmaster2_p & v1405a86 | !hmaster2_p & v1405a88;
assign d30843 = hbusreq2 & d3083f | !hbusreq2 & d30842;
assign d30860 = hbusreq2_p & v84554e | !hbusreq2_p & d3085f;
assign v166959a = hmaster1_p & v1669598 | !hmaster1_p & v1669599;
assign v121659e = hlock0_p & v1216a8d | !hlock0_p & v121659d;
assign v1552da2 = jx2_p & v1552d79 | !jx2_p & v1552da1;
assign v1446016 = hgrant5_p & v845542 | !hgrant5_p & v1446015;
assign a6470b = hmaster0_p & a66287 | !hmaster0_p & a65b13;
assign v1215c84 = hmaster1_p & v1215c7d | !hmaster1_p & v1215c83;
assign v134d36b = stateA1_p & v134d1e7 | !stateA1_p & v134d1e6;
assign v14460ff = hlock3 & v14460f4 | !hlock3 & v14460fe;
assign a662b9 = hgrant2_p & v845542 | !hgrant2_p & a662b8;
assign v138a010 = hbusreq3 & v138a008 | !hbusreq3 & v138a404;
assign f2f370 = hmaster2_p & f2f358 | !hmaster2_p & f2f234;
assign d3080d = hmaster1_p & d3080c | !hmaster1_p & d306f9;
assign v1214e0d = hmaster2_p & v1216ad6 | !hmaster2_p & v1214e0c;
assign v1215095 = hgrant4_p & v845542 | !hgrant4_p & v1215094;
assign f2f4a9 = hbusreq1_p & f2f4a8 | !hbusreq1_p & !v845542;
assign v12162b7 = hmaster0_p & f2f2a8 | !hmaster0_p & v12161f7;
assign v1445a58 = hgrant5_p & v1445907 | !hgrant5_p & v1445a57;
assign d3085c = hmaster2_p & d30654 | !hmaster2_p & !v845542;
assign v1405aa1 = stateA1_p & v1405aa0 | !stateA1_p & v845582;
assign v16a1974 = hgrant5_p & v845542 | !hgrant5_p & v16a1973;
assign v1445fdc = hmaster2_p & v1445fd4 | !hmaster2_p & v1445fdb;
assign v144623c = hbusreq2_p & v1446237 | !hbusreq2_p & v144623b;
assign v16a196f = hgrant4_p & v845559 | !hgrant4_p & !v16a196e;
assign a66278 = hbusreq4_p & a66276 | !hbusreq4_p & !v845542;
assign v15168fe = hbusreq2_p & v15168fd | !hbusreq2_p & !v845542;
assign v1214d1b = hgrant5_p & v1214d1a | !hgrant5_p & !v1214cf6;
assign v134d43e = hmaster2_p & v845542 | !hmaster2_p & v134d43d;
assign v1446726 = hmaster1_p & v1446725 | !hmaster1_p & v1446436;
assign v10d40a4 = decide_p & v10d409e | !decide_p & !v10d40a3;
assign v15167ff = hlock2_p & v845570 | !hlock2_p & !v845542;
assign v134d234 = hlock2_p & v134d233 | !hlock2_p & v134d22f;
assign bf1f5b = hgrant5_p & v845570 | !hgrant5_p & d3064a;
assign v10d3fd6 = stateA1_p & v845542 | !stateA1_p & !v88d3e4;
assign v12af225 = hgrant5_p & d30690 | !hgrant5_p & v12af224;
assign v11e596d = hgrant2_p & v11e5942 | !hgrant2_p & v11e596c;
assign v143fd7d = hgrant3_p & v143fd77 | !hgrant3_p & v143fd7c;
assign d307a5 = hbusreq5_p & d307a4 | !hbusreq5_p & !d307a3;
assign v1445798 = hlock2 & v1445786 | !hlock2 & v1445796;
assign v10d428a = hgrant4_p & v10d3fdb | !hgrant4_p & v10d4289;
assign v1446729 = hgrant2_p & v1446726 | !hgrant2_p & v1446728;
assign v134d44a = hmaster2_p & v134d43d | !hmaster2_p & v845542;
assign d3011d = hbusreq5_p & d3011c | !hbusreq5_p & !d3011b;
assign v16a2063 = hbusreq2 & v16a2062 | !hbusreq2 & v16a1f9b;
assign d300b4 = hlock2_p & d300b3 | !hlock2_p & !d2fea3;
assign v121537d = hmaster2_p & d2fbe5 | !hmaster2_p & v121537c;
assign v134d4fc = hgrant4_p & v134d4fb | !hgrant4_p & v845542;
assign v1446005 = hlock3 & v1445ff3 | !hlock3 & v1446004;
assign v10d403a = hgrant1_p & v10d4039 | !hgrant1_p & v10d4030;
assign v14460f0 = hmaster1_p & v14460ef | !hmaster1_p & v1445fae;
assign v1216a98 = hlock0_p & v16a1bc6 | !hlock0_p & v1216a97;
assign v16a1bf7 = hmaster1_p & v16a1bf2 | !hmaster1_p & v16a1bf6;
assign v14458bf = hbusreq0 & v1445878 | !hbusreq0 & v14458be;
assign v12166f8 = hmaster0_p & v12166c8 | !hmaster0_p & v12166f7;
assign bf1f81 = hgrant4_p & bf1f52 | !hgrant4_p & !v84556a;
assign v1405b5a = decide_p & v1405b54 | !decide_p & v1405b59;
assign d2fc50 = hbusreq0_p & v845570 | !hbusreq0_p & !v845542;
assign v12153fe = hbusreq2_p & v12153fd | !hbusreq2_p & v12153fc;
assign v12162e2 = hgrant3_p & v121627f | !hgrant3_p & !v12162e1;
assign v1216052 = hlock1_p & v1216050 | !hlock1_p & v1216051;
assign v12161ce = hbusreq1 & v1216587 | !hbusreq1 & v845542;
assign v1216102 = hgrant5_p & v1215ff2 | !hgrant5_p & v1216101;
assign v1216122 = hgrant0_p & v1216121 | !hgrant0_p & v1215ff6;
assign v1515840 = hbusreq2_p & v151583f | !hbusreq2_p & !v845542;
assign v134cee0 = hbusreq2_p & v134cedf | !hbusreq2_p & v134d276;
assign d30265 = hmaster0_p & v1668da6 | !hmaster0_p & v1668c17;
assign v1445800 = hbusreq2 & v14457ec | !hbusreq2 & v14457ff;
assign v144629b = hbusreq2 & v1446299 | !hbusreq2 & v144629a;
assign v1446079 = hlock0 & v1446078 | !hlock0 & v1446076;
assign v1405857 = hmaster0_p & v1405855 | !hmaster0_p & v1405856;
assign v1445ffa = hbusreq0 & v1445ff9 | !hbusreq0 & v1445fd1;
assign v1215d7a = hmaster1_p & v1215d6e | !hmaster1_p & v1215d79;
assign d3090d = hmaster2_p & d30718 | !hmaster2_p & d305ea;
assign v140590c = hmaster1_p & v140590b | !hmaster1_p & v140584d;
assign v12ad5c9 = hbusreq1 & v12ad4f6 | !hbusreq1 & v845542;
assign f2f446 = hbusreq5_p & f2f3d2 | !hbusreq5_p & !f2f445;
assign v1445ecb = hbusreq0 & v1445eca | !hbusreq0 & v1445eb8;
assign d300fe = hgrant1_p & d300fa | !hgrant1_p & d300fd;
assign v1446320 = hgrant5_p & v1446445 | !hgrant5_p & v144631f;
assign v134d500 = hbusreq0_p & v134d273 | !hbusreq0_p & v134d4e6;
assign v144663e = hbusreq1 & v14465c9 | !hbusreq1 & v144663d;
assign v14457cf = hlock3 & v1445786 | !hlock3 & v14457ce;
assign v1446050 = hmaster2_p & v144604f | !hmaster2_p & v14465db;
assign v1553217 = locked_p & v1553140 | !locked_p & v845542;
assign v144575e = hmaster1_p & v1445f35 | !hmaster1_p & v1445dd1;
assign v1446430 = hlock0_p & v1446403 | !hlock0_p & v144642f;
assign d307af = hlock4_p & d307ae | !hlock4_p & v1668d48;
assign v121538d = hbusreq2_p & v1215389 | !hbusreq2_p & v121538c;
assign v1445f71 = hgrant2_p & v1446747 | !hgrant2_p & v1445f70;
assign v12af58e = hgrant1_p & v845542 | !hgrant1_p & v12af58d;
assign f2f280 = hgrant3_p & f2f225 | !hgrant3_p & f2f27f;
assign v1215b8d = hbusreq2_p & v1215b89 | !hbusreq2_p & v1215b8c;
assign v16a13e6 = hmaster1_p & v16a13e5 | !hmaster1_p & v16a1d6d;
assign d30692 = hbusreq5_p & d305fd | !hbusreq5_p & d30691;
assign v1215cad = hgrant4_p & v12160f3 | !hgrant4_p & v845542;
assign v16a1d3d = hmaster2_p & v16a1d3c | !hmaster2_p & v16a208a;
assign v1214f54 = hmaster0_p & v1215d88 | !hmaster0_p & v1215d6c;
assign v1216552 = hlock4_p & v1216551 | !hlock4_p & v845547;
assign v16a267b = hmaster1_p & v16a2675 | !hmaster1_p & !v16a2672;
assign v10d404c = hgrant5_p & v10d3fe8 | !hgrant5_p & v10d404b;
assign v1445a00 = hlock1 & v14459cb | !hlock1 & v14459f8;
assign v1446662 = hbusreq0 & v1446661 | !hbusreq0 & v1446648;
assign v1284c98 = hmaster2_p & v140588d | !hmaster2_p & v1284c8e;
assign a65892 = hmaster2_p & v845542 | !hmaster2_p & a6587e;
assign v845568 = hmaster2_p & v845542 | !hmaster2_p & !v845542;
assign v144579a = hlock3 & v1445788 | !hlock3 & v1445799;
assign d301b1 = hbusreq2 & d301aa | !hbusreq2 & d301b0;
assign v1445fef = hmaster0_p & v1445fd1 | !hmaster0_p & v1445fd9;
assign v12ad0b6 = hbusreq1_p & v12afdab | !hbusreq1_p & v12afdac;
assign d301b8 = hlock3_p & d308fa | !hlock3_p & d301b7;
assign v1445b9b = hlock2 & v1445b92 | !hlock2 & v1445b95;
assign v16a1db8 = hbusreq5 & v16a1db7 | !hbusreq5 & v16a1aee;
assign v14460db = hlock2 & v14460a1 | !hlock2 & v14460da;
assign a658d6 = hlock0_p & a658b5 | !hlock0_p & a658d5;
assign a653f4 = hmaster1_p & a653ec | !hmaster1_p & a653f3;
assign d30137 = hbusreq0 & d30132 | !hbusreq0 & d30136;
assign v1216aa8 = hmastlock_p & v1216aa7 | !hmastlock_p & v845542;
assign v1553102 = hbusreq3 & v1553101 | !hbusreq3 & v155321a;
assign a6537a = hgrant5_p & a65360 | !hgrant5_p & a65378;
assign v1445f19 = hbusreq2 & v1445f15 | !hbusreq2 & v1445f18;
assign v121658f = hmastlock_p & v121658e | !hmastlock_p & !v845542;
assign v12ad13c = hlock2_p & v12aec0a | !hlock2_p & v12aec49;
assign v14466b1 = hmaster1_p & v14466b0 | !hmaster1_p & v14466a9;
assign v12150c5 = hbusreq1 & v12153d3 | !hbusreq1 & v12150c4;
assign v14458ac = hmaster1_p & v14458ab | !hmaster1_p & v144589f;
assign v10d4299 = hmaster2_p & v10d4298 | !hmaster2_p & !v10d4295;
assign v1445ea7 = hgrant5_p & v1445e05 | !hgrant5_p & v1445ea6;
assign v1515800 = hbusreq0 & v15157fd | !hbusreq0 & v15157ff;
assign v1215be2 = hmaster0_p & v1215be0 | !hmaster0_p & v1215be1;
assign v1445fea = hlock0 & v1445fe9 | !hlock0 & v1445fe8;
assign v1214c78 = hgrant5_p & v1215345 | !hgrant5_p & v1214c77;
assign v144673d = hmaster1_p & v1446648 | !hmaster1_p & v144666a;
assign v14459a6 = hmastlock_p & v14459a5 | !hmastlock_p & !v845542;
assign v12150f9 = hmaster0_p & v121543b | !hmaster0_p & v12150f8;
assign v1216227 = hmaster2_p & v12160d1 | !hmaster2_p & !v121620e;
assign v1446638 = hbusreq5_p & v144639c | !hbusreq5_p & v1446636;
assign d807a0 = hmaster0_p & v845542 | !hmaster0_p & d8079f;
assign v1214c17 = hmaster1_p & v1214c00 | !hmaster1_p & v1214bcf;
assign v16a1cca = hbusreq1_p & v16a1afa | !hbusreq1_p & !v845542;
assign v1445b76 = hgrant5_p & v1445b73 | !hgrant5_p & v1445b75;
assign v1446327 = hlock2 & v1446316 | !hlock2 & v1446326;
assign v14466a4 = hbusreq0 & v14466a3 | !hbusreq0 & v1446617;
assign v12acfe7 = hmaster1_p & v12acfce | !hmaster1_p & v12ad54f;
assign v12150f0 = hmaster1_p & v1215443 | !hmaster1_p & v12150ef;
assign v1445bca = decide_p & v1445bc9 | !decide_p & v1446564;
assign v1445eb9 = hbusreq0 & v1445eb5 | !hbusreq0 & v1445eb8;
assign v12150a3 = hmaster2_p & v845542 | !hmaster2_p & v12150a2;
assign v10d40ab = hmaster0_p & v10d3ffd | !hmaster0_p & v10d400e;
assign v121612e = hgrant4_p & v1216120 | !hgrant4_p & v845542;
assign v1405893 = hgrant5_p & v1405841 | !hgrant5_p & v1405892;
assign v144625d = hbusreq3 & v1446229 | !hbusreq3 & v144625c;
assign v906a5a = hburst0_p & v893df7 | !hburst0_p & v8a9c96;
assign v155350c = hready_p & v1553306 | !hready_p & v155350b;
assign v121607e = hmaster2_p & v1216067 | !hmaster2_p & v845542;
assign d30741 = hbusreq1 & d30740 | !hbusreq1 & v845542;
assign v12ad67a = hbusreq5_p & v12ad527 | !hbusreq5_p & v12ad679;
assign a65656 = hbusreq2_p & a65619 | !hbusreq2_p & a65655;
assign v1216588 = hgrant1_p & v845570 | !hgrant1_p & v1216587;
assign d2f97d = hmaster0_p & d2f978 | !hmaster0_p & d2f97c;
assign v12ad61d = hbusreq0 & v12ad61c | !hbusreq0 & v12afe63;
assign f2f2e6 = hbusreq1 & a658ca | !hbusreq1 & !v845542;
assign v14465d5 = hmaster2_p & v14465bb | !hmaster2_p & v1446412;
assign f2f34f = hbusreq1 & v10d3fd8 | !hbusreq1 & v845542;
assign v1214e40 = hmaster1_p & v1214e1a | !hmaster1_p & !v12163a9;
assign v1515807 = hbusreq5 & v15157d6 | !hbusreq5 & v1515806;
assign v12152f8 = hmaster1_p & v12157a4 | !hmaster1_p & v121579f;
assign bf1f7b = hgrant5_p & bf1f53 | !hgrant5_p & bf1f7a;
assign a658db = hburst0 & v845542 | !hburst0 & a658da;
assign v1215458 = hlock2_p & v1215456 | !hlock2_p & v1215457;
assign d307e9 = hgrant4_p & d307d3 | !hgrant4_p & d307e8;
assign v1216203 = hbusreq1 & v845542 | !hbusreq1 & v845547;
assign v1284d40 = decide_p & v1284d3f | !decide_p & !v1284cbf;
assign v14461b9 = hmaster1_p & v144616d | !hmaster1_p & v14460b6;
assign v1216708 = hmaster0_p & v1216702 | !hmaster0_p & v12166c8;
assign v1445f8c = hbusreq5_p & v1445f85 | !hbusreq5_p & v1445f8b;
assign v1668c64 = hbusreq1_p & v1668c62 | !hbusreq1_p & !v1668c63;
assign v14460c7 = hlock3 & v14460a1 | !hlock3 & v14460c6;
assign a65919 = hmaster1_p & a658ea | !hmaster1_p & !a65916;
assign f2f2a2 = hmaster0_p & f2f29c | !hmaster0_p & f2f2a1;
assign v1515778 = hbusreq5_p & v1515776 | !hbusreq5_p & v1515777;
assign v1216064 = hbusreq1 & v1216aea | !hbusreq1 & v845542;
assign d3065f = hlock5_p & v845542 | !hlock5_p & d3065e;
assign v12164c7 = hmaster1_p & v12164c6 | !hmaster1_p & v1216af8;
assign v1668de3 = hgrant2_p & v1668dad | !hgrant2_p & !v1668ddf;
assign v1445754 = hlock3 & v1445f42 | !hlock3 & v1445753;
assign v1445a11 = hlock0_p & v1445a0f | !hlock0_p & v1445a10;
assign f2f3d1 = hgrant2_p & f2f344 | !hgrant2_p & f2f3d0;
assign d308bf = hgrant5_p & d3085c | !hgrant5_p & d3089a;
assign v1445edf = hlock0 & v1445ede | !hlock0 & v1445edd;
assign v144538c = hbusreq2 & v1445387 | !hbusreq2 & v144538b;
assign v16a2678 = hbusreq2 & v16a2673 | !hbusreq2 & v16a2677;
assign v166939d = hmaster0_p & v166939c | !hmaster0_p & v845570;
assign v134d374 = hgrant1_p & v134d373 | !hgrant1_p & v845542;
assign v1668ce4 = hmaster2_p & v1668cd0 | !hmaster2_p & !v1668ce3;
assign v12ad326 = hgrant5_p & d30690 | !hgrant5_p & v12ad325;
assign v15157be = hlock0_p & v151561c | !hlock0_p & !v845542;
assign v16a1db3 = hgrant2_p & v845542 | !hgrant2_p & v16a1db2;
assign v10d4048 = hgrant0_p & v10d4047 | !hgrant0_p & v10d3ff9;
assign v121571e = hlock4_p & v121571c | !hlock4_p & v121571d;
assign v1214cb9 = hmaster0_p & v121537e | !hmaster0_p & v121537b;
assign v1215c00 = hbusreq5_p & v1215bfe | !hbusreq5_p & !v1215bff;
assign a662bb = decide_p & a662ba | !decide_p & a662a2;
assign d301ef = hgrant5_p & d301c6 | !hgrant5_p & d301ed;
assign v14463ce = hmaster1_p & v144639c | !hmaster1_p & v14463cd;
assign v1445a9d = hgrant2_p & v1445a74 | !hgrant2_p & v1445a9c;
assign v16a1e6f = hmaster1_p & v16a1e5f | !hmaster1_p & !v16a1f96;
assign d2f998 = hlock2_p & d2f996 | !hlock2_p & d2f997;
assign v12ad521 = hbusreq0_p & v1668c6c | !hbusreq0_p & v845542;
assign v12ad4fd = hmaster2_p & v12ad4fc | !hmaster2_p & v845542;
assign v1214db7 = hgrant2_p & v1214da8 | !hgrant2_p & v1214db6;
assign v16a2671 = hbusreq0 & v16a266f | !hbusreq0 & v16a2670;
assign v134d395 = hmaster2_p & v134d383 | !hmaster2_p & v134d394;
assign f2f3c8 = hgrant5_p & f2f2a8 | !hgrant5_p & !f2f37f;
assign d3088b = hmaster2_p & d30888 | !hmaster2_p & d3088a;
assign v14459ef = hgrant5_p & v14459ea | !hgrant5_p & v14459ee;
assign v144576a = hmaster1_p & v1445db8 | !hmaster1_p & v1445dd1;
assign v16a1a96 = hmaster2_p & v16a1a92 | !hmaster2_p & v845542;
assign v1445810 = hmaster1_p & v1445ecc | !hmaster1_p & v1445eaa;
assign v1668c1a = hmaster1_p & v1668c19 | !hmaster1_p & v845570;
assign v1405b28 = hgrant5_p & v1405ac7 | !hgrant5_p & v1405b27;
assign v1214ee5 = hgrant5_p & v1216a5a | !hgrant5_p & v121655a;
assign v1445a2a = hgrant4_p & v1445a25 | !hgrant4_p & v1445a29;
assign v1445fa6 = hbusreq1_p & v14463a2 | !hbusreq1_p & v144639e;
assign v10d4063 = hmaster2_p & v10d405f | !hmaster2_p & v10d4062;
assign v15157ed = hgrant5_p & v15157e7 | !hgrant5_p & !v1515758;
assign v1668c37 = hready_p & v845542 | !hready_p & v1668c36;
assign d30661 = hgrant4_p & d30660 | !hgrant4_p & v845542;
assign d3066e = hmaster1_p & d3064d | !hmaster1_p & d3066d;
assign d30276 = hgrant5_p & d30274 | !hgrant5_p & d30275;
assign v1214c5e = hgrant5_p & v1214c57 | !hgrant5_p & v1214c5d;
assign v1215c67 = hgrant5_p & v845542 | !hgrant5_p & v1215c2a;
assign v12ad5c2 = hgrant4_p & v12ad5c0 | !hgrant4_p & !v12ad5c1;
assign v1215086 = hgrant2_p & v1215024 | !hgrant2_p & v1215085;
assign v14453e8 = hlock3 & v14453e4 | !hlock3 & v14453e7;
assign v12160aa = hlock2_p & v12160a7 | !hlock2_p & v12160a9;
assign v134ce9a = hbusreq5_p & v134ce99 | !hbusreq5_p & v134d1fd;
assign v1445405 = hgrant5_p & v1445404 | !hgrant5_p & v1446472;
assign v12161f3 = hgrant5_p & v1216040 | !hgrant5_p & v12161f2;
assign v1284cff = hgrant2_p & v1284cc3 | !hgrant2_p & v1284cfe;
assign v12150ee = hbusreq5_p & v12150ed | !hbusreq5_p & v12150c9;
assign v16a1aeb = hbusreq2_p & v16a209d | !hbusreq2_p & v16a1aea;
assign d80753 = hburst0_p & v845542 | !hburst0_p & !v84556c;
assign f2f539 = hgrant5_p & v845542 | !hgrant5_p & !f2f538;
assign v1445767 = hmaster1_p & v1445f47 | !hmaster1_p & v1445dd1;
assign v16a19b7 = hgrant2_p & v16a205b | !hgrant2_p & v16a19b6;
assign v12166fe = hmaster0_p & v12164d7 | !hmaster0_p & v12166fd;
assign v1215436 = hbusreq4 & v1216048 | !hbusreq4 & v1215435;
assign v1405b62 = hbusreq2_p & v1405b5f | !hbusreq2_p & v1405b61;
assign v15533a2 = hgrant1_p & v845542 | !hgrant1_p & v15533a1;
assign v121631e = hlock2_p & v121631c | !hlock2_p & v121631d;
assign d30607 = hbusreq0 & d305ff | !hbusreq0 & d30606;
assign v1445e90 = hgrant1_p & v1445dfe | !hgrant1_p & v1445e8f;
assign v1668d07 = hbusreq2_p & v1668cfe | !hbusreq2_p & v1668d06;
assign v121531b = hgrant2_p & v1215319 | !hgrant2_p & v121531a;
assign v14463ca = hmaster0_p & v144639c | !hmaster0_p & v14463c9;
assign v1215c33 = hbusreq5_p & v1215c31 | !hbusreq5_p & v1215c32;
assign d2fea4 = hmaster2_p & d2fe9a | !hmaster2_p & !d2fe9c;
assign f2e713 = hgrant1_p & f2e712 | !hgrant1_p & !v845542;
assign v1445b09 = hlock2 & v1445b05 | !hlock2 & v1445b08;
assign v1445e52 = decide_p & v1445e51 | !decide_p & v1446564;
assign v1445a13 = hbusreq4_p & v14465b1 | !hbusreq4_p & v1445a12;
assign v121605d = hmaster0_p & v121604f | !hmaster0_p & v121605c;
assign v121618f = hmaster2_p & v1216017 | !hmaster2_p & v845542;
assign v1215378 = hready & v1215377 | !hready & v845542;
assign v12161d4 = hmaster2_p & v1216034 | !hmaster2_p & v845542;
assign d8079d = hmaster1_p & d8076f | !hmaster1_p & !d8079c;
assign v121623b = hbusreq2 & v121622f | !hbusreq2 & v121623a;
assign v144591c = hmaster1_p & v14458d5 | !hmaster1_p & v144591b;
assign v1445acb = hbusreq2 & v1445ac9 | !hbusreq2 & v1445aca;
assign v14463a1 = hlock1 & v144639c | !hlock1 & v14463a0;
assign d8073b = hmaster2_p & d8073a | !hmaster2_p & d80732;
assign v14463be = hmaster2_p & v144639c | !hmaster2_p & v14463b5;
assign v1215c8f = hgrant5_p & v845542 | !hgrant5_p & !v1215c8d;
assign v134d4cf = hmaster2_p & v134d4ca | !hmaster2_p & v845542;
assign v1215109 = hbusreq2 & v12150f3 | !hbusreq2 & v1215108;
assign v14460b1 = stateG10_5_p & v1446041 | !stateG10_5_p & v14460b0;
assign v1389f87 = hmaster1_p & v845542 | !hmaster1_p & !v1389f86;
assign v1515732 = hbusreq0 & v1515727 | !hbusreq0 & v1515731;
assign v1516998 = hmaster2_p & v845542 | !hmaster2_p & v16693aa;
assign d2fae7 = hgrant4_p & v845558 | !hgrant4_p & d2fae6;
assign d3014d = hbusreq0 & d30148 | !hbusreq0 & d3014c;
assign v138a02c = hgrant5_p & v138a02b | !hgrant5_p & v845542;
assign v12ad55c = hmaster1_p & v12ad52d | !hmaster1_p & v12ad54f;
assign v1284c9c = hmaster2_p & v14463b1 | !hmaster2_p & !v1284c9a;
assign v138a3ad = hbusreq2 & v138a3a5 | !hbusreq2 & v138a3ac;
assign v114a232 = hgrant5_p & v845542 | !hgrant5_p & !v114a231;
assign v14459c3 = hlock4 & v144639c | !hlock4 & v14465ad;
assign v1214d9e = hmaster0_p & v1214ce0 | !hmaster0_p & v1214cc1;
assign v144672e = hbusreq2_p & v1446729 | !hbusreq2_p & v144672d;
assign v14058ea = hgrant1_p & v140587c | !hgrant1_p & v14058e9;
assign f2f394 = hmaster1_p & f2f35d | !hmaster1_p & f2f393;
assign v14058a4 = hgrant5_p & v14058a2 | !hgrant5_p & v14058a3;
assign d2fe9c = hlock4_p & a65861 | !hlock4_p & !v845542;
assign v10d4080 = hmaster0_p & v10d3fdc | !hmaster0_p & v10d407f;
assign v16a1326 = hgrant1_p & v845542 | !hgrant1_p & v16a1325;
assign v16a208c = hbusreq5_p & v16a2088 | !hbusreq5_p & v16a208b;
assign v121572d = hgrant5_p & v1215b7e | !hgrant5_p & v121572c;
assign v1445fb3 = hlock2 & v1445fb2 | !hlock2 & v1445fac;
assign v144671e = hbusreq3 & v1446711 | !hbusreq3 & v144671d;
assign v134d45d = hready_p & v134d34f | !hready_p & v134d45c;
assign f2f346 = hbusreq1_p & f2f345 | !hbusreq1_p & v845542;
assign v1405b0c = hmaster1_p & v1405af8 | !hmaster1_p & v1405b09;
assign v16a143e = hgrant2_p & v845542 | !hgrant2_p & !v16a143c;
assign v144661e = hlock1 & v1446600 | !hlock1 & v144661d;
assign v1552f7c = hbusreq0 & v1552f7b | !hbusreq0 & v1553395;
assign v1405aee = hmaster2_p & v1405ae8 | !hmaster2_p & v1405aed;
assign v1216793 = hmaster1_p & v1216792 | !hmaster1_p & v1216a9b;
assign v1214f57 = hbusreq2_p & v1214f56 | !hbusreq2_p & v12164e7;
assign v121624d = hgrant2_p & v1216202 | !hgrant2_p & v121624c;
assign d2fc5f = hgrant1_p & d2fbdf | !hgrant1_p & d2fc55;
assign v14461bf = hbusreq2_p & v144619e | !hbusreq2_p & v14461be;
assign v1405912 = hlock0_p & v1405860 | !hlock0_p & v1405911;
assign v134d1f5 = hgrant4_p & v134d1f4 | !hgrant4_p & v134d1e8;
assign v1445902 = hlock0 & v1445901 | !hlock0 & v14458ff;
assign v14459bb = hlock0_p & v144640c | !hlock0_p & v14459ba;
assign v12ad0bd = hbusreq2_p & v12ad0bc | !hbusreq2_p & v12afe3d;
assign f2f32a = hbusreq2_p & f2f327 | !hbusreq2_p & f2f329;
assign d2fd43 = hready_p & d2fd3b | !hready_p & d2fd42;
assign v1445457 = hmaster1_p & v1445443 | !hmaster1_p & v1446250;
assign d300de = hbusreq1_p & d300c3 | !hbusreq1_p & d300dd;
assign v1552963 = hbusreq3_p & v15530f5 | !hbusreq3_p & v1552962;
assign v1553413 = hmaster2_p & v845542 | !hmaster2_p & v1553412;
assign v14460aa = hlock2 & v14460a1 | !hlock2 & v14460a9;
assign d2fbfd = hmaster0_p & d2fbf2 | !hmaster0_p & d2fbfc;
assign v1445fcf = hbusreq1_p & v1446407 | !hbusreq1_p & v1446406;
assign v1215782 = hbusreq2_p & v1215772 | !hbusreq2_p & !v1215781;
assign v121613d = hbusreq4_p & v121613c | !hbusreq4_p & !v845542;
assign v1215ff3 = hmaster0_p & v1215ff0 | !hmaster0_p & v1215ff2;
assign v1284ca9 = hmaster2_p & v140588d | !hmaster2_p & !v14463b1;
assign v1445aff = hbusreq2 & v1445afd | !hbusreq2 & v1445afe;
assign a654ac = hbusreq3 & a65492 | !hbusreq3 & a654ab;
assign v12160dd = hbusreq1 & v12164de | !hbusreq1 & v845542;
assign v16a1ca7 = hmaster1_p & v16a1c9f | !hmaster1_p & !v16a2672;
assign v1216703 = hmaster0_p & v12166c8 | !hmaster0_p & v1216702;
assign v1552d4c = hmaster0_p & v1552d48 | !hmaster0_p & v1552d4b;
assign v10d40c0 = hbusreq1_p & v10d401d | !hbusreq1_p & v10d40bf;
assign v1214da1 = hmaster0_p & v121538a | !hmaster0_p & v1214cdc;
assign v12ad667 = hmaster1_p & v12ad662 | !hmaster1_p & v12ad666;
assign v11f33c6 = jx1_p & v11f33c5 | !jx1_p & v8b6f6c;
assign v16a224e = hmaster1_p & v16a2246 | !hmaster1_p & !v16a2672;
assign v16a1ce5 = hbusreq2 & v16a1ce2 | !hbusreq2 & v16a1ce4;
assign v1446008 = hlock5 & v1445ff3 | !hlock5 & v1446006;
assign v134d4c7 = hbusreq3_p & v134d4bc | !hbusreq3_p & v134d4c6;
assign v144535d = hlock2 & v1445354 | !hlock2 & v1445358;
assign v8b8a8c = stateG2_p & v845542 | !stateG2_p & v936735;
assign d2fd3c = hbusreq2_p & d2fd10 | !hbusreq2_p & d302da;
assign d30748 = hmaster1_p & d30747 | !hmaster1_p & d3072c;
assign v1446103 = hmaster1_p & v1445fa2 | !hmaster1_p & v1445fbd;
assign v1216235 = hmaster2_p & v1216207 | !hmaster2_p & v12161da;
assign d3082e = hbusreq5_p & d3082d | !hbusreq5_p & d3082c;
assign v1214df7 = hbusreq5_p & v1214df6 | !hbusreq5_p & v1214df5;
assign v12ad5b8 = hbusreq1 & a653c8 | !hbusreq1 & !v12ad506;
assign v134ceb8 = hmaster1_p & v134d20a | !hmaster1_p & v134ce9d;
assign v1445ae2 = hlock5 & v1445ace | !hlock5 & v1445ae1;
assign v155351a = hgrant3_p & v1553517 | !hgrant3_p & v1553519;
assign v10d427a = stateG2_p & v88d3e4 | !stateG2_p & !v10d4264;
assign v16a1e50 = hmaster1_p & v16a1e2c | !hmaster1_p & v16a1f96;
assign v1216abb = hgrant4_p & v1216aba | !hgrant4_p & v1216ab8;
assign v1445dc3 = hmaster1_p & v144639c | !hmaster1_p & v1445dc2;
assign a65b12 = hmaster2_p & a66286 | !hmaster2_p & a6628b;
assign f2f34a = hbusreq1 & v1668d35 | !hbusreq1 & v845542;
assign v14453bd = hlock2 & v1445354 | !hlock2 & v14453bc;
assign v121617e = hmaster0_p & v1216116 | !hmaster0_p & v121617d;
assign v14453a7 = hmaster1_p & v1445a43 | !hmaster1_p & v1445a9b;
assign a65691 = hmaster0_p & a658f1 | !hmaster0_p & a658ee;
assign v1216016 = hlock1_p & v1216012 | !hlock1_p & v1216015;
assign v1445bc3 = hmaster0_p & v1445bc2 | !hmaster0_p & v144649f;
assign v140592d = hgrant1_p & v1405889 | !hgrant1_p & v140592c;
assign v1445d80 = hbusreq4_p & v1445d7f | !hbusreq4_p & v144639e;
assign a6586a = hbusreq0_p & a65851 | !hbusreq0_p & a65862;
assign v12166df = hmaster2_p & v12166d9 | !hmaster2_p & v12166de;
assign v12160c6 = hbusreq2_p & v12160c5 | !hbusreq2_p & v12160c4;
assign d2fcb2 = hlock5_p & d2fcb0 | !hlock5_p & !d2fcb1;
assign v1445b44 = hlock2 & v1445b3d | !hlock2 & v1445b43;
assign v138a440 = hbusreq2_p & v138a438 | !hbusreq2_p & v138a43f;
assign v1445f86 = hbusreq1 & v14463a0 | !hbusreq1 & v14463f1;
assign v1405843 = stateA1_p & v845542 | !stateA1_p & v845588;
assign v134d4a5 = hlock2 & v134d49c | !hlock2 & v134d4a4;
assign v1216525 = hlock0_p & v1216a5a | !hlock0_p & v845547;
assign v1215038 = hgrant4_p & v845542 | !hgrant4_p & v1215037;
assign v1445885 = hbusreq1_p & v144639c | !hbusreq1_p & v1445884;
assign v1214c65 = hbusreq0 & v1214c64 | !hbusreq0 & v845542;
assign v1214f05 = hgrant5_p & v1215c5b | !hgrant5_p & v1214eda;
assign d30105 = hbusreq4_p & d30104 | !hbusreq4_p & v845542;
assign f2f399 = hbusreq1 & a65861 | !hbusreq1 & !v845542;
assign v14461c2 = hmaster1_p & v1446182 | !hmaster1_p & v1445ffc;
assign v1214d55 = hmaster0_p & v1214d50 | !hmaster0_p & v12153ab;
assign v16a1d46 = hbusreq0 & v16a207a | !hbusreq0 & v16a1d45;
assign v16a13de = hbusreq0 & v16a2071 | !hbusreq0 & v16a13dd;
assign v16a1cf3 = hgrant2_p & v845542 | !hgrant2_p & !v16a1cf0;
assign v155314c = hlock0_p & v1553140 | !hlock0_p & v845542;
assign v1214daf = hgrant2_p & v1214dad | !hgrant2_p & v1214dae;
assign f2e3fb = hgrant2_p & v845542 | !hgrant2_p & f2e3fa;
assign v16a1b64 = hmaster1_p & v16a1afb | !hmaster1_p & !v16a1f96;
assign v14453c3 = hbusreq5 & v14453a4 | !hbusreq5 & v14453c2;
assign v14459de = hbusreq1 & v14459c2 | !hbusreq1 & v14459dd;
assign f2f335 = hmaster1_p & f2f2e9 | !hmaster1_p & !f2f330;
assign v11e5971 = decide_p & bf1f4f | !decide_p & v11e593d;
assign v1215cdd = hgrant2_p & v1215cdc | !hgrant2_p & v1215cc9;
assign d30725 = hbusreq1_p & d30724 | !hbusreq1_p & v845542;
assign v16a1e20 = hgrant4_p & v845547 | !hgrant4_p & v16a1e1f;
assign v15168f6 = hbusreq1 & d305de | !hbusreq1 & d30645;
assign v14466be = hlock3 & v1446676 | !hlock3 & v14466bd;
assign v1445447 = hmaster0_p & v1446239 | !hmaster0_p & v144639c;
assign v144660e = hgrant4_p & v1446429 | !hgrant4_p & v144660d;
assign f2f354 = hbusreq1_p & f2f353 | !hbusreq1_p & v845542;
assign v14457eb = hbusreq2_p & v14457dc | !hbusreq2_p & v14457ea;
assign v12ad01c = hmaster0_p & v12ad661 | !hmaster0_p & v12ad660;
assign v16a1b65 = hmaster1_p & v16a1afe | !hmaster1_p & !v16a1f96;
assign v16a1bbe = hgrant1_p & v84554d | !hgrant1_p & v16a1bbd;
assign f2f288 = hgrant5_p & v845542 | !hgrant5_p & !f2f287;
assign v1389fba = hmaster0_p & v1389fb9 | !hmaster0_p & v845542;
assign v134d4a8 = hbusreq3 & v134d4a7 | !hbusreq3 & v134d3b5;
assign f2f3d8 = hbusreq0 & f2f3d4 | !hbusreq0 & f2f3d7;
assign v138a07f = decide_p & v138a07e | !decide_p & v138a406;
assign v138a365 = hbusreq2 & v138a35d | !hbusreq2 & v138a364;
assign v1215475 = decide_p & v121545d | !decide_p & v1215474;
assign d306f7 = hmaster2_p & d306d0 | !hmaster2_p & !d306f6;
assign v1215c41 = hmaster2_p & v1215bf6 | !hmaster2_p & v1215c1f;
assign hmastlock = bf1fab;
assign v134d445 = hlock2 & v134d434 | !hlock2 & v134d444;
assign v10d409c = hmaster0_p & v10d4052 | !hmaster0_p & v10d3ffd;
assign v16a1381 = hready_p & v16a12f9 | !hready_p & !v16a1380;
assign d30782 = hlock4_p & d30780 | !hlock4_p & !d30781;
assign v121620d = hbusreq1 & v12166ce | !hbusreq1 & !v845542;
assign v12ad567 = hmaster1_p & v12ad566 | !hmaster1_p & !v12ad525;
assign v1446049 = hmaster2_p & v1446048 | !hmaster2_p & v14465db;
assign v1445365 = hmaster1_p & v1445364 | !hmaster1_p & v14458fd;
assign v1215021 = hbusreq2_p & v1215018 | !hbusreq2_p & v1215020;
assign v14460c2 = hmaster1_p & v14460a6 | !hmaster1_p & v1445ffc;
assign v1214ca1 = hbusreq2 & v1214c9a | !hbusreq2 & v1214ca0;
assign v1215bf6 = hgrant1_p & v1215bf0 | !hgrant1_p & v1216105;
assign v14458fe = hmaster1_p & v14458d5 | !hmaster1_p & v14458fd;
assign f2f2d5 = hbusreq1_p & f2f2d4 | !hbusreq1_p & v845542;
assign v12ad00f = hbusreq4_p & v12ad5ae | !hbusreq4_p & v12ad000;
assign v1445ac7 = hmaster1_p & v14458aa | !hmaster1_p & v144589f;
assign v16a1d50 = hgrant2_p & v845542 | !hgrant2_p & !v16a1d4c;
assign v121570e = hbusreq1_p & v121570c | !hbusreq1_p & !v121570d;
assign v1216253 = hbusreq2_p & v1216252 | !hbusreq2_p & v121624f;
assign v1668d56 = hgrant5_p & v1668d50 | !hgrant5_p & !v1668d55;
assign v1215d8a = hmaster1_p & v1215d89 | !hmaster1_p & v1215d79;
assign a6538a = hmaster2_p & a65381 | !hmaster2_p & a65389;
assign v134cd69 = hbusreq0 & v134cd68 | !hbusreq0 & v134d38b;
assign v134ce61 = hbusreq0 & v134ce60 | !hbusreq0 & v134d379;
assign a653cf = hgrant4_p & v845570 | !hgrant4_p & !a653cd;
assign f2e3f8 = hbusreq5_p & f2e731 | !hbusreq5_p & f2e3f7;
assign v1445ddb = hlock2 & v1445dc6 | !hlock2 & v1445dd9;
assign d300cc = hgrant4_p & v845542 | !hgrant4_p & d300cb;
assign v1214c4e = hbusreq1 & v1215364 | !hbusreq1 & v845542;
assign v1389451 = hbusreq2_p & v1389450 | !hbusreq2_p & v138a391;
assign d2fc8f = decide_p & d2fc8e | !decide_p & v845570;
assign v14466db = hbusreq2_p & v14466d9 | !hbusreq2_p & v14466da;
assign v1445368 = hgrant2_p & v1445365 | !hgrant2_p & v1445367;
assign v1214c88 = hbusreq0 & v1214c87 | !hbusreq0 & v845542;
assign v1216195 = hlock5_p & v1216194 | !hlock5_p & v121612c;
assign v12ad595 = hready_p & v12ad50d | !hready_p & !v12ad594;
assign v1445a07 = hbusreq0 & v14459e3 | !hbusreq0 & v1445a06;
assign v12afe3b = hbusreq0 & v12afda4 | !hbusreq0 & v12afdb1;
assign v1668d90 = hmaster2_p & v10d3fd8 | !hmaster2_p & v1668d4f;
assign v14463a4 = hmaster2_p & v144639c | !hmaster2_p & v14463a3;
assign v134cd7d = hbusreq5_p & v134cd5c | !hbusreq5_p & v134cd7c;
assign v1552fd2 = hbusreq5 & v1552fd0 | !hbusreq5 & v1552fd1;
assign v121657e = hlock2_p & v121657b | !hlock2_p & v121657d;
assign v12ad005 = hmaster2_p & v12acffe | !hmaster2_p & v12ad004;
assign v10d400b = hmaster2_p & v10d3fd4 | !hmaster2_p & !v10d3fdb;
assign f2f362 = hbusreq1_p & f2f361 | !hbusreq1_p & !v845542;
assign v16a1bef = hbusreq1_p & v16a1bee | !hbusreq1_p & v16a2089;
assign v134d34f = decide_p & v134d309 | !decide_p & v134d316;
assign v144648a = hmaster2_p & v144647f | !hmaster2_p & v1446485;
assign d301e5 = hmaster0_p & d301dd | !hmaster0_p & d301e4;
assign v134d27c = hgrant0_p & v845542 | !hgrant0_p & v134d1dd;
assign v14460cc = hbusreq5_p & v1446042 | !hbusreq5_p & v14460cb;
assign v1515740 = hlock1_p & v151573e | !hlock1_p & v151573f;
assign v1284cc0 = decide_p & v1284cb8 | !decide_p & !v1284cbf;
assign f2f23b = hgrant5_p & v845542 | !hgrant5_p & !v845574;
assign v1445af7 = hmaster0_p & v1445a4f | !hmaster0_p & v1445902;
assign d2fb2c = hgrant2_p & d2fad6 | !hgrant2_p & !d2fb2b;
assign a658e5 = hmaster0_p & a658d1 | !hmaster0_p & !a658e3;
assign v144619d = hmaster1_p & v1446163 | !hmaster1_p & v14460b6;
assign v10d40d6 = hmaster0_p & v10d400e | !hmaster0_p & v10d3ffd;
assign v144604d = hmaster2_p & v14465d9 | !hmaster2_p & v1446412;
assign v144613f = hlock3 & v1446125 | !hlock3 & v144613e;
assign v14458b4 = hlock2 & v14458b3 | !hlock2 & v14458ad;
assign v1668da5 = hbusreq2_p & v1668d8d | !hbusreq2_p & v1668da4;
assign v1215d3c = hgrant2_p & v1215d2c | !hgrant2_p & v1215d3b;
assign v84555e = hlock5_p & v845542 | !hlock5_p & !v845542;
assign v1214bd0 = hmaster1_p & v1215396 | !hmaster1_p & v1214bcf;
assign v1445ea1 = hbusreq4_p & v1446626 | !hbusreq4_p & v144660d;
assign v1389de5 = hgrant5_p & v1389de4 | !hgrant5_p & !v845542;
assign v138a3da = hlock5_p & v138a3d9 | !hlock5_p & !v15157c2;
assign v134d26a = hbusreq2 & v134d260 | !hbusreq2 & v134d269;
assign d2fb94 = hmaster1_p & d2fb93 | !hmaster1_p & d2fb7b;
assign v12ad0cb = decide_p & v12ad0ca | !decide_p & v845542;
assign v1445f58 = hbusreq2_p & v144674a | !hbusreq2_p & v1445f57;
assign v1214e81 = hlock2_p & v1214e7f | !hlock2_p & !v1214e80;
assign v16a2090 = hbusreq5_p & v16a208f | !hbusreq5_p & v16a208b;
assign a6561c = hmaster1_p & a6561a | !hmaster1_p & a653f3;
assign v121532b = hmaster1_p & v121532a | !hmaster1_p & v1215054;
assign v1284d3e = hmaster1_p & v1284d3d | !hmaster1_p & v1284ca7;
assign v1215fb2 = hmaster1_p & v12167af | !hmaster1_p & v12164e1;
assign d308ca = hbusreq2_p & d308b7 | !hbusreq2_p & !d308c9;
assign v1446455 = hbusreq2_p & v144644e | !hbusreq2_p & v1446450;
assign v1445d97 = hlock0_p & v144639c | !hlock0_p & !v1445d96;
assign v138a482 = hgrant2_p & v138a3f5 | !hgrant2_p & !v138a47b;
assign v134d3ab = hbusreq5_p & v134d3aa | !hbusreq5_p & v134d274;
assign v12152e7 = hmaster1_p & v12152e6 | !hmaster1_p & !v1215ba1;
assign v144669b = hbusreq1 & v1446699 | !hbusreq1 & v144669a;
assign d3087d = hmaster0_p & d306e6 | !hmaster0_p & d306ce;
assign v10d40a0 = hmaster1_p & v10d409f | !hmaster1_p & v10d3fe9;
assign a654c5 = hbusreq3 & a654b9 | !hbusreq3 & a654c3;
assign v1668c9e = hmaster2_p & a65469 | !hmaster2_p & !v1668c77;
assign v1445f60 = hlock3 & v1446745 | !hlock3 & v1445f5f;
assign v1445533 = hlock3 & v144552e | !hlock3 & v1445532;
assign v121608d = hmaster1_p & v1216073 | !hmaster1_p & v1216082;
assign d306fb = hbusreq3 & d306e9 | !hbusreq3 & d306fa;
assign v1445dd9 = hbusreq2_p & v1445dd2 | !hbusreq2_p & v1445dd8;
assign d807a6 = hmaster1_p & d807a5 | !hmaster1_p & !v845542;
assign v1445914 = hbusreq2 & v144590d | !hbusreq2 & v1445913;
assign v1445e33 = hlock5 & v1445e23 | !hlock5 & v1445e32;
assign v1214d54 = hbusreq2 & v1214d4d | !hbusreq2 & v1214d53;
assign v1552d97 = decide_p & v1553216 | !decide_p & v155341e;
assign v1284d17 = hbusreq5_p & v1284d12 | !hbusreq5_p & v1284d16;
assign v12157a7 = hgrant2_p & v1215775 | !hgrant2_p & !v12157a6;
assign v16a1a8d = decide_p & v16a1a8c | !decide_p & v16a1984;
assign d2fd20 = hgrant5_p & v1668da6 | !hgrant5_p & d2fd1f;
assign v138980f = hlock5_p & v138980e | !hlock5_p & !v845542;
assign v1405909 = hmaster1_p & v1405908 | !hmaster1_p & v140584d;
assign v134cf40 = hready_p & v134d3e5 | !hready_p & v134cf3f;
assign v144608a = hlock0 & v1446089 | !hlock0 & v1446088;
assign v1445388 = hmaster1_p & v1445355 | !hmaster1_p & v144591b;
assign v16a1983 = hbusreq2 & v16a1981 | !hbusreq2 & !v16a1982;
assign v15157a7 = hbusreq1 & v151561c | !hbusreq1 & v1515630;
assign d30753 = hbusreq5_p & d30752 | !hbusreq5_p & v84554e;
assign v12157a0 = hmaster1_p & v121578e | !hmaster1_p & v121579f;
assign v12166ea = hgrant1_p & v12164de | !hgrant1_p & v12166e9;
assign a65ae2 = hbusreq1_p & a66285 | !hbusreq1_p & a662aa;
assign v1214ed9 = hmaster2_p & v1216a61 | !hmaster2_p & v1216a5a;
assign v1668dd7 = hgrant5_p & v845570 | !hgrant5_p & v1668d98;
assign d2f9a5 = hbusreq1_p & d2f992 | !hbusreq1_p & d2f9a4;
assign v1668c3b = hbusreq1_p & a66295 | !hbusreq1_p & v845570;
assign v14454f2 = hgrant2_p & v14454e9 | !hgrant2_p & v14454f1;
assign v138a2f8 = hbusreq5_p & v138a2f7 | !hbusreq5_p & v845542;
assign d3086e = hbusreq0 & d3086a | !hbusreq0 & d3086d;
assign d3084b = hbusreq1_p & d307ad | !hbusreq1_p & !v845542;
assign v138a3c1 = decide_p & v138a3c0 | !decide_p & !v845542;
assign a646d9 = jx2_p & a656b9 | !jx2_p & a646d8;
assign v1214c89 = hmaster2_p & v121535e | !hmaster2_p & v845542;
assign v12acff9 = hlock0_p & v12ad5a3 | !hlock0_p & !v12acff8;
assign v1215066 = hmaster0_p & v1215030 | !hmaster0_p & v1215065;
assign v1389e2b = hgrant5_p & v1389e2a | !hgrant5_p & !v845542;
assign v1552d78 = hgrant3_p & v1552d75 | !hgrant3_p & v1552d77;
assign v12ad5e0 = hbusreq0 & v12ad5df | !hbusreq0 & v12afe63;
assign v144647e = hgrant4_p & v144647d | !hgrant4_p & v845542;
assign v1216acf = hlock1_p & v1216ace | !hlock1_p & !v845542;
assign v12ad22e = decide_p & v12ad22d | !decide_p & v12afe76;
assign v12ad4e8 = hbusreq0 & v12ad4e7 | !hbusreq0 & v845542;
assign v10d428f = hmastlock_p & v10d428e | !hmastlock_p & v845542;
assign v14459b9 = hbusreq1_p & v144639c | !hbusreq1_p & v14459b8;
assign d30165 = hgrant3_p & d2ff0d | !hgrant3_p & d30164;
assign d306f0 = hburst1 & d306ee | !hburst1 & d306ef;
assign d307ba = hbusreq5_p & d307ab | !hbusreq5_p & d307b9;
assign v10d4075 = hbusreq0_p & v10d3fd9 | !hbusreq0_p & !v10d3fdf;
assign v144582b = hbusreq2_p & v144581f | !hbusreq2_p & v144582a;
assign f2f4bf = hmaster1_p & v845542 | !hmaster1_p & f2f4be;
assign v1284cd5 = hlock4_p & v1284c8f | !hlock4_p & !v1405854;
assign v1214eb2 = hbusreq2 & v1214e82 | !hbusreq2 & v845542;
assign v1214e7c = hlock2_p & v1214e74 | !hlock2_p & !v1214e7b;
assign v1215726 = hgrant0_p & v845542 | !hgrant0_p & !v1215710;
assign v1445823 = hbusreq2_p & v144581f | !hbusreq2_p & v1445822;
assign v1446196 = hbusreq2_p & v1446186 | !hbusreq2_p & v1446195;
assign v16a1be5 = hgrant5_p & v845542 | !hgrant5_p & !v16a1bd7;
assign v16a1f95 = hmaster2_p & v845542 | !hmaster2_p & !v84554d;
assign v12af98e = hmaster1_p & v12af7f7 | !hmaster1_p & v12af98d;
assign v144578d = hmaster1_p & v144578c | !hmaster1_p & v1445e07;
assign v14462e7 = hmaster2_p & v14465ae | !hmaster2_p & v144639c;
assign v1284d61 = hgrant2_p & v1284d5c | !hgrant2_p & v1284d60;
assign v1214d7f = hbusreq2_p & v1214d7d | !hbusreq2_p & v1214d7e;
assign v1216afd = hmaster1_p & v1216afc | !hmaster1_p & v1216af8;
assign v12160bc = hlock2_p & v12160ba | !hlock2_p & v12160bb;
assign v134ce9b = hbusreq0 & v134ce9a | !hbusreq0 & v134d23b;
assign d307f5 = hmaster1_p & d307a6 | !hmaster1_p & d307f4;
assign v121651d = hlock5_p & v845547 | !hlock5_p & !v845542;
assign d3061a = hlock5_p & v845542 | !hlock5_p & !d30619;
assign v144614b = hbusreq2_p & v1446149 | !hbusreq2_p & v144614a;
assign d3023f = hgrant5_p & v845542 | !hgrant5_p & d301d8;
assign f2f4ab = hmaster0_p & f2f4aa | !hmaster0_p & v845542;
assign d80746 = hmaster0_p & d80741 | !hmaster0_p & d80745;
assign v1445f0d = hgrant2_p & v1445ef3 | !hgrant2_p & v1445f0c;
assign v1446148 = hbusreq2 & v1446146 | !hbusreq2 & v1446147;
assign v138a44b = hmaster1_p & v138a44a | !hmaster1_p & v138a341;
assign v1553056 = hlock0_p & v1553399 | !hlock0_p & v1553055;
assign v12ad00a = hgrant1_p & v12ad5bd | !hgrant1_p & v12ad009;
assign v1445bcb = hmaster0_p & v144643b | !hmaster0_p & v144639c;
assign v121600e = hmaster2_p & v1215fea | !hmaster2_p & v1215ffa;
assign v1216a67 = hready & v1216a66 | !hready & a66294;
assign f2f427 = hbusreq0 & f2f421 | !hbusreq0 & f2f426;
assign v12150e3 = hbusreq2 & v12150dd | !hbusreq2 & v12150e2;
assign v1552f89 = hlock5 & v155341e | !hlock5 & v1552f78;
assign v144552a = hlock5 & v1445512 | !hlock5 & v1445529;
assign v16a1afb = hmaster2_p & v16a1afa | !hmaster2_p & v845542;
assign d3067e = hgrant2_p & v845542 | !hgrant2_p & d3067d;
assign v1215fb9 = hgrant2_p & v1215fb7 | !hgrant2_p & v1215fb8;
assign v12af73d = hready_p & v12afe77 | !hready_p & v12af73c;
assign v1214c47 = hlock0_p & v1216523 | !hlock0_p & v845542;
assign v11e5950 = hlock5_p & v11e594e | !hlock5_p & v11e594f;
assign v10d4277 = hmaster1_p & v10d4276 | !hmaster1_p & !v10d404f;
assign v1216b15 = hbusreq2_p & v1216b14 | !hbusreq2_p & v1216b10;
assign a6543d = hgrant5_p & a6587e | !hgrant5_p & a653f5;
assign v1446333 = hmaster0_p & v14462e6 | !hmaster0_p & v1446332;
assign v12163a4 = hbusreq4 & v1216ac7 | !hbusreq4 & !v1216acd;
assign v138953a = hbusreq5_p & v1389539 | !hbusreq5_p & !v845542;
assign v1215c22 = hbusreq5_p & v1215c1e | !hbusreq5_p & v1215c21;
assign v16a2074 = hgrant0_p & v845542 | !hgrant0_p & !v16a2073;
assign d30703 = hlock0_p & v845542 | !hlock0_p & d30702;
assign f2f33f = hbusreq3 & f2f337 | !hbusreq3 & f2f33e;
assign v14058b5 = hmaster0_p & v1405856 | !hmaster0_p & v14058b4;
assign v1216711 = hbusreq2_p & v1216710 | !hbusreq2_p & v121670d;
assign v134d1ee = hgrant4_p & v134d1ed | !hgrant4_p & v134d1e8;
assign v1553142 = hbusreq1_p & v1553141 | !hbusreq1_p & v845542;
assign a65395 = hbusreq4_p & a65394 | !hbusreq4_p & !v845542;
assign v12ad510 = stateA1_p & v12ad50f | !stateA1_p & a658a5;
assign v1445528 = hlock3 & v14454fa | !hlock3 & v1445524;
assign v1215339 = hmaster1_p & v1215338 | !hmaster1_p & !v12150a6;
assign d30619 = hmaster2_p & v16693aa | !hmaster2_p & d305f2;
assign v1215cbc = hgrant1_p & v1215cbb | !hgrant1_p & v1216152;
assign f2f455 = hmaster1_p & f2f449 | !hmaster1_p & f2f454;
assign d2f96c = hbusreq1_p & d2fe9a | !hbusreq1_p & d2f96b;
assign v14466d3 = hbusreq2_p & v14466d1 | !hbusreq2_p & v14466d2;
assign v1405878 = hmaster1_p & v1405871 | !hmaster1_p & v140586f;
assign v138a43d = hbusreq5_p & v138a313 | !hbusreq5_p & v845542;
assign v1405b1a = hbusreq1_p & v845542 | !hbusreq1_p & v1405b19;
assign v1445e94 = hmaster2_p & v1446609 | !hmaster2_p & v1445e93;
assign v121540d = hlock5_p & v121540c | !hlock5_p & v12153de;
assign v1215d68 = hmaster0_p & v1215d67 | !hmaster0_p & v12164df;
assign d307d6 = hgrant0_p & d307d5 | !hgrant0_p & v845542;
assign v138a334 = hbusreq4_p & v1668cc4 | !hbusreq4_p & v1668cdd;
assign v134d285 = hmaster2_p & v845542 | !hmaster2_p & v134d284;
assign v14465c3 = hlock4 & v144639c | !hlock4 & v14465bb;
assign v1553435 = hbusreq5 & v1553434 | !hbusreq5 & v155321a;
assign v1668d16 = hmaster2_p & a65851 | !hmaster2_p & a6585c;
assign v12166c2 = hmaster1_p & v12166c1 | !hmaster1_p & v12164e1;
assign v12162f6 = hmaster2_p & v1216048 | !hmaster2_p & v845547;
assign v1215462 = hmaster2_p & v121545f | !hmaster2_p & v1215461;
assign d2fafe = hbusreq0 & d2faf9 | !hbusreq0 & d2fafd;
assign d300e0 = hmaster2_p & d300c4 | !hmaster2_p & d300df;
assign v1215d2f = hgrant5_p & v1668da6 | !hgrant5_p & v1215d2e;
assign v1668c48 = decide_p & v1668c47 | !decide_p & v845542;
assign v1215381 = hmaster2_p & v121537c | !hmaster2_p & v1215380;
assign v1215cd0 = hmaster2_p & v1215c8c | !hmaster2_p & v1215cb4;
assign d8073e = hmaster2_p & d80732 | !hmaster2_p & d8073d;
assign v1216172 = hmaster2_p & v121601c | !hmaster2_p & !v121611d;
assign v1214d13 = hmaster2_p & v1214c29 | !hmaster2_p & !v1214d12;
assign v1445ef6 = hbusreq2_p & v1445ef2 | !hbusreq2_p & v1445ef5;
assign v12aeb1c = hmaster2_p & v845542 | !hmaster2_p & v12afda7;
assign a66281 = hready_p & v845542 | !hready_p & a66280;
assign v1515632 = hmaster0_p & v1515631 | !hmaster0_p & v1668da6;
assign v14465f0 = hgrant4_p & v14465ed | !hgrant4_p & v14465ef;
assign v15532ca = hgrant5_p & v845542 | !hgrant5_p & v15532c9;
assign v1515652 = hburst1 & d305ee | !hburst1 & v1515651;
assign v14464a5 = hmaster2_p & v845542 | !hmaster2_p & v1446476;
assign v121627c = hmaster1_p & v121627b | !hmaster1_p & v12160e0;
assign d302dd = hready_p & d302d4 | !hready_p & !d302dc;
assign v1215beb = hmaster0_p & v1215be9 | !hmaster0_p & v1215bea;
assign d2f9b5 = hbusreq2_p & d2f998 | !hbusreq2_p & d2f9aa;
assign v10d42e1 = jx2_p & v10d40de | !jx2_p & v10d42e0;
assign v138a31c = hmaster1_p & v138a31b | !hmaster1_p & v845542;
assign v12153bd = hbusreq4_p & v12153bc | !hbusreq4_p & v845542;
assign v121579d = hgrant5_p & v845542 | !hgrant5_p & v121576b;
assign v1446284 = hbusreq2_p & v144627f | !hbusreq2_p & v1446283;
assign v16a1cd9 = hbusreq2_p & v16a1b03 | !hbusreq2_p & v16a1cd8;
assign v1445ae9 = hbusreq2_p & v1445ae6 | !hbusreq2_p & v1445ae8;
assign v144599e = hmaster2_p & v144599d | !hmaster2_p & v14465b3;
assign v1284d41 = hready_p & v1284d31 | !hready_p & !v1284d40;
assign d80762 = hmaster2_p & d80760 | !hmaster2_p & !v845542;
assign v1668e0e = hbusreq3_p & v1668e0d | !hbusreq3_p & !v1668c39;
assign v12161fd = hmaster1_p & v12161fc | !hmaster1_p & v12161f4;
assign v14466a9 = hmaster0_p & v1446695 | !hmaster0_p & v14466a8;
assign v14465ef = hbusreq4_p & v14465b1 | !hbusreq4_p & v14465ee;
assign v12160f1 = hbusreq1 & v12160f0 | !hbusreq1 & v845542;
assign v1284d05 = hbusreq2_p & v1284cff | !hbusreq2_p & v1284d04;
assign a653e4 = hgrant5_p & a653d4 | !hgrant5_p & a653e2;
assign v12165a2 = hmaster2_p & v121659c | !hmaster2_p & v12165a1;
assign v1445e12 = hbusreq0 & v1445e11 | !hbusreq0 & v1445e0a;
assign v1445b18 = hbusreq2_p & v1445b16 | !hbusreq2_p & v1445b17;
assign v134ce91 = hmaster1_p & v134ce90 | !hmaster1_p & v134d23c;
assign v140585f = stateA1_p & v85e70d | !stateA1_p & !v146b550;
assign d30802 = hlock5_p & d30800 | !hlock5_p & !d30801;
assign v1668d5d = hgrant1_p & v1668d53 | !hgrant1_p & v1668d58;
assign v1214d19 = hbusreq2 & v1214d11 | !hbusreq2 & v1214d18;
assign v12162d8 = hmaster1_p & v12162d7 | !hmaster1_p & !v121624b;
assign v15168b8 = hready_p & v845542 | !hready_p & v15168b7;
assign v144536b = hmaster1_p & v144536a | !hmaster1_p & v14458fd;
assign v1216208 = hmaster2_p & v1216207 | !hmaster2_p & v12161d0;
assign f2e4fc = hmaster1_p & f2e4fb | !hmaster1_p & f2f52c;
assign v14459c8 = hgrant4_p & v14458df | !hgrant4_p & v14459c7;
assign v1445db7 = hbusreq0 & v1445db6 | !hbusreq0 & v1445da7;
assign v1214d39 = hbusreq2_p & v1215372 | !hbusreq2_p & v1216a81;
assign v12163a5 = hlock4_p & v12163a4 | !hlock4_p & !v845542;
assign v121570d = hbusreq1 & v12160ec | !hbusreq1 & !v845542;
assign v134d38e = hbusreq0_p & v134d273 | !hbusreq0_p & v134d370;
assign f2e732 = hmaster0_p & f2e715 | !hmaster0_p & f2e731;
assign v14457c8 = hlock2 & v14457c5 | !hlock2 & v14457c7;
assign v10d4270 = hmaster1_p & v10d426f | !hmaster1_p & !v10d404f;
assign v1515653 = hburst0 & d305ee | !hburst0 & v1515652;
assign v1216291 = hmaster0_p & v12161a1 | !hmaster0_p & v121618e;
assign v1215033 = hbusreq4_p & v1215032 | !hbusreq4_p & !v845542;
assign d80737 = hlock3_p & d80736 | !hlock3_p & v845542;
assign d2fb53 = hmaster2_p & d2fb4d | !hmaster2_p & v845542;
assign f2f3a1 = hmaster2_p & f2f350 | !hmaster2_p & !f2f39a;
assign d2fc14 = hgrant2_p & v84554a | !hgrant2_p & d2fc12;
assign v12153e3 = hlock4_p & v12153e1 | !hlock4_p & v12153e2;
assign v14465ac = stateA1_p & v146d169 | !stateA1_p & v845542;
assign v121614e = hbusreq0_p & v1216523 | !hbusreq0_p & v12160f2;
assign v1445a6e = hgrant2_p & v1445a6d | !hgrant2_p & v1445a5c;
assign d2fd0b = hbusreq2_p & d2fd0a | !hbusreq2_p & d302d6;
assign v121627d = hbusreq2_p & v121627a | !hbusreq2_p & v121627c;
assign v12afe62 = hgrant1_p & v845542 | !hgrant1_p & v12afe61;
assign v134cd73 = hmaster1_p & v134cd72 | !hmaster1_p & v845542;
assign v1445881 = hbusreq0_p & v14463d8 | !hbusreq0_p & v144639e;
assign v1284d0f = hmaster2_p & v1284c8f | !hmaster2_p & v1446412;
assign v121536a = hbusreq4_p & v1215364 | !hbusreq4_p & v845547;
assign v1214c8f = hbusreq0 & v1214c8e | !hbusreq0 & v845542;
assign d305dd = hmastlock_p & v1552d7a | !hmastlock_p & !v845542;
assign v1284d4d = hmaster2_p & v1284d4c | !hmaster2_p & v1405844;
assign v12160c0 = hlock2_p & v12160be | !hlock2_p & v12160bf;
assign v138944e = hmaster0_p & v138944d | !hmaster0_p & v845542;
assign d2fba6 = hmaster1_p & d2fb8d | !hmaster1_p & d2fb9d;
assign v16a1d12 = hbusreq5 & v16a1d10 | !hbusreq5 & v16a1d11;
assign v138a305 = hmaster0_p & v138a2f8 | !hmaster0_p & v138a304;
assign v1515c83 = hmaster1_p & v1515c82 | !hmaster1_p & v845542;
assign v14460d3 = hgrant2_p & v14460b9 | !hgrant2_p & v14460d2;
assign v1668d1a = hmaster2_p & a65862 | !hmaster2_p & v1668d18;
assign d80781 = hmaster2_p & d8077c | !hmaster2_p & d80780;
assign v1214e7b = hmaster1_p & v1214e1a | !hmaster1_p & v1215bc2;
assign v1668c56 = hready_p & v845542 | !hready_p & v1668c55;
assign v144641a = hlock4 & v1446408 | !hlock4 & v1446406;
assign v1215bf1 = hgrant1_p & v1215bf0 | !hgrant1_p & v12160f0;
assign v12162ef = hmaster2_p & v845547 | !hmaster2_p & v12162ed;
assign v1668d6f = hbusreq4 & a65394 | !hbusreq4 & a65396;
assign v1445b4e = hmaster0_p & v1445900 | !hmaster0_p & v1445a36;
assign v16695a4 = decide_p & v16695a3 | !decide_p & !v845542;
assign v1446152 = hmaster1_p & v1446134 | !hmaster1_p & v1445ffc;
assign v138a3e2 = hgrant2_p & v138a3c4 | !hgrant2_p & !v138a3e1;
assign v1445425 = hbusreq2 & v144541c | !hbusreq2 & v1445424;
assign a65401 = hbusreq0 & a653fc | !hbusreq0 & a65400;
assign v166959e = hmaster0_p & v1668c28 | !hmaster0_p & v845542;
assign v16a16b5 = hbusreq3_p & v16a1e59 | !hbusreq3_p & v16a16b4;
assign d80732 = hmastlock_p & d80731 | !hmastlock_p & !v845542;
assign v1214c2a = hbusreq0_p & v12164d3 | !hbusreq0_p & v845542;
assign v16a1c9f = hgrant5_p & v845542 | !hgrant5_p & v16a1c9e;
assign v1445490 = hbusreq2_p & v144548f | !hbusreq2_p & v1445bba;
assign v1405867 = hmaster2_p & v1405844 | !hmaster2_p & v1405863;
assign v134d3de = hgrant1_p & v845542 | !hgrant1_p & v134d3dd;
assign v1216114 = hgrant5_p & v121601e | !hgrant5_p & !v1216112;
assign v14454e9 = hmaster1_p & v14454e8 | !hmaster1_p & v144626a;
assign v134d23a = hlock5_p & v134d1ff | !hlock5_p & v134d1fd;
assign a6548b = hmaster2_p & a658b0 | !hmaster2_p & !a6546a;
assign v138a075 = decide_p & v138a074 | !decide_p & v845542;
assign v1405884 = hmaster1_p & v1405883 | !hmaster1_p & v140584d;
assign v144576e = hbusreq2 & v144576c | !hbusreq2 & v144576d;
assign v1445e8d = hgrant4_p & v1445dfc | !hgrant4_p & v1445e8c;
assign v14457af = hmaster1_p & v144577b | !hmaster1_p & v1445e28;
assign d2fb01 = hbusreq4_p & d300fb | !hbusreq4_p & d306a3;
assign v16a1da1 = hgrant3_p & v16a1d37 | !hgrant3_p & v16a1da0;
assign v1668db7 = hgrant5_p & v845542 | !hgrant5_p & !v1668d30;
assign v14463ab = hbusreq4_p & v144639c | !hbusreq4_p & v14463a0;
assign bf1fa3 = hbusreq5_p & bf1f6d | !hbusreq5_p & !bf1fa2;
assign v14453eb = hlock2 & v14453e4 | !hlock2 & v14453ea;
assign v14462ed = stateG10_5_p & v14465d3 | !stateG10_5_p & v14462ec;
assign d2fbac = hbusreq2_p & d2fbab | !hbusreq2_p & d2fba7;
assign v12ad4c5 = hbusreq2_p & v12adf65 | !hbusreq2_p & v12ad4c4;
assign v84554e = hlock1_p & v845542 | !hlock1_p & !v845542;
assign v1216047 = hmastlock_p & v144646d | !hmastlock_p & v845542;
assign v1215b82 = hmaster2_p & v1215b7d | !hmaster2_p & v1215b81;
assign v15157de = hgrant5_p & v1668da6 | !hgrant5_p & v1515733;
assign bf1f50 = hlock3_p & v845570 | !hlock3_p & !bf1f4f;
assign d2fb20 = hgrant5_p & d3068e | !hgrant5_p & d2faf7;
assign v1284ca3 = hlock4_p & v1284c8e | !hlock4_p & !v14463b1;
assign v1668d77 = hlock0_p & v1668d24 | !hlock0_p & v1668d76;
assign d300f8 = hbusreq1 & d2fea1 | !hbusreq1 & v84555a;
assign v144662a = hgrant1_p & v1446432 | !hgrant1_p & v1446629;
assign d80774 = hmaster2_p & v845542 | !hmaster2_p & !d80773;
assign v1214f06 = hgrant5_p & v16a2243 | !hgrant5_p & v1214eda;
assign v138a351 = hmaster1_p & v138a350 | !hmaster1_p & v138a341;
assign v16a2234 = hmaster2_p & v845547 | !hmaster2_p & !v845542;
assign v134ce76 = hlock3 & v134d276 | !hlock3 & v134ce75;
assign v1215d32 = hmaster2_p & v1216a8d | !hmaster2_p & v1216a93;
assign v1215744 = hbusreq1 & v1215b80 | !hbusreq1 & v845542;
assign v1214d67 = hbusreq0 & v1214d50 | !hbusreq0 & v845542;
assign f2f3a8 = hbusreq0 & f2f3a3 | !hbusreq0 & f2f3a7;
assign d2faf7 = hmaster2_p & d2fae2 | !hmaster2_p & d2faf6;
assign v138a311 = hmaster2_p & v845542 | !hmaster2_p & v10d3ff3;
assign v14458d4 = hmaster2_p & v14458d2 | !hmaster2_p & v1446403;
assign v14462ea = hgrant5_p & v1446688 | !hgrant5_p & v14465d3;
assign v140583b = stateA1_p & v845542 | !stateA1_p & v140583a;
assign v16a1a78 = hgrant1_p & v84554d | !hgrant1_p & v16a1a77;
assign v12ad4c6 = decide_p & v12ad4c5 | !decide_p & v12afe76;
assign v134d213 = hbusreq2_p & v134d212 | !hbusreq2_p & v134d211;
assign v1214f62 = hbusreq3 & v1214f5d | !hbusreq3 & v1214f61;
assign f2f3cc = hgrant5_p & v84554c | !hgrant5_p & f2f38e;
assign v1215d38 = hbusreq5_p & v1215d34 | !hbusreq5_p & !v1215d37;
assign v16a205c = hmaster1_p & v845542 | !hmaster1_p & !v16a2672;
assign v144542b = hmaster1_p & v14465aa | !hmaster1_p & v1446290;
assign v12ad577 = hmaster0_p & v12ad531 | !hmaster0_p & v12ad52d;
assign v14463c0 = hbusreq0 & v14463bd | !hbusreq0 & v14463bf;
assign v15155f1 = hbusreq0 & v1668c17 | !hbusreq0 & v845570;
assign v16a16ae = hbusreq2_p & v16a1e0c | !hbusreq2_p & v16a16ad;
assign v16a19df = hbusreq5_p & v16a1842 | !hbusreq5_p & v16a19de;
assign d30225 = hlock5_p & d30222 | !hlock5_p & !d30224;
assign v12150f4 = hmaster1_p & v12150df | !hmaster1_p & v12150ef;
assign v1405870 = hmaster1_p & v1405861 | !hmaster1_p & v140586f;
assign v1446137 = hmaster1_p & v1446136 | !hmaster1_p & v1445fde;
assign v1445f97 = hbusreq1_p & v144639c | !hbusreq1_p & v14463b9;
assign v144609e = hmaster0_p & v144603f | !hmaster0_p & v144607f;
assign v1445e78 = hbusreq5_p & v1445e6e | !hbusreq5_p & v1445e77;
assign v1445adc = hlock2 & v1445ad9 | !hlock2 & v1445adb;
assign d3028e = hbusreq3 & d3028d | !hbusreq3 & v845542;
assign v10d4091 = hmaster2_p & v10d3fd4 | !hmaster2_p & !v10d406d;
assign v138a451 = hmaster1_p & v138a450 | !hmaster1_p & v138a341;
assign v1214d75 = hmaster1_p & v1214d74 | !hmaster1_p & v1215357;
assign v1214ff0 = hbusreq4_p & v1214fef | !hbusreq4_p & !v845542;
assign v1216028 = hmaster1_p & v121601e | !hmaster1_p & !v1216027;
assign d3010b = hlock5_p & d30109 | !hlock5_p & d3010a;
assign v12af9d5 = hbusreq5_p & v12afe5f | !hbusreq5_p & v12af9d4;
assign v1216002 = hbusreq1_p & v1216001 | !hbusreq1_p & v845542;
assign v1445f90 = hbusreq0 & v1445f8c | !hbusreq0 & v1445f8f;
assign v134d3d2 = hlock2 & v134d276 | !hlock2 & v134d3d1;
assign v10d4269 = hgrant0_p & v10d401b | !hgrant0_p & !v10d4268;
assign v16a1f9e = hbusreq5 & v16a1f94 | !hbusreq5 & !v16a1f9d;
assign v121535c = hbusreq2_p & v1215358 | !hbusreq2_p & v121535b;
assign d2fc54 = hgrant4_p & d2fbce | !hgrant4_p & d2fc53;
assign v1668d8f = hmaster0_p & v1668d2b | !hmaster0_p & v1668d8e;
assign d2fb72 = hmaster2_p & v84554a | !hmaster2_p & d2fb70;
assign v1214d18 = hbusreq2_p & v1214d17 | !hbusreq2_p & v1214d10;
assign v1445882 = hlock0_p & v14463d8 | !hlock0_p & v1445881;
assign v1445df6 = hmaster2_p & v1446403 | !hmaster2_p & v1445df5;
assign d807ba = hmaster1_p & d807b9 | !hmaster1_p & !v845542;
assign v1445e3e = hgrant5_p & v1445e3d | !hgrant5_p & v1445e3b;
assign v1215050 = hgrant1_p & v121546d | !hgrant1_p & v121504f;
assign d2fc76 = hmaster1_p & d2fc5a | !hmaster1_p & d2fc75;
assign d307b7 = hgrant1_p & v845542 | !hgrant1_p & d307b6;
assign v1553511 = hbusreq2 & v155350f | !hbusreq2 & v1553510;
assign v16a1445 = hbusreq2 & v16a1443 | !hbusreq2 & !v16a1444;
assign d2fb2f = hgrant2_p & d2f984 | !hgrant2_p & d2fb2b;
assign f2f3dc = hbusreq2_p & f2f3d1 | !hbusreq2_p & f2f3db;
assign v1445f7d = hlock3 & v144673f | !hlock3 & v1445f7b;
assign v1214cff = hgrant4_p & v1214cfe | !hgrant4_p & v845572;
assign v134d3e7 = hready_p & v134d3e5 | !hready_p & v134d3e6;
assign v14457d5 = hready_p & v1445f26 | !hready_p & v14457d4;
assign v121503d = hmaster2_p & v1215033 | !hmaster2_p & !v1215467;
assign f2e3fd = decide_p & f2e3fc | !decide_p & f2f23c;
assign d30250 = hmaster0_p & d3024c | !hmaster0_p & d3024f;
assign v10d401b = hlock0_p & v10d3fd5 | !hlock0_p & !v10d3fd4;
assign v1445f3a = hmaster1_p & v1445f39 | !hmaster1_p & v1445dc2;
assign a65920 = hbusreq2 & a6591b | !hbusreq2 & a6591f;
assign v14465b9 = hbusreq1_p & v1446403 | !hbusreq1_p & v1446444;
assign v134d392 = hlock1 & v134d385 | !hlock1 & v134d391;
assign v11f3405 = jx0_p & v11f33c6 | !jx0_p & v8b6f6c;
assign v1445e7c = hgrant1_p & v1445e7a | !hgrant1_p & v1445e7b;
assign v1445e0a = hmaster2_p & v1445de5 | !hmaster2_p & v1445dec;
assign v1445847 = hbusreq2_p & v1445844 | !hbusreq2_p & v1445846;
assign v16a1e2c = hmaster0_p & v16a1e27 | !hmaster0_p & v16a1e23;
assign v1216020 = hbusreq5_p & v121601d | !hbusreq5_p & v121601f;
assign v1215d75 = hbusreq5_p & v1215d71 | !hbusreq5_p & !v1215d74;
assign v134d382 = hbusreq1 & v134d37f | !hbusreq1 & v134d381;
assign v138a39a = hmaster0_p & v138a394 | !hmaster0_p & v138a34f;
assign d3022a = hlock5_p & d30228 | !hlock5_p & !d30229;
assign v1215793 = hlock5_p & v1215790 | !hlock5_p & v1215792;
assign d301d6 = hbusreq5_p & d301d5 | !hbusreq5_p & !d301d4;
assign v1668d2f = hgrant1_p & v1668d23 | !hgrant1_p & v1668d2e;
assign v134d275 = hmaster0_p & v134d274 | !hmaster0_p & v845542;
assign v12166e4 = locked_p & v12166e3 | !locked_p & v845542;
assign a656cb = hbusreq5_p & a656be | !hbusreq5_p & a656ca;
assign v1214d5c = hmaster2_p & v1214d4e | !hmaster2_p & v1214d42;
assign v16a1d65 = hgrant2_p & v845542 | !hgrant2_p & v16a1d63;
assign v10d42aa = decide_p & v10d4279 | !decide_p & v10d42a9;
assign v1405b14 = hgrant1_p & v1405abb | !hgrant1_p & v1405b13;
assign v16a140b = hbusreq2_p & v16a140a | !hbusreq2_p & v16a2058;
assign v1216133 = hgrant5_p & v121611d | !hgrant5_p & v1216132;
assign v1216186 = hmaster1_p & v1216185 | !hmaster1_p & v845542;
assign d305fb = hlock0_p & d305ea | !hlock0_p & !v845542;
assign d807af = hmaster0_p & d80762 | !hmaster0_p & d807ae;
assign v1215c9e = hbusreq0 & v1215c98 | !hbusreq0 & v1215c9d;
assign v1446651 = hbusreq2_p & v1446632 | !hbusreq2_p & v144664d;
assign v1445bf9 = hbusreq3_p & v1445be9 | !hbusreq3_p & v1445bf8;
assign v1389fcc = hlock3_p & v1389fb4 | !hlock3_p & v1389fcb;
assign v16a12f3 = hbusreq0 & v16a12f2 | !hbusreq0 & v16a209b;
assign v134d20a = hmaster2_p & v134d1e8 | !hmaster2_p & v845542;
assign f2f3fe = hmaster0_p & f2f2e8 | !hmaster0_p & f2f2e3;
assign v14454a8 = hready_p & v1445442 | !hready_p & v14454a7;
assign d300d3 = hbusreq0 & d300c9 | !hbusreq0 & d300d2;
assign v14463bc = hmaster2_p & v14463b9 | !hmaster2_p & v14463bb;
assign f2f2e1 = hbusreq1 & a658bd | !hbusreq1 & !v845542;
assign v14457b0 = hbusreq2_p & v14457ae | !hbusreq2_p & v14457af;
assign v1445afc = hbusreq2_p & v1445af6 | !hbusreq2_p & v1445afb;
assign v134d309 = hbusreq2_p & v134d296 | !hbusreq2_p & v134d308;
assign v14460d1 = hgrant2_p & v14460ae | !hgrant2_p & v14460d0;
assign v1215c91 = hbusreq0 & v1215c8b | !hbusreq0 & v1215c90;
assign v1214eb6 = hmaster1_p & v1214eb5 | !hmaster1_p & v1214e0f;
assign v12ad537 = hmaster0_p & v12ad517 | !hmaster0_p & v12ad536;
assign v12ad4d5 = hbusreq1_p & v12ad4d0 | !hbusreq1_p & v12ad4d4;
assign v138a4a1 = hgrant3_p & v138a477 | !hgrant3_p & v138a4a0;
assign v1445ff5 = hbusreq2 & v1445fee | !hbusreq2 & v1445ff4;
assign v1405aeb = hgrant0_p & v1405aea | !hgrant0_p & !v1405a92;
assign v1446347 = hmaster1_p & v1446323 | !hmaster1_p & v1446341;
assign v1215b9d = hmaster2_p & v1215b99 | !hmaster2_p & v1215b9c;
assign v1445a8d = hlock2 & v1445a88 | !hlock2 & v1445a8c;
assign v12afda6 = hlock0_p & v15168ad | !hlock0_p & v845542;
assign d30835 = hlock5_p & d30833 | !hlock5_p & d30834;
assign v144551b = hbusreq2 & v1445515 | !hbusreq2 & v144551a;
assign v1446665 = hmaster1_p & v1446664 | !hmaster1_p & v1446630;
assign v16a1a7a = hgrant5_p & v845542 | !hgrant5_p & v16a1a79;
assign f2f3f4 = hmaster1_p & f2f3f3 | !hmaster1_p & f2f2db;
assign v138a463 = hbusreq2 & v138a45b | !hbusreq2 & v138a462;
assign v1215798 = hlock5_p & v1215796 | !hlock5_p & v1215797;
assign v134d202 = hbusreq0 & v134d1fe | !hbusreq0 & v134d201;
assign v15157f7 = hbusreq5_p & v15157f5 | !hbusreq5_p & !v15157f6;
assign v1668d64 = hbusreq1 & v1668d63 | !hbusreq1 & !v845542;
assign v15156f9 = hbusreq2 & v15156f8 | !hbusreq2 & v15167ed;
assign v1445b9d = hbusreq2_p & v1445b8f | !hbusreq2_p & v1445b9c;
assign v15161d7 = hbusreq3 & v15161d6 | !hbusreq3 & v1516804;
assign v1214d41 = hbusreq1 & v845547 | !hbusreq1 & v121536a;
assign d2fee6 = hmaster1_p & d2feb5 | !hmaster1_p & d2fee5;
assign d2fceb = hlock2_p & v845542 | !hlock2_p & !d2fcea;
assign v134d312 = hmaster2_p & v134d30e | !hmaster2_p & v134d311;
assign v10d40bb = hbusreq0_p & v10d3fd4 | !hbusreq0_p & v10d40ba;
assign v1445a0c = hlock0_p & v1445a0a | !hlock0_p & v1445a0b;
assign v1405b3c = hready_p & v1405b3a | !hready_p & v1405b3b;
assign a65384 = hbusreq4_p & a65382 | !hbusreq4_p & v845542;
assign v12166d9 = hgrant1_p & v12164dc | !hgrant1_p & v12166d8;
assign d308b9 = hbusreq5_p & d30835 | !hbusreq5_p & d308b8;
assign a6587e = hbusreq4_p & v845570 | !hbusreq4_p & v845542;
assign v1446117 = hbusreq5 & v1446115 | !hbusreq5 & v1446116;
assign v10d3fde = stateA1_p & v845542 | !stateA1_p & v88d3e4;
assign v14460bd = hmaster1_p & v144608b | !hmaster1_p & v1445ffc;
assign a654c0 = hbusreq2_p & a654bd | !hbusreq2_p & a654be;
assign d308e3 = hlock1_p & d308e2 | !hlock1_p & v845542;
assign v1445e53 = hmaster1_p & v14465aa | !hmaster1_p & v1445e07;
assign v12153df = hlock5_p & v12153dd | !hlock5_p & v12153de;
assign v1216afa = hmaster2_p & v1216aa9 | !hmaster2_p & v845547;
assign v1553418 = hmaster1_p & v1553417 | !hmaster1_p & v845542;
assign v1216323 = hmaster1_p & v12162f7 | !hmaster1_p & v1216322;
assign v1216a78 = hmaster2_p & v845542 | !hmaster2_p & v1216a77;
assign v134cedc = hlock5 & v134d3ce | !hlock5 & v134cedb;
assign v144633b = hgrant5_p & v14462eb | !hgrant5_p & v144633a;
assign v1445e38 = hbusreq4_p & v144646e | !hbusreq4_p & v1446476;
assign v1446433 = hmaster2_p & v144641f | !hmaster2_p & v1446432;
assign v1515725 = hgrant5_p & v151570f | !hgrant5_p & v1515724;
assign v11e5947 = hmaster2_p & v11e5946 | !hmaster2_p & v845542;
assign d30887 = hbusreq1_p & d30791 | !hbusreq1_p & d306a5;
assign v1668dca = hbusreq0 & v1668dc6 | !hbusreq0 & v1668dc9;
assign d30242 = hmaster2_p & d3070c | !hmaster2_p & !v845542;
assign a65490 = hmaster1_p & a6548f | !hmaster1_p & a65476;
assign v15532cd = hgrant2_p & v155321e | !hgrant2_p & v15532cc;
assign d30648 = hgrant1_p & f2f227 | !hgrant1_p & d30647;
assign d305f5 = hbusreq1_p & d305f4 | !hbusreq1_p & !v845542;
assign v12aeb82 = hbusreq3 & v12aeb7c | !hbusreq3 & v12afe3d;
assign v15168f1 = hburst1 & a66293 | !hburst1 & v15168f0;
assign f2f42e = hbusreq0 & f2f42a | !hbusreq0 & f2f42d;
assign a656a9 = hmaster1_p & a65495 | !hmaster1_p & !a65916;
assign d30113 = hmaster1_p & d30112 | !hmaster1_p & !d2fea2;
assign v12160b0 = hmaster1_p & v12160af | !hmaster1_p & v121605d;
assign v1668d44 = hbusreq1 & a6585c | !hbusreq1 & a6588d;
assign v138a455 = hbusreq2_p & v138a452 | !hbusreq2_p & v138a454;
assign v1668cd8 = hmaster2_p & a658ad | !hmaster2_p & !v845542;
assign v11e5965 = hgrant1_p & v845542 | !hgrant1_p & !v11e5964;
assign v14838b7 = hgrant4_p & v845542 | !hgrant4_p & v845558;
assign v14459f7 = hgrant0_p & v14459f6 | !hgrant0_p & v14459c0;
assign d2fb85 = hbusreq0 & d2fb84 | !hbusreq0 & v845542;
assign v16a1bce = hbusreq0 & v16a1bc0 | !hbusreq0 & v16a1bcd;
assign v12af9c2 = hgrant5_p & d30690 | !hgrant5_p & v12af9c1;
assign a65929 = hbusreq5 & a65911 | !hbusreq5 & a65928;
assign v12ad5b9 = hlock1_p & v12ad5b7 | !hlock1_p & v12ad5b8;
assign v12160c3 = hmaster1_p & v12160ad | !hmaster1_p & v1216082;
assign a65af9 = jx2_p & a662be | !jx2_p & a65af8;
assign v1552d58 = hlock2 & v155341e | !hlock2 & v1552d4e;
assign v121579a = hbusreq5_p & v1215798 | !hbusreq5_p & v1215799;
assign v14058c5 = locked_p & v140583e | !locked_p & v1405844;
assign v134d4c2 = decide_p & v134d3ce | !decide_p & v134d276;
assign v1552d51 = hbusreq0 & v1553413 | !hbusreq0 & v1553218;
assign v16a207c = hgrant0_p & v845542 | !hgrant0_p & !v16a206a;
assign v16a1e8f = hgrant1_p & v84554d | !hgrant1_p & v16a1e8e;
assign v12147ef = hgrant2_p & v845542 | !hgrant2_p & v12147ee;
assign v12af5a6 = hgrant4_p & v845542 | !hgrant4_p & v12af5a5;
assign v138a327 = hburst1 & v138a324 | !hburst1 & v138a326;
assign v12ad52e = hmaster0_p & v12ad517 | !hmaster0_p & v12ad52d;
assign v1445f04 = hmaster2_p & v1445edc | !hmaster2_p & v1445def;
assign v16695a1 = hmaster1_p & v16695a0 | !hmaster1_p & v845542;
assign v14458f8 = hbusreq1 & v14458f5 | !hbusreq1 & v14458f7;
assign v12ad8e5 = hmaster2_p & d30690 | !hmaster2_p & !v12ad8e4;
assign v1552d89 = hgrant0_p & v1552d88 | !hgrant0_p & v845542;
assign v1215c45 = hbusreq0 & v1215c40 | !hbusreq0 & v1215c44;
assign v15157f2 = hgrant5_p & v845570 | !hgrant5_p & v1515775;
assign v1552d8f = hmaster1_p & v1553224 | !hmaster1_p & v1552d8e;
assign v15167eb = hbusreq2_p & v15167ea | !hbusreq2_p & v845542;
assign v15534fa = hgrant5_p & v15534f9 | !hgrant5_p & v1553394;
assign v1405b43 = hmaster1_p & v1405b42 | !hmaster1_p & v1405af0;
assign a654b1 = hmaster1_p & a65465 | !hmaster1_p & !a654b0;
assign v845584 = stateG3_0_p & v845542 | !stateG3_0_p & !v845542;
assign d30211 = hgrant1_p & d30209 | !hgrant1_p & d307e9;
assign f2f328 = hmaster0_p & f2f2e3 | !hmaster0_p & f2f2e8;
assign d30768 = hmaster1_p & d30767 | !hmaster1_p & d3072c;
assign v1216587 = hgrant4_p & v845570 | !hgrant4_p & v1216586;
assign v12afa0f = hbusreq2_p & v12afe72 | !hbusreq2_p & v12afa0e;
assign d302ed = decide_p & d302ec | !decide_p & v845570;
assign v12ad007 = hbusreq5_p & v12ad5e9 | !hbusreq5_p & v12ad006;
assign v12ad5bb = hlock0_p & a65396 | !hlock0_p & v845542;
assign v14453e5 = hbusreq2_p & v1446237 | !hbusreq2_p & v14453e2;
assign v1405ae8 = hgrant1_p & v1405a90 | !hgrant1_p & !v1405ae7;
assign v121631c = hmaster1_p & v12162ea | !hmaster1_p & v121631b;
assign v10d42dd = decide_p & v10d40a8 | !decide_p & v10d42dc;
assign v1215cd9 = hmaster2_p & v845542 | !hmaster2_p & v1216014;
assign v1215bfa = hbusreq5_p & v1215bf8 | !hbusreq5_p & !v1215bf9;
assign d2fb9b = hbusreq5_p & d2fb9a | !hbusreq5_p & d2fb72;
assign v144605f = hmaster2_p & v144605a | !hmaster2_p & v144605e;
assign v12af21e = hgrant5_p & d30690 | !hgrant5_p & v12af21d;
assign v16a16a3 = hbusreq2_p & v16a1e08 | !hbusreq2_p & v16a16a2;
assign v14461f1 = hbusreq2_p & v14461ee | !hbusreq2_p & v14461f0;
assign v1214fed = hgrant5_p & v12153b5 | !hgrant5_p & v1214fec;
assign v14454fd = hmaster1_p & v14454f0 | !hmaster1_p & v1446341;
assign v1214e72 = hbusreq5_p & v1214e71 | !hbusreq5_p & v1214df5;
assign v14458c7 = hlock2 & v14458c4 | !hlock2 & v14458c6;
assign v144552f = hmaster1_p & v1445506 | !hmaster1_p & v1445b8d;
assign v1552f63 = hbusreq1 & v1552f61 | !hbusreq1 & v1552f62;
assign v12acffd = hbusreq1_p & v12ad5a7 | !hbusreq1_p & v12acffc;
assign d8078d = hmaster2_p & v845542 | !hmaster2_p & !d8078c;
assign v16a1cc9 = hgrant3_p & v16a1bb3 | !hgrant3_p & v16a1cc8;
assign v1216550 = hready & v1216a60 | !hready & a66294;
assign v1216adb = hmaster2_p & v1216ad6 | !hmaster2_p & v1216ada;
assign v12162a1 = hbusreq5 & v1216290 | !hbusreq5 & v12162a0;
assign v12ad5a7 = hgrant4_p & v12ad59e | !hgrant4_p & !v12ad5a6;
assign v1668dc4 = hmaster2_p & a65396 | !hmaster2_p & v845542;
assign v12162bb = hbusreq2_p & v12162b6 | !hbusreq2_p & v12162ba;
assign v10d4022 = hgrant0_p & v10d4021 | !hgrant0_p & !v10d3fd8;
assign v138a45d = hmaster1_p & v138a45c | !hmaster1_p & v138a341;
assign v1445fb6 = hbusreq3 & v1445fb4 | !hbusreq3 & v1445fb5;
assign v144577b = hmaster0_p & v1445778 | !hmaster0_p & v1445e0c;
assign v134cd59 = hbusreq1_p & v134d273 | !hbusreq1_p & v134cd58;
assign v121617d = hbusreq0 & v1216178 | !hbusreq0 & v121617c;
assign v14466f8 = hlock2 & v14466f4 | !hlock2 & v14466f7;
assign v15532c9 = hmaster2_p & v15532c5 | !hmaster2_p & v15532c8;
assign v1445556 = jx2_p & v144553d | !jx2_p & v1445555;
assign v16a1e79 = hbusreq3 & v16a1e73 | !hbusreq3 & v16a1e78;
assign f2f2a8 = hbusreq1_p & f2f233 | !hbusreq1_p & v845542;
assign a65622 = hbusreq1_p & a653a1 | !hbusreq1_p & a65621;
assign v1215399 = hlock0_p & v1216ab8 | !hlock0_p & !v1215398;
assign v1216036 = hbusreq1 & v16a1bc6 | !hbusreq1 & v845542;
assign f2f3ac = hbusreq2_p & f2f395 | !hbusreq2_p & f2f3ab;
assign f2f2db = hmaster0_p & f2f2d1 | !hmaster0_p & f2f2da;
assign d301c1 = hmaster0_p & d301bf | !hmaster0_p & d301c0;
assign v14460f6 = hmaster1_p & v14460f5 | !hmaster1_p & v1445f9e;
assign v15160fc = hbusreq2_p & v15160fb | !hbusreq2_p & v845542;
assign v1445da0 = hlock1 & v1445d99 | !hlock1 & v1445d9f;
assign v1214c7e = hgrant2_p & v121536e | !hgrant2_p & v1214c7d;
assign v1445b45 = hmaster0_p & v1445900 | !hmaster0_p & v14458d3;
assign f2f290 = hgrant3_p & f2f225 | !hgrant3_p & f2f28f;
assign v15156f0 = hbusreq5 & v15156ce | !hbusreq5 & v15156ef;
assign v1445b6e = hmaster1_p & v1446333 | !hmaster1_p & v1446290;
assign v144655e = hgrant4_p & v845542 | !hgrant4_p & v144655d;
assign v1216123 = hgrant4_p & v1216120 | !hgrant4_p & v1216122;
assign d3072b = hbusreq0 & d30726 | !hbusreq0 & d3072a;
assign v1446271 = hmaster0_p & v1446265 | !hmaster0_p & v144642c;
assign v1445e91 = hmaster2_p & v1446609 | !hmaster2_p & v1445e90;
assign d807aa = hmaster2_p & d807a9 | !hmaster2_p & !v845542;
assign d30217 = hbusreq0 & d3020f | !hbusreq0 & d30216;
assign v14466fd = hmaster1_p & v14466f9 | !hmaster1_p & v144644d;
assign v1215c08 = hbusreq1 & v1216a61 | !hbusreq1 & v1216568;
assign a6535e = hbusreq1 & a65852 | !hbusreq1 & a6587e;
assign d2fbfe = hmaster1_p & d2fbdb | !hmaster1_p & d2fbfd;
assign d2fea1 = hlock4_p & d30703 | !hlock4_p & !v845542;
assign v14459a2 = hgrant5_p & v14458d4 | !hgrant5_p & v14459a1;
assign v1552f7f = hmaster1_p & v1553385 | !hmaster1_p & v1552f7e;
assign v1216a7e = hbusreq5 & v1216a7d | !hbusreq5 & v845542;
assign v1445a5d = hgrant2_p & v1445a51 | !hgrant2_p & v1445a5c;
assign v15157fe = hgrant5_p & v15157fb | !hgrant5_p & v15157af;
assign v1215be9 = hbusreq5_p & v1215be7 | !hbusreq5_p & v1215be8;
assign v12153fd = hlock2_p & v12153fa | !hlock2_p & v12153fc;
assign v16a1ad2 = hbusreq2_p & v16a1f9a | !hbusreq2_p & v16a1ad1;
assign v14457e3 = hmaster1_p & v14457e2 | !hmaster1_p & v1445e07;
assign v1216a5f = hmastlock_p & v1216a5e | !hmastlock_p & v845542;
assign v16a1a7f = hbusreq2_p & v16a195d | !hbusreq2_p & v16a1a7e;
assign v151580f = hlock2_p & v151580e | !hlock2_p & !v845542;
assign d3029d = hlock3_p & d30264 | !hlock3_p & d3029c;
assign v12ad584 = hlock2_p & v12ad582 | !hlock2_p & v12ad583;
assign v121510f = hmaster1_p & v121510e | !hmaster1_p & v121546f;
assign v12166d2 = hgrant1_p & v12166cf | !hgrant1_p & v12166d1;
assign v134d30d = hgrant4_p & v134d1dd | !hgrant4_p & v845542;
assign v12150df = hmaster0_p & v12153ee | !hmaster0_p & v12150de;
assign v1445875 = hmaster2_p & v14463b1 | !hmaster2_p & !v1445872;
assign v121625b = hbusreq1_p & v121625a | !hbusreq1_p & v1216715;
assign v14460e0 = hbusreq5 & v14460c9 | !hbusreq5 & v14460df;
assign v12afe77 = decide_p & v12afe73 | !decide_p & v12afe76;
assign d3088d = hbusreq5_p & d307fd | !hbusreq5_p & !d3088c;
assign v1445a84 = hgrant2_p & v1445a74 | !hgrant2_p & v1445a83;
assign v121609f = hbusreq3 & v121608b | !hbusreq3 & v121609e;
assign v138a3d5 = hgrant5_p & v845542 | !hgrant5_p & v138a3d4;
assign v12161dd = hbusreq5_p & v12161d6 | !hbusreq5_p & !v12161dc;
assign v121654b = hmaster2_p & v845542 | !hmaster2_p & v121654a;
assign v12afe3e = hbusreq5 & v12afdb5 | !hbusreq5 & v12afe3d;
assign v1215476 = hready_p & v12153c4 | !hready_p & v1215475;
assign v1668cd3 = hlock0_p & v1668cc4 | !hlock0_p & v845542;
assign v1215d39 = hgrant5_p & v1216a99 | !hgrant5_p & v12165a2;
assign v16a1d4b = hmaster0_p & v16a1d46 | !hmaster0_p & v16a1d4a;
assign v144611d = hmaster0_p & v1446079 | !hmaster0_p & v1445fea;
assign d30754 = hmaster0_p & d30753 | !hmaster0_p & d3072b;
assign a653bd = hgrant5_p & a653ab | !hgrant5_p & !a653bc;
assign d2fb0d = hgrant5_p & d2f97b | !hgrant5_p & !d2fb0c;
assign d308b1 = hgrant2_p & d30810 | !hgrant2_p & d30883;
assign v14459cc = hlock1 & v14459cb | !hlock1 & v14459c8;
assign v12150c8 = hmaster2_p & v12153d3 | !hmaster2_p & v12150c7;
assign v16a19b3 = hgrant2_p & v16a2059 | !hgrant2_p & v16a19b2;
assign d3076e = hlock2_p & d3076d | !hlock2_p & d30769;
assign v12ad8ed = hmaster1_p & v12af7f7 | !hmaster1_p & v12ad8ec;
assign v138a3fa = hgrant2_p & v138a3f9 | !hgrant2_p & v138a3ee;
assign v1446715 = hmaster1_p & v1446714 | !hmaster1_p & v1446436;
assign v12160d6 = hmaster0_p & v12160d4 | !hmaster0_p & v12160d5;
assign v134cd5f = hbusreq0_p & v134d273 | !hbusreq0_p & v134cd55;
assign v1215059 = hmaster1_p & v1215058 | !hmaster1_p & v121546f;
assign v1553238 = hmaster0_p & v155322d | !hmaster0_p & v1553237;
assign v134d1f0 = hbusreq1 & v134d1e8 | !hbusreq1 & v134d1ef;
assign v140586a = hbusreq5_p & v1405866 | !hbusreq5_p & v1405869;
assign v1553398 = hlock0 & v1553397 | !hlock0 & v1553396;
assign a656d2 = hready_p & a656d1 | !hready_p & a65b20;
assign v1445a21 = hlock4 & v14459a8 | !hlock4 & v14459a7;
assign v13897df = hlock5_p & v13897de | !hlock5_p & !v845542;
assign d3076f = hbusreq2_p & d3076e | !hbusreq2_p & d30769;
assign v1445e05 = hmaster2_p & v1446427 | !hmaster2_p & v1445e04;
assign v12161f7 = hmaster2_p & f2f2a8 | !hmaster2_p & !v12161d8;
assign v12160e8 = hmaster0_p & v1215ff2 | !hmaster0_p & v1215ff0;
assign v12acff7 = hmaster1_p & v12acff6 | !hmaster1_p & v12ad65b;
assign v15168a5 = hmaster0_p & v845542 | !hmaster0_p & v1668c4a;
assign d3064e = hbusreq1 & a66295 | !hbusreq1 & !d305de;
assign v131be8d = hgrant2_p & v84555c | !hgrant2_p & v131be8a;
assign v12ad509 = hmaster0_p & v12ad508 | !hmaster0_p & v845542;
assign f2f458 = hgrant2_p & f2f3ae | !hgrant2_p & f2f443;
assign a6566e = hgrant5_p & a65424 | !hgrant5_p & !a6563c;
assign v134d52c = hready_p & v134d4e4 | !hready_p & v134d52b;
assign v121612d = hlock5_p & v121612b | !hlock5_p & v121612c;
assign v16a1ada = hbusreq1_p & v16a206e | !hbusreq1_p & v16a1ad9;
assign v144601a = hmaster2_p & v845542 | !hmaster2_p & v144600d;
assign d30651 = hgrant1_p & d30650 | !hgrant1_p & d30649;
assign v134cf6a = decide_p & v134d3fa | !decide_p & v134d3b5;
assign v12162cb = hgrant2_p & v12162c8 | !hgrant2_p & v12162ca;
assign v121652b = hgrant1_p & v1216522 | !hgrant1_p & v121652a;
assign v1215065 = hgrant5_p & v1215463 | !hgrant5_p & v1215064;
assign v134ce47 = hmaster1_p & v134d369 | !hmaster1_p & v134ce46;
assign v15156fb = hmaster0_p & v15156fa | !hmaster0_p & v151564f;
assign a653a3 = hgrant1_p & a6539b | !hgrant1_p & !a653a2;
assign v1446052 = hgrant5_p & v144604d | !hgrant5_p & v1446051;
assign v16a1a83 = hgrant5_p & v845542 | !hgrant5_p & !v16a1a79;
assign v1215ba5 = hmaster1_p & v1215ba4 | !hmaster1_p & !v1215ba1;
assign f2f2ae = hmaster0_p & f2f2ad | !hmaster0_p & f2f2a8;
assign d2feb9 = hlock1_p & d2feb8 | !hlock1_p & v84555a;
assign a65637 = hgrant1_p & a6539b | !hgrant1_p & !a65636;
assign v12160ad = hmaster0_p & v121606b | !hmaster0_p & v121604c;
assign a65630 = hmaster2_p & a6562a | !hmaster2_p & a6562e;
assign d302d4 = decide_p & v845542 | !decide_p & !v845570;
assign v12ad527 = hmaster2_p & v12ad514 | !hmaster2_p & a658c6;
assign v10d407b = hgrant5_p & v10d3fe8 | !hgrant5_p & v10d407a;
assign v14460fc = hlock2 & v14460f9 | !hlock2 & v14460fb;
assign v134d205 = hbusreq4_p & v134d204 | !hbusreq4_p & v845542;
assign v1552f79 = hmaster2_p & v1552f6c | !hmaster2_p & v845542;
assign v138a008 = hgrant2_p & v845542 | !hgrant2_p & !v138a007;
assign v1446675 = hgrant2_p & v1446672 | !hgrant2_p & v1446674;
assign v1284cf5 = hgrant1_p & v1405849 | !hgrant1_p & !v1284cf4;
assign v12ad53a = hbusreq2 & v12ad52b | !hbusreq2 & v12ad539;
assign a658f6 = hbusreq2_p & a658f0 | !hbusreq2_p & a658f4;
assign v1215010 = hgrant0_p & v121500f | !hgrant0_p & !v845559;
assign v16a1955 = hgrant1_p & v84554d | !hgrant1_p & v16a1954;
assign v15530b7 = jx2_p & v1552fd8 | !jx2_p & v15530b6;
assign v11e5941 = hmaster0_p & v845542 | !hmaster0_p & v11e593b;
assign v1284ccf = hgrant5_p & v1284cca | !hgrant5_p & !v1284cce;
assign v1215762 = hgrant5_p & v1215ba0 | !hgrant5_p & v1215760;
assign v1668cc1 = stateA1_p & v156645f | !stateA1_p & v1668cc0;
assign v134d3cd = hmaster1_p & v134d3c3 | !hmaster1_p & v134d23c;
assign v1446218 = hlock0 & v1446217 | !hlock0 & v14463b8;
assign v12acff0 = hready_p & v12ad66a | !hready_p & !v12acfef;
assign v15167fc = hgrant2_p & v15167fb | !hgrant2_p & !v845542;
assign v1668c76 = hbusreq1 & a658b5 | !hbusreq1 & !a65469;
assign a6562a = hgrant1_p & a65362 | !hgrant1_p & !a65628;
assign d2f9c8 = hmaster2_p & d2f9b7 | !hmaster2_p & d2f98c;
assign v1446278 = hmaster2_p & v1446439 | !hmaster2_p & v1446410;
assign v138a47b = hmaster1_p & v138a47a | !hmaster1_p & v138a3e0;
assign v14457b9 = hbusreq2 & v14457b3 | !hbusreq2 & v14457b4;
assign v1445a40 = hmaster2_p & v14459a0 | !hmaster2_p & v1445a02;
assign v12153f5 = hmaster1_p & v12153f4 | !hmaster1_p & v12153ec;
assign v1446118 = hmaster0_p & v1446079 | !hmaster0_p & v1446404;
assign v1668c43 = hmaster2_p & v1668c3f | !hmaster2_p & v845542;
assign v10d402d = hbusreq4_p & v10d3fe0 | !hbusreq4_p & v10d3fdf;
assign v1445ab0 = hmaster0_p & v14458a6 | !hmaster0_p & v144639c;
assign v144605c = hbusreq1_p & v144605b | !hbusreq1_p & v1446429;
assign v1284cc5 = hgrant0_p & v140583c | !hgrant0_p & !v140588e;
assign v1445a45 = hmaster1_p & v1445a44 | !hmaster1_p & v1445a32;
assign d2fc07 = hmaster1_p & d2fc06 | !hmaster1_p & d2fb55;
assign v1214c0d = hmaster1_p & v1214bb7 | !hmaster1_p & v12153a9;
assign a658c1 = hburst1 & v10d3fde | !hburst1 & !v845542;
assign v12153d5 = hready & v845542 | !hready & !v15168aa;
assign v14459b0 = hbusreq0_p & v14459af | !hbusreq0_p & v14465bb;
assign v14453fd = hlock3 & v14453f5 | !hlock3 & v14453fc;
assign v1552d9c = decide_p & v845542 | !decide_p & v1552d9b;
assign v14459fb = hbusreq1_p & v14465b2 | !hbusreq1_p & v14459fa;
assign a65670 = hbusreq0 & a6566d | !hbusreq0 & a6566f;
assign v138a3a9 = hlock2_p & v138a3a7 | !hlock2_p & v138a3a8;
assign v1216ac3 = hmaster2_p & v845542 | !hmaster2_p & v1216abe;
assign v12ad621 = hbusreq2_p & v12ad619 | !hbusreq2_p & v12ad620;
assign v1214f5a = hmaster1_p & v1214f4e | !hmaster1_p & !v1215d9b;
assign v13895a5 = decide_p & v13895a4 | !decide_p & v845542;
assign v1446074 = hmaster1_p & v144603f | !hmaster1_p & v1446073;
assign v1214cc9 = hbusreq1_p & v1214cbd | !hbusreq1_p & v1214cbb;
assign v1445845 = hmaster1_p & v1445eba | !hmaster1_p & v1445f09;
assign v1215041 = hbusreq5_p & v121503c | !hbusreq5_p & !v1215040;
assign v15534eb = hbusreq1 & v155338c | !hbusreq1 & v1553217;
assign v1668cc6 = hbusreq1_p & v1668cc5 | !hbusreq1_p & !v845542;
assign v1446608 = hgrant4_p & v1446606 | !hgrant4_p & v1446607;
assign v16a193f = hbusreq4_p & v16a193e | !hbusreq4_p & v845542;
assign v121546d = hbusreq4_p & v121546c | !hbusreq4_p & v845542;
assign v121679f = decide_p & v12164cd | !decide_p & v121679e;
assign d2fbe4 = hlock5_p & d2fbe2 | !hlock5_p & d2fbe3;
assign v1445f70 = hmaster1_p & v1446748 | !hmaster1_p & v14466a9;
assign v1446421 = hlock0_p & v1446403 | !hlock0_p & v1446420;
assign v14465ce = hgrant4_p & v1446407 | !hgrant4_p & v14465cd;
assign v10d40cc = hmaster1_p & v10d40cb | !hmaster1_p & v10d3fe9;
assign v1445db8 = hlock0 & v1445db7 | !hlock0 & v1445db6;
assign d30897 = hmaster2_p & d3088a | !hmaster2_p & d306aa;
assign v1405b2c = hmaster2_p & v1405b14 | !hmaster2_p & !v1405b1e;
assign v144551c = hmaster1_p & v1445506 | !hmaster1_p & v1445b5f;
assign v14461e0 = hmaster1_p & v1446163 | !hmaster1_p & v14460cf;
assign v16a1bfc = hbusreq0 & v16a209a | !hbusreq0 & v16a1bfb;
assign v138a330 = hbusreq1 & a658b5 | !hbusreq1 & !v138a32f;
assign v14466b8 = hmaster1_p & v1446664 | !hmaster1_p & v14466a9;
assign d2fe8d = hmaster1_p & d2fe82 | !hmaster1_p & d2fe8c;
assign v12ad1ff = hready_p & v12af7e2 | !hready_p & v12ad1fe;
assign v1445781 = hlock2 & v144577d | !hlock2 & v1445780;
assign v1553225 = hmaster2_p & v1553138 | !hmaster2_p & v845542;
assign v16a1e5c = hbusreq4_p & v845542 | !hbusreq4_p & v16a1e5b;
assign v138a3a0 = hbusreq2 & v138a397 | !hbusreq2 & v138a39f;
assign v1445b89 = hgrant5_p & v1445b73 | !hgrant5_p & v1445b57;
assign v15157fc = hgrant5_p & v15157fb | !hgrant5_p & v15157aa;
assign v1445bb9 = hmaster0_p & v1446636 | !hmaster0_p & v144643b;
assign v138a3f5 = hlock2_p & v138a3f2 | !hlock2_p & !v138a3f4;
assign v16a1a88 = hbusreq2_p & v16a196a | !hbusreq2_p & v16a1a87;
assign a6585f = hmaster0_p & a6585e | !hmaster0_p & a65852;
assign v16693a2 = hmaster1_p & v16693a1 | !hmaster1_p & a65893;
assign v14465e7 = hbusreq4_p & v1446403 | !hbusreq4_p & v144640c;
assign v1445f77 = hgrant2_p & v1445f5b | !hgrant2_p & v1445f76;
assign v10d40a1 = hmaster0_p & v10d407f | !hmaster0_p & v10d3feb;
assign v14459d3 = hbusreq1 & v14459ac | !hbusreq1 & v14459d2;
assign v16a1ac3 = hbusreq2 & v16a1abf | !hbusreq2 & v16a1ac2;
assign v16a1a75 = hbusreq4_p & v16a193e | !hbusreq4_p & v845572;
assign v134d463 = hlock3 & v134d276 | !hlock3 & v134d462;
assign d3012a = hlock2_p & d30127 | !hlock2_p & d30129;
assign d308fa = hbusreq3 & d308eb | !hbusreq3 & d308f7;
assign v15530ff = hbusreq2_p & v15530fe | !hbusreq2_p & v155321a;
assign v1214c12 = hmaster1_p & v1214bf9 | !hmaster1_p & v1214bcf;
assign v1284ca0 = stateG10_5_p & v1284c9f | !stateG10_5_p & !v1284c9e;
assign v1445f39 = hmaster0_p & v1445da7 | !hmaster0_p & v144639c;
assign v1446340 = hlock0 & v144633f | !hlock0 & v14466a6;
assign v1445511 = hlock3 & v14454fa | !hlock3 & v144550f;
assign d2fede = hlock2_p & d2fedd | !hlock2_p & d2fed9;
assign v12161f2 = hmaster2_p & v12161ee | !hmaster2_p & v12161f1;
assign v16a1af7 = hburst1 & v16a1af6 | !hburst1 & v845542;
assign d2fbcd = hlock4_p & d2fb4d | !hlock4_p & v84554a;
assign v134d396 = hgrant5_p & v845542 | !hgrant5_p & v134d395;
assign d2faf4 = hbusreq1_p & d300d7 | !hbusreq1_p & d2faf3;
assign v144610a = hmaster1_p & v14460f5 | !hmaster1_p & v1445fbd;
assign v1216a80 = hmaster0_p & v1216a7f | !hmaster0_p & v845542;
assign v1405a96 = hmaster2_p & v1405a86 | !hmaster2_p & v1405a87;
assign v1214ebd = hbusreq2 & v1214ebc | !hbusreq2 & v845542;
assign v16a1e28 = hmaster0_p & v16a1e23 | !hmaster0_p & v16a1e27;
assign v134ce94 = hbusreq2 & v134ce93 | !hbusreq2 & v134d240;
assign v1515628 = hmaster2_p & v845570 | !hmaster2_p & !v1515627;
assign v14459e1 = stateG10_5_p & v14459dc | !stateG10_5_p & v14459e0;
assign v134d22b = hlock0 & v134d22a | !hlock0 & v134d229;
assign v144622e = hbusreq5_p & v14463dc | !hbusreq5_p & v144622d;
assign v144539d = hgrant2_p & v144539c | !hgrant2_p & v1445398;
assign v1215cf4 = hbusreq0 & v1215cf0 | !hbusreq0 & v1215cf3;
assign a65624 = hmaster2_p & a65620 | !hmaster2_p & a65623;
assign v1553396 = hbusreq5_p & v1553392 | !hbusreq5_p & v1553395;
assign v12164d9 = hbusreq1_p & v845570 | !hbusreq1_p & v12164cf;
assign d2fc31 = hbusreq0 & d2fc30 | !hbusreq0 & d3069a;
assign v1445771 = hbusreq3 & v144576f | !hbusreq3 & v1445770;
assign v12ad543 = hlock2_p & v12ad540 | !hlock2_p & v12ad542;
assign v1284d27 = hbusreq2_p & v1284d21 | !hbusreq2_p & v1284d26;
assign d2f9d3 = hmaster1_p & d2f9b9 | !hmaster1_p & d2f9cb;
assign d301f1 = hmaster2_p & d307ac | !hmaster2_p & d301c5;
assign v134d1e2 = decide_p & v134d1e1 | !decide_p & v134d1e0;
assign v12150b7 = hmaster0_p & v1215773 | !hmaster0_p & v1215ba3;
assign v1515751 = hmaster2_p & v1515750 | !hmaster2_p & v1515749;
assign v134d3e8 = hgrant3_p & v134d3d8 | !hgrant3_p & v134d3e7;
assign v14461bb = hbusreq2_p & v144619e | !hbusreq2_p & v14461ba;
assign v16a1bb7 = hmastlock_p & v16a1bb6 | !hmastlock_p & v845542;
assign v1445370 = hmaster0_p & v1445909 | !hmaster0_p & v1445a6b;
assign v121653d = hbusreq0 & v1216533 | !hbusreq0 & v121653c;
assign d30790 = hbusreq1 & d3078f | !hbusreq1 & v845542;
assign v1405b34 = hgrant3_p & v1405acf | !hgrant3_p & v1405b33;
assign v16a169d = hbusreq5_p & v16a1d6b | !hbusreq5_p & v16a169c;
assign f2f461 = hbusreq3_p & f2f3e5 | !hbusreq3_p & f2f460;
assign v16a1dd2 = hbusreq2 & v16a1dc0 | !hbusreq2 & v16a1dc1;
assign d30680 = hbusreq5 & d30679 | !hbusreq5 & d3067f;
assign v10d42af = hlock0_p & v10d42ae | !hlock0_p & v10d3fd4;
assign v10d42bd = decide_p & v10d4009 | !decide_p & v10d42bc;
assign d3083a = hbusreq5_p & d30839 | !hbusreq5_p & d30838;
assign v121506b = hmaster0_p & v1215065 | !hmaster0_p & v1215030;
assign d30682 = hready_p & d30681 | !hready_p & d3063f;
assign v144641d = hbusreq4_p & v1446403 | !hbusreq4_p & v1446407;
assign v144642b = hbusreq5_p & v1446426 | !hbusreq5_p & v144642a;
assign v10d403e = hbusreq1_p & v10d3fe5 | !hbusreq1_p & !v10d3ff7;
assign d30761 = hmaster1_p & d3074b | !hmaster1_p & d30754;
assign d2fe96 = hmaster2_p & v845542 | !hmaster2_p & d2fe80;
assign v10d4060 = hgrant0_p & v10d3fdb | !hgrant0_p & !v10d3fd8;
assign v12acfe2 = hbusreq2_p & v12acfe0 | !hbusreq2_p & v12acfe1;
assign d308c0 = hbusreq5_p & d30821 | !hbusreq5_p & d308bf;
assign v1215778 = hgrant5_p & v1215ba3 | !hgrant5_p & !v1215776;
assign v12161a5 = hbusreq2_p & v121619e | !hbusreq2_p & !v12161a4;
assign v1445b26 = hbusreq2 & v1445b24 | !hbusreq2 & v1445b25;
assign v121600d = hmaster1_p & v1215ff3 | !hmaster1_p & v121600c;
assign v16a1387 = hmaster1_p & v16a1386 | !hmaster1_p & !v16a2672;
assign v1214bf0 = hmaster1_p & v12153b1 | !hmaster1_p & v1214bcf;
assign v1445516 = hmaster1_p & v14454fb | !hmaster1_p & v1446290;
assign v138a445 = hmaster1_p & v138a444 | !hmaster1_p & v84555c;
assign v1215042 = hbusreq0_p & v1215460 | !hbusreq0_p & !v1215032;
assign d3089d = hbusreq0 & d30899 | !hbusreq0 & d3089c;
assign v12160d8 = hbusreq1_p & v12160d7 | !hbusreq1_p & v845542;
assign v1389e37 = decide_p & v1389e36 | !decide_p & v138a406;
assign v15167ef = hbusreq5 & v15167c4 | !hbusreq5 & v15167ee;
assign v1215c2d = hbusreq5_p & v1215c2b | !hbusreq5_p & v1215c2c;
assign v144620b = jx2_p & v1445f84 | !jx2_p & v144620a;
assign v12acd06 = jx1_p & v12ad03d | !jx1_p & v12acd05;
assign v14460b6 = hmaster0_p & v14460b5 | !hmaster0_p & v1446072;
assign v14463b5 = hlock0_p & v144639c | !hlock0_p & !v14463b4;
assign v138a3ee = hmaster1_p & v138a3ed | !hmaster1_p & v138a3e0;
assign d308a8 = hgrant1_p & v84554c | !hgrant1_p & d308a7;
assign v1445f7f = hlock5 & v144673f | !hlock5 & v1445f7e;
assign v1216099 = hmaster2_p & v1216092 | !hmaster2_p & v121602d;
assign v10d4282 = hlock0_p & v10d4280 | !hlock0_p & v10d4281;
assign v12ad019 = hgrant2_p & v12acff7 | !hgrant2_p & v12ad018;
assign v144622c = stateG10_5_p & v144622b | !stateG10_5_p & !v144622a;
assign v16a1bc6 = hready & v845570 | !hready & v845542;
assign d306a7 = hgrant1_p & v84554c | !hgrant1_p & d306a6;
assign v16a1d91 = hgrant5_p & v845542 | !hgrant5_p & v16a2244;
assign v1446061 = hbusreq1_p & v14465f2 | !hbusreq1_p & v1446608;
assign bf1f5a = hlock2_p & v845570 | !hlock2_p & !bf1f59;
assign v1446748 = hmaster0_p & v1446663 | !hmaster0_p & v14465b8;
assign v155342c = hbusreq5_p & v1553150 | !hbusreq5_p & v155342b;
assign v1445866 = hlock5 & v14457f6 | !hlock5 & v1445865;
assign d2fec3 = hbusreq4_p & d2fec2 | !hbusreq4_p & v845542;
assign v1215b8c = hmaster1_p & v1215b8b | !hmaster1_p & v1215b88;
assign v121537c = hbusreq0_p & v16a1bc6 | !hbusreq0_p & v845542;
assign v1445fe0 = hmaster2_p & v144639c | !hmaster2_p & v1445fcc;
assign v16a1acd = hmaster1_p & v16a1acc | !hmaster1_p & !v16a1f96;
assign v1214da6 = decide_p & v1214d8b | !decide_p & v1214da5;
assign v134d428 = hmaster2_p & v134d427 | !hmaster2_p & v134d386;
assign v16a1bd2 = hgrant0_p & v845542 | !hgrant0_p & v16a1bc6;
assign v1446397 = hmastlock_p & v1446396 | !hmastlock_p & v845542;
assign v16a205f = hmaster1_p & v845568 | !hmaster1_p & v16a1f96;
assign v12ad953 = hready_p & v12af7e2 | !hready_p & v12ad952;
assign d3086c = hmaster2_p & d30867 | !hmaster2_p & d3086b;
assign v1214de1 = hbusreq2_p & v1214de0 | !hbusreq2_p & v845542;
assign v1445a1b = hmaster2_p & v1445a1a | !hmaster2_p & v144660f;
assign v1445481 = hbusreq2_p & v1445480 | !hbusreq2_p & v1445bba;
assign v1668d4a = hgrant4_p & v1668d49 | !hgrant4_p & a65862;
assign v1214f0c = hbusreq5_p & v1214f0b | !hbusreq5_p & v1214f0a;
assign v16a209f = hbusreq2 & v16a209d | !hbusreq2 & !v16a209e;
assign v14457dc = hgrant2_p & v14457d9 | !hgrant2_p & v14457db;
assign a64707 = decide_p & a64705 | !decide_p & a662a2;
assign v1446471 = hgrant1_p & v144646f | !hgrant1_p & v845542;
assign d30147 = hlock5_p & d30145 | !hlock5_p & d30146;
assign v1445817 = hbusreq2_p & v1445807 | !hbusreq2_p & v1445816;
assign a653c4 = hlock0_p & v10d3fd8 | !hlock0_p & a653c3;
assign v14463ef = hmaster0_p & v14463df | !hmaster0_p & v14463ee;
assign v134d4d2 = hbusreq4_p & v134d1dd | !hbusreq4_p & v134d4ca;
assign v1445991 = stateA1_p & v146d169 | !stateA1_p & v1445990;
assign v1405b24 = hgrant1_p & v1405ac4 | !hgrant1_p & !v1405b23;
assign v121576e = hbusreq5_p & v121576c | !hbusreq5_p & v121576d;
assign v121509e = hbusreq5_p & v121509a | !hbusreq5_p & v121509d;
assign v134d45e = hgrant3_p & v134d3fc | !hgrant3_p & v134d45d;
assign v121501e = hmaster0_p & v1214fed | !hmaster0_p & v121501d;
assign v134cd6f = hmaster2_p & v845542 | !hmaster2_p & v134cd6e;
assign v1215d97 = hmaster2_p & v12166e5 | !hmaster2_p & !v12164d9;
assign v121626d = hmaster0_p & v1216172 | !hmaster0_p & v121601e;
assign v1216068 = hmaster2_p & v1216049 | !hmaster2_p & v1216067;
assign v14058d8 = hmaster0_p & v14058cd | !hmaster0_p & v14058d7;
assign v151580e = hmaster1_p & v151580d | !hmaster1_p & v10d3ffb;
assign v1284d1b = hgrant4_p & v1446429 | !hgrant4_p & v1284d1a;
assign v1445a72 = hlock3 & v1445a69 | !hlock3 & v1445a71;
assign f2f45f = hready_p & f2f45d | !hready_p & f2f45e;
assign v14465ad = hmastlock_p & v14465ac | !hmastlock_p & v845542;
assign v16a1d03 = hgrant3_p & v16a1ce9 | !hgrant3_p & v16a1d02;
assign d3020c = hgrant5_p & d301c0 | !hgrant5_p & d3020b;
assign v144603b = hgrant4_p & v144639c | !hgrant4_p & v144603a;
assign v14453f9 = hbusreq3 & v14453f7 | !hbusreq3 & v14453f8;
assign v140586b = hlock4_p & v140583e | !hlock4_p & v14463b1;
assign v1389ffd = hbusreq5_p & v1389ffc | !hbusreq5_p & !v845542;
assign v1516801 = hbusreq2_p & v1516800 | !hbusreq2_p & !v845542;
assign v1445e68 = hgrant4_p & v1445dec | !hgrant4_p & v1445e67;
assign v1668d35 = hgrant4_p & v1668d26 | !hgrant4_p & a65851;
assign v1445a6d = hmaster1_p & v1445a6c | !hmaster1_p & v14458fd;
assign v15167f8 = hbusreq5_p & v15167f7 | !hbusreq5_p & v845542;
assign v1445919 = hbusreq0 & v1445918 | !hbusreq0 & v14458ee;
assign v12ad65b = hmaster0_p & v12ad643 | !hmaster0_p & v12ad65a;
assign v12af229 = hmaster1_p & v12af9c3 | !hmaster1_p & v12af228;
assign v151699e = hlock3_p & v1516988 | !hlock3_p & v151699d;
assign d2fbd2 = hgrant1_p & d2fbcb | !hgrant1_p & d2fbd1;
assign d2fbb3 = hlock2_p & d2fbb1 | !hlock2_p & d2fbb2;
assign v14453ff = hlock5 & v14453f9 | !hlock5 & v14453fe;
assign v121607b = hbusreq2_p & v121607a | !hbusreq2_p & v1216079;
assign v144621c = hlock0 & v144621b | !hlock0 & v14463c4;
assign a65433 = hbusreq5_p & a6542f | !hbusreq5_p & a65431;
assign v134d514 = hmaster1_p & v134d369 | !hmaster1_p & v134d513;
assign v15156ef = hbusreq3 & v15156e9 | !hbusreq3 & v15156ee;
assign v1445374 = hlock2 & v1445354 | !hlock2 & v1445373;
assign v1445385 = hgrant2_p & v1445383 | !hgrant2_p & v1445384;
assign v134d42b = hbusreq1 & v134d391 | !hbusreq1 & v134d385;
assign a66297 = hbusreq4_p & a66296 | !hbusreq4_p & !v845542;
assign v1552f6e = hbusreq0 & v1552f6d | !hbusreq0 & v1553218;
assign v155304d = hlock0_p & v155338c | !hlock0_p & v155304c;
assign v155350b = decide_p & v1553216 | !decide_p & v155350a;
assign v1445e26 = hbusreq0 & v1445e25 | !hbusreq0 & v1445df8;
assign v1216249 = hgrant5_p & v1216248 | !hgrant5_p & !v12161db;
assign v14460ea = hbusreq2_p & v14460e8 | !hbusreq2_p & v14460e9;
assign v12166f4 = hmaster0_p & v12164d7 | !hmaster0_p & v12166f3;
assign v16a1d59 = hgrant5_p & v845542 | !hgrant5_p & !v16a1d3d;
assign v1405922 = hgrant2_p & v140591f | !hgrant2_p & v1405921;
assign d308f4 = hlock5_p & d308f3 | !hlock5_p & v84554e;
assign v1389fb9 = hbusreq5_p & v1389fb8 | !hbusreq5_p & v845542;
assign d2fbdc = hmaster2_p & d2fb4e | !hmaster2_p & d2fb4d;
assign v14458ab = hmaster0_p & v144639c | !hmaster0_p & v14458aa;
assign v15530b2 = hready_p & v1553427 | !hready_p & v15530b1;
assign v12ad51d = hmaster2_p & v12ad515 | !hmaster2_p & v12ad51c;
assign d30123 = hlock4_p & v845542 | !hlock4_p & !v1668c1c;
assign v15530ac = hbusreq2 & v15530aa | !hbusreq2 & v15530ab;
assign v1445e24 = hmaster2_p & v1445e10 | !hmaster2_p & v1445def;
assign v144554b = hready_p & v1446564 | !hready_p & v144554a;
assign v14457db = hmaster1_p & v14457da | !hmaster1_p & v1445eaa;
assign v1445439 = hbusreq3 & v1445437 | !hbusreq3 & v1445438;
assign v16a1405 = hgrant2_p & v845542 | !hgrant2_p & !v16a1404;
assign f2e4da = hbusreq5_p & f2f539 | !hbusreq5_p & f2e4d9;
assign d80770 = hmaster2_p & d80733 | !hmaster2_p & !v845542;
assign v15534d4 = hbusreq1 & v15533ad | !hbusreq1 & v15533a1;
assign v10d42d7 = hmaster0_p & v10d42b8 | !hmaster0_p & v10d42b4;
assign v1668da0 = hbusreq5_p & v1668d9e | !hbusreq5_p & v1668d9f;
assign v1445fd7 = hbusreq1_p & v144641d | !hbusreq1_p & v1446427;
assign v1214ec3 = hmaster1_p & v1214ec2 | !hmaster1_p & v1215d68;
assign v155308e = hgrant2_p & v155308d | !hgrant2_p & v1553060;
assign v1446087 = hbusreq1_p & v1446086 | !hbusreq1_p & v14465bb;
assign v15534f9 = hmaster2_p & v15534ec | !hmaster2_p & v845542;
assign v12ad5a0 = busreq_p & v10d4264 | !busreq_p & !v12ad59f;
assign v15167f1 = hready_p & v845542 | !hready_p & v15167f0;
assign v144586e = hbusreq0_p & v144639c | !hbusreq0_p & v144639e;
assign v144664c = hmaster1_p & v144664b | !hmaster1_p & v1446630;
assign v1284c9d = hlock5_p & v1284c9b | !hlock5_p & !v1284c9c;
assign v14465d9 = hbusreq1_p & v144639c | !hbusreq1_p & v14465bb;
assign v1515711 = hbusreq1 & v10d3fd4 | !hbusreq1 & !v845542;
assign v10d4035 = hmaster2_p & v10d3fef | !hmaster2_p & v10d3ff3;
assign v14466f9 = hmaster0_p & v1446638 | !hmaster0_p & v1446404;
assign a65437 = hbusreq5_p & a65434 | !hbusreq5_p & a65436;
assign v1446634 = hbusreq1 & v14465be | !hbusreq1 & v1446633;
assign v1215302 = hbusreq5 & v12152f4 | !hbusreq5 & v1215301;
assign v14463e8 = hbusreq1 & v14463e6 | !hbusreq1 & v14463e7;
assign v1445b6f = hgrant2_p & v1445b6e | !hgrant2_p & v1445b6a;
assign d3029a = hbusreq2 & d30297 | !hbusreq2 & d30299;
assign v14463f7 = hmaster0_p & v144639c | !hmaster0_p & v14463f6;
assign v1516200 = hlock3_p & v15161d7 | !hlock3_p & v15161ff;
assign v1389372 = hbusreq5 & v1389f87 | !hbusreq5 & v1389371;
assign v1445876 = stateG10_5_p & v1445875 | !stateG10_5_p & !v1445874;
assign v12ad5f8 = hbusreq0 & v12ad5f7 | !hbusreq0 & !v845542;
assign v1214efe = hbusreq2_p & v1214efd | !hbusreq2_p & v845542;
assign v1284d2e = hmaster0_p & v1284d00 | !hmaster0_p & v1405859;
assign v1445e71 = hmaster2_p & v1445e70 | !hmaster2_p & v1445def;
assign v1668cec = hbusreq2_p & v1668cd7 | !hbusreq2_p & v1668ceb;
assign v1216289 = hmaster1_p & v1216288 | !hmaster1_p & !v1216027;
assign d2fc81 = hbusreq3_p & d2fc22 | !hbusreq3_p & d2fc80;
assign v12162c8 = hmaster1_p & v12162c7 | !hmaster1_p & v12160e0;
assign v16a2099 = hbusreq2 & v16a2097 | !hbusreq2 & !v16a2098;
assign d307cb = hlock1_p & d307ca | !hlock1_p & d30658;
assign v16695c4 = decide_p & v16695bb | !decide_p & v845542;
assign v16a1ca8 = hgrant2_p & v16a205c | !hgrant2_p & v16a1ca7;
assign d2fd10 = hlock2_p & v845542 | !hlock2_p & !d2fd0f;
assign f2ed97 = hmaster0_p & f2ed96 | !hmaster0_p & f2ed95;
assign v134d227 = hbusreq2_p & v134d226 | !hbusreq2_p & v134d225;
assign v1445fbe = hmaster1_p & v144639c | !hmaster1_p & v1445fbd;
assign d30636 = hlock2_p & d30634 | !hlock2_p & d30635;
assign v12ad5e3 = hgrant2_p & v12ad597 | !hgrant2_p & v12ad5e2;
assign d305d7 = hbusreq5_p & d305d6 | !hbusreq5_p & v845542;
assign v1445fa9 = hlock0 & v1445fa8 | !hlock0 & v1445fa7;
assign v1216072 = hmaster1_p & v1216071 | !hmaster1_p & v121605d;
assign v1445bb1 = hmaster0_p & v1445bb0 | !hmaster0_p & v14463bc;
assign v12166c9 = hmastlock_p & d30788 | !hmastlock_p & !v845542;
assign bf1f94 = hbusreq5_p & bf1f5d | !hbusreq5_p & !bf1f93;
assign v12ad13f = hbusreq2 & v12ad13e | !hbusreq2 & v12afe72;
assign v1405ac3 = hbusreq5_p & v1405ac1 | !hbusreq5_p & v1405ac2;
assign a658bc = hburst0 & v156645f | !hburst0 & a658bb;
assign v121628a = hmaster1_p & v121617d | !hmaster1_p & v121616f;
assign v121658c = stateG3_2_p & v845542 | !stateG3_2_p & v1216a86;
assign v1214fff = hmaster2_p & v1214ffe | !hmaster2_p & v1214ff7;
assign v16a19c2 = hgrant2_p & v16a205f | !hgrant2_p & v16a19c1;
assign v1389448 = hbusreq5_p & v1389447 | !hbusreq5_p & v845542;
assign v134d1df = hmaster0_p & v134d1de | !hmaster0_p & v845542;
assign v121656d = hmaster2_p & v1216566 | !hmaster2_p & v121656c;
assign v1216af9 = hmaster1_p & v1216ab3 | !hmaster1_p & v1216af8;
assign d2fc60 = hmaster2_p & d2fc5e | !hmaster2_p & d2fc5f;
assign v134d389 = hgrant1_p & v845542 | !hgrant1_p & v134d380;
assign d3069e = hmaster1_p & d3069a | !hmaster1_p & d3069d;
assign f2e4d2 = hgrant2_p & v845542 | !hgrant2_p & f2e4d1;
assign v1215758 = hbusreq0_p & v845547 | !hbusreq0_p & v1216136;
assign v12ad5dc = hmaster2_p & v12ad5db | !hmaster2_p & v12afe46;
assign v1405879 = hlock2_p & v1405877 | !hlock2_p & v1405878;
assign v1214d70 = hmaster1_p & v1214d6f | !hmaster1_p & v1214c39;
assign f2f2d0 = hmaster2_p & f2f2cf | !hmaster2_p & f2f21f;
assign v1215da8 = hbusreq2_p & v1215da5 | !hbusreq2_p & v1215da1;
assign v12152ee = hmaster1_p & v121577e | !hmaster1_p & v1215770;
assign v1445b85 = hbusreq2 & v1445b83 | !hbusreq2 & v1445b84;
assign d2f994 = hbusreq0 & d2fec1 | !hbusreq0 & d2f993;
assign v1445b3f = hmaster1_p & v1445b3e | !hmaster1_p & v14458fd;
assign v1445abd = hmaster1_p & v1445abc | !hmaster1_p & v14458af;
assign v1214d0b = hmaster2_p & v1214cec | !hmaster2_p & v1214cf9;
assign v12af220 = hbusreq1_p & v12afe45 | !hbusreq1_p & v12af9d1;
assign d307f1 = hlock5_p & d307ef | !hlock5_p & d307f0;
assign v1214d4b = hmaster0_p & v1214d45 | !hmaster0_p & v1214d4a;
assign v1215330 = hgrant2_p & v121531f | !hgrant2_p & v121532f;
assign v1216a60 = locked_p & v1216a5f | !locked_p & v845542;
assign v1445fc4 = hlock2 & v1445fb2 | !hlock2 & v1445fc2;
assign v12ad03c = hbusreq3_p & v12ad630 | !hbusreq3_p & v12ad03b;
assign v138a461 = hmaster1_p & v138a354 | !hmaster1_p & v138a341;
assign v1445a5a = hlock0 & v1445a56 | !hlock0 & v1445a59;
assign v166939c = hmaster2_p & v845570 | !hmaster2_p & v166939b;
assign v1215d8e = hbusreq2_p & v1215d8b | !hbusreq2_p & v1215d83;
assign v121482d = jx1_p & v1214dcb | !jx1_p & v121482c;
assign v1216a99 = hmaster2_p & v1216a96 | !hmaster2_p & v1216a98;
assign v134ce8b = hbusreq1_p & v134d1e8 | !hbusreq1_p & v134ce8a;
assign d2fb7c = hmaster1_p & d2fb6c | !hmaster1_p & d2fb7b;
assign d2fed7 = hmaster1_p & d2fed6 | !hmaster1_p & d2fec6;
assign v1668dba = hgrant5_p & v845570 | !hgrant5_p & v1668d37;
assign v12ad558 = hbusreq2 & v12ad552 | !hbusreq2 & v12ad557;
assign v1552f8c = hready_p & v1553306 | !hready_p & v1552f8b;
assign v1445836 = hmaster1_p & v1445ecc | !hmaster1_p & v1445ef0;
assign v12160fc = hgrant4_p & v12160fa | !hgrant4_p & v12160fb;
assign v1405ab2 = hmaster1_p & v1405ab1 | !hmaster1_p & v1405aae;
assign v1445fa0 = hmaster2_p & v144639c | !hmaster2_p & v1445f87;
assign v1515600 = hlock2_p & v15155ff | !hlock2_p & !v845542;
assign v15155f6 = hbusreq2_p & v15155f5 | !hbusreq2_p & !v845542;
assign v1553239 = hmaster1_p & v1553224 | !hmaster1_p & v1553238;
assign v121630f = hlock2_p & v121630e | !hlock2_p & v12162f8;
assign d306ec = hburst1_p & v845542 | !hburst1_p & d306eb;
assign v15156ea = hmaster1_p & v15156bd | !hmaster1_p & !v15156da;
assign v1216707 = hbusreq2 & v12166fb | !hbusreq2 & v1216706;
assign d2fb90 = hmaster1_p & d2fb8f | !hmaster1_p & d2fb7b;
assign v15168ee = hgrant2_p & v15168ed | !hgrant2_p & !v845542;
assign v10d40b2 = hmaster0_p & v10d3ffd | !hmaster0_p & v10d3ff0;
assign d307a0 = hgrant1_p & v845542 | !hgrant1_p & d3079f;
assign v10a1542 = hready_p & v10a1541 | !hready_p & !v845564;
assign d2fc48 = hready_p & d2fc2a | !hready_p & d2fc47;
assign v1216537 = hgrant4_p & v1216524 | !hgrant4_p & v845542;
assign d300eb = hgrant5_p & d300e4 | !hgrant5_p & d300ea;
assign v1445ee4 = hlock2 & v1445edb | !hlock2 & v1445ee3;
assign v1215750 = hgrant1_p & v1215746 | !hgrant1_p & v845542;
assign v12ad575 = hmaster1_p & v12ad574 | !hmaster1_p & !v12ad525;
assign v134cea0 = hbusreq2_p & v134ce9f | !hbusreq2_p & v134d23e;
assign v144630b = hgrant5_p & v144643a | !hgrant5_p & v144630a;
assign a64719 = jx0_p & a65b40 | !jx0_p & a64717;
assign f2f385 = hmaster2_p & f2f382 | !hmaster2_p & f2f384;
assign v1446229 = hbusreq2 & v1446222 | !hbusreq2 & v1446228;
assign v1445453 = hmaster1_p & v1445447 | !hmaster1_p & v1446250;
assign v1215b7b = hbusreq4_p & v1215b7a | !hbusreq4_p & v845542;
assign v134d373 = hbusreq1_p & v134d273 | !hbusreq1_p & v134d372;
assign v1445aa7 = hlock2 & v1445a69 | !hlock2 & v1445aa6;
assign d2feed = hbusreq2 & d2fee9 | !hbusreq2 & d2feec;
assign v16a16aa = hmaster1_p & v16a16a9 | !hmaster1_p & v16a209c;
assign v14463d7 = hlock4 & v144639c | !hlock4 & v14463d6;
assign v1389458 = hbusreq2 & v1389451 | !hbusreq2 & v138a391;
assign v144618d = hmaster0_p & v1445fea | !hmaster0_p & v144608a;
assign v121534d = hbusreq0 & v121534c | !hbusreq0 & v845542;
assign v121604b = hbusreq1_p & v121604a | !hbusreq1_p & v845542;
assign v1446017 = hmaster0_p & v1446010 | !hmaster0_p & v1446016;
assign v134d534 = hmaster1_p & v134d533 | !hmaster1_p & v845542;
assign v16a1ca1 = hmaster1_p & v16a1ca0 | !hmaster1_p & !v16a2672;
assign v1445a17 = hgrant4_p & v1445a15 | !hgrant4_p & v1445a16;
assign v134cdc5 = hbusreq2 & v134cdc3 | !hbusreq2 & v134cdc4;
assign v134d391 = hgrant4_p & v845542 | !hgrant4_p & v134d390;
assign v1214f19 = hbusreq2_p & v1214f18 | !hbusreq2_p & v845542;
assign v12af9b6 = hbusreq2_p & v12afe3d | !hbusreq2_p & v12af9b5;
assign v134cd8c = hbusreq5 & v134cd8a | !hbusreq5 & v134cd8b;
assign v15534d8 = hgrant5_p & v845542 | !hgrant5_p & v15534d7;
assign v1214d4e = hbusreq1_p & v1215364 | !hbusreq1_p & v121536a;
assign v14458f6 = hbusreq4_p & v1446403 | !hbusreq4_p & v14458e2;
assign d302f6 = hgrant3_p & d302f2 | !hgrant3_p & d302f5;
assign v121618b = hbusreq2 & v1216181 | !hbusreq2 & v121618a;
assign v138938b = hgrant5_p & v138938a | !hgrant5_p & v845542;
assign v1668ca7 = hbusreq2_p & v1668c9d | !hbusreq2_p & v1668ca6;
assign v12165ac = hmaster2_p & v1216588 | !hmaster2_p & v845570;
assign v16693aa = hmastlock_p & a658a5 | !hmastlock_p & v845542;
assign d30114 = hmaster2_p & d300be | !hmaster2_p & d300e9;
assign v14463eb = hbusreq0 & v14463ea | !hbusreq0 & v14463bf;
assign v12af1bd = hmaster2_p & d30690 | !hmaster2_p & v12af1bc;
assign a653ec = hmaster0_p & a65360 | !hmaster0_p & a653ea;
assign v1216244 = hgrant2_p & v1216234 | !hgrant2_p & v1216243;
assign v134d242 = hmaster0_p & v134d20a | !hmaster0_p & v134d1e8;
assign v1668e03 = hgrant3_p & v1668d14 | !hgrant3_p & !v1668e02;
assign v121639a = hbusreq5 & v1216314 | !hbusreq5 & v1216399;
assign v1445361 = hmaster0_p & v1445a5a | !hmaster0_p & v14459a3;
assign v12160d1 = hbusreq1_p & v12160d0 | !hbusreq1_p & v845547;
assign v16a1e93 = hgrant0_p & v845542 | !hgrant0_p & !v16a1e5b;
assign v1215419 = hmaster1_p & v12153fb | !hmaster1_p & v121540f;
assign v12ad57d = hbusreq2_p & v12ad57a | !hbusreq2_p & v12ad57c;
assign v121539f = hmaster2_p & v845547 | !hmaster2_p & v121539d;
assign d2ff04 = hlock2_p & d2ff02 | !hlock2_p & d2ff03;
assign v1405abe = hmaster0_p & v1405abc | !hmaster0_p & v1405abd;
assign d30730 = hmaster1_p & d3072f | !hmaster1_p & d3072c;
assign v1389e26 = hlock5_p & v1389e25 | !hlock5_p & !v845542;
assign v151582d = hbusreq2 & v151582c | !hbusreq2 & v15167ed;
assign v134ce66 = hbusreq2_p & v134ce64 | !hbusreq2_p & v134ce65;
assign v10d40c5 = hmaster1_p & v10d40c4 | !hmaster1_p & !v10d404f;
assign v1405938 = hmaster1_p & v1405937 | !hmaster1_p & v140584d;
assign v1389f8c = hlock5_p & v1389f8b | !hlock5_p & v845542;
assign v16a1d44 = hmaster0_p & v16a1d3f | !hmaster0_p & v16a1d43;
assign a65893 = hmaster0_p & a6587e | !hmaster0_p & a65892;
assign v10d42c0 = hmaster0_p & v10d4275 | !hmaster0_p & v10d426f;
assign v11e5982 = hgrant3_p & v11e5972 | !hgrant3_p & v11e5981;
assign v16a1e65 = hmaster1_p & v16a1e64 | !hmaster1_p & v16a2672;
assign d300e5 = hbusreq1 & d2fe84 | !hbusreq1 & d2fe80;
assign a653f0 = hbusreq5_p & a653ed | !hbusreq5_p & !a653ef;
assign v134cea9 = hbusreq5 & v134ce96 | !hbusreq5 & v134cea8;
assign v134cecb = hlock5 & v134cec6 | !hlock5 & v134ceca;
assign v134d4dc = hmaster0_p & v134d4d1 | !hmaster0_p & v134d4db;
assign v16a1840 = hmaster2_p & v16a183f | !hmaster2_p & v845542;
assign a654b2 = hmaster1_p & a658e8 | !hmaster1_p & !a654b0;
assign v14058d5 = hgrant1_p & v140584b | !hgrant1_p & v14058d4;
assign v12af3a7 = hlock1_p & v12af3a6 | !hlock1_p & d30727;
assign v14458cd = hlock3 & v14458b3 | !hlock3 & v14458cc;
assign v14462f5 = hlock0 & v14462f4 | !hlock0 & v14462ef;
assign v1214f5e = hmaster1_p & v1214f54 | !hmaster1_p & !v1215d9b;
assign v1214c75 = hmaster1_p & v1214c56 | !hmaster1_p & v1214c74;
assign v1446308 = hmaster0_p & v14462e6 | !hmaster0_p & v1446304;
assign a65af3 = hgrant2_p & v845542 | !hgrant2_p & a65af2;
assign v16a1437 = hgrant4_p & v845559 | !hgrant4_p & v845572;
assign v16a1e04 = decide_p & v16a1dda | !decide_p & !v16a1e03;
assign v121616e = hbusreq0 & v121615a | !hbusreq0 & v121616d;
assign v1215321 = hmaster1_p & v1215320 | !hmaster1_p & v1215054;
assign a654b6 = hmaster1_p & a6548f | !hmaster1_p & !a654b0;
assign v12162fb = hlock1_p & v12162fa | !hlock1_p & v845547;
assign v12153ce = hlock4_p & v12153cd | !hlock4_p & !v845542;
assign v15157e6 = hgrant5_p & v1668dc2 | !hgrant5_p & v151574a;
assign a658cb = hbusreq4_p & a658ca | !hbusreq4_p & !v845542;
assign d300d1 = hlock5_p & d300cf | !hlock5_p & !d300d0;
assign v144543f = hmaster0_p & v14464a4 | !hmaster0_p & v845542;
assign v134d22f = hmaster1_p & v134d22e | !hmaster1_p & v134d208;
assign d2fb25 = hgrant5_p & d2f981 | !hgrant5_p & !d2fb05;
assign v138a091 = hready_p & v138a07f | !hready_p & v138a090;
assign v14463a5 = hbusreq1_p & v144639c | !hbusreq1_p & v144639e;
assign v16a1942 = hmaster2_p & v16a1941 | !hmaster2_p & v16a206f;
assign v16a1bdb = hmaster0_p & v16a1bd1 | !hmaster0_p & v16a1bda;
assign f2f294 = hbusreq1 & a6585c | !hbusreq1 & v845542;
assign v1445544 = hmaster0_p & v1445543 | !hmaster0_p & v1446616;
assign v1553096 = hgrant5_p & v1553095 | !hgrant5_p & v1553052;
assign v1215da4 = hmaster1_p & v1215d89 | !hmaster1_p & !v1215d9b;
assign v14058e3 = hbusreq2_p & v14058da | !hbusreq2_p & v14058e2;
assign v134ce40 = hlock1 & v134d380 | !hlock1 & v134ce3f;
assign v144668d = hmaster2_p & v14465b3 | !hmaster2_p & v144668c;
assign d308af = hgrant2_p & d30886 | !hgrant2_p & !d308ae;
assign bf1f60 = hmaster2_p & d3064a | !hmaster2_p & bf1f5f;
assign d2fad1 = hlock2_p & d2face | !hlock2_p & !d2fad0;
assign d30604 = hmaster2_p & a66278 | !hmaster2_p & !d30603;
assign v14465b3 = hgrant1_p & v1446403 | !hgrant1_p & v14465b2;
assign d30773 = hlock2_p & d30771 | !hlock2_p & d30772;
assign v12160fd = hbusreq1 & v12160fc | !hbusreq1 & v845542;
assign v16a13f0 = hmaster0_p & v16a13ed | !hmaster0_p & v16a13ef;
assign d2fef3 = hlock2_p & d2fef2 | !hlock2_p & d2feef;
assign d30641 = hmaster0_p & d305d7 | !hmaster0_p & d305d5;
assign d300be = hgrant1_p & d300b8 | !hgrant1_p & d300bd;
assign v1216234 = hmaster1_p & v1216233 | !hmaster1_p & v12160e0;
assign v1668c6b = hmastlock_p & v1668c6a | !hmastlock_p & !v845542;
assign v1284cda = hgrant0_p & v1284cd9 | !hgrant0_p & !v140584b;
assign f2e504 = jx2_p & f2e503 | !jx2_p & f2eda3;
assign v12afe5b = hgrant4_p & v845542 | !hgrant4_p & v12afe5a;
assign v1445a37 = hbusreq0 & v1445a35 | !hbusreq0 & v1445a36;
assign v134d3c3 = hbusreq5_p & v134d20a | !hbusreq5_p & v134d3c2;
assign v134d1d9 = stateG3_0_p & v845542 | !stateG3_0_p & !v845586;
assign v1445a55 = hgrant5_p & v1445907 | !hgrant5_p & v1445a54;
assign a65910 = hbusreq2 & a658ff | !hbusreq2 & a6590f;
assign v1445b5c = hbusreq5_p & v14462ea | !hbusreq5_p & v1445b58;
assign v134ce81 = hbusreq1_p & v134d1e8 | !hbusreq1_p & v134d1ea;
assign v134d37b = hbusreq0 & v134d37a | !hbusreq0 & v134d379;
assign v12af9d2 = hbusreq1_p & v12afe61 | !hbusreq1_p & v12af9d1;
assign d2fb3b = hbusreq0 & d2f9a3 | !hbusreq0 & d2fb3a;
assign v16a19a5 = hbusreq4_p & v16a19a4 | !hbusreq4_p & v845542;
assign v12162f1 = hbusreq5_p & v12162f0 | !hbusreq5_p & v12162ef;
assign v12ad020 = hbusreq2 & v12ad01a | !hbusreq2 & v12ad01f;
assign v1215445 = hmaster1_p & v12153ee | !hmaster1_p & v12153ec;
assign d2f974 = hbusreq5_p & d2fea4 | !hbusreq5_p & d2f973;
assign d2fef6 = hbusreq3 & d2feed | !hbusreq3 & d2fef5;
assign a656be = hgrant5_p & v845542 | !hgrant5_p & a656bd;
assign v12152f9 = hgrant2_p & v12152ed | !hgrant2_p & !v12152f8;
assign v114a233 = hgrant2_p & v845542 | !hgrant2_p & !v114a232;
assign v10d42a9 = hbusreq2_p & v10d42a3 | !hbusreq2_p & v10d42a8;
assign v134d296 = hgrant2_p & v134d27b | !hgrant2_p & v134d295;
assign v1214ef6 = hbusreq5_p & v1214ef5 | !hbusreq5_p & v1216562;
assign v1445ec1 = hmaster2_p & v144639c | !hmaster2_p & v1445ec0;
assign v1445bbc = decide_p & v1445bb4 | !decide_p & v1445bbb;
assign v13891a3 = hbusreq5_p & v13891a2 | !hbusreq5_p & v845542;
assign v12aec49 = hmaster1_p & v12afe47 | !hmaster1_p & v12aec48;
assign v1216a74 = hmaster2_p & v845542 | !hmaster2_p & v1216a73;
assign v12ad5d3 = hbusreq0_p & v15157ba | !hbusreq0_p & v845542;
assign v1668d7a = hbusreq4_p & v1668d77 | !hbusreq4_p & v1668d79;
assign v121612a = hmaster2_p & v1216111 | !hmaster2_p & v845542;
assign v1445bea = hready_p & v1445bac | !hready_p & v1445be1;
assign v1446182 = hmaster0_p & v1445fea | !hmaster0_p & v144639c;
assign v1445927 = hlock5 & v1445912 | !hlock5 & v1445925;
assign v1214c91 = hbusreq0 & v1214c90 | !hbusreq0 & v845542;
assign v12ad532 = hmaster0_p & v12ad517 | !hmaster0_p & v12ad531;
assign v12ad5fd = hbusreq2 & v12ad5f0 | !hbusreq2 & v12ad5fc;
assign v1216106 = hbusreq1 & v1216105 | !hbusreq1 & v845542;
assign v10d4089 = hmaster0_p & v10d400b | !hmaster0_p & v10d400a;
assign d301bf = hbusreq5_p & d301bd | !hbusreq5_p & d301be;
assign v1445eaf = hbusreq0 & v1445ead | !hbusreq0 & v1445eae;
assign v12162b4 = hmaster0_p & v12161fb | !hmaster0_p & v12161d3;
assign v1215c51 = hbusreq2 & v1215c49 | !hbusreq2 & v1215c50;
assign v1214cd2 = hbusreq4_p & v1215379 | !hbusreq4_p & !v1214cc7;
assign v1216b0e = hmaster1_p & v1216b0d | !hmaster1_p & v1216af8;
assign v1446266 = hbusreq0 & v1446263 | !hbusreq0 & v1446265;
assign d3013a = hmaster2_p & d2fea8 | !hmaster2_p & !v84555a;
assign v1405aac = hlock0_p & v1405a87 | !hlock0_p & !v1405a91;
assign v1515623 = stateA1_p & v1553934 | !stateA1_p & !a65884;
assign v12150cf = hmaster2_p & v845542 | !hmaster2_p & v12150ce;
assign d2fb4d = hlock0_p & v845542 | !hlock0_p & v845570;
assign v121656b = hgrant4_p & v1216524 | !hgrant4_p & v121656a;
assign a658fc = hmaster1_p & a658fb | !hmaster1_p & a658e5;
assign v1216215 = hbusreq5_p & v121620c | !hbusreq5_p & !v1216214;
assign v1216aae = hmaster2_p & v1216aa9 | !hmaster2_p & v1216aad;
assign a7c7c1 = hmaster1_p & v9337f3 | !hmaster1_p & v845542;
assign v144598f = hmaster1_p & v144598e | !hmaster1_p & v14458fd;
assign d80796 = hlock0_p & d80733 | !hlock0_p & d80795;
assign v1284d51 = hgrant2_p & v1405924 | !hgrant2_p & v1284d50;
assign v1215d01 = hgrant5_p & v845542 | !hgrant5_p & v1215cd0;
assign v14462f4 = hbusreq0 & v14462ef | !hbusreq0 & v14462f3;
assign v1284caf = hmaster1_p & v1284cae | !hmaster1_p & v1284ca7;
assign v1515705 = hbusreq2 & v1515704 | !hbusreq2 & v15167ed;
assign v1214dd8 = hlock2_p & v1214dd5 | !hlock2_p & v1214dd7;
assign v121505c = hmaster0_p & v1215030 | !hmaster0_p & v121505b;
assign v1445906 = hbusreq1 & v14458df | !hbusreq1 & v14458e3;
assign v1446446 = hbusreq5_p & v1446445 | !hbusreq5_p & v144643b;
assign v138a31d = hbusreq3 & v138a319 | !hbusreq3 & !v138a31c;
assign v12ad4d9 = hbusreq0 & v12ad4d8 | !hbusreq0 & v845542;
assign v155304e = hlock1 & v1553217 | !hlock1 & v155304d;
assign v138a48e = decide_p & v138a48d | !decide_p & v138a406;
assign f2f28c = hgrant2_p & v845542 | !hgrant2_p & f2f28b;
assign d3060b = hlock5_p & v845542 | !hlock5_p & !d3060a;
assign v1515637 = hbusreq3 & v1515622 | !hbusreq3 & v1515636;
assign d2f9bd = hbusreq2 & d2f9b5 | !hbusreq2 & d2f9bc;
assign a6564e = hgrant5_p & a653d4 | !hgrant5_p & a6564d;
assign v12adbec = hgrant3_p & v12adf67 | !hgrant3_p & v12adbeb;
assign v12af987 = hbusreq5_p & v12afda2 | !hbusreq5_p & v12af986;
assign v15168b1 = hmaster2_p & v845542 | !hmaster2_p & v15168b0;
assign v12ad635 = hmaster0_p & v12ad633 | !hmaster0_p & v12ad634;
assign v1445504 = hbusreq0 & v1445503 | !hbusreq0 & v14454ed;
assign v121654f = hbusreq0 & v1216549 | !hbusreq0 & v121654e;
assign v1552fd7 = hgrant3_p & v1552fd4 | !hgrant3_p & v1552fd6;
assign v144655b = hgrant4_p & v1446398 | !hgrant4_p & v845542;
assign v16a12ed = hbusreq0 & v16a12ec | !hbusreq0 & v16a208b;
assign v12164df = hmaster2_p & v12164dc | !hmaster2_p & v12164de;
assign f2f389 = hbusreq1_p & f2f388 | !hbusreq1_p & v845542;
assign d2fb1a = hgrant2_p & d2fad1 | !hgrant2_p & d2fb19;
assign v1445499 = hbusreq2_p & v1445498 | !hbusreq2_p & v1445bba;
assign v1445886 = hmaster2_p & v144639c | !hmaster2_p & v1445885;
assign v1445da9 = hlock0 & v1445da8 | !hlock0 & v1445da6;
assign v12afe51 = hgrant5_p & v845542 | !hgrant5_p & v12afe50;
assign v15157b6 = hburst1 & a66293 | !hburst1 & v15157b5;
assign v12150ba = hbusreq3 & v12150b9 | !hbusreq3 & !v1215ba9;
assign v12166ef = hmaster0_p & v12166d5 | !hmaster0_p & v12166ee;
assign v12160cb = hbusreq2_p & v12160ca | !hbusreq2_p & v12160c9;
assign v1215c82 = hmaster2_p & v1215fff | !hmaster2_p & v1216007;
assign v138a33b = hbusreq5_p & v1668c6f | !hbusreq5_p & v845542;
assign v16695a8 = hgrant3_p & v16695a5 | !hgrant3_p & !v16695a7;
assign v12150f3 = hbusreq2_p & v12150f2 | !hbusreq2_p & v12150f1;
assign d2f977 = hmaster2_p & d2f972 | !hmaster2_p & d2f976;
assign v144607c = hmaster2_p & v144603d | !hmaster2_p & v1446048;
assign v1214d2e = hbusreq2_p & v1214d29 | !hbusreq2_p & v1214d2d;
assign v1553158 = hlock2_p & v1553156 | !hlock2_p & v1553157;
assign v12ad5ab = hlock0_p & v1668d24 | !hlock0_p & d2fbe5;
assign v1215bc0 = hlock5_p & v1215bbf | !hlock5_p & v12163a1;
assign v1445a32 = hmaster0_p & v1445a08 | !hmaster0_p & v1445a31;
assign v12acfea = hmaster1_p & v12acfc4 | !hmaster1_p & v12acfdb;
assign v16a267a = hmaster1_p & v16a2679 | !hmaster1_p & !v16a2672;
assign v1214f10 = hmaster1_p & v1214f04 | !hmaster1_p & v1214f0f;
assign v16a1e59 = hgrant3_p & v16a1e05 | !hgrant3_p & v16a1e58;
assign v16a1ac0 = hmaster0_p & v16a1abd | !hmaster0_p & v16a2675;
assign v121610b = hgrant1_p & v845542 | !hgrant1_p & v121610a;
assign f2f32b = hbusreq2 & f2f2f1 | !hbusreq2 & f2f32a;
assign v10d4083 = hgrant5_p & v10d3feb | !hgrant5_p & v10d4082;
assign v1214c7c = hmaster0_p & v1214c56 | !hmaster0_p & v1214c7b;
assign v12ad31c = hbusreq1_p & v12ae1f0 | !hbusreq1_p & v12ad31b;
assign v15157b8 = hmastlock_p & v15157b7 | !hmastlock_p & v845542;
assign v1445efb = hlock2 & v1445ef6 | !hlock2 & v1445efa;
assign v16a13cf = hlock2_p & v16a13cd | !hlock2_p & !v16a13ce;
assign f2f420 = hgrant5_p & f2f3a1 | !hgrant5_p & !f2f41f;
assign d2fb5a = hbusreq0 & d2fb59 | !hbusreq0 & v845542;
assign d30714 = stateG2_p & v845542 | !stateG2_p & v156645f;
assign v121544a = hlock2_p & v1215449 | !hlock2_p & v1215445;
assign f2f3ec = hmaster1_p & f2f3eb | !hmaster1_p & ae2496;
assign v15533b0 = hgrant1_p & v845542 | !hgrant1_p & v15533af;
assign v12aeb18 = hmaster2_p & v845542 | !hmaster2_p & v12afda6;
assign v14463b4 = hbusreq0_p & v14463b1 | !hbusreq0_p & !v144639c;
assign a65b3b = hready_p & a65b3a | !hready_p & a65b30;
assign a65886 = hburst1 & a66293 | !hburst1 & a65885;
assign c50efd = hready_p & v845550 | !hready_p & c50efc;
assign v1445a7d = stateG10_5_p & v14459ff | !stateG10_5_p & v1445a7c;
assign v14458cf = hlock5 & v14458b7 | !hlock5 & v14458ce;
assign v1445e9e = hgrant1_p & v1445e04 | !hgrant1_p & v1445e9d;
assign v15155ed = hbusreq2_p & v15155ec | !hbusreq2_p & v845542;
assign v144540b = decide_p & v144540a | !decide_p & v1446564;
assign v1215712 = hlock0_p & v12160f2 | !hlock0_p & !v845542;
assign v12167ac = decide_p & v1216583 | !decide_p & v12167ab;
assign v1405aa0 = busreq_p & v845542 | !busreq_p & v845582;
assign v16a1391 = hmaster1_p & v16a1386 | !hmaster1_p & v16a1f96;
assign d306cb = hbusreq1_p & d306ca | !hbusreq1_p & v845542;
assign v12160e3 = hmaster0_p & v12160d4 | !hmaster0_p & v12160e2;
assign v121658e = stateA1_p & v121658d | !stateA1_p & v1216a89;
assign v1284ce5 = hmaster0_p & v1284cc9 | !hmaster0_p & v1284ce3;
assign v14466cf = hbusreq2_p & v14466cd | !hbusreq2_p & v14466ce;
assign v16695ba = hbusreq3 & v16695b2 | !hbusreq3 & v16695b9;
assign v14058f3 = hgrant4_p & v14058f1 | !hgrant4_p & v14058f2;
assign v1445903 = hmaster0_p & v14458d3 | !hmaster0_p & v1445902;
assign v1215d27 = hmaster0_p & v1668da6 | !hmaster0_p & v1216a8e;
assign v1214ee9 = hgrant5_p & v845547 | !hgrant5_p & v121656d;
assign v12ad4f9 = hmaster2_p & v12ad4f6 | !hmaster2_p & !v12ad4f7;
assign d306b9 = hbusreq2_p & d3066f | !hbusreq2_p & d306b8;
assign v121670e = hbusreq2_p & v121670a | !hbusreq2_p & v121670d;
assign v1445434 = hmaster1_p & v1445414 | !hmaster1_p & v1445b8d;
assign f2f2cc = hmaster2_p & f2f2c9 | !hmaster2_p & f2f2cb;
assign v16a1d5e = hgrant5_p & v845542 | !hgrant5_p & !v16a1d40;
assign v134d51c = hgrant2_p & v134d51b | !hgrant2_p & v134d514;
assign v1445ece = hmaster1_p & v1445ecd | !hmaster1_p & v1445eaa;
assign v134d4ab = hbusreq5_p & v134d376 | !hbusreq5_p & v134d4aa;
assign v1214dc1 = hmaster1_p & v1214d2a | !hmaster1_p & !v1214d1e;
assign v12ad676 = hlock0_p & a658c6 | !hlock0_p & v845542;
assign a6586d = hmaster2_p & v845542 | !hmaster2_p & a6586c;
assign v14460d8 = hlock2 & v14460d4 | !hlock2 & v14460d7;
assign v14457fe = hbusreq2_p & v14457dc | !hbusreq2_p & v14457fd;
assign v12157b1 = hgrant1_p & v121570e | !hgrant1_p & v12157b0;
assign v1215d43 = hmaster1_p & v1215d42 | !hmaster1_p & v1215d3a;
assign v1668e0a = hready_p & v1668c5b | !hready_p & !v1668e09;
assign v121609b = hmaster1_p & v121609a | !hmaster1_p & v1216097;
assign d2f99f = hbusreq5_p & d2f98f | !hbusreq5_p & d2f99e;
assign v151577e = hgrant0_p & v151577d | !hgrant0_p & v1515614;
assign v1515675 = hmastlock_p & v1515674 | !hmastlock_p & v845542;
assign v1516853 = decide_p & v15167ef | !decide_p & !v845576;
assign v16a2080 = hgrant1_p & v84554d | !hgrant1_p & v16a207f;
assign d30899 = hbusreq5_p & d307ab | !hbusreq5_p & d30898;
assign v12ad4ee = hmaster1_p & v12ad4ea | !hmaster1_p & v12ad4ed;
assign v1216567 = hmastlock_p & v15168f0 | !hmastlock_p & v845542;
assign d3072f = hmaster0_p & d3071e | !hmaster0_p & d3072e;
assign v1445b0d = hbusreq3 & v1445b00 | !hbusreq3 & v1445b0c;
assign v14058cb = hmaster2_p & v1405844 | !hmaster2_p & v14058c7;
assign v1215317 = hgrant2_p & v1215314 | !hgrant2_p & v1215316;
assign a65466 = stateA1_p & v1566987 | !stateA1_p & !v110b6cc;
assign v1405a8c = hbusreq1_p & v845542 | !hbusreq1_p & !v1405a87;
assign v1214ff9 = hgrant5_p & v1214fee | !hgrant5_p & v1214ff8;
assign d30720 = hlock5_p & d3071f | !hlock5_p & v84554e;
assign v16a2066 = decide_p & v16a1f9e | !decide_p & v16a2065;
assign v1515765 = hbusreq4_p & v1515763 | !hbusreq4_p & !v1515764;
assign v1214dbb = hgrant2_p & v1214db2 | !hgrant2_p & v1214db6;
assign v151562e = hburst0 & a66293 | !hburst0 & v151562d;
assign v1515609 = locked_p & v845542 | !locked_p & v10d3fd4;
assign v1445be7 = decide_p & v1446224 | !decide_p & v1445be6;
assign v1215be5 = hmaster0_p & v121601c | !hmaster0_p & v1215be4;
assign d2fc25 = hbusreq5_p & v84554a | !hbusreq5_p & d2fc24;
assign v1515659 = hmaster2_p & a658b5 | !hmaster2_p & v1515658;
assign v14058eb = hmaster2_p & v14058ea | !hmaster2_p & !v14465b3;
assign v1445e64 = hbusreq4_p & v14465ca | !hbusreq4_p & v14465d6;
assign v15160fa = hmaster1_p & v15160f9 | !hmaster1_p & v845542;
assign f2f374 = hgrant1_p & v845570 | !hgrant1_p & !f2f373;
assign v12ae1fb = hgrant1_p & v845542 | !hgrant1_p & v12ae1fa;
assign f2f402 = hbusreq2 & f2f3fd | !hbusreq2 & f2f401;
assign v1446612 = hbusreq5_p & v1446605 | !hbusreq5_p & v1446611;
assign v1216270 = hmaster1_p & v121626f | !hmaster1_p & !v1216027;
assign v1284d36 = hlock2_p & v1284d33 | !hlock2_p & v1284d35;
assign v16a1399 = decide_p & v16a1398 | !decide_p & v16a2065;
assign v1446274 = hmaster1_p & v1446273 | !hmaster1_p & v1446271;
assign v10d4055 = hmaster2_p & v10d401e | !hmaster2_p & v10d403a;
assign v14058f7 = hgrant5_p & v14058ed | !hgrant5_p & !v14058f6;
assign d2fe86 = hmaster2_p & d2fe80 | !hmaster2_p & d2fe85;
assign v1214d33 = hready_p & v1214ce5 | !hready_p & v1214d32;
assign v1214dd2 = hbusreq2_p & v1214dd1 | !hbusreq2_p & v845542;
assign v121618c = hgrant5_p & v845542 | !hgrant5_p & v1216101;
assign v15157ca = hgrant4_p & a662a9 | !hgrant4_p & v15157c9;
assign f2f3ef = hmaster0_p & f2f2dd | !hmaster0_p & f2f2cc;
assign v1668c89 = hmaster2_p & a658ad | !hmaster2_p & !a658ca;
assign v1445ed3 = hmaster0_p & v1445e84 | !hmaster0_p & v1445e95;
assign v12ad02c = hbusreq0 & v12ad02b | !hbusreq0 & v12afa0a;
assign a6568e = hmaster1_p & a65493 | !hmaster1_p & a658e5;
assign v1284cf8 = hgrant0_p & v1284cf7 | !hgrant0_p & !v140584b;
assign v134d4ee = hgrant5_p & v134d4ed | !hgrant5_p & v134d4eb;
assign v12153ad = hmaster1_p & v12153ac | !hmaster1_p & v12153a9;
assign v14058ee = hgrant1_p & v140583f | !hgrant1_p & !v14465b2;
assign f2e4e1 = hgrant3_p & f2e4cd | !hgrant3_p & f2e4e0;
assign d305e5 = hbusreq5 & d305e4 | !hbusreq5 & v845542;
assign v1445b20 = hmaster1_p & v1445b03 | !hmaster1_p & v144591b;
assign v121621c = hmaster2_p & v1216218 | !hmaster2_p & v121621b;
assign v16a13fb = hbusreq2_p & v16a13fa | !hbusreq2_p & v16a209d;
assign v10d4289 = hgrant0_p & v10d3fdb | !hgrant0_p & !v10d4288;
assign v1215ca5 = hgrant1_p & v1215ca3 | !hgrant1_p & v1215ca4;
assign a65b23 = hgrant3_p & a65b07 | !hgrant3_p & a65b21;
assign v12ad4bf = hbusreq1_p & v12adf61 | !hbusreq1_p & v12ad4be;
assign v1214c3d = hmaster0_p & v1214c2c | !hmaster0_p & v1214c3c;
assign v134d222 = hmaster0_p & v134d221 | !hmaster0_p & v134d1e8;
assign v16a2239 = hmastlock_p & v16a2238 | !hmastlock_p & !v845542;
assign a65479 = hmaster1_p & a658e8 | !hmaster1_p & a65476;
assign v1216163 = hbusreq1 & v1216162 | !hbusreq1 & v845542;
assign v138937f = hmaster1_p & v1389de1 | !hmaster1_p & v138937e;
assign d2fb38 = hbusreq1_p & d2fec3 | !hbusreq1_p & d2fb37;
assign v1553432 = hbusreq2 & v1553430 | !hbusreq2 & v1553431;
assign v1405b55 = hmaster1_p & v1405b42 | !hmaster1_p & v1405b09;
assign v1215707 = hmaster0_p & v1215b7e | !hmaster0_p & v1215b7c;
assign v1445e1d = hmaster0_p & v1445de6 | !hmaster0_p & v1445e0a;
assign a653d7 = hburst1 & v845542 | !hburst1 & !v88d3e4;
assign d300c9 = hbusreq5_p & d300c8 | !hbusreq5_p & !d300c7;
assign v12ad5c3 = hbusreq1_p & v12ad5af | !hbusreq1_p & v12ad5c2;
assign v134d238 = hlock3 & v134d227 | !hlock3 & v134d237;
assign d2fbee = hmaster2_p & d2fbed | !hmaster2_p & d2fbe0;
assign v138a396 = hmaster1_p & v138a395 | !hmaster1_p & v138a341;
assign v12ad4f0 = hlock0_p & v10d3fd4 | !hlock0_p & !v845542;
assign v144608e = hgrant1_p & v1445fe7 | !hgrant1_p & v144608d;
assign v12167a1 = hmaster0_p & v1668c1f | !hmaster0_p & v1216a8f;
assign d2fc2c = hlock0_p & v845542 | !hlock0_p & !d2fc2b;
assign v12ad4db = hmaster2_p & v12ad4da | !hmaster2_p & v845542;
assign v1389e25 = hgrant5_p & v1668c3f | !hgrant5_p & !v845542;
assign v1216179 = hmaster2_p & v121610b | !hmaster2_p & v1216131;
assign v12ad67e = hbusreq1 & v12ad677 | !hbusreq1 & v12ad67d;
assign v12ad60e = hlock5_p & v12ad60b | !hlock5_p & v12ad60d;
assign v15156da = hmaster0_p & v15156d9 | !hmaster0_p & !v151566a;
assign d305f1 = hbusreq4_p & d305ef | !hbusreq4_p & d305f0;
assign d30771 = hmaster1_p & d30767 | !hmaster1_p & d30754;
assign v16a1ce0 = hbusreq2 & v16a1cdd | !hbusreq2 & v16a1cdf;
assign v1214ddb = hbusreq3 & v1214dd3 | !hbusreq3 & v1214dda;
assign d2fc5b = hbusreq4_p & d2fbeb | !hbusreq4_p & d2fc52;
assign v121628b = hgrant2_p & v1216289 | !hgrant2_p & !v121628a;
assign v1215c27 = hbusreq1 & v1216024 | !hbusreq1 & v845542;
assign v12160a6 = hmaster0_p & v121605f | !hmaster0_p & v1216068;
assign v14462e6 = hmaster2_p & v14465ae | !hmaster2_p & v1446403;
assign d306e5 = hmaster1_p & d306d2 | !hmaster1_p & d306e4;
assign v1214bc4 = hmaster0_p & v12153b1 | !hmaster0_p & v1214bb7;
assign v134d521 = hmaster0_p & v845542 | !hmaster0_p & v134d517;
assign v1445b11 = hmaster1_p & v1445aea | !hmaster1_p & v144591b;
assign v1405880 = hmaster1_p & v140587f | !hmaster1_p & !v1446403;
assign v1553427 = decide_p & v845542 | !decide_p & v155313b;
assign v1214cf2 = hbusreq1_p & v1214c2a | !hbusreq1_p & !v1214cf1;
assign v1284d00 = hmaster2_p & v140583c | !hmaster2_p & !v1284ce9;
assign v151584f = hbusreq5 & v1515841 | !hbusreq5 & v151584e;
assign v14464a6 = hbusreq5_p & v14464a4 | !hbusreq5_p & v14464a5;
assign v1405848 = hbusreq5_p & v1405846 | !hbusreq5_p & v1405847;
assign v138a3c6 = hlock5_p & v138a3c5 | !hlock5_p & !v1515796;
assign v12acfe3 = hbusreq2 & v12acfdd | !hbusreq2 & v12acfe2;
assign v10d4066 = hgrant0_p & v10d3fe0 | !hgrant0_p & v10d3fdf;
assign v1215baa = hbusreq3 & v1215ba6 | !hbusreq3 & !v1215ba9;
assign v1668de8 = decide_p & v1668de7 | !decide_p & v845542;
assign d2fae2 = hgrant1_p & d2fade | !hgrant1_p & d2fae1;
assign d307c8 = hbusreq4_p & v845542 | !hbusreq4_p & d307b2;
assign bf1f6e = hbusreq5_p & bf1f6d | !hbusreq5_p & !bf1f6c;
assign v12ad010 = hgrant4_p & v12ad5d8 | !hgrant4_p & !v12ad00f;
assign d306e0 = hbusreq1 & d306df | !hbusreq1 & v845542;
assign v1405b66 = hbusreq3_p & v1405b34 | !hbusreq3_p & v1405b65;
assign d3065b = hgrant0_p & d3065a | !hgrant0_p & v845570;
assign v155309f = hlock2 & v155341e | !hlock2 & v155309b;
assign v144626c = hbusreq0 & v1446445 | !hbusreq0 & v144643d;
assign v1215fe3 = hbusreq5 & v1215fc1 | !hbusreq5 & v1215fe2;
assign d307ed = hgrant1_p & v845542 | !hgrant1_p & d307ec;
assign f2f436 = hmaster2_p & f2f434 | !hmaster2_p & f2f435;
assign v16a13ee = hgrant5_p & v845542 | !hgrant5_p & !v16a13dc;
assign f2e4c9 = hbusreq3_p & f2e884 | !hbusreq3_p & f2e4c8;
assign v1446174 = hmaster0_p & v144607f | !hmaster0_p & v144603f;
assign v1445bc4 = hmaster1_p & v1446466 | !hmaster1_p & v1445bc3;
assign v12162db = hgrant2_p & v12162c3 | !hgrant2_p & v12162da;
assign d3091a = hmaster1_p & d3090c | !hmaster1_p & d30918;
assign v16a142b = hready_p & v845555 | !hready_p & v16a142a;
assign d301dc = hbusreq5_p & d301db | !hbusreq5_p & !d301da;
assign v1515718 = stateA1_p & v845542 | !stateA1_p & !v1515717;
assign v1445b7c = hgrant2_p & v144634f | !hgrant2_p & v1445b7b;
assign v1214efc = hlock2_p & v1214eed | !hlock2_p & v1214efb;
assign f2f3e8 = hmaster0_p & f2f396 | !hmaster0_p & f2f3a1;
assign v12ad51f = hbusreq5_p & v12ad51d | !hbusreq5_p & !v12ad51e;
assign v1405897 = hmaster2_p & v140583f | !hmaster2_p & v1405845;
assign v134ce56 = hmaster1_p & v134ce55 | !hmaster1_p & v845542;
assign v16a19d2 = hmaster2_p & v16a19d1 | !hmaster2_p & v845542;
assign v1668d47 = hbusreq4 & a65862 | !hbusreq4 & v845570;
assign f2e4e8 = decide_p & f2e4e7 | !decide_p & v845542;
assign v1445dca = hbusreq3 & v1445dc8 | !hbusreq3 & v1445dc9;
assign v16a12f6 = hgrant2_p & v845542 | !hgrant2_p & v16a12f4;
assign d30846 = hready_p & d30845 | !hready_p & d3077b;
assign v1552f6a = hmaster1_p & v1553385 | !hmaster1_p & v1552f69;
assign v1216231 = hbusreq1_p & v1216230 | !hbusreq1_p & !v845542;
assign v15157e8 = hgrant5_p & v15157e7 | !hgrant5_p & !v151574a;
assign d306e7 = hmaster0_p & d306ce | !hmaster0_p & d306e6;
assign a65648 = hbusreq5_p & a653d3 | !hbusreq5_p & a65647;
assign v16695b2 = hbusreq2_p & v166959f | !hbusreq2_p & v1668e06;
assign v12ad0bb = hmaster1_p & v845542 | !hmaster1_p & v12ad0ba;
assign v12af7f4 = hbusreq4_p & v845542 | !hbusreq4_p & v1405a7d;
assign v16a1e4a = hbusreq3 & v16a1e2b | !hbusreq3 & v16a1e49;
assign v14459bf = hbusreq0_p & v14459be | !hbusreq0_p & v144639e;
assign v16a1e6c = hbusreq2_p & v16a1dc1 | !hbusreq2_p & v16a1e6b;
assign v1405916 = hbusreq5_p & v1405871 | !hbusreq5_p & v1405915;
assign v14459a7 = locked_p & v144639c | !locked_p & !v14459a6;
assign d2f980 = hbusreq5_p & v84555a | !hbusreq5_p & d3068e;
assign v12aead5 = hgrant3_p & v12af1c4 | !hgrant3_p & v12aead4;
assign f2f3c4 = hgrant5_p & f2f3bf | !hgrant5_p & !f2f370;
assign v1445e2c = hmaster1_p & v1445e17 | !hmaster1_p & v1445e28;
assign v1445e04 = hbusreq1 & v1445e02 | !hbusreq1 & v1445e03;
assign v16693b2 = hready_p & v16693a5 | !hready_p & !v16693b1;
assign f2f220 = hmaster2_p & v845542 | !hmaster2_p & !f2f21f;
assign v14458a1 = hmaster2_p & v144639c | !hmaster2_p & v1445871;
assign d302e1 = hgrant5_p & v845542 | !hgrant5_p & d30663;
assign v1445eb5 = hgrant5_p & v1445eb3 | !hgrant5_p & v1445eb4;
assign v1216a9c = hmaster1_p & v1216a92 | !hmaster1_p & v1216a9b;
assign v1446068 = hbusreq1 & v144661d | !hbusreq1 & v1446628;
assign v1215344 = hbusreq3_p & v12150b4 | !hbusreq3_p & !v1215343;
assign v10d40af = hready_p & v10d40a4 | !hready_p & v10d40ae;
assign v1445fc9 = hlock5 & v1445fb2 | !hlock5 & v1445fc7;
assign v1216011 = hbusreq2_p & v121600d | !hbusreq2_p & v1216010;
assign v1214db3 = hgrant2_p & v1214db2 | !hgrant2_p & v1214daa;
assign d2fd40 = hbusreq2 & d2fd3f | !hbusreq2 & d2fd3d;
assign v155321c = hready_p & v155313d | !hready_p & v155321b;
assign v14457ee = hmaster1_p & v14457ed | !hmaster1_p & v1445e1b;
assign v1445edb = hbusreq2_p & v1445ed5 | !hbusreq2_p & v1445eda;
assign v138a346 = hmaster1_p & v138a345 | !hmaster1_p & v138a341;
assign d2fce7 = hgrant1_p & d2fce6 | !hgrant1_p & d305ef;
assign v1215c04 = hbusreq5_p & v1215c02 | !hbusreq5_p & !v1215c03;
assign v1216aa6 = stateG2_p & v845542 | !stateG2_p & v1216aa5;
assign v1515791 = hgrant0_p & a6537d | !hgrant0_p & !v1515790;
assign v1668dc6 = hbusreq5_p & v1668dc3 | !hbusreq5_p & !v1668dc5;
assign a65451 = hbusreq2_p & a6544c | !hbusreq2_p & !a65450;
assign a662b2 = hbusreq5_p & a66290 | !hbusreq5_p & a662ad;
assign v144673c = hmaster1_p & v144673b | !hmaster1_p & v144644d;
assign v1553444 = decide_p & v1553443 | !decide_p & v15532cd;
assign v12166fd = hbusreq5_p & v12166fc | !hbusreq5_p & v16a2243;
assign v1445b72 = hbusreq2 & v1445b6d | !hbusreq2 & v1445b71;
assign v12164e2 = hmaster1_p & v12164d8 | !hmaster1_p & v12164e1;
assign d306bb = hbusreq2 & d306b9 | !hbusreq2 & d306ba;
assign v1446080 = hbusreq0 & v144607d | !hbusreq0 & v144607f;
assign v12166e7 = hlock0_p & v12166e5 | !hlock0_p & v12166e6;
assign v15534da = hlock0 & v15534d3 | !hlock0 & v15534d9;
assign v1515ae0 = hmaster1_p & v1515adf | !hmaster1_p & v845570;
assign v1445b05 = hbusreq2_p & v1445b02 | !hbusreq2_p & v1445b04;
assign v15156d8 = hmaster2_p & a658ca | !hmaster2_p & !v1515658;
assign v84554d = hbusreq1 & v845542 | !hbusreq1 & !v845542;
assign v1445826 = hgrant2_p & v1445824 | !hgrant2_p & v1445825;
assign v1445814 = hmaster0_p & v1445802 | !hmaster0_p & v1445edf;
assign v1668ccc = hburst1 & a66272 | !hburst1 & v1668ccb;
assign v1215d2a = hbusreq5_p & v1215d28 | !hbusreq5_p & v1215d29;
assign bf1f7f = hgrant4_p & v84556a | !hgrant4_p & !bf1f77;
assign d3024e = hgrant5_p & v845542 | !hgrant5_p & d30212;
assign v12162ea = hmaster0_p & v12162e8 | !hmaster0_p & v12162e9;
assign v12afda3 = hlock0_p & v84556a | !hlock0_p & !v845542;
assign a6565f = hbusreq2 & a65656 | !hbusreq2 & a6565c;
assign v16a1e53 = hgrant2_p & v16a1e00 | !hgrant2_p & v16a1e52;
assign v144661b = hlock0_p & v14463b1 | !hlock0_p & v14463b2;
assign v144579e = hmaster0_p & v144579d | !hmaster0_p & v1445de7;
assign d307e5 = hgrant1_p & v845542 | !hgrant1_p & d307e4;
assign v1668c68 = stateA1_p & a66272 | !stateA1_p & ab83a0;
assign v1389f83 = hmaster2_p & a66275 | !hmaster2_p & !v845542;
assign v14466a7 = hbusreq5_p & v14466a6 | !hbusreq5_p & v1446611;
assign v1445421 = hmaster1_p & v1445414 | !hmaster1_p & v1446341;
assign v15157ba = hbusreq4 & v151561c | !hbusreq4 & v15157b9;
assign v1215ff7 = locked_p & v845542 | !locked_p & v1215ff6;
assign a65896 = hbusreq3 & a6587b | !hbusreq3 & a65894;
assign v16a1421 = hbusreq2_p & v16a13c9 | !hbusreq2_p & !v16a1da9;
assign a65460 = hmaster0_p & a6540c | !hmaster0_p & v845558;
assign f2f3e9 = hmaster1_p & f2f3e8 | !hmaster1_p & f2f39d;
assign v12aeb19 = hbusreq0 & v12afda2 | !hbusreq0 & v12aeb18;
assign a6629f = hgrant2_p & v845542 | !hgrant2_p & a6629e;
assign v155341f = hlock2 & v155341e | !hlock2 & v15533b8;
assign d30295 = hgrant2_p & d30267 | !hgrant2_p & d30294;
assign v1445419 = hmaster0_p & v14465b7 | !hmaster0_p & v1446643;
assign v1553384 = hmaster2_p & v1553383 | !hmaster2_p & v845542;
assign v1215454 = hbusreq2 & v1215450 | !hbusreq2 & v1215453;
assign v1214bfb = hmaster1_p & v12153ab | !hmaster1_p & v12153a9;
assign v16a1db0 = hbusreq5_p & v16a207a | !hbusreq5_p & v16a1add;
assign d30620 = hlock2_p & d3061d | !hlock2_p & d3061f;
assign v144627c = hbusreq0 & v1446426 | !hbusreq0 & v144642c;
assign v16a13d4 = hlock2_p & v16a13d2 | !hlock2_p & !v16a13d3;
assign v15533a1 = hgrant4_p & v845542 | !hgrant4_p & v15533a0;
assign v121507c = hmaster1_p & v1215030 | !hmaster1_p & !v121507b;
assign v121574b = hgrant1_p & v1215736 | !hgrant1_p & v845542;
assign v15157d0 = hbusreq0 & v15157c5 | !hbusreq0 & v15157cf;
assign v151564d = hmastlock_p & v151564c | !hmastlock_p & v10d3fd3;
assign v1446682 = hgrant2_p & v1446681 | !hgrant2_p & v1446665;
assign v1215c55 = hgrant5_p & v845542 | !hgrant5_p & v1215bf7;
assign f2e882 = decide_p & f2ec25 | !decide_p & f2f23c;
assign v1668cac = hmaster1_p & v1668c8a | !hmaster1_p & !v1668c9c;
assign f2f34b = hbusreq1_p & f2f34a | !hbusreq1_p & v845542;
assign v1446623 = hbusreq5_p & v1446622 | !hbusreq5_p & v1446611;
assign v1214dcc = hmaster2_p & v1216a5a | !hmaster2_p & v845542;
assign v1553501 = hgrant2_p & v15534f1 | !hgrant2_p & v15534ff;
assign v12acfcc = hmaster1_p & v12acfcb | !hmaster1_p & !v12acfb9;
assign d308c4 = hgrant5_p & d30654 | !hgrant5_p & d308a9;
assign v1216578 = hgrant2_p & v845547 | !hgrant2_p & v1216576;
assign v16a1aef = hbusreq5 & v16a1ae5 | !hbusreq5 & v16a1aee;
assign v11e594f = hgrant5_p & bf1f62 | !hgrant5_p & !v11e594d;
assign d2f982 = hbusreq5_p & v84555a | !hbusreq5_p & !d2f981;
assign d2fd47 = hbusreq2 & d2fd46 | !hbusreq2 & d302ec;
assign v134d365 = hgrant0_p & v845542 | !hgrant0_p & v134d273;
assign bf1f86 = hmaster1_p & bf1f7b | !hmaster1_p & bf1f85;
assign v144625e = hlock5 & v1446246 | !hlock5 & v144625d;
assign v1515802 = hmaster1_p & v15157a5 | !hmaster1_p & v1515801;
assign d308d5 = decide_p & v845556 | !decide_p & v845570;
assign v14459ae = hlock4 & v144639c | !hlock4 & v14459ad;
assign v12ad582 = hmaster1_p & v12ad569 | !hmaster1_p & v12ad54f;
assign v12ae1f7 = hgrant0_p & v12ae1f6 | !hgrant0_p & v845542;
assign v1446417 = hbusreq5_p & v1446416 | !hbusreq5_p & v1446413;
assign v14453e7 = hbusreq2 & v14453e3 | !hbusreq2 & v14453e6;
assign v1446162 = hmaster1_p & v1446161 | !hmaster1_p & v1445fde;
assign v8b6f6c = jx2_p & v845542 | !jx2_p & !v845542;
assign v1215733 = hlock1_p & v1215732 | !hlock1_p & v1215b97;
assign d3085d = hbusreq5_p & v84554e | !hbusreq5_p & d3085c;
assign v144660d = hgrant0_p & v144660b | !hgrant0_p & !v144660c;
assign v1445ba6 = hbusreq5 & v1445b88 | !hbusreq5 & v1445ba5;
assign v1214c5a = hlock1_p & v1214c58 | !hlock1_p & v1214c59;
assign v12ad66d = busreq_p & v151566d | !busreq_p & v12ad50e;
assign d3066b = hbusreq5_p & d3066a | !hbusreq5_p & d30663;
assign v12161d0 = hgrant1_p & v845542 | !hgrant1_p & v12161cf;
assign v1445eee = hbusreq0 & v1445eed | !hbusreq0 & v1445e84;
assign v1216223 = hbusreq0 & v121621d | !hbusreq0 & v1216222;
assign v134d3e3 = hgrant2_p & v845542 | !hgrant2_p & v134d3e2;
assign v10d406a = hmaster2_p & v10d4062 | !hmaster2_p & !v10d4069;
assign v1445a78 = hgrant5_p & v1445a75 | !hgrant5_p & v1445a77;
assign a658b2 = stateA1_p & v845542 | !stateA1_p & !ab8d68;
assign v16a140f = hgrant2_p & v16a1dec | !hgrant2_p & v16a140e;
assign v1216107 = hgrant4_p & v12160f3 | !hgrant4_p & v845572;
assign v12ad663 = hmaster2_p & v845542 | !hmaster2_p & !d30690;
assign v1446290 = hmaster0_p & v144628f | !hmaster0_p & v144627d;
assign v1446280 = hbusreq0 & v144643a | !hbusreq0 & v144643d;
assign d2fb75 = hbusreq0 & d2fb74 | !hbusreq0 & v845542;
assign v14461f5 = hlock2 & v14461f1 | !hlock2 & v14461f4;
assign v1215b91 = hlock4_p & v1215b8f | !hlock4_p & v1215b90;
assign d2fd01 = hbusreq2_p & d2fd00 | !hbusreq2_p & d302d6;
assign v1215374 = hlock3_p & v1215363 | !hlock3_p & v1215373;
assign v12150c1 = hready & v845542 | !hready & !f2f4ad;
assign v16a1aec = hgrant2_p & v845542 | !hgrant2_p & v16a1ae9;
assign d30744 = hmaster2_p & d3071b | !hmaster2_p & d30743;
assign v1668d71 = hgrant4_p & v1668d70 | !hgrant4_p & v1668d1c;
assign v1215738 = hbusreq4 & v1215ff6 | !hbusreq4 & v845542;
assign v138a3de = hbusreq5_p & v138a3dd | !hbusreq5_p & !v845542;
assign d2fc10 = hbusreq0 & d2fc0f | !hbusreq0 & d302e0;
assign v1445a86 = hmaster1_p & v1445a44 | !hmaster1_p & v1445a82;
assign a65add = decide_p & a662c3 | !decide_p & a662a2;
assign v1553151 = hmaster0_p & v1553140 | !hmaster0_p & v1553150;
assign v14465e0 = hbusreq1_p & v14465b2 | !hbusreq1_p & v14465ce;
assign d2fb84 = hmaster2_p & d2fb69 | !hmaster2_p & d2fb83;
assign v1445ab7 = hbusreq2_p & v1445ab1 | !hbusreq2_p & v1445ab6;
assign v1216a87 = hburst0_p & v118e18f | !hburst0_p & !v845542;
assign v14460df = hlock5 & v14460a1 | !hlock5 & v14460de;
assign d30665 = hlock0_p & v1668c1c | !hlock0_p & v845542;
assign v1668ce0 = hmaster2_p & v1668cbd | !hmaster2_p & v1668cdf;
assign v16a2244 = hmaster2_p & v16a223d | !hmaster2_p & v845542;
assign v1214cbf = hmaster2_p & v1214cbc | !hmaster2_p & v1214cbe;
assign v12ad562 = hbusreq3 & v12ad558 | !hbusreq3 & v12ad561;
assign a6586e = hmaster0_p & a65869 | !hmaster0_p & a6586d;
assign v1215fee = hlock1_p & v1215feb | !hlock1_p & v1215fed;
assign v134ce38 = hgrant1_p & v134ce37 | !hgrant1_p & v845542;
assign v1668dde = hmaster0_p & v1668db9 | !hmaster0_p & v1668ddd;
assign v1445acc = hlock3 & v1445ac1 | !hlock3 & v1445acb;
assign v134d52f = hmaster1_p & v134d52e | !hmaster1_p & v845542;
assign v1216529 = hgrant0_p & v1216525 | !hgrant0_p & !v1216528;
assign v16a1ce9 = hready_p & v845555 | !hready_p & v16a1ce8;
assign v1445dde = hbusreq3 & v1445ddc | !hbusreq3 & v1445ddd;
assign v151570c = hlock3_p & v15156f0 | !hlock3_p & v151570b;
assign v1668c32 = hbusreq3 & v1668c2c | !hbusreq3 & v1668c31;
assign v1216591 = stateA1_p & d30788 | !stateA1_p & !v845542;
assign a65863 = hbusreq4_p & a65862 | !hbusreq4_p & v845542;
assign v144612f = hbusreq2_p & v1446129 | !hbusreq2_p & v144612e;
assign v16a197a = hbusreq2 & v16a1978 | !hbusreq2 & !v16a1979;
assign v155305c = hmaster2_p & v155305b | !hmaster2_p & v15533a2;
assign d30881 = hlock2_p & d3087e | !hlock2_p & !d30880;
assign v1445ac1 = hbusreq2 & v1445abb | !hbusreq2 & v1445ac0;
assign v1668e02 = hready_p & v1668de8 | !hready_p & v1668e01;
assign d30915 = hbusreq5_p & d30914 | !hbusreq5_p & !d30913;
assign v10d40c4 = hbusreq5_p & v10d4056 | !hbusreq5_p & !v10d40c3;
assign v1446127 = hbusreq2 & v1446120 | !hbusreq2 & v1446126;
assign v12afe6f = hbusreq0 & v12afe47 | !hbusreq0 & v12afe63;
assign v134d1f1 = hlock1_p & v134d1f0 | !hlock1_p & v845542;
assign d308b4 = hbusreq2 & d308b0 | !hbusreq2 & d308b3;
assign v1445f11 = hbusreq2_p & v1445f0b | !hbusreq2_p & v1445f0d;
assign v138a435 = hready_p & v138a407 | !hready_p & !v138a434;
assign v16a1d32 = hmaster1_p & v16a1d2d | !hmaster1_p & v16a1f96;
assign v144631f = hmaster2_p & v144639c | !hmaster2_p & v144665b;
assign a656ae = hbusreq2_p & a656ac | !hbusreq2_p & a656ad;
assign v134d4a9 = hmaster2_p & v134d3a9 | !hmaster2_p & v845542;
assign v1446396 = stateG2_p & v845542 | !stateG2_p & v1446395;
assign v15157e1 = hgrant5_p & v1668da6 | !hgrant5_p & v1515737;
assign d3068c = hmaster2_p & v845542 | !hmaster2_p & !d30654;
assign d306c7 = hbusreq3_p & d30683 | !hbusreq3_p & d306c6;
assign v144671b = hlock2 & v1446700 | !hlock2 & v1446719;
assign v1389390 = hmaster0_p & v138938e | !hmaster0_p & !v138938f;
assign v1214d7c = hbusreq2_p & v1214d79 | !hbusreq2_p & v1214d7b;
assign f2f3f3 = hmaster0_p & f2f2dd | !hmaster0_p & f2f2e3;
assign v15533a5 = hgrant1_p & v845542 | !hgrant1_p & v155339c;
assign d2fb0e = hbusreq5_p & d3010b | !hbusreq5_p & !d2fb0d;
assign v134d50b = hmaster2_p & v134d4ff | !hmaster2_p & v134d50a;
assign f2f390 = hgrant5_p & f2f385 | !hgrant5_p & !f2f38e;
assign v14466ca = hmaster1_p & v14466c9 | !hmaster1_p & v845542;
assign v1215c79 = hbusreq2 & v1215c75 | !hbusreq2 & v1215c78;
assign v1215ce5 = hbusreq5_p & v1215ce4 | !hbusreq5_p & v1215c8d;
assign v14058ff = hgrant5_p & v1446403 | !hgrant5_p & v14058fe;
assign v144616c = hmaster1_p & v144616b | !hmaster1_p & v1445fde;
assign v1216086 = hbusreq2_p & v1216085 | !hbusreq2_p & v1216084;
assign d2fcb6 = hmaster1_p & d2fcac | !hmaster1_p & !d2fcb5;
assign v13897f1 = hgrant2_p & v845542 | !hgrant2_p & !v13897f0;
assign v1445f21 = hmaster0_p & v1445e4d | !hmaster0_p & v845542;
assign v1214817 = hbusreq5 & v12147f1 | !hbusreq5 & v1214816;
assign f2f342 = hready_p & f2f2b1 | !hready_p & f2f341;
assign v1445f93 = hbusreq1_p & v1445f92 | !hbusreq1_p & v14463b9;
assign f2f4b0 = hmastlock_p & f2f4af | !hmastlock_p & v845542;
assign v14461d7 = hmaster1_p & v1446193 | !hmaster1_p & v1445ffc;
assign v1216a94 = hmaster2_p & v845542 | !hmaster2_p & v1216a93;
assign v1668dd4 = hgrant2_p & v1668d1f | !hgrant2_p & v1668dd3;
assign v16a19aa = hgrant1_p & v845542 | !hgrant1_p & v16a19a9;
assign v84556e = decide_p & v845542 | !decide_p & !v845542;
assign v1215ddf = jx1_p & v12162e4 | !jx1_p & v1215dde;
assign d30797 = hmaster2_p & d30793 | !hmaster2_p & d30796;
assign v144609a = hmaster1_p & v144603f | !hmaster1_p & v1446099;
assign v12ad032 = hgrant2_p & v12ad01d | !hgrant2_p & !v12ad02e;
assign v12164ca = hbusreq2 & v12164c5 | !hbusreq2 & v12164c9;
assign v16a143b = hbusreq0 & v16a143a | !hbusreq0 & v16a208b;
assign v16a1ae2 = hbusreq2_p & v16a2097 | !hbusreq2_p & v16a1ae1;
assign v16a1419 = hbusreq2 & v16a1418 | !hbusreq2 & v16a1f9b;
assign v1668cbd = hmastlock_p & v1668cbc | !hmastlock_p & !v845542;
assign d30190 = hlock2_p & d3018f | !hlock2_p & d3091a;
assign v12ad62e = decide_p & v12ad593 | !decide_p & !v12afe76;
assign v15161cd = hlock2_p & v15161cc | !hlock2_p & !v845542;
assign d30696 = hmaster1_p & d3068b | !hmaster1_p & d30695;
assign v1446450 = hmaster1_p & v144644f | !hmaster1_p & v144644d;
assign v1214bf9 = hmaster0_p & v12153ab | !hmaster0_p & v1215396;
assign v1215bd9 = hready_p & v845542 | !hready_p & v1215bd8;
assign v1405874 = hlock2_p & v1405870 | !hlock2_p & v1405873;
assign v1446704 = hmaster1_p & v1446703 | !hmaster1_p & v1446436;
assign v1445df1 = hlock1 & v1445dec | !hlock1 & v1445de9;
assign v134d3b6 = hlock2 & v134d3b5 | !hlock2 & v134d39c;
assign v134ce71 = hgrant3_p & v134d3fc | !hgrant3_p & v134ce70;
assign v1214d59 = hbusreq2_p & v1214c0e | !hbusreq2_p & v1214d58;
assign v12adf60 = hlock4_p & v12adf5f | !hlock4_p & d30727;
assign v15534cf = hbusreq1_p & v15534ce | !hbusreq1_p & v155339c;
assign v15157c3 = hgrant5_p & v845570 | !hgrant5_p & v15157c2;
assign v1445ffe = hmaster1_p & v1445fe4 | !hmaster1_p & v1445ffc;
assign a6545b = hmaster0_p & a653ea | !hmaster0_p & a653f9;
assign v1215c7d = hmaster0_p & v1668da6 | !hmaster0_p & v1215c7c;
assign v1446076 = hmaster2_p & v144639c | !hmaster2_p & v1446043;
assign v151560c = hmaster0_p & v151560a | !hmaster0_p & v151560b;
assign v12acfd7 = hmaster1_p & v12ad66b | !hmaster1_p & v12ad54f;
assign v16a1448 = hgrant3_p & v16a1436 | !hgrant3_p & v16a1447;
assign v1445804 = hmaster1_p & v1445803 | !hmaster1_p & v1445e07;
assign v12ad5c5 = hmaster2_p & v12ad5b0 | !hmaster2_p & v12ad5c4;
assign v16a1bf3 = hmaster2_p & v16a1bf0 | !hmaster2_p & v16a208a;
assign v155313e = stateG3_2_p & v845542 | !stateG3_2_p & !v845586;
assign v1215c1f = hgrant1_p & v1215c14 | !hgrant1_p & v121612e;
assign v138a3aa = hmaster0_p & v138a34f | !hmaster0_p & v138a354;
assign v12af22b = hbusreq2_p & v12af5b0 | !hbusreq2_p & v12af22a;
assign v12147e6 = hmaster1_p & v12147e5 | !hmaster1_p & v1215d3a;
assign v144613b = hbusreq2_p & v1446135 | !hbusreq2_p & v144613a;
assign v12ad545 = hmaster1_p & v12ad544 | !hmaster1_p & !v12ad525;
assign v10d3fee = hbusreq2_p & v10d3fea | !hbusreq2_p & v10d3fed;
assign v1445a93 = hlock3 & v1445a69 | !hlock3 & v1445a92;
assign v1405a86 = hmastlock_p & v1405a85 | !hmastlock_p & !v845542;
assign v14453aa = hmaster1_p & v1445b40 | !hmaster1_p & v1445a9b;
assign v1284c93 = hmaster0_p & v1284c90 | !hmaster0_p & v1405859;
assign v1445d9d = hmaster2_p & v14463b9 | !hmaster2_p & v1445d99;
assign v1445f1b = hbusreq3 & v1445f19 | !hbusreq3 & v1445f1a;
assign v151571b = hmastlock_p & v151571a | !hmastlock_p & v845542;
assign v1446688 = hmaster2_p & v144639c | !hmaster2_p & v1446410;
assign v1668c8a = hmaster0_p & v1668c5f | !hmaster0_p & v1668c89;
assign v14838bc = hgrant2_p & v845558 | !hgrant2_p & v14838bb;
assign v121578c = hgrant5_p & v845542 | !hgrant5_p & v1215722;
assign v16a1c99 = hgrant1_p & v16a1c96 | !hgrant1_p & v16a1c98;
assign v12acfc7 = hbusreq2_p & v12acfc0 | !hbusreq2_p & v12acfc6;
assign v16a1d2f = hbusreq2 & v16a1d2c | !hbusreq2 & v16a1d2e;
assign v1446734 = hbusreq2_p & v1446729 | !hbusreq2_p & v1446733;
assign v10d426c = hmaster2_p & v10d426b | !hmaster2_p & v10d4024;
assign d8074d = hmaster0_p & d80748 | !hmaster0_p & d8073b;
assign f2f29e = hbusreq1_p & f2f29d | !hbusreq1_p & v845542;
assign v1215075 = hbusreq2 & v1215071 | !hbusreq2 & v1215074;
assign v14465cb = hgrant4_p & v144640c | !hgrant4_p & v14465ca;
assign v121531e = hmaster0_p & v1215471 | !hmaster0_p & v1215462;
assign v12adf5e = hmaster2_p & v845542 | !hmaster2_p & !v12adf5d;
assign v1668cf1 = hmaster0_p & a658ad | !hmaster0_p & v1668cf0;
assign v1214ecd = hbusreq5_p & v1214ecb | !hbusreq5_p & v1214ecc;
assign v118e18f = stateG3_0_p & v845586 | !stateG3_0_p & v845542;
assign d302eb = hgrant2_p & v845542 | !hgrant2_p & !d302ea;
assign v1215c4f = hgrant2_p & v121657d | !hgrant2_p & v1215c47;
assign v10d3fe6 = hbusreq0_p & v10d3fdb | !hbusreq0_p & v10d3fe0;
assign v151584e = hbusreq2 & v151584d | !hbusreq2 & v1516803;
assign v10d3fda = hmaster2_p & v10d3fd5 | !hmaster2_p & !v10d3fd9;
assign v1445861 = hlock2 & v14457f6 | !hlock2 & v1445860;
assign d2fb17 = hbusreq2 & d2fb13 | !hbusreq2 & d2fb16;
assign v1215c0a = hbusreq1 & v121611d | !hbusreq1 & v845547;
assign v121532f = hmaster1_p & v1215320 | !hmaster1_p & !v121507b;
assign v1445862 = hbusreq2 & v144585b | !hbusreq2 & v1445861;
assign v138a350 = hmaster0_p & v138a32d | !hmaster0_p & v138a34f;
assign v134d4e9 = hbusreq1_p & v134d273 | !hbusreq1_p & v134d4e8;
assign v1214fc4 = hbusreq0 & v12157a2 | !hbusreq0 & v1214fc3;
assign v10d42a8 = hgrant2_p & v10d4081 | !hgrant2_p & v10d42a7;
assign v16a1ad9 = hgrant4_p & v845559 | !hgrant4_p & v16a1ad8;
assign d2fc67 = hbusreq1_p & d2fbf5 | !hbusreq1_p & d2fc66;
assign v15155f2 = hmaster0_p & v845570 | !hmaster0_p & v15155f1;
assign v14459f0 = hbusreq5_p & v14459e9 | !hbusreq5_p & v14459ef;
assign v14460ef = hmaster0_p & v1445f85 | !hmaster0_p & v144639c;
assign v12afe54 = hgrant0_p & v12afe53 | !hgrant0_p & !v845542;
assign v121602e = hmaster2_p & v845542 | !hmaster2_p & v121602d;
assign v1214c54 = hgrant5_p & v1215365 | !hgrant5_p & v1214c52;
assign v1215cc6 = hbusreq5_p & v1215cc4 | !hbusreq5_p & !v1215cc5;
assign v1216547 = hmaster2_p & v845542 | !hmaster2_p & v1216546;
assign v1216ad5 = hlock4_p & v1216ad4 | !hlock4_p & v845547;
assign v1446441 = hmaster0_p & v144639c | !hmaster0_p & v1446440;
assign d30851 = hmaster0_p & d3084d | !hmaster0_p & d30850;
assign d2fb4e = hlock0_p & v845542 | !hlock0_p & a66295;
assign v1445e4d = hmaster2_p & v845542 | !hmaster2_p & v1445e38;
assign v16a1376 = hmaster1_p & v16a132f | !hmaster1_p & v16a1f96;
assign d3094a = hburst1_p & v845542 | !hburst1_p & v893df7;
assign d306d0 = hbusreq1_p & d306cf | !hbusreq1_p & v845542;
assign v14458da = hbusreq0_p & v14458d9 | !hbusreq0_p & v1446406;
assign v1215084 = hbusreq2 & v1215080 | !hbusreq2 & v1215083;
assign d306d9 = hbusreq5_p & d306d3 | !hbusreq5_p & d306d8;
assign d2fd1c = hgrant5_p & v845542 | !hgrant5_p & !d3064b;
assign v15533a6 = hmaster2_p & v15533a5 | !hmaster2_p & v15533a2;
assign d2fec0 = hbusreq4_p & d2febf | !hbusreq4_p & v845542;
assign v1445d85 = hbusreq1_p & v144639c | !hbusreq1_p & v1445d84;
assign d2f96e = hbusreq1_p & d300d8 | !hbusreq1_p & d2f96d;
assign a65616 = hmaster1_p & a65615 | !hmaster1_p & a653e7;
assign v16a13da = hready_p & v845555 | !hready_p & v16a13d9;
assign v16a2665 = busreq_p & v16a2664 | !busreq_p & v845542;
assign d308de = hmaster1_p & v845542 | !hmaster1_p & d308dd;
assign v1445a92 = hbusreq2 & v1445a8d | !hbusreq2 & v1445a91;
assign v134d3bd = hgrant3_p & v134d278 | !hgrant3_p & v134d3bc;
assign v16a1cc0 = hmaster1_p & v16a1ca4 | !hmaster1_p & v16a1f96;
assign v144546b = hlock0 & v1445469 | !hlock0 & v1446635;
assign v1216ab9 = hready & v1446397 | !hready & !f2f4ad;
assign v12afe65 = hbusreq0 & v12afe52 | !hbusreq0 & v12afe64;
assign v1445b2a = hlock5 & v1445af2 | !hlock5 & v1445b28;
assign v1214d62 = hmaster1_p & v1214d51 | !hmaster1_p & v1214d5f;
assign v1553386 = hmaster2_p & v1553217 | !hmaster2_p & v845542;
assign v1668c52 = hlock3_p & v1668c51 | !hlock3_p & v845542;
assign v1445b01 = hmaster0_p & v1445a6b | !hmaster0_p & v14458d4;
assign v134d504 = hbusreq0_p & v134d273 | !hbusreq0_p & v134d36d;
assign d2fefb = hlock2_p & d2fef9 | !hlock2_p & d2fefa;
assign a656c8 = hbusreq0 & a66287 | !hbusreq0 & a65b2b;
assign v14463df = hlock0 & v14463de | !hlock0 & v14463dd;
assign v1445fd1 = hbusreq5_p & v1445fcb | !hbusreq5_p & v1445fd0;
assign v12ad60b = hgrant5_p & v12ad609 | !hgrant5_p & !v12ad5c5;
assign v16a138c = hbusreq2_p & v16a129e | !hbusreq2_p & v16a138b;
assign v1446741 = hmaster1_p & v1446740 | !hmaster1_p & v1446436;
assign v121622d = hmaster1_p & v121622c | !hmaster1_p & v1216224;
assign v134d279 = hmaster0_p & v845542 | !hmaster0_p & v134d1de;
assign v1668d05 = hmaster1_p & v1668cd9 | !hmaster1_p & !v1668cfd;
assign v15157da = hgrant5_p & v845570 | !hgrant5_p & v151572e;
assign v16a19e6 = hbusreq2_p & v16a1847 | !hbusreq2_p & v16a19e5;
assign v1216158 = hgrant5_p & v121600b | !hgrant5_p & v1216157;
assign v15156b3 = hlock2_p & v151566c | !hlock2_p & !v15156b2;
assign v16a196b = hgrant2_p & v845542 | !hgrant2_p & v16a1969;
assign v1215c88 = hmaster2_p & v1215c87 | !hmaster2_p & v845542;
assign v10d4001 = hlock3_p & v10d3fee | !hlock3_p & !v10d4000;
assign v1389fb3 = hbusreq3 & v1389f98 | !hbusreq3 & v138a391;
assign v1445857 = hbusreq2_p & v1445854 | !hbusreq2_p & v1445856;
assign v155308d = hmaster1_p & v155308c | !hmaster1_p & v845542;
assign v121652f = hmaster2_p & v121652b | !hmaster2_p & v121652e;
assign v144624e = hbusreq0 & v144624d | !hbusreq0 & v1446214;
assign v144603e = hmaster2_p & v144603d | !hmaster2_p & v14465b3;
assign v1215d7d = hmaster1_p & v1215d7c | !hmaster1_p & v1215d68;
assign a65458 = hgrant3_p & a6592b | !hgrant3_p & a65457;
assign v10d4008 = hmaster1_p & v10d4007 | !hmaster1_p & v10d3ffb;
assign v12150ce = hbusreq4_p & v12150cd | !hbusreq4_p & v845542;
assign d305eb = hmaster2_p & v16693aa | !hmaster2_p & !d305ea;
assign a6628b = hgrant1_p & v845542 | !hgrant1_p & !a66289;
assign v1216056 = hmaster2_p & v1216053 | !hmaster2_p & v1216055;
assign v144607e = hmaster2_p & v144603d | !hmaster2_p & v144604f;
assign v16a1da8 = hbusreq2 & v16a1da4 | !hbusreq2 & v16a1da7;
assign v16a1a93 = hmaster2_p & v16a1a92 | !hmaster2_p & !v845542;
assign d30858 = hmaster0_p & d30853 | !hmaster0_p & d30857;
assign v10d42c1 = hmaster1_p & v10d42c0 | !hmaster1_p & !v10d404f;
assign v151699b = hlock2_p & v151699a | !hlock2_p & v845542;
assign v1214e65 = hbusreq2_p & v1214e64 | !hbusreq2_p & v845542;
assign f2f442 = hmaster0_p & f2f3d8 | !hmaster0_p & f2f3be;
assign v10d3ffd = hmaster2_p & v10d3fd4 | !hmaster2_p & !v10d3fdf;
assign v1389de1 = hbusreq5_p & v1389de0 | !hbusreq5_p & !v845542;
assign d3070e = hmaster2_p & v84554e | !hmaster2_p & !d3070d;
assign v10d3ff5 = hmaster2_p & v10d3fdf | !hmaster2_p & !v10d3ff3;
assign v121623c = hmaster0_p & v1216236 | !hmaster0_p & v1216209;
assign f2f39c = hbusreq5_p & f2f398 | !hbusreq5_p & !f2f39b;
assign v16a1965 = hgrant5_p & v845542 | !hgrant5_p & !v16a1956;
assign v1515614 = hlock0_p & a65851 | !hlock0_p & v1515613;
assign v1515827 = hlock2_p & v1515826 | !hlock2_p & !v1515702;
assign f2f230 = hgrant1_p & f2f22f | !hgrant1_p & !v845542;
assign v144623f = hlock2 & v144623c | !hlock2 & v144623e;
assign v12afdb1 = hmaster2_p & v845542 | !hmaster2_p & !v84554a;
assign v12ad0b1 = hgrant1_p & v12ad0b0 | !hgrant1_p & v12afda6;
assign d302f2 = hready_p & d308d5 | !hready_p & d302f1;
assign v134cec5 = hlock3 & v134d3b5 | !hlock3 & v134cec4;
assign v1445a61 = hmaster0_p & v14459f0 | !hmaster0_p & v1445a1f;
assign bf1f77 = hgrant0_p & bf1f52 | !hgrant0_p & !v84556a;
assign v10d42c5 = hgrant0_p & v10d401b | !hgrant0_p & !v10d42c4;
assign v1552da3 = jx1_p & v155351c | !jx1_p & v1552da2;
assign v1284d5b = hmaster0_p & v1284cbc | !hmaster0_p & v1284cb9;
assign v1214f3c = hbusreq2 & v1214f3b | !hbusreq2 & v845542;
assign v12ad5cb = hgrant1_p & v12ad5ca | !hgrant1_p & v12ad5c2;
assign v16a1a2b = hmaster1_p & v16a19df | !hmaster1_p & !v16a1f96;
assign a6590e = hmaster1_p & a6590b | !hmaster1_p & a658e5;
assign v1405abd = hmaster2_p & v1405abb | !hmaster2_p & !v845542;
assign v1515786 = hmaster0_p & v151575e | !hmaster0_p & v1515785;
assign d2fc88 = hmaster0_p & d305df | !hmaster0_p & v1668da6;
assign v121502c = hbusreq4_p & v121502b | !hbusreq4_p & v845542;
assign v14460a7 = hmaster1_p & v14460a6 | !hmaster1_p & v1445fde;
assign v12157ab = hbusreq4 & v1216528 | !hbusreq4 & !v12157aa;
assign v1214c22 = hlock2_p & v1214c20 | !hlock2_p & v1214c21;
assign d2fc3e = hbusreq2_p & d2fbb7 | !hbusreq2_p & d2fc3c;
assign v1445492 = hbusreq2 & v1445490 | !hbusreq2 & v1445491;
assign v1216a5a = hready & v845542 | !hready & v845570;
assign v12af98a = hmaster2_p & d30690 | !hmaster2_p & !v12af989;
assign v1668d3b = hgrant4_p & v1668d26 | !hgrant4_p & a65382;
assign d2ff02 = hmaster1_p & d2fef8 | !hmaster1_p & d2fee5;
assign v1446059 = hbusreq1_p & v1446058 | !hbusreq1_p & v1446608;
assign v1215c15 = hgrant1_p & v1215c14 | !hgrant1_p & v1216123;
assign v1405afe = hgrant5_p & v1405ad9 | !hgrant5_p & !v1405afd;
assign v1446325 = hgrant2_p & v144631e | !hgrant2_p & v1446324;
assign v14466c4 = hlock5 & v1446676 | !hlock5 & v14466bf;
assign v1445ae5 = hmaster0_p & v1445a38 | !hmaster0_p & v14458d4;
assign v12aed9e = decide_p & v12af9b6 | !decide_p & v845542;
assign v1446233 = hlock0 & v1446232 | !hlock0 & v144622e;
assign v10d4010 = hmaster1_p & v10d400f | !hmaster1_p & !v10d3fe9;
assign v155338c = hbusreq4 & v155338a | !hbusreq4 & v155338b;
assign v15530ec = hbusreq2_p & v1552d62 | !hbusreq2_p & v155341e;
assign v1215713 = hgrant0_p & v1215712 | !hgrant0_p & !v845542;
assign v14463d8 = hbusreq4 & v14463d6 | !hbusreq4 & v14463d7;
assign v1515aea = hmaster1_p & v1515ae9 | !hmaster1_p & a65893;
assign d3077e = hmaster1_p & d3077d | !hmaster1_p & d306e4;
assign v10d4273 = hgrant5_p & v10d3feb | !hgrant5_p & v10d4272;
assign v1445dc6 = hbusreq2_p & v1445dc3 | !hbusreq2_p & v1445dc5;
assign v1445f5c = hgrant2_p & v1445f5b | !hgrant2_p & v1445f56;
assign v1214ccd = hmaster2_p & v1214cc7 | !hmaster2_p & !v1215380;
assign v1668c38 = hgrant3_p & v1668c35 | !hgrant3_p & !v1668c37;
assign v1446260 = hbusreq5 & v144625e | !hbusreq5 & v144625f;
assign bf1f5f = hgrant1_p & v845570 | !hgrant1_p & d30649;
assign v1445d89 = hmaster2_p & v1445d88 | !hmaster2_p & v1445d85;
assign d307fd = hlock5_p & d307fb | !hlock5_p & !d307fc;
assign v12162d6 = hbusreq2 & v12162d2 | !hbusreq2 & v12162d5;
assign v1405a7e = hmaster2_p & v1405a7d | !hmaster2_p & !v845542;
assign d307a9 = hgrant5_p & d307a7 | !hgrant5_p & d307a8;
assign v16a1978 = hgrant2_p & v845542 | !hgrant2_p & v16a1977;
assign d30856 = hmaster2_p & d30854 | !hmaster2_p & d30855;
assign v121575e = hgrant4_p & v845542 | !hgrant4_p & v121575d;
assign v1405b5f = hgrant2_p & v1405b5c | !hgrant2_p & v1405b5e;
assign d2fbf4 = hbusreq4_p & d2fbf3 | !hbusreq4_p & v84554a;
assign v1215366 = hbusreq1_p & v1215364 | !hbusreq1_p & v845547;
assign v16a1337 = hgrant2_p & v16a205c | !hgrant2_p & v16a1336;
assign v144615a = hlock3 & v1446125 | !hlock3 & v1446159;
assign v1516804 = hbusreq2 & v1516801 | !hbusreq2 & v1516803;
assign v12164d0 = stateA1_p & v1216aaf | !stateA1_p & !a66292;
assign a65378 = hmaster2_p & a65372 | !hmaster2_p & a65377;
assign v15530a6 = decide_p & v1553216 | !decide_p & v15530a5;
assign d30804 = hbusreq0 & d307fe | !hbusreq0 & d30803;
assign v1214ee3 = hbusreq5_p & v1214ee2 | !hbusreq5_p & v1214ee1;
assign v134d21c = hbusreq2_p & v134d21b | !hbusreq2_p & v134d20c;
assign v1214ec6 = decide_p & v1214ec1 | !decide_p & v1214ec5;
assign v14457a7 = hmaster1_p & v14457a6 | !hmaster1_p & v1445e07;
assign v1515672 = stateA1_p & v1515670 | !stateA1_p & v1515671;
assign d301eb = hbusreq1_p & v845542 | !hbusreq1_p & d307b3;
assign bf1f62 = hmaster2_p & v845570 | !hmaster2_p & !v845542;
assign v1515823 = hbusreq2_p & v1515822 | !hbusreq2_p & v845542;
assign ab8d68 = stateG3_2_p & v88d3e4 | !stateG3_2_p & !afe156;
assign v1216ad0 = hlock5_p & v1216ac3 | !hlock5_p & v1216acf;
assign f2f284 = hbusreq5_p & f2f229 | !hbusreq5_p & f2f283;
assign v144581f = hgrant2_p & v144581d | !hgrant2_p & v144581e;
assign v1445f40 = hbusreq2_p & v1445f3a | !hbusreq2_p & v1445f3f;
assign v1216051 = hbusreq1 & v1216adf | !hbusreq1 & v845542;
assign v1214c1a = hbusreq2 & v1214c15 | !hbusreq2 & v1214c19;
assign d2fb8a = hbusreq2 & d2fb82 | !hbusreq2 & d2fb89;
assign v155337f = hmaster0_p & v845542 | !hmaster0_p & v1553218;
assign v1405ad7 = hmaster2_p & v1405ad6 | !hmaster2_p & !v845542;
assign v1405861 = hmaster2_p & v1405860 | !hmaster2_p & v140583e;
assign v121577b = hgrant5_p & v1215b8a | !hgrant5_p & v121577a;
assign v12ad321 = hbusreq4_p & v12ae1f8 | !hbusreq4_p & v12af9cf;
assign v144550c = hgrant2_p & v144550a | !hgrant2_p & v144550b;
assign v1215d6c = hgrant5_p & v1215d63 | !hgrant5_p & v1215d6b;
assign v1446108 = hlock2 & v14460f2 | !hlock2 & v1446106;
assign v121573d = hgrant1_p & v1215736 | !hgrant1_p & v121573c;
assign v16a137e = hbusreq3 & v16a1378 | !hbusreq3 & v16a137d;
assign v16a1bf6 = hmaster0_p & v16a1bf5 | !hmaster0_p & v16a1bf2;
assign v138a3ab = hmaster1_p & v138a3aa | !hmaster1_p & v138a341;
assign v1446236 = hmaster0_p & v1446233 | !hmaster0_p & v1446235;
assign v1445379 = hmaster1_p & v1445b31 | !hmaster1_p & v144591b;
assign v16a1d80 = hbusreq3 & v16a1d7f | !hbusreq3 & v16a209f;
assign v134cd8a = hlock5 & v134cd7a | !hlock5 & v134cd89;
assign v138938d = hbusreq5_p & v138938c | !hbusreq5_p & v845542;
assign v16a1ac2 = hbusreq2_p & v16a2677 | !hbusreq2_p & v16a1ac1;
assign d2fc4d = hgrant4_p & d2fbce | !hgrant4_p & d2fc4c;
assign d3067b = hbusreq5_p & v845542 | !hbusreq5_p & d30663;
assign v12afe44 = hgrant0_p & a6537d | !hgrant0_p & !v845542;
assign v10d42c3 = hbusreq0_p & v10d4267 | !hbusreq0_p & v10d40ba;
assign d308aa = hgrant5_p & d30856 | !hgrant5_p & d308a9;
assign v1216049 = hlock1_p & v1216048 | !hlock1_p & !v845542;
assign v1215c3e = hgrant5_p & v1215c3c | !hgrant5_p & v1215c3d;
assign v1446107 = hlock2 & v1446104 | !hlock2 & v1446106;
assign v12153b5 = hmaster2_p & v1215bac | !hmaster2_p & v12153b4;
assign v16a131c = busreq_p & d80758 | !busreq_p & !d80757;
assign v1445a03 = hmaster2_p & v1445a02 | !hmaster2_p & v14459fc;
assign v12aee5d = hready_p & v12aedde | !hready_p & v12aee5c;
assign v1445f74 = hgrant2_p & v144674c | !hgrant2_p & v1445f73;
assign v1446733 = hgrant2_p & v1446730 | !hgrant2_p & v1446732;
assign v121600a = hbusreq1_p & v1216009 | !hbusreq1_p & v845542;
assign d305ed = hbusreq5_p & d305ec | !hbusreq5_p & v845542;
assign d30838 = hgrant5_p & v84554e | !hgrant5_p & d307ff;
assign v121659d = hbusreq0_p & v1216a8d | !hbusreq0_p & !v1216594;
assign v12161cf = hbusreq1_p & v12161ce | !hbusreq1_p & v845542;
assign v134d4b7 = hlock5 & v134d4a8 | !hlock5 & v134d4b6;
assign v14458be = hbusreq5_p & v1445886 | !hbusreq5_p & v14458bd;
assign v151576c = hlock0_p & v1668d24 | !hlock0_p & v151576b;
assign v16a1ad6 = decide_p & v16a1ad5 | !decide_p & v16a2065;
assign v1284cc9 = hgrant5_p & v1405856 | !hgrant5_p & v1284cc8;
assign a64704 = hbusreq2_p & a65b0d | !hbusreq2_p & a65b29;
assign v14459fc = hgrant1_p & v14459f4 | !hgrant1_p & v14459fb;
assign d308b3 = hbusreq2_p & d308b1 | !hbusreq2_p & d308b2;
assign v1445a68 = hgrant2_p & v1445a65 | !hgrant2_p & v1445a67;
assign d300b5 = hbusreq1 & d2fe7b | !hbusreq1 & d2fe80;
assign v1216b13 = hmaster1_p & v1216b03 | !hmaster1_p & v1216af8;
assign v1405864 = hmaster2_p & v140583e | !hmaster2_p & v1405863;
assign v12166e9 = hgrant4_p & v12164de | !hgrant4_p & !v12166e8;
assign d30630 = hmaster0_p & d30628 | !hmaster0_p & d3062c;
assign v1215d7b = hgrant2_p & v1215d69 | !hgrant2_p & v1215d7a;
assign v12ad573 = hmaster1_p & v12ad572 | !hmaster1_p & !v12ad525;
assign v1216b06 = hlock2_p & v1216b05 | !hlock2_p & v1216afd;
assign v1553059 = hlock1 & v155339c | !hlock1 & v1553058;
assign v12acfdf = hmaster1_p & v12acfbe | !hmaster1_p & v12ad54f;
assign v134d38a = hmaster2_p & v134d389 | !hmaster2_p & v134d386;
assign v1445f41 = hlock2 & v1445f40 | !hlock2 & v1445f37;
assign v1445a9e = hmaster1_p & v1445a44 | !hmaster1_p & v1445a9b;
assign f2e3f7 = hgrant5_p & v845542 | !hgrant5_p & !f2e3f6;
assign v1446723 = decide_p & v14466ef | !decide_p & v1446722;
assign v16a143c = hmaster1_p & v16a143b | !hmaster1_p & v16a1d53;
assign v14466c6 = decide_p & v1446402 | !decide_p & v14466c5;
assign v1445d90 = hmaster2_p & v14463b1 | !hmaster2_p & !v1445f97;
assign v134d460 = hmaster1_p & v134d45f | !hmaster1_p & v845542;
assign v84554c = hbusreq1_p & v845542 | !hbusreq1_p & !v845542;
assign v10d403b = hmaster2_p & v10d403a | !hmaster2_p & !v10d4032;
assign a6567c = hbusreq2_p & a65665 | !hbusreq2_p & a6567b;
assign v1446094 = hmaster1_p & v1446093 | !hmaster1_p & v1446073;
assign v155322d = hbusreq5_p & v155322c | !hbusreq5_p & v155322b;
assign d2fb99 = hmaster2_p & d2fb83 | !hmaster2_p & d2fb70;
assign v12166f9 = hmaster1_p & v12166f8 | !hmaster1_p & v12166ef;
assign v16a1959 = hgrant5_p & v845542 | !hgrant5_p & v16a1958;
assign v16a1a98 = hmaster0_p & v16a1a94 | !hmaster0_p & v16a1a97;
assign d305e7 = decide_p & d305e6 | !decide_p & v845570;
assign v1284d3b = hbusreq1_p & v140588d | !hbusreq1_p & v1284d3a;
assign a654af = hbusreq5_p & a654ad | !hbusreq5_p & a654ae;
assign v134d3c6 = hmaster1_p & v134d3c3 | !hmaster1_p & v134d20f;
assign v140589c = hgrant1_p & v140589b | !hgrant1_p & v1405845;
assign v1214e0e = hbusreq0 & v1216adb | !hbusreq0 & v1214e0d;
assign v134cd62 = hbusreq4_p & v134cd61 | !hbusreq4_p & v134d384;
assign v1668c79 = hmaster2_p & a658c6 | !hmaster2_p & !v1668c77;
assign v1216566 = hgrant1_p & v1216522 | !hgrant1_p & v1216565;
assign v1405a90 = hbusreq4_p & v845542 | !hbusreq4_p & !v1405a87;
assign v10d407c = hmaster0_p & v10d4070 | !hmaster0_p & !v10d407b;
assign a66275 = hmastlock_p & a66273 | !hmastlock_p & !v845542;
assign v155322e = hlock4_p & v1553138 | !hlock4_p & v845542;
assign d301df = hlock5_p & d301d3 | !hlock5_p & !d301de;
assign v138a0c7 = jx1_p & v1389f82 | !jx1_p & v138a0c6;
assign v85e75f = hmaster1_p & v84555c | !hmaster1_p & !v90d5cd;
assign d2fcec = hbusreq2_p & d2fceb | !hbusreq2_p & d302d6;
assign v1215c56 = hbusreq0 & v1215c54 | !hbusreq0 & v1215c55;
assign d30734 = hbusreq1_p & d30733 | !hbusreq1_p & v845542;
assign v1515816 = hbusreq2 & v1515815 | !hbusreq2 & !v845542;
assign v16a1d3c = hgrant1_p & v84554d | !hgrant1_p & v16a1bc2;
assign v1552da0 = hgrant3_p & v1552d9d | !hgrant3_p & v1552d9f;
assign a64709 = hready_p & a64707 | !hready_p & a64708;
assign v1445755 = hlock3 & v1445f40 | !hlock3 & v1445753;
assign d2fea5 = hmaster0_p & d2fe9b | !hmaster0_p & d2fea4;
assign d2fd0f = hmaster1_p & d3060a | !hmaster1_p & !d2fcb5;
assign v140591d = hmaster0_p & v1405859 | !hmaster0_p & v1405855;
assign d30953 = hmaster2_p & d305ea | !hmaster2_p & d30952;
assign v121502e = hgrant1_p & v1215bac | !hgrant1_p & v121502d;
assign v1215cda = hmaster0_p & v845542 | !hmaster0_p & v1215cd9;
assign v12ad618 = hmaster1_p & v12ad602 | !hmaster1_p & !v12ad617;
assign v1445fdd = hlock0 & v1445fda | !hlock0 & v1445fdc;
assign v1515856 = jx1_p & v1515608 | !jx1_p & v1515855;
assign v12ad627 = decide_p & v12ad626 | !decide_p & v12afe76;
assign v1445ad2 = hmaster1_p & v1445ab8 | !hmaster1_p & v14458c1;
assign v1215469 = hmaster2_p & v1215466 | !hmaster2_p & v1215467;
assign a656c0 = hmaster0_p & a656bc | !hmaster0_p & a656be;
assign d30674 = hmaster0_p & d305d7 | !hmaster0_p & d30673;
assign v151583f = hgrant2_p & v15167ff | !hgrant2_p & !v151583e;
assign v16a1952 = hgrant0_p & v845542 | !hgrant0_p & v16a1948;
assign a658c3 = hburst0 & v10d3fde | !hburst0 & a658c1;
assign v138a3f8 = hmaster0_p & v845542 | !hmaster0_p & v138a3f7;
assign v1445a57 = hmaster2_p & v14459a0 | !hmaster2_p & v1445a53;
assign v12161ec = hbusreq1 & v121659b | !hbusreq1 & v845542;
assign v1214dc3 = hbusreq2_p & v1214dc0 | !hbusreq2_p & v1214dc2;
assign v1389d74 = hmaster0_p & v1389d73 | !hmaster0_p & v845542;
assign d3020e = hlock5_p & d3020c | !hlock5_p & d3020d;
assign v1515749 = hgrant1_p & v1515743 | !hgrant1_p & v1515748;
assign v121546c = hlock0_p & v12160f2 | !hlock0_p & v121546b;
assign d30257 = hbusreq0 & d30255 | !hbusreq0 & d30256;
assign v14465f8 = hlock0_p & v14463b1 | !hlock0_p & v14463e5;
assign d301bd = hmaster2_p & v845542 | !hmaster2_p & d301bc;
assign v10d4044 = hbusreq1_p & v10d3fe7 | !hbusreq1_p & !v10d3ff9;
assign v121536b = hmaster0_p & v1215369 | !hmaster0_p & v121536a;
assign v1553221 = hgrant4_p & v845542 | !hgrant4_p & v1553220;
assign v134d43f = hbusreq0 & v134d43e | !hbusreq0 & v134d274;
assign v1515c7e = hbusreq4 & v1515c7d | !hbusreq4 & d3094f;
assign v134d3cb = hlock3 & v134d3c7 | !hlock3 & v134d3ca;
assign v11e5962 = hmaster2_p & v845542 | !hmaster2_p & !v11e5961;
assign v134cd5b = hmaster2_p & v845542 | !hmaster2_p & v134cd5a;
assign v1668cc3 = hburst0 & v156645f | !hburst0 & v1668cc2;
assign v1445925 = hbusreq3 & v1445923 | !hbusreq3 & v1445924;
assign v1552d8a = hgrant4_p & v845542 | !hgrant4_p & v1552d89;
assign d307bd = hlock1_p & d307bc | !hlock1_p & d30649;
assign v144546e = hbusreq2_p & v144546d | !hbusreq2_p & v1445bba;
assign f2e4d7 = hbusreq0 & f2f51a | !hbusreq0 & f2ed96;
assign v1215cfb = hmaster1_p & v1215cec | !hmaster1_p & v1215cfa;
assign d30125 = hmaster2_p & d2fe80 | !hmaster2_p & d30124;
assign v12aec47 = hbusreq0 & v12afe51 | !hbusreq0 & v12afe5e;
assign v12ad325 = hmaster2_p & v12af9d3 | !hmaster2_p & v12ad324;
assign v144640c = hbusreq4 & v1446406 | !hbusreq4 & v144640b;
assign d308c1 = hbusreq0 & d308be | !hbusreq0 & d308c0;
assign v1215111 = decide_p & v121510b | !decide_p & v1215110;
assign a65625 = hgrant5_p & a653f9 | !hgrant5_p & a65624;
assign f2f45c = hbusreq5 & f2f441 | !hbusreq5 & f2f45b;
assign v1214da2 = hmaster1_p & v1214da1 | !hmaster1_p & v1215388;
assign v144589f = hmaster0_p & v144588f | !hmaster0_p & v144589e;
assign v140586d = hlock0_p & v140583e | !hlock0_p & v14463b1;
assign v14453f7 = hbusreq2 & v14453f4 | !hbusreq2 & v14453f6;
assign d30139 = hgrant5_p & d30138 | !hgrant5_p & d300e0;
assign v138a45f = hmaster1_p & v138a45e | !hmaster1_p & v138a341;
assign v1389380 = hgrant2_p & v845542 | !hgrant2_p & !v138937f;
assign d8074e = hmaster1_p & d8074d | !hmaster1_p & d80746;
assign v121506f = hmaster1_p & v121506e | !hmaster1_p & v1215054;
assign d2fcb8 = hbusreq2_p & d2fcb7 | !hbusreq2_p & d302d6;
assign v1284d1e = hgrant5_p & v144642a | !hgrant5_p & v1284d1d;
assign v1445551 = hbusreq2_p & v144554e | !hbusreq2_p & v1445550;
assign v134d44b = hgrant5_p & v134d44a | !hgrant5_p & v134d378;
assign v1215be3 = hmaster1_p & v1215bdc | !hmaster1_p & v1215be2;
assign v1215c99 = hgrant1_p & v1215c93 | !hgrant1_p & v121610d;
assign v1553392 = hgrant5_p & v1553386 | !hgrant5_p & v1553391;
assign v12161a0 = hgrant5_p & v845542 | !hgrant5_p & v1216179;
assign v14462a0 = hbusreq3 & v1446277 | !hbusreq3 & v144629f;
assign v1445e3a = hgrant1_p & v1445e39 | !hgrant1_p & v845542;
assign v12166d3 = hmaster2_p & v845542 | !hmaster2_p & v12166d2;
assign v12166cd = locked_p & v12166cc | !locked_p & v845542;
assign v12ad5ac = hlock0_p & v1668d25 | !hlock0_p & !v845542;
assign v16a1382 = hgrant3_p & v16a12e5 | !hgrant3_p & v16a1381;
assign v1446658 = hmaster0_p & v1446404 | !hmaster0_p & v1446657;
assign v144670e = hlock2 & v1446707 | !hlock2 & v144670d;
assign d2fb40 = hbusreq2 & d2fb3e | !hbusreq2 & d2fb3f;
assign v151563a = hmaster0_p & v1515638 | !hmaster0_p & v1515639;
assign v16a16a8 = hbusreq5_p & v16a1d77 | !hbusreq5_p & v16a16a7;
assign v1446428 = hbusreq0_p & v1446403 | !hbusreq0_p & v1446406;
assign v1445420 = hmaster1_p & v14465aa | !hmaster1_p & v144627e;
assign d2fefa = hmaster1_p & d2fec8 | !hmaster1_p & d2fec6;
assign v1668cdb = hburst1 & v156645f | !hburst1 & v1668cda;
assign v1445b66 = hmaster1_p & v1446313 | !hmaster1_p & v1445b5f;
assign v15157b5 = stateA1_p & v845542 | !stateA1_p & !v15157b4;
assign v10d3ff1 = hmaster2_p & v10d3fd4 | !hmaster2_p & v10d3fd8;
assign v1445472 = hbusreq0 & v1446654 | !hbusreq0 & v144639c;
assign f2ed94 = hgrant2_p & v845542 | !hgrant2_p & f2ed93;
assign v10d3fd7 = hmastlock_p & v10d3fd6 | !hmastlock_p & !v845542;
assign v16a1bc9 = hbusreq1 & v16a1bc8 | !hbusreq1 & v16a2089;
assign v12acfd2 = hlock2_p & v12acfcf | !hlock2_p & v12acfd1;
assign v1445471 = hbusreq2 & v144546e | !hbusreq2 & v1445470;
assign v1216548 = hlock5_p & v1216543 | !hlock5_p & v1216547;
assign v1516900 = decide_p & v15168ff | !decide_p & v845576;
assign v1445e08 = hmaster1_p & v1445de8 | !hmaster1_p & v1445e07;
assign bf1f54 = hmaster0_p & v84556a | !hmaster0_p & bf1f53;
assign v1445863 = hlock3 & v1445852 | !hlock3 & v1445862;
assign v1668cf2 = hmaster1_p & v1668cf1 | !hmaster1_p & v1668cd6;
assign v121576a = hgrant1_p & v1215757 | !hgrant1_p & v1215769;
assign v1215c28 = hbusreq1_p & v1216005 | !hbusreq1_p & v1215c27;
assign v16a1bd0 = hgrant5_p & v845542 | !hgrant5_p & v16a1bcf;
assign d3025e = hbusreq2_p & d3025c | !hbusreq2_p & d3025d;
assign v1445489 = hbusreq2 & v144547c | !hbusreq2 & v1445482;
assign v1214816 = hbusreq3 & v1214800 | !hbusreq3 & v1214815;
assign v10d429a = hgrant5_p & v10d406c | !hgrant5_p & v10d4299;
assign d305f0 = hmastlock_p & f2f4ad | !hmastlock_p & v845542;
assign v1284d20 = hmaster1_p & v1284d0e | !hmaster1_p & !v1284d1f;
assign d30143 = hbusreq5_p & d30141 | !hbusreq5_p & d30142;
assign d3069c = hbusreq5_p & v845542 | !hbusreq5_p & d30691;
assign d30251 = hmaster1_p & d30240 | !hmaster1_p & d30250;
assign v10d4073 = hgrant4_p & v10d4071 | !hgrant4_p & !v10d4072;
assign v14463f5 = hbusreq0 & v14463f4 | !hbusreq0 & v14463c7;
assign d308cf = hbusreq5 & d308b4 | !hbusreq5 & d308ce;
assign v10d3ff8 = hbusreq0_p & v10d3fd8 | !hbusreq0_p & !v10d3fdf;
assign v1446661 = hbusreq5_p & v1446660 | !hbusreq5_p & v1446643;
assign v1405aa3 = hmaster2_p & v1405aa2 | !hmaster2_p & v1405a87;
assign v12ad5a9 = hbusreq1 & v12ad4d0 | !hbusreq1 & v12ad4e4;
assign v16a1e74 = hmaster1_p & v16a1e68 | !hmaster1_p & !v16a1f96;
assign v121543d = hmaster1_p & v121543c | !hmaster1_p & v121540f;
assign v1445ef1 = hmaster1_p & v14465b7 | !hmaster1_p & v1445ef0;
assign v12afa0c = hmaster0_p & v12af9c3 | !hmaster0_p & v12afa0b;
assign v1446004 = hbusreq2 & v1446002 | !hbusreq2 & v1446003;
assign v134d3d6 = hbusreq5 & v134d3d5 | !hbusreq5 & v134d276;
assign v10d4025 = hmaster2_p & v10d401e | !hmaster2_p & v10d4024;
assign v12ad31a = hbusreq4_p & v12afe4d | !hbusreq4_p & v12af9bd;
assign v16a2667 = stateA1_p & v16a2665 | !stateA1_p & v16a2666;
assign v12162c1 = hgrant2_p & v12162be | !hgrant2_p & v12162c0;
assign v16a1d94 = hgrant2_p & v16a2059 | !hgrant2_p & v16a1d93;
assign v1668de7 = hbusreq5 & v1668db1 | !hbusreq5 & v1668de6;
assign v1215b98 = hmaster2_p & v12160ec | !hmaster2_p & !v1215b97;
assign d308a1 = hgrant1_p & v84554c | !hgrant1_p & d308a0;
assign a653fc = hbusreq5_p & a653f8 | !hbusreq5_p & a653fa;
assign v1214cdb = hmaster2_p & d2fbe5 | !hmaster2_p & !v1214cc7;
assign d30273 = hmaster0_p & d3026d | !hmaster0_p & d30272;
assign d2fe99 = hbusreq3 & d2fe91 | !hbusreq3 & d2fe98;
assign v134d452 = hgrant2_p & v134d442 | !hgrant2_p & v134d450;
assign v1446475 = stateA1_p & v144646d | !stateA1_p & v1446468;
assign v1445f7a = hlock2 & v144673f | !hlock2 & v1445f78;
assign v144543c = decide_p & v14453f1 | !decide_p & v144543b;
assign bf1fa6 = hgrant2_p & bf1f59 | !hgrant2_p & !bf1fa5;
assign v144588f = hlock0 & v1445880 | !hlock0 & v144588e;
assign v16693a5 = decide_p & v16693a4 | !decide_p & v845542;
assign v151621d = jx2_p & v151621c | !jx2_p & v151621b;
assign d8078a = locked_p & d80789 | !locked_p & v845542;
assign bf1f5e = hbusreq5_p & bf1f5d | !hbusreq5_p & !bf1f5c;
assign v134d525 = hlock2 & v134d524 | !hlock2 & v134d51d;
assign v15167fe = hbusreq2 & v15167f6 | !hbusreq2 & v15167fd;
assign v16a169f = hmaster1_p & v16a169e | !hmaster1_p & v16a1d53;
assign d30685 = hbusreq2_p & v84555e | !hbusreq2_p & d30684;
assign d30707 = hmaster1_p & d306fd | !hmaster1_p & !d30706;
assign v16a194d = hmaster2_p & v16a1947 | !hmaster2_p & v16a194c;
assign v16a206a = hready & v16a2069 | !hready & v845542;
assign v134cf6d = hbusreq3_p & v134cf6c | !hbusreq3_p & v134d4c6;
assign v134ce7a = decide_p & v134d3ce | !decide_p & v134ce79;
assign v1214d60 = hmaster1_p & v12153ab | !hmaster1_p & v1214d5f;
assign v14466f2 = hmaster0_p & v144663a | !hmaster0_p & v1446440;
assign v1284d24 = hmaster0_p & v1284d0e | !hmaster0_p & v1284d23;
assign v1405b01 = hbusreq5_p & v1405afe | !hbusreq5_p & v1405b00;
assign v1552f70 = hmaster0_p & v845542 | !hmaster0_p & v1552f6f;
assign a65360 = hbusreq4_p & v10d3fd8 | !hbusreq4_p & v845542;
assign d30222 = hgrant5_p & d30220 | !hgrant5_p & d30221;
assign v12aeb22 = hgrant2_p & v12aeb1f | !hgrant2_p & v12aeb1b;
assign d2faf0 = hbusreq5_p & d3011c | !hbusreq5_p & !d2faef;
assign v14458c2 = hmaster1_p & v144639c | !hmaster1_p & v14458c1;
assign v15157bf = hgrant0_p & v15157be | !hgrant0_p & v845570;
assign v12160c9 = hmaster1_p & v1216099 | !hmaster1_p & v1216097;
assign v1405942 = jx1_p & v140582a | !jx1_p & v1405941;
assign a658e2 = hmaster2_p & a6627b | !hmaster2_p & a658e1;
assign v138945c = hbusreq2_p & v1389fe9 | !hbusreq2_p & v1389ff2;
assign v1214edc = hgrant5_p & v845547 | !hgrant5_p & v1214eda;
assign v1445b1f = hmaster1_p & v1445b01 | !hmaster1_p & v144591b;
assign v1215c94 = hgrant1_p & v1215c93 | !hgrant1_p & v12160fc;
assign v121614a = hlock0_p & v1216a61 | !hlock0_p & v1216149;
assign v12ad952 = decide_p & v12ad951 | !decide_p & v845542;
assign v1215379 = hbusreq0_p & v1215378 | !hbusreq0_p & v845542;
assign d2fc5e = hgrant1_p & d2fbe8 | !hgrant1_p & d2fc5d;
assign v16a1327 = hmaster2_p & v16a1326 | !hmaster2_p & !v845542;
assign v1445bf0 = hmaster1_p & v1446310 | !hmaster1_p & v1446329;
assign v1216319 = hlock5_p & v1216318 | !hlock5_p & v12162ef;
assign v12ad4d0 = hbusreq0_p & a65851 | !hbusreq0_p & v845542;
assign v13893b6 = hready_p & v1389394 | !hready_p & v13893b5;
assign v845588 = stateG3_2_p & v845542 | !stateG3_2_p & !v845542;
assign v121509a = hgrant5_p & v1215077 | !hgrant5_p & !v1215099;
assign v16a1ade = hbusreq5_p & v16a2079 | !hbusreq5_p & v16a1add;
assign v12153a7 = hmaster2_p & v12153a6 | !hmaster2_p & v845542;
assign v1215039 = hbusreq1_p & v1215035 | !hbusreq1_p & v1215038;
assign f2f37b = hgrant1_p & v845570 | !hgrant1_p & !f2f37a;
assign v138a2fd = hlock5_p & v138a2fc | !hlock5_p & v1668c21;
assign v1215cd6 = hmaster1_p & v1215cd5 | !hmaster1_p & v1215cc8;
assign v9f3194 = hburst1_p & v845542 | !hburst1_p & a67ea5;
assign v1215c66 = hbusreq0 & v1215c60 | !hbusreq0 & v1215c65;
assign v1445a52 = hbusreq1 & v14459c8 | !hbusreq1 & v14459cc;
assign v1446342 = hmaster1_p & v14465b7 | !hmaster1_p & v1446341;
assign v12ad000 = hgrant0_p & v12af9bc | !hgrant0_p & !v12acfff;
assign d2fee8 = hlock2_p & d2fee6 | !hlock2_p & d2fee7;
assign v1445995 = hlock4 & v144639c | !hlock4 & v1445994;
assign v12162c6 = hbusreq2_p & v12162c1 | !hbusreq2_p & v12162c5;
assign f2f283 = hgrant5_p & v845542 | !hgrant5_p & !f2f282;
assign v12ad4ec = hbusreq0 & v12ad4eb | !hbusreq0 & v845542;
assign v134d218 = hlock0 & v134d217 | !hlock0 & v134d216;
assign v1215d9b = hmaster0_p & v1215d9a | !hmaster0_p & !v1215d78;
assign v1668dc9 = hbusreq5_p & v1668dc7 | !hbusreq5_p & !v1668dc8;
assign v1445f6f = hbusreq2 & v1445f6d | !hbusreq2 & v1445f6e;
assign v134cd7a = hbusreq3 & v134cd78 | !hbusreq3 & v134cd79;
assign v1668cd5 = hbusreq0 & v1668cd2 | !hbusreq0 & v1668cd4;
assign v12165a9 = hbusreq5_p & v12165a8 | !hbusreq5_p & v845542;
assign d3081c = hbusreq5_p & d3081b | !hbusreq5_p & d3081a;
assign v1214e73 = hmaster0_p & v1214e72 | !hmaster0_p & v1214e0e;
assign v14463ed = hbusreq5_p & v14463ec | !hbusreq5_p & v14463bc;
assign d3074c = hmaster1_p & d3074b | !hmaster1_p & d3072c;
assign v144584d = hbusreq2_p & v1445844 | !hbusreq2_p & v144584c;
assign v1215714 = hlock4_p & v1215711 | !hlock4_p & v1215713;
assign v1552f68 = hlock0 & v15533a7 | !hlock0 & v1552f67;
assign v1445776 = hmaster2_p & v1445de5 | !hmaster2_p & v1446606;
assign d2fe7b = hbusreq4_p & d2fe7a | !hbusreq4_p & v845542;
assign v134d210 = hmaster1_p & v134d1e8 | !hmaster1_p & v134d20f;
assign v16a1d62 = hmaster0_p & v16a1d5f | !hmaster0_p & v16a1d61;
assign a662c1 = hmaster2_p & a662c0 | !hmaster2_p & !v845542;
assign d30245 = hgrant5_p & v845542 | !hgrant5_p & d301f5;
assign v1216330 = hbusreq2 & v1216327 | !hbusreq2 & v121632f;
assign v11ac6ca = hgrant3_p & v11ac67b | !hgrant3_p & v11ac6c9;
assign v16a224d = hgrant2_p & v16a205b | !hgrant2_p & v16a224c;
assign v16a13d5 = hbusreq2_p & v16a13d4 | !hbusreq2_p & !v16a1f9a;
assign v134ce68 = hlock2 & v134d3b5 | !hlock2 & v134ce64;
assign bf1faa = hgrant3_p & bf1f8c | !hgrant3_p & !bf1fa9;
assign v12ad534 = hlock2_p & v12ad52f | !hlock2_p & v12ad533;
assign v1216192 = hgrant5_p & v121601d | !hgrant5_p & v1216127;
assign f2f400 = hmaster1_p & f2f2e8 | !hmaster1_p & f2f2db;
assign v138a02d = hlock5_p & v138a02c | !hlock5_p & v845542;
assign v1215b95 = hmaster1_p & v1215b94 | !hmaster1_p & v845542;
assign v12ad583 = hmaster1_p & v12ad56b | !hmaster1_p & v12ad54f;
assign v14459e5 = hbusreq1_p & v144639c | !hbusreq1_p & v144660b;
assign d2f97c = hbusreq5_p & d2fea1 | !hbusreq5_p & !d2f97b;
assign v1515781 = hmaster2_p & v151577b | !hmaster2_p & v1515780;
assign v1216261 = hmaster2_p & v121625c | !hmaster2_p & v1216212;
assign v1445524 = hbusreq2 & v144551e | !hbusreq2 & v1445523;
assign v134ceda = hlock3 & v134d3ce | !hlock3 & v134ced9;
assign v1516988 = hbusreq3 & v1516982 | !hbusreq3 & v15167ee;
assign v1446132 = hbusreq2 & v1446130 | !hbusreq2 & v1446131;
assign v1445f20 = hgrant3_p & v1445e37 | !hgrant3_p & v1445f1f;
assign v12ad5ec = hbusreq0 & v12ad5eb | !hbusreq0 & v12afe63;
assign v1215cc0 = hbusreq5_p & v1215cbe | !hbusreq5_p & !v1215cbf;
assign v1552d85 = hgrant4_p & v1552d84 | !hgrant4_p & v845542;
assign v134d363 = hmaster0_p & v845542 | !hmaster0_p & v134d274;
assign v1215b9a = hmaster2_p & v12160ec | !hmaster2_p & !v1215b99;
assign d2fc36 = hbusreq5_p & d2fb79 | !hbusreq5_p & d2fc35;
assign v15156fd = hlock2_p & v15156fc | !hlock2_p & !v15156f6;
assign v121534b = hlock0_p & v1216a5a | !hlock0_p & v121534a;
assign v1389de0 = hlock5_p & v1389ddf | !hlock5_p & !v845542;
assign v16a19b4 = hbusreq2 & v16a19ae | !hbusreq2 & v16a19b3;
assign v12ae1f1 = hgrant1_p & v845542 | !hgrant1_p & v12ae1f0;
assign v151562c = stateA1_p & v845542 | !stateA1_p & !v151562b;
assign v134ce6b = hbusreq3 & v134ce69 | !hbusreq3 & v134ce6a;
assign a65b25 = hmaster0_p & v845542 | !hmaster0_p & !a6627c;
assign v1445b41 = hmaster1_p & v1445b40 | !hmaster1_p & v1445a32;
assign v1216030 = hmaster1_p & v121602f | !hmaster1_p & v845542;
assign v134d30b = hmaster2_p & v845542 | !hmaster2_p & v134d30a;
assign f2f23a = hgrant2_p & v845542 | !hgrant2_p & f2f239;
assign d30299 = hbusreq2_p & d30298 | !hbusreq2_p & !d30296;
assign v1216143 = hgrant1_p & v845542 | !hgrant1_p & v1216142;
assign v121504c = hlock0_p & v121504a | !hlock0_p & v121504b;
assign v1515755 = hgrant4_p & v1515746 | !hgrant4_p & v1515754;
assign v12ad5b5 = hbusreq0 & v12ad5b4 | !hbusreq0 & v12afe63;
assign d30836 = hbusreq5_p & d30835 | !hbusreq5_p & d30834;
assign v1215c49 = hbusreq2_p & v1215c37 | !hbusreq2_p & !v1215c48;
assign v12ad1b0 = decide_p & v12ad0ca | !decide_p & v12afe76;
assign v1215ba7 = hmaster2_p & v845542 | !hmaster2_p & v1215b97;
assign v1445b8c = hlock0 & v1445b8b | !hlock0 & v1445b8a;
assign v12ad13e = hbusreq2_p & v12ad13d | !hbusreq2_p & v12afe72;
assign v14460ac = hlock3 & v14460a1 | !hlock3 & v14460ab;
assign v1445392 = hgrant2_p & v144538d | !hgrant2_p & v1445391;
assign v1216a7b = hmaster0_p & v1216a7a | !hmaster0_p & v845542;
assign v151581a = hmaster0_p & v1515819 | !hmaster0_p & v151564f;
assign v16a16a1 = hbusreq2_p & v16a1e07 | !hbusreq2_p & v16a16a0;
assign d2feb0 = hbusreq4 & d30718 | !hbusreq4 & !v16693aa;
assign v1215054 = hmaster0_p & v1215041 | !hmaster0_p & v1215053;
assign v1284cca = hmaster2_p & v1284c8f | !hmaster2_p & !v1405845;
assign v12aeb70 = hmaster2_p & v845542 | !hmaster2_p & d30727;
assign v134d280 = hgrant5_p & v845542 | !hgrant5_p & v134d27f;
assign v1284d69 = jx0_p & v1284d68 | !jx0_p & v8b6f6a;
assign a6542b = hgrant5_p & a65424 | !hgrant5_p & !a653bc;
assign v1215ce7 = hgrant5_p & v845542 | !hgrant5_p & v1215c95;
assign v14460a6 = hmaster0_p & v1446404 | !hmaster0_p & v14460a5;
assign v12161f6 = hgrant2_p & v12161cd | !hgrant2_p & v12161f5;
assign v134d3d1 = hmaster1_p & v134d3d0 | !hmaster1_p & v845542;
assign v1405aca = hmaster2_p & v1405abb | !hmaster2_p & !v1405abf;
assign a658a8 = stateG3_2_p & v845542 | !stateG3_2_p & !afe156;
assign v1553231 = hgrant1_p & v845542 | !hgrant1_p & v1553230;
assign v144580e = hmaster0_p & v1445802 | !hmaster0_p & v1445ec3;
assign f2f42a = hbusreq5_p & f2f360 | !hbusreq5_p & !f2f429;
assign v151570a = hbusreq3 & v1515705 | !hbusreq3 & v1515709;
assign v1553930 = stateG3_0_p & v845586 | !stateG3_0_p & !acd334;
assign v1668c6d = hbusreq4 & a658c6 | !hbusreq4 & a658ca;
assign v1215774 = hmaster0_p & v1215b9a | !hmaster0_p & v1215773;
assign v10d401e = hgrant1_p & v10d4019 | !hgrant1_p & v10d401d;
assign d3083d = hmaster1_p & d3083c | !hmaster1_p & d30830;
assign v1214eb9 = hbusreq2 & v1214eb8 | !hbusreq2 & v845542;
assign d807be = hready_p & d807a4 | !hready_p & !d807bd;
assign v10d404f = hmaster0_p & v10d403d | !hmaster0_p & !v10d404e;
assign v16a2670 = hmaster2_p & v845559 | !hmaster2_p & !v845542;
assign v1668c63 = hbusreq1 & a658c6 | !hbusreq1 & a658ca;
assign v121571a = hbusreq1_p & v1215718 | !hbusreq1_p & v1215719;
assign v1216268 = hbusreq3 & v1216254 | !hbusreq3 & v1216267;
assign v16a16b1 = decide_p & v16a16b0 | !decide_p & v16a1e0e;
assign v134cd81 = hmaster1_p & v134d369 | !hmaster1_p & v134cd80;
assign v16695b0 = hlock3_p & v16695af | !hlock3_p & !v845542;
assign d300bc = hbusreq4_p & d300bb | !hbusreq4_p & v845542;
assign v16a12bf = hbusreq3 & v16a129c | !hbusreq3 & v16a12be;
assign v1445b7d = hmaster1_p & v1446313 | !hmaster1_p & v1445b7a;
assign v1445a25 = hbusreq4_p & v144639c | !hbusreq4_p & v1445a24;
assign v1445a79 = hbusreq5_p & v14459d1 | !hbusreq5_p & v1445a78;
assign v12aedde = decide_p & v12afa0f | !decide_p & v12afe76;
assign v12ad66e = stateA1_p & v12ad66d | !stateA1_p & a658a5;
assign v14460c8 = hbusreq3 & v14460c6 | !hbusreq3 & v14460c7;
assign d30762 = hlock2_p & d30761 | !hlock2_p & d3075e;
assign v1215b80 = hbusreq4_p & v121611e | !hbusreq4_p & v845542;
assign v1445456 = hbusreq2 & v1445445 | !hbusreq2 & v1445455;
assign v138a000 = hgrant5_p & v1389fff | !hgrant5_p & !v845542;
assign v134d45c = decide_p & v134d3fa | !decide_p & v134d45b;
assign v12152f3 = hbusreq2_p & v12152f1 | !hbusreq2_p & v12152f2;
assign v1389373 = decide_p & v1389372 | !decide_p & v845542;
assign v1515722 = hgrant4_p & v1515715 | !hgrant4_p & v1515721;
assign v1446670 = hgrant2_p & v1446669 | !hgrant2_p & v144666f;
assign v1445fb2 = hbusreq2_p & v1445faf | !hbusreq2_p & v1445fb1;
assign f2f2df = hmaster1_p & f2f2de | !hmaster1_p & f2f2db;
assign v1446067 = hbusreq0 & v1446060 | !hbusreq0 & v1446066;
assign v16a1b02 = hmaster1_p & v16a1b01 | !hmaster1_p & v16a2672;
assign v1445383 = hmaster1_p & v1445b3e | !hmaster1_p & v144591b;
assign v1445fe4 = hmaster0_p & v144639c | !hmaster0_p & v1445fe3;
assign d3064b = hmaster2_p & d30648 | !hmaster2_p & d3064a;
assign d2fc2a = decide_p & d2fc29 | !decide_p & v845570;
assign v138a3cf = hgrant5_p & v845542 | !hgrant5_p & v138a3ce;
assign a65470 = hmaster2_p & a658c7 | !hmaster2_p & !a6546d;
assign v1214d6c = hbusreq5 & v1214d5b | !hbusreq5 & v1214d6b;
assign v10d4016 = hmaster0_p & v10d3ff1 | !hmaster0_p & v10d3ff0;
assign v1668de2 = hgrant2_p & v1668da9 | !hgrant2_p & v1668dd3;
assign v14460de = hbusreq3 & v14460dc | !hbusreq3 & v14460dd;
assign d30284 = hmaster1_p & d30273 | !hmaster1_p & d30283;
assign v1445d9f = hbusreq4_p & v14463b3 | !hbusreq4_p & v14463bb;
assign v1216033 = hbusreq1 & v1216a8d | !hbusreq1 & v845542;
assign d30656 = hmaster2_p & v845542 | !hmaster2_p & d30655;
assign v12acff2 = hmaster1_p & v12acff1 | !hmaster1_p & v12ad4dd;
assign v1216a61 = hready & v1216a60 | !hready & a66295;
assign v1515700 = hbusreq3 & v15156f9 | !hbusreq3 & v15156ff;
assign v1445bc2 = hbusreq5_p & v144600c | !hbusreq5_p & v144647b;
assign a658f1 = hmaster2_p & a658b0 | !hmaster2_p & !a658cb;
assign v14460e5 = hmaster1_p & v14460e4 | !hmaster1_p & v845542;
assign d2fb4b = hbusreq3_p & d30165 | !hbusreq3_p & !d2fb4a;
assign v14466b6 = hgrant2_p & v144663c | !hgrant2_p & v14466b1;
assign d30815 = hgrant5_p & d306d0 | !hgrant5_p & d30797;
assign v1515812 = hmaster0_p & v1668dab | !hmaster0_p & v845542;
assign v144627f = hmaster1_p & v1446405 | !hmaster1_p & v144627e;
assign v1668d49 = hbusreq4_p & v1668d47 | !hbusreq4_p & !v1668d48;
assign f2f2e3 = hmaster2_p & f2f2c9 | !hmaster2_p & !f2f2e2;
assign v144631a = hmaster2_p & v14465ae | !hmaster2_p & v1446653;
assign v1445eef = hlock0 & v1445eee | !hlock0 & v1445eed;
assign v14058b6 = hmaster1_p & v14058b5 | !hmaster1_p & v140584d;
assign v155339a = hbusreq4_p & v1553217 | !hbusreq4_p & v1553399;
assign a65653 = hmaster1_p & a65635 | !hmaster1_p & a65652;
assign d3084f = hmaster2_p & d3084a | !hmaster2_p & !d3084e;
assign v138a448 = hbusreq5 & v138a447 | !hbusreq5 & v845542;
assign d2fafa = hgrant1_p & d2faf4 | !hgrant1_p & d2faec;
assign v1668c36 = decide_p & v1668c33 | !decide_p & v845542;
assign a6546a = hbusreq4_p & a65469 | !hbusreq4_p & !v845542;
assign v1446627 = hgrant4_p & v1446430 | !hgrant4_p & v1446626;
assign v1405af4 = hmaster0_p & v1405a8a | !hmaster0_p & v1405af3;
assign v1215346 = hbusreq0_p & v1215fec | !hbusreq0_p & v845542;
assign d807ad = hgrant2_p & d807a6 | !hgrant2_p & d807ac;
assign v12163a2 = hlock5_p & v12163a0 | !hlock5_p & !v12163a1;
assign v121631f = hmaster2_p & v1216ab9 | !hmaster2_p & v12162fc;
assign v15157f4 = hbusreq5_p & v15157f2 | !hbusreq5_p & !v15157f3;
assign v140585a = hmaster0_p & v1405855 | !hmaster0_p & v1405859;
assign v12af9c0 = hbusreq1_p & v12afe45 | !hbusreq1_p & v12af9bf;
assign v16a195f = hbusreq2 & v16a195d | !hbusreq2 & !v16a195e;
assign f2f376 = hgrant5_p & f2f363 | !hgrant5_p & f2f375;
assign v12af3aa = hbusreq0 & v12af3a5 | !hbusreq0 & v12af3a9;
assign v16a139d = hgrant3_p & v16a139a | !hgrant3_p & v16a139c;
assign v12ad4d7 = hmaster2_p & v12ad4d4 | !hmaster2_p & v12ad4d5;
assign d3091b = hlock2_p & d30919 | !hlock2_p & d3091a;
assign v1215407 = hmaster1_p & v12153f3 | !hmaster1_p & v12153ec;
assign v134d4e7 = hlock1 & v134d36d | !hlock1 & v134d4e6;
assign v1216082 = hmaster0_p & v1216081 | !hmaster0_p & v121605c;
assign v134d26d = hmaster1_p & v134d242 | !hmaster1_p & v134d23c;
assign a65891 = hmaster0_p & a65890 | !hmaster0_p & a6587e;
assign v16a1a8f = hready_p & v16a1a8d | !hready_p & v16a1a8e;
assign v1214ed1 = hgrant5_p & v845547 | !hgrant5_p & v1214ecf;
assign v14461d6 = hlock2 & v14461cd | !hlock2 & v14461d5;
assign v1445dbb = hbusreq2_p & v1445da5 | !hbusreq2_p & v1445dba;
assign a65676 = hbusreq5_p & a65434 | !hbusreq5_p & a65674;
assign v12150ae = hbusreq2_p & v12150a8 | !hbusreq2_p & v12150ad;
assign v1284c97 = decide_p & v1284c96 | !decide_p & v1284c95;
assign v12ad4fe = hbusreq0 & v12ad4fd | !hbusreq0 & v845542;
assign v14457ab = hbusreq2 & v14457a9 | !hbusreq2 & v14457aa;
assign v1405af7 = hgrant5_p & v1405a96 | !hgrant5_p & v1405af6;
assign v1445bed = hmaster0_p & v1446310 | !hmaster0_p & v14465b7;
assign v1405ae5 = hlock4_p & v1405a88 | !hlock4_p & !v845542;
assign v144577c = hmaster1_p & v144577b | !hmaster1_p & v1445e07;
assign d300dd = hgrant4_p & v845542 | !hgrant4_p & d300dc;
assign d2f9a9 = hmaster0_p & d2f99f | !hmaster0_p & d2f9a8;
assign v121625e = hgrant5_p & v12160d5 | !hgrant5_p & v121625d;
assign v1668d86 = hmaster2_p & v1668d83 | !hmaster2_p & v1668d85;
assign v144625b = hbusreq2 & v1446259 | !hbusreq2 & v144625a;
assign v1446010 = hbusreq5_p & v144600c | !hbusreq5_p & v144600f;
assign d2fe90 = hmaster1_p & d2fe8f | !hmaster1_p & d2fe8c;
assign v1215c8e = hgrant5_p & v1668da6 | !hgrant5_p & v1215c8d;
assign v1405892 = hmaster2_p & v1405891 | !hmaster2_p & v14463b1;
assign v134d4bb = hready_p & v134d34f | !hready_p & v134d4ba;
assign v1445d8e = hmaster2_p & v144639c | !hmaster2_p & v1445f97;
assign v1668cdd = hmastlock_p & v1668cdc | !hmastlock_p & v845542;
assign v1445df9 = hbusreq0 & v1445df4 | !hbusreq0 & v1445df8;
assign v1284d0c = hgrant1_p & v140587c | !hgrant1_p & v1284d0b;
assign d302e0 = hbusreq5_p & d302df | !hbusreq5_p & d30656;
assign v134ce59 = hlock2 & v134ce48 | !hlock2 & v134ce58;
assign v1284ce0 = hmaster1_p & v1284cc9 | !hmaster1_p & !v1284cdf;
assign v1446210 = hbusreq5_p & v14463a4 | !hbusreq5_p & v144620f;
assign v134d209 = hmaster1_p & v134d1e8 | !hmaster1_p & v134d208;
assign v12150c2 = hbusreq4 & v1216ab9 | !hbusreq4 & v12150c1;
assign v1214c6a = hlock0_p & v1216551 | !hlock0_p & v1214c69;
assign v12166db = hlock0_p & v12164d3 | !hlock0_p & v12166da;
assign v12160f5 = hbusreq1 & v12160f4 | !hbusreq1 & v845542;
assign v12153f9 = hmaster0_p & v12153f3 | !hmaster0_p & v12153d4;
assign d2fc1a = decide_p & d2fc19 | !decide_p & v845570;
assign v12152fd = hgrant2_p & v1215787 | !hgrant2_p & v12152fc;
assign v14459c4 = hbusreq4 & v14465ad | !hbusreq4 & v14459c3;
assign v12153e2 = hlock0_p & v12153d1 | !hlock0_p & !v845542;
assign v1668d91 = hmaster2_p & a65861 | !hmaster2_p & !v1668d4f;
assign a6568a = hmaster1_p & a6548f | !hmaster1_p & a658e5;
assign v1445ea4 = hbusreq1 & v1445ea2 | !hbusreq1 & v1445ea3;
assign v12ad279 = decide_p & v12ad1fd | !decide_p & v12afe76;
assign v1215d3b = hmaster1_p & v1215d31 | !hmaster1_p & v1215d3a;
assign v1284d02 = hmaster1_p & v1284d01 | !hmaster1_p & v140584d;
assign v151566f = stateA1_p & v151566e | !stateA1_p & a658a5;
assign v1552f54 = hbusreq4_p & v1552f53 | !hbusreq4_p & v1553217;
assign d807a5 = hmaster0_p & d80762 | !hmaster0_p & d80761;
assign v1216302 = hbusreq0 & v1216adb | !hbusreq0 & v1216301;
assign v1214d38 = hbusreq2_p & v1214d36 | !hbusreq2_p & v1214d37;
assign v110b6cc = stateG3_2_p & v88d3e4 | !stateG3_2_p & v9f3194;
assign v121539b = hbusreq1 & v845547 | !hbusreq1 & v1215364;
assign v1516102 = hmaster1_p & v1516101 | !hmaster1_p & v845542;
assign f2f3fb = hmaster0_p & f2f2e8 | !hmaster0_p & f2f2dd;
assign v1214c49 = hlock0_p & v1216528 | !hlock0_p & v845542;
assign v12160e0 = hmaster0_p & v12160da | !hmaster0_p & v12160df;
assign v1446244 = hbusreq2 & v144623f | !hbusreq2 & v1446243;
assign a6564a = hgrant4_p & a662a9 | !hgrant4_p & !a653de;
assign d80733 = locked_p & d80732 | !locked_p & !v845542;
assign v1668c9c = hmaster0_p & v1668c9b | !hmaster0_p & !v1668c71;
assign v12165b3 = hbusreq5 & v12165b2 | !hbusreq5 & v845542;
assign v1405b20 = hgrant5_p & v1405b17 | !hgrant5_p & !v1405b1f;
assign v15156b1 = hmaster0_p & v1668cc9 | !hmaster0_p & v15156b0;
assign v1445786 = hbusreq2_p & v1445783 | !hbusreq2_p & v1445785;
assign d300d2 = hbusreq5_p & d300d1 | !hbusreq5_p & !d300d0;
assign f2f415 = hready_p & f2f3ee | !hready_p & f2f414;
assign d301ea = hbusreq1_p & d301e8 | !hbusreq1_p & d301e9;
assign v1515657 = hlock1_p & v1515655 | !hlock1_p & v1515656;
assign v134d4b4 = hlock2 & v134d3b5 | !hlock2 & v134d4b0;
assign v12161d7 = hbusreq1 & v1216594 | !hbusreq1 & !v845542;
assign v1668d67 = hburst1_p & v845542 | !hburst1_p & v1668d66;
assign v144628f = hlock0 & v144628e | !hlock0 & v144628d;
assign v12164d2 = locked_p & v12164d1 | !locked_p & !v845542;
assign v9109e4 = hmaster0_p & v845542 | !hmaster0_p & v845568;
assign v121621e = hbusreq1 & v12166e9 | !hbusreq1 & v845542;
assign v15530a4 = hlock5 & v155341e | !hlock5 & v1553094;
assign v14465f4 = hbusreq1 & v14465f0 | !hbusreq1 & v14465f3;
assign v1214dce = hmaster1_p & v1214dcd | !hmaster1_p & v1216a5a;
assign v12ad4e2 = hmaster1_p & v12ad4e1 | !hmaster1_p & v12ad4dd;
assign v16a13c7 = hmaster0_p & v16a2674 | !hmaster0_p & v16a2669;
assign v1284cf9 = hgrant4_p & v140584b | !hgrant4_p & !v1284cf8;
assign v1668d9c = hbusreq5_p & v1668d99 | !hbusreq5_p & v1668d9b;
assign v1216298 = hgrant2_p & v12161a8 | !hgrant2_p & v1216297;
assign v1216043 = hmaster0_p & v1216035 | !hmaster0_p & f2f2a8;
assign v16a13c4 = hmaster2_p & v16a13a7 | !hmaster2_p & !v845542;
assign v144645a = hbusreq3 & v1446457 | !hbusreq3 & v1446459;
assign v134cd71 = hlock0 & v134cd70 | !hlock0 & v134cd6f;
assign v16a1a80 = hgrant2_p & v845542 | !hgrant2_p & !v16a1a7d;
assign d301ae = hmaster1_p & d3018e | !hmaster1_p & !d3019e;
assign v16a1980 = hmaster1_p & v16a197c | !hmaster1_p & v16a197f;
assign v12167a0 = hready_p & v1216796 | !hready_p & v121679f;
assign v1214e1a = hmaster0_p & v121639e | !hmaster0_p & v845542;
assign v14eb679 = hbusreq3_p & v845542 | !hbusreq3_p & v845578;
assign a6568b = hbusreq2_p & a65688 | !hbusreq2_p & a6568a;
assign v1284cec = hmaster2_p & v14463b1 | !hmaster2_p & !v1284ceb;
assign a65493 = hmaster0_p & a658f1 | !hmaster0_p & a658b7;
assign d80785 = hgrant2_p & d80769 | !hgrant2_p & d80784;
assign v1515767 = hgrant1_p & v1515761 | !hgrant1_p & v1515766;
assign v1446258 = hbusreq2_p & v1446254 | !hbusreq2_p & v1446257;
assign v140593c = decide_p & v1405933 | !decide_p & v140593b;
assign d2fbe0 = hgrant1_p & d2fbdf | !hgrant1_p & d2fbd4;
assign v121611e = hbusreq4 & v1215ff8 | !hbusreq4 & v845542;
assign a65924 = hmaster1_p & a658ee | !hmaster1_p & !a65916;
assign v138a485 = hgrant2_p & v138a484 | !hgrant2_p & v138a47f;
assign v144599d = hgrant1_p & v14458d2 | !hgrant1_p & v144599c;
assign d30785 = hgrant0_p & d30784 | !hgrant0_p & v845542;
assign v12ad4ce = hbusreq0 & v12ad4cd | !hbusreq0 & v845542;
assign v16695bd = hready_p & v16695b1 | !hready_p & !v16695bc;
assign v1445ee5 = hbusreq2 & v1445ed1 | !hbusreq2 & v1445ee4;
assign v1216135 = hbusreq0 & v1216129 | !hbusreq0 & v1216134;
assign f2f405 = hmaster1_p & f2f2dd | !hmaster1_p & !f2f330;
assign v1214ce9 = hlock0_p & v845542 | !hlock0_p & v1214ce8;
assign v138a3a4 = hmaster1_p & v138a3a3 | !hmaster1_p & v138a341;
assign v1446643 = hgrant5_p & v144643b | !hgrant5_p & v1446642;
assign v10d405b = hgrant2_p & v10d4054 | !hgrant2_p & !v10d405a;
assign v12162d4 = hgrant2_p & v12162c8 | !hgrant2_p & v12162d3;
assign v1405adf = hgrant5_p & v1405a8d | !hgrant5_p & v1405add;
assign f2f3d6 = hgrant5_p & v84554c | !hgrant5_p & f2f3a4;
assign v1216581 = hbusreq2_p & v121657f | !hbusreq2_p & v1216580;
assign d8075f = hmastlock_p & d8075e | !hmastlock_p & !v845542;
assign v121609a = hmaster0_p & v1216093 | !hmaster0_p & v1216099;
assign v14459d7 = hbusreq0_p & v845542 | !hbusreq0_p & !v14463b1;
assign v15155e6 = hbusreq0_p & d305ef | !hbusreq0_p & v16693aa;
assign v1445f9a = hbusreq0 & v1445f96 | !hbusreq0 & v1445f99;
assign v144600e = hmaster2_p & v144600d | !hmaster2_p & v845542;
assign v1215b8f = hbusreq4 & v1216568 | !hbusreq4 & v1215b8e;
assign d30264 = hbusreq5 & d3023c | !hbusreq5 & d30263;
assign v1216294 = hmaster1_p & v12161a1 | !hmaster1_p & v121619c;
assign v16a1abb = hready_p & v16a20a6 | !hready_p & !v16a1aba;
assign d2fbab = hlock2_p & d2fbaa | !hlock2_p & d2fba7;
assign v1215ca8 = hgrant5_p & v845542 | !hgrant5_p & !v1215ca6;
assign v1668d79 = hlock0_p & v1668d25 | !hlock0_p & v1668d78;
assign f2f3a2 = hgrant5_p & f2f3a1 | !hgrant5_p & !f2f39f;
assign v1215db0 = hgrant3_p & v1215bd9 | !hgrant3_p & v1215daf;
assign v14463a6 = hmaster2_p & v144639e | !hmaster2_p & v14463a5;
assign v1216187 = hlock2_p & v1216183 | !hlock2_p & v1216186;
assign v1215014 = hmaster2_p & v845542 | !hmaster2_p & v1215013;
assign v1405889 = hbusreq1_p & v1405888 | !hbusreq1_p & v140583c;
assign d3022e = hmaster1_p & d3022d | !hmaster1_p & d30218;
assign v12163a9 = hmaster0_p & v12163a3 | !hmaster0_p & v12163a8;
assign v121655e = hgrant4_p & v121655d | !hgrant4_p & v845542;
assign v1445536 = hlock5 & v14454fa | !hlock5 & v1445535;
assign v144647b = hgrant5_p & v1446477 | !hgrant5_p & v144647a;
assign v1215418 = hmaster1_p & v12153f9 | !hmaster1_p & v121540f;
assign v144617d = hmaster1_p & v144617c | !hmaster1_p & v1445fde;
assign f2f35d = hbusreq0 & f2f352 | !hbusreq0 & f2f35c;
assign d300c7 = hgrant5_p & d2fe9b | !hgrant5_p & !d300c5;
assign v134cebd = hbusreq3 & v134cebb | !hbusreq3 & v134cebc;
assign v1552d53 = hmaster0_p & v845542 | !hmaster0_p & v1552d52;
assign a653e8 = hmaster1_p & a6538f | !hmaster1_p & a653e7;
assign v10d409e = hbusreq2_p & v10d409b | !hbusreq2_p & v10d409d;
assign a65b38 = hbusreq3_p & a65b23 | !hbusreq3_p & a65b32;
assign v16a206e = hgrant4_p & v845559 | !hgrant4_p & v845542;
assign d807bc = hready_p & d807b8 | !hready_p & !d807bb;
assign a65b31 = hready_p & a65b2f | !hready_p & a65b30;
assign d30658 = hgrant4_p & a66297 | !hgrant4_p & a65382;
assign v14058df = hgrant5_p & v140584f | !hgrant5_p & v14058de;
assign a65456 = decide_p & a65929 | !decide_p & a662a2;
assign v134d21e = hbusreq2 & v134d20e | !hbusreq2 & v134d21d;
assign v10d40a6 = hmaster1_p & v10d40a5 | !hmaster1_p & v10d3ffb;
assign v10d4274 = hgrant5_p & v10d3ffd | !hgrant5_p & !v10d4272;
assign v1445e1f = hbusreq2_p & v1445e1c | !hbusreq2_p & v1445e1e;
assign d2f9cc = hmaster1_p & d2fef8 | !hmaster1_p & d2f9cb;
assign v12af3ad = decide_p & v12af3ac | !decide_p & v845542;
assign v1214ce0 = hbusreq0 & v1214cdf | !hbusreq0 & v845542;
assign v15156ae = hgrant1_p & v15156ad | !hgrant1_p & v1668cd3;
assign d2fb06 = hgrant5_p & d2f97b | !hgrant5_p & !d2fb05;
assign a6585b = hmastlock_p & a65859 | !hmastlock_p & v845542;
assign v11e5981 = hready_p & v11e5980 | !hready_p & !v845542;
assign v1445bd1 = hmaster0_p & v1446643 | !hmaster0_p & v14465b7;
assign v121536e = hmaster1_p & v121536d | !hmaster1_p & v121536b;
assign d2fc4a = hlock0_p & v845542 | !hlock0_p & !d2fc49;
assign v1445d87 = hlock1 & v14463b9 | !hlock1 & v1445d80;
assign v11e5957 = hgrant0_p & v11e5956 | !hgrant0_p & !v845542;
assign v16a1e05 = hready_p & v845555 | !hready_p & v16a1e04;
assign v1445e7b = hbusreq1_p & v14465b2 | !hbusreq1_p & v1445e68;
assign d2fb2b = hmaster1_p & d2fb1f | !hmaster1_p & d2fb2a;
assign v1216025 = hlock1_p & v1216024 | !hlock1_p & !v845542;
assign v15167b6 = hmaster0_p & v845542 | !hmaster0_p & v1668c2a;
assign v138a323 = busreq_p & v138a322 | !busreq_p & a658a5;
assign v14458b1 = hmaster0_p & v144639c | !hmaster0_p & v14458a2;
assign v1446610 = hmaster2_p & v1446609 | !hmaster2_p & v144660f;
assign d2faf3 = hbusreq1 & d2f96d | !hbusreq1 & d30660;
assign v14463ff = hlock3 & v14463d1 | !hlock3 & v14463fe;
assign d301ba = hready_p & d308d5 | !hready_p & d301b9;
assign v1445821 = hmaster1_p & v1445eba | !hmaster1_p & v1445ef0;
assign v1215749 = hgrant5_p & v1215743 | !hgrant5_p & v1215748;
assign v121501d = hgrant5_p & v1215bac | !hgrant5_p & v121501c;
assign v1216ad4 = hbusreq4 & v1216aad | !hbusreq4 & v1216ad3;
assign v16a1deb = hmaster0_p & v16a2243 | !hmaster0_p & v16a2234;
assign f2f22f = hbusreq1_p & f2f22e | !hbusreq1_p & !v845542;
assign v121615b = hgrant4_p & v1216137 | !hgrant4_p & v845542;
assign v1214d3d = hmaster0_p & v1214cdc | !hmaster0_p & v121538a;
assign d307c6 = hbusreq4 & d307ac | !hbusreq4 & v845542;
assign v134cdcd = hready_p & v134d3e5 | !hready_p & v134cdcc;
assign a662a2 = hgrant2_p & v845542 | !hgrant2_p & a662a1;
assign d30799 = hgrant5_p & d306fd | !hgrant5_p & !d30797;
assign v1445fcc = hbusreq1_p & v1446439 | !hbusreq1_p & v1446406;
assign d2fc3b = hmaster0_p & d2fc34 | !hmaster0_p & d2fc3a;
assign v134d23e = hmaster1_p & v134d20b | !hmaster1_p & v134d23c;
assign v14457d8 = hmaster0_p & v14457d7 | !hmaster0_p & v144639c;
assign d30207 = hbusreq1 & d30703 | !hbusreq1 & v845542;
assign v134cd6a = hlock0 & v134d38b | !hlock0 & v134cd69;
assign v1215bcd = hbusreq2 & v1215bc6 | !hbusreq2 & v1215bcc;
assign d3027b = hgrant5_p & v845542 | !hgrant5_p & !d3065e;
assign v1214d5e = hbusreq0 & v1214d5d | !hbusreq0 & v845542;
assign v16a141c = decide_p & v16a13d8 | !decide_p & !v16a141b;
assign d2fc7b = hbusreq5 & d2fc72 | !hbusreq5 & d2fc7a;
assign v1405913 = hbusreq4_p & v1405860 | !hbusreq4_p & v1405912;
assign v1445502 = hmaster2_p & v1445412 | !hmaster2_p & v144665b;
assign v134d295 = hmaster1_p & v134d280 | !hmaster1_p & v134d294;
assign d2fbc3 = hlock3_p & d2fbaf | !hlock3_p & d2fbc2;
assign v16a1841 = hmaster1_p & v16a1840 | !hmaster1_p & v16a2672;
assign v1445f94 = hbusreq1 & v14463b3 | !hbusreq1 & v14463e7;
assign v121601b = hbusreq3 & v1216011 | !hbusreq3 & v121601a;
assign v15161fe = hbusreq2 & v15161cf | !hbusreq2 & v15161fd;
assign v144600a = decide_p & v1445fca | !decide_p & v1446009;
assign v121545c = hbusreq5 & v121544c | !hbusreq5 & v121545b;
assign d2fbbd = hbusreq2_p & d2fbbc | !hbusreq2_p & d2fbbb;
assign v12ad4c2 = hbusreq0 & v12ad8e6 | !hbusreq0 & v12ad4c1;
assign v12161b2 = hgrant2_p & v12161a7 | !hgrant2_p & v12161b1;
assign v15157c1 = hgrant1_p & f2f281 | !hgrant1_p & v15157c0;
assign v11e5969 = hmaster2_p & v11e5965 | !hmaster2_p & v11e5968;
assign v12ad52b = hbusreq2_p & v12ad526 | !hbusreq2_p & v12ad52a;
assign v16a1322 = hbusreq0_p & v16a1321 | !hbusreq0_p & !v845542;
assign v1214ecc = hgrant5_p & v845547 | !hgrant5_p & v1216539;
assign v1214c63 = hgrant5_p & v1215368 | !hgrant5_p & v1214c62;
assign v1405b56 = hgrant2_p & v1405b3e | !hgrant2_p & v1405b55;
assign v1668c47 = hlock3_p & v1668c46 | !hlock3_p & !v845542;
assign f2ec25 = hmaster1_p & v845542 | !hmaster1_p & f2ec24;
assign v1214bd6 = hlock2_p & v1214bd4 | !hlock2_p & v1214bd5;
assign v1445795 = hmaster1_p & v1445791 | !hmaster1_p & v1445e07;
assign v1445a7a = hbusreq0 & v1445a79 | !hbusreq0 & v14459f0;
assign d80791 = hbusreq5_p & d8078e | !hbusreq5_p & !d80790;
assign v1214d9c = hmaster0_p & v121538a | !hmaster0_p & v121537b;
assign d807b4 = hready_p & d807a4 | !hready_p & !d807b3;
assign v1405a9c = hmaster1_p & v1405a9b | !hmaster1_p & !v1405a94;
assign v144618f = hmaster1_p & v1446092 | !hmaster1_p & v1446073;
assign v12147ea = decide_p & v1214f1b | !decide_p & v12147e9;
assign v10d4078 = hgrant4_p & v10d3fe7 | !hgrant4_p & !v10d4077;
assign v1446629 = hbusreq1 & v1446627 | !hbusreq1 & v1446628;
assign v1552fd5 = decide_p & v155342e | !decide_p & v1552f8a;
assign v12ad5b4 = hbusreq5_p & v12ad5b2 | !hbusreq5_p & v12ad5b3;
assign v10d42b5 = hmaster1_p & v10d42b4 | !hmaster1_p & v10d407c;
assign v1445a16 = hbusreq4_p & v14465b1 | !hbusreq4_p & v14459ca;
assign v1445ac4 = hmaster0_p & v14458aa | !hmaster0_p & v14458a6;
assign v1405b17 = hmaster2_p & v1405a88 | !hmaster2_p & !v1405ac0;
assign v144640f = hbusreq1 & v144640d | !hbusreq1 & v144640e;
assign v1445e98 = hlock0_p & v144639c | !hlock0_p & v1445e97;
assign v1215cf0 = hbusreq5_p & v1215cef | !hbusreq5_p & !v1215cab;
assign v12ad27c = hbusreq3_p & v12ad1b3 | !hbusreq3_p & v12ad27b;
assign v134d4f1 = hgrant1_p & v134d4f0 | !hgrant1_p & v845542;
assign d3010f = hmaster1_p & d300d3 | !hmaster1_p & d3010e;
assign v15155f7 = hbusreq0 & v845570 | !hbusreq0 & v845542;
assign v16a1d28 = hbusreq2 & v16a1d26 | !hbusreq2 & v16a1d27;
assign v1445efd = hgrant2_p & v1445efc | !hgrant2_p & v1445ef8;
assign v1445e8f = hbusreq1 & v1445e8b | !hbusreq1 & v1445e8e;
assign a65363 = hlock0_p & a65851 | !hlock0_p & v10d3fd8;
assign v1405a7d = hlock0_p & v845542 | !hlock0_p & v845548;
assign v151578d = hburst1 & v151578c | !hburst1 & v1515672;
assign v1445907 = hmaster2_p & v14458d2 | !hmaster2_p & v1445906;
assign v1445494 = hbusreq2_p & v1445493 | !hbusreq2_p & v1445bba;
assign v144661d = hgrant4_p & v1446430 | !hgrant4_p & v144661c;
assign v16a2097 = hgrant2_p & v845542 | !hgrant2_p & v16a2096;
assign v12ad01a = hbusreq2_p & v12acff5 | !hbusreq2_p & v12ad019;
assign v121572a = hgrant1_p & v121570e | !hgrant1_p & v1215729;
assign v121541a = hlock2_p & v1215418 | !hlock2_p & v1215419;
assign d2fbe7 = hlock1_p & d2fbe6 | !hlock1_p & v84554a;
assign f2f425 = hgrant5_p & f2f3a1 | !hgrant5_p & !f2f424;
assign v1216259 = hbusreq2_p & v1216256 | !hbusreq2_p & v1216258;
assign v16a13ec = hgrant5_p & v845542 | !hgrant5_p & !v16a2081;
assign d2fe7e = hmaster2_p & d2fe7b | !hmaster2_p & d2fe7d;
assign v144586d = hlock0_p & v14463a0 | !hlock0_p & v144586c;
assign v1216182 = hmaster0_p & v845542 | !hmaster0_p & v1216018;
assign a662cb = hgrant5_p & v845542 | !hgrant5_p & a662ca;
assign v1445bb0 = hbusreq5_p & v1445f85 | !hbusreq5_p & v1445baf;
assign v1214c42 = hmaster0_p & v121534d | !hmaster0_p & v1215349;
assign v138a308 = hlock5_p & v1515628 | !hlock5_p & v1515631;
assign v12af9da = hbusreq2_p & v12afe68 | !hbusreq2_p & v12af9d9;
assign v16a1d74 = hbusreq2 & v16a1d70 | !hbusreq2 & !v16a1d73;
assign v1668c50 = hmaster1_p & v1668c4f | !hmaster1_p & v845542;
assign v14459e0 = hmaster2_p & v14459df | !hmaster2_p & v14459cf;
assign v1216216 = hbusreq1 & v12166d8 | !hbusreq1 & v845542;
assign v1445406 = hbusreq5_p & v1446473 | !hbusreq5_p & v1445405;
assign v16a1e0b = hgrant2_p & v845542 | !hgrant2_p & !v16a1e0a;
assign v12af1b9 = hbusreq1_p & v12afda1 | !hbusreq1_p & v12af984;
assign v1405adc = hgrant1_p & v1405adb | !hgrant1_p & !v1405a8c;
assign v1668dac = hmaster0_p & v845542 | !hmaster0_p & v1668dab;
assign v1445b23 = hbusreq2_p & v1445b1f | !hbusreq2_p & v1445b22;
assign v12ad600 = hgrant5_p & v845542 | !hgrant5_p & !v12ad5b1;
assign d305e0 = hlock5_p & v845542 | !hlock5_p & d305df;
assign f2f40f = hmaster1_p & f2f2e8 | !hmaster1_p & !f2f330;
assign v12af3a5 = hmaster2_p & v845542 | !hmaster2_p & !v12af3a4;
assign v12157a9 = hmastlock_p & a65366 | !hmastlock_p & v845542;
assign v1553306 = decide_p & v15532bf | !decide_p & v15532cd;
assign v1215b78 = hbusreq4 & v1216a61 | !hbusreq4 & v1215b77;
assign v12153d4 = hmaster2_p & v12153ce | !hmaster2_p & v12153d3;
assign v10d4049 = hgrant4_p & v10d4045 | !hgrant4_p & !v10d4048;
assign v1445aa6 = hbusreq2_p & v1445a9d | !hbusreq2_p & v1445aa5;
assign v14453a5 = hmaster1_p & v1445b33 | !hmaster1_p & v1445a9b;
assign v15155f4 = hlock2_p & v15155f3 | !hlock2_p & !v845542;
assign f2f2d1 = hbusreq5_p & f2f2cd | !hbusreq5_p & !f2f2d0;
assign v121539e = hmaster2_p & v1215394 | !hmaster2_p & v121539d;
assign v1214c40 = decide_p & v1214c27 | !decide_p & v1214c3f;
assign v1215790 = hgrant5_p & v121578f | !hgrant5_p & v121573e;
assign a658d0 = hmaster2_p & a658c7 | !hmaster2_p & !a658ce;
assign v151563c = hlock2_p & v151563b | !hlock2_p & !v845542;
assign d301f8 = hbusreq1_p & v845542 | !hbusreq1_p & d307bb;
assign v138a392 = hbusreq5 & v138a366 | !hbusreq5 & !v138a391;
assign v14453c7 = hbusreq3_p & v1445aaf | !hbusreq3_p & v14453c6;
assign d80771 = hlock1_p & d80733 | !hlock1_p & !v845542;
assign a65389 = hgrant1_p & a65362 | !hgrant1_p & !a65387;
assign a65685 = hmaster1_p & a658e8 | !hmaster1_p & a658e5;
assign a658d7 = hbusreq4_p & a658d6 | !hbusreq4_p & v845542;
assign v1214c07 = hmaster0_p & v1214bb7 | !hmaster0_p & v12153ab;
assign v1214d1a = hmaster2_p & v1214d12 | !hmaster2_p & !v1214c31;
assign f2f351 = hgrant5_p & f2f350 | !hgrant5_p & !f2f34d;
assign v1668d14 = hready_p & v1668c5b | !hready_p & !v1668d13;
assign v16a1e24 = hmaster1_p & v16a1e23 | !hmaster1_p & !v16a2672;
assign v1445b0e = hmaster1_p & v1445ae5 | !hmaster1_p & v144591b;
assign v1445396 = hbusreq2_p & v1445392 | !hbusreq2_p & v1445395;
assign d2fb82 = hbusreq2_p & d2fb81 | !hbusreq2_p & d2fb80;
assign v1214db1 = hmaster0_p & v1214c3c | !hmaster0_p & v1214d14;
assign v1216092 = hbusreq1_p & v1216091 | !hbusreq1_p & v845542;
assign v11e5979 = hgrant1_p & v845542 | !hgrant1_p & v11e5978;
assign v1214f00 = hbusreq0 & v1216530 | !hbusreq0 & v121653a;
assign v12164da = hmaster2_p & v845542 | !hmaster2_p & v12164d9;
assign v1446336 = hbusreq2_p & v1446301 | !hbusreq2_p & v1446335;
assign v1214800 = hbusreq2 & v12147ff | !hbusreq2 & v12164e7;
assign v1214bb8 = hmaster0_p & v1215396 | !hmaster0_p & v1214bb7;
assign d30679 = hbusreq2 & d30671 | !hbusreq2 & d30678;
assign v1216160 = hbusreq1_p & v121615f | !hbusreq1_p & v845542;
assign v155341b = hlock2 & v15533b8 | !hlock2 & v155341a;
assign v1446200 = hbusreq3 & v14461fe | !hbusreq3 & v14461ff;
assign v1214c4b = hgrant4_p & v1214c48 | !hgrant4_p & v1214c4a;
assign v12ad00e = hbusreq0 & v12ad00d | !hbusreq0 & v12afa0a;
assign a656b9 = hbusreq3_p & a65458 | !hbusreq3_p & a656b8;
assign v134d449 = hbusreq3 & v134d447 | !hbusreq3 & v134d448;
assign v1668d1f = hmaster1_p & v1668d17 | !hmaster1_p & v1668d1e;
assign v1216b00 = hmaster2_p & v1216aa9 | !hmaster2_p & v1216abb;
assign v138980d = hmaster2_p & v1515ae7 | !hmaster2_p & a6587e;
assign v144606e = hgrant1_p & v1445fdb | !hgrant1_p & v144606d;
assign v1445de7 = hmaster2_p & v1445de5 | !hmaster2_p & v1446403;
assign v155309b = hgrant2_p & v1553380 | !hgrant2_p & v155309a;
assign a653dc = hlock0_p & a6588d | !hlock0_p & !a653da;
assign v1215ce6 = hbusreq0 & v1215ce3 | !hbusreq0 & v1215ce5;
assign v151581d = hbusreq2_p & v151581c | !hbusreq2_p & v845542;
assign v14460b3 = hbusreq5_p & v1446042 | !hbusreq5_p & v14460b2;
assign v14058e5 = hmaster0_p & v140587e | !hmaster0_p & v140587d;
assign v138a47f = hmaster1_p & v138a3ec | !hmaster1_p & v138a3e0;
assign a65636 = hbusreq1_p & a65376 | !hbusreq1_p & a65621;
assign v15156db = hmaster1_p & v1515650 | !hmaster1_p & !v15156da;
assign v1552d93 = hmaster1_p & v1552d92 | !hmaster1_p & v845542;
assign a653c2 = hbusreq1 & a6586c | !hbusreq1 & a6587e;
assign v1214d83 = hgrant2_p & v1214d76 | !hgrant2_p & v1214d82;
assign d307dc = hmaster2_p & d307cd | !hmaster2_p & d307db;
assign v12af985 = hbusreq1_p & v12afda3 | !hbusreq1_p & v12af984;
assign v16a2058 = hmaster1_p & v845568 | !hmaster1_p & !v16a2672;
assign v140591e = hmaster1_p & v140591d | !hmaster1_p & v140584d;
assign v12157a2 = hgrant5_p & v845542 | !hgrant5_p & v1215776;
assign v1215799 = hgrant5_p & v1215791 | !hgrant5_p & v1215751;
assign d3012b = hgrant2_p & d3012a | !hgrant2_p & d3010f;
assign v134d37a = hbusreq5_p & v134d376 | !hbusreq5_p & v134d379;
assign v1445b29 = hlock5 & v1445b0d | !hlock5 & v1445b28;
assign v1515621 = hbusreq2_p & v1515620 | !hbusreq2_p & v845542;
assign d30831 = hmaster1_p & d3081d | !hmaster1_p & d30830;
assign v1445de0 = hlock5 & v1445dc6 | !hlock5 & v1445dde;
assign f2f2c9 = hbusreq1_p & f2f2c8 | !hbusreq1_p & v845542;
assign v1215cd5 = hmaster0_p & v1215c91 | !hmaster0_p & v1215cd4;
assign d3019c = hlock5_p & d3019b | !hlock5_p & d30913;
assign v1553091 = hlock2 & v155341e | !hlock2 & v1553061;
assign v1445509 = hbusreq2_p & v1445508 | !hbusreq2_p & v1445bdb;
assign a65ae6 = hbusreq5_p & a662cb | !hbusreq5_p & a65ae5;
assign v12af5c4 = decide_p & v12af5b0 | !decide_p & v12afe76;
assign v1445b17 = hmaster1_p & v1445af7 | !hmaster1_p & v144591b;
assign v1216a75 = stateA1_p & v845542 | !stateA1_p & !a65854;
assign v14460fa = hmaster1_p & v1445fa9 | !hmaster1_p & v1445f9e;
assign v14058a2 = hmaster2_p & v140589a | !hmaster2_p & v1405845;
assign v1214ceb = hgrant4_p & v1214c29 | !hgrant4_p & v1214cea;
assign v12160b9 = hbusreq3 & v12160ac | !hbusreq3 & v12160b8;
assign v1215328 = hmaster0_p & v1215471 | !hmaster0_p & v1215061;
assign v14460cf = hmaster0_p & v14460ce | !hmaster0_p & v1446072;
assign v12ad50f = busreq_p & v138a322 | !busreq_p & v12ad50e;
assign v1668c7e = hmaster1_p & v1668c75 | !hmaster1_p & v1668c7d;
assign v1284d48 = hgrant0_p & v140583c | !hgrant0_p & !v1405928;
assign d307b8 = hmaster2_p & d307b7 | !hmaster2_p & d30655;
assign v1215fb6 = hmaster0_p & v12164e3 | !hmaster0_p & v12166f3;
assign d306a0 = hbusreq5 & d30699 | !hbusreq5 & d3069f;
assign v12150e1 = hlock2_p & v12150e0 | !hlock2_p & v12150d3;
assign v1215fed = hbusreq1 & v1215fec | !hbusreq1 & v845542;
assign d30100 = hgrant5_p & d2fe8b | !hgrant5_p & d300ff;
assign v10d42ce = hgrant2_p & v10d40b9 | !hgrant2_p & !v10d42cd;
assign d30699 = hbusreq2 & d30697 | !hbusreq2 & d30698;
assign d307f2 = hbusreq5_p & d307f1 | !hbusreq5_p & d307f0;
assign v16a1d54 = hgrant2_p & v845542 | !hgrant2_p & v16a1d53;
assign v14461de = hbusreq3 & v14461dc | !hbusreq3 & v14461dd;
assign v144536c = hmaster1_p & v1445a5a | !hmaster1_p & v1445a32;
assign v10d40cf = hbusreq2_p & v10d40ca | !hbusreq2_p & v10d40ce;
assign v121579e = hbusreq0 & v121579c | !hbusreq0 & v121579d;
assign v12aeb40 = hbusreq3 & v12aeb23 | !hbusreq3 & v12afe3d;
assign v14458fa = hmaster2_p & v14458f6 | !hmaster2_p & v1446429;
assign v1515ae3 = hbusreq2_p & v1515ae2 | !hbusreq2_p & !v845542;
assign v144645e = decide_p & v1446402 | !decide_p & v144645d;
assign v16a197f = hmaster0_p & v16a197c | !hmaster0_p & v16a197e;
assign v144548f = hmaster1_p & v144546c | !hmaster1_p & v1446290;
assign v1552f5c = hlock0 & v1552f5b | !hlock0 & v1552f5a;
assign v1445bba = hmaster1_p & v1445bb9 | !hmaster1_p & v1445bb7;
assign v138a459 = hmaster0_p & v138a354 | !hmaster0_p & v138a344;
assign v16a1416 = hmaster1_p & v16a140d | !hmaster1_p & v16a1f96;
assign v1446111 = hbusreq2 & v144610f | !hbusreq2 & v1446110;
assign f2f3f1 = hmaster1_p & f2f2dd | !hmaster1_p & f2f2db;
assign stateG10_3 = !v14eb679;
assign v1215d72 = hmaster2_p & v12166ce | !hmaster2_p & !v12164d9;
assign d2febc = hmaster2_p & v84555a | !hmaster2_p & d2feba;
assign f2f3ce = hbusreq0 & f2f3ca | !hbusreq0 & f2f3cd;
assign f2f438 = hbusreq5_p & f2f38f | !hbusreq5_p & f2f437;
assign d30898 = hgrant5_p & d30896 | !hgrant5_p & d30897;
assign v1515848 = hbusreq0 & v1515844 | !hbusreq0 & v1515847;
assign v11e593b = hmaster2_p & v845542 | !hmaster2_p & !v11e593a;
assign v1215026 = hbusreq4_p & v1215025 | !hbusreq4_p & v845547;
assign v1553147 = hlock4_p & v1553140 | !hlock4_p & v845542;
assign v144614e = hlock2 & v144614b | !hlock2 & v144614d;
assign a658fb = hmaster0_p & a658ee | !hmaster0_p & a658b7;
assign v12ad563 = hbusreq5 & v12ad548 | !hbusreq5 & v12ad562;
assign v14454f0 = hmaster0_p & v14454ef | !hmaster0_p & v1445414;
assign v121535a = hmaster0_p & v1215349 | !hmaster0_p & v1215359;
assign v12af9d0 = hbusreq4_p & v12afe60 | !hbusreq4_p & v12af9cf;
assign v1668c72 = hmaster0_p & v1668c67 | !hmaster0_p & v1668c71;
assign d300cd = hgrant1_p & d300b8 | !hgrant1_p & d300cc;
assign d30152 = hgrant5_p & v84555a | !hgrant5_p & d30114;
assign d3063f = decide_p & d3063e | !decide_p & v845570;
assign v1215721 = hgrant1_p & v121571a | !hgrant1_p & v1215720;
assign v1445455 = hlock2 & v1445446 | !hlock2 & v1445454;
assign v144590b = hmaster1_p & v144590a | !hmaster1_p & v14458fd;
assign v151575a = hgrant1_p & v151574f | !hgrant1_p & v1515755;
assign v1214ed5 = hgrant5_p & v845547 | !hgrant5_p & v1214ed3;
assign f2e4d1 = hmaster1_p & f2f229 | !hmaster1_p & f2e4d0;
assign v1445af2 = hbusreq2_p & v1445aef | !hbusreq2_p & v1445af1;
assign v12166ee = hbusreq0 & v12166e1 | !hbusreq0 & v12166ed;
assign v1214dab = hgrant2_p & v1214da8 | !hgrant2_p & v1214daa;
assign v12af5b0 = hgrant2_p & v845542 | !hgrant2_p & v12af5af;
assign v1216071 = hmaster0_p & v1216068 | !hmaster0_p & v121604c;
assign v138a443 = hbusreq5_p & v138a3f7 | !hbusreq5_p & !v845542;
assign v144578c = hmaster0_p & v144578b | !hmaster0_p & v1445de7;
assign d306ae = hgrant4_p & d30660 | !hgrant4_p & d306a4;
assign v1214dbc = hbusreq2_p & v1214dbb | !hbusreq2_p & v1214db9;
assign v12acfc9 = hmaster0_p & v12ad536 | !hmaster0_p & v12ad517;
assign v15530ae = hbusreq3 & v15530ad | !hbusreq3 & v155321a;
assign v1215cf7 = hgrant5_p & v845542 | !hgrant5_p & v1215cc3;
assign v15156ce = hbusreq3 & v15156b5 | !hbusreq3 & v15156cd;
assign v1446457 = hbusreq2 & v144644c | !hbusreq2 & v1446456;
assign v12152fa = hbusreq2_p & v12152f7 | !hbusreq2_p & !v12152f9;
assign v1405905 = hgrant3_p & v1405882 | !hgrant3_p & v1405904;
assign d308d1 = hready_p & d308d0 | !hready_p & d3087b;
assign v1214c19 = hbusreq2_p & v1214c18 | !hbusreq2_p & v1214c17;
assign d305de = locked_p & d305dd | !locked_p & v845542;
assign v15156e6 = hmaster1_p & v151567f | !hmaster1_p & v15156e5;
assign v134d4ef = hbusreq5_p & v134d4ec | !hbusreq5_p & v134d4ee;
assign a66291 = hbusreq5_p & a66290 | !hbusreq5_p & a6628c;
assign v12166c8 = hbusreq5_p & v12166c7 | !hbusreq5_p & v16a2243;
assign v1445877 = hgrant5_p & v1445874 | !hgrant5_p & !v1445876;
assign v16a266a = hbusreq5_p & v16a2669 | !hbusreq5_p & !v845542;
assign v1214dad = hmaster1_p & v1214dac | !hmaster1_p & v1214c39;
assign v144639e = hmastlock_p & v144639d | !hmastlock_p & v845542;
assign f2e500 = decide_p & f2e4ff | !decide_p & f2f23c;
assign v1446394 = stateG3_0_p & v845586 | !stateG3_0_p & !v845542;
assign d2fd17 = hbusreq5 & d2fd12 | !hbusreq5 & d2fd16;
assign v134ce43 = hmaster2_p & v134ce42 | !hmaster2_p & v134d386;
assign v138a05a = hready_p & v138a03a | !hready_p & v138a059;
assign v1405b49 = hlock0_p & v1405ad3 | !hlock0_p & v1405b48;
assign v1668c95 = hbusreq3 & v1668c8f | !hbusreq3 & a7c7c1;
assign v1446193 = hmaster0_p & v1445fea | !hmaster0_p & v14460a5;
assign v1216117 = hmaster2_p & v1215fef | !hmaster2_p & v845542;
assign v1284d13 = hmaster2_p & v14058f4 | !hmaster2_p & v1284d10;
assign v16a19c5 = hbusreq2 & v16a19c2 | !hbusreq2 & v16a19c4;
assign d2fd30 = decide_p & d2fd2f | !decide_p & v845570;
assign v134d262 = hmaster1_p & v134d20a | !hmaster1_p & v134d20f;
assign v16a19cb = hbusreq3 & v16a19c5 | !hbusreq3 & v16a19ca;
assign a65853 = hburst0_p & v155392f | !hburst0_p & !v845542;
assign v16695a0 = hmaster0_p & v1668c2e | !hmaster0_p & v845542;
assign a65658 = hgrant2_p & a6540a | !hgrant2_p & a65616;
assign v12162ff = hlock5_p & v12162fd | !hlock5_p & v12162fe;
assign f2f29c = hbusreq5_p & f2f298 | !hbusreq5_p & f2f29b;
assign v121621b = hgrant1_p & v845542 | !hgrant1_p & v121621a;
assign v12166ce = hready & v12166ca | !hready & v12166cd;
assign v1445e95 = hgrant5_p & v1445e00 | !hgrant5_p & v1445e94;
assign v12adbeb = hready_p & v12ae209 | !hready_p & v12adbea;
assign v1445828 = hlock2 & v1445823 | !hlock2 & v1445827;
assign v1215baf = hmaster2_p & v1215bac | !hmaster2_p & v1215bae;
assign v15530b0 = hbusreq5 & v15530ae | !hbusreq5 & v15530af;
assign v134cd55 = hbusreq4 & v134d36e | !hbusreq4 & v134d273;
assign a65380 = hgrant4_p & v845570 | !hgrant4_p & !a6537f;
assign v12160bf = hmaster1_p & v12160a8 | !hmaster1_p & v1216082;
assign v1214c82 = hlock2_p & v1214c81 | !hlock2_p & v121657d;
assign v138a44c = hmaster1_p & v138a344 | !hmaster1_p & v138a341;
assign v14464a8 = hmaster1_p & v14464a7 | !hmaster1_p & v845542;
assign v1216aa4 = hburst1_p & v845584 | !hburst1_p & v1216aa3;
assign v14460a5 = hlock0 & v14460a4 | !hlock0 & v14460a3;
assign d2fade = hbusreq1_p & d300e7 | !hbusreq1_p & d2fadd;
assign d2fbfa = hlock5_p & d2fbf8 | !hlock5_p & d2fbf9;
assign v1445442 = decide_p & v1445441 | !decide_p & v144639b;
assign v1445e73 = hbusreq1 & v1445e60 | !hbusreq1 & v1445e72;
assign v1515716 = hlock0_p & v1515609 | !hlock0_p & v10d3fd4;
assign d2fd1a = hready_p & d2fc8f | !hready_p & d2fd19;
assign a662cc = hmaster2_p & a662ca | !hmaster2_p & a6628b;
assign a6565c = hbusreq2_p & a65658 | !hbusreq2_p & !a6565a;
assign v16a1cdf = hbusreq2_p & v16a1b65 | !hbusreq2_p & v16a1cde;
assign v1215466 = hbusreq4_p & v1215465 | !hbusreq4_p & v845542;
assign v12147f1 = hbusreq2 & v12147f0 | !hbusreq2 & v12164e7;
assign d307d2 = hlock4_p & d307cf | !hlock4_p & d307d1;
assign v1214bcb = hmaster2_p & v1215364 | !hmaster2_p & v121539d;
assign v12ad597 = hmaster1_p & v12ad596 | !hmaster1_p & v12ad4dd;
assign v1216557 = hgrant0_p & v1216556 | !hgrant0_p & v845542;
assign v14457f5 = hgrant2_p & v14457f3 | !hgrant2_p & v14457f4;
assign v14466d7 = hbusreq3 & v14466d5 | !hbusreq3 & v14466d6;
assign v10d426e = hgrant5_p & v10d3ff1 | !hgrant5_p & !v10d426c;
assign v12ad548 = hbusreq3 & v12ad53a | !hbusreq3 & v12ad547;
assign v12ae6db = hready_p & v845542 | !hready_p & v12ae6da;
assign v10d40c9 = hmaster1_p & v10d40c8 | !hmaster1_p & !v10d407c;
assign v144629a = hlock2 & v1446275 | !hlock2 & v1446298;
assign v1446198 = hbusreq2 & v1446192 | !hbusreq2 & v1446197;
assign d306f1 = hburst0 & d306ee | !hburst0 & d306f0;
assign v12afda1 = hlock0_p & a66275 | !hlock0_p & !v845542;
assign v14460e7 = hmaster0_p & v1445fa2 | !hmaster0_p & v144639c;
assign d30616 = hlock2_p & d30615 | !hlock2_p & d3060e;
assign v144643e = hbusreq5_p & v144643d | !hbusreq5_p & v144643b;
assign v1216007 = hlock0_p & v1216a5a | !hlock0_p & v1216006;
assign v1216148 = hbusreq4_p & v1216145 | !hbusreq4_p & v1216147;
assign v1446719 = hbusreq2_p & v1446713 | !hbusreq2_p & v1446718;
assign v14838b9 = hready_p & v845558 | !hready_p & v14838b8;
assign v14460d9 = hgrant2_p & v14460c2 | !hgrant2_p & v14460d5;
assign v14457fd = hgrant2_p & v14457f8 | !hgrant2_p & v14457e9;
assign d2fbd5 = hgrant1_p & d2fbcb | !hgrant1_p & d2fbd4;
assign v12ad32d = decide_p & v12ad32c | !decide_p & v12afe76;
assign v14466df = hlock2 & v14466db | !hlock2 & v14466de;
assign v1446743 = hbusreq2_p & v1446729 | !hbusreq2_p & v1446742;
assign v1389816 = hbusreq5_p & v1389815 | !hbusreq5_p & !v845542;
assign v144621a = hmaster1_p & v144639c | !hmaster1_p & v1446219;
assign v144548e = hbusreq3 & v144548a | !hbusreq3 & v144548d;
assign f2f337 = hbusreq2 & f2f333 | !hbusreq2 & f2f336;
assign d2fba1 = hbusreq2_p & d2fba0 | !hbusreq2_p & d2fb9f;
assign v12153ea = hmaster2_p & v845542 | !hmaster2_p & v12153e9;
assign v1284d2d = hmaster1_p & v1284d2c | !hmaster1_p & v140584d;
assign d30109 = hgrant5_p & d2fe8b | !hgrant5_p & d30108;
assign v16a19e3 = hbusreq2 & v16a19dd | !hbusreq2 & v16a19e2;
assign v134d3ba = hbusreq5 & v134d3b9 | !hbusreq5 & v134d3b5;
assign v1515760 = hbusreq1 & v10d3ff7 | !hbusreq1 & !v845542;
assign v1215d35 = hmaster2_p & v1216594 | !hmaster2_p & !v1216a93;
assign v138a407 = decide_p & v138a405 | !decide_p & v138a406;
assign v14454a3 = hlock5 & v144548e | !hlock5 & v144549f;
assign v1215d89 = hmaster0_p & v1215d6c | !hmaster0_p & v1215d88;
assign v11e595a = hmaster2_p & v11e5955 | !hmaster2_p & v11e5959;
assign v16a138e = hbusreq3 & v16a1389 | !hbusreq3 & v16a138d;
assign v1552d6d = hready_p & v1553306 | !hready_p & v1552d6c;
assign v12ad617 = hmaster0_p & v12ad612 | !hmaster0_p & !v12ad616;
assign v1445924 = hlock3 & v1445912 | !hlock3 & v1445923;
assign v134d4d3 = hgrant4_p & v134d4d2 | !hgrant4_p & v845542;
assign v16a1432 = decide_p & v16a1429 | !decide_p & !v16a141b;
assign f2f2ee = hmaster1_p & f2f2ed | !hmaster1_p & f2f2db;
assign v1215110 = hbusreq2_p & v121510d | !hbusreq2_p & v121510f;
assign v134d4f9 = hbusreq4_p & v134d273 | !hbusreq4_p & v134d4e6;
assign d2fb10 = hmaster0_p & d2fafe | !hmaster0_p & d2fb0f;
assign v16a1bc5 = hgrant1_p & v84554d | !hgrant1_p & v16a1bc4;
assign v134d1e8 = hmastlock_p & v134d1e7 | !hmastlock_p & v845542;
assign v138a34f = hbusreq5_p & v138a34e | !hbusreq5_p & !v845542;
assign v134ce37 = hbusreq1_p & v134d273 | !hbusreq1_p & v134ce36;
assign v1215093 = hgrant0_p & v1215465 | !hgrant0_p & !v845559;
assign a65b2b = hbusreq5_p & a6628c | !hbusreq5_p & a662ad;
assign v12ad5f1 = hmaster0_p & v12ad4e9 | !hmaster0_p & v12ad4e8;
assign v114a231 = hgrant1_p & v845542 | !hgrant1_p & !v114a230;
assign v144539f = hlock2 & v1445354 | !hlock2 & v144539e;
assign d30712 = hlock3_p & d306fb | !hlock3_p & !d30711;
assign d2fb13 = hbusreq2_p & d2fad4 | !hbusreq2_p & !d2fb12;
assign v1515850 = decide_p & v151584f | !decide_p & v845576;
assign d306c1 = hgrant2_p & v845542 | !hgrant2_p & !d306c0;
assign v155342b = hmaster2_p & v155342a | !hmaster2_p & v845542;
assign v10d4062 = hgrant1_p & v10d3fdb | !hgrant1_p & v10d4061;
assign bf1f80 = hgrant1_p & bf1f52 | !hgrant1_p & !bf1f7f;
assign v1215ddb = hready_p & v845542 | !hready_p & v1215dda;
assign v14459ec = hgrant1_p & v14458e2 | !hgrant1_p & v14459cb;
assign v1669595 = hmaster0_p & v1668c17 | !hmaster0_p & v845570;
assign v1215410 = hmaster1_p & v12153d4 | !hmaster1_p & v121540f;
assign d30828 = hgrant5_p & v84554e | !hgrant5_p & d307dc;
assign v16a1a25 = hbusreq2_p & v16a1889 | !hbusreq2_p & v16a1a24;
assign v16a1cd3 = hbusreq2_p & v16a1aff | !hbusreq2_p & v16a1cd2;
assign v134d3b2 = hlock2 & v134d39c | !hlock2 & v134d3b1;
assign d2faed = hgrant1_p & d2fade | !hgrant1_p & d2faec;
assign d30130 = hgrant5_p & v84555a | !hgrant5_p & d300c5;
assign d3089b = hgrant5_p & d30896 | !hgrant5_p & d3089a;
assign d305f7 = hbusreq5_p & d305f6 | !hbusreq5_p & v84554e;
assign v1216a90 = hmaster2_p & v845570 | !hmaster2_p & v16a1bc6;
assign v14453f1 = hbusreq5 & v14453ef | !hbusreq5 & v14453f0;
assign v1668d75 = hbusreq1_p & v1668d73 | !hbusreq1_p & v1668d74;
assign v16a1ac9 = hbusreq5_p & v845542 | !hbusreq5_p & !v845568;
assign v12164c8 = hlock2_p & v12164c7 | !hlock2_p & v12164c3;
assign d2fb16 = hbusreq2_p & d2fb14 | !hbusreq2_p & d2fb15;
assign v1668d1b = hbusreq5_p & v1668d19 | !hbusreq5_p & v1668d1a;
assign v1215071 = hbusreq2_p & v121506d | !hbusreq2_p & v1215070;
assign v14461f0 = hgrant2_p & v14461c5 | !hgrant2_p & v14461ef;
assign v14453b8 = hgrant2_p & v1445397 | !hgrant2_p & v14453b7;
assign v1552f74 = hlock2 & v1552f6b | !hlock2 & v1552f73;
assign v1445423 = hbusreq2_p & v1445422 | !hbusreq2_p & v144541b;
assign v10d4283 = hgrant0_p & v10d3fd5 | !hgrant0_p & !v10d4282;
assign v144537f = hbusreq2_p & v144537b | !hbusreq2_p & v144537e;
assign v134d1dc = hmastlock_p & v134d1db | !hmastlock_p & v845542;
assign v1215cc9 = hmaster1_p & v1215c9f | !hmaster1_p & v1215cc8;
assign v14465d2 = hgrant1_p & v14465c7 | !hgrant1_p & v14465d1;
assign v12153c2 = hmaster1_p & v12153c1 | !hmaster1_p & v12153bf;
assign v12adf67 = hready_p & v845542 | !hready_p & v12adf66;
assign v16a2248 = hmaster1_p & v16a2247 | !hmaster1_p & !v16a2672;
assign v134d3fb = decide_p & v134d3fa | !decide_p & v134d276;
assign v10d4296 = hmaster2_p & v10d428b | !hmaster2_p & !v10d4295;
assign v16a1adb = hgrant1_p & v84554d | !hgrant1_p & v16a1ada;
assign v121575a = hgrant0_p & v1215759 | !hgrant0_p & v845542;
assign v12afa32 = decide_p & v12af9b7 | !decide_p & v12afe76;
assign v15168a9 = stateA1_p & d30714 | !stateA1_p & v156645f;
assign v121626c = hgrant3_p & v12160e7 | !hgrant3_p & v121626b;
assign d2ff07 = hlock2_p & d2ff06 | !hlock2_p & d2ff03;
assign d2f999 = hbusreq4_p & d2feb1 | !hbusreq4_p & v845548;
assign v16a1be3 = hgrant5_p & v845542 | !hgrant5_p & !v16a1bcf;
assign v12ad529 = hmaster0_p & v12ad517 | !hmaster0_p & v12ad528;
assign d2feaa = hmaster0_p & d2fea9 | !hmaster0_p & v84555a;
assign v12adf64 = hmaster0_p & v845542 | !hmaster0_p & v12adf63;
assign v131be8c = hready_p & v84555c | !hready_p & v131be8b;
assign v10d42bc = hbusreq2_p & v10d42b6 | !hbusreq2_p & v10d42bb;
assign v144632c = hmaster0_p & v14465b7 | !hmaster0_p & v1446310;
assign v121577d = hbusreq5_p & v121577b | !hbusreq5_p & !v121577c;
assign v1553218 = hmaster2_p & v845542 | !hmaster2_p & v1553217;
assign v1446463 = hgrant4_p & v845542 | !hgrant4_p & v1446462;
assign d305fd = hlock5_p & v845542 | !hlock5_p & d305fc;
assign d30218 = hmaster0_p & d30202 | !hmaster0_p & d30217;
assign v1214d40 = decide_p & v1214d3a | !decide_p & v1214d3f;
assign f2f28e = decide_p & f2f28d | !decide_p & f2f23c;
assign v10d42b4 = hgrant5_p & v10d400b | !hgrant5_p & v10d42b3;
assign v10d400e = hmaster2_p & v10d3fd4 | !hmaster2_p & !v10d3fe0;
assign d2fc74 = hbusreq0 & d2fc73 | !hbusreq0 & d302e7;
assign d30854 = hbusreq1_p & d30701 | !hbusreq1_p & !v845542;
assign v1515c85 = hbusreq2_p & v1515c84 | !hbusreq2_p & v845542;
assign v144581b = hlock3 & v14457f6 | !hlock3 & v1445819;
assign v1405b38 = hmaster1_p & v1405b37 | !hmaster1_p & !v1405a94;
assign v14457bd = hmaster1_p & v1445791 | !hmaster1_p & v1445e28;
assign d2fb0c = hmaster2_p & d306b0 | !hmaster2_p & d2fb0b;
assign v1284cbf = hbusreq2_p & v1284cbb | !hbusreq2_p & v1284cbe;
assign v14453a6 = hgrant2_p & v1445379 | !hgrant2_p & v14453a5;
assign v1214f7e = hready_p & v1214f6b | !hready_p & v1214f7d;
assign v140590d = hmaster0_p & v14058db | !hmaster0_p & v140584f;
assign f2f41b = hmaster0_p & f2f3a1 | !hmaster0_p & f2f396;
assign v1215bc4 = hmaster1_p & v845542 | !hmaster1_p & v1215bc2;
assign v1446484 = hgrant4_p & v845542 | !hgrant4_p & v1446483;
assign v1445a4f = hlock0 & v1445a4b | !hlock0 & v1445a4e;
assign v1515611 = hbusreq5_p & v151560f | !hbusreq5_p & v1515610;
assign v14458ec = hmaster2_p & v1446403 | !hmaster2_p & v14458eb;
assign v1215080 = hbusreq2_p & v121507d | !hbusreq2_p & v121507f;
assign v1446747 = hmaster1_p & v1446746 | !hmaster1_p & v1446436;
assign d807b1 = hgrant2_p & d807b0 | !hgrant2_p & d807ac;
assign v1446694 = hbusreq0 & v1446693 | !hbusreq0 & v14465e4;
assign a65371 = hgrant4_p & v845570 | !hgrant4_p & !a65370;
assign v1216053 = hbusreq1_p & v1216052 | !hbusreq1_p & v845542;
assign v1405b2d = hgrant5_p & v1405aca | !hgrant5_p & v1405b2c;
assign v1668cfd = hmaster0_p & v1668cfc | !hmaster0_p & !v1668cd5;
assign v134d46c = hbusreq3_p & v134d45e | !hbusreq3_p & v134d46b;
assign v1214d77 = hmaster0_p & v1214c7b | !hmaster0_p & v1214c56;
assign v1215c4b = hmaster0_p & v845542 | !hmaster0_p & v1215c4a;
assign v1216058 = hbusreq1 & v1216af3 | !hbusreq1 & !v845542;
assign v1215fea = hbusreq1_p & v1215fe9 | !hbusreq1_p & v845542;
assign v1214e62 = hmaster0_p & v1216b01 | !hmaster0_p & v845542;
assign v12afe3d = hmaster1_p & v845542 | !hmaster1_p & v12afe3c;
assign v1215ce2 = hgrant5_p & v845542 | !hgrant5_p & v1215c88;
assign v1668cb6 = hbusreq5 & v1668c95 | !hbusreq5 & v1668cb5;
assign v144655f = hgrant1_p & v845542 | !hgrant1_p & v144655e;
assign v134d535 = hlock2 & v134d534 | !hlock2 & v134d532;
assign d306d5 = hbusreq1 & d306d4 | !hbusreq1 & v845542;
assign v121500f = hlock0_p & v1215bad | !hlock0_p & v121500e;
assign v12150f7 = hbusreq2 & v12150f3 | !hbusreq2 & v12150f6;
assign v121602c = hbusreq2_p & v1216028 | !hbusreq2_p & v121602b;
assign v16a1bd7 = hmaster2_p & v16a206f | !hmaster2_p & v16a1bd6;
assign a653a2 = hbusreq1_p & a65376 | !hbusreq1_p & a653a1;
assign v12166e2 = stateA1_p & v1446394 | !stateA1_p & a66292;
assign v1446467 = hmaster2_p & v1446398 | !hmaster2_p & v845542;
assign f2f44c = hgrant5_p & f2f3c1 | !hgrant5_p & f2f42b;
assign v12152f2 = hgrant2_p & v1215786 | !hgrant2_p & v12152ee;
assign v144612b = hmaster1_p & v144612a | !hmaster1_p & v1445fde;
assign v134ce7f = hbusreq3_p & v134ce71 | !hbusreq3_p & v134ce7e;
assign v134d530 = decide_p & v845542 | !decide_p & v134d52f;
assign v14461e4 = hbusreq2_p & v14461e1 | !hbusreq2_p & v14461e3;
assign v16a1c9a = hmaster2_p & v16a1c99 | !hmaster2_p & !v845542;
assign d301cb = hmaster1_p & d301c4 | !hmaster1_p & !d301ca;
assign v1515745 = hbusreq4 & v10d3fdf | !hbusreq4 & v845542;
assign v1446116 = hlock5 & v14460f2 | !hlock5 & v1446114;
assign d30691 = hmaster2_p & d3068e | !hmaster2_p & d30690;
assign v1216067 = hbusreq1_p & v1216066 | !hbusreq1_p & v845542;
assign v15155e5 = hbusreq3_p & v1515bb0 | !hbusreq3_p & v15155e4;
assign v1215c38 = hmaster0_p & v121601c | !hmaster0_p & v1216172;
assign v1216522 = hbusreq1_p & v1216521 | !hbusreq1_p & v16a1c95;
assign v1552fcc = hmaster1_p & v1552fcb | !hmaster1_p & v845542;
assign v1445db6 = hmaster2_p & v144639c | !hmaster2_p & v1445db5;
assign f2f43f = hgrant2_p & f2f3b4 | !hgrant2_p & !f2f43b;
assign v134ce84 = hmaster0_p & v134ce83 | !hmaster0_p & v134d20a;
assign v1445430 = hbusreq2 & v144542a | !hbusreq2 & v144542f;
assign v13891a8 = hready_p & v845542 | !hready_p & v13891a7;
assign v1405858 = hmaster1_p & v1405857 | !hmaster1_p & v140584d;
assign v134d233 = hmaster1_p & v134d232 | !hmaster1_p & v134d208;
assign v14461cc = hgrant2_p & v14461c5 | !hgrant2_p & v14461c6;
assign v144633f = hbusreq0 & v14466a2 | !hbusreq0 & v1446616;
assign v15168ff = hbusreq2 & v15168ef | !hbusreq2 & v15168fe;
assign v1445f67 = hgrant2_p & v144672b | !hgrant2_p & v1445f66;
assign d2fb6a = hlock0_p & v845542 | !hlock0_p & d305ea;
assign v14453bf = hlock3 & v14453b1 | !hlock3 & v14453be;
assign v16a1a31 = hready_p & v845555 | !hready_p & v16a1a30;
assign v1446321 = hbusreq0 & v1446320 | !hbusreq0 & v1446310;
assign v1214f09 = hgrant5_p & v1215c5b | !hgrant5_p & v1214edf;
assign v12164ce = hlock3_p & v12164c0 | !hlock3_p & v12164cd;
assign v14463fa = hmaster1_p & v14463ca | !hmaster1_p & v14463ef;
assign v12ad613 = hgrant5_p & v12ad4eb | !hgrant5_p & v12ad5dc;
assign v138a074 = hbusreq5 & v138a06a | !hbusreq5 & v138a391;
assign d3080b = hmaster2_p & d306d0 | !hmaster2_p & d3080a;
assign d30895 = hbusreq0 & d3088d | !hbusreq0 & d30894;
assign d30625 = hbusreq2_p & d30624 | !hbusreq2_p & d3061f;
assign d3082f = hbusreq0 & d3082a | !hbusreq0 & d3082e;
assign v1446322 = hlock0 & v1446321 | !hlock0 & v1446320;
assign v16a1c02 = hgrant2_p & v845542 | !hgrant2_p & v16a1c00;
assign v16a1d0f = hbusreq2 & v16a1d0e | !hbusreq2 & v16a205c;
assign d2fc29 = hbusreq2_p & v84554a | !hbusreq2_p & d2fc28;
assign v155321a = hmaster1_p & v1553219 | !hmaster1_p & v845542;
assign v1445bb7 = hmaster0_p & v1445bb6 | !hmaster0_p & v144642a;
assign v1216acc = stateA1_p & v845542 | !stateA1_p & afe156;
assign v1446158 = hlock2 & v1446125 | !hlock2 & v1446156;
assign v140592a = hbusreq4_p & v140588f | !hbusreq4_p & v1405929;
assign v15157b2 = hbusreq5_p & v15157b0 | !hbusreq5_p & !v15157b1;
assign v1446314 = hmaster1_p & v1446313 | !hmaster1_p & v14462ff;
assign d302f5 = hready_p & d302f4 | !hready_p & d302f1;
assign v1215c9c = hgrant5_p & v845542 | !hgrant5_p & !v1215c9a;
assign v138a3ca = hbusreq5_p & v138a3c9 | !hbusreq5_p & !v845542;
assign v1405b5b = hmaster0_p & v1405aca | !hmaster0_p & v1405abc;
assign v14058cf = hgrant4_p & v14058ce | !hgrant4_p & v1405849;
assign v1216543 = hgrant5_p & v845542 | !hgrant5_p & v1216542;
assign d2fbea = hbusreq4_p & d2fbe9 | !hbusreq4_p & v84554a;
assign a6545a = hmaster1_p & a65459 | !hmaster1_p & a653f3;
assign v151572f = hgrant5_p & v151570f | !hgrant5_p & v151572e;
assign d30918 = hmaster0_p & d30915 | !hmaster0_p & d30917;
assign v12162ce = hmaster1_p & v12162bf | !hmaster1_p & !v121624b;
assign v1216aef = hmaster2_p & v1216ad6 | !hmaster2_p & v1216aee;
assign v1445f8b = hgrant5_p & v1445f88 | !hgrant5_p & !v1445f8a;
assign v14460d5 = hmaster1_p & v1446093 | !hmaster1_p & v14460cf;
assign f2f447 = hgrant5_p & v84554c | !hgrant5_p & f2f424;
assign v1445806 = hmaster1_p & v1445805 | !hmaster1_p & v1445eaa;
assign v1215fe8 = hready & d306c8 | !hready & v845570;
assign v1214cc4 = hmastlock_p & v1214cc3 | !hmastlock_p & !v845542;
assign v16a1dfd = hbusreq2 & v16a1dec | !hbusreq2 & v16a1ded;
assign a65857 = stateA1_p & v845542 | !stateA1_p & !a65856;
assign v15167e8 = hmaster0_p & v845542 | !hmaster0_p & v1668c29;
assign v12af222 = hbusreq1_p & v12af5a8 | !hbusreq1_p & v12af9d1;
assign a654bd = hmaster1_p & a65499 | !hmaster1_p & !a654b0;
assign v134cd8f = hgrant3_p & v134d3fc | !hgrant3_p & v134cd8e;
assign v1214cf7 = hgrant5_p & v1214cf0 | !hgrant5_p & v1214cf6;
assign v1446002 = hlock2 & v1445fff | !hlock2 & v1446001;
assign v1446123 = hmaster0_p & v1446077 | !hmaster0_p & v1445fe1;
assign v1553104 = hbusreq5 & v1553102 | !hbusreq5 & v1553103;
assign v1215ffa = hbusreq1_p & v1215ff9 | !hbusreq1_p & v845542;
assign v12ae1fe = hbusreq0 & v12ae1f3 | !hbusreq0 & v12ae1fd;
assign v16a1d39 = hgrant1_p & v84554d | !hgrant1_p & v16a1bbb;
assign v14466ec = hlock3 & v14466d3 | !hlock3 & v14466ea;
assign a65455 = decide_p & a65454 | !decide_p & a662a2;
assign v1446267 = hlock0 & v1446266 | !hlock0 & v1446263;
assign v1445e84 = hbusreq5_p & v1445e7e | !hbusreq5_p & v1445e83;
assign f2f225 = hready_p & v845542 | !hready_p & f2f224;
assign v1446053 = hbusreq5_p & v1446042 | !hbusreq5_p & v1446052;
assign v12acfb5 = hbusreq1_p & v12ad522 | !hbusreq1_p & v12acfb4;
assign v138a362 = hmaster0_p & v138a34b | !hmaster0_p & v138a354;
assign v134d507 = hgrant4_p & v845542 | !hgrant4_p & v134d506;
assign v1445e18 = hmaster1_p & v1445e17 | !hmaster1_p & v1445e07;
assign d306db = hbusreq1 & d306da | !hbusreq1 & v845542;
assign v1214df1 = hbusreq1 & v1216aad | !hbusreq1 & v1216ab8;
assign v1668cf7 = hbusreq3 & v1668cf6 | !hbusreq3 & v845542;
assign v1215094 = hbusreq4_p & v1215093 | !hbusreq4_p & v845542;
assign d3085b = hbusreq5_p & v84554e | !hbusreq5_p & d30654;
assign v1445dce = hbusreq5_p & v1445d86 | !hbusreq5_p & v1445dcd;
assign v1515738 = hgrant5_p & v151560b | !hgrant5_p & v1515737;
assign d302d5 = hmaster0_p & d308f5 | !hmaster0_p & d305fe;
assign v14454a7 = decide_p & v1445468 | !decide_p & v14454a6;
assign v144605e = hgrant1_p & v144605c | !hgrant1_p & v144605d;
assign d301b0 = hbusreq2_p & d301af | !hbusreq2_p & d301a9;
assign v1215cb1 = hgrant5_p & v1215ca0 | !hgrant5_p & v1215cb0;
assign v1284cef = hmaster2_p & v1405844 | !hmaster2_p & !v1284ceb;
assign v151584c = hgrant2_p & v15167ff | !hgrant2_p & !v151584b;
assign a6470c = hmaster1_p & a6470b | !hmaster1_p & a65b09;
assign v1553500 = hgrant2_p & v1553380 | !hgrant2_p & v15534ff;
assign v1446293 = hbusreq2_p & v1446291 | !hbusreq2_p & v1446292;
assign v1553423 = hbusreq5 & v1553422 | !hbusreq5 & v155341e;
assign v16a1e97 = hgrant1_p & v84554d | !hgrant1_p & v16a1e96;
assign v12153e5 = hmaster2_p & v845542 | !hmaster2_p & v12153e4;
assign v166959b = hbusreq3 & v1669596 | !hbusreq3 & v166959a;
assign v1445e6f = hlock1 & v1446606 | !hlock1 & v1445e55;
assign d301f4 = hgrant1_p & d301f3 | !hgrant1_p & d307b3;
assign d30840 = hgrant2_p & d30810 | !hgrant2_p & d30831;
assign v1668c23 = hmaster0_p & v1668c22 | !hmaster0_p & v1668c1f;
assign v1445d83 = hlock1 & v14463b9 | !hlock1 & v1445d81;
assign d2fc22 = hgrant3_p & d2fbc5 | !hgrant3_p & d2fc21;
assign v138a3d1 = hbusreq5_p & v138a3d0 | !hbusreq5_p & !v845542;
assign v140593f = hgrant3_p & v140591a | !hgrant3_p & v140593e;
assign v10d3fdf = hmastlock_p & v10d3fde | !hmastlock_p & v845542;
assign v11e5940 = hready_p & v11e593f | !hready_p & !v845542;
assign v1214bbf = hmaster0_p & v12153b1 | !hmaster0_p & v12153ab;
assign d3073e = hburst1 & d3073c | !hburst1 & d3073d;
assign d302e7 = hbusreq5_p & d302df | !hbusreq5_p & !d306ac;
assign v16a196d = hbusreq5 & v16a195f | !hbusreq5 & v16a196c;
assign v16a1d1e = hmaster2_p & v16a1d19 | !hmaster2_p & !v845542;
assign v12aec09 = hmaster0_p & v12afe47 | !hmaster0_p & v12aec08;
assign v1405b27 = hmaster2_p & v1405b24 | !hmaster2_p & v1405b26;
assign v16a1ce2 = hbusreq2_p & v16a1b67 | !hbusreq2_p & v16a1ce1;
assign v1446171 = hlock2 & v144616a | !hlock2 & v1446170;
assign v121652a = hgrant4_p & v1216524 | !hgrant4_p & v1216529;
assign v12afda5 = hbusreq5_p & v12afda2 | !hbusreq5_p & v12afda4;
assign v12153ef = hmaster0_p & v12153d4 | !hmaster0_p & v12153ee;
assign v16a1961 = hgrant5_p & v845542 | !hgrant5_p & !v16a194d;
assign bf1f89 = hready_p & bf1f74 | !hready_p & bf1f88;
assign bf1f67 = hgrant1_p & f2f227 | !hgrant1_p & bf1f66;
assign v12ad536 = hbusreq0 & v12ad535 | !hbusreq0 & !v845542;
assign v1445469 = hbusreq0 & v1446635 | !hbusreq0 & v144639c;
assign v1446438 = hlock1 & v1446407 | !hlock1 & v144640a;
assign v1445e60 = hgrant4_p & v1445e5e | !hgrant4_p & v1445e5f;
assign v12162d9 = hgrant2_p & v12162c8 | !hgrant2_p & v12162d8;
assign f2ed9e = hgrant3_p & f2ed91 | !hgrant3_p & f2ed9d;
assign d30861 = hbusreq3 & d3085a | !hbusreq3 & !d30860;
assign v14463dc = hmaster2_p & v144639c | !hmaster2_p & v14463db;
assign v134d38f = hlock0_p & v134d273 | !hlock0_p & v134d38e;
assign v1668c7a = hbusreq5_p & v1668c78 | !hbusreq5_p & !v1668c79;
assign v1515727 = hbusreq5_p & v1515725 | !hbusreq5_p & v1515726;
assign v1445790 = hbusreq2_p & v144578d | !hbusreq2_p & v144578f;
assign bf1f4f = hmaster1_p & bf1f4e | !hmaster1_p & v845542;
assign v16a1d92 = hmaster0_p & v16a1d8c | !hmaster0_p & v16a1d91;
assign v1215459 = hbusreq2_p & v1215458 | !hbusreq2_p & v1215457;
assign d306bf = hmaster0_p & d306bd | !hmaster0_p & d306be;
assign v1216aa7 = stateA1_p & v1216aa2 | !stateA1_p & v1216aa6;
assign v1389e36 = hbusreq5 & v1389dfb | !hbusreq5 & v1389e33;
assign v1215c5c = hgrant5_p & v1215c5b | !hgrant5_p & v1215c0e;
assign v1216202 = hmaster1_p & v1216201 | !hmaster1_p & v12160e0;
assign v1445f47 = hmaster0_p & v1445db8 | !hmaster0_p & v144639c;
assign v1445a3f = hbusreq0 & v1445a3c | !hbusreq0 & v1445a3e;
assign v1668de0 = hgrant2_p & v1668d94 | !hgrant2_p & v1668ddf;
assign v1405a87 = hmastlock_p & v845580 | !hmastlock_p & !v845542;
assign d3029c = hbusreq5 & d3028e | !hbusreq5 & d3029b;
assign v1214da7 = hmaster0_p & v1214c3c | !hmaster0_p & v1214c2c;
assign d30911 = hbusreq1_p & d30910 | !hbusreq1_p & !v845542;
assign a658da = hburst1 & v845542 | !hburst1 & v10d3fd6;
assign a662ba = hbusreq2_p & a6629f | !hbusreq2_p & a662b9;
assign bf1f6f = hmaster0_p & bf1f65 | !hmaster0_p & bf1f6e;
assign f2f3e4 = hready_p & f2f3e2 | !hready_p & f2f3e3;
assign v1515808 = decide_p & v1515807 | !decide_p & v845576;
assign v12160d2 = hbusreq1 & v12164d3 | !hbusreq1 & v845542;
assign f2f2da = hbusreq0 & f2f2d6 | !hbusreq0 & f2f2d9;
assign d807a8 = hgrant4_p & d80760 | !hgrant4_p & d807a7;
assign v1216709 = hmaster1_p & v1216708 | !hmaster1_p & v12166ef;
assign v140584d = hmaster0_p & v1405848 | !hmaster0_p & v140584c;
assign v15156d7 = hmaster2_p & v15156d6 | !hmaster2_p & !v1515658;
assign d30234 = hlock2_p & v845542 | !hlock2_p & d30233;
assign d8074a = hmaster1_p & d80749 | !hmaster1_p & d80746;
assign f2f2a5 = hmaster0_p & f2f296 | !hmaster0_p & f2f2a4;
assign f2e275 = hlock1_p & f2e274 | !hlock1_p & !v845542;
assign v1214c9f = hgrant2_p & v1214c9c | !hgrant2_p & v1214c98;
assign f2f3c7 = hbusreq0 & f2f3c3 | !hbusreq0 & f2f3c6;
assign v144671c = hbusreq2 & v144671a | !hbusreq2 & v144671b;
assign v845560 = hburst0_p & v845542 | !hburst0_p & !v845542;
assign v1214c03 = hbusreq2_p & v1214c02 | !hbusreq2_p & v1214c01;
assign v14457e1 = hbusreq2_p & v14457dc | !hbusreq2_p & v14457e0;
assign v16a1425 = hbusreq2 & v16a1424 | !hbusreq2 & v16a1ace;
assign v1445f8d = stateG10_5_p & v1445f89 | !stateG10_5_p & !v14463a5;
assign v121613c = hlock4_p & v121613b | !hlock4_p & !v845542;
assign v1445897 = hbusreq0_p & v14463e1 | !hbusreq0_p & v144639e;
assign v1668d00 = hbusreq5_p & v1668cff | !hbusreq5_p & v1668ce1;
assign v155305e = hbusreq0 & v155305d | !hbusreq0 & v15533a7;
assign v12acffe = hgrant1_p & v12ad59a | !hgrant1_p & v12acffd;
assign v1214f6f = hmaster1_p & v1214f6e | !hmaster1_p & v1215d68;
assign f2f4ad = stateA1_p & v146af2e | !stateA1_p & a658a3;
assign v1214c5c = hgrant1_p & v1214c5b | !hgrant1_p & v1214c50;
assign v134cdce = hgrant3_p & v134cdcb | !hgrant3_p & v134cdcd;
assign v12160b5 = hmaster1_p & v121606b | !hmaster1_p & v121605d;
assign v12162bd = hmaster0_p & v12160e2 | !hmaster0_p & v12160d4;
assign v134ce86 = hlock2_p & v134d23d | !hlock2_p & v134ce85;
assign v134d36d = locked_p & v134d36c | !locked_p & v845542;
assign bf1f7e = hgrant5_p & bf1f53 | !hgrant5_p & !bf1f7d;
assign v10d406c = hmaster2_p & v10d3fdf | !hmaster2_p & v10d3fe1;
assign v12afe74 = hgrant1_p & v845542 | !hgrant1_p & v114a230;
assign d305d8 = hmaster0_p & d305d5 | !hmaster0_p & d305d7;
assign v134d462 = hbusreq2 & v134d460 | !hbusreq2 & v134d461;
assign bf1f72 = hgrant2_p & bf1f59 | !hgrant2_p & !bf1f70;
assign v12ad520 = hbusreq0 & v12ad51f | !hbusreq0 & v845542;
assign v14463cf = hmaster0_p & v144639c | !hmaster0_p & v14463c7;
assign v1445e89 = hbusreq4_p & v1445e88 | !hbusreq4_p & v1446429;
assign v16a1db6 = hbusreq2_p & v16a1d55 | !hbusreq2_p & v16a1db5;
assign v1214ee8 = hgrant5_p & v1216a5a | !hgrant5_p & v121656d;
assign v1216285 = hmaster0_p & v121617d | !hmaster0_p & v1216116;
assign v144671f = hlock3 & v1446702 | !hlock3 & v144671c;
assign v121605e = hmaster1_p & v121604c | !hmaster1_p & v121605d;
assign v151574a = hmaster2_p & v1668d36 | !hmaster2_p & v1515749;
assign v121503f = hmaster2_p & v121503e | !hmaster2_p & v121503a;
assign v1446637 = hbusreq5_p & v1446635 | !hbusreq5_p & v1446636;
assign v121619b = hbusreq0 & v1216199 | !hbusreq0 & v121619a;
assign d306e1 = hlock1_p & d306e0 | !hlock1_p & v845570;
assign v16a19ad = hmaster1_p & v16a19ac | !hmaster1_p & !v16a2672;
assign v134ce5b = hbusreq2 & v134ce59 | !hbusreq2 & v134ce5a;
assign d2fcb1 = hmaster2_p & v845542 | !hmaster2_p & !d2fcaf;
assign v12af98f = hbusreq2_p & v12afdb5 | !hbusreq2_p & v12af98e;
assign v121606a = hmaster1_p & v1216069 | !hmaster1_p & v121605d;
assign v16a2069 = hmastlock_p & v16a2068 | !hmastlock_p & v845542;
assign v16a1f9c = hbusreq2 & v16a1f9a | !hbusreq2 & v16a1f9b;
assign v15534f5 = hlock2 & v155341e | !hlock2 & v15534dd;
assign v1215398 = hbusreq0_p & v1216acd | !hbusreq0_p & !v845542;
assign v1214c18 = hlock2_p & v1214c16 | !hlock2_p & v1214c17;
assign v134d20f = hmaster0_p & v134d201 | !hmaster0_p & v134d207;
assign v1216aff = hbusreq2_p & v1216afe | !hbusreq2_p & v1216afd;
assign v12150f8 = hmaster2_p & v1215438 | !hmaster2_p & v12150c4;
assign v15168ac = hburst0 & v15168a9 | !hburst0 & v15168ab;
assign v121617f = hmaster1_p & v121617e | !hmaster1_p & v121616f;
assign v1668e06 = hmaster1_p & v1668e05 | !hmaster1_p & v845542;
assign d2fc87 = hbusreq2 & d2fc86 | !hbusreq2 & v845542;
assign d30268 = hgrant1_p & f2f227 | !hgrant1_p & d3078f;
assign v1389460 = hmaster1_p & v138945e | !hmaster1_p & !v138a032;
assign v1515788 = hburst0_p & v155392f | !hburst0_p & !v893df7;
assign v14465dc = hmaster2_p & v14465d8 | !hmaster2_p & v14465db;
assign v14466a3 = hbusreq5_p & v14466a2 | !hbusreq5_p & v1446611;
assign v1552d4b = hlock0 & v1552d49 | !hlock0 & v1552d4a;
assign v14461b3 = hbusreq2_p & v144619e | !hbusreq2_p & v14461b2;
assign v15157c5 = hbusreq5_p & v15157c3 | !hbusreq5_p & !v15157c4;
assign v1446402 = hbusreq5 & v14463d5 | !hbusreq5 & v1446401;
assign v14460a1 = hbusreq2_p & v144609b | !hbusreq2_p & v14460a0;
assign d2feb7 = hbusreq4_p & d2feb6 | !hbusreq4_p & v845542;
assign v121612f = hbusreq1 & v121612e | !hbusreq1 & v845542;
assign v1446412 = hbusreq1_p & v1446403 | !hbusreq1_p & v1446406;
assign v144674d = hmaster0_p & v1446663 | !hmaster0_p & v144664a;
assign v1445e20 = hlock2 & v1445e1f | !hlock2 & v1445e19;
assign v16a1cc3 = hgrant2_p & v16a1f9b | !hgrant2_p & v16a1cc2;
assign v10d40aa = hmaster1_p & v10d40a9 | !hmaster1_p & !v10d3fe9;
assign v16a13d8 = hbusreq5 & v16a13cc | !hbusreq5 & v16a13d7;
assign v138a32e = hbusreq4_p & v1515654 | !hbusreq4_p & v15156b9;
assign v1284ce1 = hgrant2_p & v1284cc4 | !hgrant2_p & v1284ce0;
assign v155343d = hgrant1_p & v845542 | !hgrant1_p & v155343c;
assign v1516975 = jx2_p & v1516855 | !jx2_p & v1516959;
assign d2fd09 = hmaster1_p & d2fce9 | !hmaster1_p & d2fcfe;
assign d2facf = hmaster0_p & d2fea4 | !hmaster0_p & d2fe9b;
assign a662aa = hgrant4_p & a662a9 | !hgrant4_p & !v845542;
assign d2fc64 = hbusreq5_p & d2fbe4 | !hbusreq5_p & d2fc63;
assign v1215ff4 = hmaster2_p & v1215ff1 | !hmaster2_p & v845542;
assign a65393 = hburst0 & v88d3e4 | !hburst0 & a65392;
assign v16a1bcf = hmaster2_p & v16a1bcb | !hmaster2_p & v16a208a;
assign v14466b9 = hgrant2_p & v1446681 | !hgrant2_p & v14466b8;
assign v12acfe1 = hmaster1_p & v12acfc5 | !hmaster1_p & v12acfdb;
assign d30758 = hbusreq2_p & d30757 | !hbusreq2_p & d30756;
assign d2fb31 = hbusreq2 & d2fb2d | !hbusreq2 & d2fb30;
assign v10d40c8 = hmaster0_p & v10d4083 | !hmaster0_p & v10d4064;
assign f2f347 = hgrant1_p & v845570 | !hgrant1_p & !f2f346;
assign v1405b63 = decide_p & v1405ab4 | !decide_p & v1405b62;
assign v121624c = hmaster1_p & v1216209 | !hmaster1_p & !v121624b;
assign d30888 = hgrant1_p & v84554c | !hgrant1_p & d30887;
assign v1552962 = hgrant3_p & v1553106 | !hgrant3_p & v1552961;
assign v1445baa = hmaster0_p & v14464a5 | !hmaster0_p & v845542;
assign f2f53a = hmaster0_p & f2f539 | !hmaster0_p & f2f229;
assign d2fec4 = hmaster2_p & v84555a | !hmaster2_p & d2fec3;
assign v1405aba = hlock3_p & v1405ab4 | !hlock3_p & v1405ab9;
assign d307ae = hbusreq4 & d306d4 | !hbusreq4 & v845542;
assign v16a1d7e = hgrant2_p & v845542 | !hgrant2_p & v16a1d7c;
assign v1668ce5 = hbusreq0 & v1668cd2 | !hbusreq0 & v1668ce4;
assign d307fc = hgrant5_p & d30708 | !hgrant5_p & !d307fa;
assign v12acfbf = hmaster1_p & v12acfbe | !hmaster1_p & !v12ad525;
assign v1405a98 = hmaster1_p & v1405a97 | !hmaster1_p & !v1405a94;
assign v1405930 = hbusreq5_p & v14058ba | !hbusreq5_p & v140592f;
assign v15168aa = stateA1_p & d30714 | !stateA1_p & a658a3;
assign v16a13f8 = hmaster1_p & v16a13f7 | !hmaster1_p & v16a1d7a;
assign d3015c = hgrant2_p & d30113 | !hgrant2_p & !d3015b;
assign v14058a5 = hbusreq5_p & v14058a1 | !hbusreq5_p & v14058a4;
assign v1216adf = hbusreq4_p & v1216ade | !hbusreq4_p & !v845542;
assign v144576b = hbusreq2_p & v1445767 | !hbusreq2_p & v144576a;
assign v14058fb = hgrant0_p & v140583f | !hgrant0_p & v14463b1;
assign a65412 = hbusreq2 & a65408 | !hbusreq2 & a65410;
assign v16a19b0 = hgrant5_p & v845542 | !hgrant5_p & v16a19af;
assign v1215c75 = hbusreq2_p & v1215c6c | !hbusreq2_p & !v1215c74;
assign v16a1ab8 = hbusreq3 & v16a224a | !hbusreq3 & v16a1ab7;
assign v1446683 = hbusreq2_p & v1446632 | !hbusreq2_p & v1446682;
assign v1445ae1 = hbusreq3 & v1445adf | !hbusreq3 & v1445ae0;
assign d2f997 = hmaster1_p & d2fec8 | !hmaster1_p & d2f995;
assign v1445aa0 = hbusreq2_p & v1445a9d | !hbusreq2_p & v1445a9f;
assign v1445f85 = hmaster2_p & v144639c | !hmaster2_p & v14463a5;
assign d307e1 = hgrant4_p & d307c7 | !hgrant4_p & v845542;
assign v12162f4 = hmaster0_p & v12162f1 | !hmaster0_p & v12162f3;
assign v1216aba = hbusreq4_p & v1216ab8 | !hbusreq4_p & v1216ab9;
assign v1214cca = hgrant1_p & v1214cc8 | !hgrant1_p & v1214cc9;
assign v16a1db7 = hbusreq2 & v16a1db4 | !hbusreq2 & !v16a1db6;
assign d30749 = hlock2_p & d30746 | !hlock2_p & d30748;
assign v1668cad = hgrant2_p & v1668cab | !hgrant2_p & v1668cac;
assign v1214bc7 = hbusreq2_p & v1214bc6 | !hbusreq2_p & v1214bc5;
assign v14058af = hmaster2_p & v14058a9 | !hmaster2_p & v14058ae;
assign v1668d70 = hbusreq4_p & v1668d6e | !hbusreq4_p & !v1668d6f;
assign v15168b3 = hmaster1_p & v15168b2 | !hmaster1_p & v845542;
assign v1668d43 = hmaster2_p & a6585c | !hmaster2_p & v1668d18;
assign stateG3_1 = !v1552990;
assign d2fb9c = hbusreq0 & d2fb9b | !hbusreq0 & v845542;
assign v12ad565 = hbusreq0 & v12ad564 | !hbusreq0 & !v845542;
assign a658bf = hbusreq1 & a658b6 | !hbusreq1 & !a658be;
assign d306d3 = hmaster2_p & d306d0 | !hmaster2_p & v845542;
assign v12160cf = hlock3_p & v12160a0 | !hlock3_p & v12160ce;
assign v134d520 = hgrant2_p & v134d364 | !hgrant2_p & v134d51f;
assign v134d4a6 = hlock2 & v134d3b5 | !hlock2 & v134d49c;
assign v11e5949 = hmaster2_p & v11e593a | !hmaster2_p & !v845542;
assign v1216592 = hmastlock_p & v1216591 | !hmastlock_p & !v845542;
assign v16a12e7 = hlock0_p & v16a206a | !hlock0_p & !v16a12e6;
assign v12160a2 = hmaster1_p & v12160a1 | !hmaster1_p & v121605d;
assign v1216a95 = hbusreq5_p & v1216a94 | !hbusreq5_p & v845542;
assign v14453be = hbusreq2 & v14453ba | !hbusreq2 & v14453bd;
assign v16a1966 = hgrant5_p & v845542 | !hgrant5_p & !v16a1958;
assign d308cc = hgrant2_p & d3085f | !hgrant2_p & d308c8;
assign v1215437 = hlock4_p & v1215436 | !hlock4_p & !v845559;
assign v12166de = hgrant1_p & v12164de | !hgrant1_p & v12166dd;
assign v138a364 = hbusreq2_p & v138a361 | !hbusreq2_p & v138a363;
assign v14463a2 = hbusreq1 & v14463a0 | !hbusreq1 & v14463a1;
assign v15157e2 = hgrant5_p & v845542 | !hgrant5_p & !v1515737;
assign d30664 = hbusreq5_p & d3065f | !hbusreq5_p & d30663;
assign v14058c2 = hgrant1_p & v140583d | !hgrant1_p & v14058c1;
assign v16a138f = hmaster1_p & v16a1383 | !hmaster1_p & v16a1f96;
assign v1445441 = hbusreq2_p & v1445440 | !hbusreq2_p & v1445bab;
assign v134d201 = hbusreq5_p & v134d200 | !hbusreq5_p & v134d1fd;
assign v1445356 = hmaster1_p & v1445355 | !hmaster1_p & v14458fd;
assign v16a188e = hbusreq2 & v16a188c | !hbusreq2 & v16a188d;
assign v12ad586 = hbusreq2_p & v12ad584 | !hbusreq2_p & v12ad585;
assign a65aeb = hgrant1_p & v845542 | !hgrant1_p & !a65aea;
assign v1214f53 = hbusreq2 & v1214f51 | !hbusreq2 & v12164e7;
assign v1445f18 = hlock2 & v1445edb | !hlock2 & v1445f17;
assign v10d428d = hgrant5_p & v10d3fdc | !hgrant5_p & v10d428c;
assign v12ae1f3 = hgrant5_p & v845542 | !hgrant5_p & v12ae1f2;
assign v12ad51a = hbusreq1 & v12ad515 | !hbusreq1 & !v12ad519;
assign v1668c8e = hbusreq2_p & v1668c88 | !hbusreq2_p & v1668c8d;
assign v1445b08 = hbusreq2_p & v1445b02 | !hbusreq2_p & v1445b07;
assign d300d5 = hbusreq1 & d2fe7d | !hbusreq1 & !d2fe93;
assign hgrant4 = !a64719;
assign v138a3e7 = hlock5_p & v138a3e6 | !hlock5_p & !v1515796;
assign f2f411 = hbusreq2 & f2f40d | !hbusreq2 & f2f410;
assign v1445768 = hmaster1_p & v1445f49 | !hmaster1_p & v1445dd1;
assign v1216228 = hmaster0_p & v12160d5 | !hmaster0_p & v1216227;
assign d8073a = hmastlock_p & d80739 | !hmastlock_p & !v845542;
assign v1214c5f = hgrant5_p & v1215367 | !hgrant5_p & v1214c5d;
assign a653cd = hbusreq4_p & a653cc | !hbusreq4_p & v845542;
assign v1445e5a = hlock1 & v1446606 | !hlock1 & v1445e59;
assign d2fecc = hbusreq2_p & d2fecb | !hbusreq2_p & d2feca;
assign v151560f = hmaster2_p & a65851 | !hmaster2_p & v151560e;
assign v138a3fb = hbusreq2_p & v138a3f6 | !hbusreq2_p & !v138a3fa;
assign v1215c74 = hgrant2_p & v1215c39 | !hgrant2_p & !v1215c73;
assign v16a266b = hmaster2_p & v845542 | !hmaster2_p & v84554d;
assign v1445eea = hmaster2_p & v1445ec8 | !hmaster2_p & v1445e6c;
assign v12ad61e = hmaster0_p & v12ad602 | !hmaster0_p & v12ad61d;
assign v1668d3f = hgrant5_p & v10d3fd8 | !hgrant5_p & v1668d3d;
assign v144582e = hmaster1_p & v1445803 | !hmaster1_p & v1445e28;
assign v121610e = hbusreq1 & v121610d | !hbusreq1 & v845542;
assign v134cd7f = hlock0 & v134cd7e | !hlock0 & v134cd7d;
assign v14463bf = hbusreq5_p & v14463be | !hbusreq5_p & v14463bc;
assign v144667d = hbusreq5_p & v1446678 | !hbusreq5_p & v1446636;
assign v14463cb = hmaster1_p & v14463ca | !hmaster1_p & v14463c2;
assign v121533c = hgrant2_p & v1215324 | !hgrant2_p & v121533b;
assign v1214ecf = hmaster2_p & v121652b | !hmaster2_p & v845542;
assign v1215c6c = hgrant2_p & v1215bed | !hgrant2_p & v1215c6b;
assign v14458a5 = hbusreq0 & v14458a1 | !hbusreq0 & v14458a4;
assign v14453b1 = hbusreq2 & v14453ad | !hbusreq2 & v14453b0;
assign v16a1e5b = hlock0_p & v845542 | !hlock0_p & v16a1e5a;
assign v1215087 = hmaster1_p & v121506e | !hmaster1_p & !v121507b;
assign v12afe58 = hgrant5_p & v845542 | !hgrant5_p & v12afe57;
assign v1445eb1 = hmaster0_p & v1446404 | !hmaster0_p & v1445eb0;
assign v15533a9 = hbusreq0 & v15533a8 | !hbusreq0 & v15533a7;
assign v1445aab = hlock5 & v1445a69 | !hlock5 & v1445aaa;
assign v1215719 = hbusreq1 & v1215b99 | !hbusreq1 & v845542;
assign v16a208d = hbusreq0 & v16a207b | !hbusreq0 & v16a208c;
assign v1214e67 = hbusreq3 & v1214e50 | !hbusreq3 & v1214e66;
assign v1389efc = decide_p & v1389d76 | !decide_p & v138a406;
assign v1216532 = hlock5_p & v1216530 | !hlock5_p & v1216531;
assign v134d4ce = hgrant5_p & v134d281 | !hgrant5_p & v134d4cd;
assign bf1f82 = hgrant1_p & bf1f52 | !hgrant1_p & bf1f81;
assign v12ad4be = hbusreq4_p & v12adf60 | !hbusreq4_p & !v845542;
assign v1515801 = hmaster0_p & v1515800 | !hmaster0_p & v15157d0;
assign v1445402 = decide_p & v14453f1 | !decide_p & v1445401;
assign v14453a1 = hlock3 & v144538c | !hlock3 & v14453a0;
assign v16a1e69 = hmaster1_p & v16a1e68 | !hmaster1_p & v16a2672;
assign v134d269 = hlock2 & v134d264 | !hlock2 & v134d268;
assign v12162b8 = hmaster1_p & v12162b7 | !hmaster1_p & v1216041;
assign a656b1 = hbusreq3 & a656a4 | !hbusreq3 & a656b0;
assign v144644c = hlock2 & v1446443 | !hlock2 & v144644b;
assign v12ad506 = hlock0_p & v151563e | !hlock0_p & v845542;
assign v14459b4 = hbusreq4 & v14459a7 | !hbusreq4 & v14459b3;
assign v1445dee = hbusreq1 & v1445deb | !hbusreq1 & v1445ded;
assign v1405846 = hmaster2_p & v14463b1 | !hmaster2_p & v1405845;
assign v15160f9 = hmaster0_p & v845542 | !hmaster0_p & v16693a7;
assign v1445e5d = hbusreq4 & v1446406 | !hbusreq4 & v1446409;
assign v16a2084 = hgrant4_p & v845559 | !hgrant4_p & !v16a2083;
assign v151573e = hbusreq1 & a6585c | !hbusreq1 & !v1515627;
assign v1216af3 = hlock0_p & v1216adc | !hlock0_p & v845542;
assign v12af9d6 = hbusreq0 & v12af9ce | !hbusreq0 & v12af9d5;
assign v1445dc4 = hmaster0_p & v144639c | !hmaster0_p & v1445da7;
assign v1445a97 = hbusreq5_p & v14459d1 | !hbusreq5_p & v1445a96;
assign f2f2ad = hmaster2_p & f2f2a8 | !hmaster2_p & v845542;
assign d30215 = hlock5_p & d30213 | !hlock5_p & d30214;
assign v12162c2 = hmaster0_p & v12160e2 | !hmaster0_p & v1216227;
assign bf1f9b = hgrant1_p & f2f227 | !hgrant1_p & bf1f9a;
assign v1284d55 = hmaster0_p & v1405859 | !hmaster0_p & v1284d00;
assign v16a13f5 = hgrant5_p & v845542 | !hgrant5_p & !v16a13e2;
assign v1445eff = hlock2 & v1445edb | !hlock2 & v1445efe;
assign v10d4090 = hmaster1_p & v10d408f | !hmaster1_p & !v10d3fe9;
assign v1445ff2 = hmaster1_p & v1445ff1 | !hmaster1_p & v1445fef;
assign v138a39e = hmaster1_p & v138a39d | !hmaster1_p & v138a341;
assign v1515709 = hbusreq2 & v1515708 | !hbusreq2 & v15167ed;
assign v134d4eb = hmaster2_p & v845542 | !hmaster2_p & v134d4ea;
assign v138a093 = hbusreq3_p & v138a05b | !hbusreq3_p & v138a092;
assign v12afa34 = hgrant3_p & v12af9b9 | !hgrant3_p & v12afa33;
assign v1214c90 = hgrant5_p & v845542 | !hgrant5_p & v1214c6f;
assign v12150b5 = hmaster0_p & v1215773 | !hmaster0_p & v1215b9a;
assign v14466eb = hlock3 & v14466e1 | !hlock3 & v14466ea;
assign v16a1af6 = stateA1_p & v84557e | !stateA1_p & !v16a1af5;
assign v1405ab7 = hmaster1_p & v1405ab0 | !hmaster1_p & v1405aae;
assign v1445dc9 = hlock3 & v1445dc6 | !hlock3 & v1445dc8;
assign v1214d03 = hbusreq0 & v1214d02 | !hbusreq0 & v845542;
assign v1668dd8 = hgrant5_p & v845542 | !hgrant5_p & !v1668d98;
assign v1284cab = hmaster1_p & v1284caa | !hmaster1_p & v1284ca7;
assign v1668d21 = hbusreq1 & a65851 | !hbusreq1 & v845570;
assign v1552d81 = hmaster2_p & v1552d7c | !hmaster2_p & v845542;
assign v12ad026 = hbusreq0 & v12ad025 | !hbusreq0 & v12afa0a;
assign a653d3 = hgrant5_p & a6586d | !hgrant5_p & a653d1;
assign v1552d66 = hlock2 & v155341e | !hlock2 & v1552d62;
assign v144634f = hmaster1_p & v14462e8 | !hmaster1_p & v1446290;
assign v144646e = locked_p & v144646d | !locked_p & v845542;
assign a65692 = hmaster1_p & a65691 | !hmaster1_p & a658e5;
assign v121632b = hmaster1_p & v121630d | !hmaster1_p & v121631b;
assign v1214d22 = hgrant2_p & v1214d0a | !hgrant2_p & v1214d21;
assign v1214f15 = hmaster0_p & v1214f14 | !hmaster0_p & v1214ef9;
assign v12150d0 = hbusreq0 & v12153e5 | !hbusreq0 & v12150cf;
assign v12ad024 = hgrant5_p & v845542 | !hgrant5_p & !v12ad005;
assign v15534d9 = hbusreq0 & v15534d8 | !hbusreq0 & v15534d2;
assign v134d27a = hmaster1_p & v134d279 | !hmaster1_p & v845542;
assign v1515644 = hbusreq3 & v151563d | !hbusreq3 & !v1515643;
assign v138a478 = hmaster0_p & v138a304 | !hmaster0_p & v138a2f8;
assign a6627f = hmaster1_p & v845542 | !hmaster1_p & a6627e;
assign v1216173 = hmaster0_p & v121601e | !hmaster0_p & v1216172;
assign v12162f9 = hlock2_p & v12162f5 | !hlock2_p & v12162f8;
assign v144587d = stateG10_5_p & v144587c | !stateG10_5_p & !v144587b;
assign v1215032 = hbusreq4 & v12166ce | !hbusreq4 & !v845542;
assign d301d2 = hmaster2_p & d301d1 | !hmaster2_p & v845542;
assign d2fb6f = hlock1_p & d2fb6e | !hlock1_p & v84554a;
assign d308a5 = hbusreq1_p & d307e3 | !hbusreq1_p & d306ae;
assign v1214f56 = hgrant2_p & v845542 | !hgrant2_p & v1214f55;
assign v16a1ae6 = hgrant5_p & v845542 | !hgrant5_p & !v16a1adc;
assign d306b4 = hbusreq5_p & d3066a | !hbusreq5_p & !d306b2;
assign v1214f68 = hmaster1_p & v1214f67 | !hmaster1_p & v1215d2b;
assign v12150be = hmaster1_p & v12150bd | !hmaster1_p & v12153bf;
assign v1445873 = hmaster2_p & v144639c | !hmaster2_p & v1445872;
assign v144547c = hbusreq2_p & v144547a | !hbusreq2_p & v1445bba;
assign d2fb3f = hbusreq2_p & d2feff | !hbusreq2_p & d2fb3d;
assign v121544e = hmaster1_p & v12153ee | !hmaster1_p & v121540f;
assign v1214fe3 = hgrant0_p & v12160f2 | !hgrant0_p & !v845559;
assign v138a3ae = hbusreq3 & v138a3a0 | !hbusreq3 & v138a3ad;
assign v16a1e4f = hbusreq2 & v16a1e4c | !hbusreq2 & v16a1e4e;
assign v1668d7f = hmaster2_p & v1668d63 | !hmaster2_p & a653c4;
assign v16a224b = hmaster0_p & v16a2246 | !hmaster0_p & v16a2240;
assign d301fa = hmaster2_p & v845542 | !hmaster2_p & d301f9;
assign v1446221 = hmaster1_p & v144621d | !hmaster1_p & v1446219;
assign v14459f9 = hlock1 & v14459f8 | !hlock1 & v14459c8;
assign v1446101 = hbusreq3 & v14460ff | !hbusreq3 & v1446100;
assign v13895a4 = hbusreq5 & v138953c | !hbusreq5 & v13895a3;
assign v1214ef9 = hbusreq0 & v1214ef6 | !hbusreq0 & v1214ef8;
assign d30200 = hgrant5_p & d301f1 | !hgrant5_p & d301ff;
assign v134d385 = hgrant4_p & v845542 | !hgrant4_p & v134d384;
assign v1516107 = hready_p & v845542 | !hready_p & v1516106;
assign v155350f = hmaster1_p & v155350e | !hmaster1_p & v845542;
assign v1446161 = hmaster0_p & v1445fe3 | !hmaster0_p & v144639c;
assign v134cf41 = hgrant3_p & v134cee7 | !hgrant3_p & v134cf40;
assign v1668d28 = hgrant1_p & v1668d23 | !hgrant1_p & v1668d27;
assign v144545d = hbusreq3 & v144545b | !hbusreq3 & v144545c;
assign v16a1d2c = hmaster1_p & v16a2234 | !hmaster1_p & !v16a2672;
assign d2fc0d = hgrant5_p & d2fc0c | !hgrant5_p & d2fbe1;
assign d2fbf7 = hmaster2_p & d2fbf6 | !hmaster2_p & v845542;
assign v1214c9c = hmaster1_p & v1214c9b | !hmaster1_p & v845542;
assign v1216017 = hbusreq1_p & v1216016 | !hbusreq1_p & v845542;
assign v12ad5d0 = hbusreq1 & v12ad4da | !hbusreq1 & v12ad4e4;
assign v1553157 = hmaster1_p & v1553150 | !hmaster1_p & v155314e;
assign v1214f16 = hmaster1_p & v1214eef | !hmaster1_p & v1214f15;
assign v1216219 = hbusreq1 & v12166dd | !hbusreq1 & v845542;
assign v134d240 = hbusreq2_p & v134d23f | !hbusreq2_p & v134d23e;
assign v14461ec = hbusreq2 & v14461e8 | !hbusreq2 & v14461eb;
assign v10d404b = hmaster2_p & v10d4043 | !hmaster2_p & v10d404a;
assign v1405a8b = hmaster0_p & v1405a89 | !hmaster0_p & v1405a8a;
assign v1445a8b = hgrant2_p & v1445a89 | !hgrant2_p & v1445a8a;
assign v1445da4 = hmaster0_p & v1445d95 | !hmaster0_p & v1445da3;
assign v14463c3 = hmaster1_p & v144639c | !hmaster1_p & v14463c2;
assign v10d42a5 = hgrant5_p & v10d3feb | !hgrant5_p & v10d42a4;
assign v1216248 = hmaster2_p & v1216231 | !hmaster2_p & !v845542;
assign v1389411 = jx2_p & v138932d | !jx2_p & v13893b7;
assign a6569c = hmaster1_p & a65465 | !hmaster1_p & !a65916;
assign v1445a6a = hbusreq0 & v1445a4d | !hbusreq0 & v1445a36;
assign d2fb1f = hbusreq0 & d2fb1c | !hbusreq0 & d2fb1e;
assign v16a143f = hbusreq2 & v16a143d | !hbusreq2 & !v16a143e;
assign acd334 = stateG3_1_p & v845542 | !stateG3_1_p & v84556c;
assign v14453ed = hlock3 & v14453e4 | !hlock3 & v14453ec;
assign v14457bc = hbusreq2_p & v14457ba | !hbusreq2_p & v14457bb;
assign v1446632 = hgrant2_p & v14465ab | !hgrant2_p & v1446631;
assign v1215c11 = hlock5_p & v1215c0f | !hlock5_p & v1215c10;
assign v10d4268 = hlock0_p & v10d4267 | !hlock0_p & v10d3fd4;
assign v14466e0 = hlock2 & v14466d3 | !hlock2 & v14466de;
assign v144664b = hmaster0_p & v14465b8 | !hmaster0_p & v144664a;
assign v1214c71 = hgrant5_p & v121536a | !hgrant5_p & v1214c6f;
assign v134d4c6 = hgrant3_p & v134d4c3 | !hgrant3_p & v134d4c5;
assign v10d4081 = hmaster1_p & v10d4080 | !hmaster1_p & v10d3fe9;
assign d2fae6 = hbusreq4_p & d300ca | !hbusreq4_p & d306a3;
assign v134d28a = hlock4_p & v134d1dd | !hlock4_p & v845542;
assign v12ad1b3 = hgrant3_p & v12ad0cc | !hgrant3_p & v12ad1b1;
assign v12af7e1 = hbusreq2_p & v845542 | !hbusreq2_p & v12af73f;
assign v1446184 = hmaster0_p & v1446092 | !hmaster0_p & v144603f;
assign d2fb89 = hbusreq2_p & d2fb88 | !hbusreq2_p & d2fb80;
assign v1284d5f = hgrant2_p & v1284d5c | !hgrant2_p & v1284d5e;
assign v1284cb0 = hbusreq2_p & v1284cac | !hbusreq2_p & v1284caf;
assign v1214ef4 = hbusreq5_p & v1214ef3 | !hbusreq5_p & v1216547;
assign v1215d46 = hbusreq3 & v1215d45 | !hbusreq3 & v845542;
assign v1553447 = hgrant3_p & v1553437 | !hgrant3_p & v1553446;
assign v16a19a6 = hbusreq4 & v16a223a | !hbusreq4 & !v845542;
assign d2f99c = hbusreq5_p & d2fec8 | !hbusreq5_p & d2f99b;
assign v1515654 = hmastlock_p & v1515653 | !hmastlock_p & v845542;
assign v16a223a = locked_p & v845542 | !locked_p & !v16a2239;
assign v1445853 = hmaster1_p & v1445805 | !hmaster1_p & v1445f09;
assign v1214fba = hgrant4_p & v845542 | !hgrant4_p & v1214fb9;
assign v1215bf0 = hbusreq1_p & v1215fe9 | !hbusreq1_p & !v1215bef;
assign v1214c32 = hmaster2_p & d2fbe5 | !hmaster2_p & v1214c31;
assign v1668c4b = hmaster0_p & v1668c4a | !hmaster0_p & v845542;
assign v1284d31 = decide_p & v140590a | !decide_p & v1284d30;
assign v16a1972 = hbusreq0 & v16a207a | !hbusreq0 & v16a1971;
assign v16a1d11 = hbusreq3 & v16a1b66 | !hbusreq3 & !v16a1f9c;
assign stateA1 = !v10d4305;
assign v1668c60 = hmaster2_p & a658ad | !hmaster2_p & a658b5;
assign v1214dd7 = hmaster1_p & v1214dd6 | !hmaster1_p & v845542;
assign f2f21b = hlock1_p & f2f21a | !hlock1_p & !v845542;
assign v1215442 = hbusreq5 & v121540b | !hbusreq5 & v1215441;
assign v134cee4 = hlock5 & v134d276 | !hlock5 & v134cee3;
assign d2fc16 = hgrant2_p & d2fc08 | !hgrant2_p & d2fc12;
assign v1445884 = hbusreq1 & v1445883 | !hbusreq1 & v1445870;
assign v134d284 = hgrant1_p & v134d283 | !hgrant1_p & v845542;
assign bf1f8e = hbusreq4_p & a65382 | !hbusreq4_p & bf1f8d;
assign v1215ca1 = hbusreq1 & v1215fec | !hbusreq1 & v1216014;
assign v1668c59 = jx2_p & v1668c3a | !jx2_p & v1668c58;
assign d30776 = hlock2_p & d30775 | !hlock2_p & d30772;
assign v1214d88 = hgrant2_p & v121657d | !hgrant2_p & v1214d84;
assign v1284cd8 = hgrant1_p & v1405849 | !hgrant1_p & !v1284cd7;
assign v1215d47 = decide_p & v1215d0d | !decide_p & v1215d46;
assign v144662e = hbusreq0 & v1446623 | !hbusreq0 & v144662d;
assign v1445e0e = hmaster1_p & v1445e0d | !hmaster1_p & v1445e07;
assign v134cec9 = hlock3 & v134d3b5 | !hlock3 & v134cec8;
assign v12acfed = hbusreq3 & v12acfe3 | !hbusreq3 & v12acfec;
assign v10d42d3 = hmaster1_p & v10d42a5 | !hmaster1_p & !v10d42a1;
assign v1668c81 = hmaster1_p & v1668c75 | !hmaster1_p & v1668c72;
assign v12afe5d = hmaster2_p & v12afe46 | !hmaster2_p & v12afe5c;
assign v1515837 = hmaster2_p & v151572a | !hmaster2_p & v151575a;
assign v138a302 = hmaster1_p & v138a2fb | !hmaster1_p & v138a301;
assign a6627c = hmaster2_p & a6627b | !hmaster2_p & !v845542;
assign d2fc6e = hmaster1_p & d2fc5a | !hmaster1_p & d2fc6d;
assign v134ce6f = decide_p & v134d3fa | !decide_p & v134ce6e;
assign v1668db6 = hgrant5_p & v1668da6 | !hgrant5_p & v1668d30;
assign v1446083 = hmaster1_p & v1446082 | !hmaster1_p & v1446073;
assign d3088a = hgrant1_p & v84554c | !hgrant1_p & d30889;
assign v13891a7 = decide_p & v13891a6 | !decide_p & v845542;
assign v14058f2 = hgrant0_p & v14058f1 | !hgrant0_p & !v1405844;
assign a6541d = hbusreq5_p & a65419 | !hbusreq5_p & !a6541b;
assign v144649e = hmaster2_p & v1446493 | !hmaster2_p & v144649d;
assign v140588e = locked_p & v140588d | !locked_p & !v140583c;
assign d8079e = hgrant2_p & d80768 | !hgrant2_p & d8079d;
assign d300f5 = hbusreq5_p & d300f1 | !hbusreq5_p & d300f4;
assign v10d3fe3 = hmaster2_p & v10d3fe0 | !hmaster2_p & v10d3fe1;
assign v1446645 = hgrant1_p & v1446407 | !hgrant1_p & v14465ce;
assign v1215da2 = hbusreq2_p & v1215d9d | !hbusreq2_p & v1215da1;
assign d30288 = hmaster0_p & v1668da6 | !hmaster0_p & v1668c1d;
assign v138a3e0 = hmaster0_p & v138a3d8 | !hmaster0_p & v138a3df;
assign v16a1c9d = hgrant2_p & v16a2058 | !hgrant2_p & v16a1c9c;
assign v14458f3 = hbusreq0_p & v14458f2 | !hbusreq0_p & v1446406;
assign v1216308 = hbusreq2_p & v12162f9 | !hbusreq2_p & v1216307;
assign d80764 = hmaster1_p & d80763 | !hmaster1_p & !v845542;
assign v1214d26 = hbusreq2 & v1214d23 | !hbusreq2 & v1214d25;
assign v16a1e09 = hbusreq2 & v16a1e07 | !hbusreq2 & !v16a1e08;
assign d2fad2 = hmaster0_p & d3011e | !hmaster0_p & d300d3;
assign d2fb3c = hmaster0_p & d2fb36 | !hmaster0_p & d2fb3b;
assign v12ad673 = hlock0_p & v12ad513 | !hlock0_p & v12ad672;
assign d2fe84 = hbusreq4_p & d2fe83 | !hbusreq4_p & v845542;
assign d2fbf0 = hgrant5_p & v84554a | !hgrant5_p & d2fbef;
assign v1214cd4 = hgrant1_p & v1215385 | !hgrant1_p & v1214cd3;
assign v1405ad3 = locked_p & v1405aa2 | !locked_p & v1405a86;
assign v1214c8d = hgrant5_p & v16a2243 | !hgrant5_p & v1214c62;
assign v15534d0 = hgrant1_p & v845542 | !hgrant1_p & v15534cf;
assign v12ad674 = hbusreq4_p & v12ad514 | !hbusreq4_p & v12ad673;
assign v138a39d = hmaster0_p & v138a394 | !hmaster0_p & v138a354;
assign v11ac67a = decide_p & v11ac602 | !decide_p & v84554c;
assign v1515790 = locked_p & v151578f | !locked_p & v845542;
assign v1214dd1 = hlock2_p & v1214dce | !hlock2_p & v1214dd0;
assign v12150a4 = hgrant5_p & v121546e | !hgrant5_p & v12150a3;
assign v12ad67b = hbusreq0 & v12ad67a | !hbusreq0 & !v12af7f7;
assign v12ad630 = hgrant3_p & v12ad595 | !hgrant3_p & v12ad62f;
assign v16a1846 = hmaster0_p & v16a1842 | !hmaster0_p & v16a1840;
assign v12ad4f2 = hbusreq0 & v12ad4f1 | !hbusreq0 & v845542;
assign v12153da = hbusreq1 & v12153d3 | !hbusreq1 & v12153d9;
assign v16a1394 = hmaster1_p & v16a138a | !hmaster1_p & v16a1f96;
assign v1216a5e = stateA1_p & v845542 | !stateA1_p & v1216a5d;
assign v144551f = hmaster1_p & v14454e8 | !hmaster1_p & v1446290;
assign v12ad5d7 = hlock0_p & v1515764 | !hlock0_p & v845542;
assign d3024b = hbusreq5_p & d30249 | !hbusreq5_p & d3024a;
assign v12167af = hmaster0_p & v12164e3 | !hmaster0_p & v12164d5;
assign v1515605 = decide_p & v15155ee | !decide_p & !v845576;
assign v1445eab = hmaster1_p & v14465b7 | !hmaster1_p & v1445eaa;
assign v14458e6 = hmaster2_p & v1446403 | !hmaster2_p & v14458e5;
assign v1668c20 = hmaster0_p & v1668c1e | !hmaster0_p & v1668c1f;
assign v12aeb85 = hready_p & v845542 | !hready_p & v12aeb84;
assign v1405b0f = decide_p & v1405afb | !decide_p & v1405b0e;
assign v1214e7d = hbusreq2_p & v1214e7c | !hbusreq2_p & v845542;
assign a658ab = hburst1 & a658aa | !hburst1 & v845542;
assign v16a1f96 = hmaster0_p & v16a1f95 | !hmaster0_p & !v16a2671;
assign v1668c83 = hbusreq2_p & v1668c73 | !hbusreq2_p & v1668c82;
assign d308ba = hgrant5_p & d30654 | !hgrant5_p & d30892;
assign v121570c = hbusreq1 & v1215b76 | !hbusreq1 & v845542;
assign v12ad576 = hbusreq2_p & v12ad573 | !hbusreq2_p & v12ad575;
assign v12160c2 = hbusreq2 & v12160bd | !hbusreq2 & v12160c1;
assign v134d1eb = hlock4 & v134d1e8 | !hlock4 & v134d1ea;
assign v14458af = hmaster0_p & v144587f | !hmaster0_p & v1445895;
assign v1216076 = hbusreq2_p & v1216075 | !hbusreq2_p & v1216074;
assign v16a1bde = hgrant2_p & v845542 | !hgrant2_p & !v16a1bdc;
assign v14466fe = hmaster0_p & v1446638 | !hmaster0_p & v144643e;
assign v12160ca = hlock2_p & v12160c8 | !hlock2_p & v12160c9;
assign v1405934 = hmaster0_p & v14058df | !hmaster0_p & v14058c4;
assign a65af4 = hbusreq2_p & a65adb | !hbusreq2_p & a65af3;
assign v10d4029 = hmaster2_p & v10d3fd9 | !hmaster2_p & !v10d3fe1;
assign v1445b6c = hbusreq2_p & v1445b64 | !hbusreq2_p & v1445b6b;
assign v16a1402 = hbusreq2 & v16a1401 | !hbusreq2 & !v16a1d55;
assign v14459db = hgrant1_p & v14459d6 | !hgrant1_p & v14459da;
assign v16a19c1 = hmaster1_p & v16a19ac | !hmaster1_p & v16a1f96;
assign v1445915 = hlock3 & v1445912 | !hlock3 & v1445914;
assign d307a4 = hlock5_p & d307a2 | !hlock5_p & !d307a3;
assign v1405ac0 = hbusreq1_p & v845542 | !hbusreq1_p & v1405abf;
assign v121538e = decide_p & v1215374 | !decide_p & v121538d;
assign v1515772 = hgrant0_p & v1515771 | !hgrant0_p & v1515614;
assign v1445fdb = hbusreq1_p & v1446432 | !hbusreq1_p & v1446429;
assign v143fd7c = hready_p & v143fd7b | !hready_p & v845566;
assign d30163 = decide_p & d30162 | !decide_p & v845570;
assign v12160ed = hbusreq4_p & v12160eb | !hbusreq4_p & !v12160ec;
assign a662be = hbusreq3_p & a662a7 | !hbusreq3_p & a662bd;
assign v16a1e8c = hbusreq4_p & v845542 | !hbusreq4_p & v16a1e8b;
assign v15157d5 = hbusreq2_p & v15157d4 | !hbusreq2_p & !v845542;
assign v12152eb = hgrant2_p & v12152e8 | !hgrant2_p & v12152ea;
assign d2fc8d = hbusreq3 & d2fc87 | !hbusreq3 & d2fc8c;
assign v16a1ceb = hgrant1_p & v84554d | !hgrant1_p & v16a1cea;
assign v1445fc1 = hmaster1_p & v1445faa | !hmaster1_p & v1445fbd;
assign v12ad643 = hbusreq0 & v12ad4fa | !hbusreq0 & v12af73f;
assign v14465bb = locked_p & v144639c | !locked_p & !v14463b1;
assign v16a1dd5 = hbusreq2 & v16a1f97 | !hbusreq2 & v16a1dd4;
assign v1215313 = hmaster0_p & v1215bac | !hmaster0_p & v1215baf;
assign v121651c = hmaster1_p & v121651b | !hmaster1_p & v1216a71;
assign v16a1dbe = hmaster1_p & v9109e4 | !hmaster1_p & v16a2672;
assign v1445ed6 = hmaster0_p & v1446404 | !hmaster0_p & v1445eae;
assign v11e597b = hgrant5_p & v845542 | !hgrant5_p & v11e597a;
assign a656a3 = hbusreq2_p & a656a1 | !hbusreq2_p & a656a2;
assign f2eda2 = hgrant3_p & f2ed91 | !hgrant3_p & f2eda1;
assign v1214d2b = hmaster0_p & v1214d27 | !hmaster0_p & v1214d2a;
assign v10d4304 = jx1_p & v10d42e1 | !jx1_p & v10d40de;
assign d300fd = hgrant4_p & v845542 | !hgrant4_p & d300fc;
assign d2fbb2 = hmaster1_p & d2fb7e | !hmaster1_p & d2fb7b;
assign v134cea4 = hbusreq2_p & v134cea3 | !hbusreq2_p & v134d23e;
assign v16a12f2 = hgrant5_p & v845542 | !hgrant5_p & !v16a12eb;
assign v1446603 = hgrant1_p & v1446425 | !hgrant1_p & v1446602;
assign v16a13ea = hbusreq2 & v16a13e9 | !hbusreq2 & !v16a1d55;
assign v1445e49 = hgrant5_p & v845542 | !hgrant5_p & v1445e48;
assign v14457e0 = hgrant2_p & v14457de | !hgrant2_p & v14457df;
assign v134d49f = hbusreq0 & v134d3aa | !hbusreq0 & v134d274;
assign v1445d8a = hmaster2_p & v14463b1 | !hmaster2_p & !v1445d85;
assign v1445415 = hmaster1_p & v1445414 | !hmaster1_p & v14462ff;
assign a653bc = hmaster2_p & a653bb | !hmaster2_p & a653b8;
assign v14463d2 = hlock2 & v14463d1 | !hlock2 & v14463cc;
assign f2f2ab = hmaster2_p & f2f2a8 | !hmaster2_p & f2f2aa;
assign v1216250 = hbusreq2_p & v121624d | !hbusreq2_p & v121624f;
assign d308b7 = hgrant2_p & d30881 | !hgrant2_p & d308b6;
assign v12161dc = hgrant5_p & v12161d9 | !hgrant5_p & !v12161db;
assign v1214c35 = hbusreq0 & v1214c34 | !hbusreq0 & v845542;
assign v12ad59a = hbusreq1_p & v12ad598 | !hbusreq1_p & v12ad599;
assign v14463aa = hlock0 & v14463a9 | !hlock0 & v14463a7;
assign v121607f = hmaster2_p & v121601d | !hmaster2_p & v845542;
assign d2feeb = hlock2_p & d2feea | !hlock2_p & d2fee7;
assign d306c8 = locked_p & v845542 | !locked_p & !v845580;
assign v138a3ec = hbusreq0 & v138a3e8 | !hbusreq0 & v138a3eb;
assign v1445bd6 = hmaster1_p & v1445bd1 | !hmaster1_p & v1445bd5;
assign v138a068 = hbusreq5_p & v138a067 | !hbusreq5_p & !v845542;
assign v16a13ce = hmaster1_p & v16a2669 | !hmaster1_p & v16a1f96;
assign v138a438 = hmaster1_p & v138a437 | !hmaster1_p & v138a314;
assign f2f33a = hbusreq2_p & f2f338 | !hbusreq2_p & f2f339;
assign v134d440 = hlock0 & v134d43f | !hlock0 & v134d43e;
assign v1445ee0 = hmaster0_p & v1446404 | !hmaster0_p & v1445edf;
assign d30670 = hgrant2_p & v84555e | !hgrant2_p & d3066e;
assign v1216a8d = hready & v1216a8c | !hready & v845542;
assign v138a35f = hmaster0_p & v138a34b | !hmaster0_p & v138a34f;
assign v16a1a23 = hbusreq3 & v16a19e3 | !hbusreq3 & v16a1a22;
assign v1215300 = hbusreq2_p & v12152fd | !hbusreq2_p & v12152ff;
assign v16a16af = hbusreq2 & v16a16ac | !hbusreq2 & !v16a16ae;
assign c50efe = hgrant3_p & c50efd | !hgrant3_p & c50efb;
assign v134d4da = hmaster2_p & v134d4d4 | !hmaster2_p & v134d4d9;
assign v15167b9 = hbusreq2_p & v15167b8 | !hbusreq2_p & v845542;
assign v144615c = hlock5 & v1446140 | !hlock5 & v144615b;
assign v12ad015 = hbusreq5_p & v12ad5dd | !hbusreq5_p & v12ad014;
assign v1215c24 = hbusreq1 & v1216021 | !hbusreq1 & v845542;
assign v15534ed = hmaster2_p & v845542 | !hmaster2_p & v15534ec;
assign v1668dc0 = hbusreq0 & v1668dbc | !hbusreq0 & v1668dbf;
assign v151697f = hmaster1_p & v151697e | !hmaster1_p & v845542;
assign v16a1d1b = hmaster1_p & v16a1d1a | !hmaster1_p & v16a2672;
assign d2fd25 = hmaster1_p & d2fd24 | !hmaster1_p & d30283;
assign v121505d = hmaster1_p & v121505c | !hmaster1_p & v1215054;
assign v1389fc3 = hgrant2_p & v1389fc0 | !hgrant2_p & v1389fbb;
assign v1214bff = hmaster1_p & v1214bfe | !hmaster1_p & v12153a9;
assign v151579d = hgrant5_p & v845570 | !hgrant5_p & v151579c;
assign v15533ab = hlock0_p & v1553217 | !hlock0_p & v15533aa;
assign v1552d7f = hmaster2_p & v845542 | !hmaster2_p & v1552d7e;
assign v1445813 = hlock2 & v144580d | !hlock2 & v1445812;
assign bf1f98 = hbusreq5_p & bf1f64 | !hbusreq5_p & bf1f97;
assign v1446045 = hbusreq1 & v144640c | !hbusreq1 & v1446438;
assign f2f369 = hgrant1_p & v845570 | !hgrant1_p & !f2f368;
assign v1284cba = hmaster0_p & v1284cb9 | !hmaster0_p & v140587e;
assign v151561b = hmastlock_p & v151561a | !hmastlock_p & v845542;
assign v11e597c = hbusreq5_p & v11e5948 | !hbusreq5_p & v11e597b;
assign v1515795 = hgrant1_p & f2f281 | !hgrant1_p & v1515794;
assign v16695ae = hbusreq2_p & v16695ad | !hbusreq2_p & v845542;
assign v10d40b8 = hmaster0_p & v10d3ffd | !hmaster0_p & v10d4052;
assign v15534f2 = hgrant2_p & v15534f1 | !hgrant2_p & v15534dc;
assign v1446559 = hmaster2_p & v845542 | !hmaster2_p & v1446558;
assign v1215387 = hbusreq0 & v1215386 | !hbusreq0 & v845542;
assign v12150ca = hlock5_p & v12150c8 | !hlock5_p & v12150c9;
assign v1445e47 = hgrant1_p & v845542 | !hgrant1_p & v1445e46;
assign v1445e11 = hmaster2_p & v1445de5 | !hmaster2_p & v1445e10;
assign d2fed2 = hlock2_p & d2fed1 | !hlock2_p & d2feca;
assign v134d3ae = hmaster0_p & v845542 | !hmaster0_p & v134d3ad;
assign v14454f9 = hgrant2_p & v1445bec | !hgrant2_p & v14454f8;
assign v1445fad = hlock2 & v1445fa5 | !hlock2 & v1445fac;
assign v134d517 = hmaster2_p & v845542 | !hmaster2_p & v134d36d;
assign d3075f = hlock2_p & d3075d | !hlock2_p & d3075e;
assign v15156c9 = hmaster0_p & v15156c8 | !hmaster0_p & v1515675;
assign v114a3bf = hgrant3_p & v114a22f | !hgrant3_p & v114a3be;
assign v14459d2 = hlock1 & v144660b | !hlock1 & v14459ac;
assign v1445a1e = hmaster2_p & v1445a1d | !hmaster2_p & v144660f;
assign v12af58f = hmaster2_p & v12afe46 | !hmaster2_p & v12af58e;
assign f2f4b3 = hbusreq1_p & f2f4b2 | !hbusreq1_p & !v845542;
assign d2fb47 = hbusreq5 & d2fb40 | !hbusreq5 & d2fb46;
assign v1216a83 = hbusreq5 & v1216a82 | !hbusreq5 & v845542;
assign f2f3cd = hbusreq5_p & f2f3cb | !hbusreq5_p & !f2f3cc;
assign v1515ae4 = hbusreq4 & v15168f4 | !hbusreq4 & !v1668c1c;
assign v14465c4 = hbusreq4 & v14465bb | !hbusreq4 & v14465c3;
assign v114a3be = hready_p & v114a233 | !hready_p & !v845568;
assign v12160a1 = hmaster0_p & v121605f | !hmaster0_p & v121604c;
assign v92fc87 = hburst1_p & v845542 | !hburst1_p & v960a34;
assign v1668da4 = hgrant2_p & v1668d94 | !hgrant2_p & v1668da3;
assign v1215787 = hlock2_p & v1215784 | !hlock2_p & v1215786;
assign v1668dbc = hbusreq5_p & v1668dba | !hbusreq5_p & !v1668dbb;
assign v1516981 = hbusreq2_p & v1516980 | !hbusreq2_p & v845542;
assign v1405ac9 = hmaster1_p & v1405abe | !hmaster1_p & !v1405ac8;
assign v134d245 = hlock2_p & v134d243 | !hlock2_p & v134d244;
assign v16695c8 = jx2_p & v16695c7 | !jx2_p & v1668e0e;
assign v16a1e5f = hbusreq5_p & v845542 | !hbusreq5_p & v16a1e5e;
assign v144642a = hmaster2_p & v1446427 | !hmaster2_p & v1446429;
assign v134cecf = hready_p & v134d34f | !hready_p & v134cece;
assign v1668e07 = hbusreq3 & v1668e06 | !hbusreq3 & a7c7c1;
assign v1215356 = hbusreq0 & v1215355 | !hbusreq0 & v845542;
assign d300e3 = hlock5_p & d300e1 | !hlock5_p & d300e2;
assign v1214d07 = hmaster2_p & v1214c29 | !hmaster2_p & !v1214cf1;
assign v12af9b1 = hbusreq5_p & v12afda4 | !hbusreq5_p & v12af986;
assign v1515aef = decide_p & v1515aee | !decide_p & v845576;
assign v1552fd3 = decide_p & v155342e | !decide_p & v1552fd2;
assign v121627e = decide_p & v12160ce | !decide_p & v121627d;
assign v151577c = hbusreq0_p & v151563e | !hbusreq0_p & a65396;
assign d2f986 = hbusreq3 & d2f97f | !hbusreq3 & !d2f985;
assign v16a20a5 = hbusreq5 & v16a20a4 | !hbusreq5 & v16a209f;
assign v1446202 = hbusreq5 & v14461df | !hbusreq5 & v1446201;
assign v1445546 = hgrant2_p & v1445be3 | !hgrant2_p & v1445545;
assign v1215753 = hbusreq5_p & v121574f | !hbusreq5_p & v1215752;
assign v1216563 = hlock5_p & v121655b | !hlock5_p & v1216562;
assign a654c9 = decide_p & a654c6 | !decide_p & v845542;
assign v1446142 = hmaster1_p & v144611a | !hmaster1_p & v1445ffc;
assign v12166d8 = hgrant4_p & v12166d6 | !hgrant4_p & v12166d7;
assign v15167fa = hmaster1_p & v15167f9 | !hmaster1_p & v1668c23;
assign v1668d42 = hmaster0_p & v1668d34 | !hmaster0_p & v1668d41;
assign v14466bc = hlock2 & v1446676 | !hlock2 & v14466ba;
assign f2f452 = hbusreq5_p & f2f3cb | !hbusreq5_p & !f2f451;
assign v1405acd = hbusreq2_p & v1405ac9 | !hbusreq2_p & v1405acc;
assign v1553053 = hgrant5_p & v1553386 | !hgrant5_p & v1553052;
assign v134d4cb = hbusreq1_p & v134d1dd | !hbusreq1_p & v134d4ca;
assign d3015d = hbusreq2_p & d30150 | !hbusreq2_p & !d3015c;
assign v16a1446 = hbusreq5 & v16a143f | !hbusreq5 & v16a1445;
assign v1445758 = hmaster1_p & v1445da9 | !hmaster1_p & v1445dd1;
assign v1445f03 = hlock5 & v1445ee7 | !hlock5 & v1445f02;
assign d30159 = hbusreq0 & d30154 | !hbusreq0 & d30158;
assign v10d3ffe = hmaster0_p & v10d3ff0 | !hmaster0_p & v10d3ffd;
assign v1214819 = hready_p & v12147ea | !hready_p & v1214818;
assign v134d223 = hmaster1_p & v134d222 | !hmaster1_p & v134d20f;
assign v15156ed = hbusreq2_p & v15156ec | !hbusreq2_p & v845542;
assign v1445b30 = hready_p & v1445bac | !hready_p & v1445b2f;
assign v1446064 = hgrant1_p & v1445fd8 | !hgrant1_p & v1446063;
assign v15533b3 = hbusreq5_p & v15533b2 | !hbusreq5_p & v15533a7;
assign v121507f = hgrant2_p & v1215059 | !hgrant2_p & v121507e;
assign v12ad590 = hbusreq2 & v12ad58a | !hbusreq2 & v12ad58f;
assign v1446431 = hlock1 & v1446423 | !hlock1 & v1446430;
assign v1405926 = locked_p & v1405925 | !locked_p & !v140583c;
assign v1445b80 = hmaster1_p & v1446323 | !hmaster1_p & v1445b7a;
assign v1215c63 = hlock5_p & v1215c61 | !hlock5_p & v1215c62;
assign v16a1b68 = hmaster1_p & v16a1afd | !hmaster1_p & !v16a1f96;
assign v14463e2 = hbusreq4_p & v144639c | !hbusreq4_p & v14463e1;
assign v134d4bc = hgrant3_p & v134d3fc | !hgrant3_p & v134d4bb;
assign a658b5 = hmastlock_p & a658b4 | !hmastlock_p & v845580;
assign v134d53a = hbusreq5 & v134d538 | !hbusreq5 & v134d539;
assign v1216151 = hlock0_p & v1215fec | !hlock0_p & !v845542;
assign v12160b2 = hbusreq2_p & v12160b1 | !hbusreq2_p & v12160b0;
assign v144548a = hlock3 & v1445471 | !hlock3 & v1445489;
assign hgrant0 = !v12acd07;
assign d307d9 = hlock1_p & d307d8 | !hlock1_p & d3065c;
assign a6628f = hmaster2_p & a6628b | !hmaster2_p & a66286;
assign v134d4c3 = hready_p & v134d3be | !hready_p & v134d4c2;
assign v138a3f3 = hmaster0_p & v845542 | !hmaster0_p & v138a31a;
assign v1216715 = hgrant4_p & v845547 | !hgrant4_p & v1216714;
assign v1445364 = hmaster0_p & v1445909 | !hmaster0_p & v1445a38;
assign d3011b = hgrant5_p & d2fea4 | !hgrant5_p & !d30119;
assign v1446166 = hmaster0_p & v1445fe3 | !hmaster0_p & v1446079;
assign v11e5956 = hlock0_p & v11e593a | !hlock0_p & v845570;
assign v1216169 = hgrant1_p & v845542 | !hgrant1_p & v1216168;
assign v1445929 = decide_p & v14458d1 | !decide_p & v1445928;
assign v1284d68 = jx1_p & v140582a | !jx1_p & !v1284d67;
assign v10d42dc = hbusreq2_p & v10d42d9 | !hbusreq2_p & v10d42db;
assign v12150af = hbusreq2 & v1215089 | !hbusreq2 & v12150ae;
assign d2fd4c = hbusreq3_p & d2fd38 | !hbusreq3_p & d2fd4b;
assign d301c3 = hmaster2_p & v845580 | !hmaster2_p & !v845542;
assign d2fb21 = hbusreq5_p & d3013c | !hbusreq5_p & d2fb20;
assign v134d4e2 = hgrant2_p & v134d4e1 | !hgrant2_p & v134d4dd;
assign v1215449 = hmaster1_p & v1215448 | !hmaster1_p & v12153ec;
assign v1405b51 = hbusreq5_p & v1405af7 | !hbusreq5_p & v1405b50;
assign v10d42cd = hmaster1_p & v10d42cc | !hmaster1_p & !v10d404f;
assign v16a12c3 = hmaster1_p & v16a129d | !hmaster1_p & v16a1f96;
assign v14458e4 = hbusreq1 & v14458e0 | !hbusreq1 & v14458e3;
assign v134ce78 = hlock5 & v134d276 | !hlock5 & v134ce77;
assign v134cd84 = hbusreq2_p & v134cd82 | !hbusreq2_p & v134cd83;
assign v1553507 = hbusreq3 & v1553505 | !hbusreq3 & v1553506;
assign d30871 = hbusreq2_p & d3076a | !hbusreq2_p & d30870;
assign v12153f7 = hbusreq2_p & v12153f6 | !hbusreq2_p & v12153f0;
assign v1446261 = hmaster2_p & v1446403 | !hmaster2_p & v14465b9;
assign v1446328 = hmaster1_p & v14462e8 | !hmaster1_p & v1446271;
assign v121614d = hbusreq1 & v121614c | !hbusreq1 & v845542;
assign v14460ce = hlock0 & v14460cd | !hlock0 & v14460cc;
assign d2feff = hlock2_p & d2fefe | !hlock2_p & d2fefa;
assign v121533a = hgrant2_p & v1215329 | !hgrant2_p & v1215339;
assign v1446652 = hlock1 & v144639c | !hlock1 & v14465c1;
assign v16a13fe = hmaster0_p & v16a1d6d | !hmaster0_p & v16a1d6c;
assign v16a1b6a = hbusreq3 & v16a1b66 | !hbusreq3 & v16a1b69;
assign v1215bdd = hbusreq1_p & v1216a5a | !hbusreq1_p & v1215ff8;
assign v1552d9f = hready_p & v1552d9e | !hready_p & v1552d76;
assign v12153a2 = hbusreq0 & v12153a1 | !hbusreq0 & v845542;
assign v12165ad = hgrant5_p & v845542 | !hgrant5_p & v12165ac;
assign d2fb96 = hbusreq2_p & d2fb95 | !hbusreq2_p & d2fb90;
assign v1216230 = hbusreq1 & v12166e5 | !hbusreq1 & !v845542;
assign v11e5974 = hlock0_p & v11e593a | !hlock0_p & v11e5973;
assign v16a1946 = hgrant4_p & v845559 | !hgrant4_p & !v16a1945;
assign v1515619 = hburst1 & v1515618 | !hburst1 & v845542;
assign v1216a6f = hlock5_p & v1216a6e | !hlock5_p & v845542;
assign v16a2093 = hbusreq5_p & v16a2092 | !hbusreq5_p & v16a208b;
assign d80761 = hmaster2_p & d80760 | !hmaster2_p & d80733;
assign v1445aec = hbusreq2_p & v1445ae6 | !hbusreq2_p & v1445aeb;
assign v16a13e9 = hbusreq2_p & v16a13e8 | !hbusreq2_p & v16a1d54;
assign v1405939 = hmaster1_p & v14058df | !hmaster1_p & v14058d8;
assign v15169a0 = hready_p & v845542 | !hready_p & v151699f;
assign v12ad552 = hbusreq2_p & v12ad550 | !hbusreq2_p & v12ad551;
assign d30866 = hbusreq5_p & d30720 | !hbusreq5_p & d30654;
assign v16a142e = hbusreq2_p & v16a13fa | !hbusreq2_p & v16a1aea;
assign v1445b37 = hmaster1_p & v1445b36 | !hmaster1_p & v14458fd;
assign f2f286 = hgrant1_p & f2f285 | !hgrant1_p & !v845542;
assign v1389394 = decide_p & v1389393 | !decide_p & v138a406;
assign v1445f53 = hbusreq2_p & v144674a | !hbusreq2_p & v1445f52;
assign v14461c4 = hgrant2_p & v14461c2 | !hgrant2_p & v14461c3;
assign v12af9d7 = hmaster0_p & v12af9c3 | !hmaster0_p & v12af9d6;
assign v1445be2 = hready_p & v144639b | !hready_p & v1445be1;
assign v1445f65 = hgrant2_p & v1446726 | !hgrant2_p & v1445f64;
assign v1215c8c = hgrant1_p & f2f285 | !hgrant1_p & v1216107;
assign v121622e = hgrant2_p & v1216229 | !hgrant2_p & v121622d;
assign f2e4fb = hmaster0_p & f2f229 | !hmaster0_p & f2f539;
assign v1445372 = hgrant2_p & v1445371 | !hgrant2_p & v144536c;
assign v1445bdd = decide_p & v1445bb4 | !decide_p & v1445bdc;
assign bf1f70 = hmaster1_p & bf1f5e | !hmaster1_p & bf1f6f;
assign v1668d51 = hbusreq1 & a65862 | !hbusreq1 & v845570;
assign d2f970 = hbusreq5_p & d30111 | !hbusreq5_p & d2f96f;
assign v12ad513 = hmastlock_p & v12ad512 | !hmastlock_p & !v138a32a;
assign v138a30b = hmaster1_p & v138a30a | !hmaster1_p & v1668c23;
assign v14459aa = hbusreq4 & v14459a8 | !hbusreq4 & v14459a9;
assign v1389168 = decide_p & v13895a4 | !decide_p & v138a406;
assign v14058b1 = hmaster0_p & v14058a5 | !hmaster0_p & v14058b0;
assign v1284cb3 = hmaster1_p & v1284ca9 | !hmaster1_p & v1284ca7;
assign v1214c57 = hmaster2_p & v1215347 | !hmaster2_p & v121534f;
assign a65913 = hmaster2_p & a658cb | !hmaster2_p & !a658ce;
assign v16a1941 = hgrant1_p & v84554d | !hgrant1_p & v16a1940;
assign v1389fcb = hbusreq5 & v1389f87 | !hbusreq5 & v1389fca;
assign d2fed1 = hmaster1_p & d2fed0 | !hmaster1_p & d2fec6;
assign v12af9b9 = hready_p & v12af7e2 | !hready_p & v12af9b8;
assign v134d268 = hbusreq2_p & v134d267 | !hbusreq2_p & v134d244;
assign v1215361 = hmaster0_p & v1215360 | !hmaster0_p & v845542;
assign v12ad22d = hbusreq2 & v12ad22c | !hbusreq2 & v12afa0f;
assign d300c0 = hbusreq1_p & d300bf | !hbusreq1_p & v84555a;
assign d2fc43 = hbusreq2_p & d2fbbc | !hbusreq2_p & d2fc42;
assign v16a139b = decide_p & v16a1398 | !decide_p & v16a137f;
assign v1445e6b = hbusreq1_p & v14465b2 | !hbusreq1_p & v1445e6a;
assign v1215d00 = hbusreq5_p & v1215cff | !hbusreq5_p & v1215c87;
assign d2fbb9 = hbusreq2 & d2fbb4 | !hbusreq2 & d2fbb8;
assign v12ad5a5 = hlock0_p & v12ad5a3 | !hlock0_p & !v12ad5a4;
assign v144631e = hmaster1_p & v144631d | !hmaster1_p & v144627e;
assign v121572e = hgrant5_p & v1215b9a | !hgrant5_p & !v121572c;
assign v15167ec = hlock2_p & v9745f6 | !hlock2_p & v845542;
assign d3086b = hbusreq1_p & d30728 | !hbusreq1_p & d3068f;
assign d30647 = hgrant4_p & a66284 | !hgrant4_p & d30646;
assign v134ce5d = hbusreq3 & v134ce5b | !hbusreq3 & v134ce5c;
assign d3066c = hbusreq0 & d30664 | !hbusreq0 & d3066b;
assign d30134 = hgrant5_p & v84555a | !hgrant5_p & d300ce;
assign d2fcfe = hmaster0_p & d2fcfd | !hmaster0_p & !d2fcb4;
assign v15157bb = hbusreq4_p & v15157ba | !hbusreq4_p & !v845542;
assign d2fc32 = hmaster2_p & v845542 | !hmaster2_p & !v84554c;
assign v138a069 = hmaster0_p & v138a068 | !hmaster0_p & !v845542;
assign v16a1aed = hbusreq2_p & v16a209e | !hbusreq2_p & v16a1aec;
assign v1668c31 = hmaster1_p & v1668c30 | !hmaster1_p & v845542;
assign v1445ff8 = hmaster2_p & v1445fe7 | !hmaster2_p & v1446412;
assign v12160dc = hbusreq1_p & v12160db | !hbusreq1_p & v845542;
assign d301f9 = hgrant1_p & d301ea | !hgrant1_p & d301f8;
assign v12150aa = hgrant5_p & v1215471 | !hgrant5_p & v12150a9;
assign d2fd3b = decide_p & d2fd3a | !decide_p & v845570;
assign v1668d8c = hmaster1_p & v1668d42 | !hmaster1_p & v1668d8b;
assign v1553237 = hgrant5_p & v845542 | !hgrant5_p & v1553236;
assign v1668cd9 = hmaster0_p & a658ad | !hmaster0_p & v1668cd8;
assign d30241 = hgrant5_p & v845542 | !hgrant5_p & d301ed;
assign v1405b42 = hmaster0_p & v1405af7 | !hmaster0_p & v1405ad8;
assign v134d1f8 = hbusreq1_p & v134d1f7 | !hbusreq1_p & v845542;
assign v10d405c = hbusreq2_p & v10d4051 | !hbusreq2_p & !v10d405b;
assign v12ad56a = hmaster1_p & v12ad569 | !hmaster1_p & !v12ad525;
assign v12ae83c = hbusreq3_p & v12ae76c | !hbusreq3_p & v12aee5e;
assign v1215c0d = hgrant1_p & v1215c0b | !hgrant1_p & v1215c0c;
assign v1215375 = stateA1_p & v845542 | !stateA1_p & !v1216a88;
assign v1214c20 = hmaster1_p & v1214c1f | !hmaster1_p & v1214bcf;
assign a65af0 = hbusreq5_p & a65ad6 | !hbusreq5_p & a65aee;
assign v15534fb = hbusreq5_p & v1553395 | !hbusreq5_p & v15534fa;
assign v1216101 = hmaster2_p & v12160f8 | !hmaster2_p & v1216100;
assign v121575f = hgrant1_p & v1215757 | !hgrant1_p & v121575e;
assign v14454fe = hgrant2_p & v14454fc | !hgrant2_p & v14454fd;
assign v12ad568 = hbusreq2_p & v12ad526 | !hbusreq2_p & v12ad567;
assign f2f329 = hmaster1_p & f2f328 | !hmaster1_p & f2f2db;
assign v134d541 = hbusreq3_p & v134d52d | !hbusreq3_p & v134d540;
assign v155305b = hgrant1_p & v845542 | !hgrant1_p & v155305a;
assign v1214c13 = hmaster1_p & v12153ab | !hmaster1_p & v1214bcf;
assign v138a3e8 = hbusreq5_p & v138a3e7 | !hbusreq5_p & !v845542;
assign v134d3d5 = hbusreq3 & v134d3d4 | !hbusreq3 & v134d276;
assign v12af21d = hmaster2_p & v12af9c1 | !hmaster2_p & v12af21c;
assign v1215057 = hmaster2_p & v121545f | !hmaster2_p & !v1215033;
assign v138944b = hmaster2_p & d2fce7 | !hmaster2_p & v845542;
assign v15534f8 = hbusreq3 & v15534f6 | !hbusreq3 & v15534f7;
assign v14458ce = hbusreq3 & v14458cc | !hbusreq3 & v14458cd;
assign v1214d7b = hgrant2_p & v1214d37 | !hgrant2_p & v1214d7a;
assign v1446126 = hlock2 & v1446125 | !hlock2 & v144611f;
assign v14463f8 = hmaster1_p & v14463f7 | !hmaster1_p & v14463ef;
assign v10d40d8 = hmaster1_p & v10d4092 | !hmaster1_p & v10d407c;
assign a656cd = hmaster0_p & a656c8 | !hmaster0_p & a656cb;
assign d30882 = hmaster0_p & d30804 | !hmaster0_p & d307a6;
assign v1552f53 = hbusreq4 & v155338a | !hbusreq4 & v1553217;
assign v1553934 = stateG2_p & v845542 | !stateG2_p & v1553933;
assign v1216264 = hmaster1_p & v1216263 | !hmaster1_p & !v121624b;
assign v15156b5 = hbusreq2 & v15156b4 | !hbusreq2 & v15167ed;
assign d2fc3f = hbusreq2 & d2fc3d | !hbusreq2 & d2fc3e;
assign v16a208a = hgrant1_p & v84554d | !hgrant1_p & v16a2089;
assign v1216034 = hbusreq1_p & v1216033 | !hbusreq1_p & v845542;
assign v1216037 = hbusreq1_p & v1216036 | !hbusreq1_p & v845542;
assign d300d4 = hmaster2_p & d2fe7d | !hmaster2_p & d2fe85;
assign v1668d9b = hgrant5_p & v1668d9a | !hgrant5_p & v1668d98;
assign v12ad55b = hbusreq2_p & v12ad559 | !hbusreq2_p & v12ad55a;
assign v16a139a = hready_p & v845555 | !hready_p & !v16a1399;
assign bf1f51 = decide_p & bf1f50 | !decide_p & v845570;
assign v14459c5 = hbusreq0_p & v14459c4 | !hbusreq0_p & v144639e;
assign v138a45c = hmaster0_p & v138a354 | !hmaster0_p & v138a34b;
assign v16a16a4 = hbusreq2 & v16a16a1 | !hbusreq2 & !v16a16a3;
assign v15155ea = hmaster0_p & v845542 | !hmaster0_p & v15155e9;
assign v1216207 = hgrant1_p & v1216204 | !hgrant1_p & v1216206;
assign v1515ae7 = hbusreq4_p & v1515ae6 | !hbusreq4_p & v845542;
assign v15157f8 = hbusreq0 & v15157f4 | !hbusreq0 & v15157f7;
assign v12ad011 = hbusreq1_p & v12ad5da | !hbusreq1_p & v12ad010;
assign f2f3b9 = hgrant5_p & v84554c | !hgrant5_p & f2f34d;
assign v16a1429 = hbusreq5 & v16a1423 | !hbusreq5 & v16a1428;
assign v1446149 = hmaster1_p & v1446128 | !hmaster1_p & v1445ffc;
assign v1515733 = hmaster2_p & v1515723 | !hmaster2_p & v845542;
assign v84557c = hgrant5_p & v845542 | !hgrant5_p & !v845542;
assign v16a1d97 = hbusreq3 & v16a1d95 | !hbusreq3 & v16a205d;
assign v12af5ad = hbusreq0 & v12af590 | !hbusreq0 & v12af5ac;
assign v10d3feb = hmaster2_p & v10d3fd5 | !hmaster2_p & v10d3fe0;
assign f2f3f5 = hmaster0_p & f2f2dd | !hmaster0_p & f2f2e8;
assign d2fee7 = hmaster1_p & d2fec9 | !hmaster1_p & d2fee5;
assign v140583c = hmastlock_p & v140583b | !hmastlock_p & !v845542;
assign v12160d7 = hbusreq1 & v12164cf | !hbusreq1 & v845542;
assign v1553426 = hgrant3_p & v155321c | !hgrant3_p & v1553425;
assign v134d497 = hbusreq0 & v134d388 | !hbusreq0 & v134d38b;
assign d2fb86 = hmaster0_p & d2fb6c | !hmaster0_p & d2fb85;
assign v1216590 = locked_p & v121658f | !locked_p & v845542;
assign v1445ebc = hmaster1_p & v1445ebb | !hmaster1_p & v1445eaa;
assign v1445afd = hlock2 & v1445af9 | !hlock2 & v1445afc;
assign v11e594b = hbusreq1_p & v11e594a | !hbusreq1_p & v845570;
assign v1668d63 = hbusreq4_p & v10d3fd8 | !hbusreq4_p & !a65861;
assign v14460e1 = decide_p & v1445fca | !decide_p & v14460e0;
assign v134ced8 = hbusreq2_p & v134ceb9 | !hbusreq2_p & v134d3cd;
assign v1214efd = hgrant2_p & v845542 | !hgrant2_p & v1214efc;
assign v12acfcf = hmaster1_p & v12acfce | !hmaster1_p & !v12ad525;
assign v121574a = hbusreq5_p & v1215742 | !hbusreq5_p & v1215749;
assign v14463bd = hbusreq5_p & v14463b8 | !hbusreq5_p & v14463bc;
assign v1446346 = hbusreq2_p & v1446343 | !hbusreq2_p & v1446345;
assign v1445429 = hgrant2_p & v1445411 | !hgrant2_p & v1445428;
assign v1214d71 = hbusreq2_p & v1214d6e | !hbusreq2_p & v1214d70;
assign v11e594c = hgrant1_p & v11e594b | !hgrant1_p & !v845542;
assign v140590e = hmaster1_p & v140590d | !hmaster1_p & v140584d;
assign v1515766 = hgrant4_p & v1515765 | !hgrant4_p & v1515612;
assign v16a1cd4 = hbusreq2 & v16a1cce | !hbusreq2 & v16a1cd3;
assign d30606 = hbusreq5_p & d30605 | !hbusreq5_p & d305fe;
assign v1215d06 = hgrant2_p & v845542 | !hgrant2_p & !v1215d05;
assign v1215770 = hmaster0_p & v1215754 | !hmaster0_p & v121576f;
assign d2fd00 = hlock2_p & v845542 | !hlock2_p & !d2fcff;
assign v134d315 = hmaster1_p & v134d280 | !hmaster1_p & v134d314;
assign v134cedd = hbusreq5 & v134d3ce | !hbusreq5 & v134cedc;
assign v15161d6 = hbusreq2 & v15161cf | !hbusreq2 & v15161d5;
assign v1668d81 = hbusreq5_p & v1668d7e | !hbusreq5_p & v1668d80;
assign v144660a = hbusreq0_p & v144639c | !hbusreq0_p & v14465bb;
assign v1216a79 = hlock5_p & v1216a74 | !hlock5_p & v1216a78;
assign v12ad52d = hbusreq0 & v12ad52c | !hbusreq0 & !v845542;
assign v16a1cbd = hmaster1_p & v16a1ca0 | !hmaster1_p & v16a1f96;
assign v14457b1 = hmaster1_p & v144577e | !hmaster1_p & v1445e28;
assign v16a1411 = hbusreq2 & v16a1410 | !hbusreq2 & v16a205c;
assign v12157b0 = hgrant4_p & v845542 | !hgrant4_p & v12157af;
assign v1405b3b = decide_p & v1405ab4 | !decide_p & v1405acd;
assign v1553228 = hgrant1_p & v1553227 | !hgrant1_p & v845542;
assign v1215ba2 = hmaster1_p & v1215b9b | !hmaster1_p & !v1215ba1;
assign v1445bf8 = hgrant3_p & v1445bea | !hgrant3_p & v1445bf7;
assign f2f3e5 = hgrant3_p & f2f342 | !hgrant3_p & f2f3e4;
assign v1215c1e = hlock5_p & v1215c1c | !hlock5_p & v1215c1d;
assign v1214f61 = hbusreq2 & v1214f60 | !hbusreq2 & v121671a;
assign v1215dac = hbusreq3 & v1215da9 | !hbusreq3 & v121678b;
assign v1216a7f = hmaster2_p & v845542 | !hmaster2_p & v845547;
assign v14459cf = hgrant1_p & v14459b9 | !hgrant1_p & v14459ce;
assign v1445fe8 = hmaster2_p & v144639c | !hmaster2_p & v1445fe7;
assign v16a1420 = hbusreq2 & v16a141f | !hbusreq2 & v16a1da7;
assign v1215108 = hbusreq2_p & v12150fc | !hbusreq2_p & v12150fb;
assign v1284c92 = hmaster1_p & v1284c91 | !hmaster1_p & v140584d;
assign v1215c7c = hmaster2_p & v845570 | !hmaster2_p & v1215fec;
assign v1445e2b = hbusreq2_p & v1445e29 | !hbusreq2_p & v1445e2a;
assign v14459f8 = hgrant4_p & v14458db | !hgrant4_p & v14459f7;
assign v16a13d0 = hbusreq2_p & v16a13cf | !hbusreq2_p & v16a1f97;
assign v1405a99 = hbusreq2_p & v1405a95 | !hbusreq2_p & v1405a98;
assign v12ad1fe = decide_p & v12ad1fd | !decide_p & v845542;
assign v144537b = hgrant2_p & v1445379 | !hgrant2_p & v144537a;
assign f2f42d = hbusreq5_p & f2f371 | !hbusreq5_p & !f2f42c;
assign v1445433 = hlock5 & v1445427 | !hlock5 & v1445432;
assign v1215c03 = hgrant5_p & v1215be4 | !hgrant5_p & !v1215c01;
assign v1516216 = decide_p & v15167ee | !decide_p & v845542;
assign v1445ec9 = hmaster2_p & v144639c | !hmaster2_p & v1445ec8;
assign v12160e9 = hmaster1_p & v12160e8 | !hmaster1_p & v121600c;
assign v1668c1b = hmastlock_p & v1553933 | !hmastlock_p & !v845542;
assign v1216579 = hbusreq2_p & v1216577 | !hbusreq2_p & v1216578;
assign v15157c2 = hmaster2_p & v15157bd | !hmaster2_p & v15157c1;
assign v1445eb6 = hmaster2_p & v144639c | !hmaster2_p & v1445dec;
assign v138a3d7 = hbusreq5_p & v138a3d6 | !hbusreq5_p & !v845542;
assign v14460e8 = hmaster1_p & v14460e7 | !hmaster1_p & v1445f9e;
assign f2f459 = hgrant2_p & f2f3b4 | !hgrant2_p & !f2f455;
assign v16a1cb9 = hbusreq2 & v16a1ca6 | !hbusreq2 & v16a1ca8;
assign v1405adb = hbusreq1_p & v1405ada | !hbusreq1_p & d3070c;
assign v12aeb74 = hlock0_p & f2f4b0 | !hlock0_p & v845542;
assign v1389f84 = hlock5_p & v1389f83 | !hlock5_p & !v845542;
assign v1515754 = hgrant0_p & a6537d | !hgrant0_p & v151560d;
assign v1446213 = hgrant5_p & v144639c | !hgrant5_p & !v1446212;
assign v16a1d4c = hmaster1_p & v16a1d44 | !hmaster1_p & v16a1d4b;
assign v1215058 = hmaster0_p & v1215463 | !hmaster0_p & v1215057;
assign v121625a = hbusreq1 & v12166c4 | !hbusreq1 & v1216715;
assign v1553441 = hmaster1_p & v1553440 | !hmaster1_p & v1553238;
assign d2fb4f = hmaster2_p & d2fb4d | !hmaster2_p & d2fb4e;
assign v134d30e = hgrant1_p & v845542 | !hgrant1_p & v134d30d;
assign d2f97b = hmaster2_p & v845542 | !hmaster2_p & !d2f97a;
assign v155341c = hmaster0_p & v1553395 | !hmaster0_p & v15533a7;
assign d30767 = hmaster0_p & d3072e | !hmaster0_p & d3071e;
assign v1284cd2 = hmaster2_p & v1405844 | !hmaster2_p & !v1284ccd;
assign d30755 = hmaster1_p & d3071e | !hmaster1_p & d30754;
assign v1389499 = hready_p & v1389466 | !hready_p & v1389498;
assign v12acff6 = hmaster0_p & v12ad634 | !hmaster0_p & v12ad633;
assign v15156ca = hmaster1_p & v15156c9 | !hmaster1_p & !v15156b1;
assign d2fc5a = hbusreq0 & d2fc59 | !hbusreq0 & d306bc;
assign v1445a2d = hgrant1_p & v14458f8 | !hgrant1_p & v1445a2c;
assign v144612e = hmaster1_p & v144612d | !hmaster1_p & v1445fde;
assign d30296 = hgrant2_p & v845542 | !hgrant2_p & !d30294;
assign a6548c = hmaster0_p & a658e8 | !hmaster0_p & a6548b;
assign v1553397 = hbusreq0 & v1553396 | !hbusreq0 & v1553395;
assign d3064f = hlock1_p & d3064e | !hlock1_p & !v845542;
assign d30633 = hmaster0_p & d3060c | !hmaster0_p & d305ed;
assign v16a138a = hmaster0_p & v16a1a97 | !hmaster0_p & v16a1383;
assign d8077c = hgrant1_p & v845542 | !hgrant1_p & !d8077b;
assign d302da = hmaster1_p & d3069a | !hmaster1_p & d302d9;
assign d2fedb = hbusreq2_p & d2feda | !hbusreq2_p & d2fed9;
assign a65af6 = hready_p & a65af5 | !hready_p & a65add;
assign v138a33a = hbusreq5_p & v138a339 | !hbusreq5_p & !v845542;
assign v121509f = hgrant0_p & v121504c | !hgrant0_p & v845559;
assign f2f223 = hmaster1_p & v845542 | !hmaster1_p & f2f222;
assign a6535d = hmaster1_p & a6535b | !hmaster1_p & a6586e;
assign v144552e = hbusreq2 & v144552d | !hbusreq2 & v144551a;
assign d30652 = hmaster2_p & v845542 | !hmaster2_p & d30651;
assign v16a1a84 = hbusreq5_p & v16a1960 | !hbusreq5_p & v16a1a83;
assign v15532cb = hmaster0_p & v15532c3 | !hmaster0_p & v15532ca;
assign v1389f97 = hgrant2_p & v1389f94 | !hgrant2_p & v1389f8f;
assign v12162e9 = hmaster2_p & v1216048 | !hmaster2_p & v1216aad;
assign v1405b4e = hgrant1_p & v1405a86 | !hgrant1_p & v1405b4d;
assign v1445ec0 = hbusreq1 & v1445e57 | !hbusreq1 & v1445ebf;
assign v1214eb5 = hmaster0_p & v12162f6 | !hmaster0_p & v12162e8;
assign v1445bc7 = hmaster1_p & v1445bc6 | !hmaster1_p & v845542;
assign v1445891 = hbusreq4_p & v144639c | !hbusreq4_p & v144586f;
assign f2f3ff = hmaster1_p & f2f3fe | !hmaster1_p & f2f2db;
assign v12160a9 = hmaster1_p & v12160a8 | !hmaster1_p & v121605d;
assign v14466f7 = hbusreq2_p & v14466f1 | !hbusreq2_p & v14466f6;
assign v138a3c7 = hbusreq5_p & v138a3c6 | !hbusreq5_p & !v845542;
assign v1405aea = hlock0_p & v1405a88 | !hlock0_p & !v1405ae9;
assign v144625f = hlock5 & v1446224 | !hlock5 & v144625d;
assign d30812 = hgrant2_p & v84554e | !hgrant2_p & d30806;
assign v1389370 = hmaster0_p & v138936f | !hmaster0_p & v845542;
assign v1445ad7 = hmaster1_p & v1445ac2 | !hmaster1_p & v14458c1;
assign v1552d88 = hlock0_p & v1553138 | !hlock0_p & v1552d87;
assign a653b9 = hmaster2_p & a65389 | !hmaster2_p & a653b8;
assign v12166fc = hmaster2_p & v12164cf | !hmaster2_p & !v12166e5;
assign v155308a = hmaster2_p & v845542 | !hmaster2_p & v1553089;
assign v134d4fa = hgrant4_p & v134d4f9 | !hgrant4_p & v845542;
assign v144661a = hlock0_p & v144639c | !hlock0_p & v1446619;
assign v1284cce = hmaster2_p & v14463b1 | !hmaster2_p & !v1284ccd;
assign v11e596b = hmaster0_p & v11e5963 | !hmaster0_p & !v11e596a;
assign a65424 = hmaster2_p & a65399 | !hmaster2_p & v845558;
assign v1445a87 = hgrant2_p & v1445a85 | !hgrant2_p & v1445a86;
assign v1214c7f = hbusreq2_p & v1214c76 | !hbusreq2_p & v1214c7e;
assign v134ce5a = hlock2 & v134d3b5 | !hlock2 & v134ce48;
assign v1668dc5 = hgrant5_p & v1668dc4 | !hgrant5_p & !v1668d55;
assign v1553417 = hmaster0_p & v845542 | !hmaster0_p & v1553416;
assign v144579d = hlock0 & v144579c | !hlock0 & v144579b;
assign v138a47c = hgrant2_p & v138a479 | !hgrant2_p & !v138a47b;
assign v138a345 = hmaster0_p & v138a32d | !hmaster0_p & v138a344;
assign v16a2062 = hmaster1_p & v9109e4 | !hmaster1_p & v16a1f96;
assign v155339d = hlock1 & v155339c | !hlock1 & v155339b;
assign v134d4fd = hlock1 & v134d4fc | !hlock1 & v134d4fa;
assign v12acfe6 = hbusreq2_p & v12acfe4 | !hbusreq2_p & v12acfe5;
assign a65afe = hmaster0_p & v845542 | !hmaster0_p & !a6627a;
assign v1405896 = hbusreq5_p & v1405895 | !hbusreq5_p & v1405894;
assign v1553514 = hlock5 & v155321a | !hlock5 & v1553513;
assign v144541c = hbusreq2_p & v1445416 | !hbusreq2_p & v144541b;
assign v1389466 = decide_p & v1389465 | !decide_p & v138a406;
assign v12ae1f8 = hlock4_p & v12ae1f5 | !hlock4_p & !v12ae1f7;
assign v15156f1 = hmaster2_p & v151564d | !hmaster2_p & a658d4;
assign v134ce55 = hmaster0_p & v845542 | !hmaster0_p & v134ce54;
assign v144606d = hbusreq1_p & v1446629 | !hbusreq1_p & v144660e;
assign v1214dda = hbusreq2 & v1214dd9 | !hbusreq2 & v845542;
assign v1445eeb = stateG10_5_p & v1445e6d | !stateG10_5_p & v1445eea;
assign v1214e59 = hmaster2_p & v1216048 | !hmaster2_p & v1214e58;
assign v1216ada = hlock0_p & v1216aad | !hlock0_p & v845547;
assign d3078c = hmastlock_p & d3078b | !hmastlock_p & v845542;
assign v144583d = hlock2 & v14457f6 | !hlock2 & v144583c;
assign v144626b = hmaster1_p & v1446405 | !hmaster1_p & v144626a;
assign v1445503 = hgrant5_p & v1446445 | !hgrant5_p & v1445502;
assign v155343b = hgrant4_p & v845542 | !hgrant4_p & v155343a;
assign v16a1a7e = hgrant2_p & v845542 | !hgrant2_p & v16a1a7d;
assign v1405af0 = hmaster0_p & v1405ae4 | !hmaster0_p & !v1405aef;
assign d301c2 = hmaster1_p & d301bb | !hmaster1_p & d301c1;
assign v14058b2 = hmaster1_p & v1405896 | !hmaster1_p & v14058b1;
assign v1215bb6 = hlock2_p & v1215bb5 | !hlock2_p & v12163ab;
assign d2fbe3 = hgrant5_p & v84554a | !hgrant5_p & d2fbe1;
assign v1215d6f = hmaster2_p & v12164d3 | !hmaster2_p & v12164d9;
assign v134d21b = hlock2_p & v134d21a | !hlock2_p & v134d20c;
assign v134d1ff = hmaster2_p & v134d1e8 | !hmaster2_p & v134d1fc;
assign a658ca = hmastlock_p & a658c9 | !hmastlock_p & v845542;
assign v12166f5 = hmaster1_p & v12166f4 | !hmaster1_p & v12164e1;
assign v134cd45 = jx1_p & v134d46d | !jx1_p & v134cd44;
assign v1445f5d = hbusreq2_p & v144674a | !hbusreq2_p & v1445f5c;
assign v1446737 = hmaster1_p & v1446736 | !hmaster1_p & v144644d;
assign d306a6 = hbusreq1_p & v845542 | !hbusreq1_p & d306a5;
assign v11e596c = hmaster1_p & v11e5948 | !hmaster1_p & !v11e596b;
assign v16a1336 = hmaster1_p & v16a132e | !hmaster1_p & !v16a2672;
assign v121679c = hmaster1_p & v121679b | !hmaster1_p & v12164e1;
assign v138a3f4 = hmaster1_p & v138a3f3 | !hmaster1_p & v845542;
assign v10d40cd = hmaster1_p & v10d4083 | !hmaster1_p & !v10d407c;
assign v1215b9f = hbusreq5_p & v1215b9d | !hbusreq5_p & v1215b9e;
assign v138a458 = hmaster1_p & v138a457 | !hmaster1_p & v138a341;
assign f2f361 = hbusreq1 & a65394 | !hbusreq1 & !v845542;
assign v1389447 = hlock5_p & v1389446 | !hlock5_p & v845542;
assign v1446727 = hmaster0_p & v144664a | !hmaster0_p & v14465b8;
assign d3023e = hgrant5_p & v845542 | !hgrant5_p & d301d2;
assign v16a1e62 = hmaster2_p & v16a1e5d | !hmaster2_p & !v845542;
assign v14457a8 = hbusreq2_p & v144579f | !hbusreq2_p & v14457a7;
assign v144648d = hgrant4_p & v144648c | !hgrant4_p & v845542;
assign v14459a3 = hbusreq0 & v144599f | !hbusreq0 & v14459a2;
assign v1445e46 = hgrant4_p & v845542 | !hgrant4_p & v1445e45;
assign v1446728 = hmaster1_p & v1446727 | !hmaster1_p & v1446630;
assign d308ae = hmaster1_p & d30895 | !hmaster1_p & d308ad;
assign f2f395 = hgrant2_p & f2f344 | !hgrant2_p & f2f394;
assign v16693a1 = hmaster0_p & v16693a0 | !hmaster0_p & a6587e;
assign v1446272 = hmaster1_p & v1446405 | !hmaster1_p & v1446271;
assign v16a1a94 = hbusreq0 & v16a1a93 | !hbusreq0 & !v845542;
assign v155338b = hlock4 & v1553217 | !hlock4 & v155338a;
assign v1446077 = hmaster2_p & v144639c | !hmaster2_p & v14465d9;
assign v1552f7b = hbusreq5_p & v1552f5a | !hbusreq5_p & v1552f7a;
assign v1552f58 = hgrant1_p & v1552f57 | !hgrant1_p & v845542;
assign v10d3fdb = locked_p & v845542 | !locked_p & !v10d3fd8;
assign v1445bb8 = hmaster1_p & v1445bb5 | !hmaster1_p & v1445bb7;
assign v1552d7d = hbusreq1_p & v1553138 | !hbusreq1_p & v1552d7c;
assign f2ed8d = decide_p & f2f4c2 | !decide_p & f2f23c;
assign d2fe95 = hmaster0_p & d2fe94 | !hmaster0_p & d2fe80;
assign v16a1ac4 = hmaster0_p & v16a2675 | !hmaster0_p & v16a1abd;
assign d2fcf4 = hbusreq3 & d2fcd9 | !hbusreq3 & d2fcf3;
assign v121600f = hmaster0_p & v1215ff0 | !hmaster0_p & v121600e;
assign v10d4047 = hlock0_p & v10d3fd9 | !hlock0_p & v10d4046;
assign v16a1377 = hgrant2_p & v16a2060 | !hgrant2_p & v16a1376;
assign v121506c = hmaster1_p & v121506b | !hmaster1_p & v1215054;
assign v12af9b5 = hmaster1_p & v12af7f7 | !hmaster1_p & v12af9b4;
assign v1405b05 = hgrant4_p & v1405a92 | !hgrant4_p & !v1405b04;
assign v1214f3d = decide_p & v1214f1b | !decide_p & v1214f3c;
assign v12acfb4 = hbusreq4_p & v12ad521 | !hbusreq4_p & !v12acfb3;
assign v15156e9 = hbusreq2 & v15156e8 | !hbusreq2 & v15167ed;
assign v1445512 = hbusreq3 & v1445510 | !hbusreq3 & v1445511;
assign d30289 = hmaster1_p & d30288 | !hmaster1_p & v845570;
assign v16a207d = hgrant4_p & v845559 | !hgrant4_p & !v16a207c;
assign a6543f = hbusreq5_p & a6543d | !hbusreq5_p & !a6543e;
assign v151583b = hbusreq0 & v1515836 | !hbusreq0 & v151583a;
assign v134d3c2 = hmaster2_p & v134d3c1 | !hmaster2_p & v845542;
assign v1668cd0 = hbusreq4_p & v1668ccf | !hbusreq4_p & !v845542;
assign v12ad526 = hmaster1_p & v12ad517 | !hmaster1_p & !v12ad525;
assign d2fafd = hbusreq5_p & d300f1 | !hbusreq5_p & d2fafc;
assign d2fb8d = hmaster0_p & d2fb8c | !hmaster0_p & d2fb6c;
assign d30659 = hgrant1_p & f2f227 | !hgrant1_p & d30658;
assign v1445ab8 = hmaster0_p & v14458a6 | !hmaster0_p & v14458aa;
assign v144601b = hmaster0_p & v845542 | !hmaster0_p & v144601a;
assign v121504a = hbusreq4 & v12166e5 | !hbusreq4 & !v845542;
assign v134d1fb = hlock1_p & v134d1e8 | !hlock1_p & v845542;
assign v15156fc = hmaster1_p & v15156fb | !hmaster1_p & v151566b;
assign v144602b = hgrant2_p & v144601c | !hgrant2_p & v1446018;
assign v1215011 = hbusreq4_p & v1215010 | !hbusreq4_p & v845542;
assign v16a1da5 = hmaster1_p & v845564 | !hmaster1_p & v16a2672;
assign v15530a1 = hlock3 & v155341e | !hlock3 & v15530a0;
assign v1446607 = hbusreq4_p & v14465b1 | !hbusreq4_p & v14465d6;
assign v121652e = hgrant1_p & v1216522 | !hgrant1_p & v121652d;
assign v155322a = hgrant5_p & v1553225 | !hgrant5_p & v1553229;
assign v1216b03 = hbusreq5_p & v1216b02 | !hbusreq5_p & v845542;
assign v12ad324 = hgrant1_p & d30690 | !hgrant1_p & v12ad323;
assign v12acfee = hbusreq5 & v12acfd6 | !hbusreq5 & v12acfed;
assign v1445f9e = hmaster0_p & v1445f91 | !hmaster0_p & v1445f9d;
assign f2f233 = hbusreq1 & v845570 | !hbusreq1 & v845542;
assign v1216161 = hgrant1_p & v845542 | !hgrant1_p & v1216160;
assign v1284cf6 = hbusreq0_p & v1284c8f | !hbusreq0_p & v1284ce9;
assign v1668c75 = hmaster0_p & v1668c5f | !hmaster0_p & v1668c74;
assign v134d3ce = hbusreq2_p & v134d26f | !hbusreq2_p & v134d3cd;
assign a65474 = hmaster2_p & a6627b | !hmaster2_p & a65473;
assign v1214c2e = hbusreq0 & v1214c2d | !hbusreq0 & v16a2243;
assign v1214cc1 = hbusreq0 & v1214cc0 | !hbusreq0 & v845542;
assign v10d4036 = hgrant5_p & v10d4035 | !hgrant5_p & !v10d4033;
assign v1389ffc = hlock5_p & v1389ffb | !hlock5_p & !v845542;
assign v14453c4 = decide_p & v1445ae4 | !decide_p & v14453c3;
assign v15161fa = hmaster1_p & v15161f9 | !hmaster1_p & v845570;
assign v16a132f = hmaster0_p & v16a1329 | !hmaster0_p & v16a132e;
assign v16a1bf2 = hbusreq0 & v16a207a | !hbusreq0 & v16a1bf1;
assign v1215761 = hgrant5_p & v1215b87 | !hgrant5_p & v1215760;
assign v10d4052 = hmaster2_p & v10d3fd4 | !hmaster2_p & !v10d402b;
assign f2f456 = hgrant2_p & f2f41c | !hgrant2_p & f2f455;
assign v16a1954 = hgrant4_p & v845559 | !hgrant4_p & v16a1953;
assign d3076d = hmaster1_p & d3076c | !hmaster1_p & d3072c;
assign v12160ae = hmaster1_p & v12160ad | !hmaster1_p & v121605d;
assign v144672d = hgrant2_p & v144672b | !hgrant2_p & v144672c;
assign v12161d3 = hgrant5_p & v1216038 | !hgrant5_p & v12161d2;
assign v12166d1 = hbusreq1_p & v12166d0 | !hbusreq1_p & v12166c4;
assign v1284cbc = hmaster2_p & v140587c | !hmaster2_p & !v1446406;
assign f2f410 = hbusreq2_p & f2f40e | !hbusreq2_p & f2f40f;
assign v1405917 = hmaster1_p & v1405916 | !hmaster1_p & v140586f;
assign v1445b77 = hbusreq5_p & v144668e | !hbusreq5_p & v1445b76;
assign a65b2f = decide_p & a65b2e | !decide_p & a662a2;
assign d301e2 = hlock5_p & d301d9 | !hlock5_p & !d301e1;
assign v1446311 = hbusreq0 & v144630b | !hbusreq0 & v1446310;
assign v1445a64 = hmaster0_p & v14458d4 | !hmaster0_p & v1445a36;
assign v1445a46 = hgrant2_p & v1445a3a | !hgrant2_p & v1445a45;
assign v144542f = hlock2 & v144541f | !hlock2 & v144542e;
assign v14460f9 = hbusreq2_p & v14460f6 | !hbusreq2_p & v14460f8;
assign v1446707 = hbusreq2_p & v1446704 | !hbusreq2_p & v1446706;
assign f2f2e7 = hbusreq1_p & f2f2e6 | !hbusreq1_p & !v845542;
assign v1552d57 = hlock2 & v1552d4e | !hlock2 & v1552d56;
assign v1215c2c = hgrant5_p & v1215bea | !hgrant5_p & v1215c2a;
assign v1553516 = decide_p & v155342e | !decide_p & v1553515;
assign d3066f = hgrant2_p & d30643 | !hgrant2_p & d3066e;
assign v144647f = hgrant1_p & v845542 | !hgrant1_p & v144647e;
assign v14461f4 = hbusreq2_p & v14461ee | !hbusreq2_p & v14461f3;
assign v1669592 = hready_p & v845542 | !hready_p & v1669591;
assign v12ad54a = hmaster2_p & a658dc | !hmaster2_p & !v12ad51c;
assign d3077d = hmaster0_p & d306d1 | !hmaster0_p & d306ce;
assign v134ce46 = hmaster0_p & v134ce3b | !hmaster0_p & v134ce45;
assign v1445842 = hlock5 & v144581c | !hlock5 & v1445841;
assign d3077b = decide_p & d3077a | !decide_p & v845570;
assign v15156f6 = hmaster1_p & v15156f5 | !hmaster1_p & !v15156b1;
assign v16a195c = hmaster1_p & v16a194f | !hmaster1_p & v16a195b;
assign v1214dc7 = decide_p & v1214d6c | !decide_p & v1214dc6;
assign v1515aeb = hlock2_p & v1515aea | !hlock2_p & !v845542;
assign v16a2664 = stateG2_p & v845542 | !stateG2_p & !d3094a;
assign v16a1887 = hbusreq2 & v16a1847 | !hbusreq2 & v16a1848;
assign v12adf5f = hlock0_p & v15160fd | !hlock0_p & v845542;
assign v1515833 = hmaster2_p & v1515723 | !hmaster2_p & v1515750;
assign v121603b = hbusreq5_p & v121603a | !hbusreq5_p & f2f2ad;
assign d3072a = hmaster2_p & d30723 | !hmaster2_p & d30729;
assign v1214cce = hmaster2_p & v1214cbc | !hmaster2_p & v1214cca;
assign v121546e = hmaster2_p & v845542 | !hmaster2_p & v121546d;
assign d308c8 = hmaster1_p & d308bc | !hmaster1_p & d308c7;
assign v1216288 = hmaster0_p & v1216029 | !hmaster0_p & v1216172;
assign v16a1acc = hmaster0_p & v16a1ac9 | !hmaster0_p & !v845542;
assign f2ec24 = hmaster0_p & f2ec23 | !hmaster0_p & v845542;
assign d307d1 = hlock0_p & v845542 | !hlock0_p & d307d0;
assign v134d1e0 = hmaster1_p & v134d1df | !hmaster1_p & v845542;
assign v1216a88 = hburst1_p & v1216a86 | !hburst1_p & v1216a87;
assign a65b29 = hgrant2_p & v845542 | !hgrant2_p & a6628c;
assign v12afda9 = hgrant4_p & v12afda8 | !hgrant4_p & v12afda6;
assign v1446398 = locked_p & v1446397 | !locked_p & v845542;
assign v1445816 = hgrant2_p & v1445815 | !hgrant2_p & v1445810;
assign v134d49c = hgrant2_p & v134d364 | !hgrant2_p & v134d49b;
assign v10d42d8 = hmaster1_p & v10d42d7 | !hmaster1_p & v10d407c;
assign v1445ffc = hmaster0_p & v1445ffb | !hmaster0_p & v1445fdd;
assign d30879 = hbusreq2 & d30877 | !hbusreq2 & d30878;
assign v1389fdb = hgrant5_p & d30274 | !hgrant5_p & !v845542;
assign v134d316 = hgrant2_p & v134d27a | !hgrant2_p & v134d315;
assign v1216544 = hbusreq1 & v1216a67 | !hbusreq1 & v1216a77;
assign v1214c27 = hlock3_p & v1214bf8 | !hlock3_p & v1214c26;
assign a65b0d = hgrant2_p & v845542 | !hgrant2_p & a65b0a;
assign d2f9c9 = hlock5_p & d2f9c8 | !hlock5_p & d2f98e;
assign v1445b00 = hlock3 & v1445af4 | !hlock3 & v1445aff;
assign v12161a4 = hgrant2_p & v1216174 | !hgrant2_p & !v12161a3;
assign d2fc39 = hbusreq5_p & v845542 | !hbusreq5_p & d2fc38;
assign v121536f = hbusreq2_p & v121536c | !hbusreq2_p & v121536e;
assign d307e8 = hgrant0_p & d307e7 | !hgrant0_p & v845542;
assign a656b4 = decide_p & a656b2 | !decide_p & a662a2;
assign d3087c = hready_p & d30862 | !hready_p & !d3087b;
assign v1284d1a = hgrant0_p & v1284c8f | !hgrant0_p & !v144660c;
assign v14058d0 = hgrant1_p & v1405849 | !hgrant1_p & v14058cf;
assign v15157fb = hmaster2_p & v1515630 | !hmaster2_p & v845570;
assign v1214bfc = hlock2_p & v1214bfa | !hlock2_p & v1214bfb;
assign d3094b = stateG3_2_p & v845542 | !stateG3_2_p & !d3094a;
assign v1445fe1 = hmaster2_p & v144639c | !hmaster2_p & v1445fcf;
assign v15168f5 = hbusreq1 & v15168f4 | !hbusreq1 & v845542;
assign v1215064 = hmaster2_p & v121502a | !hmaster2_p & v1214ffe;
assign v1446740 = hmaster0_p & v1446440 | !hmaster0_p & v144667f;
assign v1446440 = hlock0 & v144643f | !hlock0 & v144643c;
assign d308dd = hmaster0_p & d308dc | !hmaster0_p & v845542;
assign d3021a = hgrant2_p & d301cc | !hgrant2_p & d30219;
assign v12153fa = hmaster1_p & v12153f9 | !hmaster1_p & v12153ec;
assign v16a1d7f = hbusreq2 & v16a1d7d | !hbusreq2 & !v16a1d7e;
assign d2fefe = hmaster1_p & d2fefd | !hmaster1_p & d2fec6;
assign v12aee5f = hbusreq3_p & v12aecdc | !hbusreq3_p & v12aee5e;
assign v14459e9 = hgrant5_p & v14459e4 | !hgrant5_p & v14459e8;
assign v1553395 = hgrant5_p & v1553386 | !hgrant5_p & v1553394;
assign v10d4021 = hlock0_p & v10d3fdb | !hlock0_p & !v10d3fd8;
assign v1214f0b = hlock5_p & v1214f09 | !hlock5_p & v1214f0a;
assign v16a13db = hbusreq0 & v16a2071 | !hbusreq0 & v16a2082;
assign v16a1cde = hmaster1_p & v16a1cd1 | !hmaster1_p & !v16a1f96;
assign v16693a9 = hmaster1_p & v16693a8 | !hmaster1_p & v845542;
assign v1552d77 = hready_p & v1553444 | !hready_p & v1552d76;
assign v12add47 = hlock4_p & v12add46 | !hlock4_p & v12aeb74;
assign v134d522 = hmaster1_p & v134d521 | !hmaster1_p & v845542;
assign v12ad4e0 = hbusreq0 & v12ad4df | !hbusreq0 & v845542;
assign v12acfd6 = hbusreq3 & v12acfc8 | !hbusreq3 & v12acfd5;
assign v144553f = hmaster1_p & v144639c | !hmaster1_p & v144553e;
assign v12ad033 = hbusreq2_p & v12ad031 | !hbusreq2_p & !v12ad032;
assign v10d42ae = locked_p & v10d3fd4 | !locked_p & v10d427c;
assign d30688 = hbusreq4_p & v845542 | !hbusreq4_p & v845548;
assign d2f9d6 = hbusreq2 & d2f9d2 | !hbusreq2 & d2f9d5;
assign v1445d7f = hbusreq4 & v144639e | !hbusreq4 & v14463d7;
assign v1216553 = hbusreq4_p & v1216552 | !hbusreq4_p & v845547;
assign v12ad5e9 = hgrant5_p & v12ad4df | !hgrant5_p & v12ad5e8;
assign v1215c34 = hbusreq0 & v1215c2d | !hbusreq0 & v1215c33;
assign v1215bf9 = hgrant5_p & v121601c | !hgrant5_p & !v1215bf7;
assign v1445ffd = hmaster1_p & v1446405 | !hmaster1_p & v1445ffc;
assign d30681 = decide_p & d30680 | !decide_p & v845570;
assign v12150cb = hbusreq5_p & v12150ca | !hbusreq5_p & v12150c9;
assign v134ce72 = hmaster0_p & v134ce54 | !hmaster0_p & v845542;
assign v1445772 = hlock5 & v1445756 | !hlock5 & v1445771;
assign f2f3b2 = hmaster2_p & v84554c | !hmaster2_p & f2f3b1;
assign v12ad5f0 = hbusreq2_p & v12ad5e3 | !hbusreq2_p & v12ad5ef;
assign v134d39a = hmaster0_p & v134d37c | !hmaster0_p & v134d399;
assign v1446007 = hlock5 & v1445ff7 | !hlock5 & v1446006;
assign v1405b35 = hmaster0_p & v1405af3 | !hmaster0_p & v1405a8a;
assign v1446456 = hlock2 & v1446455 | !hlock2 & v144644b;
assign v121576f = hbusreq0 & v1215763 | !hbusreq0 & v121576e;
assign f2e278 = hmaster0_p & f2e277 | !hmaster0_p & v845542;
assign a646dc = hready_p & v845542 | !hready_p & a646db;
assign v10d3ff4 = hmaster2_p & v10d3fd8 | !hmaster2_p & v10d3ff3;
assign d30791 = hlock1_p & d30787 | !hlock1_p & d30790;
assign v1445b69 = hmaster1_p & v144631d | !hmaster1_p & v1446290;
assign f2f3d9 = hmaster0_p & f2f3be | !hmaster0_p & f2f3d8;
assign v14461e8 = hlock2 & v14461e4 | !hlock2 & v14461e7;
assign v14454ed = hgrant5_p & v144643d | !hgrant5_p & v14454ec;
assign d2fbbc = hlock2_p & d2fbba | !hlock2_p & d2fbbb;
assign f2e730 = hmaster2_p & f2f22a | !hmaster2_p & f2f228;
assign v16a1406 = hbusreq2_p & v16a1405 | !hbusreq2_p & v16a209d;
assign v144539a = hbusreq2_p & v1445392 | !hbusreq2_p & v1445399;
assign d3065e = hmaster2_p & d30659 | !hmaster2_p & d3065d;
assign v1215fff = hbusreq4_p & v1216a5a | !hbusreq4_p & v845570;
assign v12164d6 = hmaster2_p & v12164cf | !hmaster2_p & v845570;
assign f2f3d2 = hgrant5_p & f2f2a8 | !hgrant5_p & !f2f39f;
assign v1215022 = decide_p & v1214fca | !decide_p & v1215021;
assign v16a1e70 = hbusreq2_p & v16a1f97 | !hbusreq2_p & v16a1e6f;
assign v1552d49 = hbusreq0 & v15533a4 | !hbusreq0 & v15533a7;
assign v1445513 = hmaster1_p & v14454f0 | !hmaster1_p & v1445b5f;
assign v1405b00 = hgrant5_p & v1405ad9 | !hgrant5_p & v1405aff;
assign v138a034 = hgrant2_p & v845542 | !hgrant2_p & !v138a033;
assign v138a331 = hlock1_p & v138a330 | !hlock1_p & v1515656;
assign v1216b16 = hbusreq2 & v1216b12 | !hbusreq2 & v1216b15;
assign v14463b6 = hlock1 & v14463b5 | !hlock1 & v14463b3;
assign v1214df6 = hlock5_p & v1214df4 | !hlock5_p & v1214df5;
assign v12ad5b0 = hgrant1_p & v12ad5aa | !hgrant1_p & v12ad5af;
assign v1516957 = decide_p & v15168b6 | !decide_p & !v845576;
assign v1445f6b = hgrant2_p & v1446741 | !hgrant2_p & v1445f6a;
assign v1445a4d = hmaster2_p & v14458d2 | !hmaster2_p & v1445a4c;
assign v144613e = hbusreq2 & v144613c | !hbusreq2 & v144613d;
assign v1216096 = hbusreq5_p & v1216095 | !hbusreq5_p & v1216094;
assign v1215043 = hlock0_p & v1215460 | !hlock0_p & v1215042;
assign v1214bc0 = hmaster1_p & v1214bbf | !hmaster1_p & v12153a9;
assign v12af1be = hbusreq5_p & v12af3a9 | !hbusreq5_p & v12af1bd;
assign d30760 = hbusreq2_p & d3075f | !hbusreq2_p & d3075e;
assign d8079a = hmaster2_p & d80794 | !hmaster2_p & d80799;
assign v1215c42 = hgrant5_p & v1215c3c | !hgrant5_p & v1215c41;
assign v134d1e1 = hlock3_p & v134d1e0 | !hlock3_p & v845542;
assign d3063b = hbusreq2_p & d3063a | !hbusreq2_p & d30635;
assign v1446420 = hbusreq0_p & v1446403 | !hbusreq0_p & v144640a;
assign v12152ef = hgrant2_p & v12152ed | !hgrant2_p & !v12152ee;
assign v1405a93 = hmaster2_p & v1405a90 | !hmaster2_p & v1405a92;
assign v15532c8 = hgrant1_p & v845542 | !hgrant1_p & v15532c7;
assign v16a12eb = hmaster2_p & v16a12ea | !hmaster2_p & v16a206f;
assign d308d4 = jx2_p & d306c7 | !jx2_p & d308d3;
assign a653ab = hmaster2_p & a65395 | !hmaster2_p & !a653aa;
assign a65364 = stateG3_2_p & v845542 | !stateG3_2_p & a65854;
assign d2feb1 = hlock4_p & v845542 | !hlock4_p & d2feb0;
assign v16a1cbc = hgrant2_p & v16a205f | !hgrant2_p & v16a1cbb;
assign v16a1bb8 = locked_p & v16a1bb7 | !locked_p & !v845542;
assign v1389f8f = hmaster1_p & v845542 | !hmaster1_p & v1389f8e;
assign v1553057 = hbusreq4_p & v1553217 | !hbusreq4_p & v1553056;
assign v144604c = hbusreq5_p & v1446042 | !hbusreq5_p & v144604b;
assign v16a1bec = hbusreq2 & v16a1bea | !hbusreq2 & !v16a1beb;
assign v14465ea = hmaster2_p & v14465e9 | !hmaster2_p & v1446432;
assign v16a16a0 = hgrant2_p & v845542 | !hgrant2_p & v16a169f;
assign v121657d = hmaster1_p & v121657c | !hmaster1_p & v845542;
assign d308cb = hgrant2_p & d30810 | !hgrant2_p & d308b6;
assign d2f98d = hmaster2_p & d2feb4 | !hmaster2_p & d2f98c;
assign v1214c4f = hbusreq1_p & v1214c4d | !hbusreq1_p & v1214c4e;
assign v138a3ed = hmaster0_p & v138a3cb | !hmaster0_p & v138a3ec;
assign f2f4aa = hmaster2_p & v845542 | !hmaster2_p & !f2f4a9;
assign v12147f0 = hbusreq2_p & v12147ef | !hbusreq2_p & v12164e7;
assign v1445f98 = hbusreq1_p & v14463b5 | !hbusreq1_p & v14463bb;
assign v1214c4c = hgrant1_p & v1214c46 | !hgrant1_p & v1214c4b;
assign v144620c = hmaster2_p & v14463a2 | !hmaster2_p & v14463a3;
assign v1445892 = hlock1 & v1445891 | !hlock1 & v1445890;
assign v12160af = hmaster0_p & v121606b | !hmaster0_p & v121605f;
assign v12161cc = hmaster0_p & v1216038 | !hmaster0_p & v1216035;
assign v134d27d = hgrant4_p & v845542 | !hgrant4_p & v134d27c;
assign v16a1436 = hready_p & v845555 | !hready_p & !v16a2065;
assign d80768 = hmaster1_p & d80767 | !hmaster1_p & v845542;
assign a658bb = hburst1 & v156645f | !hburst1 & a658ba;
assign v1216029 = hmaster2_p & v121601c | !hmaster2_p & !v121601f;
assign v10d40d7 = hmaster1_p & v10d40d6 | !hmaster1_p & !v10d3fe9;
assign v12ad004 = hgrant1_p & v12ad5ca | !hgrant1_p & v12ad003;
assign v144590f = hmaster1_p & v14458d5 | !hmaster1_p & v144590e;
assign v1214e42 = hbusreq2_p & v1214e41 | !hbusreq2_p & v845542;
assign v16a1bf9 = hgrant2_p & v845542 | !hgrant2_p & !v16a1bf7;
assign a656ab = hbusreq2_p & a656a5 | !hbusreq2_p & a656a9;
assign a658ff = hbusreq2_p & a658fc | !hbusreq2_p & a658fe;
assign v1215746 = hbusreq1_p & v1215744 | !hbusreq1_p & v1215745;
assign v1552d69 = hlock5 & v1552d5a | !hlock5 & v1552d68;
assign v12ad8e6 = hbusreq5_p & v12adf5e | !hbusreq5_p & v12ad8e5;
assign v1446633 = hlock1 & v144639c | !hlock1 & v14465be;
assign d300e8 = hbusreq1_p & d300e7 | !hbusreq1_p & d300e6;
assign v144619c = hmaster1_p & v1446161 | !hmaster1_p & v1445ffc;
assign v10d4097 = decide_p & v10d4009 | !decide_p & v10d4096;
assign v1215794 = hgrant5_p & v1215791 | !hgrant5_p & v1215748;
assign v144639b = hmaster1_p & v144639a | !hmaster1_p & v845542;
assign v14465b2 = hgrant4_p & v1446403 | !hgrant4_p & v14465b1;
assign v1284d44 = hlock2_p & v1284d43 | !hlock2_p & v140591e;
assign v16a1ccf = hmaster2_p & v16a1cca | !hmaster2_p & !v845542;
assign v1389fe7 = hmaster0_p & v1389fdd | !hmaster0_p & v1389de1;
assign v1445e34 = hlock5 & v1445e1f | !hlock5 & v1445e32;
assign v12ad50a = hmaster1_p & v12ad509 | !hmaster1_p & v845542;
assign v1445ea2 = hgrant4_p & v1445e02 | !hgrant4_p & v1445ea1;
assign a6536e = hgrant0_p & a65363 | !hgrant0_p & a6536d;
assign v12aeb23 = hbusreq2_p & v12aeb1b | !hbusreq2_p & v12aeb22;
assign v1216021 = hbusreq4_p & v845547 | !hbusreq4_p & v121601f;
assign v12afe66 = hmaster0_p & v12afe47 | !hmaster0_p & v12afe65;
assign v1389de4 = hmaster2_p & v1668c3b | !hmaster2_p & v845570;
assign v1445992 = hmastlock_p & v1445991 | !hmastlock_p & v845542;
assign v12157a5 = hmaster0_p & v121578e | !hmaster0_p & v12157a4;
assign v144544a = hlock2 & v1445446 | !hlock2 & v1445449;
assign v138a2f7 = hlock5_p & v151560a | !hlock5_p & v151561d;
assign v134d37e = hbusreq4_p & v134d273 | !hbusreq4_p & v134d37d;
assign v155298d = hbusreq3_p & v155298c | !hbusreq3_p & v1552d78;
assign d308f5 = hbusreq5_p & d308f4 | !hbusreq5_p & v84554e;
assign d300bf = hlock1_p & d2fe80 | !hlock1_p & v84555a;
assign f2f293 = hbusreq1_p & f2f292 | !hbusreq1_p & v845542;
assign f2e3fc = hbusreq2_p & f2e734 | !hbusreq2_p & f2e3fb;
assign v12157a8 = hbusreq2_p & v12157a1 | !hbusreq2_p & !v12157a7;
assign v1515780 = hgrant1_p & v151576a | !hgrant1_p & v151577f;
assign v134cd7e = hbusreq0 & v134cd7d | !hbusreq0 & v134d379;
assign v134d4df = hmaster2_p & v845542 | !hmaster2_p & v134d4ca;
assign v144606a = hgrant1_p & v1445fdb | !hgrant1_p & v1446069;
assign v12160bb = hmaster1_p & v121605f | !hmaster1_p & v1216082;
assign v14458d7 = hready & v14458d6 | !hready & v1446407;
assign v1214d53 = hbusreq2_p & v1214c02 | !hbusreq2_p & v1214d52;
assign v1552d98 = hready_p & v1552d96 | !hready_p & v1552d97;
assign d807a7 = hgrant0_p & d80760 | !hgrant0_p & d8073a;
assign v1445ede = hbusreq0 & v1445edd | !hbusreq0 & v1445eae;
assign v134ce97 = hbusreq3 & v134d240 | !hbusreq3 & v134ce88;
assign v134d372 = hbusreq1 & v134d371 | !hbusreq1 & v134d273;
assign v1216164 = hlock0_p & v1216014 | !hlock0_p & !v845542;
assign v16a1bbf = hmaster2_p & v16a1bbe | !hmaster2_p & v16a206f;
assign v14457c1 = hbusreq2 & v14457bf | !hbusreq2 & v14457c0;
assign v1445ddc = hbusreq2 & v1445dda | !hbusreq2 & v1445ddb;
assign v1214d56 = hmaster1_p & v1214d55 | !hmaster1_p & v1214d4b;
assign a656c5 = hgrant3_p & a65b07 | !hgrant3_p & a656c4;
assign v1216134 = hbusreq5_p & v121612d | !hbusreq5_p & v1216133;
assign f2f355 = hgrant1_p & v845570 | !hgrant1_p & !f2f354;
assign v1553094 = hbusreq3 & v1553092 | !hbusreq3 & v1553093;
assign d30104 = hlock4_p & d307e8 | !hlock4_p & !d30666;
assign v1214d8b = hbusreq5 & v1214d80 | !hbusreq5 & v1214d8a;
assign v12ae76c = hgrant3_p & v12ae6db | !hgrant3_p & v12ae76b;
assign v15161ff = hbusreq3 & v15161fe | !hbusreq3 & v1516804;
assign f2f2cd = hmaster2_p & f2f2cb | !hmaster2_p & !f2f21f;
assign v12165a5 = hmaster0_p & v1216599 | !hmaster0_p & v12165a4;
assign a66298 = hgrant4_p & a66297 | !hgrant4_p & !v845542;
assign d30612 = hlock5_p & v845542 | !hlock5_p & !d30611;
assign v12ad01b = hgrant2_p & v12ad5f5 | !hgrant2_p & v12acff4;
assign v1445360 = hmaster1_p & v144535f | !hmaster1_p & v14458fd;
assign f2e712 = hbusreq1_p & f2e711 | !hbusreq1_p & !v845542;
assign v138a44e = hmaster0_p & v138a344 | !hmaster0_p & v138a34b;
assign v121629c = hmaster0_p & v121629b | !hmaster0_p & v121619b;
assign v144660f = hgrant1_p & v1446429 | !hgrant1_p & v144660e;
assign v11e595f = hgrant2_p & bf1f59 | !hgrant2_p & v11e595d;
assign v121624b = hmaster0_p & v121624a | !hmaster0_p & !v1216223;
assign v11e593f = decide_p & v11e593e | !decide_p & v11e593d;
assign a65681 = hbusreq5 & a6565f | !hbusreq5 & a65680;
assign v134d446 = hlock2 & v134d3b5 | !hlock2 & v134d434;
assign f2f52c = hmaster0_p & f2f51a | !hmaster0_p & f2f229;
assign v1216712 = hbusreq2 & v121670e | !hbusreq2 & v1216711;
assign v1216241 = hgrant2_p & v1216229 | !hgrant2_p & v1216240;
assign v1553095 = hmaster2_p & v1553089 | !hmaster2_p & v845542;
assign v151571c = stateG2_p & v845542 | !stateG2_p & v88d3e4;
assign v1405ace = decide_p & v1405aba | !decide_p & v1405acd;
assign v10d409d = hmaster1_p & v10d409c | !hmaster1_p & v10d3ffb;
assign d2fc77 = hgrant2_p & d2fc28 | !hgrant2_p & d2fc76;
assign v12aec4a = hgrant2_p & v845542 | !hgrant2_p & v12aec49;
assign v1445fba = hbusreq5_p & v1445f85 | !hbusreq5_p & v1445fb9;
assign v16a1d58 = hgrant5_p & v845542 | !hgrant5_p & !v16a1d3a;
assign v1214de0 = hmaster1_p & v1214ddf | !hmaster1_p & v1215d2b;
assign d30781 = hbusreq4 & v845580 | !hbusreq4 & !v845542;
assign v1445fe3 = hlock0 & v1445fe2 | !hlock0 & v1445fe0;
assign v144535f = hmaster0_p & v1445909 | !hmaster0_p & v14458d3;
assign v12ad4ed = hmaster0_p & v12ad4e9 | !hmaster0_p & v12ad4ec;
assign v14458bd = hgrant5_p & v14458b8 | !hgrant5_p & !v14458b9;
assign v16a1d79 = hgrant5_p & v845542 | !hgrant5_p & !v16a2080;
assign v1214ff8 = hmaster2_p & v1214feb | !hmaster2_p & v1214ff7;
assign v1214fc3 = hgrant5_p & v845542 | !hgrant5_p & v1214fc2;
assign v138a07e = hbusreq5 & v1389ff2 | !hbusreq5 & v138a404;
assign v121655f = hgrant1_p & v845542 | !hgrant1_p & v121655e;
assign v1214f04 = hmaster0_p & v1214f00 | !hmaster0_p & v1214f03;
assign d3014c = hbusreq5_p & d3014b | !hbusreq5_p & d3014a;
assign v1215324 = hmaster1_p & v1215323 | !hmaster1_p & v121546f;
assign v14458fd = hmaster0_p & v14458f0 | !hmaster0_p & v14458fc;
assign bf1f76 = hmaster1_p & bf1f75 | !hmaster1_p & !bf1f52;
assign v134ce9c = hlock0 & v134ce9b | !hlock0 & v134ce9a;
assign d2fee2 = hmaster2_p & d2fece | !hmaster2_p & d2feba;
assign d306f8 = hmaster0_p & d306f7 | !hmaster0_p & d306d0;
assign a654ba = hmaster1_p & a65493 | !hmaster1_p & !a654b0;
assign d300fb = hlock4_p & d307d6 | !hlock4_p & d3065b;
assign v144589d = hbusreq0 & v1445894 | !hbusreq0 & v144589c;
assign v144614a = hmaster1_p & v144612a | !hmaster1_p & v1445ffc;
assign v16a19cf = hgrant3_p & v16a18de | !hgrant3_p & v16a19ce;
assign v1215725 = hbusreq5_p & v1215723 | !hbusreq5_p & !v1215724;
assign v16a2083 = hgrant0_p & v845542 | !hgrant0_p & v16a2073;
assign f2e4d5 = hready_p & f2e4d3 | !hready_p & f2e4d4;
assign v1215d2e = hmaster2_p & v1216588 | !hmaster2_p & v845542;
assign v14461ff = hlock3 & v144617b | !hlock3 & v14461fd;
assign v1668d6c = hmastlock_p & v1668d6b | !hmastlock_p & v845542;
assign v1445399 = hgrant2_p & v1445397 | !hgrant2_p & v1445398;
assign v1515704 = hbusreq2_p & v1515703 | !hbusreq2_p & v845542;
assign v1215b8a = hmaster2_p & v1215b76 | !hmaster2_p & v1215b80;
assign v144591b = hmaster0_p & v144591a | !hmaster0_p & v14458fc;
assign v1405b1d = hgrant5_p & v1405b17 | !hgrant5_p & !v1405b1c;
assign v12150ab = hmaster0_p & v1215092 | !hmaster0_p & v12150aa;
assign v121616d = hbusreq5_p & v121616b | !hbusreq5_p & v121616c;
assign v1215331 = hmaster1_p & v121505b | !hmaster1_p & !v121507b;
assign v144643a = hmaster2_p & v144639c | !hmaster2_p & v1446439;
assign v12af73c = decide_p & v12afe3e | !decide_p & v12afe76;
assign v1215bac = hbusreq4_p & v12160f2 | !hbusreq4_p & v845542;
assign v14462e8 = hmaster0_p & v14462e6 | !hmaster0_p & v14462e7;
assign v1214ede = hbusreq5_p & v1214edd | !hbusreq5_p & v1214edc;
assign v1215cbb = hbusreq1_p & v1216008 | !hbusreq1_p & !v845542;
assign a656a4 = hbusreq2 & a656a0 | !hbusreq2 & a656a3;
assign v16695c5 = hready_p & v845542 | !hready_p & v16695c4;
assign v1553143 = hmaster2_p & v1553140 | !hmaster2_p & v1553142;
assign v1215bfb = hbusreq0 & v1215bf5 | !hbusreq0 & v1215bfa;
assign v16a1d6a = hmaster2_p & v16a2080 | !hmaster2_p & v16a208a;
assign v16a1a22 = hbusreq2 & v16a19e6 | !hbusreq2 & v16a1a21;
assign v1405901 = hmaster1_p & v14058ec | !hmaster1_p & v1405900;
assign v16a1ae1 = hgrant2_p & v845542 | !hgrant2_p & v16a1ae0;
assign d30701 = hlock1_p & d30700 | !hlock1_p & !v845542;
assign v14461da = hlock2 & v144617b | !hlock2 & v14461d9;
assign v10d407e = hgrant2_p & v10d4015 | !hgrant2_p & v10d407d;
assign v16a1cdb = hbusreq3 & v16a1cd4 | !hbusreq3 & v16a1cda;
assign v134cd75 = hbusreq2_p & v134cd6d | !hbusreq2_p & v134cd74;
assign v1552f83 = hlock2 & v1552f80 | !hlock2 & v1552f82;
assign f2f352 = hbusreq5_p & f2f34e | !hbusreq5_p & f2f351;
assign v1215d85 = hmaster0_p & v1215d63 | !hmaster0_p & v12166fc;
assign v1389815 = hlock5_p & v1389814 | !hlock5_p & !v845542;
assign v1214d7e = hgrant2_p & v121657d | !hgrant2_p & v1214d7a;
assign v1552f80 = hgrant2_p & v1553380 | !hgrant2_p & v1552f7f;
assign d80789 = hmastlock_p & d80788 | !hmastlock_p & v845542;
assign v155350a = hbusreq5 & v1553508 | !hbusreq5 & v1553509;
assign f2f3a7 = hbusreq5_p & f2f3a5 | !hbusreq5_p & f2f3a6;
assign v12ad518 = hbusreq0_p & v1668cc4 | !hbusreq0_p & !v845542;
assign f2f3b3 = hmaster0_p & v84554c | !hmaster0_p & f2f3b2;
assign d30649 = hgrant4_p & a66284 | !hgrant4_p & a65382;
assign v12ad5e4 = hmaster2_p & v12ad4f0 | !hmaster2_p & !v12ad5ba;
assign d2fbd1 = hgrant4_p & d2fbce | !hgrant4_p & d2fbd0;
assign v15157d6 = hbusreq2 & v15157d5 | !hbusreq2 & v1516803;
assign d306ed = stateG3_2_p & v845542 | !stateG3_2_p & d306ec;
assign v138a3db = hbusreq5_p & v138a3da | !hbusreq5_p & !v845542;
assign v1445387 = hlock2 & v144537f | !hlock2 & v1445386;
assign v12164e7 = hmaster1_p & v16a2243 | !hmaster1_p & v845542;
assign d2fd13 = hmaster1_p & d3060a | !hmaster1_p & d2fcfe;
assign v1216267 = hbusreq2 & v1216259 | !hbusreq2 & v1216266;
assign v140587b = hlock3_p & v1405875 | !hlock3_p & v140587a;
assign v121607c = hbusreq2 & v1216076 | !hbusreq2 & v121607b;
assign v134d272 = hlock3_p & v134d241 | !hlock3_p & v134d271;
assign v1214f5f = hgrant2_p & v845542 | !hgrant2_p & v1214f5e;
assign v12ad544 = hmaster0_p & v12ad52d | !hmaster0_p & v12ad536;
assign d3087f = hmaster0_p & d30708 | !hmaster0_p & d306fd;
assign f2f4b6 = hmaster1_p & v845542 | !hmaster1_p & f2f4b5;
assign v12afe40 = hready_p & v845542 | !hready_p & v12afe3f;
assign v14453f8 = hlock3 & v14453f5 | !hlock3 & v14453f7;
assign v1515634 = hlock2_p & v151562a | !hlock2_p & v1515633;
assign v1215c70 = hgrant5_p & v845542 | !hgrant5_p & v1215c41;
assign v1445550 = hgrant2_p & v1445bec | !hgrant2_p & v144554f;
assign v1405850 = hmaster0_p & v1405840 | !hmaster0_p & v140584f;
assign v16a1a8a = hbusreq2_p & v16a196b | !hbusreq2_p & v16a1a89;
assign v16a1982 = hgrant2_p & v845542 | !hgrant2_p & v16a1980;
assign d3061b = hbusreq5_p & d3061a | !hbusreq5_p & v845542;
assign v1445fb1 = hmaster1_p & v1445fb0 | !hmaster1_p & v1445fae;
assign v134ceba = hbusreq2_p & v134ceb9 | !hbusreq2_p & v134d26e;
assign v151576b = hbusreq0_p & v1668d24 | !hbusreq0_p & v1515744;
assign v1445b2f = decide_p & v1445ae4 | !decide_p & v1445b2b;
assign v1405860 = hmastlock_p & v140585f | !hmastlock_p & !v845542;
assign d3020b = hmaster2_p & d30206 | !hmaster2_p & d3020a;
assign v1515622 = hbusreq2 & v1515621 | !hbusreq2 & v845542;
assign v15157ac = hgrant5_p & v845542 | !hgrant5_p & !v15157aa;
assign a6629d = hmaster0_p & a66291 | !hmaster0_p & a6629c;
assign v12ad4e9 = hbusreq0 & v12ad4e4 | !hbusreq0 & v845542;
assign v1405921 = hmaster1_p & v1405920 | !hmaster1_p & v14058b1;
assign a6546d = hbusreq1_p & a6546c | !hbusreq1_p & !a658cc;
assign v12af5a4 = hbusreq1 & v12afe55 | !hbusreq1 & v12afe61;
assign v1515712 = hbusreq1_p & v1515710 | !hbusreq1_p & v1515711;
assign v1445839 = hlock2 & v1445834 | !hlock2 & v1445838;
assign v1445446 = hbusreq2_p & v1446224 | !hbusreq2_p & v1445bb3;
assign d2fd44 = hbusreq2_p & d2fd27 | !hbusreq2_p & !d302eb;
assign d3079b = hbusreq5_p & d3079a | !hbusreq5_p & !d30799;
assign v1284c9e = hmaster2_p & v144639e | !hmaster2_p & v1284c9a;
assign v1515777 = hgrant5_p & v10d3ffa | !hgrant5_p & v1515775;
assign a646d8 = hbusreq3_p & a656c5 | !hbusreq3_p & a656d3;
assign v1215389 = hmaster1_p & v121537f | !hmaster1_p & v1215388;
assign v1216089 = hlock2_p & v1216087 | !hlock2_p & v1216088;
assign v138a316 = hlock5_p & v10d3ffd | !hlock5_p & !v845542;
assign d2fba5 = hbusreq2 & d2fba1 | !hbusreq2 & d2fba4;
assign v1405aad = hmaster2_p & v1405aab | !hmaster2_p & v1405aac;
assign v1214c85 = hbusreq2_p & v1214c83 | !hbusreq2_p & v1214c84;
assign v1389e2c = hlock5_p & v1389e2b | !hlock5_p & !v845542;
assign v1668c3c = hmaster2_p & v845570 | !hmaster2_p & v1668c3b;
assign v1445375 = hbusreq2 & v144536f | !hbusreq2 & v1445374;
assign v1216aa0 = hbusreq5 & v1216a9f | !hbusreq5 & v845542;
assign v134d4f5 = hgrant5_p & v134d4f4 | !hgrant5_p & v134d4f2;
assign a6540c = hmaster2_p & v845558 | !hmaster2_p & a65399;
assign f2f3bd = hbusreq5_p & f2f3bb | !hbusreq5_p & !f2f3bc;
assign v1215c18 = hbusreq5_p & v1215c11 | !hbusreq5_p & v1215c17;
assign v1446197 = hlock2 & v144617b | !hlock2 & v1446196;
assign f2f401 = hbusreq2_p & f2f3ff | !hbusreq2_p & f2f400;
assign d305e4 = hbusreq3 & d305dc | !hbusreq3 & d305e3;
assign v12153e4 = hbusreq4_p & v12153e3 | !hbusreq4_p & v845542;
assign v10d429e = hgrant1_p & v10d3fe5 | !hgrant1_p & !v10d429d;
assign v14463c8 = hbusreq0 & v14463c6 | !hbusreq0 & v14463c7;
assign v1445a6f = hbusreq2_p & v1445a34 | !hbusreq2_p & v1445a6e;
assign v14459c0 = hlock0_p & v14459be | !hlock0_p & v14459bf;
assign d3067f = hbusreq2_p & d3067e | !hbusreq2_p & d3067d;
assign v12af3ae = hready_p & v845542 | !hready_p & v12af3ad;
assign v1405b52 = hmaster1_p & v1405b51 | !hmaster1_p & v1405af0;
assign v144587a = hmaster2_p & v144639c | !hmaster2_p & v1445879;
assign v14465ab = hmaster1_p & v14465aa | !hmaster1_p & v1446436;
assign v1446640 = hmaster2_p & v14465b0 | !hmaster2_p & v144663f;
assign v121618d = hgrant5_p & v845542 | !hgrant5_p & v1216112;
assign v10d4278 = hgrant2_p & v10d4054 | !hgrant2_p & !v10d4277;
assign v15157fd = hbusreq5_p & v15157fc | !hbusreq5_p & !v15157ac;
assign v151562d = hburst1 & a66293 | !hburst1 & v151562c;
assign v1214f65 = hready_p & v1214f3d | !hready_p & v1214f64;
assign v16a13c8 = hmaster1_p & v16a13c7 | !hmaster1_p & !v16a2672;
assign f2eda0 = decide_p & f2ed94 | !decide_p & f2f23c;
assign v16a1d70 = hgrant2_p & v845542 | !hgrant2_p & v16a1d6f;
assign v1216273 = hmaster0_p & v12161f7 | !hmaster0_p & v1216038;
assign f2f3a0 = hgrant5_p & f2f2a4 | !hgrant5_p & !f2f39f;
assign v16a12ec = hgrant5_p & v845542 | !hgrant5_p & v16a12eb;
assign v138a397 = hbusreq2_p & v138a342 | !hbusreq2_p & v138a396;
assign v1446494 = hbusreq0_p & v1446480 | !hbusreq0_p & v1446476;
assign v16a1da2 = hmaster1_p & v845542 | !hmaster1_p & v16a2672;
assign a6561d = hgrant4_p & a662a9 | !hgrant4_p & !a65370;
assign v144649a = hlock0_p & v1446398 | !hlock0_p & v1446494;
assign v1445889 = hmaster2_p & v1445888 | !hmaster2_p & v1445885;
assign v1405ae0 = hlock5_p & v1405ade | !hlock5_p & !v1405adf;
assign v1552fd8 = hbusreq3_p & v1552f8d | !hbusreq3_p & v1552fd7;
assign v1445498 = hmaster1_p & v144547f | !hmaster1_p & v1446290;
assign v12162d0 = hmaster1_p & v121622b | !hmaster1_p & !v121624b;
assign v1445928 = hbusreq5 & v1445926 | !hbusreq5 & v1445927;
assign d2fb02 = hgrant4_p & v845558 | !hgrant4_p & d2fb01;
assign v1389d77 = decide_p & v1389d76 | !decide_p & v845542;
assign v1446131 = hlock2 & v1446125 | !hlock2 & v144612f;
assign v134d4b0 = hgrant2_p & v134d364 | !hgrant2_p & v134d4af;
assign d30957 = hlock0_p & d3094f | !hlock0_p & v845542;
assign v12162fc = hbusreq1_p & v12162fb | !hbusreq1_p & v845547;
assign v134cd66 = hgrant1_p & v845542 | !hgrant1_p & v134cd65;
assign v1215743 = hmaster2_p & v1215734 | !hmaster2_p & v1215b9c;
assign v138937d = hbusreq0 & v1389fdd | !hbusreq0 & v1389de1;
assign v134d42f = hgrant5_p & v845542 | !hgrant5_p & v134d42e;
assign d3070a = hmaster1_p & d30709 | !hmaster1_p & !d30706;
assign v1446151 = hlock3 & v1446148 | !hlock3 & v1446150;
assign v1668c67 = hbusreq5_p & v1668c65 | !hbusreq5_p & !v1668c66;
assign v1214ce5 = decide_p & v1214ca2 | !decide_p & v1214ce4;
assign v1445e5e = hbusreq4_p & v1445e5d | !hbusreq4_p & v1446406;
assign v1215368 = hmaster2_p & v845547 | !hmaster2_p & v1215366;
assign v12160e4 = hmaster1_p & v12160e3 | !hmaster1_p & v12160e0;
assign f2f421 = hbusreq5_p & f2f3a0 | !hbusreq5_p & f2f420;
assign v1215cae = hbusreq1_p & v121610d | !hbusreq1_p & v1215cad;
assign v15157a4 = hbusreq5_p & v15157a2 | !hbusreq5_p & !v15157a3;
assign v1446613 = hgrant1_p & v144641d | !hgrant1_p & v14465f2;
assign v1284d4c = hgrant1_p & v140583c | !hgrant1_p & v1284d4b;
assign v1445b4f = hmaster1_p & v1445b4e | !hmaster1_p & v144590e;
assign d3090e = hmaster0_p & d3090c | !hmaster0_p & d3090d;
assign v1445a41 = hgrant5_p & v14458ff | !hgrant5_p & v1445a40;
assign v121611a = hgrant5_p & v121601d | !hgrant5_p & v1216118;
assign v1215ca4 = hbusreq1_p & v12160fc | !hbusreq1_p & v12160f4;
assign v1446275 = hbusreq2_p & v1446272 | !hbusreq2_p & v1446274;
assign v144611e = hmaster1_p & v144611d | !hmaster1_p & v1445fde;
assign v1445a06 = hbusreq5_p & v14459fe | !hbusreq5_p & v1445a05;
assign v1516106 = decide_p & v1516105 | !decide_p & v845542;
assign v16a1c9e = hmaster2_p & v16a1c99 | !hmaster2_p & v845542;
assign v12147fd = hmaster1_p & v12147ed | !hmaster1_p & !v1215d9b;
assign v1214cbb = hgrant4_p & d2fbe5 | !hgrant4_p & v845572;
assign a65928 = hbusreq3 & a65920 | !hbusreq3 & a65927;
assign v121659c = hgrant1_p & v1216a96 | !hgrant1_p & v121659b;
assign v134d28d = hgrant1_p & v845542 | !hgrant1_p & v134d28c;
assign v1445a7e = hgrant5_p & v1445a7b | !hgrant5_p & v1445a7d;
assign d2fb5d = hbusreq3 & d2fb56 | !hbusreq3 & d2fb5c;
assign v1405885 = hmaster0_p & v1405856 | !hmaster0_p & v1405855;
assign v1445af6 = hmaster1_p & v1445af5 | !hmaster1_p & v14458fd;
assign v1445efa = hbusreq2_p & v1445ef2 | !hbusreq2_p & v1445ef9;
assign v151573c = hmaster0_p & v1515732 | !hmaster0_p & v151573b;
assign f2ec21 = hlock1_p & f2ec20 | !hlock1_p & !v845542;
assign d3018f = hmaster1_p & d3018e | !hmaster1_p & d30918;
assign v16a16ab = hgrant2_p & v845542 | !hgrant2_p & !v16a16aa;
assign v1515834 = hgrant5_p & v1515832 | !hgrant5_p & v1515833;
assign v1445904 = hmaster1_p & v1445903 | !hmaster1_p & v14458fd;
assign d8077b = hgrant4_p & d8077a | !hgrant4_p & !v845542;
assign v10d4271 = hgrant2_p & v10d4018 | !hgrant2_p & v10d4270;
assign d2f9a2 = hmaster2_p & d3068e | !hmaster2_p & d2f9a1;
assign v121609e = hbusreq2 & v121608f | !hbusreq2 & v121609d;
assign v15530ea = hlock3 & v155341e | !hlock3 & v15530e9;
assign d2fbff = hgrant2_p & d2fbc9 | !hgrant2_p & d2fbfe;
assign a65b3c = hgrant3_p & a65b28 | !hgrant3_p & a65b3b;
assign f2e505 = jx1_p & f2e4e3 | !jx1_p & f2e504;
assign v1215cd1 = hgrant5_p & v845570 | !hgrant5_p & v1215cd0;
assign v14464a4 = hmaster2_p & v845542 | !hmaster2_p & v144646e;
assign f2f332 = hmaster1_p & f2f2de | !hmaster1_p & !f2f330;
assign v1214c2b = hmaster2_p & v1214c29 | !hmaster2_p & v1214c2a;
assign v138a481 = hbusreq2_p & v138a47c | !hbusreq2_p & v138a480;
assign v1284cc4 = hlock2_p & v1284cc3 | !hlock2_p & v1405886;
assign d8075b = stateA1_p & d80756 | !stateA1_p & d8075a;
assign v121604c = hmaster2_p & v1216049 | !hmaster2_p & v121604b;
assign v12160f0 = hgrant4_p & v12160ed | !hgrant4_p & v12160ef;
assign d3025b = hbusreq2_p & d30252 | !hbusreq2_p & !d3025a;
assign v16a1d04 = hbusreq3_p & v16a1cc9 | !hbusreq3_p & v16a1d03;
assign v12153bc = hlock0_p & v1215bb0 | !hlock0_p & v12153bb;
assign v1214d14 = hbusreq0 & v1214d13 | !hbusreq0 & v16a2243;
assign v16693a0 = hmaster2_p & a6587e | !hmaster2_p & !v166939f;
assign v12161fc = hmaster0_p & v12161d3 | !hmaster0_p & v12161fb;
assign a653e3 = hgrant5_p & a6586d | !hgrant5_p & a653e2;
assign v144628b = hbusreq3 & v1446277 | !hbusreq3 & v144628a;
assign v1446285 = hmaster1_p & v144626e | !hmaster1_p & v144627e;
assign v138a3e3 = hlock5_p & v151580c | !hlock5_p & !v845542;
assign v1445a0b = hbusreq0_p & v1445a0a | !hbusreq0_p & v14465bb;
assign d307ce = hbusreq0_p & v845542 | !hbusreq0_p & d307ae;
assign a653ac = hbusreq1 & a65863 | !hbusreq1 & a6587e;
assign v140585e = decide_p & v140585d | !decide_p & v1405852;
assign v14058db = hmaster2_p & v140583d | !hmaster2_p & v14058c5;
assign v144634a = hlock2 & v1446346 | !hlock2 & v1446349;
assign v1216290 = hbusreq2 & v121628c | !hbusreq2 & v121628f;
assign f2f39f = hmaster2_p & f2f347 | !hmaster2_p & f2f369;
assign v1445ba7 = decide_p & v1446260 | !decide_p & v1445ba6;
assign d301aa = hbusreq2_p & d301a1 | !hbusreq2_p & d301a9;
assign v10d4288 = hlock0_p & v10d4287 | !hlock0_p & v10d3fd8;
assign d301a3 = hlock5_p & d301a2 | !hlock5_p & d30954;
assign v14458dd = hbusreq4 & v14458d6 | !hbusreq4 & v14458dc;
assign v1668c2a = hbusreq5_p & v1668c28 | !hbusreq5_p & v1668c29;
assign d2fea2 = hmaster0_p & d2fea0 | !hmaster0_p & d2fea1;
assign d307c3 = hbusreq0 & d307ba | !hbusreq0 & d307c2;
assign f2e4de = hbusreq2_p & f2e4d2 | !hbusreq2_p & f2e4dd;
assign v151575e = hbusreq0 & v1515753 | !hbusreq0 & v151575d;
assign v1405ae9 = hbusreq0_p & v845542 | !hbusreq0_p & !d3070c;
assign v12153bf = hmaster0_p & v12153ba | !hmaster0_p & v12153be;
assign v1216ae3 = hlock0_p & v1216ab0 | !hlock0_p & !v845542;
assign a65465 = hmaster0_p & a658e8 | !hmaster0_p & a658b7;
assign d301db = hlock5_p & d301d9 | !hlock5_p & !d301da;
assign v1445e77 = hgrant5_p & v1445e71 | !hgrant5_p & v1445e76;
assign v144624c = hgrant5_p & v144624a | !hgrant5_p & !v144624b;
assign v1216314 = hbusreq3 & v1216313 | !hbusreq3 & v845542;
assign v14058bc = hmaster0_p & v1405896 | !hmaster0_p & v14058bb;
assign v151578a = stateG3_2_p & v845542 | !stateG3_2_p & v1515789;
assign v151566b = hmaster0_p & v151565b | !hmaster0_p & v151566a;
assign v12162c9 = hmaster0_p & v121622b | !hmaster0_p & v1216236;
assign v1214d76 = hlock2_p & v1214d75 | !hlock2_p & v1214d36;
assign d306ce = hmaster2_p & d306cb | !hmaster2_p & d306cd;
assign d2fb2e = hgrant2_p & d3012a | !hgrant2_p & d2fb19;
assign d30203 = hbusreq1 & d30700 | !hbusreq1 & v845542;
assign v16a1d2d = hmaster0_p & v16a2234 | !hmaster0_p & v16a2243;
assign f2f40b = hmaster1_p & f2f3f9 | !hmaster1_p & !f2f330;
assign v1215b97 = hlock4_p & v845547 | !hlock4_p & !v845542;
assign v1214c21 = hmaster1_p & v1214bf1 | !hmaster1_p & v1214bcf;
assign v12163a6 = hmaster2_p & v12163a5 | !hmaster2_p & v1216ac7;
assign v12164de = hlock0_p & v845570 | !hlock0_p & v12164dd;
assign v1446485 = hgrant1_p & v845542 | !hgrant1_p & v1446484;
assign v1445e7f = hmaster2_p & v1446606 | !hmaster2_p & v1445df5;
assign v14458e9 = hmaster2_p & v14458e8 | !hmaster2_p & v14458e5;
assign v1214c66 = hbusreq1 & v1215354 | !hbusreq1 & v845542;
assign d30717 = hburst0 & d30715 | !hburst0 & d30716;
assign v121615f = hlock1_p & v121615c | !hlock1_p & v121615e;
assign v1552d62 = hgrant2_p & v1553380 | !hgrant2_p & v1552d61;
assign v16a19de = hmaster2_p & v16a19d1 | !hmaster2_p & !v845542;
assign v14459e4 = hmaster2_p & v144639c | !hmaster2_p & v14458eb;
assign v10d4092 = hgrant5_p & v10d400e | !hgrant5_p & v10d4091;
assign v1668d17 = hmaster0_p & v1668d15 | !hmaster0_p & v1668d16;
assign v1446409 = hlock4 & v1446407 | !hlock4 & v1446408;
assign d2f9cf = hbusreq5_p & d2f9c9 | !hbusreq5_p & d2f99e;
assign a654a9 = hbusreq2_p & a6549a | !hbusreq2_p & a6549b;
assign v1446136 = hmaster0_p & v14460a5 | !hmaster0_p & v1445fe3;
assign v1445abc = hmaster0_p & v14458a2 | !hmaster0_p & v144639c;
assign v1215415 = hlock2_p & v1215414 | !hlock2_p & v1215411;
assign a65443 = hbusreq5_p & a65440 | !hbusreq5_p & !a65441;
assign d3010c = hbusreq5_p & d3010b | !hbusreq5_p & d3010a;
assign v12160df = hmaster2_p & v12160dc | !hmaster2_p & v12160de;
assign d2fb5e = hlock3_p & d2fb5d | !hlock3_p & v84554a;
assign d807b8 = decide_p & v845542 | !decide_p & d807b7;
assign d2fb71 = hmaster2_p & d2fb6a | !hmaster2_p & d2fb70;
assign v16a2098 = hgrant2_p & v845542 | !hgrant2_p & !v16a2096;
assign v1216113 = hgrant5_p & v1215ff2 | !hgrant5_p & v1216112;
assign v134d276 = hmaster1_p & v134d275 | !hmaster1_p & v845542;
assign d307b4 = hbusreq1 & d307b3 | !hbusreq1 & v845542;
assign f2f3df = hbusreq2_p & f2f3dd | !hbusreq2_p & !f2f3de;
assign v134d393 = hbusreq1 & v134d391 | !hbusreq1 & v134d392;
assign d80795 = hbusreq0_p & d80733 | !hbusreq0_p & !d8078a;
assign v12163aa = hmaster1_p & v121639f | !hmaster1_p & !v12163a9;
assign v11e5966 = hgrant0_p & v11e593a | !hgrant0_p & !v845542;
assign d301d3 = hgrant5_p & d301bb | !hgrant5_p & d301d2;
assign d30121 = hgrant2_p & d30113 | !hgrant2_p & !d30120;
assign v1445dfd = hlock1 & v1445dfc | !hlock1 & v1445dfb;
assign v10d401a = hbusreq4_p & v10d3fd5 | !hbusreq4_p & !v10d3fd4;
assign v134d425 = hbusreq1 & v134d37f | !hbusreq1 & v134d380;
assign v1446664 = hmaster0_p & v14465b8 | !hmaster0_p & v1446663;
assign v1405b13 = hgrant4_p & v1405abb | !hgrant4_p & v1405b12;
assign v1668d2e = hgrant4_p & v1668d26 | !hgrant4_p & a6537e;
assign v16695a9 = hbusreq3_p & v16695a8 | !hbusreq3_p & !v1668c39;
assign v1445424 = hlock2 & v144541f | !hlock2 & v1445423;
assign v1214d17 = hgrant2_p & v1214d16 | !hgrant2_p & v1214d05;
assign v1214c80 = hmaster0_p & v845542 | !hmaster0_p & v1215360;
assign v14463b1 = hmastlock_p & v845588 | !hmastlock_p & !v845542;
assign v1214d5d = hbusreq5_p & v1214bcc | !hbusreq5_p & v1214d5c;
assign d2fba8 = hlock2_p & d2fba6 | !hlock2_p & d2fba7;
assign v12ad60f = hmaster2_p & v12ad5bb | !hmaster2_p & v845542;
assign v12acfc5 = hmaster0_p & v12ad67b | !hmaster0_p & v12acfc4;
assign v12ad501 = hmaster2_p & v12ad4f0 | !hmaster2_p & !v12ad4f6;
assign v12ad65f = hmaster1_p & v12ad65e | !hmaster1_p & v845542;
assign v1215cb9 = hbusreq1_p & v1216000 | !hbusreq1_p & !v845542;
assign d2fbc0 = hbusreq2_p & d2fbbf | !hbusreq2_p & d2fbbb;
assign v134d3e6 = decide_p & v134d3cf | !decide_p & v134d3ba;
assign v1214cfe = hbusreq4_p & v1214c2a | !hbusreq4_p & !v1214cf1;
assign v1284d06 = decide_p & v1284ce8 | !decide_p & v1284d05;
assign d30280 = hlock5_p & d3027e | !hlock5_p & !d3027f;
assign v10d42a3 = hgrant2_p & v10d4015 | !hgrant2_p & v10d42a2;
assign v1445ac0 = hlock2 & v1445abf | !hlock2 & v1445aba;
assign v16a1845 = hbusreq2 & v16a1841 | !hbusreq2 & v16a1844;
assign v1405b16 = hgrant5_p & v1405abd | !hgrant5_p & v1405b15;
assign v121532c = hgrant2_p & v1215329 | !hgrant2_p & v121532b;
assign d305fc = hmaster2_p & a66278 | !hmaster2_p & d305fb;
assign v14458d5 = hmaster0_p & v14458d3 | !hmaster0_p & v14458d4;
assign v134cf70 = jx0_p & v134cd45 | !jx0_p & v134cf6f;
assign bf1fa2 = hgrant5_p & v845542 | !hgrant5_p & !bf1fa1;
assign v144633a = stateG10_5_p & v144668d | !stateG10_5_p & v1446339;
assign v12ad1b1 = hready_p & v12ad140 | !hready_p & v12ad1b0;
assign v14460ed = hbusreq2_p & v14460e8 | !hbusreq2_p & v14460ec;
assign v16a1acb = hbusreq2_p & v16a1f97 | !hbusreq2_p & v16a1aca;
assign v16a12c2 = hbusreq2 & v16a12c0 | !hbusreq2 & v16a12c1;
assign v13891a2 = hlock5_p & v13891a1 | !hlock5_p & v845542;
assign v12161ad = hbusreq0 & v1216193 | !hbusreq0 & v12161ac;
assign v15157dd = hbusreq0 & v15157d9 | !hbusreq0 & v15157dc;
assign v15161d1 = hmaster0_p & v1668da6 | !hmaster0_p & v15161d0;
assign v144580b = hmaster1_p & v144580a | !hmaster1_p & v1445eaa;
assign v15157ad = hbusreq5_p & v15157ab | !hbusreq5_p & !v15157ac;
assign v1668d36 = hgrant1_p & v1668d23 | !hgrant1_p & v1668d35;
assign v1445dd8 = hmaster1_p & v1445db9 | !hmaster1_p & v1445dd1;
assign f2f22a = hgrant1_p & v845570 | !hgrant1_p & !v845542;
assign v1215c90 = hbusreq5_p & v1215c8e | !hbusreq5_p & !v1215c8f;
assign v1445a24 = hlock0_p & v1445a22 | !hlock0_p & v1445a23;
assign v16a1e00 = hmaster1_p & v16a2243 | !hmaster1_p & v16a1f96;
assign v16a1cf2 = hbusreq2_p & v16a1bdd | !hbusreq2_p & v16a1cf1;
assign d301be = hmaster2_p & d306d4 | !hmaster2_p & d301bc;
assign f2f419 = hmaster1_p & f2f418 | !hmaster1_p & f2f393;
assign v14462ec = hmaster2_p & v144663f | !hmaster2_p & v14465d2;
assign v1284ca4 = hbusreq4_p & v1284ca3 | !hbusreq4_p & v144639e;
assign d2fbaf = hbusreq5 & d2fb98 | !hbusreq5 & d2fbae;
assign v12aeb1d = hbusreq0 & v12afda2 | !hbusreq0 & v12aeb1c;
assign d2fc13 = hgrant2_p & d2fbc9 | !hgrant2_p & d2fc12;
assign v14462eb = hmaster2_p & v1446634 | !hmaster2_p & v1446410;
assign v12ad006 = hgrant5_p & v12ad501 | !hgrant5_p & v12ad005;
assign d2fbdd = hbusreq1 & d2fb4e | !hbusreq1 & d2fb58;
assign f2e279 = hmaster1_p & v845542 | !hmaster1_p & f2e278;
assign d2fb09 = hgrant4_p & v845558 | !hgrant4_p & d2fb08;
assign bf1f53 = hmaster2_p & v84556a | !hmaster2_p & !bf1f52;
assign v12afe63 = hgrant5_p & v845542 | !hgrant5_p & v12afe62;
assign v1668dd1 = hbusreq0 & v1668dcd | !hbusreq0 & v1668dd0;
assign v134cd6e = hbusreq1 & v134cd56 | !hbusreq1 & v134cd57;
assign v12ad4c7 = hready_p & v12ad32d | !hready_p & v12ad4c6;
assign v16a19d3 = hbusreq5_p & v16a1840 | !hbusreq5_p & v16a19d2;
assign v1214cdf = hgrant5_p & d2fbe5 | !hgrant5_p & v1214cbc;
assign v16a1d40 = hgrant1_p & v84554d | !hgrant1_p & v16a1bc8;
assign v10d40ba = locked_p & v10d3fd2 | !locked_p & v10d3fd4;
assign d2fcd8 = hbusreq2_p & v845542 | !hbusreq2_p & d302d6;
assign v134d214 = hbusreq1 & v134d1ee | !hbusreq1 & v134d1ef;
assign v1216046 = decide_p & v1216032 | !decide_p & v1216045;
assign v134ce77 = hbusreq3 & v134ce76 | !hbusreq3 & v134d276;
assign v151572c = hgrant4_p & v1668d26 | !hgrant4_p & v151572b;
assign v1668d6a = hburst1 & a66293 | !hburst1 & v1668d69;
assign v1445e3f = hbusreq5_p & v1445e3c | !hbusreq5_p & v1445e3e;
assign v1214c46 = hbusreq1_p & v1214c45 | !hbusreq1_p & v16a1c95;
assign v1446091 = hbusreq0 & v1446090 | !hbusreq0 & v144607f;
assign v14466da = hmaster1_p & v14463f6 | !hmaster1_p & v14463ef;
assign v1215fbc = hmaster1_p & v1215fbb | !hmaster1_p & v12164e1;
assign v14457c0 = hlock2 & v1445786 | !hlock2 & v14457be;
assign v144542c = hmaster1_p & v1445414 | !hmaster1_p & v1445b7a;
assign f2f2a9 = hbusreq1 & a6588d | !hbusreq1 & v845542;
assign v12153d8 = hlock4_p & v12153d6 | !hlock4_p & !v12153d7;
assign v1445827 = hbusreq2_p & v144581f | !hbusreq2_p & v1445826;
assign v10d406b = hgrant5_p & v10d4029 | !hgrant5_p & !v10d406a;
assign a6586c = hbusreq4_p & a6586b | !hbusreq4_p & v845542;
assign a6629e = hmaster1_p & a6628e | !hmaster1_p & a6629d;
assign a65461 = hmaster1_p & a65460 | !hmaster1_p & a1db63;
assign v14458a2 = hmaster2_p & v144639c | !hmaster2_p & v144586f;
assign v1553230 = hgrant4_p & v155322f | !hgrant4_p & v845542;
assign v1214fec = hmaster2_p & v1214fe6 | !hmaster2_p & v1214feb;
assign v1445f07 = hbusreq0 & v1445f06 | !hbusreq0 & v1445e84;
assign v1216012 = hbusreq1 & v1216568 | !hbusreq1 & v845542;
assign v1216aa5 = stateG3_2_p & v845542 | !stateG3_2_p & !v1216aa4;
assign v121619f = hgrant5_p & v845542 | !hgrant5_p & v1216175;
assign v1445a3b = hmaster2_p & v144599d | !hmaster2_p & v14459df;
assign v1214fe4 = hbusreq4_p & v1214fe3 | !hbusreq4_p & v845542;
assign v12164e3 = hbusreq5_p & v12164cf | !hbusreq5_p & v16a2243;
assign v1216558 = hgrant4_p & v1216524 | !hgrant4_p & v1216557;
assign v16693b1 = decide_p & v16693b0 | !decide_p & !v845542;
assign v12ad585 = hmaster1_p & v12ad56e | !hmaster1_p & v12ad54f;
assign v138a35a = hmaster1_p & v138a359 | !hmaster1_p & v138a341;
assign v1445d8f = hmaster2_p & v14463b9 | !hmaster2_p & v1445f97;
assign v15157a0 = hbusreq0 & v1515799 | !hbusreq0 & v151579f;
assign v1445bad = hmaster0_p & v14463c5 | !hmaster0_p & v144639c;
assign v1284ca8 = hmaster1_p & v1284c98 | !hmaster1_p & v1284ca7;
assign v14464a0 = hbusreq5_p & v144648b | !hbusreq5_p & v144649f;
assign v14465dd = hgrant5_p & v14465d5 | !hgrant5_p & v14465dc;
assign v16a2675 = hbusreq5_p & v16a2674 | !hbusreq5_p & v845542;
assign v1445a69 = hbusreq2_p & v1445a63 | !hbusreq2_p & v1445a68;
assign v1445ed2 = hmaster1_p & v14465aa | !hmaster1_p & v1445e1b;
assign d2fbef = stateG10_5_p & d2fbee | !stateG10_5_p & d2fbe1;
assign v121481b = hbusreq3_p & v1214f66 | !hbusreq3_p & v121481a;
assign v12160ce = hbusreq5 & v12160b9 | !hbusreq5 & v12160cd;
assign v144669c = hgrant1_p & v144641f | !hgrant1_p & v144669b;
assign a658d3 = hburst0 & v10d3fd6 | !hburst0 & a658d2;
assign v1216aad = hready & v1446397 | !hready & v1216aac;
assign v10d3fd4 = hmastlock_p & v10d3fd2 | !hmastlock_p & v10d3fd3;
assign v14453ec = hbusreq2 & v14453e3 | !hbusreq2 & v14453eb;
assign v15157a9 = hgrant1_p & v15157a8 | !hgrant1_p & v1515794;
assign v1215dde = jx2_p & v1215ddd | !jx2_p & v845542;
assign v1445eba = hlock0 & v1445eb9 | !hlock0 & v1445eb5;
assign v121670b = hmaster0_p & v1216702 | !hmaster0_p & v12166f7;
assign d2fd41 = hbusreq5 & d2fd3e | !hbusreq5 & d2fd40;
assign v12af5a5 = hgrant0_p & d30645 | !hgrant0_p & v845542;
assign v12ad4c0 = hmaster2_p & d30690 | !hmaster2_p & v12ad4bf;
assign v134cd5e = hlock0 & v134cd5d | !hlock0 & v134cd5c;
assign v15156ba = hbusreq1_p & v1515654 | !hbusreq1_p & v15156b9;
assign v1445feb = hmaster0_p & v144639c | !hmaster0_p & v1445fea;
assign v12166e8 = hgrant0_p & v12166e7 | !hgrant0_p & v845542;
assign f2f440 = hbusreq2_p & f2f43e | !hbusreq2_p & !f2f43f;
assign v1215c46 = hmaster0_p & v1215bfb | !hmaster0_p & v1215c45;
assign v16a1e52 = hmaster1_p & v16a1e27 | !hmaster1_p & v16a1f96;
assign v1445a5e = hbusreq2_p & v1445a34 | !hbusreq2_p & v1445a5d;
assign v1215372 = hmaster1_p & v1215371 | !hmaster1_p & v845542;
assign v1668ccb = stateA1_p & a66272 | !stateA1_p & !v1668cca;
assign v12ad531 = hbusreq0 & v12ad530 | !hbusreq0 & !v845542;
assign v1445bab = hmaster1_p & v1445baa | !hmaster1_p & v845542;
assign f2f229 = hgrant5_p & v845542 | !hgrant5_p & !f2f228;
assign d307a8 = hmaster2_p & d30796 | !hmaster2_p & d30655;
assign v1215343 = hgrant3_p & v1215112 | !hgrant3_p & !v1215342;
assign a65885 = stateA1_p & v845542 | !stateA1_p & a65884;
assign a65459 = hmaster0_p & a653ea | !hmaster0_p & a65360;
assign stateG3_2 = !v1445558;
assign v12af1ba = hmaster2_p & d30690 | !hmaster2_p & !v12af1b9;
assign v1389fb8 = hlock5_p & d3060a | !hlock5_p & v845542;
assign v1553101 = hlock3 & v155321a | !hlock3 & v1553100;
assign v845564 = hmaster0_p & v845542 | !hmaster0_p & !v845542;
assign v1553383 = hgrant1_p & v845542 | !hgrant1_p & v1553382;
assign f2f340 = hbusreq5 & f2f32c | !hbusreq5 & f2f33f;
assign v1215455 = hmaster0_p & v121543b | !hmaster0_p & v1215439;
assign v12162ba = hgrant2_p & v12162b8 | !hgrant2_p & v12162b9;
assign d2fd48 = hbusreq5 & d2fd45 | !hbusreq5 & d2fd47;
assign v16a1bbc = hbusreq1 & v16a1bbb | !hbusreq1 & v16a206e;
assign v12acffa = hgrant0_p & v12af9bc | !hgrant0_p & !v12acff9;
assign d3068d = hbusreq5_p & d305f6 | !hbusreq5_p & !d3068c;
assign v14459bc = hready & v14465ad | !hready & v144639c;
assign v1214d6b = hbusreq3 & v1214d64 | !hbusreq3 & v1214d6a;
assign v1216afb = hlock5_p & v1216afa | !hlock5_p & !v845542;
assign v1552f64 = hgrant1_p & v845542 | !hgrant1_p & v1552f63;
assign v1445555 = hbusreq3_p & v144554c | !hbusreq3_p & v1445554;
assign v134cd87 = hbusreq2 & v134cd85 | !hbusreq2 & v134cd86;
assign v12162a0 = hbusreq2 & v1216296 | !hbusreq2 & v121629f;
assign v138a326 = stateA1_p & v138a325 | !stateA1_p & !v1180b7b;
assign v16a1daa = hbusreq2_p & v16a1d0e | !hbusreq2_p & v16a1da9;
assign d306e6 = hmaster2_p & d306cb | !hmaster2_p & d306d7;
assign d2fae3 = hmaster2_p & d2fadc | !hmaster2_p & d2fae2;
assign v134d4aa = hgrant5_p & v134d4a9 | !hgrant5_p & v134d375;
assign v134d36a = hmaster2_p & v134d273 | !hmaster2_p & v845542;
assign v1445a8c = hbusreq2_p & v1445a84 | !hbusreq2_p & v1445a8b;
assign v121628c = hbusreq2_p & v1216287 | !hbusreq2_p & !v121628b;
assign v1405847 = hmaster2_p & v1405844 | !hmaster2_p & v1405845;
assign v134d51d = hbusreq2_p & v134d515 | !hbusreq2_p & v134d51c;
assign v1445803 = hmaster0_p & v1445802 | !hmaster0_p & v144639c;
assign v14463d9 = hlock1 & v14463d8 | !hlock1 & v14463a0;
assign v1405b67 = jx2_p & v85e750 | !jx2_p & v1405b66;
assign f2f453 = hbusreq0 & f2f450 | !hbusreq0 & f2f452;
assign v134cdca = decide_p & v134d3ce | !decide_p & v134cdc9;
assign v16a1332 = hbusreq2 & v16a132b | !hbusreq2 & v16a1331;
assign d308b2 = hgrant2_p & d3085f | !hgrant2_p & d308ae;
assign v15157d1 = hmaster0_p & v15157b3 | !hmaster0_p & v15157d0;
assign v16a1d7a = hbusreq0 & v16a209a | !hbusreq0 & v16a1d79;
assign v1214d6e = hmaster1_p & v1214d6d | !hmaster1_p & v1214c39;
assign v15534ee = hbusreq0 & v15534ed | !hbusreq0 & v1553218;
assign v12af98b = hbusreq5_p & v12afdb0 | !hbusreq5_p & v12af98a;
assign v138a32a = stateA1_p & v138a329 | !stateA1_p & !v845542;
assign v1446416 = hmaster2_p & v1446403 | !hmaster2_p & v1446415;
assign v1552d82 = hgrant5_p & v1552d81 | !hgrant5_p & v1552d7f;
assign bf1f6b = hgrant5_p & v845570 | !hgrant5_p & bf1f6a;
assign v1389464 = hbusreq2 & v1389463 | !hbusreq2 & v138a404;
assign v16695c9 = jx1_p & v16695aa | !jx1_p & v16695c8;
assign v16a132e = hbusreq0 & v16a132d | !hbusreq0 & v845542;
assign v144582f = hmaster1_p & v1445805 | !hmaster1_p & v1445ef0;
assign v12ad0b3 = hbusreq0 & v12afda2 | !hbusreq0 & v12ad0b2;
assign v1216126 = hgrant1_p & v845542 | !hgrant1_p & v1216125;
assign v121654c = hgrant5_p & v845542 | !hgrant5_p & v121654b;
assign v12164d1 = hmastlock_p & v12164d0 | !hmastlock_p & v845542;
assign v1445fb5 = hlock3 & v1445fb2 | !hlock3 & v1445fb4;
assign v121534e = hmaster0_p & v1215349 | !hmaster0_p & v121534d;
assign v1668ddf = hmaster1_p & v1668dde | !hmaster1_p & v1668dd2;
assign v134d288 = hlock5_p & v134d286 | !hlock5_p & v134d287;
assign v1215394 = hbusreq0_p & v1216aad | !hbusreq0_p & v845542;
assign v15157e9 = hlock5_p & v15157e6 | !hlock5_p & !v15157e8;
assign v14453ba = hlock2 & v14453b6 | !hlock2 & v14453b9;
assign v12ad0ba = hmaster0_p & v845542 | !hmaster0_p & v12ad0b9;
assign d30238 = hbusreq2 & d30230 | !hbusreq2 & d30237;
assign d2fb44 = hbusreq2_p & d2ff04 | !hbusreq2_p & d2fb43;
assign f2f3ad = hmaster0_p & f2f2a8 | !hmaster0_p & f2f2ab;
assign v1445fa2 = hlock0 & v1445fa1 | !hlock0 & v1445fa0;
assign d305d4 = hlock5_p & v845542 | !hlock5_p & v1668c17;
assign v15168f0 = stateA1_p & v845542 | !stateA1_p & !v1553933;
assign d306e8 = hmaster1_p & d306e7 | !hmaster1_p & d306e4;
assign v134cd56 = hbusreq4_p & v134cd55 | !hbusreq4_p & v134d273;
assign v1445e03 = hlock1 & v1445dfc | !hlock1 & v1445e02;
assign v1515724 = hmaster2_p & v1515723 | !hmaster2_p & v1668d36;
assign v12acfeb = hbusreq2_p & v12acfe9 | !hbusreq2_p & v12acfea;
assign v15533a4 = hgrant5_p & v845542 | !hgrant5_p & v15533a3;
assign v1516217 = hready_p & v845542 | !hready_p & v1516216;
assign v121510c = hmaster0_p & v1215057 | !hmaster0_p & v1215463;
assign d30112 = hmaster0_p & d2fe9b | !hmaster0_p & d30111;
assign d30745 = hmaster0_p & d30744 | !hmaster0_p & d3071e;
assign v1215c81 = hbusreq5_p & v1215c7f | !hbusreq5_p & v1215c80;
assign v1445f3f = hmaster1_p & v1445da7 | !hmaster1_p & v1445dc2;
assign v1668ce1 = hmaster2_p & v845542 | !hmaster2_p & !v1668cdf;
assign v1668d74 = hbusreq1 & a653c4 | !hbusreq1 & !v845542;
assign v14459c9 = hlock1 & v14459c2 | !hlock1 & v14459c8;
assign d307b3 = hgrant4_p & d307b0 | !hgrant4_p & d307b2;
assign d302ee = hready_p & d302ed | !hready_p & d302dc;
assign v151560b = hmaster2_p & v1515609 | !hmaster2_p & v845542;
assign a6539b = hbusreq1_p & a65391 | !hbusreq1_p & !a6539a;
assign v1214bf4 = hlock2_p & v1214bf0 | !hlock2_p & v1214bf3;
assign v12157ae = hlock4_p & v12157ac | !hlock4_p & v12157ad;
assign v1216193 = hbusreq5_p & v1216191 | !hbusreq5_p & v1216192;
assign v12150c9 = hmaster2_p & v1215b97 | !hmaster2_p & v12150c7;
assign v14058ab = hlock0_p & v140583f | !hlock0_p & v14058aa;
assign a6538d = hgrant5_p & a65360 | !hgrant5_p & a6538a;
assign v12160b1 = hlock2_p & v12160ae | !hlock2_p & v12160b0;
assign v1446060 = hgrant5_p & v1445fd6 | !hgrant5_p & v144605f;
assign v151570b = hbusreq5 & v1515700 | !hbusreq5 & v151570a;
assign v16a19ac = hgrant5_p & v845568 | !hgrant5_p & v16a19ab;
assign v14458a9 = hbusreq2_p & v14458a0 | !hbusreq2_p & v14458a8;
assign v10d406e = hmaster2_p & v10d406d | !hmaster2_p & !v10d4069;
assign v1553138 = locked_p & v1553137 | !locked_p & v845542;
assign d30272 = hbusreq5_p & d30271 | !hbusreq5_p & !d30270;
assign v121608c = hmaster1_p & v1216071 | !hmaster1_p & v1216082;
assign v16a1be0 = hgrant5_p & v845542 | !hgrant5_p & !v16a1bbf;
assign v12ad5bc = hbusreq1 & v12ad5ba | !hbusreq1 & v12ad5bb;
assign v1445bc9 = hbusreq2_p & v1445bc5 | !hbusreq2_p & v1445bc8;
assign v1215c87 = hgrant1_p & f2f285 | !hgrant1_p & v12160f4;
assign v16a1d5b = hgrant5_p & v845542 | !hgrant5_p & !v16a1d41;
assign d2fcb5 = hmaster0_p & d2fcb3 | !hmaster0_p & d2fcb4;
assign a66283 = hlock4_p & v845570 | !hlock4_p & !v845542;
assign v1445b04 = hmaster1_p & v1445b03 | !hmaster1_p & v14458fd;
assign v144576f = hlock3 & v1445766 | !hlock3 & v144576e;
assign f2f373 = hbusreq1_p & f2f372 | !hbusreq1_p & v845542;
assign v134d20b = hmaster0_p & v134d1e8 | !hmaster0_p & v134d20a;
assign v1215027 = hgrant0_p & v121545e | !hgrant0_p & !v845542;
assign v1445da8 = hbusreq0 & v1445da6 | !hbusreq0 & v1445da7;
assign a65613 = hmaster0_p & a65878 | !hmaster0_p & a6585e;
assign v10d408e = hgrant2_p & v10d408a | !hgrant2_p & v10d408d;
assign v12ad5d6 = hlock4_p & v12ad5d4 | !hlock4_p & v12ad5d5;
assign d80750 = hlock2_p & d8074e | !hlock2_p & d8074f;
assign v16a1ad3 = hbusreq2 & v16a1ad2 | !hbusreq2 & v16a1f9b;
assign v1668e01 = decide_p & v1668d12 | !decide_p & v845542;
assign a658aa = stateA1_p & a658a7 | !stateA1_p & !a658a9;
assign d307ee = hmaster2_p & d307e5 | !hmaster2_p & d307ed;
assign v1215456 = hmaster1_p & v1215455 | !hmaster1_p & v121540f;
assign v134d232 = hmaster0_p & v134d22b | !hmaster0_p & v134d218;
assign a65408 = hbusreq2_p & a653e9 | !hbusreq2_p & a65407;
assign f2f53e = decide_p & f2f53d | !decide_p & f2f23c;
assign v1446288 = hlock2 & v1446275 | !hlock2 & v1446286;
assign v14466a8 = hlock0 & v14466a4 | !hlock0 & v14466a7;
assign v12acfc8 = hbusreq2 & v12acfbb | !hbusreq2 & v12acfc7;
assign v134d379 = hgrant5_p & v134d36a | !hgrant5_p & v134d378;
assign d306ca = hlock1_p & d306c9 | !hlock1_p & v845570;
assign a658a7 = busreq_p & v845542 | !busreq_p & !a658a5;
assign v1446624 = hbusreq0_p & v144639c | !hbusreq0_p & v14465c4;
assign v1215ff8 = hready & v1215ff7 | !hready & v845570;
assign a65650 = hbusreq0 & a65648 | !hbusreq0 & a6564f;
assign a6627b = hbusreq4_p & v84556a | !hbusreq4_p & !v845542;
assign v1445e39 = hbusreq1_p & v1446398 | !hbusreq1_p & v1445e38;
assign v1445ff6 = hlock3 & v1445ff3 | !hlock3 & v1445ff5;
assign v11ac6a3 = hgrant2_p & v84554c | !hgrant2_p & v11ac67c;
assign v12166fb = hbusreq2_p & v12166f1 | !hbusreq2_p & v12166fa;
assign v15168a6 = hmaster1_p & v15168a5 | !hmaster1_p & v845542;
assign v16a1cc8 = hready_p & v16a1c05 | !hready_p & v16a1cc7;
assign v16a1ce1 = hmaster1_p & v16a1cd5 | !hmaster1_p & !v16a1f96;
assign v16a12e6 = hbusreq0_p & v16a2073 | !hbusreq0_p & v845542;
assign v10d40d3 = hmaster0_p & v10d4092 | !hmaster0_p & v10d408c;
assign f2f3c3 = hbusreq5_p & f2f3c0 | !hbusreq5_p & !f2f3c2;
assign v1216551 = hbusreq4 & v1216a61 | !hbusreq4 & v1216550;
assign v12ad320 = hbusreq5_p & v12ae1f3 | !hbusreq5_p & v12ad31f;
assign v121507b = hmaster0_p & v121507a | !hmaster0_p & !v1215053;
assign v1445ef0 = hmaster0_p & v1445eef | !hmaster0_p & v1445ea9;
assign v1216584 = hmaster0_p & v1216a91 | !hmaster0_p & v1216a8f;
assign v12aec0b = hgrant2_p & v845542 | !hgrant2_p & v12aec0a;
assign v16a1ca3 = hbusreq2 & v16a1c9d | !hbusreq2 & v16a1ca2;
assign v1668c2d = hmastlock_p & a658a3 | !hmastlock_p & v845542;
assign v1668d7b = hgrant4_p & v1668d7a | !hgrant4_p & a653cc;
assign v1668d4e = hgrant5_p & v1668d43 | !hgrant5_p & v1668d4d;
assign d2fea7 = hbusreq2_p & d2fea3 | !hbusreq2_p & d2fea6;
assign v144582a = hgrant2_p & v1445829 | !hgrant2_p & v1445825;
assign v1215fe4 = decide_p & v12164cd | !decide_p & v1215fe3;
assign v1445e56 = hbusreq4 & v14465bf | !hbusreq4 & v14465c3;
assign v12152e6 = hmaster0_p & v1215ba3 | !hmaster0_p & v1215b98;
assign a656d1 = decide_p & a656d0 | !decide_p & a662a2;
assign v15533a0 = hgrant0_p & v1553217 | !hgrant0_p & v845542;
assign v134d364 = hmaster1_p & v134d363 | !hmaster1_p & v845542;
assign v15168b7 = decide_p & v15168b6 | !decide_p & v845542;
assign v134cd80 = hmaster0_p & v134cd7f | !hmaster0_p & v134cd6a;
assign v14457df = hmaster1_p & v1445eba | !hmaster1_p & v1445eaa;
assign v1215b90 = hbusreq4 & v1216014 | !hbusreq4 & v845542;
assign v16a2065 = hbusreq5 & v16a205e | !hbusreq5 & v16a2064;
assign v121612b = hgrant5_p & v1216117 | !hgrant5_p & v121612a;
assign v138a464 = hbusreq3 & v138a456 | !hbusreq3 & v138a463;
assign d2fc08 = hlock2_p & d2fc07 | !hlock2_p & v84554a;
assign v11e5945 = hgrant4_p & v845542 | !hgrant4_p & v11e5944;
assign v12af1c1 = hmaster1_p & v12af7f7 | !hmaster1_p & v12af1c0;
assign v1446175 = hmaster1_p & v1446174 | !hmaster1_p & v1446099;
assign v1389de7 = hbusreq5_p & v1389de6 | !hbusreq5_p & !v845542;
assign v15167fb = hlock2_p & v15167fa | !hlock2_p & !v845542;
assign v14453b5 = hgrant2_p & v1445393 | !hgrant2_p & v14453b4;
assign v16a13a7 = hready & v16a1d16 | !hready & v845542;
assign v1445b46 = hmaster1_p & v1445b45 | !hmaster1_p & v144590e;
assign v12ad66a = decide_p & v12ad669 | !decide_p & v845542;
assign v12ad4d2 = hbusreq0 & v12ad4d1 | !hbusreq0 & v845542;
assign a65416 = hgrant5_p & v845558 | !hgrant5_p & !a65378;
assign v1668d0e = hbusreq2_p & v1668d0b | !hbusreq2_p & v1668d06;
assign v1446680 = hmaster0_p & v1446404 | !hmaster0_p & v144667f;
assign v1515803 = hlock2_p & v15157fa | !hlock2_p & v1515802;
assign v12150a6 = hmaster0_p & v121509e | !hmaster0_p & !v12150a5;
assign v16a131d = stateA1_p & v16a2237 | !stateA1_p & v16a131c;
assign v1445532 = hbusreq2 & v1445531 | !hbusreq2 & v1445523;
assign v16a1cf6 = hgrant5_p & v845542 | !hgrant5_p & !v16a1cec;
assign v15530f2 = hbusreq5 & v15530f0 | !hbusreq5 & v15530f1;
assign v1216224 = hmaster0_p & v1216215 | !hmaster0_p & v1216223;
assign v14058c6 = hbusreq1_p & v140583f | !hbusreq1_p & v14058c5;
assign v14460bc = hbusreq2_p & v14460b8 | !hbusreq2_p & v14460bb;
assign v12aead4 = hready_p & v12af22c | !hready_p & v12aead3;
assign v134ce62 = hmaster0_p & v134ce61 | !hmaster0_p & v134ce45;
assign v1215ca0 = hmaster2_p & v1215fec | !hmaster2_p & v1215c7e;
assign v1214ef5 = hgrant5_p & v845542 | !hgrant5_p & v1216562;
assign d30884 = hgrant2_p & d30881 | !hgrant2_p & d30883;
assign v1446668 = hlock2 & v1446651 | !hlock2 & v1446667;
assign v14458d1 = hbusreq5 & v14458cf | !hbusreq5 & v14458d0;
assign v1284c9a = hbusreq1_p & v1284c99 | !hbusreq1_p & v144639e;
assign a65878 = hmaster2_p & a65852 | !hmaster2_p & a65863;
assign d301c7 = hmaster2_p & a65861 | !hmaster2_p & d301c5;
assign f2f2e2 = hbusreq1_p & f2f2e1 | !hbusreq1_p & !v845542;
assign v1445400 = hlock5 & v14453f5 | !hlock5 & v14453fe;
assign d3071e = hmaster2_p & d3071b | !hmaster2_p & d3071d;
assign v134d1f9 = hmaster2_p & v845542 | !hmaster2_p & v134d1f8;
assign v16a1b69 = hbusreq2 & v16a1b67 | !hbusreq2 & v16a1b68;
assign v1445a76 = hmaster2_p & v1445a53 | !hmaster2_p & v14459cf;
assign v10d3fe7 = hlock0_p & v10d3fdb | !hlock0_p & v10d3fe6;
assign v121602d = hlock1_p & v16a1c95 | !hlock1_p & !v845542;
assign v14461e3 = hgrant2_p & v14461b0 | !hgrant2_p & v14461e2;
assign v138953b = hmaster0_p & v138953a | !hmaster0_p & !v845542;
assign v1215097 = hbusreq1_p & v1215035 | !hbusreq1_p & v1215096;
assign f2f34e = hgrant5_p & f2f293 | !hgrant5_p & !f2f34d;
assign v1215076 = hbusreq3 & v121506a | !hbusreq3 & v1215075;
assign a81304 = stateG3_1_p & v845542 | !stateG3_1_p & !v84556c;
assign d306de = hbusreq0_p & v845542 | !hbusreq0_p & d306d4;
assign v1216518 = hbusreq5 & v12164e6 | !hbusreq5 & v12164e7;
assign v16a1bca = hbusreq1_p & v16a1bc9 | !hbusreq1_p & v16a2089;
assign v14465cc = hlock1 & v14465c9 | !hlock1 & v14465cb;
assign v12ad57e = hbusreq2 & v12ad576 | !hbusreq2 & v12ad57d;
assign v134cea8 = hlock5 & v134ce97 | !hlock5 & v134cea7;
assign d3094f = hmastlock_p & d3094e | !hmastlock_p & v845542;
assign v138a34b = hbusreq5_p & v138a34a | !hbusreq5_p & !v845542;
assign v1215350 = hmaster2_p & v121534b | !hmaster2_p & v121534f;
assign a656c9 = hmaster2_p & a66299 | !hmaster2_p & a662ac;
assign v151580a = hready_p & v1515808 | !hready_p & !v1515809;
assign v1214c53 = hgrant5_p & v121534c | !hgrant5_p & v1214c52;
assign v1215786 = hmaster1_p & v1215785 | !hmaster1_p & v845542;
assign a654c3 = hbusreq2 & a654bc | !hbusreq2 & a654c0;
assign a653c3 = hbusreq0_p & v10d3fd8 | !hbusreq0_p & !a65861;
assign v15157e7 = hmaster2_p & v151563e | !hmaster2_p & v845542;
assign d2f9b7 = hbusreq4_p & d2f9b6 | !hbusreq4_p & v845542;
assign d2fec8 = hmaster2_p & d2feb2 | !hmaster2_p & v84555a;
assign v1215085 = hmaster1_p & v121506b | !hmaster1_p & !v121507b;
assign v10d400a = hmaster2_p & v10d3fd4 | !hmaster2_p & v10d3fd9;
assign v1215c39 = hmaster1_p & v1215c38 | !hmaster1_p & !v1215beb;
assign d30256 = hgrant5_p & v845542 | !hgrant5_p & d30227;
assign v1214d61 = hbusreq2_p & v1214c14 | !hbusreq2_p & v1214d60;
assign v121622a = hmaster2_p & v1216207 | !hmaster2_p & v1216212;
assign v12ad60c = hmaster2_p & v12ad506 | !hmaster2_p & v845542;
assign v121531f = hmaster1_p & v121531e | !hmaster1_p & v121546f;
assign v12164c4 = hlock2_p & v12164c2 | !hlock2_p & v12164c3;
assign v10d42d2 = hgrant2_p & v10d40b1 | !hgrant2_p & v10d42d1;
assign v1445867 = hbusreq5 & v1445842 | !hbusreq5 & v1445866;
assign v1214c6f = hmaster2_p & v1214c6e | !hmaster2_p & v845542;
assign v138a3d4 = hmaster2_p & v845542 | !hmaster2_p & v15157ae;
assign v1515615 = hmaster2_p & v1515612 | !hmaster2_p & v1515614;
assign v1446720 = hbusreq3 & v144671f | !hbusreq3 & v144671d;
assign v1446685 = hbusreq2 & v1446668 | !hbusreq2 & v1446684;
assign f2f3d3 = hgrant5_p & v84554c | !hgrant5_p & f2f39f;
assign d30850 = hbusreq5_p & d30708 | !hbusreq5_p & d3084f;
assign d301d7 = hgrant1_p & d301d0 | !hgrant1_p & d3079c;
assign v12ad016 = hbusreq0 & v12ad015 | !hbusreq0 & v12afa0a;
assign v10d42b0 = hgrant0_p & v10d3fd4 | !hgrant0_p & v10d42af;
assign d301f0 = hlock5_p & d301ee | !hlock5_p & d301ef;
assign d30148 = hbusreq5_p & d30147 | !hbusreq5_p & d30146;
assign v16a206f = hgrant1_p & v84554d | !hgrant1_p & v16a206e;
assign d308eb = hbusreq2_p & d308de | !hbusreq2_p & d308ea;
assign v16a1bd6 = hgrant1_p & v84554d | !hgrant1_p & v16a1bd5;
assign v134d3be = decide_p & v845542 | !decide_p & v134d1e0;
assign d306d8 = hmaster2_p & d306d7 | !hmaster2_p & v845542;
assign bf1fa9 = hready_p & bf1fa8 | !hready_p & bf1f88;
assign v1553385 = hgrant5_p & v845542 | !hgrant5_p & v1553384;
assign v1445a54 = hmaster2_p & v144599d | !hmaster2_p & v1445a53;
assign v155321e = hmaster1_p & v155321d | !hmaster1_p & v845542;
assign v1215cb5 = hmaster2_p & v1215cb4 | !hmaster2_p & v1215caf;
assign d30223 = hmaster2_p & v845580 | !hmaster2_p & !a65861;
assign v1214ec5 = hbusreq2 & v1214ec4 | !hbusreq2 & v12164e7;
assign v16a1bd3 = hgrant4_p & v845559 | !hgrant4_p & v16a1bd2;
assign v12acfbb = hbusreq2_p & v12ad66c | !hbusreq2_p & v12acfba;
assign v1405842 = hmaster0_p & v1405840 | !hmaster0_p & v1405841;
assign d306cf = hlock1_p & v845542 | !hlock1_p & v845570;
assign v1515741 = locked_p & a658c3 | !locked_p & v10d3fdf;
assign v12aecdc = hgrant3_p & v12aeb85 | !hgrant3_p & v12aecdb;
assign a65909 = hmaster1_p & a658ee | !hmaster1_p & a658e5;
assign v14459b8 = hbusreq1 & v14459b2 | !hbusreq1 & v14459b7;
assign v16a1a29 = hmaster1_p & v16a19e4 | !hmaster1_p & !v16a1f96;
assign d8078c = hgrant1_p & d8078b | !hgrant1_p & !v845542;
assign v1214e66 = hbusreq2 & v1214e65 | !hbusreq2 & v845542;
assign v14461bc = hlock2 & v14461b3 | !hlock2 & v14461bb;
assign v1446659 = hmaster1_p & v1446658 | !hmaster1_p & v1446436;
assign v1405854 = locked_p & v1405853 | !locked_p & v14463b1;
assign v12147e5 = hmaster0_p & v1215d41 | !hmaster0_p & v1215d2f;
assign v12aed9f = hready_p & v12af7e2 | !hready_p & v12aed9e;
assign v144609b = hgrant2_p & v1446098 | !hgrant2_p & v144609a;
assign d30668 = hgrant1_p & f2f227 | !hgrant1_p & d30667;
assign v1215c14 = hbusreq1_p & v1215ff9 | !hbusreq1_p & v1215c13;
assign v14453e2 = hmaster1_p & v14453e1 | !hmaster1_p & v1445bb1;
assign v14460fd = hlock2 & v14460f2 | !hlock2 & v14460fb;
assign f2f343 = hmaster0_p & f2f293 | !hmaster0_p & f2f296;
assign v1446217 = hbusreq0 & v14463b8 | !hbusreq0 & v14463be;
assign d301cf = hlock1_p & d306c9 | !hlock1_p & !d301ce;
assign v1215cea = hbusreq5_p & v1215ce9 | !hbusreq5_p & v1215c9a;
assign v1669598 = hmaster0_p & v1668c1d | !hmaster0_p & v845570;
assign v15534ce = hbusreq1 & v155339b | !hbusreq1 & v155339c;
assign v14462a1 = hlock5 & v144628b | !hlock5 & v14462a0;
assign d30789 = stateA1_p & v845542 | !stateA1_p & !d30788;
assign v1668c17 = hmaster2_p & v845570 | !hmaster2_p & a66295;
assign v12ad574 = hmaster0_p & v12ad531 | !hmaster0_p & v12ad528;
assign v12ad329 = hmaster0_p & v12af9c3 | !hmaster0_p & v12ad328;
assign v1445df0 = hmaster2_p & v1446403 | !hmaster2_p & v1445def;
assign v134cd8b = hlock5 & v134d3b5 | !hlock5 & v134cd7a;
assign v144588b = stateG10_5_p & v144588a | !stateG10_5_p & !v1445889;
assign v16a1dbd = hbusreq3_p & v16a1da1 | !hbusreq3_p & v16a1dbc;
assign d3073a = hbusreq2 & d30732 | !hbusreq2 & d30739;
assign a6545c = hmaster1_p & a6545b | !hmaster1_p & a653f3;
assign v1214cfb = hgrant5_p & v1214cf8 | !hgrant5_p & !v1214cfa;
assign v12150fa = hmaster1_p & v12150f9 | !hmaster1_p & v12150ef;
assign d306c2 = hbusreq2_p & d3067e | !hbusreq2_p & !d306c1;
assign v1405873 = hmaster1_p & v1405872 | !hmaster1_p & v140586f;
assign v1214d44 = hbusreq5_p & v12153a0 | !hbusreq5_p & v1214d43;
assign v1216599 = hbusreq5_p & v1216598 | !hbusreq5_p & v845542;
assign v9a051b = hburst1_p & v906a5a | !hburst1_p & v893df7;
assign d3089e = hbusreq1_p & d307cb | !hbusreq1_p & d306ae;
assign v10d40db = decide_p & v10d40a8 | !decide_p & v10d40da;
assign v12150b0 = hbusreq3 & v1215084 | !hbusreq3 & v12150af;
assign v16a1bc2 = hgrant4_p & v845559 | !hgrant4_p & !v16a1bc1;
assign f2eda3 = hbusreq3_p & f2eda2 | !hbusreq3_p & f2ed9e;
assign d3025d = hgrant2_p & v845542 | !hgrant2_p & d30259;
assign v14463f1 = hlock1 & v144639c | !hlock1 & v14463d8;
assign v1668d87 = hgrant5_p & v1668d1d | !hgrant5_p & v1668d86;
assign v1445b78 = hbusreq0 & v1445b77 | !hbusreq0 & v14462f3;
assign d2fe8c = hmaster0_p & d2fe88 | !hmaster0_p & d2fe8b;
assign v155313d = decide_p & v155313c | !decide_p & v155313b;
assign f2f41f = hmaster2_p & f2f41d | !hmaster2_p & f2f41e;
assign v1216075 = hlock2_p & v1216072 | !hlock2_p & v1216074;
assign v1389ffe = hmaster0_p & v1389ffd | !hmaster0_p & v1389de1;
assign v1405b5c = hmaster1_p & v1405b5b | !hmaster1_p & !v1405ac8;
assign v144600d = hbusreq1_p & v144646e | !hbusreq1_p & v1446476;
assign d3011a = hgrant5_p & d2fe8e | !hgrant5_p & d30119;
assign v14465e6 = hlock0 & v14465e5 | !hlock0 & v14465de;
assign v1446697 = hbusreq4 & v1446696 | !hbusreq4 & v14465c3;
assign v121503a = hgrant1_p & v1215034 | !hgrant1_p & v1215039;
assign v1216796 = decide_p & v1216a82 | !decide_p & v1216795;
assign d2fbf3 = hlock4_p & d2fb4e | !hlock4_p & v84554a;
assign v121578d = hgrant5_p & v845542 | !hgrant5_p & v121572c;
assign v12162d7 = hmaster0_p & v1216262 | !hmaster0_p & v121625e;
assign d302e6 = hgrant2_p & v845542 | !hgrant2_p & d302e5;
assign d305f4 = hlock1_p & d305f3 | !hlock1_p & !v845542;
assign d3078a = hburst1 & d30789 | !hburst1 & v845542;
assign v144605b = hbusreq1 & v1446430 | !hbusreq1 & v1446424;
assign v15530eb = hbusreq3 & v15530e9 | !hbusreq3 & v15530ea;
assign v134d457 = hlock3 & v134d3b5 | !hlock3 & v134d456;
assign v16a2077 = hmaster2_p & v16a2076 | !hmaster2_p & v16a206f;
assign v16a1f9a = hmaster1_p & v845564 | !hmaster1_p & v16a1f96;
assign v144550d = hbusreq2_p & v144550c | !hbusreq2_p & v1445bdb;
assign v138936f = hbusreq0 & v138936e | !hbusreq0 & !v138a38f;
assign v15534fe = hmaster0_p & v15534fd | !hmaster0_p & v15534da;
assign v12ad5db = hgrant1_p & v12ad5d2 | !hgrant1_p & v12ad5da;
assign v155321d = hmaster0_p & v845542 | !hmaster0_p & v1553139;
assign v16a137c = hgrant2_p & v16a1f9b | !hgrant2_p & v16a137b;
assign v1553416 = hlock0 & v1553415 | !hlock0 & v1553414;
assign d30737 = hmaster1_p & d30736 | !hmaster1_p & d3072c;
assign v12af226 = hbusreq5_p & v12af5ac | !hbusreq5_p & v12af225;
assign v134d3b7 = hbusreq2 & v134d3b2 | !hbusreq2 & v134d3b6;
assign v1553506 = hlock3 & v155341e | !hlock3 & v1553505;
assign v134d466 = hbusreq5 & v134d464 | !hbusreq5 & v134d465;
assign a65379 = hgrant5_p & a65852 | !hgrant5_p & a65378;
assign d302f1 = decide_p & d302d6 | !decide_p & v845570;
assign v1446618 = hbusreq0 & v1446612 | !hbusreq0 & v1446617;
assign v12ad5c6 = hgrant5_p & v12ad5b6 | !hgrant5_p & v12ad5c5;
assign v1214eff = hbusreq2 & v1214efe | !hbusreq2 & v845542;
assign v1668cb5 = hbusreq3 & v1668caf | !hbusreq3 & a7c7c1;
assign v1215caa = hmaster2_p & v1215c87 | !hmaster2_p & v1215ca5;
assign v16a1e29 = hmaster1_p & v16a1e28 | !hmaster1_p & !v16a2672;
assign v12153b4 = hbusreq4_p & v1215bb0 | !hbusreq4_p & v845542;
assign d3070b = hbusreq2_p & d30707 | !hbusreq2_p & d3070a;
assign v134d503 = hgrant4_p & v845542 | !hgrant4_p & v134d502;
assign v1216704 = hmaster1_p & v1216703 | !hmaster1_p & v12166ef;
assign v144624f = hlock0 & v144624e | !hlock0 & v144624d;
assign v1214cf3 = hgrant4_p & v1214c30 | !hgrant4_p & v845572;
assign bf1f63 = hgrant5_p & bf1f62 | !hgrant5_p & bf1f60;
assign v1668ce6 = hmaster0_p & v1668ce2 | !hmaster0_p & v1668ce5;
assign v1515855 = jx2_p & v1515854 | !jx2_p & v151621b;
assign v1445e4a = hmaster0_p & v1445e3f | !hmaster0_p & v1445e49;
assign v12162b3 = hmaster1_p & v12162b2 | !hmaster1_p & v1216041;
assign v144622d = hgrant5_p & v144622a | !hgrant5_p & !v144622c;
assign v1214e82 = hbusreq2_p & v1214e81 | !hbusreq2_p & v845542;
assign v16a16b0 = hbusreq5 & v16a16a4 | !hbusreq5 & v16a16af;
assign d2f983 = hmaster0_p & d2f980 | !hmaster0_p & d2f982;
assign v1389430 = hbusreq2_p & v1389f87 | !hbusreq2_p & v138a06a;
assign v14461c3 = hmaster1_p & v1446184 | !hmaster1_p & v14460b6;
assign v1445f36 = hmaster1_p & v1445f35 | !hmaster1_p & v1445da4;
assign v1216063 = hbusreq2_p & v1216062 | !hbusreq2_p & v1216061;
assign v140592e = hmaster2_p & v140592d | !hmaster2_p & v1405844;
assign v144550a = hmaster1_p & v14454e8 | !hmaster1_p & v144627e;
assign v1445d88 = hbusreq1 & v1445d80 | !hbusreq1 & v1445d87;
assign d2fb78 = hbusreq4_p & d2fb77 | !hbusreq4_p & v84554a;
assign v16a1a85 = hbusreq0 & v16a1a84 | !hbusreq0 & v16a1961;
assign v1216a68 = hmaster2_p & v845542 | !hmaster2_p & v1216a67;
assign v16a1e76 = hmaster1_p & v16a1e63 | !hmaster1_p & !v16a1f96;
assign f2f398 = hmaster2_p & f2f350 | !hmaster2_p & v845542;
assign v1515822 = hlock2_p & v1515821 | !hlock2_p & !v15156f6;
assign v1445799 = hbusreq2 & v1445797 | !hbusreq2 & v1445798;
assign d2fe9f = hmaster2_p & d2fe9c | !hmaster2_p & d2fe9d;
assign v134d3b1 = hbusreq2_p & v134d39c | !hbusreq2_p & v134d3b0;
assign v1445f76 = hmaster1_p & v1446663 | !hmaster1_p & v14466a9;
assign v14466e9 = hlock2 & v14466d3 | !hlock2 & v14466e7;
assign v144623a = hmaster0_p & v144639c | !hmaster0_p & v1446239;
assign v10d42c6 = hbusreq4_p & v10d4269 | !hbusreq4_p & v10d42c5;
assign v1445ed9 = hmaster1_p & v1445ed8 | !hmaster1_p & v1445ed3;
assign d305ec = hlock5_p & v845542 | !hlock5_p & !d305eb;
assign v15156b2 = hmaster1_p & v151567f | !hmaster1_p & !v15156b1;
assign v1445a33 = hmaster1_p & v14459a3 | !hmaster1_p & v1445a32;
assign v1215357 = hmaster0_p & v1215353 | !hmaster0_p & v1215356;
assign d300b8 = hbusreq1_p & d300b7 | !hbusreq1_p & !d300b6;
assign v1216085 = hlock2_p & v1216083 | !hlock2_p & v1216084;
assign v1214ebc = hbusreq2_p & v1214ebb | !hbusreq2_p & v845542;
assign v151699a = hmaster1_p & v1516999 | !hmaster1_p & v845542;
assign v1445a81 = hlock0 & v1445a7a | !hlock0 & v1445a80;
assign v1214c0c = hmaster1_p & v1214c0b | !hmaster1_p & v12153a9;
assign v1445f35 = hmaster0_p & v1445da9 | !hmaster0_p & v1445db8;
assign v16a1cfe = hbusreq2 & v16a1cfb | !hbusreq2 & !v16a1cfd;
assign d2fb12 = hgrant2_p & d2fad6 | !hgrant2_p & !d2fb11;
assign d3080a = hbusreq1_p & d30809 | !hbusreq1_p & v845542;
assign v1214d0a = hmaster1_p & v1214d09 | !hmaster1_p & v1214c39;
assign f2f287 = hmaster2_p & f2f282 | !hmaster2_p & f2f286;
assign v12ad5ca = hbusreq1_p & v12ad5c8 | !hbusreq1_p & !v12ad5c9;
assign d2f971 = hbusreq4_p & d2fe9c | !hbusreq4_p & !v845542;
assign v1515826 = hmaster1_p & v151581a | !hmaster1_p & !v15156da;
assign v1668caf = hbusreq2 & v1668ca7 | !hbusreq2 & v1668cae;
assign v1552f78 = hbusreq3 & v1552f76 | !hbusreq3 & v1552f77;
assign v121623d = hmaster1_p & v121623c | !hmaster1_p & v1216224;
assign d30695 = hmaster0_p & d3068d | !hmaster0_p & d30694;
assign v144670d = hbusreq2_p & v1446704 | !hbusreq2_p & v144670c;
assign v1284cdc = hgrant1_p & v140584b | !hgrant1_p & v1284cdb;
assign v1216057 = hbusreq1 & v1216aeb | !hbusreq1 & v845542;
assign v1445f17 = hbusreq2_p & v1445f0b | !hbusreq2_p & v1445f16;
assign d30622 = hmaster0_p & d3061b | !hmaster0_p & d30613;
assign v121601f = hready & v1215ff6 | !hready & !v845542;
assign v1668c27 = decide_p & v1668c26 | !decide_p & v845542;
assign v10d4007 = hmaster0_p & v10d3ff1 | !hmaster0_p & v10d3ffd;
assign v12ad5b1 = hmaster2_p & v12ad5a8 | !hmaster2_p & v12ad5b0;
assign v134d513 = hmaster0_p & v134d4f8 | !hmaster0_p & v134d512;
assign d2fc53 = hbusreq4_p & d2fbd3 | !hbusreq4_p & d2fc52;
assign v12153de = hmaster2_p & v1215b97 | !hmaster2_p & v12153dc;
assign v1446695 = hlock0 & v1446694 | !hlock0 & v1446693;
assign v1446434 = hbusreq5_p & v1446433 | !hbusreq5_p & v144642a;
assign a6548d = hmaster1_p & a6548c | !hmaster1_p & a65476;
assign v12ad622 = hgrant2_p & v12ad5f5 | !hgrant2_p & v12ad618;
assign v16a1a2a = hbusreq2_p & v16a188c | !hbusreq2_p & v16a1a29;
assign v1552f6d = hmaster2_p & v845542 | !hmaster2_p & v1552f6c;
assign a65671 = hgrant5_p & v949cd9 | !hgrant5_p & a65646;
assign a1db63 = hmaster0_p & v845558 | !hmaster0_p & !v949cd9;
assign v12afdb2 = hbusreq5_p & v12afdb0 | !hbusreq5_p & v12afdb1;
assign d2fce8 = hmaster2_p & v16693aa | !hmaster2_p & d2fce7;
assign f2f43c = hgrant2_p & f2f41c | !hgrant2_p & f2f43b;
assign v16a140c = hbusreq2 & v16a140b | !hbusreq2 & v16a2059;
assign v121653e = hbusreq1 & v1216a61 | !hbusreq1 & v1216a73;
assign f2f38d = hgrant1_p & v845570 | !hgrant1_p & !f2f38c;
assign d2fb19 = hmaster1_p & d2fb18 | !hmaster1_p & d3014e;
assign v1214cc8 = hbusreq1_p & v1215379 | !hbusreq1_p & !v1214cc7;
assign v1215cc5 = hgrant5_p & v845542 | !hgrant5_p & !v1215cc3;
assign d30191 = hbusreq2_p & d30190 | !hbusreq2_p & d30188;
assign v1445f29 = hmaster1_p & v1445da9 | !hmaster1_p & v1445da4;
assign v1445e23 = hbusreq3 & v1445e21 | !hbusreq3 & v1445e22;
assign v1668d3a = hbusreq5_p & v1668d38 | !hbusreq5_p & v1668d39;
assign d2fc80 = hgrant3_p & d2fc48 | !hgrant3_p & d2fc7f;
assign v1553504 = hlock2 & v155341e | !hlock2 & v1553500;
assign f2f237 = hbusreq5_p & f2f232 | !hbusreq5_p & f2f236;
assign v16a1e2d = hmaster1_p & v16a1e2c | !hmaster1_p & !v16a2672;
assign d30847 = hgrant3_p & d3077c | !hgrant3_p & d30846;
assign d30122 = hbusreq2_p & d30110 | !hbusreq2_p & !d30121;
assign v1446071 = hbusreq0 & v144606c | !hbusreq0 & v1446070;
assign v10d4000 = hbusreq2_p & v10d3ffc | !hbusreq2_p & v10d3fff;
assign v16a1e98 = hmaster2_p & v16a1e97 | !hmaster2_p & v16a208a;
assign v1446669 = hmaster1_p & v14465aa | !hmaster1_p & v144644d;
assign v144646d = stateG2_p & v845542 | !stateG2_p & v1446468;
assign v1445ae6 = hmaster1_p & v1445ae5 | !hmaster1_p & v14458fd;
assign v12ad53b = hmaster0_p & v12ad52d | !hmaster0_p & v12ad517;
assign v1214cbe = hgrant1_p & v121537c | !hgrant1_p & v1214cbd;
assign v1214bbc = hbusreq2 & v12153af | !hbusreq2 & v1214bbb;
assign v14460b7 = hmaster1_p & v144603f | !hmaster1_p & v14460b6;
assign v14465d6 = hgrant0_p & v1446406 | !hgrant0_p & v144639e;
assign v1446086 = hbusreq1 & v14465c1 | !hbusreq1 & v14465c5;
assign v144591f = hmaster1_p & v144590a | !hmaster1_p & v144591b;
assign v1445aac = hbusreq5 & v1445a95 | !hbusreq5 & v1445aab;
assign v1445e88 = hlock0_p & v1446403 | !hlock0_p & v1445e87;
assign v144603a = hgrant0_p & v14465ae | !hgrant0_p & v144639c;
assign f2e506 = jx0_p & f2eda5 | !jx0_p & f2e505;
assign v1284d5a = decide_p & v1284d52 | !decide_p & v1284d59;
assign v12153f4 = hmaster0_p & v12153d4 | !hmaster0_p & v12153f3;
assign v14463d1 = hbusreq2_p & v14463ce | !hbusreq2_p & v14463d0;
assign v1445b5f = hmaster0_p & v1445b5e | !hmaster0_p & v14462fe;
assign v15167bd = hmaster2_p & v845542 | !hmaster2_p & d305f2;
assign v16a194a = hbusreq4_p & v16a1949 | !hbusreq4_p & v845542;
assign v10d427e = stateA1_p & v84557e | !stateA1_p & v10d427d;
assign v845542 = 1;
assign v1552f88 = hlock5 & v1552f78 | !hlock5 & v1552f87;
assign v12162cf = hgrant2_p & v12162be | !hgrant2_p & v12162ce;
assign d2fd37 = hready_p & d2fd30 | !hready_p & d2fd19;
assign v1668d55 = hmaster2_p & v1668d54 | !hmaster2_p & v1668d4c;
assign v1214ec4 = hbusreq2_p & v1214ec3 | !hbusreq2_p & v12164e7;
assign v121507e = hmaster1_p & v121505c | !hmaster1_p & !v121507b;
assign v1445fc5 = hbusreq2 & v1445fc3 | !hbusreq2 & v1445fc4;
assign v1668da8 = hmaster0_p & v1668da6 | !hmaster0_p & v1668da7;
assign d2fe87 = hmaster2_p & d2fe84 | !hmaster2_p & d2fe85;
assign v16a19ca = hbusreq2 & v16a19c7 | !hbusreq2 & v16a19c9;
assign v1515667 = hbusreq1_p & a658e0 | !hbusreq1_p & a65472;
assign v12ad0b2 = hmaster2_p & v845542 | !hmaster2_p & v12ad0b1;
assign v1445bd2 = stateG10_5_p & v1446041 | !stateG10_5_p & v14465dc;
assign v10d42df = hgrant3_p & v10d40af | !hgrant3_p & !v10d42de;
assign v151697b = hlock2_p & v151697a | !hlock2_p & v845542;
assign v1405ac4 = hbusreq4_p & v845542 | !hbusreq4_p & v1405abf;
assign a65aff = hmaster1_p & v845542 | !hmaster1_p & a65afe;
assign v1445b3e = hmaster0_p & v1445902 | !hmaster0_p & v1445a4f;
assign v1214d4f = hmaster2_p & v1215392 | !hmaster2_p & v1214d4e;
assign d307ca = hbusreq1 & d307c9 | !hbusreq1 & v845542;
assign v1668d54 = hgrant1_p & v1668d53 | !hgrant1_p & v1668d4a;
assign v14058ed = hmaster2_p & v140583f | !hmaster2_p & !v1446403;
assign d307f9 = hmaster1_p & d307f8 | !hmaster1_p & !d30706;
assign v1214bd3 = hbusreq2_p & v1214bd2 | !hbusreq2_p & v1214bd1;
assign d3026a = hgrant5_p & v1668da6 | !hgrant5_p & d30269;
assign v1215bf5 = hbusreq5_p & v1215bf3 | !hbusreq5_p & !v1215bf4;
assign v16a144a = jx1_p & v16a139f | !jx1_p & v16a1449;
assign v12ad5f7 = hmaster2_p & v845542 | !hmaster2_p & v12ad5bb;
assign d307f6 = hgrant2_p & d3077f | !hgrant2_p & d307f5;
assign v134d228 = hlock5_p & v134d215 | !hlock5_p & v134d21f;
assign d2fef2 = hmaster1_p & d2fedc | !hmaster1_p & d2fee5;
assign v12afe5c = hgrant1_p & v845542 | !hgrant1_p & v12afe5b;
assign v1215da9 = hbusreq2 & v1215da2 | !hbusreq2 & v1215da8;
assign v14460f5 = hmaster0_p & v1445fa9 | !hmaster0_p & v144639c;
assign v1445543 = hbusreq5_p & v14465e3 | !hbusreq5_p & v1445542;
assign v1215c1a = hgrant1_p & v1215c0b | !hgrant1_p & v1215c19;
assign d2fef9 = hmaster1_p & d2fef8 | !hmaster1_p & d2fec6;
assign f2e4f3 = hbusreq2 & f2e4f2 | !hbusreq2 & f2ed94;
assign v12add4c = hmaster1_p & v845542 | !hmaster1_p & v12add4b;
assign d30704 = hlock1_p & d30703 | !hlock1_p & !v845542;
assign v1216129 = hbusreq5_p & v121611b | !hbusreq5_p & v1216128;
assign v1445f0c = hmaster1_p & v1445ebb | !hmaster1_p & v1445f09;
assign v1215bda = hmaster2_p & v1215fe8 | !hmaster2_p & v845542;
assign v12ad59e = hbusreq4_p & v12ad59c | !hbusreq4_p & v12ad59d;
assign f2f384 = hbusreq1_p & f2f383 | !hbusreq1_p & v845542;
assign v1214d4a = hbusreq0 & v1214d49 | !hbusreq0 & v845542;
assign v16a1cce = hbusreq2_p & v16a1afc | !hbusreq2_p & v16a1ccd;
assign v1214db4 = hbusreq2_p & v1214db3 | !hbusreq2_p & v1214daf;
assign v12ad03d = jx2_p & v12ad4c9 | !jx2_p & v12ad03c;
assign v1445761 = hlock2 & v1445f40 | !hlock2 & v144575f;
assign v12153e9 = hbusreq4_p & v12153e8 | !hbusreq4_p & v845542;
assign d306a2 = hready_p & d30687 | !hready_p & d306a1;
assign d2f96b = hbusreq4_p & d2fe9a | !hbusreq4_p & v845542;
assign v134ce8c = hgrant1_p & v134ce8b | !hgrant1_p & v134d1e8;
assign v134d1ef = hlock1 & v134d1e8 | !hlock1 & v134d1ee;
assign d30226 = hbusreq5_p & d30225 | !hbusreq5_p & !d30224;
assign v11e5951 = hbusreq5_p & v11e5950 | !hbusreq5_p & v11e594f;
assign v15168b0 = hbusreq1_p & v15168af | !hbusreq1_p & !v845542;
assign f2f33e = hbusreq2 & f2f33a | !hbusreq2 & f2f33d;
assign v14459d6 = hlock0_p & v845542 | !hlock0_p & v14459d5;
assign v16a1390 = hbusreq2_p & v16a12c0 | !hbusreq2_p & v16a138f;
assign v1445fa1 = hbusreq0 & v1445fa0 | !hbusreq0 & v1445f85;
assign v1215d8f = hbusreq2 & v1215d84 | !hbusreq2 & v1215d8e;
assign v134d3aa = hmaster2_p & v845542 | !hmaster2_p & v134d3a9;
assign v1215382 = hmaster2_p & d2fbe5 | !hmaster2_p & v1215380;
assign v1445e67 = hbusreq4_p & v14465cd | !hbusreq4_p & v14465d6;
assign v14457ec = hlock2 & v14457e1 | !hlock2 & v14457eb;
assign d307a1 = hmaster2_p & d307a0 | !hmaster2_p & d30796;
assign v16a1424 = hbusreq2_p & v16a13cf | !hbusreq2_p & v16a1aca;
assign v155304c = hbusreq0_p & v155338c | !hbusreq0_p & v1553217;
assign v1214ddf = hmaster0_p & v1216a8e | !hmaster0_p & v1668da6;
assign v12ad67f = hbusreq1_p & v12ad51b | !hbusreq1_p & !v12ad67e;
assign v16a13e5 = hmaster0_p & v16a13e1 | !hmaster0_p & v16a13e4;
assign a65436 = hgrant5_p & v949cd9 | !hgrant5_p & a653e2;
assign f2f21f = hbusreq1_p & f2f21e | !hbusreq1_p & !v845542;
assign d2fed6 = hmaster0_p & d2fed5 | !hmaster0_p & d2feb5;
assign v1215060 = hbusreq4_p & v121504a | !hbusreq4_p & !v845542;
assign v1216b0f = hmaster0_p & v1216b03 | !hmaster0_p & v1216afb;
assign v1445faa = hmaster0_p & v144639c | !hmaster0_p & v1445fa9;
assign v1445b0a = hlock2 & v1445af2 | !hlock2 & v1445b08;
assign v1216526 = stateA1_p & v845542 | !stateA1_p & !v134d1db;
assign v12ad58b = hmaster1_p & v12ad577 | !hmaster1_p & v12ad54f;
assign v1216281 = hmaster1_p & v1216280 | !hmaster1_p & v121600c;
assign v16a2240 = hbusreq5_p & v16a223f | !hbusreq5_p & v845568;
assign v14460af = hmaster2_p & v1446087 | !hmaster2_p & v1446412;
assign v1215cd2 = hgrant5_p & v845542 | !hgrant5_p & !v1215cd0;
assign d3079d = hbusreq1 & d3079c | !hbusreq1 & v845542;
assign a65643 = hgrant4_p & a662a9 | !hgrant4_p & !a653cd;
assign f2f443 = hmaster1_p & f2f442 | !hmaster1_p & f2f3cf;
assign v1214c09 = hlock2_p & v1214c06 | !hlock2_p & v1214c08;
assign v134d3e9 = hbusreq3_p & v134d3bd | !hbusreq3_p & v134d3e8;
assign v1445e25 = hbusreq5_p & v1445df0 | !hbusreq5_p & v1445e24;
assign v12ad609 = hmaster2_p & v12ad4e6 | !hmaster2_p & !v12ad4e4;
assign v138937e = hmaster0_p & v138937d | !hmaster0_p & v1389de1;
assign v1215cf5 = hgrant5_p & v845542 | !hgrant5_p & v1215cbd;
assign v1215461 = hbusreq4_p & v1215460 | !hbusreq4_p & v845542;
assign v16a1e23 = hgrant5_p & v16a2234 | !hgrant5_p & v16a1e22;
assign v134d53f = hready_p & v134d53d | !hready_p & v134d53e;
assign v1446330 = hmaster2_p & v14465ae | !hmaster2_p & v1446677;
assign v1515785 = hbusreq0 & v1515778 | !hbusreq0 & v1515784;
assign v1445fd6 = hmaster2_p & v1445fd4 | !hmaster2_p & v1445fd5;
assign v16a1bda = hbusreq0 & v16a1bd8 | !hbusreq0 & v16a1bd9;
assign v14058e0 = hmaster0_p & v14058c4 | !hmaster0_p & v14058df;
assign f2f36f = hbusreq5_p & f2f360 | !hbusreq5_p & !f2f36e;
assign v1405ad8 = hgrant5_p & v1405a8a | !hgrant5_p & v1405ad7;
assign v16695aa = jx2_p & v1669594 | !jx2_p & v16695a9;
assign v1215783 = hmaster0_p & v845542 | !hmaster0_p & v1215b93;
assign v134d241 = hbusreq5 & v134d239 | !hbusreq5 & v134d240;
assign v16693ab = hbusreq4_p & v16693aa | !hbusreq4_p & !v845542;
assign v15534d3 = hbusreq0 & v15534d2 | !hbusreq0 & v15533a7;
assign d30155 = hgrant5_p & d2fe80 | !hgrant5_p & d30119;
assign v14463e9 = hmaster2_p & v14463e4 | !hmaster2_p & v14463e8;
assign a65884 = stateG3_2_p & v88d3e4 | !stateG3_2_p & a65883;
assign v14453fc = hbusreq2 & v14453fa | !hbusreq2 & v14453fb;
assign v1445999 = hgrant4_p & v14458d2 | !hgrant4_p & v1445998;
assign d306fa = hmaster1_p & d306f8 | !hmaster1_p & d306f9;
assign v1389f94 = hmaster1_p & v845542 | !hmaster1_p & v1389f93;
assign v1445438 = hlock3 & v144541f | !hlock3 & v1445437;
assign d30832 = hgrant2_p & d3077f | !hgrant2_p & d30831;
assign v121620e = hbusreq1_p & v121620d | !hbusreq1_p & !v845542;
assign v134d42a = hbusreq0 & v134d429 | !hbusreq0 & v134d38b;
assign a66299 = hgrant1_p & v845542 | !hgrant1_p & !a66298;
assign d2fbb6 = hmaster1_p & d2fbb5 | !hmaster1_p & d2fb7b;
assign d3061c = hmaster0_p & d3061b | !hmaster0_p & d305ed;
assign v1215069 = hbusreq2_p & v1215068 | !hbusreq2_p & v121505e;
assign v12ad57f = hbusreq3 & v12ad571 | !hbusreq3 & v12ad57e;
assign v14458e0 = hlock1 & v14458db | !hlock1 & v14458df;
assign f2e4ff = hbusreq2 & f2e4fe | !hbusreq2 & f2ed9a;
assign v134cecc = hlock5 & v134d3b5 | !hlock5 & v134cec6;
assign v131be8f = hready_p & v131be8d | !hready_p & v131be8e;
assign v134d4af = hmaster1_p & v134d369 | !hmaster1_p & v134d4ae;
assign d30292 = hbusreq5_p & d30291 | !hbusreq5_p & d30277;
assign v16a1afc = hmaster1_p & v16a1afb | !hmaster1_p & v16a2672;
assign v1215444 = hmaster1_p & v1215443 | !hmaster1_p & v12153ec;
assign v1445f1c = hlock5 & v1445edb | !hlock5 & v1445f1b;
assign d30731 = hlock2_p & d3072d | !hlock2_p & d30730;
assign v1446480 = locked_p & v1446468 | !locked_p & v845542;
assign v151561f = hmaster1_p & v151561e | !hmaster1_p & v845570;
assign v12150e2 = hbusreq2_p & v12150e1 | !hbusreq2_p & v12150d3;
assign v12166c1 = hmaster0_p & v12164d7 | !hmaster0_p & v12164d5;
assign v134d444 = hbusreq2_p & v134d434 | !hbusreq2_p & v134d443;
assign d3075c = hbusreq2 & d30758 | !hbusreq2 & d3075b;
assign v121543a = hmaster1_p & v1215439 | !hmaster1_p & v121540f;
assign v121603e = hbusreq1 & v1216a98 | !hbusreq1 & v845542;
assign v134d22e = hmaster0_p & v134d22b | !hmaster0_p & v134d20a;
assign v121656e = hgrant5_p & v845542 | !hgrant5_p & v121656d;
assign v12153cf = hready & v845542 | !hready & v1668cba;
assign v134ce67 = hlock2 & v134ce64 | !hlock2 & v134ce66;
assign v1215757 = hbusreq1_p & v1215755 | !hbusreq1_p & v1215756;
assign v14462f6 = hgrant5_p & v1446426 | !hgrant5_p & v1446604;
assign d30738 = hlock2_p & d30737 | !hlock2_p & d30730;
assign v14465c0 = hlock4 & v144639c | !hlock4 & v14465bf;
assign v14460ca = hmaster2_p & v14460a2 | !hmaster2_p & v1446412;
assign v1446309 = hmaster1_p & v1446308 | !hmaster1_p & v144627e;
assign d2fd1d = hlock5_p & d2fd1b | !hlock5_p & !d2fd1c;
assign d30603 = hlock0_p & v1668c2d | !hlock0_p & v845542;
assign v12af1c4 = hready_p & v12af7e2 | !hready_p & v12af1c3;
assign v1214d89 = hbusreq2_p & v1214d87 | !hbusreq2_p & v1214d88;
assign v138a43e = hmaster0_p & v138a43c | !hmaster0_p & v138a43d;
assign v12160fe = hlock1_p & v12160f9 | !hlock1_p & v12160fd;
assign v12af3a8 = hbusreq1_p & v12af3a7 | !hbusreq1_p & !v84554a;
assign v1405aed = hgrant1_p & v1405a92 | !hgrant1_p & v1405aec;
assign d306ba = hbusreq2_p & d30677 | !hbusreq2_p & d306b8;
assign v12165a3 = hgrant5_p & v845542 | !hgrant5_p & v12165a2;
assign v1284d64 = hready_p & v1284d5a | !hready_p & !v1284d63;
assign a658c7 = hbusreq4_p & a658c6 | !hbusreq4_p & !v845542;
assign d30235 = hgrant2_p & d30234 | !hgrant2_p & d30219;
assign v12acfd0 = hmaster0_p & v12ad536 | !hmaster0_p & v12ad531;
assign v134ce80 = jx2_p & v134cdcf | !jx2_p & v134ce7f;
assign v12162f0 = hlock5_p & v12162ee | !hlock5_p & v12162ef;
assign d307d5 = hlock0_p & v845542 | !hlock0_p & d307d4;
assign v1216155 = hbusreq1_p & v1216154 | !hbusreq1_p & v845542;
assign v16a138b = hmaster1_p & v16a138a | !hmaster1_p & !v16a2672;
assign v1215da5 = hgrant2_p & v1215d86 | !hgrant2_p & v1215da4;
assign v1284d18 = hgrant4_p & v1284c8f | !hgrant4_p & v1446607;
assign v14058d4 = hgrant4_p & v140584b | !hgrant4_p & v14058d3;
assign v12ad5fe = hgrant5_p & v12ad4e4 | !hgrant5_p & v12ad5b1;
assign v12ad594 = decide_p & v12ad593 | !decide_p & !v845542;
assign v1405859 = hmaster2_p & v140583c | !hmaster2_p & v1405844;
assign d3028a = hlock2_p & d30289 | !hlock2_p & !v845542;
assign v1445f61 = hlock3 & v144673f | !hlock3 & v1445f5f;
assign v16a1962 = hbusreq0 & v16a1960 | !hbusreq0 & v16a1961;
assign a65369 = hmastlock_p & a65368 | !hmastlock_p & v845542;
assign v1668c6c = hbusreq4 & a658b5 | !hbusreq4 & v1668c6b;
assign v11ac6c9 = hready_p & v11ac6a3 | !hready_p & v11ac6c8;
assign v121540e = hbusreq5_p & v121540d | !hbusreq5_p & v12153de;
assign v1445d84 = hbusreq1 & v1445d82 | !hbusreq1 & v1445d83;
assign v14458cc = hbusreq2 & v14458c7 | !hbusreq2 & v14458cb;
assign v14460c5 = hlock2 & v14460a1 | !hlock2 & v14460c4;
assign v144608b = hmaster0_p & v1446404 | !hmaster0_p & v144608a;
assign v1552f8b = decide_p & v1553216 | !decide_p & v1552f8a;
assign v14463ec = hmaster2_p & v14463e4 | !hmaster2_p & v14463b7;
assign v1284cd4 = hbusreq5_p & v1284cd1 | !hbusreq5_p & !v1284cd3;
assign d308d0 = decide_p & d308cf | !decide_p & v845570;
assign v12166ed = hbusreq5_p & v12166ec | !hbusreq5_p & v845542;
assign v10d40b3 = hmaster1_p & v10d40b2 | !hmaster1_p & v10d3ffb;
assign v144618c = hbusreq2_p & v1446186 | !hbusreq2_p & v144618b;
assign v16a13f1 = hmaster1_p & v16a13f0 | !hmaster1_p & v16a1d7a;
assign v14459df = hgrant1_p & v14458e8 | !hgrant1_p & v14459de;
assign v1215b87 = hmaster2_p & v845542 | !hmaster2_p & v1215b86;
assign v121610a = hbusreq1_p & v1216109 | !hbusreq1_p & v845542;
assign v14457d1 = hlock5 & v14457ad | !hlock5 & v14457d0;
assign v1216521 = hbusreq1 & v1216a5a | !hbusreq1 & v845542;
assign v16a1ca0 = hmaster0_p & v16a1c9b | !hmaster0_p & v16a1c9f;
assign v1445f57 = hgrant2_p & v1445f55 | !hgrant2_p & v1445f56;
assign d2fc47 = decide_p & d2fc46 | !decide_p & v845570;
assign v1552d9b = hmaster1_p & v1552d9a | !hmaster1_p & v845542;
assign v1445452 = hbusreq3 & v1445450 | !hbusreq3 & v1445451;
assign v1215cdc = hlock2_p & v1215cdb | !hlock2_p & !v845542;
assign v15533af = hbusreq1 & v15533ad | !hbusreq1 & v15533ae;
assign d301e9 = hbusreq1 & d307ac | !hbusreq1 & v845542;
assign d2fd18 = hlock3_p & d2fd0e | !hlock3_p & d2fd17;
assign v15168ef = hbusreq2_p & v15168ee | !hbusreq2_p & !v845542;
assign v11e5970 = hgrant3_p & v11e5940 | !hgrant3_p & v11e596f;
assign d300d9 = hbusreq1 & d300d8 | !hbusreq1 & v84555a;
assign d2fb35 = hmaster2_p & d3068e | !hmaster2_p & d2fb34;
assign v1668c3d = hmaster0_p & v1668c3c | !hmaster0_p & v845570;
assign v1445911 = hmaster1_p & v1445910 | !hmaster1_p & v144590e;
assign v16a1b63 = hbusreq3 & v16a1b00 | !hbusreq3 & v16a1b62;
assign v14058ca = hmaster2_p & v14058c5 | !hmaster2_p & v1405845;
assign a65916 = hmaster0_p & a65915 | !hmaster0_p & a658e3;
assign v134d531 = hmaster0_p & v134d519 | !hmaster0_p & v845542;
assign v1445a5b = hmaster0_p & v14459a3 | !hmaster0_p & v1445a5a;
assign v1445b34 = hmaster1_p & v1445b33 | !hmaster1_p & v1445a32;
assign v1216536 = hgrant1_p & v1216522 | !hgrant1_p & v1216535;
assign v1445b84 = hlock2 & v144632f | !hlock2 & v1445b82;
assign v1446424 = hlock1 & v1446423 | !hlock1 & v1446421;
assign v16a1943 = hgrant5_p & v845542 | !hgrant5_p & v16a1942;
assign a662d2 = hmaster2_p & a662d0 | !hmaster2_p & a662ca;
assign v15168eb = hmaster0_p & v845570 | !hmaster0_p & v1668c3c;
assign v15530b3 = decide_p & v155342e | !decide_p & v15530a5;
assign v1215c78 = hbusreq2_p & v1215c76 | !hbusreq2_p & v1215c77;
assign a653ed = hmaster2_p & a65360 | !hmaster2_p & a653aa;
assign v1445adb = hbusreq2_p & v1445ad7 | !hbusreq2_p & v1445ada;
assign d30896 = hmaster2_p & d3084b | !hmaster2_p & !v845542;
assign v16a1e92 = hbusreq5_p & v16a207a | !hbusreq5_p & v16a1e91;
assign v10d428e = stateA1_p & v845542 | !stateA1_p & !v10d4264;
assign v15167f0 = decide_p & v15167ef | !decide_p & v845542;
assign v134d204 = hlock4_p & v134d1e8 | !hlock4_p & v845542;
assign v14463d6 = hready & v144639e | !hready & v144639c;
assign v144629f = hlock3 & v1446275 | !hlock3 & v144629b;
assign v12ad51e = hmaster2_p & a658c6 | !hmaster2_p & !v12ad51c;
assign v1446449 = hmaster0_p & v144639c | !hmaster0_p & v1446448;
assign v1214c39 = hmaster0_p & v1214c35 | !hmaster0_p & v1214c38;
assign v138945d = hbusreq2 & v138945c | !hbusreq2 & v1389ff2;
assign v144642e = hbusreq0 & v144642b | !hbusreq0 & v144642d;
assign v15533b8 = hgrant2_p & v1553380 | !hgrant2_p & v15533b7;
assign v10d3ffa = hmaster2_p & v10d3ff7 | !hmaster2_p & v10d3ff9;
assign d8076d = hgrant1_p & v845542 | !hgrant1_p & d8076c;
assign a653f8 = hgrant5_p & a65878 | !hgrant5_p & a653f5;
assign v14460b4 = hbusreq0 & v14460b3 | !hbusreq0 & v1446053;
assign bf1f95 = hgrant1_p & v845570 | !hgrant1_p & bf1f90;
assign v16a1cef = hbusreq0 & v16a1cee | !hbusreq0 & v16a1bcd;
assign v1445900 = hmaster2_p & v14458d2 | !hmaster2_p & v14458e2;
assign v138a434 = decide_p & v138a3c0 | !decide_p & !v138a406;
assign v1214df2 = hlock1_p & v1214df1 | !hlock1_p & v845547;
assign v1215365 = hmaster2_p & v845547 | !hmaster2_p & v1215364;
assign v1215cca = hgrant2_p & v1215c85 | !hgrant2_p & v1215cc9;
assign v14058a1 = hlock5_p & v140589e | !hlock5_p & v14058a0;
assign v1284cb7 = hbusreq2_p & v1284cb4 | !hbusreq2_p & v1284cb6;
assign v1445367 = hmaster1_p & v1445366 | !hmaster1_p & v1445a32;
assign v1445b65 = hmaster1_p & v1446308 | !hmaster1_p & v1446290;
assign v1214bb5 = hmaster0_p & v1215396 | !hmaster0_p & v12153b1;
assign v134ceca = hbusreq3 & v134cec8 | !hbusreq3 & v134cec9;
assign v12af9bc = hlock0_p & v845570 | !hlock0_p & v845542;
assign a65b40 = jx1_p & a65af9 | !jx1_p & a65b3f;
assign d30240 = hbusreq0 & d3023e | !hbusreq0 & d3023f;
assign v1284d59 = hbusreq2_p & v1284d54 | !hbusreq2_p & v1284d58;
assign v1515735 = hgrant5_p & v1515639 | !hgrant5_p & v1515733;
assign v134ce90 = hmaster0_p & v134ce8f | !hmaster0_p & v134d1e8;
assign v151697c = hbusreq2_p & v151697b | !hbusreq2_p & v845542;
assign d30796 = hgrant1_p & v845542 | !hgrant1_p & d30795;
assign d2ff03 = hmaster1_p & d2fec8 | !hmaster1_p & d2fee5;
assign v1446405 = hmaster0_p & v144639c | !hmaster0_p & v1446404;
assign d3060a = hmaster2_p & v16693aa | !hmaster2_p & v845542;
assign v1215d78 = hbusreq0 & v1215d76 | !hbusreq0 & v1215d77;
assign v1445b9e = hlock2 & v144632f | !hlock2 & v1445b9d;
assign f2f388 = hbusreq1 & v1668d82 | !hbusreq1 & v845542;
assign a6564d = hmaster2_p & a662ac | !hmaster2_p & a6564c;
assign a64713 = hready_p & a64712 | !hready_p & a64708;
assign d2f9d2 = hbusreq2_p & d2f9ce | !hbusreq2_p & d2f9d1;
assign v1215001 = hbusreq5_p & v1214ff9 | !hbusreq5_p & !v1215000;
assign v1214f11 = hmaster2_p & v1216a77 | !hmaster2_p & v845542;
assign v16693b0 = hlock3_p & v16693af | !hlock3_p & v845542;
assign v1216257 = hmaster1_p & v121623f | !hmaster1_p & !v121624b;
assign v1215036 = hgrant0_p & v1215465 | !hgrant0_p & !v845542;
assign v1445d94 = hbusreq0 & v1445d8d | !hbusreq0 & v1445d93;
assign v14457f8 = hmaster1_p & v14457f7 | !hmaster1_p & v1445e07;
assign v144554c = hgrant3_p & v1445541 | !hgrant3_p & v144554b;
assign v1445df5 = hbusreq1_p & v1446403 | !hbusreq1_p & v1445dec;
assign bf1f9f = hbusreq1_p & bf1f68 | !hbusreq1_p & bf1f9e;
assign v1215bc1 = hbusreq5_p & v1215bc0 | !hbusreq5_p & !v1216acf;
assign v14459f5 = hbusreq0_p & v144640a | !hbusreq0_p & v1446406;
assign v1515647 = stateG2_p & v845542 | !stateG2_p & ab8d68;
assign v1214c5b = hbusreq1_p & v1214c5a | !hbusreq1_p & v845547;
assign v138a306 = hmaster1_p & v138a305 | !hmaster1_p & v138a301;
assign v12ad557 = hbusreq2_p & v12ad555 | !hbusreq2_p & v12ad556;
assign v16a1d6d = hbusreq0 & v16a207a | !hbusreq0 & v16a2092;
assign v1553150 = hmaster2_p & v1553140 | !hmaster2_p & v845542;
assign d2fc70 = hbusreq2_p & d2fbff | !hbusreq2_p & d2fc6f;
assign v12aec16 = hbusreq3 & v12aec0b | !hbusreq3 & v12afe72;
assign d2f978 = hbusreq5_p & d2fe9e | !hbusreq5_p & d2f977;
assign v12162da = hmaster1_p & v1216262 | !hmaster1_p & !v121624b;
assign v12af988 = hbusreq4_p & v84554a | !hbusreq4_p & v845542;
assign d2fb1b = hgrant5_p & d3068e | !hgrant5_p & d2fae3;
assign d306b8 = hgrant2_p & d30684 | !hgrant2_p & d306b7;
assign d2fd2c = hgrant2_p & v845542 | !hgrant2_p & d2fd2b;
assign v1445e0b = hbusreq0 & v1445e09 | !hbusreq0 & v1445e0a;
assign v1445e8a = hbusreq4_p & v14465f9 | !hbusreq4_p & v144660d;
assign d30824 = hgrant5_p & v84554e | !hgrant5_p & d307c0;
assign v1214c7d = hmaster1_p & v1214c7c | !hmaster1_p & v1214c74;
assign v144662b = hmaster2_p & v14465f5 | !hmaster2_p & v144662a;
assign v1445aa1 = hmaster1_p & v1445a5b | !hmaster1_p & v1445a9b;
assign v166959f = hmaster1_p & v166959e | !hmaster1_p & v845542;
assign v12ad31d = hgrant1_p & d30690 | !hgrant1_p & v12ad31c;
assign v155304f = hbusreq1 & v155304e | !hbusreq1 & v1553217;
assign v10d4086 = hgrant2_p & v10d4081 | !hgrant2_p & v10d4085;
assign v1553510 = hlock2 & v155321a | !hlock2 & v155350f;
assign v1216af8 = hmaster0_p & v1216ad1 | !hmaster0_p & v1216af7;
assign v1515c80 = hbusreq4_p & v1515c7f | !hbusreq4_p & !v845542;
assign a65864 = hbusreq1_p & a65852 | !hbusreq1_p & a65863;
assign v16a1398 = hbusreq5 & v16a138e | !hbusreq5 & v16a1397;
assign v1446098 = hmaster1_p & v14465aa | !hmaster1_p & v1445fef;
assign v1214c50 = hgrant4_p & v1214c48 | !hgrant4_p & v845542;
assign v121533f = hbusreq3 & v1215337 | !hbusreq3 & v121533e;
assign v1445d9c = hmaster2_p & v14463b9 | !hmaster2_p & v1445d9b;
assign a6563e = hgrant5_p & a653ab | !hgrant5_p & !a6563c;
assign v16a1f9d = hbusreq3 & v16a1f99 | !hbusreq3 & !v16a1f9c;
assign a65394 = locked_p & a65393 | !locked_p & a65861;
assign v138a037 = hbusreq3 & v138a034 | !hbusreq3 & v138a404;
assign v151572a = hgrant1_p & v1515712 | !hgrant1_p & v1515729;
assign v1284ceb = hgrant1_p & v1284cea | !hgrant1_p & !v1405845;
assign v15155ec = hlock2_p & v15155eb | !hlock2_p & v845542;
assign v16a129e = hmaster1_p & v16a129d | !hmaster1_p & !v16a2672;
assign d2fad7 = hbusreq1 & d2f96b | !hbusreq1 & !d30660;
assign v1214dcb = jx2_p & v1215344 | !jx2_p & v1214dca;
assign v13897de = hgrant5_p & v13897dd | !hgrant5_p & !v845542;
assign v1215053 = hbusreq0 & v1215049 | !hbusreq0 & v1215052;
assign d30210 = hgrant1_p & d30205 | !hgrant1_p & d307e1;
assign v121535f = hmaster2_p & v845542 | !hmaster2_p & v121535e;
assign v1284cf0 = hgrant5_p & v1284cee | !hgrant5_p & !v1284cef;
assign v1446445 = hmaster2_p & v144639c | !hmaster2_p & v1446444;
assign d2fc01 = hbusreq2_p & d2fbff | !hbusreq2_p & d2fc00;
assign v134d516 = hmaster2_p & v845542 | !hmaster2_p & v134d4e8;
assign v16a1e4b = hmaster1_p & v16a1e23 | !hmaster1_p & v16a1f96;
assign v1446183 = hmaster1_p & v1446182 | !hmaster1_p & v1445fde;
assign d80775 = hgrant5_p & d80770 | !hgrant5_p & !d80774;
assign f2f35c = hbusreq5_p & f2f35a | !hbusreq5_p & f2f35b;
assign v1214ef0 = hmaster2_p & v1216a67 | !hmaster2_p & v845542;
assign f2f3e1 = hbusreq5 & f2f3b7 | !hbusreq5 & f2f3e0;
assign v1214cd3 = hgrant4_p & v1214cd2 | !hgrant4_p & v845572;
assign v1284ce8 = hbusreq2_p & v1284ce1 | !hbusreq2_p & v1284ce7;
assign v14453f4 = hbusreq2_p & v144627f | !hbusreq2_p & v14453f3;
assign v1215c52 = hbusreq3 & v1215c51 | !hbusreq3 & v845542;
assign v121656c = hgrant1_p & v1216522 | !hgrant1_p & v121656b;
assign v12ad5a2 = hmastlock_p & v12ad5a1 | !hmastlock_p & v10d3fd3;
assign v144549b = hbusreq2 & v1445494 | !hbusreq2 & v144549a;
assign v1216177 = hgrant5_p & v1216029 | !hgrant5_p & !v1216175;
assign v1445eae = hmaster2_p & v144639c | !hmaster2_p & v1446606;
assign v14465f7 = hlock0_p & v144639c | !hlock0_p & v14465f6;
assign f2f37f = hmaster2_p & f2f37b | !hmaster2_p & f2f37e;
assign v1215d28 = hmaster2_p & v16a1bc6 | !hmaster2_p & v1216a93;
assign v14466e4 = hmaster1_p & v14466e3 | !hmaster1_p & v14463ef;
assign v16a1373 = hbusreq3 & v16a1332 | !hbusreq3 & v16a1372;
assign v16a1af2 = hready_p & v16a1af0 | !hready_p & !v16a1af1;
assign v1214f0a = hgrant5_p & v16a2243 | !hgrant5_p & v1214edf;
assign v138a312 = hlock5_p & v138a311 | !hlock5_p & !v845542;
assign v16a223e = hmaster2_p & v16a223d | !hmaster2_p & !v845542;
assign v1284d52 = hbusreq2_p & v1284d47 | !hbusreq2_p & v1284d51;
assign v1214d66 = hbusreq2_p & v1214c1d | !hbusreq2_p & v1214d65;
assign v15167c2 = hlock2_p & v15167c1 | !hlock2_p & v845542;
assign v1446165 = hgrant2_p & v1446162 | !hgrant2_p & v1446164;
assign v12af7f7 = hbusreq5_p & v845542 | !hbusreq5_p & v12af7f6;
assign d2faea = hbusreq4_p & d300c1 | !hbusreq4_p & d306a3;
assign v1214d47 = hbusreq1_p & v12153a6 | !hbusreq1_p & v1214d46;
assign d2fe80 = hbusreq4_p & d2fe7f | !hbusreq4_p & v845542;
assign d30874 = hbusreq5_p & d30752 | !hbusreq5_p & d30654;
assign v12ad5d4 = hlock0_p & v1668d6e | !hlock0_p & v12ad5d3;
assign v155308f = hbusreq2_p & v1553061 | !hbusreq2_p & v155308e;
assign d2fd26 = hlock2_p & v845542 | !hlock2_p & d2fd25;
assign v14457e4 = hmaster0_p & v1445eba | !hmaster0_p & v1445ecc;
assign v12150d4 = hlock2_p & v12150d2 | !hlock2_p & v12150d3;
assign v1446245 = hlock3 & v1446224 | !hlock3 & v1446244;
assign v12ad02b = hbusreq5_p & v12ad613 | !hbusreq5_p & !v12ad02a;
assign a65686 = hbusreq2_p & a65684 | !hbusreq2_p & a65685;
assign f2e4e0 = hready_p & f2e4df | !hready_p & f2e4d4;
assign v1216abe = hbusreq1_p & v1216abd | !hbusreq1_p & v845547;
assign v12ad634 = hbusreq0 & v12ad501 | !hbusreq0 & v12af73f;
assign v10d4056 = hgrant5_p & v10d3feb | !hgrant5_p & v10d4055;
assign v138a354 = hbusreq5_p & v138a353 | !hbusreq5_p & !v845542;
assign f2f2d6 = hmaster2_p & f2f2d3 | !hmaster2_p & f2f2d5;
assign v15157b1 = hgrant5_p & v845542 | !hgrant5_p & !v15157af;
assign f2ed98 = hmaster1_p & f2ed95 | !hmaster1_p & f2ed97;
assign v15155e9 = hbusreq0 & v15155e8 | !hbusreq0 & v845568;
assign v1214f3a = hgrant2_p & v845542 | !hgrant2_p & v1214f39;
assign d2fcac = hmaster0_p & d305eb | !hmaster0_p & v16693aa;
assign v1284d35 = hmaster1_p & v1284d34 | !hmaster1_p & v1284ca7;
assign d2fb52 = hmaster0_p & d2fb50 | !hmaster0_p & d2fb51;
assign v138981c = hbusreq5 & v13897f1 | !hbusreq5 & v1389819;
assign v1445824 = hmaster1_p & v14457e2 | !hmaster1_p & v1445e28;
assign v1215d64 = hmaster0_p & v1215d63 | !hmaster0_p & v12164d4;
assign d2fc26 = hbusreq0 & d2fc25 | !hbusreq0 & !v845542;
assign v16a19e0 = hmaster0_p & v16a19d3 | !hmaster0_p & v16a19df;
assign d30728 = hlock1_p & v845542 | !hlock1_p & !d30727;
assign v1668d9f = hgrant5_p & v1668d9a | !hgrant5_p & v1668d9d;
assign v121601c = hready & v845580 | !hready & v845542;
assign v134d3db = hbusreq4_p & v134d27c | !hbusreq4_p & v134d3da;
assign v1215336 = hbusreq2_p & v1215335 | !hbusreq2_p & v1215332;
assign v12ad023 = hgrant2_p & v12acff2 | !hgrant2_p & v12ad022;
assign v12167a9 = hgrant2_p & v12167a7 | !hgrant2_p & v12167a8;
assign v1668c88 = hmaster1_p & v1668c87 | !hmaster1_p & v1668c72;
assign v1445880 = hbusreq0 & v1445878 | !hbusreq0 & v144587f;
assign v1668d24 = hbusreq4 & a65851 | !hbusreq4 & v845570;
assign v1216239 = hgrant2_p & v1216234 | !hgrant2_p & v1216238;
assign v1216ab3 = hbusreq5_p & v1216ab2 | !hbusreq5_p & v845542;
assign v138a359 = hmaster0_p & v138a34b | !hmaster0_p & v138a32d;
assign v144607d = hgrant5_p & v1445fe0 | !hgrant5_p & v144607c;
assign v134d381 = hlock1 & v134d380 | !hlock1 & v134d37f;
assign v144610e = hbusreq2_p & v144610a | !hbusreq2_p & v144610d;
assign v12ad4f6 = hlock0_p & v10d3fdf | !hlock0_p & v845542;
assign a653f9 = hmaster2_p & a65360 | !hmaster2_p & !a653a9;
assign v16a13fa = hgrant2_p & v845542 | !hgrant2_p & !v16a13f9;
assign d30618 = hbusreq2 & d30610 | !hbusreq2 & d30617;
assign v1405b31 = hbusreq2_p & v1405b2b | !hbusreq2_p & v1405b30;
assign v12153ae = hlock2_p & v12153aa | !hlock2_p & v12153ad;
assign v12ad5fc = hbusreq2_p & v12ad5f6 | !hbusreq2_p & !v12ad5fb;
assign d2fc6b = hbusreq5_p & d2fbfa | !hbusreq5_p & d2fc6a;
assign d3024f = hbusreq0 & d3024d | !hbusreq0 & d3024e;
assign d2fc2d = hbusreq4_p & d2fb69 | !hbusreq4_p & d2fc2c;
assign d80757 = stateG3_2_p & v845542 | !stateG3_2_p & !v84556c;
assign d8073d = hbusreq1_p & d8073c | !hbusreq1_p & !v845542;
assign d3027f = hgrant5_p & v845542 | !hgrant5_p & !d30669;
assign v1284d3f = hbusreq2_p & v1284d36 | !hbusreq2_p & v1284d3e;
assign v12ad4f1 = hmaster2_p & v12ad4f0 | !hmaster2_p & a653c8;
assign v16a1ac8 = hbusreq3 & v16a1ac3 | !hbusreq3 & v16a1ac7;
assign v16a2238 = stateA1_p & v16a2237 | !stateA1_p & d8075a;
assign d307ab = hlock5_p & d307a9 | !hlock5_p & d307aa;
assign v140588a = hlock4_p & v140583d | !hlock4_p & v140583c;
assign v1405b46 = hmaster1_p & v1405b45 | !hmaster1_p & !v1405a94;
assign v10d40de = hbusreq3_p & v10d4099 | !hbusreq3_p & !v10d40dd;
assign v1516854 = hready_p & v1516806 | !hready_p & !v1516853;
assign v16a1d64 = hgrant2_p & v845542 | !hgrant2_p & !v16a1d63;
assign v138a462 = hbusreq2_p & v138a460 | !hbusreq2_p & v138a461;
assign a653d9 = locked_p & a653d8 | !locked_p & v845542;
assign v1515c7f = hlock4_p & v1515c7e | !hlock4_p & f2f4b0;
assign bf1f58 = hmaster0_p & v845542 | !hmaster0_p & bf1f4d;
assign a653d8 = hburst0 & v845542 | !hburst0 & a653d7;
assign v1216196 = hgrant5_p & v121601d | !hgrant5_p & v1216132;
assign v10d402c = hbusreq1_p & v10d402a | !hbusreq1_p & !v10d402b;
assign v138a4a2 = hbusreq3_p & v138a436 | !hbusreq3_p & v138a4a1;
assign d30891 = hgrant1_p & v84554c | !hgrant1_p & d30890;
assign v138a399 = hmaster1_p & v138a398 | !hmaster1_p & v138a341;
assign a65478 = hmaster1_p & a65465 | !hmaster1_p & a65476;
assign v1445418 = hmaster1_p & v1445417 | !hmaster1_p & v1445bb7;
assign d2fb6d = hlock0_p & v845542 | !hlock0_p & !d305ef;
assign v151574e = hbusreq1 & v10d3fdf | !hbusreq1 & v845542;
assign v1446012 = hgrant1_p & v845542 | !hgrant1_p & v1446011;
assign d2fc4e = hbusreq1_p & d2fbd1 | !hbusreq1_p & d2fc4d;
assign v12ad666 = hmaster0_p & v12ad661 | !hmaster0_p & v12ad665;
assign v12ad4de = hmaster1_p & v12ad4d3 | !hmaster1_p & v12ad4dd;
assign v16a1e58 = hready_p & v16a1e0e | !hready_p & v16a1e57;
assign v1446712 = hmaster0_p & v144667f | !hmaster0_p & v1446404;
assign v14058f6 = stateG10_5_p & v14058f5 | !stateG10_5_p & v14058ef;
assign v14466bd = hbusreq2 & v14466bb | !hbusreq2 & v14466bc;
assign v16a2088 = hlock5_p & v16a2082 | !hlock5_p & v16a2087;
assign v1446649 = hbusreq0 & v1446644 | !hbusreq0 & v1446648;
assign v1668d5a = hgrant1_p & v1668d46 | !hgrant1_p & v1668d59;
assign v15157ec = hgrant5_p & v1668dc2 | !hgrant5_p & v1515758;
assign v1668c55 = decide_p & v1668c52 | !decide_p & v845542;
assign v15532c4 = hgrant4_p & v1553138 | !hgrant4_p & v845542;
assign v1216105 = hgrant4_p & v12160ed | !hgrant4_p & v1216534;
assign v138a338 = hmaster2_p & v845542 | !hmaster2_p & v138a337;
assign v1214c92 = hmaster0_p & v1214c8f | !hmaster0_p & v1214c91;
assign v16a1d47 = hgrant1_p & v84554d | !hgrant1_p & v16a1bd3;
assign v1552d5d = hbusreq5_p & v1553392 | !hbusreq5_p & v1552d5c;
assign v14462fe = hlock0 & v14462f7 | !hlock0 & v14462fa;
assign v134cdc8 = hlock5 & v134d276 | !hlock5 & v134cdc7;
assign v12ad678 = hbusreq1_p & a658c6 | !hbusreq1_p & v12ad677;
assign v1214f12 = hgrant5_p & v1214f11 | !hgrant5_p & v1216547;
assign v134d50c = hgrant5_p & v845542 | !hgrant5_p & v134d50b;
assign v10a1541 = hgrant2_p & v845542 | !hgrant2_p & !v10a1540;
assign v1668c4f = hmaster0_p & v1668c4e | !hmaster0_p & v845542;
assign v1214cd8 = hmaster0_p & v1214cd1 | !hmaster0_p & v1214cd7;
assign v1214fb4 = hmaster2_p & v12157b1 | !hmaster2_p & v121572b;
assign v1215b9e = hmaster2_p & v121611f | !hmaster2_p & v1215b9c;
assign v1515792 = hgrant4_p & a662a9 | !hgrant4_p & v1515791;
assign d2fc42 = hmaster1_p & d2fc31 | !hmaster1_p & d2fc41;
assign v1215765 = hgrant0_p & v1215764 | !hgrant0_p & v845542;
assign v134d38b = hgrant5_p & v845542 | !hgrant5_p & v134d38a;
assign v1214dc0 = hgrant2_p & v1214db2 | !hgrant2_p & v1214dbf;
assign v12ad677 = hbusreq4_p & a658c6 | !hbusreq4_p & v12ad676;
assign v14465f1 = hbusreq4_p & v14465b1 | !hbusreq4_p & v14465cd;
assign v12afe50 = hmaster2_p & v12afe46 | !hmaster2_p & v12afe4f;
assign v16a1ce6 = hbusreq3 & v16a1ce0 | !hbusreq3 & v16a1ce5;
assign v1405b23 = hgrant4_p & v1405a88 | !hgrant4_p & !v1405b22;
assign d30917 = hbusreq0 & d305fc | !hbusreq0 & d30916;
assign v12153a4 = hlock0_p & v1216ad4 | !hlock0_p & v12153a3;
assign d30801 = hgrant5_p & d30708 | !hgrant5_p & !d307ff;
assign v16a13ef = hbusreq0 & v16a13eb | !hbusreq0 & v16a13ee;
assign v1215be6 = hbusreq1_p & v845547 | !hbusreq1_p & v121601f;
assign v14462f3 = hbusreq5_p & v14465e3 | !hbusreq5_p & v14462f2;
assign a662a9 = hbusreq4_p & v845570 | !hbusreq4_p & !v845542;
assign v1214d29 = hgrant2_p & v1214d16 | !hgrant2_p & v1214d28;
assign f2f433 = hbusreq5_p & f2f380 | !hbusreq5_p & f2f432;
assign v140593b = hbusreq2_p & v1405936 | !hbusreq2_p & v140593a;
assign v14457c7 = hbusreq2_p & v14457c3 | !hbusreq2_p & v14457c6;
assign d80780 = hgrant1_p & v845542 | !hgrant1_p & d8077f;
assign v1446188 = hmaster1_p & v1446187 | !hmaster1_p & v1445fde;
assign d300c1 = hlock4_p & v845542 | !hlock4_p & a65382;
assign v15160fb = hlock2_p & v15160fa | !hlock2_p & v845542;
assign a65856 = stateG3_2_p & v88d3e4 | !stateG3_2_p & a65854;
assign d30277 = hgrant5_p & v845542 | !hgrant5_p & !d30275;
assign v1445ef7 = hmaster1_p & v1445ec4 | !hmaster1_p & v1445e28;
assign d3022d = hmaster0_p & d301dd | !hmaster0_p & d3022c;
assign d30230 = hbusreq2_p & d3021a | !hbusreq2_p & !d3022f;
assign v1215d82 = hmaster1_p & v1215d81 | !hmaster1_p & v1215d79;
assign v1515658 = hbusreq1_p & v1515657 | !hbusreq1_p & !v1668c63;
assign d8075e = busreq_p & d80756 | !busreq_p & !d8075d;
assign v1445acd = hlock3 & v1445abf | !hlock3 & v1445acb;
assign f2f21a = hbusreq1 & a66275 | !hbusreq1 & !v1668c2d;
assign v138a309 = hbusreq5_p & v138a308 | !hbusreq5_p & v845542;
assign v134cea3 = hlock2_p & v134ce91 | !hlock2_p & v134cea2;
assign v16a1ce8 = decide_p & v16a1ce7 | !decide_p & !v16a2065;
assign d30779 = hbusreq5 & d30770 | !hbusreq5 & d30778;
assign v1445e6c = hgrant1_p & v1445e5c | !hgrant1_p & v1445e6b;
assign d2fc6d = hmaster0_p & d2fc65 | !hmaster0_p & d2fc6c;
assign v16695bc = decide_p & v16695bb | !decide_p & !v845542;
assign v1446411 = hmaster2_p & v1446403 | !hmaster2_p & v1446410;
assign v1446644 = hbusreq5_p & v1446641 | !hbusreq5_p & v1446643;
assign d2fb83 = hlock0_p & v845542 | !hlock0_p & !v1668c2d;
assign v1445ed5 = hgrant2_p & v1445ed2 | !hgrant2_p & v1445ed4;
assign v14453c8 = jx2_p & v144586b | !jx2_p & v14453c7;
assign f2f391 = hbusreq5_p & f2f38f | !hbusreq5_p & f2f390;
assign v12153ac = hmaster0_p & v1215396 | !hmaster0_p & v12153ab;
assign v14463a7 = hbusreq5_p & v14463a4 | !hbusreq5_p & v14463a6;
assign v12ae6da = decide_p & v12afe3d | !decide_p & v845542;
assign v1284d14 = hmaster2_p & v14465d8 | !hmaster2_p & v1284d10;
assign v1216019 = hmaster0_p & v1216018 | !hmaster0_p & v845542;
assign v14466cd = hmaster1_p & v14466cc | !hmaster1_p & v14463c2;
assign v1216569 = hlock0_p & v1216568 | !hlock0_p & v845547;
assign v144646f = hbusreq1_p & v1446398 | !hbusreq1_p & v144646e;
assign v1445777 = hbusreq0 & v1445775 | !hbusreq0 & v1445776;
assign v1405b57 = hmaster1_p & v1405af7 | !hmaster1_p & v1405b09;
assign v12ad679 = hmaster2_p & v12ad675 | !hmaster2_p & v12ad678;
assign v10d42c7 = hgrant4_p & v10d401a | !hgrant4_p & v10d42c6;
assign d80734 = hmaster2_p & v845542 | !hmaster2_p & !d80733;
assign v1214fea = hgrant4_p & v845542 | !hgrant4_p & v12153b4;
assign d2fb3d = hmaster1_p & d2f99c | !hmaster1_p & d2fb3c;
assign v121621d = hgrant5_p & v12160df | !hgrant5_p & v121621c;
assign v1214f17 = hlock2_p & v1214f10 | !hlock2_p & v1214f16;
assign v1515843 = hgrant5_p & v845542 | !hgrant5_p & !v1515833;
assign v11e5958 = hgrant4_p & v845542 | !hgrant4_p & !v11e5957;
assign v12167aa = hbusreq2_p & v12167a5 | !hbusreq2_p & v12167a9;
assign v1668d22 = hbusreq1 & v10d3fd8 | !hbusreq1 & !v845542;
assign d30263 = hbusreq3 & d3025f | !hbusreq3 & v845542;
assign a656b0 = hbusreq2 & a656ab | !hbusreq2 & a656ae;
assign d307ad = hlock1_p & d307ac | !hlock1_p & !v845542;
assign v1405b60 = hmaster1_p & v1405b2d | !hmaster1_p & v1405b29;
assign v138a356 = hmaster1_p & v138a355 | !hmaster1_p & v138a341;
assign v155309c = hgrant2_p & v155308d | !hgrant2_p & v155309a;
assign v1445d86 = hmaster2_p & v144639c | !hmaster2_p & v1445d85;
assign v16a2096 = hmaster1_p & v16a208d | !hmaster1_p & v16a2095;
assign d3024c = hbusreq0 & d30246 | !hbusreq0 & d3024b;
assign v1389efe = hgrant3_p & v1389d78 | !hgrant3_p & v1389efd;
assign v1445a15 = hbusreq4_p & v144639c | !hbusreq4_p & v144660b;
assign v1215413 = hbusreq2_p & v1215412 | !hbusreq2_p & v1215411;
assign v16a1d33 = hbusreq2 & v16a1d31 | !hbusreq2 & v16a1d32;
assign v138a393 = hmaster2_p & v138a32b | !hmaster2_p & !a658d4;
assign d2fd16 = hbusreq2 & d2fd15 | !hbusreq2 & d2fcd8;
assign v12162d5 = hbusreq2_p & v12162d4 | !hbusreq2_p & v12162d1;
assign a653d5 = hgrant5_p & a653d4 | !hgrant5_p & a653d1;
assign v1445e1c = hmaster1_p & v1445de8 | !hmaster1_p & v1445e1b;
assign d2fc4b = hgrant0_p & v84554a | !hgrant0_p & d2fc4a;
assign d2fb39 = hmaster2_p & d3068e | !hmaster2_p & d2fb38;
assign v1516805 = hbusreq5 & v15167fe | !hbusreq5 & v1516804;
assign v14457c4 = hmaster1_p & v14457a3 | !hmaster1_p & v1445e28;
assign d2f9bb = hlock2_p & d2f9ba | !hlock2_p & d2f997;
assign v12ad5d8 = hbusreq4_p & v12ad5d6 | !hbusreq4_p & !v12ad5d7;
assign v1214d27 = hbusreq0 & v1214cee | !hbusreq0 & v1216718;
assign v1668dce = hgrant5_p & v845570 | !hgrant5_p & v1668d86;
assign v1214c3c = hbusreq0 & v1214c3b | !hbusreq0 & v16a2243;
assign v14457bb = hmaster1_p & v144578e | !hmaster1_p & v1445e28;
assign d300f0 = hgrant5_p & d2fe9e | !hgrant5_p & d300ee;
assign v14465eb = hlock4 & v14465bc | !hlock4 & v14465bf;
assign f2f3fc = hmaster1_p & f2f3fb | !hmaster1_p & f2f2db;
assign v151575b = hmaster2_p & v151575a | !hmaster2_p & v1515757;
assign v134cd82 = hgrant2_p & v134d364 | !hgrant2_p & v134cd81;
assign v134ce42 = hgrant1_p & v845542 | !hgrant1_p & v134ce41;
assign a65677 = hbusreq0 & a65672 | !hbusreq0 & a65676;
assign f2f39b = hmaster2_p & f2f39a | !hmaster2_p & !v845542;
assign v12166da = hbusreq0_p & v12164d3 | !hbusreq0_p & !v12166ce;
assign v121620a = hmaster2_p & v12160d3 | !hmaster2_p & v845542;
assign v16a13c5 = hmaster0_p & v16a13c4 | !hmaster0_p & v16a13a8;
assign v1668c39 = hgrant3_p & v84556e | !hgrant3_p & v845542;
assign v1445dc8 = hbusreq2 & v1445dc1 | !hbusreq2 & v1445dc7;
assign a653d4 = hmaster2_p & v845542 | !hmaster2_p & a653c5;
assign v16695b1 = decide_p & v16695b0 | !decide_p & v845542;
assign v1214ef3 = hlock5_p & v1214ef1 | !hlock5_p & !v1214ef2;
assign v1446243 = hlock2 & v1446224 | !hlock2 & v144623e;
assign d30914 = hlock5_p & d30912 | !hlock5_p & !d30913;
assign v121505a = hmaster2_p & v121502a | !hmaster2_p & v121503e;
assign v1389d59 = hlock5_p & v1389d58 | !hlock5_p & !v845542;
assign v134d51e = hmaster0_p & v134d4f6 | !hmaster0_p & v134d510;
assign v1446046 = hbusreq1_p & v1446045 | !hbusreq1_p & v1446406;
assign v16a1971 = hgrant5_p & v845542 | !hgrant5_p & v16a1970;
assign v1516101 = hmaster0_p & v845542 | !hmaster0_p & v1516100;
assign v12ad5fb = hgrant2_p & v12ad5fa | !hgrant2_p & !v12ad5ee;
assign d2fc23 = hbusreq0 & v84554a | !hbusreq0 & !v845542;
assign v134cec4 = hbusreq2 & v134cec3 | !hbusreq2 & v134d3b5;
assign v12afdaa = hmaster2_p & v845542 | !hmaster2_p & v12afda9;
assign v12160e1 = hmaster1_p & v12160d6 | !hmaster1_p & v12160e0;
assign d3082a = hbusreq5_p & d30829 | !hbusreq5_p & d30828;
assign v1214e6f = hgrant1_p & v1214e6e | !hgrant1_p & v1216aea;
assign c50efb = hbusreq2_p & v845542 | !hbusreq2_p & v845576;
assign v1668d41 = hbusreq0 & v1668d3a | !hbusreq0 & v1668d40;
assign v1214c8a = hgrant5_p & v1214c89 | !hgrant5_p & v1214c5d;
assign v1445a39 = hmaster0_p & v14458d4 | !hmaster0_p & v1445a38;
assign d3026b = hgrant5_p & v845542 | !hgrant5_p & !d30269;
assign v1553519 = hready_p & v1553444 | !hready_p & v1553518;
assign d307e4 = hbusreq1_p & d307e3 | !hbusreq1_p & d30661;
assign v16a16b4 = hgrant3_p & v16a1e8a | !hgrant3_p & v16a16b3;
assign v144649d = hgrant1_p & v845542 | !hgrant1_p & v144649c;
assign f2f3ed = hbusreq3 & f2f3ea | !hbusreq3 & !f2f3ec;
assign v845552 = hlock2_p & v845542 | !hlock2_p & !v845542;
assign v1216301 = hmaster2_p & v1216ad6 | !hmaster2_p & v1216aec;
assign v15156b0 = hbusreq0 & v1668cd2 | !hbusreq0 & v15156af;
assign v12ad5a1 = stateA1_p & v84557e | !stateA1_p & v12ad5a0;
assign v1216300 = hbusreq5_p & v12162ff | !hbusreq5_p & v12162fe;
assign v14463c9 = hlock0 & v14463c8 | !hlock0 & v14463c6;
assign v1214e10 = hmaster1_p & v1214dea | !hmaster1_p & v1214e0f;
assign v16a1397 = hbusreq3 & v16a1393 | !hbusreq3 & v16a1396;
assign v14058ec = hgrant5_p & v140587e | !hgrant5_p & v14058eb;
assign d2fc0e = hlock5_p & d2fc0d | !hlock5_p & d2fbe3;
assign v10d402f = hgrant0_p & v10d402e | !hgrant0_p & v10d3fdf;
assign v1284d30 = hbusreq2_p & v1284d2d | !hbusreq2_p & v1284d2f;
assign v1445be8 = hready_p & v1445bca | !hready_p & v1445be7;
assign v138a4a0 = hready_p & v138a48e | !hready_p & !v138a49f;
assign f2e502 = hgrant3_p & f2e4e9 | !hgrant3_p & f2e501;
assign v1445a56 = hbusreq0 & v1445a55 | !hbusreq0 & v1445a3e;
assign v16a1e02 = hbusreq3 & v16a1d33 | !hbusreq3 & v16a1e01;
assign d3081d = hbusreq0 & d30818 | !hbusreq0 & d3081c;
assign v12153a1 = hbusreq5_p & v12153a0 | !hbusreq5_p & v121539f;
assign v1216165 = hgrant4_p & v1216150 | !hgrant4_p & v1216164;
assign d3075e = hmaster1_p & d30747 | !hmaster1_p & d30754;
assign v14457e9 = hmaster1_p & v14457e4 | !hmaster1_p & v1445eaa;
assign v1284d34 = hmaster0_p & v1284cad | !hmaster0_p & v1284ca9;
assign v134d3e2 = hmaster1_p & v134d3e1 | !hmaster1_p & v134d294;
assign d80784 = hmaster1_p & d8076f | !hmaster1_p & !d80783;
assign v16a131f = locked_p & v845542 | !locked_p & !v16a131e;
assign a65923 = hbusreq2_p & a65921 | !hbusreq2_p & a65922;
assign d306b3 = hbusreq5_p & d3065f | !hbusreq5_p & !d306b2;
assign v16a183f = hbusreq4 & v16a1afa | !hbusreq4 & !v845542;
assign a65647 = hgrant5_p & a653d4 | !hgrant5_p & a65646;
assign v1445a7b = hmaster2_p & v1445a4c | !hmaster2_p & v14458e5;
assign f2f2e4 = hmaster0_p & f2f2cc | !hmaster0_p & f2f2e3;
assign v16a12f5 = hgrant2_p & v845542 | !hgrant2_p & !v16a12f4;
assign v1446716 = hbusreq2_p & v1446713 | !hbusreq2_p & v1446715;
assign v121610d = hgrant4_p & v12160fa | !hgrant4_p & v845542;
assign v1445b22 = hmaster1_p & v1445b06 | !hmaster1_p & v144591b;
assign v12afe57 = hmaster2_p & v12afe46 | !hmaster2_p & v12afe56;
assign d2fe81 = hmaster2_p & d2fe7b | !hmaster2_p & d2fe80;
assign v12acfdc = hmaster1_p & v12ad67b | !hmaster1_p & v12acfdb;
assign stateG2 = !d807c0;
assign d80790 = hgrant5_p & d8078f | !hgrant5_p & d8078d;
assign a6562e = hgrant1_p & a653ae | !hgrant1_p & !a6562d;
assign v14459e8 = hmaster2_p & v14465b3 | !hmaster2_p & v14459e7;
assign v12ad4f3 = hmaster2_p & v12ad4f0 | !hmaster2_p & v10d3fd8;
assign d80772 = hbusreq1_p & d80771 | !hbusreq1_p & !v845542;
assign a6588f = hbusreq4_p & a6588d | !hbusreq4_p & v845542;
assign d807b5 = hgrant3_p & d80766 | !hgrant3_p & d807b4;
assign a65644 = hbusreq1_p & a653cf | !hbusreq1_p & a65643;
assign hgrant3 = v16695ca;
assign v155341a = hbusreq2_p & v15533b8 | !hbusreq2_p & v1553419;
assign a65869 = hbusreq5_p & a65866 | !hbusreq5_p & a65867;
assign a65883 = hburst1_p & v845542 | !hburst1_p & a6587f;
assign v1445908 = hbusreq0 & v1445907 | !hbusreq0 & v1445900;
assign v1445efc = hmaster1_p & v1445ee0 | !hmaster1_p & v1445e28;
assign v1215cf8 = hbusreq5_p & v1215cf7 | !hbusreq5_p & v1215cc3;
assign v1445b73 = hmaster2_p & v1446677 | !hmaster2_p & v1446410;
assign v1668c53 = decide_p & v1668c52 | !decide_p & !v845542;
assign a65457 = hready_p & a65455 | !hready_p & a65456;
assign v144664a = hlock0 & v1446649 | !hlock0 & v1446644;
assign v1445ac3 = hmaster1_p & v1445ac2 | !hmaster1_p & v144589f;
assign v1216181 = hbusreq2_p & v1216171 | !hbusreq2_p & !v1216180;
assign v1553429 = hbusreq4_p & v1553140 | !hbusreq4_p & v1553428;
assign v1445549 = hbusreq2_p & v1445546 | !hbusreq2_p & v1445548;
assign v144598e = hmaster0_p & v14458d4 | !hmaster0_p & v14458d3;
assign v14058fe = hmaster2_p & v14058fa | !hmaster2_p & v14058fd;
assign v1214c74 = hmaster0_p & v1214c65 | !hmaster0_p & v1214c73;
assign d2fbf6 = hgrant1_p & d2fbcb | !hgrant1_p & d2fbf5;
assign a65af5 = decide_p & a65af4 | !decide_p & a662a2;
assign v12ad4d1 = hmaster2_p & v12ad4ca | !hmaster2_p & v12ad4d0;
assign v1445da3 = hlock0 & v1445d9e | !hlock0 & v1445da2;
assign f2f40e = hmaster1_p & f2f3fe | !hmaster1_p & !f2f330;
assign v15168f9 = hmaster2_p & v1668c3f | !hmaster2_p & v15168f8;
assign v1215d71 = hgrant5_p & v1215d6f | !hgrant5_p & v1215d70;
assign v14460ad = hbusreq3 & v14460ab | !hbusreq3 & v14460ac;
assign v1445a51 = hmaster1_p & v1445a50 | !hmaster1_p & v14458fd;
assign v144554d = hmaster1_p & v1445bed | !hmaster1_p & v1445544;
assign v16a205d = hbusreq2 & v16a205b | !hbusreq2 & v16a205c;
assign a64712 = decide_p & a6470f | !decide_p & a662a2;
assign v1445451 = hlock3 & v1445446 | !hlock3 & v144544f;
assign f2f3f2 = hbusreq2_p & f2f3f0 | !hbusreq2_p & f2f3f1;
assign v1215cf1 = hgrant5_p & v1215ced | !hgrant5_p & v1215cb0;
assign v14465f5 = hgrant1_p & v144641f | !hgrant1_p & v14465f4;
assign v13895a3 = hmaster1_p & v845542 | !hmaster1_p & v13895a2;
assign v1216217 = hbusreq1_p & v1216216 | !hbusreq1_p & v845542;
assign v151578e = hburst0 & v151578c | !hburst0 & v151578d;
assign v134ce6e = hbusreq5 & v134ce6c | !hbusreq5 & v134ce6d;
assign v1552fd6 = hready_p & v1553444 | !hready_p & v1552fd5;
assign v1553931 = hburst0_p & v155392f | !hburst0_p & v1553930;
assign v16a1d27 = hmaster1_p & v16a1d1f | !hmaster1_p & !v16a1f96;
assign v16a12ef = hgrant2_p & v845542 | !hgrant2_p & v16a12ee;
assign f2f426 = hbusreq5_p & f2f3a5 | !hbusreq5_p & f2f425;
assign v1216af6 = hbusreq5_p & v1216af5 | !hbusreq5_p & v845542;
assign d3061d = hmaster1_p & d3061c | !hmaster1_p & d30608;
assign d2fbb5 = hmaster0_p & d2fb7e | !hmaster0_p & d2fb85;
assign d2fc83 = hmaster0_p & v1668c17 | !hmaster0_p & v1668da6;
assign d2fb6e = hbusreq1 & d2fb6a | !hbusreq1 & d2fb6d;
assign v1445deb = hlock1 & v1445de9 | !hlock1 & v1445dea;
assign v1214d23 = hbusreq2_p & v1214d20 | !hbusreq2_p & v1214d22;
assign v1445b1a = hbusreq2_p & v1445b16 | !hbusreq2_p & v1445b19;
assign d30798 = hgrant5_p & d306d1 | !hgrant5_p & d30797;
assign v1445abb = hlock2 & v1445ab7 | !hlock2 & v1445aba;
assign v1214bc5 = hmaster1_p & v1214bc4 | !hmaster1_p & v12153a9;
assign v1668d99 = hgrant5_p & v1668d97 | !hgrant5_p & v1668d98;
assign v16a1ccd = hmaster1_p & v16a1ccc | !hmaster1_p & v16a2672;
assign v138a442 = hmaster1_p & v138a441 | !hmaster1_p & v845542;
assign v144630a = hmaster2_p & v144639c | !hmaster2_p & v144663f;
assign v14458e5 = hbusreq1_p & v1446403 | !hbusreq1_p & v14458e4;
assign d308e5 = hmaster2_p & v845542 | !hmaster2_p & d308e4;
assign v144620e = stateG10_5_p & v144620d | !stateG10_5_p & !v144620c;
assign v1284d19 = hgrant1_p & v1446427 | !hgrant1_p & v1284d18;
assign d2fb56 = hmaster1_p & d2fb52 | !hmaster1_p & d2fb55;
assign v12ad5ae = hgrant0_p & a6537d | !hgrant0_p & !v12ad4d0;
assign v1445398 = hmaster1_p & v1445a5a | !hmaster1_p & v1445a82;
assign v1214d02 = hgrant5_p & v1214c37 | !hgrant5_p & v1214d01;
assign v1214c93 = hmaster1_p & v1214c88 | !hmaster1_p & v1214c92;
assign v12aeb7b = hgrant2_p & v12aeb78 | !hgrant2_p & v12aeb73;
assign v1216ad3 = hready & v1216ad2 | !hready & !v156645f;
assign v14466e1 = hbusreq2 & v14466df | !hbusreq2 & v14466e0;
assign v1405840 = hmaster2_p & v140583d | !hmaster2_p & v140583f;
assign d2febd = hlock5_p & d2febb | !hlock5_p & d2febc;
assign v1446406 = locked_p & v845542 | !locked_p & v144639e;
assign d3065a = hlock0_p & a66295 | !hlock0_p & !v845542;
assign v134d3bb = decide_p & v134d272 | !decide_p & v134d3ba;
assign f2f430 = hgrant1_p & f2f281 | !hgrant1_p & !f2f37d;
assign v138a332 = hbusreq1_p & v138a331 | !hbusreq1_p & !v1668c63;
assign v144613a = hmaster1_p & v1446139 | !hmaster1_p & v1445fde;
assign d3027a = hgrant5_p & v845570 | !hgrant5_p & d3065e;
assign v10d4085 = hmaster1_p & v10d4084 | !hmaster1_p & !v10d407c;
assign v12ad55a = hmaster1_p & v12ad53d | !hmaster1_p & v12ad54f;
assign v1214c7a = hbusreq5_p & v1214c78 | !hbusreq5_p & v1214c79;
assign v16a142a = decide_p & v16a1429 | !decide_p & !v16a2065;
assign v1215ca7 = hgrant5_p & v1215ca0 | !hgrant5_p & v1215ca6;
assign v138a328 = hburst0 & v138a324 | !hburst0 & v138a327;
assign v144588d = hbusreq5_p & v1445886 | !hbusreq5_p & v144588c;
assign v1214f67 = hmaster0_p & v12165a8 | !hmaster0_p & v1668da6;
assign v1445878 = hbusreq5_p & v1445873 | !hbusreq5_p & v1445877;
assign v1446185 = hmaster1_p & v1446184 | !hmaster1_p & v1446073;
assign v12164d3 = hready & v12164d2 | !hready & v845542;
assign v121601a = hmaster1_p & v1216019 | !hmaster1_p & v845542;
assign v14465bc = hready & v14465bb | !hready & v144639c;
assign v1445a96 = hgrant5_p & v1445a7b | !hgrant5_p & v1445a77;
assign d2faf2 = hmaster2_p & d2f96e | !hmaster2_p & d2f976;
assign v1214dbd = hbusreq2 & v1214dba | !hbusreq2 & v1214dbc;
assign v16a1dbf = hbusreq2 & v16a1da2 | !hbusreq2 & v16a1dbe;
assign v10d42d4 = hgrant2_p & v10d40cc | !hgrant2_p & v10d42d3;
assign v12add4b = hmaster0_p & v845542 | !hmaster0_p & v12add4a;
assign v10d40b4 = hlock2_p & v10d40b1 | !hlock2_p & !v10d40b3;
assign v1552d5a = hbusreq3 & v1552d59 | !hbusreq3 & v155341e;
assign v14058a3 = hmaster2_p & v1405844 | !hmaster2_p & v140589c;
assign v144536d = hgrant2_p & v144536b | !hgrant2_p & v144536c;
assign v16a1947 = hgrant1_p & v84554d | !hgrant1_p & v16a1946;
assign v14463d5 = hbusreq3 & v14463d3 | !hbusreq3 & v14463d4;
assign f2f387 = hbusreq5_p & f2f380 | !hbusreq5_p & f2f386;
assign v1214cd5 = hmaster2_p & v1214cd4 | !hmaster2_p & v845542;
assign f2f29f = hbusreq1 & a6586b | !hbusreq1 & v845542;
assign v1215327 = hbusreq2_p & v1215322 | !hbusreq2_p & v1215326;
assign v1553412 = hbusreq1 & v155338c | !hbusreq1 & v155338d;
assign v15534ec = hbusreq1_p & v15534eb | !hbusreq1_p & v1553217;
assign v12af9b8 = decide_p & v12af9b7 | !decide_p & v845542;
assign v10d42cf = hbusreq2_p & v10d42c2 | !hbusreq2_p & !v10d42ce;
assign bf1f92 = hmaster2_p & d3064a | !hmaster2_p & bf1f91;
assign v1214d84 = hmaster1_p & v1214c96 | !hmaster1_p & v1214c92;
assign v16a1d4d = hgrant2_p & v845542 | !hgrant2_p & v16a1d4c;
assign v10d4069 = hgrant1_p & v10d4065 | !hgrant1_p & !v10d4068;
assign v1214ff7 = hgrant1_p & v1214ff1 | !hgrant1_p & v1214ff6;
assign v12acfd1 = hmaster1_p & v12acfd0 | !hmaster1_p & !v12ad525;
assign v12ad029 = hbusreq0 & v12ad028 | !hbusreq0 & !v12afa0a;
assign v121604d = hmaster2_p & v121604b | !hmaster2_p & v845542;
assign v1553224 = hgrant5_p & v845542 | !hgrant5_p & v1553223;
assign v1446292 = hmaster1_p & v1446282 | !hmaster1_p & v1446290;
assign d3063e = hlock3_p & d30632 | !hlock3_p & d3063d;
assign v134d224 = hmaster0_p & v134d221 | !hmaster0_p & v134d20a;
assign v16a13f6 = hbusreq0 & v16a13f2 | !hbusreq0 & v16a13f5;
assign v1215bde = hmaster2_p & v1216a5a | !hmaster2_p & v1215bdd;
assign v12150e0 = hmaster1_p & v12150df | !hmaster1_p & v12150d1;
assign d30153 = hlock5_p & d30151 | !hlock5_p & d30152;
assign v1215fec = hready & v1216a66 | !hready & a66295;
assign v14459af = hbusreq4 & v14459ad | !hbusreq4 & v14459ae;
assign v1445e17 = hmaster0_p & v1445de6 | !hmaster0_p & v1445e13;
assign v1216a6e = hmaster2_p & v845542 | !hmaster2_p & v1216a5a;
assign v10d426d = hgrant5_p & v10d3fdc | !hgrant5_p & v10d426c;
assign v144543d = hready_p & v144540b | !hready_p & v144543c;
assign v16a1d45 = hgrant5_p & v845542 | !hgrant5_p & v16a1d40;
assign v1284cb6 = hmaster1_p & v1284cb5 | !hmaster1_p & v1284ca7;
assign v1214c38 = hbusreq0 & v1214c37 | !hbusreq0 & v845542;
assign d2fed0 = hmaster0_p & d2feb5 | !hmaster0_p & d2fecf;
assign v146b550 = stateG2_p & v845542 | !stateG2_p & !v85e70d;
assign v1445b0b = hbusreq2 & v1445b09 | !hbusreq2 & v1445b0a;
assign v1216327 = hbusreq2_p & v121631e | !hbusreq2_p & v1216326;
assign bf1f90 = hbusreq1_p & d30649 | !hbusreq1_p & bf1f8f;
assign v1552f8a = hbusreq5 & v1552f88 | !hbusreq5 & v1552f89;
assign v14453f6 = hlock2 & v14453f5 | !hlock2 & v14453f4;
assign v12160c5 = hlock2_p & v12160c3 | !hlock2_p & v12160c4;
assign v138a2fe = hbusreq5_p & v138a2fd | !hbusreq5_p & v845542;
assign v12ad03a = hready_p & v12ad036 | !hready_p & !v12ad039;
assign v1668d0f = hbusreq2 & v1668d07 | !hbusreq2 & v1668d0e;
assign v16a1e5e = hmaster2_p & v16a1e5d | !hmaster2_p & v845542;
assign v1216147 = hlock0_p & v16a19a4 | !hlock0_p & v1216146;
assign f2f3cf = hmaster0_p & f2f3c7 | !hmaster0_p & f2f3ce;
assign v1445542 = hgrant5_p & v14465df | !hgrant5_p & v14462f0;
assign v16a1944 = hgrant0_p & v845542 | !hgrant0_p & !v16a193d;
assign v151579e = hgrant5_p & v845542 | !hgrant5_p & !v151579c;
assign d2fc8a = hlock2_p & v845542 | !hlock2_p & d2fc89;
assign v10d42c2 = hgrant2_p & v10d40b4 | !hgrant2_p & v10d42c1;
assign d2fc19 = hbusreq5 & d2fc0b | !hbusreq5 & d2fc18;
assign v1445fd0 = hmaster2_p & v1445fcf | !hmaster2_p & v1446412;
assign v16a2071 = hgrant5_p & v845542 | !hgrant5_p & v16a2070;
assign d30111 = hmaster2_p & d2fe9a | !hmaster2_p & !d300d8;
assign v1389459 = hbusreq5 & v1389430 | !hbusreq5 & v1389458;
assign d2fef1 = hbusreq2_p & d2fef0 | !hbusreq2_p & d2feef;
assign v12af9d1 = hgrant4_p & d3068f | !hgrant4_p & !v12af9d0;
assign v16a1431 = decide_p & v16a1430 | !decide_p & v16a1408;
assign a65859 = hburst0 & a65857 | !hburst0 & a65858;
assign v144590a = hmaster0_p & v14458d3 | !hmaster0_p & v1445909;
assign f2e4db = hmaster0_p & f2e4d7 | !hmaster0_p & f2e4da;
assign v1215736 = hbusreq1_p & v1215733 | !hbusreq1_p & v1215735;
assign v1445759 = hbusreq2_p & v1445757 | !hbusreq2_p & v1445758;
assign v15155f5 = hgrant2_p & v15155f4 | !hgrant2_p & !v845542;
assign v12ad00b = hmaster2_p & v12ad004 | !hmaster2_p & v12ad00a;
assign v1446143 = hbusreq2_p & v1446141 | !hbusreq2_p & v1446142;
assign v1445b5e = hlock0 & v1445b5d | !hlock0 & v1445b5c;
assign v121539d = hbusreq1_p & v121539c | !hbusreq1_p & v121539b;
assign v14459c1 = hgrant0_p & v14459bb | !hgrant0_p & v14459c0;
assign v16a140e = hmaster1_p & v16a140d | !hmaster1_p & !v16a2672;
assign v121540c = hmaster2_p & v12153d9 | !hmaster2_p & v12153dc;
assign v1446157 = hlock2 & v1446154 | !hlock2 & v1446156;
assign v11e5978 = hbusreq1_p & v11e5945 | !hbusreq1_p & v11e5977;
assign v16a12f0 = hgrant2_p & v845542 | !hgrant2_p & !v16a12ee;
assign v1445aa5 = hgrant2_p & v1445a8e | !hgrant2_p & v1445aa1;
assign v15533b1 = hmaster2_p & v155339f | !hmaster2_p & v15533b0;
assign v14453a4 = hlock5 & v1445378 | !hlock5 & v14453a3;
assign v1668dd3 = hmaster1_p & v1668dc1 | !hmaster1_p & v1668dd2;
assign v1216093 = hmaster2_p & v1216092 | !hmaster2_p & v1216067;
assign v151561e = hmaster0_p & v151561d | !hmaster0_p & v1668da6;
assign v16a1e27 = hgrant5_p & v16a2243 | !hgrant5_p & v16a1e26;
assign d308b6 = hmaster1_p & d308b5 | !hmaster1_p & d30830;
assign v1445407 = hmaster0_p & v1445406 | !hmaster0_p & v144648b;
assign v15167f3 = hmaster1_p & v15167f2 | !hmaster1_p & v845570;
assign v1215b79 = hbusreq4 & v1215fec | !hbusreq4 & v845542;
assign v1405b3f = hmaster0_p & v1405a96 | !hmaster0_p & v1405a8a;
assign v1215c62 = hgrant5_p & v16a2243 | !hgrant5_p & v1215c1b;
assign v1445de6 = hmaster2_p & v1445de5 | !hmaster2_p & v144639c;
assign v15534d5 = hbusreq1_p & v15534d4 | !hbusreq1_p & v15533a1;
assign v1445910 = hmaster0_p & v14458d3 | !hmaster0_p & v1445900;
assign d2feee = hmaster1_p & d2fed6 | !hmaster1_p & d2fee5;
assign v16a1964 = hbusreq0 & v16a209a | !hbusreq0 & v16a1963;
assign d2ff0b = hlock3_p & d2fef7 | !hlock3_p & d2ff0a;
assign a654b4 = hbusreq2_p & a654b1 | !hbusreq2_p & a654b2;
assign a654b8 = hbusreq2_p & a654b5 | !hbusreq2_p & a654b6;
assign v146af2e = stateG2_p & v845542 | !stateG2_p & v1566987;
assign v1515620 = hlock2_p & v1515617 | !hlock2_p & v151561f;
assign v10d40c3 = hgrant5_p & v10d3ffd | !hgrant5_p & !v10d40c2;
assign v140590a = hbusreq2_p & v1405907 | !hbusreq2_p & v1405909;
assign v138a2fa = hbusreq5_p & v138a2f9 | !hbusreq5_p & v845542;
assign v144672c = hmaster1_p & v144664a | !hmaster1_p & v1446630;
assign v1215c57 = hgrant5_p & v845542 | !hgrant5_p & v1215bfd;
assign v1553098 = hbusreq0 & v1553097 | !hbusreq0 & v1553395;
assign v1405aa6 = hmaster2_p & v1405a87 | !hmaster2_p & v1405aa5;
assign d30615 = hmaster1_p & d30614 | !hmaster1_p & d30608;
assign v1214c3e = hmaster1_p & v1214c3d | !hmaster1_p & v1214c39;
assign v134d265 = hmaster0_p & v134d20a | !hmaster0_p & v134d218;
assign a653bb = hgrant1_p & a653ae | !hgrant1_p & !a65387;
assign v1515730 = hgrant5_p & v10d3ff1 | !hgrant5_p & v151572e;
assign v1214c08 = hmaster1_p & v1214c07 | !hmaster1_p & v12153a9;
assign v1446281 = hlock0 & v1446280 | !hlock0 & v144643a;
assign d307db = hgrant1_p & v845542 | !hgrant1_p & d307da;
assign v144670f = hlock2 & v1446700 | !hlock2 & v144670d;
assign a65684 = hmaster1_p & a65465 | !hmaster1_p & a658e5;
assign v1445395 = hgrant2_p & v1445393 | !hgrant2_p & v1445394;
assign v1446302 = hmaster2_p & v14465ae | !hmaster2_p & v1446634;
assign v134ce64 = hgrant2_p & v134d364 | !hgrant2_p & v134ce63;
assign v1216716 = hgrant1_p & v845547 | !hgrant1_p & v1216715;
assign v14465b1 = hgrant0_p & v1446403 | !hgrant0_p & !v14463b1;
assign v16a2245 = hgrant5_p & v16a2243 | !hgrant5_p & v16a2244;
assign v14457f6 = hbusreq2_p & v14457f1 | !hbusreq2_p & v14457f5;
assign v10d3fef = locked_p & v10d3fd6 | !locked_p & v10d3fd8;
assign v1445fbf = hmaster1_p & v1445fa3 | !hmaster1_p & v1445fbd;
assign v14458eb = hbusreq1_p & v1446403 | !hbusreq1_p & v14458e2;
assign v16a1428 = hbusreq3 & v16a1425 | !hbusreq3 & v16a1427;
assign a662cd = hgrant5_p & v845542 | !hgrant5_p & a662cc;
assign v14458cb = hlock2 & v14458b3 | !hlock2 & v14458c6;
assign v15533b2 = hgrant5_p & v845542 | !hgrant5_p & v15533b1;
assign v12165ab = hmaster1_p & v12165aa | !hmaster1_p & v1216a9b;
assign v1445e66 = hlock1 & v1445e60 | !hlock1 & v1445e65;
assign v15156cd = hbusreq2 & v15156cc | !hbusreq2 & v15167ed;
assign v14454ea = hmaster2_p & v1445412 | !hmaster2_p & v144663f;
assign v1215bc5 = hlock2_p & v1215bc3 | !hlock2_p & v1215bc4;
assign bf1f99 = hgrant4_p & v845570 | !hgrant4_p & bf1f8e;
assign v12ad616 = hbusreq0 & v12ad615 | !hbusreq0 & v12afe63;
assign v1445f4d = hbusreq2_p & v1445f48 | !hbusreq2_p & v1445f4c;
assign v1515717 = stateG2_p & v845542 | !stateG2_p & a65856;
assign v1215788 = hgrant2_p & v1215787 | !hgrant2_p & v1215771;
assign d30144 = hbusreq0 & d3013e | !hbusreq0 & d30143;
assign v1216aa3 = hburst0_p & v845584 | !hburst0_p & !v845542;
assign v121656f = hgrant4_p & v845542 | !hgrant4_p & v1216a77;
assign v1445829 = hmaster1_p & v14457f7 | !hmaster1_p & v1445e28;
assign v16a1cee = hbusreq5_p & v16a1bc0 | !hbusreq5_p & v16a1ced;
assign v138a475 = hbusreq5 & v138a464 | !hbusreq5 & !v138a391;
assign v1445eda = hgrant2_p & v1445ed7 | !hgrant2_p & v1445ed9;
assign a65450 = hgrant2_p & a6540e | !hgrant2_p & !a65446;
assign v134d294 = hmaster0_p & v134d289 | !hmaster0_p & v134d293;
assign v1445fc6 = hlock3 & v1445fb2 | !hlock3 & v1445fc5;
assign v151581e = hbusreq2 & v151581d | !hbusreq2 & v15167ed;
assign v15534db = hmaster0_p & v1553395 | !hmaster0_p & v15534da;
assign v121502f = hmaster2_p & v121502a | !hmaster2_p & v121502e;
assign d2fd1b = hgrant5_p & v845570 | !hgrant5_p & d3064b;
assign d2fbd4 = hgrant4_p & d2fbce | !hgrant4_p & d2fbd3;
assign d2fbde = hlock1_p & d2fbdd | !hlock1_p & v84554a;
assign v10d42d9 = hgrant2_p & v10d40d2 | !hgrant2_p & v10d42d8;
assign v1215fb5 = hgrant2_p & v1215fb2 | !hgrant2_p & v1215fb4;
assign d2ff0d = hready_p & d2feae | !hready_p & d2ff0c;
assign v14460ec = hmaster1_p & v14460eb | !hmaster1_p & v1445f9e;
assign v1405ad9 = hmaster2_p & v1405a88 | !hmaster2_p & !v1405a8c;
assign v12ad555 = hlock2_p & v12ad553 | !hlock2_p & v12ad554;
assign v1552961 = hready_p & v1553444 | !hready_p & v1552960;
assign v16a194c = hgrant1_p & v84554d | !hgrant1_p & v16a194b;
assign v1552d9a = hmaster0_p & v1552d91 | !hmaster0_p & v845542;
assign v1214ec1 = hlock3_p & v1214eb4 | !hlock3_p & v1214ec0;
assign f2f43e = hgrant2_p & f2f3ae | !hgrant2_p & f2f419;
assign f2e501 = hready_p & f2e500 | !hready_p & f2e4f8;
assign d2fed5 = hmaster2_p & d2feb2 | !hmaster2_p & d2feb7;
assign d2fbfb = hbusreq5_p & d2fbfa | !hbusreq5_p & d2fbf9;
assign v1215c8b = hbusreq5_p & v1215c89 | !hbusreq5_p & !v1215c8a;
assign v1445fd9 = hmaster2_p & v1445fd7 | !hmaster2_p & v1445fd8;
assign d80747 = hmaster1_p & d8073b | !hmaster1_p & d80746;
assign v1552d6e = hgrant3_p & v155321c | !hgrant3_p & v1552d6d;
assign v1445fac = hbusreq2_p & v1445f9f | !hbusreq2_p & v1445fab;
assign v14463e0 = hlock4 & v14463d6 | !hlock4 & v144639e;
assign v134d4d4 = hgrant1_p & v845542 | !hgrant1_p & v134d4d3;
assign v14058ce = hbusreq4_p & v140583f | !hbusreq4_p & v14058c5;
assign v1216531 = hmaster2_p & v143fd79 | !hmaster2_p & v845542;
assign v15167bf = hbusreq5_p & v15167be | !hbusreq5_p & v845568;
assign v1405aae = hmaster0_p & v1405aa9 | !hmaster0_p & v1405aad;
assign v121573c = hbusreq1_p & v1215720 | !hbusreq1_p & v121573b;
assign v1446636 = hmaster2_p & v144639c | !hmaster2_p & v14465bb;
assign v138a3d9 = hgrant5_p & v845570 | !hgrant5_p & !v1515775;
assign d306bc = hbusreq5_p & v845542 | !hbusreq5_p & !d306a8;
assign v1445f0a = hmaster1_p & v14465b7 | !hmaster1_p & v1445f09;
assign v1215d88 = hgrant5_p & v12164d6 | !hgrant5_p & v1216700;
assign v16a2677 = hmaster1_p & v16a2676 | !hmaster1_p & !v16a2672;
assign v138932c = hgrant3_p & v13891a8 | !hgrant3_p & v1389169;
assign v12ad670 = hburst0 & v12ad66e | !hburst0 & v12ad66f;
assign v1515635 = hbusreq2_p & v1515634 | !hbusreq2_p & v845542;
assign v12afe72 = hgrant2_p & v845542 | !hgrant2_p & v12afe71;
assign d2fadd = hbusreq1 & d2f971 | !hbusreq1 & d30660;
assign a64714 = hgrant3_p & a646dc | !hgrant3_p & a64713;
assign v12ad633 = hbusreq0 & v12ad5e4 | !hbusreq0 & v12af73f;
assign v134d42c = hbusreq1_p & v134d42b | !hbusreq1_p & v134d385;
assign v1214ed8 = hmaster0_p & v1214ece | !hmaster0_p & v1214ed7;
assign v151699d = hbusreq2 & v151697c | !hbusreq2 & v151699c;
assign v12ad5df = hbusreq5_p & v12ad5dd | !hbusreq5_p & v12ad5de;
assign v12166c7 = hgrant5_p & v845542 | !hgrant5_p & v12166c6;
assign v1214f39 = hmaster1_p & v1214f38 | !hmaster1_p & v1215d3a;
assign v1405ac1 = hmaster2_p & v845542 | !hmaster2_p & v1405ac0;
assign v1214bb9 = hmaster1_p & v1214bb8 | !hmaster1_p & v12153a9;
assign v16a19c4 = hgrant2_p & v16a2060 | !hgrant2_p & v16a19c3;
assign v1215756 = hbusreq1 & v1215ba0 | !hbusreq1 & v845542;
assign d30713 = decide_p & d30712 | !decide_p & v845570;
assign d2ff01 = hbusreq2 & d2fefc | !hbusreq2 & d2ff00;
assign v16a13ed = hbusreq0 & v16a13eb | !hbusreq0 & v16a13ec;
assign f2e4d0 = hmaster0_p & f2e4cf | !hmaster0_p & f2f539;
assign f2f2ed = hmaster0_p & f2f2e3 | !hmaster0_p & f2f2cc;
assign v121603f = hbusreq1_p & v121603e | !hbusreq1_p & v845542;
assign v138945f = hmaster1_p & v138945e | !hmaster1_p & v138a006;
assign v1445858 = hmaster1_p & v1445ecc | !hmaster1_p & v1445f09;
assign v14458f0 = hlock0 & v14458ef | !hlock0 & v14458ea;
assign v15156c6 = hbusreq1_p & v1668cc4 | !hbusreq1_p & v1668cdd;
assign v12ad51b = hlock1_p & v12ad51a | !hlock1_p & v1515656;
assign v10d4040 = hbusreq4_p & v10d403f | !hbusreq4_p & !v10d402b;
assign v1214d4d = hbusreq2_p & v1214bfc | !hbusreq2_p & v1214d4c;
assign v1552f84 = hlock2 & v155341e | !hlock2 & v1552f80;
assign a662b7 = hmaster0_p & a662b2 | !hmaster0_p & a662b4;
assign f2ed95 = hbusreq5_p & f2f22b | !hbusreq5_p & f2f283;
assign v1216a62 = hmaster2_p & v1216a5a | !hmaster2_p & v1216a61;
assign v12aec08 = hbusreq0 & v12afe51 | !hbusreq0 & v12afe58;
assign v1445aea = hmaster0_p & v1445a38 | !hmaster0_p & v1445909;
assign v1214d06 = hgrant2_p & v1214ce7 | !hgrant2_p & v1214d05;
assign v12ad53d = hmaster0_p & v12ad52d | !hmaster0_p & v12ad528;
assign v1446337 = hlock2 & v144632f | !hlock2 & v1446336;
assign v16a19c7 = hgrant2_p & v16a2062 | !hgrant2_p & v16a19c6;
assign v1214db2 = hmaster1_p & v1214db1 | !hmaster1_p & v1214c39;
assign v1216008 = hbusreq1 & v1216007 | !hbusreq1 & v845542;
assign v1405908 = hmaster0_p & v14058b4 | !hmaster0_p & v1405859;
assign v1445fda = hbusreq0 & v1445fd6 | !hbusreq0 & v1445fd9;
assign d2fb42 = hmaster0_p & d2fb41 | !hmaster0_p & d2fb3b;
assign d2fc71 = hbusreq2_p & d2fc09 | !hbusreq2_p & d2fc6f;
assign v1284d2c = hmaster0_p & v1284d00 | !hmaster0_p & v1405856;
assign v16a1dd4 = hmaster1_p & v9109e4 | !hmaster1_p & !v16a1f96;
assign v16a1ae5 = hbusreq2 & v16a1ae2 | !hbusreq2 & !v16a1ae4;
assign v10d3fe0 = locked_p & v845542 | !locked_p & v10d3fdf;
assign d307f3 = hbusreq0 & d307e0 | !hbusreq0 & d307f2;
assign v1216a72 = hmaster1_p & v1216a6d | !hmaster1_p & v1216a71;
assign v12acd07 = jx0_p & v12ae83e | !jx0_p & v12acd06;
assign f2e4fa = hgrant3_p & f2e4e9 | !hgrant3_p & f2e4f9;
assign v1405881 = decide_p & v140587b | !decide_p & v1405880;
assign v12adbea = decide_p & v12adf65 | !decide_p & v12afe76;
assign a656a0 = hbusreq2_p & a6569c | !hbusreq2_p & a6569e;
assign v1214bd5 = hmaster1_p & v1214bb8 | !hmaster1_p & v1214bcf;
assign v134d53d = decide_p & v134d3e4 | !decide_p & v134d4e3;
assign d30770 = hbusreq2 & d3076b | !hbusreq2 & d3076f;
assign v1405b48 = hbusreq0_p & v1405ad3 | !hbusreq0_p & v1405b47;
assign v1216af7 = hbusreq0 & v1216ae6 | !hbusreq0 & v1216af6;
assign a654bc = hbusreq2_p & a654ba | !hbusreq2_p & a654bb;
assign v16a2059 = hmaster1_p & v9337f3 | !hmaster1_p & !v16a2672;
assign v14457d9 = hmaster1_p & v14457d8 | !hmaster1_p & v1445e07;
assign v1445493 = hmaster1_p & v1445479 | !hmaster1_p & v1446290;
assign v1216070 = hbusreq2 & v1216063 | !hbusreq2 & v121606f;
assign v15534f1 = hmaster1_p & v15534f0 | !hmaster1_p & v845542;
assign v14460d6 = hgrant2_p & v14460bd | !hgrant2_p & v14460d5;
assign v134d4f0 = hbusreq1_p & v134d273 | !hbusreq1_p & v134d36d;
assign v15530ab = hlock2 & v155321a | !hlock2 & v15530aa;
assign v12157ac = hgrant0_p & v845542 | !hgrant0_p & !v12157ab;
assign v1446427 = hbusreq4_p & v1446403 | !hbusreq4_p & v1446406;
assign v10d42db = hgrant2_p & v10d40d7 | !hgrant2_p & v10d42da;
assign v12acfb8 = hbusreq0 & v12acfb7 | !hbusreq0 & v12af9b2;
assign v1445508 = hgrant2_p & v14454e9 | !hgrant2_p & v1445507;
assign d302de = hgrant5_p & v845542 | !hgrant5_p & d30656;
assign v12ad5dd = hgrant5_p & v12ad4db | !hgrant5_p & v12ad5dc;
assign v134d448 = hlock3 & v134d3b5 | !hlock3 & v134d447;
assign v14462a5 = hready_p & v144639b | !hready_p & v14462a4;
assign v16a19cc = hbusreq5 & v16a19c0 | !hbusreq5 & v16a19cb;
assign v138a3df = hbusreq0 & v138a3db | !hbusreq0 & v138a3de;
assign v14463e3 = hlock1 & v144639c | !hlock1 & v14463e2;
assign v12166cf = hbusreq1_p & v12164d3 | !hbusreq1_p & !v12166ce;
assign v16a1a99 = hmaster1_p & v16a1a98 | !hmaster1_p & !v16a2672;
assign v12ad596 = hmaster0_p & v12ad4d2 | !hmaster0_p & v12ad4ce;
assign v1214ec8 = hgrant5_p & v1216a5a | !hgrant5_p & v121652f;
assign a66276 = hlock4_p & a66275 | !hlock4_p & !v845542;
assign bf1f75 = hmaster0_p & bf1f53 | !hmaster0_p & v84556a;
assign v155313c = hlock3_p & v155313b | !hlock3_p & v845542;
assign d30735 = hmaster2_p & d3071b | !hmaster2_p & d30734;
assign bf1f8f = hgrant4_p & a66284 | !hgrant4_p & bf1f8e;
assign v1216061 = hmaster1_p & v1216060 | !hmaster1_p & v121605d;
assign v14458e3 = hlock1 & v14458e2 | !hlock1 & v14458df;
assign d308c2 = hgrant5_p & d30654 | !hgrant5_p & d308a2;
assign v134d4b8 = hlock5 & v134d3b5 | !hlock5 & v134d4a8;
assign v1515821 = hmaster1_p & v1515820 | !hmaster1_p & v151566b;
assign d30698 = hbusreq2_p & d3063a | !hbusreq2_p & d30696;
assign d30862 = decide_p & d30861 | !decide_p & !v845570;
assign v1668c7b = hmaster2_p & v1668c6e | !hmaster2_p & !a65472;
assign d3085a = hbusreq2_p & d30849 | !hbusreq2_p & d30859;
assign v1668caa = hmaster1_p & v1668c87 | !hmaster1_p & !v1668c9c;
assign v1445a9f = hgrant2_p & v1445a85 | !hgrant2_p & v1445a9e;
assign v1553437 = hready_p & v1553427 | !hready_p & v1553436;
assign v1445e83 = hgrant5_p & v1445e7f | !hgrant5_p & v1445e82;
assign v1445d82 = hlock1 & v1445d80 | !hlock1 & v1445d81;
assign v12af73e = hgrant3_p & v12afe40 | !hgrant3_p & v12af73d;
assign d301e7 = hbusreq1 & v845542 | !hbusreq1 & !d3070c;
assign v15157d2 = hmaster1_p & v15157a5 | !hmaster1_p & v15157d1;
assign d3080f = hmaster1_p & d3080e | !hmaster1_p & v84554e;
assign v1445473 = hlock0 & v1445472 | !hlock0 & v1446654;
assign v12ad5c4 = hgrant1_p & v12ad5bd | !hgrant1_p & v12ad5c3;
assign v1515601 = hgrant2_p & v1515600 | !hgrant2_p & !v845542;
assign v1446172 = hmaster0_p & v1445fe1 | !hmaster0_p & v144639c;
assign v121537f = hmaster0_p & v121537b | !hmaster0_p & v121537e;
assign v1216ac7 = hready & v1216aaf | !hready & a66272;
assign v121500e = hbusreq0_p & v1215bad | !hbusreq0_p & !v1214fef;
assign d2fb26 = hbusreq5_p & d30147 | !hbusreq5_p & !d2fb25;
assign v1216050 = hbusreq1 & v1216ad6 | !hbusreq1 & v845542;
assign v12ad624 = hbusreq2_p & v12ad622 | !hbusreq2_p & !v12ad623;
assign v1216523 = hbusreq4 & v1216a5a | !hbusreq4 & v845542;
assign v144668c = hgrant1_p & v144668b | !hgrant1_p & v14465d1;
assign v1284cfd = hmaster0_p & v1284cf2 | !hmaster0_p & !v1284cfc;
assign v1214f5d = hbusreq2 & v1214f5c | !hbusreq2 & v12164e7;
assign d30853 = hbusreq5_p & v84554e | !hbusreq5_p & d30852;
assign v151621e = jx1_p & v1516975 | !jx1_p & v151621d;
assign v121577a = hmaster2_p & v121572a | !hmaster2_p & v1215750;
assign v1445aaa = hbusreq3 & v1445aa8 | !hbusreq3 & v1445aa9;
assign d30841 = hgrant2_p & v84554e | !hgrant2_p & d3083d;
assign v134d44c = hbusreq5_p & v134d379 | !hbusreq5_p & v134d44b;
assign v1445e00 = hmaster2_p & v1446427 | !hmaster2_p & v1445dfc;
assign v1284c95 = hbusreq2_p & v1284c92 | !hbusreq2_p & v1284c94;
assign v15530f1 = hlock5 & v155341e | !hlock5 & v15530eb;
assign v12161ed = hbusreq1_p & v12161ec | !hbusreq1_p & v845542;
assign v1445b67 = hgrant2_p & v1445b65 | !hgrant2_p & v1445b66;
assign v1445f73 = hmaster1_p & v1445f72 | !hmaster1_p & v14466a9;
assign a658c9 = hburst0 & v845542 | !hburst0 & a658c8;
assign v134d533 = hmaster0_p & v134d517 | !hmaster0_p & v845542;
assign v1446724 = hready_p & v14466cb | !hready_p & v1446723;
assign v10d3fd8 = hmastlock_p & v10d3fd6 | !hmastlock_p & v845580;
assign v1446235 = hlock0 & v1446234 | !hlock0 & v14463ec;
assign v1445e86 = hlock0 & v1445e85 | !hlock0 & v1445e78;
assign bf1f5d = hlock5_p & bf1f5b | !hlock5_p & !bf1f5c;
assign v1215b7c = hmaster2_p & v1215b76 | !hmaster2_p & v1215b7b;
assign v1215099 = hmaster2_p & v1214ffe | !hmaster2_p & v1215098;
assign a65431 = hgrant5_p & v949cd9 | !hgrant5_p & a653d1;
assign d30727 = hlock0_p & v16693aa | !hlock0_p & v845542;
assign v12164c2 = hmaster1_p & v12164c1 | !hmaster1_p & v1216af8;
assign f2e3f6 = hmaster2_p & f2f282 | !hmaster2_p & f2f228;
assign v10d4057 = hgrant5_p & v10d3ffd | !hgrant5_p & !v10d4055;
assign d306f2 = hmastlock_p & d306f1 | !hmastlock_p & !v845542;
assign v1668d3e = hgrant5_p & a65851 | !hgrant5_p & v1668d3d;
assign a658d1 = hbusreq5_p & a658cf | !hbusreq5_p & !a658d0;
assign v10d40b5 = hmaster0_p & v10d4058 | !hmaster0_p & v10d4028;
assign d2f987 = decide_p & d2f986 | !decide_p & !v845570;
assign v14058a8 = hgrant4_p & v14058a7 | !hgrant4_p & v1405849;
assign v1446732 = hmaster1_p & v1446731 | !hmaster1_p & v1446630;
assign v1214da3 = hmaster1_p & v1214ce0 | !hmaster1_p & v1214cd8;
assign v1446742 = hgrant2_p & v1446741 | !hgrant2_p & v1446732;
assign v12ad0b4 = hmaster0_p & v845542 | !hmaster0_p & v12ad0b3;
assign v140592b = hgrant4_p & v140588b | !hgrant4_p & v140592a;
assign f2f448 = hbusreq5_p & f2f3d5 | !hbusreq5_p & !f2f447;
assign d2fb80 = hmaster1_p & d2fb7f | !hmaster1_p & d2fb7b;
assign v134d45b = hbusreq5 & v134d459 | !hbusreq5 & v134d45a;
assign v1214c24 = hbusreq2 & v1214c1e | !hbusreq2 & v1214c23;
assign v1668d73 = hbusreq1 & a6586b | !hbusreq1 & v845570;
assign v1405abf = locked_p & v845542 | !locked_p & !v1405a87;
assign v1446323 = hmaster0_p & v14465b7 | !hmaster0_p & v1446322;
assign d300b6 = hbusreq1 & d2fe9a | !hbusreq1 & !v84555a;
assign d308e0 = hburst0 & d3073c | !hburst0 & d308df;
assign v1446106 = hbusreq2_p & v1446102 | !hbusreq2_p & v1446105;
assign v1215c3f = hgrant5_p & v1216029 | !hgrant5_p & !v1215c3d;
assign v144550b = hmaster1_p & v1445506 | !hmaster1_p & v1446341;
assign v12164c0 = hbusreq5 & v1216b17 | !hbusreq5 & v845542;
assign v16a1d3b = hgrant5_p & v845542 | !hgrant5_p & v16a1d3a;
assign v15530ee = hlock3 & v155341e | !hlock3 & v15530ed;
assign v14460dd = hlock3 & v14460a1 | !hlock3 & v14460dc;
assign d2fc68 = hgrant1_p & d2fbcb | !hgrant1_p & d2fc67;
assign v151697e = hmaster0_p & v845542 | !hmaster0_p & v151697d;
assign v15157e3 = hbusreq5_p & v15157e1 | !hbusreq5_p & !v15157e2;
assign v1553215 = hbusreq2_p & v1553158 | !hbusreq2_p & v1553157;
assign v1445e5b = hbusreq1 & v1445e58 | !hbusreq1 & v1445e5a;
assign v12af221 = hgrant1_p & d30690 | !hgrant1_p & v12af220;
assign v1214e0f = hmaster0_p & v1214df7 | !hmaster0_p & v1214e0e;
assign d30252 = hgrant2_p & d301cc | !hgrant2_p & d30251;
assign v134d369 = hgrant5_p & v845542 | !hgrant5_p & v134d368;
assign v1445db5 = hbusreq1 & v1445d81 | !hbusreq1 & v1445d83;
assign v1215318 = hmaster0_p & v1215bac | !hmaster0_p & v1215019;
assign d307a3 = hgrant5_p & d306fd | !hgrant5_p & !d307a1;
assign d2fc59 = hbusreq5_p & d2fbd9 | !hbusreq5_p & d2fc58;
assign v1216a8e = hmaster2_p & v845570 | !hmaster2_p & v1216a8d;
assign v16a1a30 = decide_p & v16a1a2f | !decide_p & !v16a2065;
assign v1215d7c = hmaster0_p & v1215d63 | !hmaster0_p & v12166f2;
assign v1405935 = hmaster1_p & v1405934 | !hmaster1_p & v14058d8;
assign v10d403c = hgrant5_p & v10d4038 | !hgrant5_p & v10d403b;
assign d306c9 = hbusreq1 & d306c8 | !hbusreq1 & v845542;
assign v121679a = hmaster1_p & v1216799 | !hmaster1_p & v12164e1;
assign f2f441 = hbusreq2 & f2f43d | !hbusreq2 & f2f440;
assign d3011f = hmaster0_p & d300d3 | !hmaster0_p & d3011e;
assign v1446739 = hmaster1_p & v1446738 | !hmaster1_p & v144666a;
assign v14461e7 = hbusreq2_p & v14461e1 | !hbusreq2_p & v14461e6;
assign v1552f73 = hbusreq2_p & v1552f6b | !hbusreq2_p & v1552f72;
assign v16a137d = hbusreq2 & v16a137a | !hbusreq2 & v16a137c;
assign v1215353 = hbusreq0 & v1215352 | !hbusreq0 & v845542;
assign f2f341 = decide_p & f2f340 | !decide_p & v845542;
assign v1284cae = hmaster0_p & v1284c98 | !hmaster0_p & v1284cad;
assign v138916a = hgrant3_p & v13895a6 | !hgrant3_p & v1389169;
assign a658b4 = hburst0 & a658b2 | !hburst0 & a658b3;
assign a65894 = hmaster1_p & a65891 | !hmaster1_p & a65893;
assign v12147e8 = hbusreq2_p & v12147e7 | !hbusreq2_p & v845542;
assign v14463f6 = hlock0 & v14463f5 | !hlock0 & v14463f4;
assign v1668d2d = hbusreq5_p & v1668d2a | !hbusreq5_p & v1668d2c;
assign v1405855 = hmaster2_p & v140583c | !hmaster2_p & v1405854;
assign v121502d = hgrant4_p & v845542 | !hgrant4_p & v121502c;
assign v16a1af4 = hbusreq3_p & v16a1abc | !hbusreq3_p & v16a1af3;
assign v1214c56 = hbusreq0 & v1214c55 | !hbusreq0 & v845542;
assign v1445a67 = hmaster1_p & v1445a66 | !hmaster1_p & v1445a61;
assign v1515612 = hbusreq4_p & a65851 | !hbusreq4_p & v151560d;
assign v12ad31b = hgrant4_p & d3068f | !hgrant4_p & !v12ad31a;
assign d306dc = hlock1_p & d306db | !hlock1_p & v845570;
assign v121543c = hmaster0_p & v1215439 | !hmaster0_p & v121543b;
assign v16a143d = hgrant2_p & v845542 | !hgrant2_p & v16a143c;
assign v16a1d95 = hbusreq2 & v16a1d8e | !hbusreq2 & v16a1d94;
assign v1214cda = hgrant2_p & v1214cba | !hgrant2_p & v1214cd9;
assign v1445e4e = hmaster0_p & v845542 | !hmaster0_p & v1445e4d;
assign v1215c80 = hmaster2_p & v845570 | !hmaster2_p & v1215c7e;
assign bf1f61 = hgrant5_p & v845570 | !hgrant5_p & bf1f60;
assign v134d451 = hgrant2_p & v134d364 | !hgrant2_p & v134d450;
assign v10d406f = hgrant5_p & v10d406c | !hgrant5_p & v10d406e;
assign v144632d = hmaster1_p & v144632c | !hmaster1_p & v1446329;
assign v1216066 = hlock1_p & v1216064 | !hlock1_p & !v1216065;
assign v1445f7b = hbusreq2 & v1445f79 | !hbusreq2 & v1445f7a;
assign v1446466 = hgrant5_p & v845542 | !hgrant5_p & v1446465;
assign d30673 = hbusreq5_p & d30672 | !hbusreq5_p & v845542;
assign d2fc61 = hmaster2_p & d2fc56 | !hmaster2_p & d2fc5f;
assign d30690 = hbusreq1_p & v845542 | !hbusreq1_p & d3068f;
assign v16a1e75 = hbusreq2_p & v16a1dd6 | !hbusreq2_p & v16a1e74;
assign v15167fd = hbusreq2_p & v15167fc | !hbusreq2_p & !v845542;
assign v16a1ce3 = hmaster1_p & v16a1cd0 | !hmaster1_p & !v16a1f96;
assign v16a196c = hbusreq2 & v16a196a | !hbusreq2 & !v16a196b;
assign v1668c71 = hbusreq0 & v1668c6f | !hbusreq0 & v1668c70;
assign v1446003 = hlock2 & v1445ff3 | !hlock2 & v1446001;
assign v1445a02 = hgrant1_p & v14458e8 | !hgrant1_p & v1445a01;
assign f2f408 = hmaster1_p & f2f3f5 | !hmaster1_p & !f2f330;
assign d2f9d0 = hmaster0_p & d2f9cf | !hmaster0_p & d2f9a8;
assign d3073d = stateA1_p & d3073b | !stateA1_p & v845542;
assign v1216059 = hlock1_p & v1216057 | !hlock1_p & !v1216058;
assign d3065d = hgrant1_p & f2f227 | !hgrant1_p & d3065c;
assign a653fd = hmaster2_p & a65381 | !hmaster2_p & a653bb;
assign d2f989 = hbusreq4_p & d2f988 | !hbusreq4_p & v845542;
assign v845576 = hgrant2_p & v845542 | !hgrant2_p & !v845542;
assign f2f4c2 = hbusreq3 & f2f4ba | !hbusreq3 & f2f4bf;
assign v1215092 = hgrant5_p & v1215463 | !hgrant5_p & v1215091;
assign d301de = hgrant5_p & d301c3 | !hgrant5_p & !d301d2;
assign v1215351 = hmaster2_p & v1215345 | !hmaster2_p & v121534f;
assign v16a1a89 = hgrant2_p & v845542 | !hgrant2_p & v16a1a86;
assign v1446110 = hlock2 & v14460f2 | !hlock2 & v144610e;
assign v10d4043 = hgrant1_p & v10d403e | !hgrant1_p & !v10d4042;
assign a658d8 = hmaster2_p & a6627b | !hmaster2_p & !a658d7;
assign v1445809 = hmaster1_p & v1445808 | !hmaster1_p & v1445e07;
assign v1215c98 = hbusreq5_p & v1215c96 | !hbusreq5_p & !v1215c97;
assign v12ad65a = hbusreq0 & v12ad645 | !hbusreq0 & v12af73f;
assign stateG10_5 = !v131be90;
assign v1445f88 = hmaster2_p & v1445f87 | !hmaster2_p & v14463a5;
assign v12ad328 = hbusreq0 & v12ad320 | !hbusreq0 & v12ad327;
assign v134cd5c = hgrant5_p & v134d36a | !hgrant5_p & v134cd5b;
assign v138a3ac = hbusreq2_p & v138a3a9 | !hbusreq2_p & v138a3ab;
assign v1215cc8 = hmaster0_p & v1215cb8 | !hmaster0_p & v1215cc7;
assign v1668cbc = hburst0 & v1668cba | !hburst0 & v1668cbb;
assign v1215c30 = hmaster2_p & v1215c2e | !hmaster2_p & v1215c2f;
assign f2f38a = hgrant1_p & v845570 | !hgrant1_p & !f2f389;
assign v14459f6 = hlock0_p & v144640a | !hlock0_p & v14459f5;
assign d30274 = hmaster2_p & a66295 | !hmaster2_p & v845570;
assign v1215072 = hmaster1_p & v1215065 | !hmaster1_p & v1215054;
assign v1446254 = hmaster1_p & v144639c | !hmaster1_p & v1446250;
assign d30848 = hmaster0_p & d307f7 | !hmaster0_p & d306fd;
assign d2fbb8 = hbusreq2_p & d2fbb7 | !hbusreq2_p & d2fbb2;
assign v16a1a28 = hbusreq2 & v16a1a25 | !hbusreq2 & v16a1a27;
assign bf1f7d = hmaster2_p & bf1f79 | !hmaster2_p & !bf1f7c;
assign v1445386 = hbusreq2_p & v144537b | !hbusreq2_p & v1445385;
assign v10d4297 = hgrant5_p & v10d4029 | !hgrant5_p & !v10d4296;
assign a65614 = hmaster1_p & a65613 | !hmaster1_p & a6586e;
assign v15156ec = hlock2_p & v15156ea | !hlock2_p & !v15156eb;
assign v144546d = hmaster1_p & v144546c | !hmaster1_p & v144627e;
assign v10d4266 = hmastlock_p & v10d4265 | !hmastlock_p & v10d3fd3;
assign v134cea1 = hbusreq2 & v134cea0 | !hbusreq2 & v134d240;
assign d308bd = hgrant5_p & d3085c | !hgrant5_p & d30897;
assign f2f34d = hmaster2_p & f2f347 | !hmaster2_p & f2f34c;
assign d2f993 = hmaster2_p & v84555a | !hmaster2_p & d2f992;
assign v1552d75 = hready_p & v1553427 | !hready_p & v1552d74;
assign v144581e = hmaster1_p & v14457da | !hmaster1_p & v1445ef0;
assign v15157b4 = stateG3_2_p & v845542 | !stateG3_2_p & !v1668d67;
assign v1216549 = hbusreq5_p & v1216548 | !hbusreq5_p & v845542;
assign d3073c = stateA1_p & d3073b | !stateA1_p & d306ed;
assign v1215c65 = hbusreq5_p & v1215c63 | !hbusreq5_p & v1215c64;
assign v12164cd = hbusreq5 & v12164ca | !hbusreq5 & v845542;
assign d8074f = hmaster1_p & d80748 | !hmaster1_p & d80746;
assign v1445e30 = hbusreq2 & v1445e2e | !hbusreq2 & v1445e2f;
assign v1215ccf = hbusreq5_p & v1215ccd | !hbusreq5_p & !v1215cce;
assign v1215340 = hbusreq5 & v121532e | !hbusreq5 & v121533f;
assign v12ad61a = hgrant5_p & v12ad4e4 | !hgrant5_p & v12ad5e8;
assign v1445a28 = hgrant0_p & v1445a27 | !hgrant0_p & v1445a11;
assign v12add48 = hbusreq4_p & v12add47 | !hbusreq4_p & !v84554a;
assign d2faef = hgrant5_p & d2f973 | !hgrant5_p & !d2faee;
assign v1445b07 = hmaster1_p & v1445b06 | !hmaster1_p & v14458fd;
assign v14453f2 = hmaster0_p & v144639c | !hmaster0_p & v144643b;
assign v1669594 = hbusreq3_p & v1669593 | !hbusreq3_p & !v1668c39;
assign d3019b = hmaster2_p & v16693aa | !hmaster2_p & !d30911;
assign v1405b39 = hbusreq2_p & v1405b36 | !hbusreq2_p & v1405b38;
assign v12164c9 = hbusreq2_p & v12164c8 | !hbusreq2_p & v12164c3;
assign d2fb15 = hgrant2_p & d2f984 | !hgrant2_p & d2fb11;
assign v14058e2 = hgrant2_p & v14058dd | !hgrant2_p & v14058e1;
assign d307e7 = hlock0_p & v845542 | !hlock0_p & d307e6;
assign d30293 = hmaster0_p & d30292 | !hmaster0_p & !d30282;
assign v10d4072 = hbusreq4_p & v10d4060 | !hbusreq4_p & v10d4066;
assign v1215fe9 = hbusreq1 & v1215fe8 | !hbusreq1 & v845542;
assign v1445864 = hlock3 & v14457f6 | !hlock3 & v1445862;
assign v1445e3b = hmaster2_p & v845542 | !hmaster2_p & v1445e3a;
assign v15167e9 = hmaster1_p & v15167e8 | !hmaster1_p & v845542;
assign v12afdb0 = hlock5_p & v12afdaa | !hlock5_p & v12afdaf;
assign v1216a91 = hbusreq5_p & v1216a90 | !hbusreq5_p & v845542;
assign v15157ef = hgrant5_p & v1668dc4 | !hgrant5_p & !v151575b;
assign v134d3b5 = hgrant2_p & v134d364 | !hgrant2_p & v134d3b4;
assign v12ad5ad = hbusreq4_p & v12ad5ab | !hbusreq4_p & v12ad5ac;
assign v1215c8d = hmaster2_p & v1215c8c | !hmaster2_p & v845542;
assign d306ee = stateA1_p & v1553934 | !stateA1_p & !d306ed;
assign v16a1acf = hbusreq2 & v16a1acb | !hbusreq2 & v16a1ace;
assign bf1f9e = hgrant4_p & a66284 | !hgrant4_p & bf1f9d;
assign v16a2668 = hready & v16a2667 | !hready & !v845542;
assign v1216a9f = hbusreq2_p & v1216a9c | !hbusreq2_p & v1216a9e;
assign v1668ce2 = hbusreq5_p & v1668ce0 | !hbusreq5_p & !v1668ce1;
assign v16a19b5 = hmaster0_p & v16a19b0 | !hmaster0_p & v16a19ac;
assign v1515638 = hmaster2_p & v10d3fd4 | !hmaster2_p & a653c8;
assign v138a3a7 = hmaster1_p & v138a3a6 | !hmaster1_p & v138a341;
assign v151582c = hbusreq2_p & v151582b | !hbusreq2_p & v845542;
assign v1215438 = hbusreq4_p & v1215437 | !hbusreq4_p & v845542;
assign d8079f = hmaster2_p & v845542 | !hmaster2_p & d8078a;
assign v134ce69 = hbusreq2 & v134ce67 | !hbusreq2 & v134ce68;
assign v1446179 = hmaster1_p & v144607f | !hmaster1_p & v1446099;
assign v121671a = hgrant2_p & v12164e7 | !hgrant2_p & v1216719;
assign v1668c6e = hbusreq4_p & v1668c6c | !hbusreq4_p & !v1668c6d;
assign d2fe7f = hlock4_p & v845542 | !hlock4_p & v845570;
assign v134d1fc = hbusreq1_p & v134d1fb | !hbusreq1_p & v845542;
assign v1668c35 = hready_p & v1668c27 | !hready_p & !v1668c34;
assign v144627e = hmaster0_p & v144627b | !hmaster0_p & v144627d;
assign v10d3ff7 = hbusreq4_p & v10d3fd8 | !hbusreq4_p & !v10d3fdf;
assign v155314f = hmaster1_p & v1553140 | !hmaster1_p & v155314e;
assign v14463cc = hbusreq2_p & v14463c3 | !hbusreq2_p & v14463cb;
assign d2fd3f = hbusreq2_p & d2fd14 | !hbusreq2_p & d302da;
assign d3068e = hbusreq1_p & v84555a | !hbusreq1_p & d30660;
assign v12161d6 = hgrant5_p & v12161d4 | !hgrant5_p & v12161d5;
assign v1446129 = hmaster1_p & v1446128 | !hmaster1_p & v1445fde;
assign a6470d = hgrant2_p & v845542 | !hgrant2_p & a6470c;
assign v12166dd = hgrant4_p & v12164de | !hgrant4_p & v12166dc;
assign v1445a89 = hmaster1_p & v1445a50 | !hmaster1_p & v144591b;
assign v1445b42 = hgrant2_p & v1445b3f | !hgrant2_p & v1445b41;
assign d2fcb0 = hmaster2_p & d305ea | !hmaster2_p & d2fcaf;
assign v14460ba = hmaster1_p & v1446082 | !hmaster1_p & v14460b6;
assign v1445391 = hmaster1_p & v1445361 | !hmaster1_p & v1445a82;
assign v1216156 = hgrant1_p & v845542 | !hgrant1_p & v1216155;
assign d300ea = hmaster2_p & d300e9 | !hmaster2_p & d300df;
assign v1445e50 = hgrant2_p & v1445e4f | !hgrant2_p & v1445e4b;
assign v144549a = hlock2 & v144546f | !hlock2 & v1445499;
assign d2fc52 = hgrant0_p & v84554a | !hgrant0_p & d2fc51;
assign v1445f16 = hgrant2_p & v1445efc | !hgrant2_p & v1445f12;
assign v1446215 = hbusreq0 & v1446210 | !hbusreq0 & v1446214;
assign v134d1f4 = hbusreq4_p & v134d1e8 | !hbusreq4_p & v134d1ea;
assign v12161f5 = hmaster1_p & v12161d3 | !hmaster1_p & v12161f4;
assign v121507a = hbusreq5_p & v1215079 | !hbusreq5_p & v1215040;
assign v1389f85 = hbusreq5_p & v1389f84 | !hbusreq5_p & !v845542;
assign v12ad5f6 = hgrant2_p & v12ad5f5 | !hgrant2_p & v12ad5e2;
assign v1215ff1 = hbusreq1_p & v1216521 | !hbusreq1_p & v845542;
assign v10a1543 = hgrant3_p & v10a153f | !hgrant3_p & !v10a1542;
assign v144661c = hgrant0_p & v144661a | !hgrant0_p & !v144661b;
assign v1445ae0 = hlock3 & v1445abf | !hlock3 & v1445ade;
assign v1215b88 = hmaster0_p & v1215b84 | !hmaster0_p & v1215b87;
assign v12164e0 = hbusreq5_p & v12164df | !hbusreq5_p & v845542;
assign v12acfe0 = hlock2_p & v12acfde | !hlock2_p & v12acfdf;
assign v12150bc = hmaster1_p & v12150bb | !hmaster1_p & v12153bf;
assign v1668e05 = hmaster0_p & v1668c29 | !hmaster0_p & v845542;
assign v16a1e66 = hbusreq2_p & v16a1dbe | !hbusreq2_p & v16a1e65;
assign v1515809 = decide_p & v151570c | !decide_p & !v845576;
assign v1446415 = hbusreq1_p & v1446403 | !hbusreq1_p & v1446407;
assign v1215c5f = hgrant5_p & v16a2243 | !hgrant5_p & v1215c16;
assign v1515784 = hbusreq5_p & v1515782 | !hbusreq5_p & v1515783;
assign v144614d = hbusreq2_p & v1446149 | !hbusreq2_p & v144614c;
assign v16a188d = hmaster1_p & v16a1842 | !hmaster1_p & !v16a1f96;
assign d3079f = hbusreq1_p & d3079e | !hbusreq1_p & v845542;
assign d3085f = hmaster1_p & d3085b | !hmaster1_p & d3085e;
assign v12ad580 = hmaster1_p & v12ad566 | !hmaster1_p & v12ad54f;
assign d306b1 = hmaster2_p & d306b0 | !hmaster2_p & d306a7;
assign v138a02b = hmaster2_p & d305de | !hmaster2_p & !v845570;
assign d2fae9 = hgrant1_p & d2fad8 | !hgrant1_p & d2fae8;
assign v1215d09 = hbusreq2_p & v1215d08 | !hbusreq2_p & !v1215d06;
assign v121572b = hgrant1_p & v121571a | !hgrant1_p & v845542;
assign bf1f85 = hmaster0_p & bf1f7e | !hmaster0_p & !bf1f84;
assign v1445357 = hgrant2_p & v1445356 | !hgrant2_p & v1445b41;
assign v134cd89 = hbusreq3 & v134cd87 | !hbusreq3 & v134cd88;
assign v1405b0e = hbusreq2_p & v1405b0b | !hbusreq2_p & v1405b0d;
assign v10d401d = hgrant4_p & v10d401a | !hgrant4_p & v10d401c;
assign v134d237 = hbusreq2 & v134d231 | !hbusreq2 & v134d236;
assign v1216795 = hbusreq5 & v1216794 | !hbusreq5 & v845542;
assign v12160c8 = hmaster1_p & v12160c7 | !hmaster1_p & v1216097;
assign v14459cb = hgrant4_p & v14458e2 | !hgrant4_p & v14459ca;
assign v144608f = hmaster2_p & v144603d | !hmaster2_p & v144608e;
assign v121575c = hlock4_p & v121575a | !hlock4_p & v121575b;
assign v144582d = hbusreq2 & v1445828 | !hbusreq2 & v144582c;
assign v16a1d61 = hbusreq0 & v16a1d60 | !hbusreq0 & v16a1d5e;
assign v1216120 = hbusreq4_p & v121611e | !hbusreq4_p & v121611f;
assign v14460a9 = hbusreq2_p & v1446075 | !hbusreq2_p & v14460a8;
assign v121670d = hgrant2_p & v12166f5 | !hgrant2_p & v121670c;
assign v121605b = hmaster2_p & v1216053 | !hmaster2_p & v121605a;
assign v121573b = hgrant4_p & v845542 | !hgrant4_p & v121573a;
assign d30208 = hlock1_p & d306e0 | !hlock1_p & d30207;
assign v12ad4dc = hbusreq0 & v12ad4db | !hbusreq0 & v845542;
assign v1215d9a = hbusreq5_p & v1215d99 | !hbusreq5_p & v1215d74;
assign v134ce58 = hbusreq2_p & v134ce48 | !hbusreq2_p & v134ce57;
assign v121655b = hgrant5_p & v845542 | !hgrant5_p & v121655a;
assign v1214f59 = hbusreq3 & v1214f53 | !hbusreq3 & v1214f58;
assign v1445756 = hbusreq3 & v1445754 | !hbusreq3 & v1445755;
assign v12ad66f = hburst1 & v12ad66e | !hburst1 & v1515672;
assign v144663c = hmaster1_p & v144663b | !hmaster1_p & v1446436;
assign v16a1adf = hbusreq0 & v16a1ade | !hbusreq0 & v16a208c;
assign v1216233 = hmaster0_p & v12160d5 | !hmaster0_p & v1216232;
assign v12150a5 = hbusreq0 & v1215049 | !hbusreq0 & v12150a4;
assign d2fc3c = hmaster1_p & d2fc31 | !hmaster1_p & d2fc3b;
assign v1552f69 = hmaster0_p & v1552f5c | !hmaster0_p & v1552f68;
assign v134d526 = hbusreq2 & v134d51d | !hbusreq2 & v134d525;
assign a6540f = hgrant2_p & a6540e | !hgrant2_p & !a65405;
assign v12ad669 = hbusreq3 & v12ad65d | !hbusreq3 & !v12ad668;
assign f2f396 = hmaster2_p & f2f350 | !hmaster2_p & !f2f362;
assign v11e596f = hready_p & v11e596e | !hready_p & !v845542;
assign v1284d63 = decide_p & v1284d3f | !decide_p & !v1284d62;
assign f2f29b = hmaster2_p & f2f29a | !hmaster2_p & v845542;
assign v1216225 = hmaster1_p & v1216209 | !hmaster1_p & v1216224;
assign d2fc5d = hbusreq1_p & d2fbec | !hbusreq1_p & d2fc5c;
assign v14463ee = hlock0 & v14463eb | !hlock0 & v14463ed;
assign v121658a = hgrant5_p & v845542 | !hgrant5_p & v1216589;
assign v134d523 = hgrant2_p & v134d522 | !hgrant2_p & v134d51f;
assign v1405914 = hbusreq1_p & v1405860 | !hbusreq1_p & v1405913;
assign v14058d7 = hgrant5_p & v140584c | !hgrant5_p & v14058d6;
assign v1405aec = hgrant4_p & v1405a92 | !hgrant4_p & !v1405aeb;
assign v1216320 = hlock5_p & v121631f | !hlock5_p & v12162fe;
assign v16a1328 = hgrant5_p & v845568 | !hgrant5_p & v16a1327;
assign v1445796 = hbusreq2_p & v144578d | !hbusreq2_p & v1445795;
assign v14453bb = hgrant2_p & v144539c | !hgrant2_p & v14453b7;
assign v1214c5d = hmaster2_p & v1214c51 | !hmaster2_p & v1214c5c;
assign d2fe9e = hmaster2_p & v84555a | !hmaster2_p & d2fe9d;
assign d30746 = hmaster1_p & d30745 | !hmaster1_p & d3072c;
assign v1216159 = hgrant5_p & v1216026 | !hgrant5_p & v1216157;
assign v1215715 = hbusreq4_p & v1215714 | !hbusreq4_p & v845542;
assign v14058ae = hgrant1_p & v140584b | !hgrant1_p & v14058ad;
assign v155321f = hlock2_p & v155321e | !hlock2_p & v845542;
assign a65396 = locked_p & a658c9 | !locked_p & v845542;
assign v1215ff9 = hbusreq1 & v1215ff8 | !hbusreq1 & v845542;
assign v14453a9 = hbusreq2_p & v14453a6 | !hbusreq2_p & v14453a8;
assign v16a224c = hmaster1_p & v16a224b | !hmaster1_p & !v16a2672;
assign v15530ef = hbusreq3 & v15530ed | !hbusreq3 & v15530ee;
assign v16a12e8 = hgrant0_p & v845542 | !hgrant0_p & v16a12e7;
assign d2fd3a = hbusreq2 & d2fd39 | !hbusreq2 & !v845542;
assign v1445ba8 = hready_p & v1446564 | !hready_p & v1445ba7;
assign v893df7 = stateG3_0_p & v845542 | !stateG3_0_p & v845586;
assign v1446238 = hbusreq0 & v14463f3 | !hbusreq0 & v144639c;
assign f2e884 = hgrant3_p & f2ec27 | !hgrant3_p & f2e883;
assign d30759 = hmaster1_p & d30736 | !hmaster1_p & d30754;
assign f2f2a0 = hbusreq1_p & f2f29f | !hbusreq1_p & v845542;
assign v15533a8 = hbusreq5_p & v15533a4 | !hbusreq5_p & v15533a7;
assign v10d40ad = hbusreq2_p & v10d40aa | !hbusreq2_p & v10d40ac;
assign v1284c96 = hlock3_p & v1284c95 | !hlock3_p & v140585c;
assign v134d289 = hbusreq5_p & v134d288 | !hbusreq5_p & v134d287;
assign v121606b = hmaster2_p & v1216049 | !hmaster2_p & v121601d;
assign v12162e4 = jx2_p & v1215fe7 | !jx2_p & v12162e3;
assign v144665b = hgrant1_p & v1446444 | !hgrant1_p & v144665a;
assign v845566 = hmaster1_p & v845542 | !hmaster1_p & !v845542;
assign v15168b2 = hmaster0_p & v845542 | !hmaster0_p & v15168b1;
assign v10d40ae = decide_p & v10d40a8 | !decide_p & v10d40ad;
assign d2fae0 = hgrant4_p & v845558 | !hgrant4_p & d2fadf;
assign v1214c15 = hbusreq2_p & v1214c14 | !hbusreq2_p & v1214c13;
assign v1446403 = locked_p & v845542 | !locked_p & !v14463b1;
assign v12150c3 = hlock4_p & v12150c2 | !hlock4_p & !v12153d7;
assign d306e2 = hbusreq1_p & d306e1 | !hbusreq1_p & v845542;
assign v144655a = hgrant5_p & v1446467 | !hgrant5_p & v1446559;
assign v1445a8f = hgrant2_p & v1445a8e | !hgrant2_p & v1445a8a;
assign v121539a = hbusreq1 & v1215394 | !hbusreq1 & v1215399;
assign f2f3c6 = hbusreq5_p & f2f3c4 | !hbusreq5_p & !f2f3c5;
assign v10d404e = hbusreq5_p & v10d404c | !hbusreq5_p & !v10d404d;
assign v1445802 = hlock0 & v1445801 | !hlock0 & v1445ec6;
assign v10d427d = busreq_p & v10d4264 | !busreq_p & !v10d427a;
assign a65390 = hmaster2_p & a6585d | !hmaster2_p & a65864;
assign v1446653 = hbusreq1 & v14465c1 | !hbusreq1 & v1446652;
assign v12ad4d8 = hbusreq5_p & v12ad4d6 | !hbusreq5_p & v12ad4d7;
assign d3078e = hgrant0_p & a6537d | !hgrant0_p & d3078d;
assign v1445a6b = hlock0 & v1445a6a | !hlock0 & v1445a4d;
assign v14466a6 = hgrant5_p & v1446433 | !hgrant5_p & v14466a5;
assign v134d26c = hbusreq3 & v134d26a | !hbusreq3 & v134d26b;
assign v10d408c = hgrant5_p & v10d400b | !hgrant5_p & v10d408b;
assign v12160cc = hbusreq2 & v12160c6 | !hbusreq2 & v12160cb;
assign f2e4c7 = hready_p & f2e3fd | !hready_p & f2e882;
assign v1215023 = hmaster0_p & v1215463 | !hmaster0_p & v1215462;
assign v1515606 = hready_p & v1515604 | !hready_p & !v1515605;
assign v13893b7 = hgrant3_p & v1389374 | !hgrant3_p & v13893b6;
assign v140584e = hmaster1_p & v1405842 | !hmaster1_p & v140584d;
assign v1405891 = hgrant1_p & v1405889 | !hgrant1_p & v1405890;
assign d2fb7d = hmaster2_p & d2fb69 | !hmaster2_p & v84554a;
assign v1215d3a = hmaster0_p & v1215d38 | !hmaster0_p & v1215d39;
assign v1284d0d = hmaster2_p & v1284d0c | !hmaster2_p & !v14465b3;
assign d300dc = hbusreq4_p & d300db | !hbusreq4_p & v845542;
assign v14465e3 = hgrant5_p & v14465df | !hgrant5_p & v14465e2;
assign f2ed8e = hready_p & f2f53e | !hready_p & f2ed8d;
assign f2e4e7 = hbusreq2_p & f2e4cb | !hbusreq2_p & f2f4bf;
assign a6537b = hbusreq5_p & a65379 | !hbusreq5_p & a6537a;
assign v12acfe9 = hlock2_p & v12acfe7 | !hlock2_p & v12acfe8;
assign v14465d7 = hgrant4_p & v1446406 | !hgrant4_p & v14465d6;
assign v16a1bf5 = hbusreq0 & v16a207a | !hbusreq0 & v16a1bf4;
assign v12ad54b = hlock5_p & v12ad549 | !hlock5_p & v12ad54a;
assign v12150f2 = hlock2_p & v12150f0 | !hlock2_p & v12150f1;
assign f2f43b = hmaster1_p & f2f427 | !hmaster1_p & f2f43a;
assign d3015b = hmaster1_p & d3015a | !hmaster1_p & d3014e;
assign f2f32c = hbusreq3 & f2f2ec | !hbusreq3 & f2f32b;
assign v1214d57 = hbusreq2_p & v1214c09 | !hbusreq2_p & v1214d56;
assign d306e9 = hbusreq2_p & d306e5 | !hbusreq2_p & d306e8;
assign v1215be4 = hmaster2_p & v121601c | !hmaster2_p & !v845547;
assign a65407 = hgrant2_p & a653f4 | !hgrant2_p & a65405;
assign v1668d85 = hgrant1_p & v1668d75 | !hgrant1_p & v1668d84;
assign bf1f68 = hgrant4_p & a66284 | !hgrant4_p & v845570;
assign v1445be4 = hgrant2_p & v1445be3 | !hgrant2_p & v144632a;
assign v1214dc2 = hgrant2_p & v1214dad | !hgrant2_p & v1214dc1;
assign v1405ab3 = hlock2_p & v1405aaf | !hlock2_p & v1405ab2;
assign v1668c62 = hbusreq1 & a658b5 | !hbusreq1 & !a658bd;
assign v121571c = hgrant0_p & v121571b | !hgrant0_p & v845542;
assign v16a12be = hbusreq2 & v16a129e | !hbusreq2 & v16a129f;
assign v144549d = hbusreq2 & v1445499 | !hbusreq2 & v144549a;
assign v1515721 = hgrant0_p & v1515716 | !hgrant0_p & v1515720;
assign v12160d3 = hbusreq1_p & v12160d2 | !hbusreq1_p & v845542;
assign ae2496 = hmaster0_p & v9dde65 | !hmaster0_p & v84554c;
assign a662ab = hbusreq1_p & a66289 | !hbusreq1_p & a662aa;
assign v1216287 = hgrant2_p & v1216284 | !hgrant2_p & v1216286;
assign v14466b7 = hbusreq2_p & v14466ab | !hbusreq2_p & v14466b6;
assign d30233 = hmaster1_p & d30232 | !hmaster1_p & v845542;
assign a658be = hbusreq4_p & a658bd | !hbusreq4_p & !v845542;
assign v12150ef = hmaster0_p & v12150ee | !hmaster0_p & v12150d0;
assign v121571b = hlock0_p & v1216523 | !hlock0_p & v16a19a4;
assign v12ad523 = hmaster2_p & v12ad522 | !hmaster2_p & !v12afda3;
assign v1445b7e = hgrant2_p & v1445b65 | !hgrant2_p & v1445b7d;
assign v1445e9d = hbusreq1 & v1445e9b | !hbusreq1 & v1445e9c;
assign v1445b8d = hmaster0_p & v1445b8c | !hmaster0_p & v14462fe;
assign v1668da7 = hmaster2_p & v845570 | !hmaster2_p & a6588d;
assign v12aead7 = jx2_p & v12afa35 | !jx2_p & v12aead6;
assign v151566e = busreq_p & v151566d | !busreq_p & a658a5;
assign v1215c02 = hgrant5_p & v1215bfc | !hgrant5_p & v1215c01;
assign v14466ea = hbusreq2 & v14466e8 | !hbusreq2 & v14466e9;
assign v14459a8 = hready & v14459a7 | !hready & v144639c;
assign v16a1e6d = hbusreq2 & v16a1e6a | !hbusreq2 & v16a1e6c;
assign v12ad533 = hmaster1_p & v12ad532 | !hmaster1_p & !v12ad525;
assign a662ac = hgrant1_p & v845542 | !hgrant1_p & !a662ab;
assign v1215452 = hlock2_p & v1215451 | !hlock2_p & v121544e;
assign v1215c25 = hbusreq1_p & v1215ffe | !hbusreq1_p & v1215c24;
assign v1446671 = hmaster0_p & v1446404 | !hmaster0_p & v1446638;
assign v1216580 = hgrant2_p & v121657d | !hgrant2_p & v1216576;
assign v1668dc8 = hgrant5_p & v1668dc4 | !hgrant5_p & !v1668d5e;
assign v14460c9 = hlock5 & v14460ad | !hlock5 & v14460c8;
assign v1445f8e = hgrant5_p & v14463a5 | !hgrant5_p & !v1445f8d;
assign v1553382 = hgrant4_p & v845542 | !hgrant4_p & v1553381;
assign v1214d6d = hmaster0_p & v1214d08 | !hmaster0_p & v1214c2e;
assign f2f4b2 = hlock1_p & f2f4b1 | !hlock1_p & !v845542;
assign v134d506 = hgrant0_p & v134d505 | !hgrant0_p & v845542;
assign v134d4fe = hbusreq1 & v134d4fa | !hbusreq1 & v134d4fd;
assign v16a1967 = hbusreq0 & v16a1965 | !hbusreq0 & v16a1966;
assign v1445d9e = hbusreq0 & v1445d9c | !hbusreq0 & v1445d9d;
assign v12166d6 = hbusreq4_p & v12164d3 | !hbusreq4_p & !v12166ce;
assign d30816 = hgrant5_p & v84554e | !hgrant5_p & d30797;
assign d2fc2b = hbusreq0_p & v16693aa | !hbusreq0_p & v845542;
assign v1405863 = hbusreq1_p & v1405862 | !hbusreq1_p & v14463b1;
assign v16a1db5 = hgrant2_p & v845542 | !hgrant2_p & !v16a1db2;
assign v16a13d2 = hmaster1_p & v16a13c5 | !hmaster1_p & !v16a1f96;
assign v1515708 = hbusreq2_p & v1515707 | !hbusreq2_p & v845542;
assign a653a8 = hgrant5_p & a65390 | !hgrant5_p & a653a7;
assign v134cee3 = hbusreq3 & v134cee2 | !hbusreq3 & v134d276;
assign v1668de1 = hbusreq2_p & v1668dd4 | !hbusreq2_p & v1668de0;
assign v1216ade = hlock4_p & v1216add | !hlock4_p & !v845542;
assign v1216220 = hgrant1_p & v845542 | !hgrant1_p & v121621f;
assign v151564a = stateA1_p & v845542 | !stateA1_p & v1515649;
assign v138a31e = hbusreq5 & v138a31d | !hbusreq5 & v845542;
assign v1216205 = hbusreq1 & v12166c4 | !hbusreq1 & v845547;
assign v12ad58a = hbusreq2_p & v12ad588 | !hbusreq2_p & v12ad589;
assign f2f22b = hgrant5_p & v845542 | !hgrant5_p & !f2f22a;
assign v12ad542 = hmaster1_p & v12ad541 | !hmaster1_p & !v12ad525;
assign v1446313 = hmaster0_p & v14465b7 | !hmaster0_p & v1446312;
assign v12ae83e = jx1_p & v12aead7 | !jx1_p & v12ae83d;
assign v121545b = hbusreq3 & v1215454 | !hbusreq3 & v121545a;
assign v134d384 = hgrant0_p & v134d273 | !hgrant0_p & v845542;
assign d2fc7c = decide_p & d2fc7b | !decide_p & v845570;
assign bf1fa5 = hmaster1_p & bf1f94 | !hmaster1_p & bf1fa4;
assign v10d42b8 = hgrant5_p & v10d400e | !hgrant5_p & v10d42b7;
assign v12161b3 = hbusreq2_p & v12161b0 | !hbusreq2_p & v12161b2;
assign f2f2eb = hbusreq2_p & f2f2e5 | !hbusreq2_p & f2f2ea;
assign v1215cf2 = hlock5_p & v1215cf1 | !hlock5_p & !v1215cb2;
assign v1668db5 = hbusreq5_p & v1668db3 | !hbusreq5_p & !v1668db4;
assign v144617c = hmaster0_p & v1445fe3 | !hmaster0_p & v14460a5;
assign v134d52d = hgrant3_p & v134d3fc | !hgrant3_p & v134d52c;
assign v1389f82 = jx2_p & v138a4a2 | !jx2_p & v1389efe;
assign v134d22a = hbusreq0 & v134d229 | !hbusreq0 & v134d221;
assign v1668cd6 = hmaster0_p & v1668cc9 | !hmaster0_p & v1668cd5;
assign v1216018 = hmaster2_p & v845542 | !hmaster2_p & v1216017;
assign v12ad22c = hbusreq2_p & v12ad13d | !hbusreq2_p & v12afa0e;
assign v1446631 = hmaster1_p & v14465b8 | !hmaster1_p & v1446630;
assign v16a1d5a = hbusreq0 & v16a1d58 | !hbusreq0 & v16a1d59;
assign v1552f7a = hgrant5_p & v1552f79 | !hgrant5_p & v1552f59;
assign d30951 = hlock1_p & d30950 | !hlock1_p & !v845542;
assign v1668e0d = hgrant3_p & v1668e0a | !hgrant3_p & !v1668e0c;
assign v1216240 = hmaster1_p & v121623f | !hmaster1_p & v1216224;
assign v1445e99 = hgrant0_p & v1445e98 | !hgrant0_p & !v144661b;
assign d3090c = hmaster2_p & d30718 | !hmaster2_p & !v845542;
assign d2fcd9 = hbusreq2 & d2fcb8 | !hbusreq2 & d2fcd8;
assign a662a6 = hready_p & a662a3 | !hready_p & a662a4;
assign v1215bd3 = hbusreq3 & v1215bcd | !hbusreq3 & !v845542;
assign d2fbe6 = hlock0_p & v845542 | !hlock0_p & d2fbe5;
assign f2f3db = hgrant2_p & f2f39e | !hgrant2_p & f2f3da;
assign v138a447 = hbusreq3 & v138a440 | !hbusreq3 & !v138a446;
assign v1405839 = hmastlock_p & v1405838 | !hmastlock_p & !v845542;
assign v15157dc = hbusreq5_p & v15157da | !hbusreq5_p & !v15157db;
assign v12152fe = hmaster1_p & v1214fc4 | !hmaster1_p & v1214fbf;
assign v14458dc = hlock4 & v1446407 | !hlock4 & v14458d6;
assign v1214d73 = hready_p & v1214d40 | !hready_p & v1214d72;
assign f2f359 = hmaster2_p & f2f355 | !hmaster2_p & f2f358;
assign v1405845 = hbusreq1_p & v14463b1 | !hbusreq1_p & v1405844;
assign v1445efe = hbusreq2_p & v1445ef2 | !hbusreq2_p & v1445efd;
assign f2f51a = hgrant5_p & v845542 | !hgrant5_p & !f2f519;
assign v1216595 = hbusreq1_p & v1216a8d | !hbusreq1_p & !v1216594;
assign v1668d18 = hbusreq1_p & a65851 | !hbusreq1_p & a65862;
assign v12ad512 = hburst0 & v12ad510 | !hburst0 & v12ad511;
assign v1216026 = hmaster2_p & v1216022 | !hmaster2_p & v1216025;
assign v1405ab8 = hlock2_p & v1405ab6 | !hlock2_p & v1405ab7;
assign v121612c = hgrant5_p & v121601d | !hgrant5_p & v121612a;
assign v138a39c = hlock2_p & v138a399 | !hlock2_p & v138a39b;
assign v1552d4a = hbusreq0 & v15533b2 | !hbusreq0 & v15533a4;
assign v1515655 = hbusreq1 & a658b5 | !hbusreq1 & !v1515654;
assign v14458f7 = hlock1 & v14458f6 | !hlock1 & v14458f5;
assign a65b28 = hready_p & v845542 | !hready_p & a65b27;
assign v12162c3 = hmaster1_p & v12162c2 | !hmaster1_p & v12160e0;
assign v144641c = hbusreq4_p & v1446403 | !hbusreq4_p & v144641b;
assign d30889 = hbusreq1_p & d307b5 | !hbusreq1_p & d306a5;
assign v1446135 = hmaster1_p & v1446134 | !hmaster1_p & v1445fde;
assign v1445df8 = hbusreq5_p & v1445df6 | !hbusreq5_p & v1445df7;
assign v1445e7d = hmaster2_p & v14465b3 | !hmaster2_p & v1445e7c;
assign v15156b9 = hmastlock_p & v15156b8 | !hmastlock_p & v845542;
assign v134d283 = hbusreq1_p & v134d282 | !hbusreq1_p & v845542;
assign v12acfc1 = hbusreq1_p & a658ca | !hbusreq1_p & v12ad67d;
assign v1445e7a = hbusreq1_p & v144639c | !hbusreq1_p & v1446606;
assign v134d23d = hmaster1_p & v134d1e8 | !hmaster1_p & v134d23c;
assign v12afa35 = hbusreq3_p & v12af73e | !hbusreq3_p & v12afa34;
assign v151573d = hmaster2_p & a6585c | !hmaster2_p & v151560e;
assign v1553054 = hbusreq0 & v1553053 | !hbusreq0 & v1553395;
assign d3010d = hbusreq0 & d30103 | !hbusreq0 & d3010c;
assign v138a390 = hmaster0_p & v138a38f | !hmaster0_p & !v845542;
assign v1214d3a = hbusreq3 & v1214d38 | !hbusreq3 & v1214d39;
assign v12150d1 = hmaster0_p & v12150cb | !hmaster0_p & v12150d0;
assign v1215bed = hlock2_p & v1215be3 | !hlock2_p & !v1215bec;
assign v1284caa = hmaster0_p & v1284c98 | !hmaster0_p & v1284ca9;
assign a65aee = hgrant5_p & v845542 | !hgrant5_p & a65aed;
assign d301ed = hmaster2_p & v845542 | !hmaster2_p & d301ec;
assign v14463fe = hbusreq2 & v14463fc | !hbusreq2 & v14463fd;
assign v1214d69 = hbusreq2_p & v1214c22 | !hbusreq2_p & v1214d68;
assign d2fbc7 = hmaster0_p & d2fb51 | !hmaster0_p & d2fb50;
assign v1668d62 = hbusreq1 & v1668d1c | !hbusreq1 & v845570;
assign v14465af = hgrant4_p & v14465ae | !hgrant4_p & v144639c;
assign v134d4d1 = hbusreq5_p & v134d4ce | !hbusreq5_p & v134d4d0;
assign v10d4275 = hbusreq5_p & v10d4273 | !hbusreq5_p & !v10d4274;
assign v1446105 = hmaster1_p & v14460eb | !hmaster1_p & v1445fbd;
assign v121620f = hmaster2_p & v121620e | !hmaster2_p & !v845542;
assign v1445e92 = hgrant5_p & v1445dff | !hgrant5_p & v1445e91;
assign v1446250 = hmaster0_p & v144624f | !hmaster0_p & v1446235;
assign d308a6 = hgrant1_p & v84554c | !hgrant1_p & d308a5;
assign v134d308 = hgrant2_p & v845542 | !hgrant2_p & v134d295;
assign v1284d4f = hbusreq5_p & v1284ce3 | !hbusreq5_p & v1284d4e;
assign v11e5948 = hgrant5_p & v845542 | !hgrant5_p & v11e5947;
assign a6627e = hmaster0_p & v845542 | !hmaster0_p & !a6627d;
assign v1445dc5 = hmaster1_p & v1445dc4 | !hmaster1_p & v1445dc2;
assign a65444 = hbusreq0 & a6543f | !hbusreq0 & a65443;
assign v1214d16 = hmaster1_p & v1214d15 | !hmaster1_p & v1214c39;
assign v1445a4b = hbusreq0 & v1445a4a | !hbusreq0 & v1445a36;
assign d2f9d5 = hbusreq2_p & d2f9d4 | !hbusreq2_p & d2f9d1;
assign v1445440 = hmaster1_p & v144543f | !hmaster1_p & v845542;
assign v1445898 = hlock0_p & v14463e1 | !hlock0_p & v1445897;
assign v1552d67 = hbusreq2 & v1552d65 | !hbusreq2 & v1552d66;
assign v151562f = hmastlock_p & v151562e | !hmastlock_p & v845542;
assign d30227 = hmaster2_p & d301d7 | !hmaster2_p & d301fe;
assign f2ec26 = decide_p & f2ec25 | !decide_p & v845542;
assign v1216116 = hbusreq0 & v1216104 | !hbusreq0 & v1216115;
assign v1445f91 = hlock0 & v1445f90 | !hlock0 & v1445f8c;
assign v134ce5c = hlock3 & v134d3b5 | !hlock3 & v134ce5b;
assign v1214d11 = hbusreq2_p & v1214d06 | !hbusreq2_p & v1214d10;
assign v1668dcb = hgrant5_p & v845570 | !hgrant5_p & v1668d7d;
assign a6541e = hbusreq0 & a65418 | !hbusreq0 & a6541d;
assign a65491 = hbusreq2_p & a6548d | !hbusreq2_p & a65490;
assign v1668d58 = hgrant4_p & v1668d49 | !hgrant4_p & a65382;
assign v144551e = hbusreq2_p & v144551d | !hbusreq2_p & v1445bdb;
assign v13891a6 = hbusreq5 & v138953c | !hbusreq5 & v13891a5;
assign v16a1abc = hgrant3_p & v16a2067 | !hgrant3_p & v16a1abb;
assign v1216307 = hgrant2_p & v1216304 | !hgrant2_p & v12162f8;
assign v1515602 = hbusreq2_p & v1515601 | !hbusreq2_p & !v845542;
assign a658eb = hmaster1_p & a658ea | !hmaster1_p & a658e5;
assign v1445b74 = hmaster2_p & v144665b | !hmaster2_p & v144668c;
assign d2fbcb = hbusreq1_p & d2fbca | !hbusreq1_p & v84554a;
assign a65b30 = decide_p & a65b26 | !decide_p & a662a2;
assign v12ad5b6 = hmaster2_p & v12ad4cc | !hmaster2_p & v12ad4d5;
assign d80763 = hmaster0_p & d80761 | !hmaster0_p & d80762;
assign v1405ade = hgrant5_p & v1405ad9 | !hgrant5_p & !v1405add;
assign f2f333 = hbusreq2_p & f2f331 | !hbusreq2_p & f2f332;
assign d2f9a6 = hmaster2_p & d3068e | !hmaster2_p & d2f9a5;
assign v16a1ae0 = hmaster1_p & v16a1adf | !hmaster1_p & v16a2095;
assign v1214ce3 = hgrant2_p & v1214cde | !hgrant2_p & v1214ce2;
assign v1446277 = hbusreq2 & v1446270 | !hbusreq2 & v1446276;
assign v15157f5 = hgrant5_p & v845570 | !hgrant5_p & v1515781;
assign v1215031 = hmaster2_p & v1215461 | !hmaster2_p & v1215467;
assign v12150bd = hmaster0_p & v1215019 | !hmaster0_p & v1215bac;
assign d300f6 = hbusreq0 & d300ec | !hbusreq0 & d300f5;
assign a65879 = hmaster0_p & a6585e | !hmaster0_p & a65878;
assign v144645d = hbusreq5 & v144645a | !hbusreq5 & v144645b;
assign a65469 = hmastlock_p & a65468 | !hmastlock_p & v845542;
assign v134ce3d = hlock0_p & v134d37d | !hlock0_p & v134ce3c;
assign v16a1d48 = hmaster2_p & v16a206f | !hmaster2_p & v16a1d47;
assign v12ad507 = hmaster2_p & v845542 | !hmaster2_p & v12ad506;
assign v1552d59 = hbusreq2 & v1552d57 | !hbusreq2 & v1552d58;
assign v134d399 = hlock0 & v134d38d | !hlock0 & v134d398;
assign a658ac = hburst0 & a658aa | !hburst0 & a658ab;
assign v1214c11 = hbusreq3 & v1214c04 | !hbusreq3 & v1214c10;
assign v1668d5e = hmaster2_p & v1668d5d | !hmaster2_p & v1668d5a;
assign v16a1443 = hgrant2_p & v845542 | !hgrant2_p & !v16a1442;
assign d807a2 = hgrant2_p & d807a1 | !hgrant2_p & d8079d;
assign v138a3a3 = hmaster0_p & v138a34f | !hmaster0_p & v138a344;
assign v14454f8 = hmaster1_p & v14454f7 | !hmaster1_p & v1446329;
assign v12152f6 = hmaster1_p & v12152f5 | !hmaster1_p & v121579f;
assign v151621a = hready_p & v1516218 | !hready_p & !v1516219;
assign d306ab = hmaster2_p & d306a7 | !hmaster2_p & d306aa;
assign d2fad3 = hmaster1_p & d2fad2 | !hmaster1_p & d3010e;
assign v1446399 = hmaster2_p & v845542 | !hmaster2_p & v1446398;
assign v10d40ca = hgrant2_p & v10d40b1 | !hgrant2_p & v10d40c9;
assign v121579b = hbusreq0 & v1215795 | !hbusreq0 & v121579a;
assign v16a2235 = stateG3_2_p & v845542 | !stateG3_2_p & d80753;
assign d305da = hbusreq5_p & d305d9 | !hbusreq5_p & v845542;
assign v1446646 = hmaster2_p & v14465b0 | !hmaster2_p & v1446645;
assign v1214c64 = hbusreq5_p & v1214c60 | !hbusreq5_p & v1214c63;
assign d2f9cd = hmaster1_p & d2fec8 | !hmaster1_p & d2f9cb;
assign v121611c = locked_p & v1215ff5 | !locked_p & v1215ff6;
assign v134ce93 = hbusreq2_p & v134ce92 | !hbusreq2_p & v134d23e;
assign v151560a = hmaster2_p & v1515609 | !hmaster2_p & a6585c;
assign v1214dc6 = hbusreq5 & v1214db5 | !hbusreq5 & v1214dc5;
assign v1214c86 = hbusreq2 & v1214c7f | !hbusreq2 & v1214c85;
assign v10d403f = hlock4_p & v10d3fd9 | !hlock4_p & v10d3fef;
assign v1445ea5 = hgrant1_p & v1445e04 | !hgrant1_p & v1445ea4;
assign a653e2 = hmaster2_p & a6628b | !hmaster2_p & a653e0;
assign v10d4267 = locked_p & v10d3fd4 | !locked_p & v10d4266;
assign v11e5968 = hgrant1_p & v845542 | !hgrant1_p & v11e5967;
assign v1214ce8 = hbusreq0_p & v845542 | !hbusreq0_p & v845547;
assign v12ad5c7 = hmaster2_p & v12ad5ba | !hmaster2_p & !v12ad4f7;
assign v1215bbf = hmaster2_p & v1216acd | !hmaster2_p & !v1216acf;
assign v1552d5f = hlock0 & v1552d5e | !hlock0 & v1552d5d;
assign v1216554 = hgrant4_p & v1216553 | !hgrant4_p & v121652c;
assign v1405ae7 = hgrant4_p & v1405ae6 | !hgrant4_p & !v1405a90;
assign v121611f = hbusreq4 & v121601f | !hbusreq4 & v845542;
assign v1445a09 = hlock4 & v14459a8 | !hlock4 & v14459ad;
assign v1216081 = hbusreq5_p & v1216080 | !hbusreq5_p & v121607f;
assign v134d4b5 = hbusreq2 & v134d4b3 | !hbusreq2 & v134d4b4;
assign v138a406 = hgrant2_p & v845542 | !hgrant2_p & !v84557c;
assign v1445e0f = hbusreq2_p & v1445e08 | !hbusreq2_p & v1445e0e;
assign v12161f1 = hgrant1_p & v845542 | !hgrant1_p & v12161f0;
assign v1284d5e = hmaster1_p & v1284d5d | !hmaster1_p & !v1284d1f;
assign v1214edd = hlock5_p & v1214edb | !hlock5_p & v1214edc;
assign v1446481 = hbusreq0_p & v1446480 | !hbusreq0_p & v144646e;
assign v1553220 = hgrant0_p & v845542 | !hgrant0_p & v1553138;
assign v144620d = hmaster2_p & v14463b1 | !hmaster2_p & !v14463a3;
assign v1445353 = hgrant2_p & v1445b4f | !hgrant2_p & v1445b50;
assign f2f3c1 = hmaster2_p & f2f3b1 | !hmaster2_p & !v845542;
assign v134d502 = hgrant0_p & v134d501 | !hgrant0_p & v845542;
assign d8076a = locked_p & d8073a | !locked_p & !v845542;
assign v1515836 = hbusreq5_p & v1515834 | !hbusreq5_p & v1515835;
assign v1215c6b = hmaster1_p & v1215c5a | !hmaster1_p & v1215c6a;
assign v1216ab0 = hready & v1216aaf | !hready & v1216aac;
assign v1284d03 = hmaster1_p & v1284ce5 | !hmaster1_p & !v1284cfd;
assign v1214cc3 = stateA1_p & v121658d | !stateA1_p & v1216a88;
assign v144673f = hbusreq2_p & v144673a | !hbusreq2_p & v144673e;
assign v138a001 = hlock5_p & v138a000 | !hlock5_p & !v845542;
assign v1214c25 = hbusreq3 & v1214c1a | !hbusreq3 & v1214c24;
assign bf1f8b = decide_p & bf1f4f | !decide_p & !v845570;
assign v1215bcc = hbusreq2_p & v1215bcb | !hbusreq2_p & v1215bc4;
assign d3028d = hbusreq2 & d30287 | !hbusreq2 & d3028c;
assign v151577b = hgrant1_p & v1515761 | !hgrant1_p & v151577a;
assign v138a303 = hlock5_p & v1515832 | !hlock5_p & v845570;
assign v1215d33 = hmaster2_p & v16a1bc6 | !hmaster2_p & v1216596;
assign v144662f = hlock0 & v1446618 | !hlock0 & v144662e;
assign v134cd74 = hgrant2_p & v134cd73 | !hgrant2_p & v134cd6c;
assign v1216175 = hmaster2_p & v12160f8 | !hmaster2_p & v1216126;
assign v12163a1 = hmaster2_p & v845542 | !hmaster2_p & !v1216acf;
assign f2f3a5 = hgrant5_p & f2f2a4 | !hgrant5_p & !f2f3a4;
assign v1668c58 = hbusreq3_p & v1668c57 | !hbusreq3_p & !v1668c39;
assign d3072c = hmaster0_p & d30721 | !hmaster0_p & d3072b;
assign v16a141b = hbusreq5 & v16a1412 | !hbusreq5 & v16a141a;
assign v1215fb4 = hmaster1_p & v1215fb3 | !hmaster1_p & v12166ef;
assign v16a18de = hready_p & v845555 | !hready_p & v16a18dd;
assign v1446259 = hlock2 & v1446256 | !hlock2 & v1446258;
assign d301a6 = hmaster1_p & d3090c | !hmaster1_p & !d301a5;
assign v1284c91 = hmaster0_p & v1284c90 | !hmaster0_p & v1405856;
assign v1284d15 = stateG10_5_p & v1284d13 | !stateG10_5_p & v1284d14;
assign v16a1dec = hmaster1_p & v16a1deb | !hmaster1_p & !v16a2672;
assign v14458d8 = hlock4 & v1446407 | !hlock4 & v14458d7;
assign v12ad593 = hlock3_p & v12ad563 | !hlock3_p & v12ad592;
assign v16a1d10 = hbusreq3 & v16a1b00 | !hbusreq3 & !v16a1d0f;
assign v1214c6d = hgrant4_p & v1214c6c | !hgrant4_p & v845542;
assign d301a5 = hmaster0_p & d301a4 | !hmaster0_p & !d30959;
assign v138a33f = hbusreq5_p & v138a33e | !hbusreq5_p & v845542;
assign v1216209 = hgrant5_p & v12160d5 | !hgrant5_p & v1216208;
assign v134cdc4 = hlock2 & v134d276 | !hlock2 & v134cdc3;
assign v1445f62 = hbusreq3 & v1445f60 | !hbusreq3 & v1445f61;
assign v16a139c = hready_p & v16a12f9 | !hready_p & !v16a139b;
assign v14454fb = hmaster0_p & v1446281 | !hmaster0_p & v144639c;
assign v12160f9 = hbusreq1 & v121652d | !hbusreq1 & v845542;
assign v1668d31 = hgrant5_p & v1668d15 | !hgrant5_p & v1668d30;
assign v1215724 = hgrant5_p & v1215b9a | !hgrant5_p & !v1215722;
assign v16a1b67 = hmaster1_p & v16a1b01 | !hmaster1_p & !v16a1f96;
assign v16a2092 = hgrant5_p & v845542 | !hgrant5_p & v16a2080;
assign v1214cf8 = hmaster2_p & v1214cf1 | !hmaster2_p & !v1214c31;
assign d2fb22 = hgrant5_p & d3068e | !hgrant5_p & d2fafb;
assign d301c4 = hmaster0_p & v845580 | !hmaster0_p & d301c3;
assign v1445445 = hbusreq2_p & v1445444 | !hbusreq2_p & v1445bb3;
assign v936735 = stateG3_2_p & v845542 | !stateG3_2_p & v86ab0d;
assign v1389f90 = hmaster2_p & v1515c7d | !hmaster2_p & v845542;
assign v1553144 = hmaster2_p & v845542 | !hmaster2_p & v1553142;
assign v14458d6 = locked_p & v845542 | !locked_p & v14465ad;
assign v1445812 = hbusreq2_p & v1445807 | !hbusreq2_p & v1445811;
assign v10d3fff = hmaster1_p & v10d3ffe | !hmaster1_p & v10d3ffb;
assign v12ad32a = hmaster1_p & v12af9c3 | !hmaster1_p & v12ad329;
assign v15533ac = hgrant0_p & v15533ab | !hgrant0_p & v845542;
assign v1515761 = hbusreq1_p & v151575f | !hbusreq1_p & v1515760;
assign v16695af = hbusreq3 & v16695ab | !hbusreq3 & v16695ae;
assign v14461df = hlock5 & v144619b | !hlock5 & v14461de;
assign d2fbae = hbusreq3 & d2fba5 | !hbusreq3 & d2fbad;
assign v1446199 = hlock3 & v1446181 | !hlock3 & v1446198;
assign v1215b8b = hmaster0_p & v1215b7c | !hmaster0_p & v1215b8a;
assign v134d3ad = hlock0 & v134d3ac | !hlock0 & v134d3ab;
assign d30877 = hbusreq2_p & d30773 | !hbusreq2_p & d30876;
assign v1216acd = hready & v1446394 | !hready & !v1216acc;
assign v14465c5 = hlock1 & v144639c | !hlock1 & v14465c4;
assign v1215dda = decide_p & v845542 | !decide_p & v121671a;
assign d2fba0 = hlock2_p & d2fb9e | !hlock2_p & d2fb9f;
assign d30106 = hgrant4_p & v845542 | !hgrant4_p & d30105;
assign v12153fc = hmaster1_p & v12153fb | !hmaster1_p & v12153ec;
assign v14466d2 = hmaster1_p & v14463c7 | !hmaster1_p & v14463cd;
assign v1553419 = hgrant2_p & v1553418 | !hgrant2_p & v15533b7;
assign v138938e = hbusreq0 & v138938d | !hbusreq0 & !v138a403;
assign v15157c9 = hgrant0_p & v15157c8 | !hgrant0_p & v845570;
assign v138a437 = hmaster0_p & v138a3e3 | !hmaster0_p & v138a30f;
assign v12ad4e6 = hlock0_p & v1515627 | !hlock0_p & !v12ad4e5;
assign f2e4cd = hready_p & v845542 | !hready_p & f2e4cc;
assign f2f368 = hbusreq1_p & f2f367 | !hbusreq1_p & v845542;
assign v134d509 = hbusreq1 & v134d503 | !hbusreq1 & v134d508;
assign v14459d1 = hgrant5_p & v14459a4 | !hgrant5_p & v14459d0;
assign v1216a82 = hbusreq3 & v845547 | !hbusreq3 & v1216a81;
assign v1389d5c = hmaster1_p & v845542 | !hmaster1_p & !v1389d5b;
assign v12153be = hmaster2_p & v845542 | !hmaster2_p & v12153bd;
assign d2fd4b = hgrant3_p & d2fd43 | !hgrant3_p & d2fd4a;
assign a65427 = hbusreq5_p & a65422 | !hbusreq5_p & !a65426;
assign v1214cde = hmaster1_p & v1214cdd | !hmaster1_p & v1215388;
assign v144592a = hready_p & v144639b | !hready_p & v1445929;
assign v14465c2 = hlock1 & v14465be | !hlock1 & v14465c1;
assign v144647c = hbusreq5_p & v1446473 | !hbusreq5_p & v144647b;
assign v1216576 = hmaster1_p & v121653d | !hmaster1_p & v1216575;
assign d30639 = hmaster1_p & d30638 | !hmaster1_p & d30608;
assign v15167b8 = hlock2_p & v15167b7 | !hlock2_p & v845542;
assign v1668da3 = hmaster1_p & v1668da2 | !hmaster1_p & v1668d8b;
assign v1389817 = hmaster0_p & v1389810 | !hmaster0_p & v1389816;
assign v121624f = hgrant2_p & v1216229 | !hgrant2_p & v121624e;
assign v16a1f97 = hmaster1_p & v845542 | !hmaster1_p & !v16a1f96;
assign v1515763 = hlock4_p & v1668d6e | !hlock4_p & v1515762;
assign d308e4 = hbusreq1_p & d308e3 | !hbusreq1_p & v845542;
assign v12166eb = hmaster2_p & v12166d9 | !hmaster2_p & v12166ea;
assign v1552f87 = hbusreq3 & v1552f85 | !hbusreq3 & v1552f86;
assign v10d409a = hmaster0_p & v10d4052 | !hmaster0_p & v10d3ff1;
assign v134ce9d = hmaster0_p & v134ce9c | !hmaster0_p & v134d207;
assign d2fbbe = hmaster1_p & d2fbb5 | !hmaster1_p & d2fb9d;
assign v1216297 = hmaster1_p & v1216291 | !hmaster1_p & v12161ae;
assign v1215380 = hbusreq1_p & v121537c | !hbusreq1_p & d2fbe5;
assign v1214daa = hmaster1_p & v1214da9 | !hmaster1_p & v1214d04;
assign v138a44d = hbusreq2_p & v138a44b | !hbusreq2_p & v138a44c;
assign v10d4028 = hbusreq5_p & v10d4026 | !hbusreq5_p & !v10d4027;
assign a65667 = hbusreq5_p & a6543d | !hbusreq5_p & !a65666;
assign f2f439 = hbusreq0 & f2f433 | !hbusreq0 & f2f438;
assign v1445b95 = hbusreq2_p & v1445b8f | !hbusreq2_p & v1445b94;
assign v1445be3 = hmaster1_p & v14465aa | !hmaster1_p & v1446271;
assign v1214d3e = hmaster1_p & v1214d3d | !hmaster1_p & v1215388;
assign v134d261 = hmaster1_p & v134d242 | !hmaster1_p & v134d20f;
assign v121538f = stateA1_p & v845542 | !stateA1_p & v1216aa6;
assign v14462e9 = hmaster1_p & v14462e8 | !hmaster1_p & v144627e;
assign v1515771 = hlock0_p & a6585c | !hlock0_p & v1515770;
assign v12160be = hmaster1_p & v12160a6 | !hmaster1_p & v1216082;
assign v144604a = stateG10_5_p & v1446041 | !stateG10_5_p & v1446049;
assign v151563f = hmaster2_p & v845542 | !hmaster2_p & v151563e;
assign v121651b = hmaster0_p & v1216a6c | !hmaster0_p & v1216a6a;
assign v1216a5d = stateG3_2_p & v845542 | !stateG3_2_p & v1216a5c;
assign v1214d1d = hbusreq0 & v1214d1c | !hbusreq0 & !v845542;
assign d2fc8e = hlock3_p & d2fc8d | !hlock3_p & v845552;
assign v1215314 = hmaster1_p & v1215313 | !hmaster1_p & v12153bf;
assign v1216098 = hmaster1_p & v1216093 | !hmaster1_p & v1216097;
assign v1216251 = hmaster1_p & v1216237 | !hmaster1_p & !v121624b;
assign d30784 = hlock0_p & d306c8 | !hlock0_p & !v845580;
assign v1405a95 = hmaster1_p & v1405a8b | !hmaster1_p & !v1405a94;
assign v16a1d00 = decide_p & v16a1cff | !decide_p & v16a1c04;
assign v134d270 = hbusreq2_p & v134d26f | !hbusreq2_p & v134d26e;
assign v1214bce = hbusreq0 & v1214bcd | !hbusreq0 & v845542;
assign v1445e0c = hlock0 & v1445e0b | !hlock0 & v1445e09;
assign v16a1bf8 = hgrant2_p & v845542 | !hgrant2_p & v16a1bf7;
assign v1668c42 = hmaster0_p & v1668c41 | !hmaster0_p & v1668c3f;
assign v166939f = hbusreq4_p & v1668c1c | !hbusreq4_p & !v845542;
assign v1446190 = hgrant2_p & v144618e | !hgrant2_p & v144618f;
assign v1445af0 = hmaster0_p & v1445a36 | !hmaster0_p & v1445900;
assign d2fd2d = hbusreq2_p & d2fd2c | !hbusreq2_p & d302e5;
assign v138a3c4 = hmaster1_p & v138a3c3 | !hmaster1_p & v138a301;
assign v16a1e2a = hgrant2_p & v16a1d2e | !hgrant2_p & v16a1e29;
assign v1216275 = hmaster0_p & v12161f7 | !hmaster0_p & f2f2a8;
assign v1216131 = hgrant1_p & v845542 | !hgrant1_p & v1216130;
assign v1215791 = hmaster2_p & v1215b97 | !hmaster2_p & v845542;
assign d300fc = hbusreq4_p & d300fb | !hbusreq4_p & v845542;
assign v11e597a = hmaster2_p & v11e5979 | !hmaster2_p & v845542;
assign v12afe47 = hgrant5_p & v845542 | !hgrant5_p & v12afe46;
assign d30678 = hbusreq2_p & d30677 | !hbusreq2_p & d30670;
assign v138a3a8 = hmaster1_p & v138a34f | !hmaster1_p & v138a341;
assign v15161d3 = hlock2_p & v15161d2 | !hlock2_p & !v845542;
assign v121679e = hbusreq5 & v121679d | !hbusreq5 & v12164e7;
assign v15530b1 = decide_p & v155342e | !decide_p & v15530b0;
assign v1216245 = hbusreq2_p & v1216244 | !hbusreq2_p & v1216241;
assign v1445bd7 = hgrant2_p & v1445bcc | !hgrant2_p & v1445bd6;
assign f2f3a6 = hgrant5_p & f2f3a1 | !hgrant5_p & !f2f3a4;
assign v12166f0 = hmaster1_p & v12166c8 | !hmaster1_p & v12166ef;
assign d2f98f = hlock5_p & d2f98d | !hlock5_p & d2f98e;
assign d307d8 = hbusreq1 & d307d7 | !hbusreq1 & v845542;
assign v1214bf1 = hbusreq0 & v1214bb7 | !hbusreq0 & v845542;
assign a6567f = hbusreq2_p & a6567d | !hbusreq2_p & !a6567e;
assign v12ad01e = hgrant2_p & v12ad01d | !hgrant2_p & !v12ad018;
assign v144666f = hmaster1_p & v14465b8 | !hmaster1_p & v144666a;
assign f2f3ba = hbusreq5_p & f2f3b8 | !hbusreq5_p & !f2f3b9;
assign v1405b50 = hgrant5_p & v1405a96 | !hgrant5_p & v1405b4f;
assign v16a13e8 = hgrant2_p & v845542 | !hgrant2_p & v16a13e7;
assign v1215bf3 = hgrant5_p & v1215bda | !hgrant5_p & v1215bf2;
assign v134d429 = hgrant5_p & v845542 | !hgrant5_p & v134d428;
assign v1389fca = hbusreq3 & v1389fc4 | !hbusreq3 & v138a391;
assign a6569a = hbusreq3 & a6568d | !hbusreq3 & a65699;
assign v144648b = hgrant5_p & v845542 | !hgrant5_p & v144648a;
assign v1214d85 = hgrant2_p & v1214d37 | !hgrant2_p & v1214d84;
assign a65ae0 = hready_p & a65adc | !hready_p & a65add;
assign v1445aed = hlock2 & v1445ae9 | !hlock2 & v1445aec;
assign v134d4e1 = hmaster1_p & v134d4e0 | !hmaster1_p & v845542;
assign v121578e = hbusreq0 & v121578c | !hbusreq0 & v121578d;
assign v1215333 = hbusreq2_p & v1215330 | !hbusreq2_p & v1215332;
assign d2fb0b = hgrant1_p & d2fb00 | !hgrant1_p & d2fb0a;
assign v1516213 = decide_p & v151699e | !decide_p & !v845576;
assign v1668d11 = hbusreq5 & v1668cf7 | !hbusreq5 & v1668d10;
assign v155338f = hbusreq1_p & v1553217 | !hbusreq1_p & v155338e;
assign v144537e = hgrant2_p & v144537c | !hgrant2_p & v144537d;
assign v14458b5 = hbusreq2 & v14458ae | !hbusreq2 & v14458b4;
assign v1446329 = hmaster0_p & v14462f3 | !hmaster0_p & v1446616;
assign v15161fd = hbusreq2_p & v15161fc | !hbusreq2_p & !v845542;
assign v12af9d8 = hmaster1_p & v12af9c3 | !hmaster1_p & v12af9d7;
assign v1216174 = hmaster1_p & v1216173 | !hmaster1_p & !v1216027;
assign v1445363 = hgrant2_p & v1445360 | !hgrant2_p & v1445362;
assign v1215745 = hbusreq1 & v121611f | !hbusreq1 & v845542;
assign v121570b = hlock2_p & v1215708 | !hlock2_p & !v121570a;
assign v1445de5 = hbusreq4_p & v14465ae | !hbusreq4_p & v144639c;
assign v12aeb1e = hmaster0_p & v845542 | !hmaster0_p & v12aeb1d;
assign v12162cd = hbusreq2 & v12162c6 | !hbusreq2 & v12162cc;
assign v16a1b6b = hbusreq5 & v16a1b63 | !hbusreq5 & v16a1b6a;
assign v16a12c4 = hmaster1_p & v16a1a97 | !hmaster1_p & v16a1f96;
assign v1214e70 = hmaster2_p & v1214e6f | !hmaster2_p & v1214df3;
assign v144599c = hbusreq1 & v1445999 | !hbusreq1 & v144599b;
assign v11e5973 = hbusreq0_p & v11e593a | !hbusreq0_p & v845570;
assign f2f356 = hbusreq1 & v1668d3b | !hbusreq1 & v845542;
assign v15156e7 = hlock2_p & v15156db | !hlock2_p & !v15156e6;
assign v1445b8e = hmaster1_p & v14465b7 | !hmaster1_p & v1445b8d;
assign v1389393 = hbusreq5 & v1389380 | !hbusreq5 & v1389392;
assign v10d405a = hmaster1_p & v10d4059 | !hmaster1_p & !v10d404f;
assign v12ad579 = hmaster1_p & v12ad531 | !hmaster1_p & !v12ad525;
assign v12ad52f = hmaster1_p & v12ad52e | !hmaster1_p & !v12ad525;
assign v10d40a2 = hmaster1_p & v10d40a1 | !hmaster1_p & v10d3fe9;
assign v10d4030 = hgrant4_p & v10d402d | !hgrant4_p & v10d402f;
assign v121622f = hbusreq2_p & v1216226 | !hbusreq2_p & v121622e;
assign v1215d69 = hmaster1_p & v1215d64 | !hmaster1_p & v1215d68;
assign v144606f = hmaster2_p & v144605a | !hmaster2_p & v144606e;
assign d30285 = hgrant2_p & d30267 | !hgrant2_p & d30284;
assign v1445f52 = hgrant2_p & v144674c | !hgrant2_p & v144674e;
assign v1445f02 = hbusreq3 & v1445f00 | !hbusreq3 & v1445f01;
assign v14454a6 = hbusreq5 & v14454a3 | !hbusreq5 & v14454a4;
assign v1284d67 = jx2_p & v85e755 | !jx2_p & v1284d66;
assign v15530e9 = hbusreq2 & v15530e8 | !hbusreq2 & v155341e;
assign v1216079 = hmaster1_p & v1216078 | !hmaster1_p & v121605d;
assign v144640d = hlock1 & v144640a | !hlock1 & v144640c;
assign a6542e = hbusreq0 & a65427 | !hbusreq0 & a6542d;
assign d30952 = hbusreq1_p & d30951 | !hbusreq1_p & !v845542;
assign v1215360 = hbusreq0 & v121535f | !hbusreq0 & v845542;
assign v1552f5b = hbusreq0 & v1552f5a | !hbusreq0 & v1553395;
assign v14465cd = hgrant0_p & v1446407 | !hgrant0_p & v144639c;
assign v1215cba = hgrant1_p & v1215cb9 | !hgrant1_p & v121613f;
assign d3069b = hbusreq5_p & v845542 | !hbusreq5_p & !d3068c;
assign v1445b88 = hlock5 & v144634e | !hlock5 & v1445b87;
assign v1445ef9 = hgrant2_p & v1445ef7 | !hgrant2_p & v1445ef8;
assign d80799 = hgrant1_p & v845542 | !hgrant1_p & d80798;
assign v1668dab = hmaster2_p & v845542 | !hmaster2_p & a65396;
assign v12ae76b = hready_p & v12ae6fe | !hready_p & v12ae76a;
assign v1215d8b = hgrant2_p & v1215d86 | !hgrant2_p & v1215d8a;
assign v1445ee1 = hmaster1_p & v1445ee0 | !hmaster1_p & v1445e07;
assign v12ad5e7 = hmaster1_p & v12ad5e6 | !hmaster1_p & v12ad4ff;
assign v14058e6 = hmaster1_p & v14058e5 | !hmaster1_p & !v1446403;
assign a6561a = hmaster0_p & a653f9 | !hmaster0_p & a653ea;
assign v1445b60 = hmaster1_p & v14465b7 | !hmaster1_p & v1445b5f;
assign v10d4098 = hready_p & v10d4088 | !hready_p & !v10d4097;
assign v16a1d6f = hmaster1_p & v16a1d6e | !hmaster1_p & v16a1d6d;
assign v16a1413 = hgrant2_p & v16a1d31 | !hgrant2_p & v16a1d98;
assign v1405acc = hmaster1_p & v1405acb | !hmaster1_p & !v1405ac8;
assign v121608f = hbusreq2_p & v121608e | !hbusreq2_p & v121608d;
assign f2f3b7 = hbusreq2 & f2f3ac | !hbusreq2 & f2f3b6;
assign v134d1e7 = stateG2_p & v845542 | !stateG2_p & v134d1e6;
assign v16a19c0 = hbusreq3 & v16a19b4 | !hbusreq3 & v16a19bf;
assign d300e2 = hgrant5_p & d2fe9e | !hgrant5_p & d300e0;
assign v1215c69 = hbusreq0 & v1215c67 | !hbusreq0 & v1215c68;
assign d2fb2a = hmaster0_p & d2fb24 | !hmaster0_p & d2fb29;
assign v1445af1 = hmaster1_p & v1445af0 | !hmaster1_p & v144590e;
assign v12166d7 = hbusreq4_p & v1216586 | !hbusreq4_p & v12166c3;
assign v121627f = hready_p & v1216278 | !hready_p & !v121627e;
assign v1445916 = hbusreq3 & v1445914 | !hbusreq3 & v1445915;
assign d306f9 = hmaster0_p & d306d3 | !hmaster0_p & d306d0;
assign v1668d30 = hmaster2_p & v1668d2f | !hmaster2_p & v845542;
assign v138a3f2 = hmaster1_p & v138a3f1 | !hmaster1_p & v1668c23;
assign v14458b7 = hbusreq3 & v14458b5 | !hbusreq3 & v14458b6;
assign v134d4ca = locked_p & v134d4c9 | !locked_p & v845542;
assign v134d536 = hbusreq2 & v134d532 | !hbusreq2 & v134d535;
assign a65873 = hmaster1_p & a6585f | !hmaster1_p & a6586e;
assign v1445f66 = hmaster1_p & v14466af | !hmaster1_p & v14466a9;
assign v11e5983 = hbusreq3_p & v11e5970 | !hbusreq3_p & v11e5982;
assign d30867 = hbusreq1_p & d30722 | !hbusreq1_p & d30660;
assign f2f23d = decide_p & f2f23a | !decide_p & f2f23c;
assign v134d4f8 = hlock0 & v134d4f7 | !hlock0 & v134d4ef;
assign v1214e7e = hbusreq2 & v1214e7d | !hbusreq2 & v845542;
assign v1215ff0 = hmaster2_p & v1215fea | !hmaster2_p & v1215fef;
assign v1214cec = hgrant1_p & v1214c29 | !hgrant1_p & v1214ceb;
assign d30188 = hgrant2_p & d3095b | !hgrant2_p & d3091a;
assign v14459b3 = hlock4 & v144639c | !hlock4 & v14459a7;
assign f2f3b0 = hbusreq1 & a65396 | !hbusreq1 & !v845542;
assign v1405925 = stateG2_p & v845542 | !stateG2_p & !v1405853;
assign v12157a6 = hmaster1_p & v12157a5 | !hmaster1_p & v121579f;
assign v121629f = hbusreq2_p & v1216298 | !hbusreq2_p & v121629e;
assign a65898 = decide_p & a65896 | !decide_p & v845542;
assign v14466bb = hlock2 & v14466b7 | !hlock2 & v14466ba;
assign d2fba7 = hmaster1_p & d2fb8f | !hmaster1_p & d2fb9d;
assign v12ad003 = hbusreq1_p & v12ad5c2 | !hbusreq1_p & v12ad002;
assign v1216197 = hbusreq5_p & v1216195 | !hbusreq5_p & v1216196;
assign v1445d91 = stateG10_5_p & v1445d90 | !stateG10_5_p & !v1445d8f;
assign v1214818 = decide_p & v1214ec0 | !decide_p & v1214817;
assign v845556 = hlock3_p & v845542 | !hlock3_p & !v845542;
assign v121614c = hgrant4_p & v1216148 | !hgrant4_p & v121614b;
assign v14453fa = hbusreq2_p & v1446291 | !hbusreq2_p & v14453f3;
assign v138a404 = hgrant2_p & v845542 | !hgrant2_p & !v138a403;
assign v1405b41 = hlock2_p & v1405b3e | !hlock2_p & v1405b40;
assign v16a1cf5 = hbusreq2 & v16a1cf2 | !hbusreq2 & !v16a1cf4;
assign v1445427 = hbusreq3 & v1445425 | !hbusreq3 & v1445426;
assign v12ae1ef = hbusreq4_p & v12afe4d | !hbusreq4_p & v12afe44;
assign v1446201 = hlock5 & v144617b | !hlock5 & v1446200;
assign v1389fc4 = hbusreq2_p & v1389fbb | !hbusreq2_p & v1389fc3;
assign v12ae200 = hmaster1_p & v12afe47 | !hmaster1_p & v12ae1ff;
assign v1445782 = hmaster0_p & v1445776 | !hmaster0_p & v1445de7;
assign a6628e = hbusreq5_p & a66287 | !hbusreq5_p & a6628c;
assign v1445535 = hbusreq3 & v1445533 | !hbusreq3 & v1445534;
assign f2f292 = hbusreq1 & a65851 | !hbusreq1 & v845542;
assign v16a13e3 = hgrant5_p & v845542 | !hgrant5_p & v16a13e2;
assign v14459fa = hbusreq1 & v14459f9 | !hbusreq1 & v14459cc;
assign v1668ca2 = hmaster1_p & v1668c75 | !hmaster1_p & !v1668ca1;
assign v121508d = hgrant1_p & v121545f | !hgrant1_p & v121508c;
assign v16a139e = hbusreq3_p & v16a1382 | !hbusreq3_p & v16a139d;
assign v134d468 = hready_p & v134d3be | !hready_p & v134d467;
assign v12162f7 = hmaster0_p & v12162e8 | !hmaster0_p & v12162f6;
assign v134cd63 = hgrant4_p & v845542 | !hgrant4_p & v134cd62;
assign d305fe = hmaster2_p & v84555a | !hmaster2_p & v845542;
assign v16a1cd2 = hmaster1_p & v16a1cd1 | !hmaster1_p & v16a2672;
assign d2fead = hlock3_p & d2fe99 | !hlock3_p & !d2feac;
assign v1445554 = hgrant3_p & v1445541 | !hgrant3_p & v1445553;
assign v144609f = hmaster1_p & v144609e | !hmaster1_p & v1446099;
assign v138944c = hlock5_p & v138944b | !hlock5_p & v845542;
assign v12acfc6 = hmaster1_p & v12acfc5 | !hmaster1_p & !v12acfb9;
assign v1445a4e = hbusreq0 & v1445a4a | !hbusreq0 & v1445a4d;
assign a6543e = hgrant5_p & v845558 | !hgrant5_p & !a653f5;
assign v1214f7d = decide_p & v1214ec0 | !decide_p & v1214f71;
assign v1445517 = hmaster1_p & v14454f0 | !hmaster1_p & v1445b7a;
assign v845572 = hgrant0_p & v845542 | !hgrant0_p & !v845542;
assign v138a325 = busreq_p & v138a322 | !busreq_p & !v845542;
assign d301f3 = hbusreq1_p & d301f2 | !hbusreq1_p & v1668d52;
assign v15157cc = hmaster2_p & v15157c7 | !hmaster2_p & v15157cb;
assign f2f41a = hgrant2_p & f2f417 | !hgrant2_p & f2f419;
assign v10a153f = hready_p & v845542 | !hready_p & v845564;
assign v1216535 = hgrant4_p & v1216524 | !hgrant4_p & v1216534;
assign v1553513 = hbusreq3 & v1553512 | !hbusreq3 & v155321a;
assign d2fec1 = hmaster2_p & v84555a | !hmaster2_p & d2fec0;
assign v12ad0ca = hbusreq2 & v12ad0bd | !hbusreq2 & v12afe3d;
assign v1553436 = decide_p & v155342e | !decide_p & v1553435;
assign v1214d78 = hmaster1_p & v1214d77 | !hmaster1_p & v1214c74;
assign v1445dfe = hbusreq1 & v1445dfb | !hbusreq1 & v1445dfd;
assign v1389fbb = hmaster1_p & v845542 | !hmaster1_p & v1389fba;
assign v1552d60 = hmaster0_p & v1552d5f | !hmaster0_p & v1552d4b;
assign v144583e = hbusreq2 & v1445839 | !hbusreq2 & v144583d;
assign v1284d28 = decide_p & v1284cb8 | !decide_p & !v1284d27;
assign v12161a3 = hmaster1_p & v12161a2 | !hmaster1_p & v121619c;
assign v14457da = hmaster0_p & v1445eba | !hmaster0_p & v14465b7;
assign d2fe98 = hmaster1_p & d2fe95 | !hmaster1_p & d2fe97;
assign v1515746 = hbusreq4_p & v1515744 | !hbusreq4_p & !v1515745;
assign v121541b = hbusreq2_p & v121541a | !hbusreq2_p & v1215419;
assign d2fd22 = hlock5_p & d2fd20 | !hlock5_p & !d2fd21;
assign v121603a = hmaster2_p & v1216037 | !hmaster2_p & v845542;
assign d30708 = hmaster2_p & d306fc | !hmaster2_p & !d306fe;
assign d30839 = hlock5_p & d30837 | !hlock5_p & d30838;
assign v1445a71 = hbusreq2 & v1445a5f | !hbusreq2 & v1445a70;
assign v10d400d = hmaster1_p & v10d400c | !hmaster1_p & !v10d3fe9;
assign v1445eb0 = hlock0 & v1445eaf | !hlock0 & v1445ead;
assign v12152f1 = hgrant2_p & v1215787 | !hgrant2_p & v12152ea;
assign v1445fca = hbusreq5 & v1445fc8 | !hbusreq5 & v1445fc9;
assign d30818 = hbusreq5_p & d30817 | !hbusreq5_p & d30816;
assign v138a335 = hgrant4_p & v138a334 | !hgrant4_p & v1668cc4;
assign v1215c35 = hmaster0_p & v1215c23 | !hmaster0_p & v1215c34;
assign v1216003 = hbusreq0_p & v1216a5a | !hbusreq0_p & v1215ff8;
assign f2f414 = decide_p & f2f413 | !decide_p & v845542;
assign v1405877 = hmaster1_p & v1405876 | !hmaster1_p & v140586f;
assign v1445ee6 = hlock3 & v1445edb | !hlock3 & v1445ee5;
assign v12166ca = locked_p & v12166c9 | !locked_p & v845542;
assign f2f42c = hgrant5_p & f2f363 | !hgrant5_p & f2f42b;
assign v1214f0e = hbusreq0 & v121655b | !hbusreq0 & v121656e;
assign d307df = hlock5_p & d307dd | !hlock5_p & d307de;
assign d30131 = hlock5_p & d3012f | !hlock5_p & d30130;
assign v1446115 = hlock5 & v1446101 | !hlock5 & v1446114;
assign v1405b02 = hgrant4_p & v1405a88 | !hgrant4_p & !v1405a90;
assign d30623 = hmaster1_p & d30622 | !hmaster1_p & d30608;
assign v1216185 = hmaster0_p & v845542 | !hmaster0_p & v1216184;
assign v121532a = hmaster0_p & v121505b | !hmaster0_p & v1215065;
assign v1552d79 = hbusreq3_p & v1552d6e | !hbusreq3_p & v1552d78;
assign v16a1bd8 = hgrant5_p & v845542 | !hgrant5_p & v16a1bd7;
assign v14460b8 = hgrant2_p & v14460ae | !hgrant2_p & v14460b7;
assign f2e4d8 = hmaster2_p & f2f228 | !hmaster2_p & f2f282;
assign v1552f7d = hlock0 & v1552f7c | !hlock0 & v1552f7b;
assign v12aee5e = hgrant3_p & v12aed9f | !hgrant3_p & v12aee5d;
assign d30870 = hmaster1_p & d30865 | !hmaster1_p & d3086f;
assign v1446063 = hbusreq1_p & v1446600 | !hbusreq1_p & v144660e;
assign d3084c = hmaster2_p & d3084a | !hmaster2_p & !d3084b;
assign d807b9 = hmaster0_p & d807ae | !hmaster0_p & d80762;
assign v15530f4 = hready_p & v1553306 | !hready_p & v15530f3;
assign f2f460 = hgrant3_p & f2f415 | !hgrant3_p & f2f45f;
assign a658f0 = hmaster1_p & a658ef | !hmaster1_p & a658e5;
assign d3087e = hmaster1_p & d3087d | !hmaster1_p & d306e4;
assign v1405b26 = hgrant1_p & v1405ac6 | !hgrant1_p & v1405b25;
assign v16a1a8e = decide_p & v16a1a2f | !decide_p & !v16a19cc;
assign a65b0a = hmaster1_p & a66287 | !hmaster1_p & a65b09;
assign v1214da8 = hmaster1_p & v1214da7 | !hmaster1_p & v1214c39;
assign v15167ea = hlock2_p & v15167e9 | !hlock2_p & v845542;
assign v1446746 = hmaster0_p & v1446448 | !hmaster0_p & v144639c;
assign v144544b = hbusreq2 & v1445445 | !hbusreq2 & v144544a;
assign v1552d86 = hgrant1_p & v845542 | !hgrant1_p & v1552d85;
assign v1668cc4 = hmastlock_p & v1668cc3 | !hmastlock_p & v845542;
assign v16a132b = hgrant2_p & v16a2058 | !hgrant2_p & v16a132a;
assign a65b06 = decide_p & a65aff | !decide_p & v845542;
assign v1445422 = hgrant2_p & v1445420 | !hgrant2_p & v1445421;
assign v12adf66 = decide_p & v12adf65 | !decide_p & v845542;
assign v16a1bfd = hgrant5_p & v845542 | !hgrant5_p & !v16a1bf3;
assign v1445f6c = hbusreq2_p & v1445f65 | !hbusreq2_p & v1445f6b;
assign v14459fd = hmaster2_p & v14465b3 | !hmaster2_p & v14459fc;
assign v1668d1c = hbusreq4_p & a65851 | !hbusreq4_p & a65862;
assign d305f6 = hlock5_p & v845542 | !hlock5_p & d305f5;
assign v14459ab = hbusreq0_p & v14459aa | !hbusreq0_p & v14465bb;
assign v1215474 = hbusreq2_p & v1215470 | !hbusreq2_p & v1215473;
assign v134ce89 = hlock1 & v134d1e8 | !hlock1 & v134d1ec;
assign v16a1c95 = hbusreq1 & v845547 | !hbusreq1 & v845542;
assign v134cd68 = hgrant5_p & v845542 | !hgrant5_p & v134cd67;
assign v1445e07 = hmaster0_p & v1445dfa | !hmaster0_p & v1445e06;
assign v10d4293 = hgrant4_p & v10d3fe0 | !hgrant4_p & v10d4292;
assign a653b7 = hbusreq5_p & a653a8 | !hbusreq5_p & !a653b6;
assign v12153c1 = hmaster0_p & v1215baf | !hmaster0_p & v1215bac;
assign d2fada = hgrant4_p & v845558 | !hgrant4_p & d2fad9;
assign v12ad58f = hbusreq2_p & v12ad58d | !hbusreq2_p & v12ad58e;
assign v1446093 = hmaster0_p & v144603f | !hmaster0_p & v1446092;
assign v1668cda = stateA1_p & v1566987 | !stateA1_p & v1668cc0;
assign a65b3d = hbusreq3_p & a65b3c | !hbusreq3_p & a65b32;
assign v121626b = hready_p & v1216200 | !hready_p & v121626a;
assign v10d3ff0 = hmaster2_p & v10d3fd4 | !hmaster2_p & v10d3fef;
assign f2f37a = hbusreq1_p & f2f379 | !hbusreq1_p & v845542;
assign v16a2249 = hgrant2_p & v16a2059 | !hgrant2_p & v16a2248;
assign v16a1be6 = hgrant5_p & v845542 | !hgrant5_p & !v16a1bcb;
assign a65ad6 = hgrant5_p & v845542 | !hgrant5_p & a662d2;
assign v1284cbb = hmaster1_p & v1284cba | !hmaster1_p & !v1445bb7;
assign v121575b = hlock0_p & v1215b79 | !hlock0_p & !v845542;
assign d3064c = hlock5_p & v845542 | !hlock5_p & d3064b;
assign v16a209a = hgrant5_p & v845542 | !hgrant5_p & !v16a206f;
assign v1446054 = hbusreq0 & v144604c | !hbusreq0 & v1446053;
assign d3070f = hmaster0_p & d3070e | !hmaster0_p & v84554e;
assign v134d3c5 = hbusreq2_p & v134d245 | !hbusreq2_p & v134d3c4;
assign v12ad662 = hmaster0_p & v12ad660 | !hmaster0_p & v12ad661;
assign v1215ba3 = hmaster2_p & v12160ec | !hmaster2_p & !v121611f;
assign v134d461 = hlock2 & v134d276 | !hlock2 & v134d460;
assign d80738 = decide_p & d80737 | !decide_p & d80736;
assign d302d6 = hmaster1_p & v845542 | !hmaster1_p & d302d5;
assign v1553424 = decide_p & v1553216 | !decide_p & v1553423;
assign v1668cc7 = hmaster2_p & v1668cbd | !hmaster2_p & v1668cc6;
assign v16a1bee = hbusreq1 & v16a207f | !hbusreq1 & v16a2089;
assign v15156b4 = hbusreq2_p & v15156b3 | !hbusreq2_p & v845542;
assign v1446124 = hmaster1_p & v1446123 | !hmaster1_p & v1445fef;
assign d306ff = hbusreq5_p & v84554e | !hbusreq5_p & d306fe;
assign v138a3d0 = hlock5_p & v138a3cd | !hlock5_p & !v138a3cf;
assign v12153e6 = hlock0_p & v12153d6 | !hlock0_p & v845547;
assign v12afe68 = hgrant2_p & v845542 | !hgrant2_p & v12afe67;
assign v10d407d = hmaster1_p & v10d4064 | !hmaster1_p & !v10d407c;
assign v155322f = hbusreq4_p & v155322e | !hbusreq4_p & v845542;
assign d3094d = hburst1 & a658a5 | !hburst1 & d3094c;
assign v1668c22 = hbusreq5_p & v1668c21 | !hbusreq5_p & v845542;
assign d3062c = hbusreq5_p & v845542 | !hbusreq5_p & d305fe;
assign v16a132a = hmaster1_p & v16a1329 | !hmaster1_p & !v16a2672;
assign v1215c21 = hgrant5_p & v1215c12 | !hgrant5_p & v1215c20;
assign v1214c83 = hgrant2_p & v1214c82 | !hgrant2_p & v1214c75;
assign v144580d = hbusreq2_p & v1445807 | !hbusreq2_p & v144580c;
assign v1284cee = hmaster2_p & v1284ce9 | !hmaster2_p & !v1405845;
assign v131be90 = hgrant3_p & v131be8c | !hgrant3_p & v131be8f;
assign v121546f = hmaster0_p & v121546a | !hmaster0_p & v121546e;
assign d301e4 = hbusreq0 & d301e0 | !hbusreq0 & d301e3;
assign v1668cea = hmaster1_p & v1668cd9 | !hmaster1_p & v1668cd6;
assign f2e733 = hmaster1_p & f2f229 | !hmaster1_p & f2e732;
assign f2ed9f = hbusreq3_p & f2ed8f | !hbusreq3_p & f2ed9e;
assign d301ca = hmaster0_p & d301c8 | !hmaster0_p & d301c9;
assign v1215c4a = hmaster2_p & v845542 | !hmaster2_p & v1216568;
assign v1215044 = hgrant0_p & v1215043 | !hgrant0_p & !v845542;
assign d30724 = hlock1_p & v845542 | !hlock1_p & d305fb;
assign v16693a8 = hmaster0_p & v16693a7 | !hmaster0_p & v845542;
assign v1445527 = hlock3 & v144551b | !hlock3 & v1445524;
assign v155342a = hbusreq1_p & v1553140 | !hbusreq1_p & v1553429;
assign v121536c = hmaster1_p & v1215365 | !hmaster1_p & v121536b;
assign v1446268 = hbusreq0 & v14465ea | !hbusreq0 & v144642c;
assign a653c9 = hbusreq0_p & a653c8 | !hbusreq0_p & !a65394;
assign v151583e = hlock2_p & v151583d | !hlock2_p & v15157d2;
assign d30809 = hlock1_p & v845542 | !hlock1_p & !v1668c1c;
assign v1668c9d = hmaster1_p & v1668c61 | !hmaster1_p & !v1668c9c;
assign v140593e = hready_p & v140593c | !hready_p & v140593d;
assign v14461b2 = hgrant2_p & v14461b0 | !hgrant2_p & v14461b1;
assign v16695a3 = hlock3_p & v16695a2 | !hlock3_p & v845542;
assign d2fcff = hmaster1_p & d2fcac | !hmaster1_p & d2fcfe;
assign a6591c = hmaster1_p & a658ef | !hmaster1_p & !a65916;
assign v1446676 = hbusreq2_p & v1446670 | !hbusreq2_p & v1446675;
assign v15156f7 = hlock2_p & v15156f3 | !hlock2_p & !v15156f6;
assign d308ad = hmaster0_p & d3089d | !hmaster0_p & d308ac;
assign d2fcf3 = hbusreq2 & d2fcec | !hbusreq2 & d2fcd8;
assign v134ce83 = hmaster2_p & v134d1e8 | !hmaster2_p & v134ce82;
assign v1515787 = hmaster1_p & v151573c | !hmaster1_p & v1515786;
assign a65b2c = hgrant2_p & v845542 | !hgrant2_p & a65b2b;
assign v1445468 = hbusreq5 & v144545e | !hbusreq5 & v144545f;
assign d30837 = hgrant5_p & d306d0 | !hgrant5_p & d307ff;
assign v134d3cf = hbusreq5 & v134d3cc | !hbusreq5 & v134d3ce;
assign v16a1bcc = hmaster2_p & v16a1bc5 | !hmaster2_p & v16a1bcb;
assign a653a1 = hgrant4_p & v845570 | !hgrant4_p & !a65863;
assign d3086d = hbusreq5_p & d3072a | !hbusreq5_p & d3086c;
assign v12150c6 = hlock1_p & v12150c5 | !hlock1_p & v1215b97;
assign v1214fc9 = hbusreq2 & v12157a8 | !hbusreq2 & v1214fc8;
assign v15155e4 = hgrant3_p & v1515c88 | !hgrant3_p & !v1515baf;
assign v1446602 = hbusreq1 & v14465fa | !hbusreq1 & v1446601;
assign d301fd = hlock5_p & d301fb | !hlock5_p & d301fc;
assign d2fbeb = hgrant0_p & v845542 | !hgrant0_p & d2fbe6;
assign a64705 = hbusreq2 & a64704 | !hbusreq2 & a65b29;
assign v1446055 = hlock0 & v1446054 | !hlock0 & v144604c;
assign v12162d1 = hgrant2_p & v12162c3 | !hgrant2_p & v12162d0;
assign v1405b07 = hmaster2_p & v1405b03 | !hmaster2_p & v1405b06;
assign v1552fcd = hlock2 & v155321a | !hlock2 & v1552fcc;
assign v1445e10 = hbusreq1 & v1445dea | !hbusreq1 & v1445ded;
assign v10d4284 = hgrant4_p & v10d3fd5 | !hgrant4_p & v10d4283;
assign d2fc46 = hbusreq5 & d2fc3f | !hbusreq5 & d2fc45;
assign v1446001 = hbusreq2_p & v1445ffd | !hbusreq2_p & v1446000;
assign v12afda8 = hbusreq4_p & v12afda6 | !hbusreq4_p & v12afda7;
assign v1445bb3 = hmaster1_p & v14463c5 | !hmaster1_p & v1445bb1;
assign v1215c2f = hgrant1_p & v1215c28 | !hgrant1_p & v1216162;
assign v10d429d = hgrant4_p & v10d4071 | !hgrant4_p & !v10d429c;
assign v1445ec8 = hgrant1_p & v1445e10 | !hgrant1_p & v1445ec7;
assign f2f2d2 = hbusreq1 & v1668c6e | !hbusreq1 & v845542;
assign v15530fd = hmaster0_p & v1552d52 | !hmaster0_p & v845542;
assign d30626 = hbusreq2 & d30621 | !hbusreq2 & d30625;
assign v1214f08 = hbusreq5_p & v1214f07 | !hbusreq5_p & v1214f06;
assign v1215cd7 = hgrant2_p & v845542 | !hgrant2_p & !v1215cd6;
assign v1668d98 = hmaster2_p & v1668d28 | !hmaster2_p & v1668d54;
assign v1405b2e = hmaster0_p & v1405b16 | !hmaster0_p & v1405b2d;
assign v138a066 = hmaster2_p & v84556a | !hmaster2_p & !v845542;
assign v1445f68 = hbusreq2_p & v1445f65 | !hbusreq2_p & v1445f67;
assign v138a34e = hmaster2_p & v138a32b | !hmaster2_p & a658dc;
assign v14466c9 = hmaster0_p & v14464a6 | !hmaster0_p & v845542;
assign v140586f = hmaster0_p & v140586a | !hmaster0_p & v140586e;
assign d30631 = hmaster1_p & v845542 | !hmaster1_p & d30630;
assign v1216542 = hmaster2_p & v845542 | !hmaster2_p & v1216541;
assign v16a1cfa = hgrant2_p & v845542 | !hgrant2_p & !v16a1cf9;
assign v14462fa = hbusreq0 & v14462f8 | !hbusreq0 & v14462f9;
assign d2fb97 = hbusreq2 & d2fb92 | !hbusreq2 & d2fb96;
assign v12153d3 = hbusreq4_p & v12153d2 | !hbusreq4_p & v845542;
assign v1216279 = hmaster0_p & v1216227 | !hmaster0_p & v12160d5;
assign v1214ccb = hmaster2_p & v1214cbe | !hmaster2_p & v1214cca;
assign v15157f0 = hbusreq5_p & v15157ee | !hbusreq5_p & !v15157ef;
assign v1445996 = hbusreq4 & v1445994 | !hbusreq4 & v1445995;
assign v1214fef = hbusreq4 & v1216594 | !hbusreq4 & !v845542;
assign v1668c78 = hmaster2_p & a658b5 | !hmaster2_p & v1668c77;
assign v14460a0 = hgrant2_p & v144609d | !hgrant2_p & v144609f;
assign v1215012 = hgrant4_p & v845542 | !hgrant4_p & v1215011;
assign v12ad5f4 = hmaster1_p & v12ad5f3 | !hmaster1_p & v845542;
assign d30766 = hbusreq5 & d30750 | !hbusreq5 & d30765;
assign v1214fbb = hgrant1_p & v1215757 | !hgrant1_p & v1214fba;
assign v1445dcd = hgrant5_p & v1445dcb | !hgrant5_p & !v1445dcc;
assign v16a1e0e = hbusreq5 & v16a1e09 | !hbusreq5 & v16a1e0d;
assign v1668c5b = decide_p & v1668c5a | !decide_p & v845542;
assign v1446219 = hmaster0_p & v1446216 | !hmaster0_p & v1446218;
assign v15157d9 = hbusreq5_p & v15157d7 | !hbusreq5_p & !v15157d8;
assign d2fc75 = hmaster0_p & d2fc74 | !hmaster0_p & d2fc6c;
assign v1215c12 = hmaster2_p & v121611d | !hmaster2_p & v1215be6;
assign v16a13dd = hgrant5_p & v845542 | !hgrant5_p & v16a13dc;
assign v12ae1ff = hmaster0_p & v12afe47 | !hmaster0_p & v12ae1fe;
assign a65852 = hbusreq4_p & a65851 | !hbusreq4_p & v845542;
assign v121619a = hgrant5_p & v845542 | !hgrant5_p & v121616a;
assign v1214bc8 = hbusreq2 & v1214bc2 | !hbusreq2 & v1214bc7;
assign d2fb9e = hmaster1_p & d2fb6c | !hmaster1_p & d2fb9d;
assign v155339b = hgrant4_p & v155339a | !hgrant4_p & v845542;
assign v1214ed4 = hgrant5_p & v1214dcc | !hgrant5_p & v1214ed3;
assign v10d4077 = hgrant0_p & v10d4076 | !hgrant0_p & v10d3ff9;
assign v1214d52 = hmaster1_p & v1214d51 | !hmaster1_p & v1214d4b;
assign v16a1ad0 = hmaster0_p & v845542 | !hmaster0_p & !v16a1ac9;
assign v12af5a9 = hbusreq1_p & v12af5a8 | !hbusreq1_p & v12afe61;
assign v16a2068 = stateA1_p & v845542 | !stateA1_p & !v845582;
assign v1445ad6 = hbusreq2 & v1445ad4 | !hbusreq2 & v1445ad5;
assign f2f296 = hmaster2_p & f2f293 | !hmaster2_p & f2f295;
assign v12aeb76 = hbusreq0 & v12afda2 | !hbusreq0 & v12aeb75;
assign f2f224 = decide_p & f2f223 | !decide_p & v845542;
assign v1446040 = hmaster2_p & v144639c | !hmaster2_p & v1446412;
assign d2feda = hlock2_p & d2fed7 | !hlock2_p & d2fed9;
assign v12ad5eb = hbusreq5_p & v12ad5e9 | !hbusreq5_p & v12ad5ea;
assign v14058fa = hgrant1_p & v1446403 | !hgrant1_p & !v14058f9;
assign v1405919 = decide_p & v1405918 | !decide_p & v1405880;
assign v1405af1 = hmaster1_p & v1405ad8 | !hmaster1_p & v1405af0;
assign d30775 = hmaster1_p & d3076c | !hmaster1_p & d30754;
assign v134d46d = jx2_p & v134d3e9 | !jx2_p & v134d46c;
assign v134d4e6 = hbusreq4 & v134d273 | !hbusreq4 & v134d4e5;
assign v14838bf = hgrant3_p & v14838b9 | !hgrant3_p & v14838be;
assign v1445e29 = hmaster1_p & v1445de8 | !hmaster1_p & v1445e28;
assign v12150ad = hgrant2_p & v1215059 | !hgrant2_p & v12150ac;
assign v1215775 = hmaster1_p & v1215774 | !hmaster1_p & !v1215ba1;
assign v14457d6 = hbusreq0 & v1445eb3 | !hbusreq0 & v1445eb6;
assign v12acfff = hlock0_p & v151560d | !hlock0_p & d2fc50;
assign v1215c3c = hmaster2_p & v1215fe8 | !hmaster2_p & v1215ff8;
assign v16a1847 = hmaster1_p & v16a1846 | !hmaster1_p & v16a2672;
assign v121503c = hgrant5_p & v1215031 | !hgrant5_p & v121503b;
assign d3076c = hmaster0_p & d3072e | !hmaster0_p & d30735;
assign a6566f = hbusreq5_p & a65429 | !hbusreq5_p & !a6566e;
assign v1445bf3 = decide_p & v1446224 | !decide_p & v1445bf2;
assign v1215bab = hlock3_p & v1215b96 | !hlock3_p & !v1215baa;
assign v134d30c = hgrant5_p & v134d281 | !hgrant5_p & v134d30b;
assign v16a19a7 = hgrant0_p & v845542 | !hgrant0_p & !v16a19a6;
assign v11ac602 = hgrant1_p & v845542 | !hgrant1_p & v84554c;
assign v1445838 = hbusreq2_p & v1445830 | !hbusreq2_p & v1445837;
assign d30765 = hbusreq3 & d3075c | !hbusreq3 & d30764;
assign v144674e = hmaster1_p & v144674d | !hmaster1_p & v1446630;
assign v12ad54d = hbusreq5_p & v12ad54b | !hbusreq5_p & v12ad54c;
assign v15157c4 = hgrant5_p & v845542 | !hgrant5_p & !v15157c2;
assign d2fb07 = hbusreq5_p & d30102 | !hbusreq5_p & !d2fb06;
assign v12af5a8 = hlock1_p & v12af5a4 | !hlock1_p & v12af5a7;
assign v14466f6 = hmaster1_p & v14466f5 | !hmaster1_p & v1446436;
assign v12166d0 = hbusreq1 & v1216587 | !hbusreq1 & v845570;
assign v1389463 = hbusreq2_p & v1389462 | !hbusreq2_p & v138a404;
assign v1214e58 = hgrant1_p & v1214e57 | !hgrant1_p & v1216ab8;
assign v14460e2 = hready_p & v1446038 | !hready_p & v14460e1;
assign v9337f3 = hmaster0_p & v845568 | !hmaster0_p & v845542;
assign v12161db = hmaster2_p & v12161da | !hmaster2_p & v845542;
assign v121615a = hbusreq5_p & v1216158 | !hbusreq5_p & v1216159;
assign d807ac = hmaster1_p & d807ab | !hmaster1_p & d8079c;
assign v121653b = hlock5_p & v121653a | !hlock5_p & v1216531;
assign v16a1d9c = hbusreq2 & v16a1d99 | !hbusreq2 & v16a1d9b;
assign v15532bf = hbusreq2_p & v155323a | !hbusreq2_p & v15532be;
assign d8078f = hmaster2_p & d8078a | !hmaster2_p & v845542;
assign v1405b4f = hmaster2_p & v1405b4e | !hmaster2_p & v1405a87;
assign v138a32f = hgrant4_p & v138a32e | !hgrant4_p & v1515654;
assign v1216afc = hmaster0_p & v1216ab3 | !hmaster0_p & v1216afb;
assign v10d42bb = hgrant2_p & v10d4090 | !hgrant2_p & v10d42ba;
assign v12153ee = hmaster2_p & v12153ce | !hmaster2_p & v1215b97;
assign d2fcb7 = hlock2_p & v845542 | !hlock2_p & !d2fcb6;
assign v155343c = hbusreq1_p & v1553221 | !hbusreq1_p & v155343b;
assign v140588f = hgrant0_p & v140588c | !hgrant0_p & !v140588e;
assign bf1f55 = hmaster1_p & bf1f54 | !hmaster1_p & !bf1f52;
assign v138a322 = stateG2_p & v845542 | !stateG2_p & !v138a321;
assign v12153dd = hmaster2_p & v12153d3 | !hmaster2_p & v12153dc;
assign v1553448 = hbusreq3_p & v1553426 | !hbusreq3_p & v1553447;
assign d2fedd = hmaster1_p & d2fedc | !hmaster1_p & d2fec6;
assign v14465db = hgrant1_p & v14465d9 | !hgrant1_p & v14465da;
assign v16a1888 = hbusreq3 & v16a1845 | !hbusreq3 & v16a1887;
assign d30910 = hlock1_p & d3090f | !hlock1_p & !v845542;
assign d807bf = hgrant3_p & d807bc | !hgrant3_p & d807be;
assign v16a1bc0 = hgrant5_p & v845542 | !hgrant5_p & v16a1bbf;
assign v140583a = busreq_p & v845588 | !busreq_p & !v146d169;
assign v1668ccf = hbusreq4 & v1668cbd | !hbusreq4 & v1668cce;
assign v14461ed = hmaster1_p & v1446184 | !hmaster1_p & v14460cf;
assign v1284cd7 = hgrant4_p & v1284cd6 | !hgrant4_p & !v1405849;
assign v10d4015 = hmaster1_p & v10d4014 | !hmaster1_p & v10d3fe9;
assign v1388ce9 = jx0_p & v138a0c7 | !jx0_p & v1388ce8;
assign v1668c4c = hmaster1_p & v1668c4b | !hmaster1_p & v845542;
assign v1445fcb = hmaster2_p & v1446403 | !hmaster2_p & v1446412;
assign d80743 = hbusreq4_p & d80742 | !hbusreq4_p & !v845542;
assign d80755 = stateG3_2_p & v845542 | !stateG3_2_p & d80754;
assign v16a1a90 = hgrant3_p & v16a1a31 | !hgrant3_p & v16a1a8f;
assign v12acff1 = hmaster0_p & v12ad4e0 | !hmaster0_p & v12ad4ce;
assign v1214c31 = hbusreq1_p & d2fbe5 | !hbusreq1_p & v1214c30;
assign v1445854 = hgrant2_p & v144582e | !hgrant2_p & v1445853;
assign v1515748 = hbusreq1_p & v1668d35 | !hbusreq1_p & v1515747;
assign f2f2a6 = hmaster1_p & f2f2a5 | !hmaster1_p & f2f2a2;
assign v12164d7 = hbusreq5_p & v12164d6 | !hbusreq5_p & v16a2243;
assign v12162bc = decide_p & v12162a1 | !decide_p & v12162bb;
assign v1668dc3 = hgrant5_p & v1668dc2 | !hgrant5_p & v1668d4d;
assign v121653a = hgrant5_p & v845542 | !hgrant5_p & v1216539;
assign v1553391 = hmaster2_p & v845542 | !hmaster2_p & v1553390;
assign v134ce5f = hgrant5_p & v134ce5e | !hgrant5_p & v134ce39;
assign d8074b = hlock2_p & d80747 | !hlock2_p & d8074a;
assign d3013f = hgrant5_p & d30138 | !hgrant5_p & d300ee;
assign v16a223d = hgrant1_p & v845542 | !hgrant1_p & v16a223c;
assign v1215b83 = hmaster2_p & v1215b80 | !hmaster2_p & v1215b81;
assign v16a1dd9 = hbusreq3 & v16a1dd5 | !hbusreq3 & v16a1dd8;
assign v12aecdb = hready_p & v12aec4f | !hready_p & v12aecda;
assign a65626 = hbusreq5_p & a653f8 | !hbusreq5_p & a65625;
assign v1445e59 = hbusreq4_p & v14465c4 | !hbusreq4_p & v14465bb;
assign d2fc37 = hbusreq1_p & v845542 | !hbusreq1_p & v845558;
assign v1216b05 = hmaster1_p & v1216b04 | !hmaster1_p & v1216af8;
assign v1284d0e = hgrant5_p & v140587e | !hgrant5_p & v1284d0d;
assign v12afe75 = hgrant5_p & v845542 | !hgrant5_p & v12afe74;
assign v1216038 = hmaster2_p & f2f2a8 | !hmaster2_p & v1216037;
assign a6546f = hmaster2_p & a658b6 | !hmaster2_p & a6546d;
assign v131be8b = decide_p & v131be8a | !decide_p & v84555c;
assign a662a1 = hgrant5_p & v845542 | !hgrant5_p & a662a0;
assign v138a3fc = hbusreq2 & v138a3f0 | !hbusreq2 & v138a3fb;
assign v121545a = hbusreq2 & v1215450 | !hbusreq2 & v1215459;
assign v15168af = hlock1_p & v15168ae | !hlock1_p & v16693aa;
assign v12ad951 = hbusreq2_p & v12add4c | !hbusreq2_p & v12ad8ed;
assign v12166c4 = hgrant4_p & v12164cf | !hgrant4_p & v12166c3;
assign v1214d0d = hbusreq0 & v1214d0c | !hbusreq0 & v16a2243;
assign v16a208e = hmaster2_p & v16a208a | !hmaster2_p & v16a2080;
assign v1215c07 = hmaster2_p & v1216a61 | !hmaster2_p & v1215bdd;
assign v1515bae = decide_p & v1516105 | !decide_p & !v845576;
assign f2f4ac = hmaster1_p & v845542 | !hmaster1_p & f2f4ab;
assign v16a1ab7 = hbusreq2 & v16a224d | !hbusreq2 & v16a224f;
assign v1216284 = hlock2_p & v1216281 | !hlock2_p & !v1216283;
assign v1445a3e = hgrant5_p & v1445900 | !hgrant5_p & v1445a3d;
assign v1216b10 = hmaster1_p & v1216b0f | !hmaster1_p & v1216af8;
assign v12ad4e1 = hmaster0_p & v12ad4ce | !hmaster0_p & v12ad4e0;
assign v1216269 = hbusreq5 & v1216247 | !hbusreq5 & v1216268;
assign d2fecd = hlock4_p & v845542 | !hlock4_p & !v16693aa;
assign v12aeb71 = hbusreq0 & v12afda2 | !hbusreq0 & v12aeb70;
assign d308cd = hbusreq2_p & d308cb | !hbusreq2_p & d308cc;
assign v134d200 = hlock5_p & v134d1ff | !hlock5_p & v134d1f9;
assign v16a16a9 = hbusreq0 & v16a16a6 | !hbusreq0 & v16a16a8;
assign v1515758 = hmaster2_p & v151572d | !hmaster2_p & v1515757;
assign v1215bf8 = hgrant5_p & v1215bda | !hgrant5_p & v1215bf7;
assign d2fee4 = hbusreq5_p & d2fee3 | !hbusreq5_p & d2febc;
assign d2fd0c = hbusreq2 & d2fd0b | !hbusreq2 & d2fcd8;
assign v1214eea = hbusreq5_p & v1214ee8 | !hbusreq5_p & v1214ee9;
assign v12ad02a = hgrant5_p & v12ad663 | !hgrant5_p & !v12ad013;
assign v14058c3 = hmaster2_p & v14058c2 | !hmaster2_p & v14463b1;
assign v151581b = hmaster1_p & v151581a | !hmaster1_p & v151566b;
assign v1446628 = hlock1 & v1446600 | !hlock1 & v1446627;
assign v14464a3 = hgrant2_p & v1446461 | !hgrant2_p & v14464a2;
assign v10d40d4 = hmaster1_p & v10d40d3 | !hmaster1_p & v10d407c;
assign a66287 = hgrant5_p & v845542 | !hgrant5_p & a66286;
assign v144577d = hbusreq2_p & v144577a | !hbusreq2_p & v144577c;
assign v1215329 = hmaster1_p & v1215328 | !hmaster1_p & v121546f;
assign v1446345 = hgrant2_p & v1446309 | !hgrant2_p & v1446344;
assign v12ad52a = hmaster1_p & v12ad529 | !hmaster1_p & !v12ad525;
assign v1445bde = hready_p & v1445bca | !hready_p & v1445bdd;
assign d30129 = hmaster1_p & d30128 | !hmaster1_p & v84555a;
assign v1215ce8 = hbusreq5_p & v1215ce7 | !hbusreq5_p & v1215c95;
assign a653cc = hgrant0_p & a653cb | !hgrant0_p & v845570;
assign v14463ba = hbusreq0_p & v14463b1 | !hbusreq0_p & !v144639e;
assign v85e750 = hbusreq2_p & v9745f6 | !hbusreq2_p & !v845542;
assign v1215015 = hgrant5_p & v12153be | !hgrant5_p & v1215014;
assign v1216031 = hbusreq3 & v121602c | !hbusreq3 & !v1216030;
assign v1284ccd = hgrant1_p & v1284ccc | !hgrant1_p & !v1405845;
assign v1215ba8 = hmaster0_p & v1215ba7 | !hmaster0_p & v845542;
assign v1405ae6 = hbusreq4_p & v1405ae5 | !hbusreq4_p & d3070c;
assign v16a1cd8 = hmaster1_p & v16a1cd0 | !hmaster1_p & v16a2672;
assign v1216a6a = hbusreq5_p & v1216a69 | !hbusreq5_p & v845542;
assign v1553515 = hbusreq5 & v1553513 | !hbusreq5 & v1553514;
assign v14453b0 = hlock2 & v1445354 | !hlock2 & v14453af;
assign v144619e = hgrant2_p & v144619c | !hgrant2_p & v144619d;
assign v1446701 = hlock2 & v1446700 | !hlock2 & v14466f7;
assign v12ae1f0 = hgrant4_p & v845542 | !hgrant4_p & !v12ae1ef;
assign v1552d8e = hmaster0_p & v1552d83 | !hmaster0_p & v1552d8d;
assign d30653 = hlock5_p & v845542 | !hlock5_p & d30652;
assign v1216146 = hbusreq0_p & v16a19a4 | !hbusreq0_p & v121611f;
assign v1389d75 = hmaster1_p & v845542 | !hmaster1_p & v1389d74;
assign v134d512 = hlock0 & v134d511 | !hlock0 & v134d50c;
assign v1445846 = hgrant2_p & v1445820 | !hgrant2_p & v1445845;
assign a656c1 = hmaster1_p & a66287 | !hmaster1_p & a656c0;
assign v1445ea0 = hgrant5_p & v1445e05 | !hgrant5_p & v1445e9f;
assign v1552f77 = hlock3 & v155341e | !hlock3 & v1552f76;
assign v1515739 = hgrant5_p & v1515639 | !hgrant5_p & v1515737;
assign v1215c9d = hbusreq5_p & v1215c9b | !hbusreq5_p & !v1215c9c;
assign v16a1e5a = hbusreq0_p & v845542 | !hbusreq0_p & !v845547;
assign v134d311 = hgrant1_p & v845542 | !hgrant1_p & v134d310;
assign v138a43a = hbusreq5_p & v138a316 | !hbusreq5_p & v845542;
assign v134d28b = hbusreq4_p & v134d28a | !hbusreq4_p & v845542;
assign d30750 = hbusreq3 & d3073a | !hbusreq3 & d3074f;
assign d3012f = hgrant5_p & d2fe80 | !hgrant5_p & d300c5;
assign v16a1cc2 = hmaster1_p & v16a1c9f | !hmaster1_p & v16a1f96;
assign a65492 = hbusreq2 & a6548a | !hbusreq2 & a65491;
assign d2fd08 = hbusreq2 & d2fd01 | !hbusreq2 & d2fcd8;
assign v1553234 = hgrant4_p & v845542 | !hgrant4_p & v1553233;
assign v16a1d7d = hgrant2_p & v845542 | !hgrant2_p & !v16a1d7c;
assign d2fc05 = hbusreq0 & d2fc04 | !hbusreq0 & v845542;
assign v134d219 = hmaster0_p & v134d1e8 | !hmaster0_p & v134d218;
assign v1215760 = hmaster2_p & v845542 | !hmaster2_p & v121575f;
assign v138a452 = hlock2_p & v138a44f | !hlock2_p & v138a451;
assign v14458c3 = hmaster1_p & v14458a7 | !hmaster1_p & v14458c1;
assign d30216 = hbusreq5_p & d30215 | !hbusreq5_p & d30214;
assign v138a033 = hmaster1_p & v1389ffe | !hmaster1_p & !v138a032;
assign v12165a6 = hmaster1_p & v121658b | !hmaster1_p & v12165a5;
assign v144612a = hmaster0_p & v144608a | !hmaster0_p & v1445fe3;
assign d2fb32 = hbusreq5 & d2fb17 | !hbusreq5 & d2fb31;
assign v12af5ae = hmaster0_p & v12afe47 | !hmaster0_p & v12af5ad;
assign v1445a8a = hmaster1_p & v1445a5b | !hmaster1_p & v1445a82;
assign v1215bcb = hlock2_p & v1215bca | !hlock2_p & v1215bc4;
assign v1668d29 = hmaster2_p & v1668d28 | !hmaster2_p & v845542;
assign v1389374 = hready_p & v845542 | !hready_p & v1389373;
assign v1215bb4 = hmaster0_p & v845542 | !hmaster0_p & v1216b01;
assign v1214ebb = hlock2_p & v1214eba | !hlock2_p & !v1215bc4;
assign v16a2087 = hgrant5_p & v845542 | !hgrant5_p & v16a2086;
assign v12ad5e1 = hmaster0_p & v12ad5cf | !hmaster0_p & v12ad5e0;
assign v1552f55 = hlock1 & v1553217 | !hlock1 & v1552f54;
assign v1405a97 = hmaster0_p & v1405a89 | !hmaster0_p & v1405a96;
assign v12ae1f4 = hlock0_p & v1515ae4 | !hlock0_p & !v845542;
assign v16a1af5 = stateG2_p & v845542 | !stateG2_p & v845588;
assign v144553e = hmaster0_p & v144639c | !hmaster0_p & v14463be;
assign v1445fe5 = hmaster1_p & v1445fe4 | !hmaster1_p & v1445fde;
assign v1445ff3 = hbusreq2_p & v1445ff0 | !hbusreq2_p & v1445ff2;
assign v1405a9f = decide_p & v1405a9e | !decide_p & v1405a99;
assign v1668c8b = hmaster1_p & v1668c8a | !hmaster1_p & v1668c7d;
assign v1215396 = hbusreq0 & v1215395 | !hbusreq0 & v845542;
assign d807a9 = hgrant1_p & d80760 | !hgrant1_p & d807a8;
assign v16a1a77 = hbusreq1_p & v16a1940 | !hbusreq1_p & v16a1a76;
assign d30646 = hgrant0_p & a6537d | !hgrant0_p & !d30645;
assign v1215c93 = hbusreq1_p & v1216521 | !hbusreq1_p & !v845542;
assign d307e0 = hbusreq5_p & d307df | !hbusreq5_p & d307de;
assign d2fee9 = hbusreq2_p & d2fee8 | !hbusreq2_p & d2fee7;
assign v1445dd3 = hmaster1_p & v1445db2 | !hmaster1_p & v1445dd1;
assign v1215cb0 = hmaster2_p & v1215c99 | !hmaster2_p & v1215caf;
assign v14465b6 = hmaster2_p & v144639c | !hmaster2_p & v14465b3;
assign v144541a = hmaster1_p & v1445419 | !hmaster1_p & v1445bd5;
assign d2fb9d = hmaster0_p & d2fb9c | !hmaster0_p & d2fb7a;
assign v1552d52 = hlock0 & v1552d51 | !hlock0 & v1553413;
assign v14458c5 = hmaster1_p & v14458ab | !hmaster1_p & v14458c1;
assign v1215732 = hbusreq1 & v1215b7b | !hbusreq1 & v1215b92;
assign v88d3e4 = hburst1_p & v845542 | !hburst1_p & v845560;
assign d307fb = hgrant5_p & d306e6 | !hgrant5_p & d307fa;
assign v134d211 = hmaster1_p & v134d20b | !hmaster1_p & v134d20f;
assign v15157fa = hmaster1_p & v15157e5 | !hmaster1_p & v15157f9;
assign v1215b94 = hmaster0_p & v1215b93 | !hmaster0_p & v845542;
assign v1214f63 = hbusreq5 & v1214f59 | !hbusreq5 & v1214f62;
assign v16a1d36 = decide_p & v16a1d2b | !decide_p & !v16a1d35;
assign d305d9 = hlock5_p & v845542 | !hlock5_p & v1668c21;
assign v16a20a6 = decide_p & v16a20a0 | !decide_p & v16a20a5;
assign v16a19af = hmaster2_p & v16a19aa | !hmaster2_p & v845542;
assign v14465e5 = hbusreq0 & v14465de | !hbusreq0 & v14465e4;
assign v12ad566 = hmaster0_p & v12ad565 | !hmaster0_p & v12ad528;
assign v12165b2 = hbusreq2_p & v12165a7 | !hbusreq2_p & v12165b1;
assign v144584c = hgrant2_p & v1445824 | !hgrant2_p & v1445848;
assign v16a19b1 = hmaster0_p & v16a19ac | !hmaster0_p & v16a19b0;
assign v1446222 = hbusreq2_p & v144621a | !hbusreq2_p & v1446221;
assign v134cedb = hbusreq3 & v134ced9 | !hbusreq3 & v134ceda;
assign v16a13f9 = hlock2_p & v16a13f1 | !hlock2_p & v16a13f8;
assign v1445773 = hlock5 & v1445f40 | !hlock5 & v1445771;
assign d2faf6 = hgrant1_p & d2faf4 | !hgrant1_p & d2faf5;
assign v1214c10 = hbusreq2 & v1214c0a | !hbusreq2 & v1214c0f;
assign v10d42b3 = hmaster2_p & v10d42b2 | !hmaster2_p & !v10d4062;
assign v121509b = hgrant1_p & v1215466 | !hgrant1_p & v1215095;
assign v16a224a = hbusreq2 & v16a2242 | !hbusreq2 & v16a2249;
assign v121624a = hbusreq5_p & v1216249 | !hbusreq5_p & v1216214;
assign v140592c = hbusreq1_p & v1405890 | !hbusreq1_p & v140592b;
assign d30663 = hmaster2_p & d30662 | !hmaster2_p & v845542;
assign v16a20a1 = hmaster1_p & v16a2094 | !hmaster1_p & v16a2095;
assign v134d53e = decide_p & v134d3ce | !decide_p & v134d52a;
assign a658a5 = stateG2_p & v845542 | !stateG2_p & a658a3;
assign d2fefd = hmaster0_p & d2fec8 | !hmaster0_p & d2fecf;
assign v1215739 = hgrant0_p & v1215737 | !hgrant0_p & v1215738;
assign v15530aa = hmaster1_p & v15530a9 | !hmaster1_p & v845542;
assign v14463b2 = hbusreq0_p & v14463b1 | !hbusreq0_p & !v14463a0;
assign v134d37d = hbusreq4 & v134d36f | !hbusreq4 & v134d273;
assign v144618b = hgrant2_p & v1446188 | !hgrant2_p & v144618a;
assign v15530f5 = hgrant3_p & v155321c | !hgrant3_p & v15530f4;
assign v15155f8 = hbusreq0_p & d305de | !hbusreq0_p & d30645;
assign v1214cef = hbusreq0 & v1214cee | !hbusreq0 & v16a2243;
assign v1515616 = hmaster0_p & v1515611 | !hmaster0_p & v1515615;
assign v1446160 = hready_p & v14460e6 | !hready_p & v144615f;
assign v155298c = hgrant3_p & v155321c | !hgrant3_p & v155298b;
assign v12ad8e7 = hbusreq4_p & v12add47 | !hbusreq4_p & !v845542;
assign a64717 = jx1_p & a646d9 | !jx1_p & a64716;
assign v14458f4 = hlock0_p & v14458f2 | !hlock0_p & v14458f3;
assign d307fa = hmaster2_p & d30793 | !hmaster2_p & d307b7;
assign v144644b = hbusreq2_p & v1446437 | !hbusreq2_p & v144644a;
assign v1552f81 = hgrant2_p & v1552f71 | !hgrant2_p & v1552f7f;
assign v1214bd9 = hmaster1_p & v1214bbd | !hmaster1_p & v1214bcf;
assign d3019f = hmaster1_p & d3090e | !hmaster1_p & !d3019e;
assign v10d42b9 = hmaster0_p & v10d42b4 | !hmaster0_p & v10d42b8;
assign v15167f7 = hlock5_p & v1668c1d | !hlock5_p & d305df;
assign v1553093 = hlock3 & v155341e | !hlock3 & v1553092;
assign f2f2ce = hbusreq1 & a658c6 | !hbusreq1 & !v845542;
assign v12150cc = hlock0_p & v12150c2 | !hlock0_p & v845547;
assign v16a1e95 = hgrant4_p & v845559 | !hgrant4_p & !v16a1e94;
assign v1445e13 = hlock0 & v1445e12 | !hlock0 & v1445e11;
assign f2f383 = hbusreq1 & a653c4 | !hbusreq1 & v845542;
assign v1445b58 = hgrant5_p & v1445b55 | !hgrant5_p & v1445b57;
assign d2fc41 = hmaster0_p & d2fc40 | !hmaster0_p & d2fc3a;
assign v15155fc = hmaster0_p & v15155f7 | !hmaster0_p & v15155fb;
assign v12af9bd = hgrant0_p & v12af9bc | !hgrant0_p & !v1405a7d;
assign a65698 = hbusreq2_p & a65692 | !hbusreq2_p & a65693;
assign v1216242 = hbusreq2_p & v121623e | !hbusreq2_p & v1216241;
assign v1214d80 = hbusreq2 & v1214d7c | !hbusreq2 & v1214d7f;
assign v16a1d41 = hmaster2_p & v16a1d3c | !hmaster2_p & v16a1d40;
assign d2fee3 = hlock5_p & d2fee2 | !hlock5_p & d2febc;
assign v12ad551 = hmaster1_p & v12ad529 | !hmaster1_p & v12ad54f;
assign v1215417 = hbusreq2 & v1215413 | !hbusreq2 & v1215416;
assign v12150b8 = hmaster1_p & v12150b7 | !hmaster1_p & !v1215ba1;
assign f2ed9a = hbusreq2_p & f2ed94 | !hbusreq2_p & f2ed99;
assign v1405a8a = hmaster2_p & v1405a86 | !hmaster2_p & !v845542;
assign v1445403 = hready_p & v144639b | !hready_p & v1445402;
assign v14457f2 = hmaster0_p & v1445eb6 | !hmaster0_p & v1445eae;
assign v1215319 = hmaster1_p & v1215318 | !hmaster1_p & v12153bf;
assign v14462a4 = decide_p & v1446260 | !decide_p & v14462a3;
assign v14462f7 = hbusreq0 & v14462f6 | !hbusreq0 & v1446616;
assign v134d1e9 = stateA1_p & v144646d | !stateA1_p & v134d1e6;
assign v1215c77 = hgrant2_p & v121657d | !hgrant2_p & v1215c73;
assign v15168ec = hmaster1_p & v15168eb | !hmaster1_p & v845570;
assign d3011e = hbusreq0 & d30118 | !hbusreq0 & d3011d;
assign v144670b = hmaster0_p & v1446657 | !hmaster0_p & v1446448;
assign v15157b0 = hgrant5_p & v15157a6 | !hgrant5_p & v15157af;
assign v1389f8e = hmaster0_p & v1389f8d | !hmaster0_p & v845542;
assign v1215323 = hmaster0_p & v1215471 | !hmaster0_p & v1215057;
assign v12153a3 = hbusreq0_p & v1216add | !hbusreq0_p & v845542;
assign v1445fbb = hbusreq0 & v1445fba | !hbusreq0 & v1445f8f;
assign d2ff06 = hmaster1_p & d2fefd | !hmaster1_p & d2fee5;
assign v12af9b4 = hmaster0_p & v12af73f | !hmaster0_p & v12af9b3;
assign v1215447 = hbusreq2_p & v1215446 | !hbusreq2_p & v1215445;
assign d30732 = hbusreq2_p & d30731 | !hbusreq2_p & d30730;
assign v12af3a9 = hmaster2_p & v845542 | !hmaster2_p & v12af3a8;
assign v144668b = hbusreq1_p & v144639c | !hbusreq1_p & v144668a;
assign v10d40c7 = hbusreq2_p & v10d40b7 | !hbusreq2_p & !v10d40c6;
assign d2fc8b = hbusreq2_p & d2fc8a | !hbusreq2_p & v845542;
assign v1516201 = decide_p & v1516200 | !decide_p & v845576;
assign v14465b5 = hgrant5_p & v1446404 | !hgrant5_p & v14465b4;
assign v134d426 = hbusreq1_p & v134d425 | !hbusreq1_p & v134d380;
assign a656bc = hbusreq0 & a66287 | !hbusreq0 & a6628c;
assign a658fe = hmaster1_p & a658fd | !hmaster1_p & a658e5;
assign v12167a3 = hmaster0_p & v12165ae | !hmaster0_p & v121658b;
assign v134d4de = hgrant2_p & v134d27a | !hgrant2_p & v134d4dd;
assign v12ad53f = hbusreq2_p & v12ad53c | !hbusreq2_p & v12ad53e;
assign v1216a8a = stateA1_p & v845542 | !stateA1_p & !v1216a89;
assign v1215752 = hgrant5_p & v1215743 | !hgrant5_p & v1215751;
assign d30719 = hbusreq1 & d30718 | !hbusreq1 & v845542;
assign d2feea = hmaster1_p & d2fed0 | !hmaster1_p & d2fee5;
assign d30878 = hbusreq2_p & d30776 | !hbusreq2_p & d30876;
assign d2f972 = hbusreq1_p & d2fe9c | !hbusreq1_p & d2f971;
assign d2fef5 = hbusreq2 & d2fef1 | !hbusreq2 & d2fef4;
assign v151697a = hmaster1_p & v1516979 | !hmaster1_p & v845542;
assign v1405aa2 = hmastlock_p & v1405aa1 | !hmastlock_p & !v845542;
assign v134d290 = hgrant4_p & v845542 | !hgrant4_p & v134d28f;
assign v144639a = hmaster0_p & v1446399 | !hmaster0_p & v845542;
assign v16a1435 = hbusreq3_p & v16a141e | !hbusreq3_p & v16a1434;
assign v1215c7f = hmaster2_p & v1216a5a | !hmaster2_p & v1215c7e;
assign v1553137 = hmastlock_p & v1553934 | !hmastlock_p & v845542;
assign v15167be = hlock5_p & v1668c2e | !hlock5_p & v15167bd;
assign v1405ad5 = hgrant4_p & v1405a86 | !hgrant4_p & v1405ad4;
assign d2fb27 = hgrant5_p & d2f981 | !hgrant5_p & !d2fb0c;
assign v1216705 = hgrant2_p & v12166ff | !hgrant2_p & v1216704;
assign v16a137b = hmaster1_p & v16a132e | !hmaster1_p & v16a1f96;
assign stateG10_2 = !c50efe;
assign v1445819 = hbusreq2 & v1445813 | !hbusreq2 & v1445818;
assign v12165aa = hmaster0_p & v1216a91 | !hmaster0_p & v12165a9;
assign v1446169 = hgrant2_p & v1446167 | !hgrant2_p & v1446168;
assign v1445e51 = hbusreq2_p & v1445e4c | !hbusreq2_p & v1445e50;
assign v1516980 = hlock2_p & v151697f | !hlock2_p & v845542;
assign v16a1948 = hbusreq4 & v16a1bc6 | !hbusreq4 & !v845542;
assign v151579a = hgrant4_p & a662a9 | !hgrant4_p & a65382;
assign v1214c04 = hbusreq2 & v1214bfd | !hbusreq2 & v1214c03;
assign a65680 = hbusreq2 & a6567c | !hbusreq2 & a6567f;
assign v1668c41 = hmaster2_p & v1668c3f | !hmaster2_p & !v1668c40;
assign v140587c = locked_p & v1405839 | !locked_p & !v144639c;
assign d2fed9 = hmaster1_p & d2fed8 | !hmaster1_p & d2fec6;
assign v10d40b9 = hmaster1_p & v10d40b8 | !hmaster1_p & v10d3ffb;
assign b09421 = hbusreq5_p & v845568 | !hbusreq5_p & v845542;
assign v12152f7 = hgrant2_p & v12152e8 | !hgrant2_p & v12152f6;
assign d300c6 = hgrant5_p & d2fe81 | !hgrant5_p & d300c5;
assign v1214dde = hlock3_p & v1214ddb | !hlock3_p & v1214ddd;
assign v1284c9b = hmaster2_p & v1284c8e | !hmaster2_p & v1284c9a;
assign v143fd7b = hgrant2_p & v845542 | !hgrant2_p & !v143fd7a;
assign v1445fd5 = hbusreq1_p & v1446425 | !hbusreq1_p & v1446429;
assign v16a1d05 = jx2_p & v16a1af4 | !jx2_p & v16a1d04;
assign v1445f84 = hbusreq3_p & v14466c8 | !hbusreq3_p & v1445f83;
assign v1216283 = hmaster1_p & v1216282 | !hmaster1_p & !v1216027;
assign v166939e = hmaster1_p & v166939d | !hmaster1_p & v845570;
assign v1515796 = hmaster2_p & v1515793 | !hmaster2_p & v1515795;
assign v10d404a = hgrant1_p & v10d4044 | !hgrant1_p & v10d4049;
assign v121625d = hmaster2_p & v121625c | !hmaster2_p & v12161da;
assign v1446089 = hbusreq0 & v1446088 | !hbusreq0 & v1446077;
assign a65439 = hmaster0_p & a6542e | !hmaster0_p & a65438;
assign v15157d7 = hgrant5_p & v845570 | !hgrant5_p & v1515724;
assign f2f32d = hmaster2_p & f2f2e2 | !hmaster2_p & f2f21f;
assign v1445b33 = hmaster0_p & v1445a43 | !hmaster0_p & v14459a3;
assign v144590e = hmaster0_p & v14458ee | !hmaster0_p & v14458fa;
assign v1216074 = hmaster1_p & v1216073 | !hmaster1_p & v121605d;
assign v16a1bf1 = hgrant5_p & v845542 | !hgrant5_p & v16a1bf0;
assign a658f4 = hmaster1_p & a658f2 | !hmaster1_p & a658e5;
assign v134d220 = hlock5_p & v134d1e8 | !hlock5_p & v134d21f;
assign v16a13f2 = hgrant5_p & v845542 | !hgrant5_p & !v16a2077;
assign v1515713 = hbusreq4 & v1515609 | !hbusreq4 & v845570;
assign v151571d = busreq_p & v88d3e4 | !busreq_p & v151571c;
assign v1446606 = hbusreq4_p & v144639c | !hbusreq4_p & v14465bb;
assign v13891a1 = hmaster2_p & v1515c80 | !hmaster2_p & v845542;
assign v144663f = hgrant1_p & v1446439 | !hgrant1_p & v144663e;
assign v14463e6 = hlock0_p & v144639c | !hlock0_p & !v14463e5;
assign d308be = hbusreq5_p & d30821 | !hbusreq5_p & d308bd;
assign a6540b = hgrant2_p & a6540a | !hgrant2_p & a653e8;
assign v134cf3f = decide_p & v134cedd | !decide_p & v134cecd;
assign v1445376 = hlock3 & v144535e | !hlock3 & v1445375;
assign v14458ad = hbusreq2_p & v14458a0 | !hbusreq2_p & v14458ac;
assign d307cd = hgrant1_p & v845542 | !hgrant1_p & d307cc;
assign v1215fbb = hmaster0_p & v12164e3 | !hmaster0_p & v12166fd;
assign v1515776 = hgrant5_p & v1515615 | !hgrant5_p & v1515775;
assign v1405929 = hgrant0_p & v140588c | !hgrant0_p & !v1405928;
assign a6629c = hbusreq5_p & a6629b | !hbusreq5_p & a6628c;
assign v10d3fe4 = hbusreq5_p & v10d3fe2 | !hbusreq5_p & v10d3fe3;
assign v1445437 = hbusreq2 & v1445436 | !hbusreq2 & v144542f;
assign v15533b7 = hmaster1_p & v1553385 | !hmaster1_p & v15533b6;
assign f2ed99 = hgrant2_p & v845542 | !hgrant2_p & f2ed98;
assign v10d4037 = hlock5_p & v10d4034 | !hlock5_p & v10d4036;
assign d3020a = hgrant1_p & d30209 | !hgrant1_p & d307d7;
assign d300e7 = hlock1_p & d300e5 | !hlock1_p & d300e6;
assign v1389446 = hmaster2_p & v1389445 | !hmaster2_p & v845542;
assign v1389fdc = hlock5_p & v1389fdb | !hlock5_p & !v845542;
assign v134d21a = hmaster1_p & v134d219 | !hmaster1_p & v134d208;
assign v138a317 = hmaster0_p & v138a30e | !hmaster0_p & v138a316;
assign a653a9 = hbusreq4_p & a65861 | !hbusreq4_p & !v845542;
assign v12af5a3 = hgrant1_p & v845542 | !hgrant1_p & v12af5a2;
assign v14058e1 = hmaster1_p & v14058e0 | !hmaster1_p & v14058d8;
assign d2fd45 = hbusreq2 & d2fd44 | !hbusreq2 & d302ec;
assign v1215784 = hmaster1_p & v1215783 | !hmaster1_p & v845542;
assign v1552d9e = decide_p & v1553443 | !decide_p & v1552d95;
assign f2f27f = hready_p & f2f23d | !hready_p & f2f27e;
assign f2f28a = hmaster0_p & f2f289 | !hmaster0_p & f2f284;
assign v134d4c5 = hready_p & v134d3e5 | !hready_p & v134d4c4;
assign d30611 = hmaster2_p & v16693aa | !hmaster2_p & v1668c2d;
assign v144586c = hbusreq0_p & v14463a0 | !hbusreq0_p & v144639e;
assign v1215c17 = hgrant5_p & v1215c12 | !hgrant5_p & v1215c16;
assign v1446736 = hmaster0_p & v144643e | !hmaster0_p & v144639c;
assign v10d42de = hready_p & v10d42d6 | !hready_p & !v10d42dd;
assign v12ae6fe = decide_p & v12afe72 | !decide_p & v12afe76;
assign v16a1403 = hmaster0_p & v16a1d7a | !hmaster0_p & v16a1d78;
assign f2e4cc = decide_p & f2e4cb | !decide_p & v845542;
assign d30634 = hmaster1_p & d30633 | !hmaster1_p & d30608;
assign v1389ddf = hgrant5_p & v845570 | !hgrant5_p & !v845542;
assign v144648c = hbusreq4_p & v1446398 | !hbusreq4_p & v1446476;
assign a65917 = hmaster1_p & a658b7 | !hmaster1_p & !a65916;
assign v16a142d = hbusreq2 & v16a142c | !hbusreq2 & !v16a1db6;
assign v1215332 = hgrant2_p & v1215324 | !hgrant2_p & v1215331;
assign v1389ffb = hgrant5_p & v1668da6 | !hgrant5_p & !v845542;
assign v10d42d5 = hbusreq2_p & v10d42d2 | !hbusreq2_p & v10d42d4;
assign v1445888 = hbusreq1 & v1445882 | !hbusreq1 & v1445887;
assign f2f2ac = hmaster0_p & f2f2ab | !hmaster0_p & f2f2a8;
assign v1668c87 = hmaster0_p & v1668c5f | !hmaster0_p & v1668c86;
assign v15530af = hlock5 & v155321a | !hlock5 & v15530ae;
assign f2e4d4 = decide_p & f2e4cb | !decide_p & f2f23c;
assign d300fa = hbusreq1_p & d300f9 | !hbusreq1_p & d300f8;
assign v1445b3d = hbusreq2_p & v1445b35 | !hbusreq2_p & v1445b39;
assign v16a12c7 = hbusreq5 & v16a12bf | !hbusreq5 & v16a12c6;
assign v1445e2f = hlock2 & v1445e1f | !hlock2 & v1445e2d;
assign d3079a = hlock5_p & d30798 | !hlock5_p & !d30799;
assign v11e595e = hgrant2_p & v11e5943 | !hgrant2_p & v11e595d;
assign v16a1a21 = hbusreq2_p & v16a1848 | !hbusreq2_p & v16a1a20;
assign d2fef8 = hmaster0_p & d2fec8 | !hmaster0_p & d2feb5;
assign v1284cf3 = hbusreq4_p & v1284c8f | !hbusreq4_p & v1284ce9;
assign v1552f6c = hbusreq1 & v1552f54 | !hbusreq1 & v1552f55;
assign v1405ac5 = hbusreq0_p & v845542 | !hbusreq0_p & v1405abf;
assign v1215bfc = hmaster2_p & v1215fe8 | !hmaster2_p & v1216a5a;
assign v134cdcf = hbusreq3_p & v134cd8f | !hbusreq3_p & v134cdce;
assign v16a1d19 = hready & v16a1d18 | !hready & v845542;
assign v16695c6 = hgrant3_p & v16695bd | !hgrant3_p & !v16695c5;
assign v1445414 = hgrant5_p & v1446404 | !hgrant5_p & v1445413;
assign d3075b = hbusreq2_p & d3075a | !hbusreq2_p & d30756;
assign v144673e = hgrant2_p & v144673c | !hgrant2_p & v144673d;
assign v1445831 = hmaster1_p & v1445808 | !hmaster1_p & v1445e28;
assign v138a439 = hbusreq5_p & v138a3e3 | !hbusreq5_p & v845542;
assign v16a2673 = hmaster1_p & v16a266a | !hmaster1_p & !v16a2672;
assign v144591a = hlock0 & v1445919 | !hlock0 & v1445918;
assign v1215c29 = hgrant1_p & v1215c28 | !hgrant1_p & v121614c;
assign v14463d0 = hmaster1_p & v14463cf | !hmaster1_p & v14463cd;
assign v134d244 = hmaster1_p & v134d20a | !hmaster1_p & v134d208;
assign v12162b6 = hgrant2_p & v12162b3 | !hgrant2_p & v12162b5;
assign v134ce8d = hmaster2_p & v134d1e8 | !hmaster2_p & v134ce8c;
assign v134cec8 = hbusreq2 & v134cec7 | !hbusreq2 & v134d3b5;
assign v134cee7 = hready_p & v134d3be | !hready_p & v134cee6;
assign v138a479 = hmaster1_p & v138a478 | !hmaster1_p & v138a301;
assign d308f6 = hmaster0_p & d308f5 | !hmaster0_p & v845542;
assign v14461fe = hlock3 & v14461ec | !hlock3 & v14461fd;
assign v134cec1 = decide_p & v134cec0 | !decide_p & v134d276;
assign v1405904 = hready_p & v14058e4 | !hready_p & v1405903;
assign d308f7 = hmaster1_p & v845542 | !hmaster1_p & d308f6;
assign v1445a30 = hbusreq0 & v1445a1c | !hbusreq0 & v1445a2f;
assign v1405ad4 = hgrant0_p & v1405a86 | !hgrant0_p & v1405ad3;
assign v134d225 = hmaster1_p & v134d224 | !hmaster1_p & v134d20f;
assign v14459b2 = hlock1 & v14459ac | !hlock1 & v14459b1;
assign v1445fa7 = hmaster2_p & v144639c | !hmaster2_p & v1445fa6;
assign v134cd85 = hlock2 & v134cd82 | !hlock2 & v134cd84;
assign v16a19c8 = hmaster1_p & v16a19b0 | !hmaster1_p & v16a1f96;
assign v12152ec = hmaster0_p & v1215ba3 | !hmaster0_p & v1215773;
assign v11ac6c8 = decide_p & v11ac602 | !decide_p & v11ac6a3;
assign v1215bdb = hmaster2_p & v1215fe8 | !hmaster2_p & v1216a61;
assign v144612d = hmaster0_p & v144608a | !hmaster0_p & v1445fea;
assign v15534f7 = hlock3 & v155341e | !hlock3 & v15534f6;
assign v12afe5e = hgrant5_p & v845542 | !hgrant5_p & v12afe5d;
assign f2f3f6 = hmaster1_p & f2f3f5 | !hmaster1_p & f2f2db;
assign v15534fc = hbusreq0 & v15534fb | !hbusreq0 & v1553395;
assign d3026e = hmaster2_p & d30268 | !hmaster2_p & d3064a;
assign v14058f1 = locked_p & v845542 | !locked_p & !v1405844;
assign v1284cc3 = hmaster1_p & v1284cc2 | !hmaster1_p & v140584d;
assign d2fb7a = hbusreq0 & d2fb79 | !hbusreq0 & v845542;
assign v144628c = hmaster2_p & v1446444 | !hmaster2_p & v1446410;
assign v155308b = hbusreq0 & v155308a | !hbusreq0 & v1553218;
assign v1446189 = hmaster0_p & v1446092 | !hmaster0_p & v1446081;
assign d2fbfc = hbusreq0 & d2fbfb | !hbusreq0 & v845542;
assign v85e75b = hmaster1_p & v845558 | !hmaster1_p & a1db63;
assign v138981d = decide_p & v138981c | !decide_p & v138a406;
assign v15533aa = hbusreq0_p & v1553217 | !hbusreq0_p & v155338c;
assign v134d375 = hmaster2_p & v845542 | !hmaster2_p & v134d374;
assign v121621a = hbusreq1_p & v1216219 | !hbusreq1_p & v845542;
assign v12150a7 = hmaster1_p & v1215092 | !hmaster1_p & !v12150a6;
assign d302f8 = jx2_p & d302f0 | !jx2_p & d302f7;
assign a65b13 = hgrant5_p & v845542 | !hgrant5_p & a65b12;
assign v1214cba = hmaster1_p & v1214cb9 | !hmaster1_p & v1215388;
assign v14058dc = hmaster0_p & v1405841 | !hmaster0_p & v14058db;
assign v12afa0d = hmaster1_p & v12af9c3 | !hmaster1_p & v12afa0c;
assign a653d0 = hgrant1_p & a653c7 | !hgrant1_p & !a653cf;
assign v1445f69 = hmaster0_p & v14466af | !hmaster0_p & v1446663;
assign v1446262 = hmaster2_p & v1446444 | !hmaster2_p & v14465b9;
assign v151576a = hbusreq1_p & v1515768 | !hbusreq1_p & v1515769;
assign v1445a7f = hbusreq5_p & v14459fe | !hbusreq5_p & v1445a7e;
assign v134d532 = hmaster1_p & v134d531 | !hmaster1_p & v845542;
assign v10d408b = hmaster2_p & v10d3fd4 | !hmaster2_p & !v10d4062;
assign d2fb6c = hbusreq0 & d2fb6b | !hbusreq0 & v845542;
assign v1216121 = hlock0_p & v1215ff8 | !hlock0_p & v121601f;
assign v1515793 = hgrant1_p & f2f281 | !hgrant1_p & v1515792;
assign a65464 = decide_p & a65463 | !decide_p & v845542;
assign a65888 = hburst0 & a66293 | !hburst0 & a65886;
assign d80788 = stateA1_p & v845542 | !stateA1_p & v936735;
assign a65861 = hmastlock_p & v88d3e4 | !hmastlock_p & v845542;
assign v10d405f = hgrant1_p & v10d3fd5 | !hgrant1_p & v10d405e;
assign v1216128 = hgrant5_p & v121611d | !hgrant5_p & v1216127;
assign d301ee = hgrant5_p & d301bd | !hgrant5_p & d301ed;
assign d30205 = hbusreq1_p & d30204 | !hbusreq1_p & d30203;
assign v134d51a = hmaster0_p & v845542 | !hmaster0_p & v134d519;
assign v1215b7d = hbusreq4_p & v1216523 | !hbusreq4_p & v845542;
assign d30739 = hbusreq2_p & d30738 | !hbusreq2_p & d30730;
assign v144641f = hbusreq1 & v144641c | !hbusreq1 & v144641e;
assign d2f99d = hbusreq1_p & d2f98b | !hbusreq1_p & d30660;
assign v121609d = hbusreq2_p & v121609c | !hbusreq2_p & v121609b;
assign v14466e5 = hbusreq2_p & v14466e2 | !hbusreq2_p & v14466e4;
assign d307ea = hbusreq1 & d307e9 | !hbusreq1 & v845542;
assign v10a1540 = hgrant5_p & v845542 | !hgrant5_p & v845574;
assign v10d427b = stateA1_p & v84557e | !stateA1_p & !v10d427a;
assign v134cd6d = hgrant2_p & v134d364 | !hgrant2_p & v134cd6c;
assign v16a1e06 = hmaster1_p & v16a1d6c | !hmaster1_p & v16a1d53;
assign v1216565 = hgrant4_p & v1216553 | !hgrant4_p & v845542;
assign v1446102 = hmaster1_p & v14460e7 | !hmaster1_p & v1445fbd;
assign v1445ecc = hlock0 & v1445ecb | !hlock0 & v1445eca;
assign v151578b = stateG2_p & v845542 | !stateG2_p & v151578a;
assign v151575f = hbusreq1 & v1515612 | !hbusreq1 & v845570;
assign v151566a = hbusreq0 & v1668c6f | !hbusreq0 & v1515669;
assign v144575f = hbusreq2_p & v1445757 | !hbusreq2_p & v144575e;
assign v1216100 = hgrant1_p & v845542 | !hgrant1_p & v12160ff;
assign d307c2 = hbusreq5_p & d307ab | !hbusreq5_p & d307c1;
assign v16a13c9 = hlock2_p & v16a13c6 | !hlock2_p & !v16a13c8;
assign v151574f = hbusreq1_p & v151574d | !hbusreq1_p & !v151574e;
assign v134d539 = hlock5 & v134d534 | !hlock5 & v134d538;
assign v12ad4f4 = hbusreq0 & v12ad4f3 | !hbusreq0 & v845542;
assign v1446239 = hlock0 & v1446238 | !hlock0 & v14463f3;
assign v1445417 = hmaster0_p & v1446404 | !hmaster0_p & v1446636;
assign v16a1393 = hbusreq2 & v16a1390 | !hbusreq2 & v16a1392;
assign v1216304 = hmaster1_p & v12162f7 | !hmaster1_p & v1216303;
assign v1405b53 = hgrant2_p & v1405b46 | !hgrant2_p & v1405b52;
assign d3088f = hgrant1_p & v84554c | !hgrant1_p & d3088e;
assign v1389d78 = hready_p & v845542 | !hready_p & v1389d77;
assign a65422 = hgrant5_p & a6541f | !hgrant5_p & a653a7;
assign v14463c5 = hmaster2_p & v144639c | !hmaster2_p & v144639e;
assign v1284cfe = hmaster1_p & v1284cc9 | !hmaster1_p & !v1284cfd;
assign v12ad022 = hmaster1_p & v12ad021 | !hmaster1_p & !v12ad617;
assign v151573b = hbusreq0 & v1515736 | !hbusreq0 & v151573a;
assign v1515847 = hbusreq5_p & v1515845 | !hbusreq5_p & !v1515846;
assign d2fc0b = hbusreq2 & d2fc01 | !hbusreq2 & d2fc0a;
assign v1216718 = hgrant5_p & v16a2243 | !hgrant5_p & v1216717;
assign v1515853 = hgrant3_p & v1515831 | !hgrant3_p & !v1515852;
assign v1445a88 = hbusreq2_p & v1445a84 | !hbusreq2_p & v1445a87;
assign v12ad02e = hmaster1_p & v12ad026 | !hmaster1_p & !v12ad02d;
assign v1216add = hbusreq4 & v1216ab0 | !hbusreq4 & !v1216adc;
assign d30956 = hbusreq5_p & d30955 | !hbusreq5_p & !d30954;
assign v1668c25 = hbusreq3 & v1668c1a | !hbusreq3 & v1668c24;
assign v16a1977 = hmaster1_p & v16a1972 | !hmaster1_p & v16a1976;
assign v14465fa = hgrant4_p & v1446421 | !hgrant4_p & v14465f9;
assign v16a1d5c = hbusreq0 & v16a1d58 | !hbusreq0 & v16a1d5b;
assign v16a2082 = hgrant5_p & v845542 | !hgrant5_p & v16a2081;
assign v1214ef8 = hbusreq5_p & v1214ef7 | !hbusreq5_p & v1216571;
assign v12160e5 = hbusreq2_p & v12160e1 | !hbusreq2_p & v12160e4;
assign v1445e69 = hlock1 & v1445e68 | !hlock1 & v1445e65;
assign d2fc2e = hbusreq1_p & d2fb69 | !hbusreq1_p & d2fc2d;
assign v1216170 = hmaster1_p & v1216116 | !hmaster1_p & v121616f;
assign v144626f = hmaster1_p & v144626e | !hmaster1_p & v144626a;
assign v1668d37 = hmaster2_p & v1668d28 | !hmaster2_p & v1668d36;
assign v1215caf = hgrant1_p & v1215ca3 | !hgrant1_p & v1215cae;
assign v1214c77 = hmaster2_p & v1214c4c | !hmaster2_p & v1214c61;
assign a66295 = locked_p & a66294 | !locked_p & !v845542;
assign d2fb36 = hbusreq5_p & d2febd | !hbusreq5_p & d2fb35;
assign v1553139 = hmaster2_p & v845542 | !hmaster2_p & v1553138;
assign v1445a42 = hbusreq0 & v1445a3c | !hbusreq0 & v1445a41;
assign v1215d45 = hbusreq2_p & v1215d3c | !hbusreq2_p & v1215d44;
assign a653f3 = hmaster0_p & a653f0 | !hmaster0_p & a653d4;
assign v16a1bdd = hgrant2_p & v845542 | !hgrant2_p & v16a1bdc;
assign v155350d = hgrant3_p & v155321c | !hgrant3_p & v155350c;
assign d30120 = hmaster1_p & d3011f | !hmaster1_p & d3010e;
assign d306b7 = hmaster1_p & d306a9 | !hmaster1_p & d306b6;
assign v1446614 = hgrant1_p & v1446423 | !hgrant1_p & v1446600;
assign v1214dd0 = hmaster1_p & v1214dcf | !hmaster1_p & v845542;
assign v138a398 = hmaster0_p & v138a394 | !hmaster0_p & v138a34b;
assign f2f40a = hbusreq2 & f2f406 | !hbusreq2 & f2f409;
assign v1445e5f = hbusreq4_p & v14465c8 | !hbusreq4_p & v14465d6;
assign v1216272 = hbusreq3 & v1216271 | !hbusreq3 & !v1216030;
assign v1215ca3 = hbusreq1_p & v1215ca2 | !hbusreq1_p & !v845542;
assign v1446015 = hmaster2_p & v1446012 | !hmaster2_p & v1446014;
assign v1516105 = hbusreq2 & v15160fc | !hbusreq2 & v1516104;
assign v121607d = hbusreq3 & v1216070 | !hbusreq3 & v121607c;
assign v16a1adc = hmaster2_p & v16a1adb | !hmaster2_p & v16a206f;
assign v12153af = hbusreq2_p & v12153ae | !hbusreq2_p & v12153ad;
assign v1446276 = hlock2 & v1446275 | !hlock2 & v1446270;
assign f2f21e = hbusreq1 & v84556a | !hbusreq1 & v845542;
assign v12ad539 = hbusreq2_p & v12ad534 | !hbusreq2_p & v12ad538;
assign v1215448 = hmaster0_p & v12153ee | !hmaster0_p & v12153f3;
assign v1445dc2 = hmaster0_p & v1445d93 | !hmaster0_p & v1445d9d;
assign v121544d = hmaster1_p & v1215443 | !hmaster1_p & v121540f;
assign v14462f2 = hgrant5_p & v14465df | !hgrant5_p & v14462f1;
assign v14459ba = hbusreq0_p & v144640c | !hbusreq0_p & v1446406;
assign v12160fa = hbusreq4_p & v1216523 | !hbusreq4_p & !v845542;
assign d3013c = hlock5_p & d30139 | !hlock5_p & !d3013b;
assign v144549c = hlock3 & v1445492 | !hlock3 & v144549b;
assign v1446444 = hbusreq1 & v144640c | !hbusreq1 & v144640e;
assign f2f239 = hmaster1_p & f2f22c | !hmaster1_p & f2f238;
assign v1214c70 = hgrant5_p & v1215355 | !hgrant5_p & v1214c6f;
assign v16a1aca = hmaster1_p & v16a1ac9 | !hmaster1_p & !v16a1f96;
assign v16a12f1 = hbusreq2 & v16a12ef | !hbusreq2 & !v16a12f0;
assign v12ad530 = hmaster2_p & v12ad514 | !hmaster2_p & a658dc;
assign v1215d05 = hmaster1_p & v1215d04 | !hmaster1_p & v1215cfa;
assign f2ed90 = decide_p & f2f4bf | !decide_p & v845542;
assign v11e593c = hmaster0_p & v11e593b | !hmaster0_p & v845542;
assign v1214cd0 = hbusreq5_p & v1214ccc | !hbusreq5_p & !v1214ccf;
assign v16a1ca6 = hgrant2_p & v16a205b | !hgrant2_p & v16a1ca5;
assign v12ad4f7 = hbusreq1_p & v10d3fd8 | !hbusreq1_p & !v12ad4f6;
assign v1214f13 = hlock5_p & v1214f12 | !hlock5_p & !v1214ef2;
assign d30204 = hlock1_p & d306db | !hlock1_p & d30203;
assign v15161d0 = hmaster2_p & v845570 | !hmaster2_p & v15168f4;
assign v12ad039 = decide_p & v12acfee | !decide_p & !v12afe76;
assign v1214d46 = hbusreq4_p & v12153a5 | !hbusreq4_p & v845547;
assign a65640 = hbusreq0 & a6563a | !hbusreq0 & a6563f;
assign a65912 = hmaster2_p & a658be | !hmaster2_p & !a658ce;
assign d307ef = hgrant5_p & d306e3 | !hgrant5_p & d307ee;
assign d2faec = hbusreq1_p & d300c3 | !hbusreq1_p & d2faeb;
assign d2fb87 = hmaster1_p & d2fb86 | !hmaster1_p & d2fb7b;
assign v16a13e1 = hbusreq0 & v16a2078 | !hbusreq0 & v16a2087;
assign v1515ae9 = hmaster0_p & a6587e | !hmaster0_p & v1515ae8;
assign v1446180 = hlock2 & v144617b | !hlock2 & v144617f;
assign f2f434 = hgrant1_p & f2f281 | !hgrant1_p & !f2f389;
assign d2fc04 = hmaster2_p & d2fb4d | !hmaster2_p & d2fc03;
assign v15157ee = hlock5_p & v15157ec | !hlock5_p & !v15157ed;
assign v1515625 = hburst0 & v1552d7a | !hburst0 & v1515624;
assign a653d1 = hmaster2_p & a6628b | !hmaster2_p & a653d0;
assign d30232 = hmaster0_p & v845542 | !hmaster0_p & d30231;
assign v1445aa9 = hlock3 & v1445a69 | !hlock3 & v1445aa8;
assign v1445def = hbusreq1_p & v1446403 | !hbusreq1_p & v1445dee;
assign v1668c74 = hmaster2_p & a658ad | !hmaster2_p & !a658c6;
assign v1216212 = hgrant1_p & v845542 | !hgrant1_p & v1216211;
assign v16a129f = hmaster1_p & v16a1a97 | !hmaster1_p & !v16a2672;
assign v1668d7c = hgrant1_p & v1668d75 | !hgrant1_p & v1668d7b;
assign bf1f7c = hgrant1_p & v84556a | !hgrant1_p & !bf1f78;
assign v1668c1d = hmaster2_p & v845570 | !hmaster2_p & !v1668c1c;
assign v1214dd6 = hmaster0_p & v1216a78 | !hmaster0_p & v845542;
assign v16a1d57 = hbusreq3 & v16a1d51 | !hbusreq3 & v16a1d56;
assign v12161ae = hmaster0_p & v12161ad | !hmaster0_p & v121619b;
assign v1284d53 = hmaster1_p & v1284d45 | !hmaster1_p & !v1284cfd;
assign v144644f = hmaster0_p & v144639c | !hmaster0_p & v144643e;
assign v1668dd2 = hmaster0_p & v1668dca | !hmaster0_p & v1668dd1;
assign v1214eb8 = hbusreq2_p & v1214eb7 | !hbusreq2_p & v845542;
assign v16a19e4 = hmaster0_p & v16a19df | !hmaster0_p & v16a19d3;
assign v1515703 = hlock2_p & v1515701 | !hlock2_p & !v1515702;
assign v1214f51 = hbusreq2_p & v1214f50 | !hbusreq2_p & v12164e7;
assign v151572d = hgrant1_p & v1668d23 | !hgrant1_p & v151572c;
assign d30716 = hburst1 & d30715 | !hburst1 & v845542;
assign v1405ab9 = hbusreq2_p & v1405ab8 | !hbusreq2_p & v1405ab6;
assign v1668ca1 = hmaster0_p & v1668ca0 | !hmaster0_p & !v1668c7c;
assign v1445506 = hmaster0_p & v1445505 | !hmaster0_p & v1445414;
assign v1216589 = hmaster2_p & v1216588 | !hmaster2_p & v16a1bc6;
assign v1552d63 = hgrant2_p & v1552d54 | !hgrant2_p & v1552d61;
assign v1445921 = hlock2 & v144591e | !hlock2 & v1445920;
assign v1214dca = hbusreq3_p & v1214d34 | !hbusreq3_p & v1214dc9;
assign v1515adf = hmaster0_p & v845570 | !hmaster0_p & v166939c;
assign v1445da7 = hmaster2_p & v144639c | !hmaster2_p & v14463b9;
assign v15160fe = hlock4_p & v15160fd | !hlock4_p & v16693aa;
assign d80767 = hmaster0_p & v845542 | !hmaster0_p & d80734;
assign v151576f = hbusreq4_p & v151576c | !hbusreq4_p & v151576e;
assign v1445b03 = hmaster0_p & v1445a6b | !hmaster0_p & v1445902;
assign d301e6 = hbusreq1 & v845542 | !hbusreq1 & !d306f3;
assign v1284d56 = hmaster1_p & v1284d55 | !hmaster1_p & v140584d;
assign v144624d = hbusreq5_p & v14463dc | !hbusreq5_p & v144624c;
assign v16a1842 = hmaster2_p & v16a183f | !hmaster2_p & !v845542;
assign v1216aac = hmastlock_p & a66272 | !hmastlock_p & !v845542;
assign v10d42a4 = hmaster2_p & v10d4285 | !hmaster2_p & v10d4298;
assign v1445ead = hmaster2_p & v144639c | !hmaster2_p & v1445e70;
assign v1214ec0 = hbusreq5 & v1214eb9 | !hbusreq5 & v1214ebd;
assign v1668c4d = hbusreq1_p & v1668c2d | !hbusreq1_p & !v845542;
assign v1405b36 = hmaster1_p & v1405b35 | !hmaster1_p & !v1405a94;
assign v138a318 = hmaster1_p & v138a317 | !hmaster1_p & v138a314;
assign v12164dd = hbusreq0_p & v845570 | !hbusreq0_p & v12164cf;
assign f2f422 = hgrant1_p & f2f281 | !hgrant1_p & !f2f354;
assign d30192 = hbusreq2 & d30189 | !hbusreq2 & d30191;
assign d30116 = hgrant5_p & d2fea4 | !hgrant5_p & !d30114;
assign v1215414 = hmaster1_p & v12153f4 | !hmaster1_p & v121540f;
assign v1445a19 = hbusreq1 & v1445a14 | !hbusreq1 & v1445a18;
assign v1445a5f = hlock2 & v1445a47 | !hlock2 & v1445a5e;
assign v1214c97 = hmaster0_p & v1214c88 | !hmaster0_p & v1214c96;
assign v138a38f = hbusreq5_p & v138a38e | !hbusreq5_p & !v845542;
assign v1445ed1 = hlock2 & v1445ebe | !hlock2 & v1445ed0;
assign v121615e = hbusreq1 & v121615d | !hbusreq1 & v845542;
assign v1553156 = hmaster1_p & v1553155 | !hmaster1_p & v155314e;
assign v16a13cd = hmaster1_p & v16a13a8 | !hmaster1_p & !v16a1f96;
assign d2fc6a = hgrant5_p & d2fc24 | !hgrant5_p & d2fc69;
assign v16a12e9 = hgrant4_p & v845559 | !hgrant4_p & v16a12e8;
assign v134d4c4 = decide_p & v134d3ce | !decide_p & v134d3b5;
assign v1445ea8 = hbusreq0 & v1445ea0 | !hbusreq0 & v1445ea7;
assign a65927 = hbusreq2 & a65923 | !hbusreq2 & a65926;
assign d3060d = hmaster0_p & d305ed | !hmaster0_p & d3060c;
assign v1445dea = hbusreq4_p & v144640c | !hbusreq4_p & v1446406;
assign f2f2aa = hbusreq1_p & f2f2a9 | !hbusreq1_p & v845542;
assign d807a1 = hmaster1_p & d807a0 | !hmaster1_p & v845542;
assign d2f975 = hmaster0_p & d2f970 | !hmaster0_p & d2f974;
assign v12ad5d1 = hbusreq1 & v12ad4fc | !hbusreq1 & !v845542;
assign v121544c = hbusreq2 & v1215447 | !hbusreq2 & v121544b;
assign v16a1890 = hbusreq5 & v16a1888 | !hbusreq5 & v16a188f;
assign v12ae1fc = hmaster2_p & v12afe62 | !hmaster2_p & v12ae1fb;
assign v1405924 = hmaster1_p & v1405923 | !hmaster1_p & v140584d;
assign v144608c = hmaster1_p & v144608b | !hmaster1_p & v1445fde;
assign v12ad31e = hmaster2_p & v12af9c1 | !hmaster2_p & v12ad31d;
assign v1445d9b = hbusreq1 & v1445d98 | !hbusreq1 & v1445d9a;
assign v1214f70 = hbusreq2_p & v1214f6f | !hbusreq2_p & v12164e7;
assign a654ab = hbusreq2 & a65498 | !hbusreq2 & a654a9;
assign d300ed = hgrant1_p & d300da | !hgrant1_p & d300c3;
assign v12ad65e = hmaster0_p & v12ad5f8 | !hmaster0_p & v845542;
assign v144639d = stateA1_p & v146d169 | !stateA1_p & !v845588;
assign v1446150 = hbusreq2 & v144614e | !hbusreq2 & v144614f;
assign v16a13a8 = hmaster2_p & v16a13a7 | !hmaster2_p & v845542;
assign v16a1d98 = hmaster1_p & v16a1d8c | !hmaster1_p & v16a1f96;
assign v134d4ad = hlock0 & v134d4ac | !hlock0 & v134d4ab;
assign v12161d2 = hmaster2_p & v12161d0 | !hmaster2_p & v12161d1;
assign d30237 = hbusreq2_p & d30235 | !hbusreq2_p & d30236;
assign v12ad665 = hbusreq0 & v12ad664 | !hbusreq0 & !v12af73f;
assign v1515734 = hgrant5_p & v151560b | !hgrant5_p & v1515733;
assign v1445769 = hbusreq2_p & v1445767 | !hbusreq2_p & v1445768;
assign bf1f88 = decide_p & v84556a | !decide_p & bf1f87;
assign v16a1cbe = hgrant2_p & v16a2060 | !hgrant2_p & v16a1cbd;
assign v1215081 = hmaster1_p & v1215066 | !hmaster1_p & !v121507b;
assign v1215088 = hgrant2_p & v1215059 | !hgrant2_p & v1215087;
assign d2fe9a = hlock4_p & v845580 | !hlock4_p & v845542;
assign v1214ee1 = hgrant5_p & v845547 | !hgrant5_p & v1214edf;
assign d80751 = hbusreq2_p & d80750 | !hbusreq2_p & d8074f;
assign bf1f7a = hmaster2_p & v84556a | !hmaster2_p & !bf1f79;
assign v138a02e = hbusreq5_p & v138a02d | !hbusreq5_p & v845542;
assign f2f344 = hmaster1_p & f2f343 | !hmaster1_p & f2f2a2;
assign d3068a = hmaster2_p & d30689 | !hmaster2_p & !v845542;
assign v1215ce3 = hbusreq5_p & v1215ce2 | !hbusreq5_p & v1215c88;
assign v1566987 = stateG3_2_p & v845542 | !stateG3_2_p & !v893df7;
assign v1515804 = hgrant2_p & v15167ff | !hgrant2_p & !v1515803;
assign d3015f = hgrant2_p & v84555a | !hgrant2_p & d3015b;
assign v1445ebd = hgrant2_p & v1445eb2 | !hgrant2_p & v1445ebc;
assign v1445a2f = hgrant5_p & v14458f9 | !hgrant5_p & v1445a2e;
assign v12ad0bc = hlock2_p & v12ad0b5 | !hlock2_p & v12ad0bb;
assign d2fb8f = hmaster0_p & d2fb8c | !hmaster0_p & d2fb7e;
assign d30742 = hlock1_p & d30741 | !hlock1_p & !d305ef;
assign v134cec3 = hbusreq2_p & v134d49c | !hbusreq2_p & v134d3b5;
assign v121574d = hgrant5_p & v1215731 | !hgrant5_p & v121574c;
assign d3094c = stateA1_p & v146af2e | !stateA1_p & d3094b;
assign v14454ef = hlock0 & v14454ee | !hlock0 & v14454eb;
assign v12147e9 = hbusreq2 & v12147e8 | !hbusreq2 & v845542;
assign v121613f = hgrant4_p & v121613d | !hgrant4_p & v121613e;
assign v16a13d6 = hbusreq2 & v16a13d5 | !hbusreq2 & !v16a1f9b;
assign v12acfce = hmaster0_p & v12ad536 | !hmaster0_p & v12ad52d;
assign v134d367 = hgrant1_p & v845542 | !hgrant1_p & v134d366;
assign v121601e = hmaster2_p & v121601c | !hmaster2_p & !v121601d;
assign v16a1bc8 = hgrant4_p & v845559 | !hgrant4_p & !v16a1bc7;
assign v1214d72 = decide_p & v1214d6c | !decide_p & v1214d71;
assign v16a1412 = hbusreq3 & v16a140c | !hbusreq3 & v16a1411;
assign v1216221 = hmaster2_p & v1216218 | !hmaster2_p & v1216220;
assign d2fb46 = hbusreq2 & d2fb44 | !hbusreq2 & d2fb45;
assign v121534f = hbusreq1_p & v121534b | !hbusreq1_p & v1215345;
assign v1445428 = hmaster1_p & v1445414 | !hmaster1_p & v1445b5f;
assign v1445eec = hgrant5_p & v1445ee9 | !hgrant5_p & v1445eeb;
assign v11e594d = hmaster2_p & v845542 | !hmaster2_p & !v11e594c;
assign d30278 = hlock5_p & d30276 | !hlock5_p & !d30277;
assign v1446689 = hlock1 & v14465be | !hlock1 & v14465c4;
assign f2f3ca = hbusreq5_p & f2f3c8 | !hbusreq5_p & !f2f3c9;
assign v1446621 = hmaster2_p & v14465f5 | !hmaster2_p & v1446620;
assign d30605 = hlock5_p & v845542 | !hlock5_p & d30604;
assign v1215ff5 = stateA1_p & v88d3e4 | !stateA1_p & v845542;
assign v1215c6f = hgrant5_p & v845542 | !hgrant5_p & v1215c3d;
assign v140583d = locked_p & v1405839 | !locked_p & v140583c;
assign v134d4b1 = hgrant2_p & v134d4a2 | !hgrant2_p & v134d4af;
assign d8079b = hgrant5_p & v845542 | !hgrant5_p & d8079a;
assign v10d3fdc = hmaster2_p & v10d3fd5 | !hmaster2_p & v10d3fdb;
assign v12153d0 = hbusreq4 & v1216aad | !hbusreq4 & v12153cf;
assign v1215342 = hready_p & v121531d | !hready_p & v1215341;
assign d306cd = hbusreq1_p & d306cc | !hbusreq1_p & v845542;
assign v144580a = hmaster0_p & v1445ecc | !hmaster0_p & v1445eba;
assign d2facd = hmaster0_p & d2fe8e | !hmaster0_p & d2fe7e;
assign v1446310 = hgrant5_p & v144643d | !hgrant5_p & v144630c;
assign a662bd = hgrant3_p & a66281 | !hgrant3_p & a662bc;
assign v1445aad = decide_p & v14458d1 | !decide_p & v1445aac;
assign v1445b1e = hlock3 & v1445b15 | !hlock3 & v1445b1d;
assign v144660b = hlock0_p & v144639c | !hlock0_p & v144660a;
assign v12af1c2 = hbusreq2_p & v12af3ac | !hbusreq2_p & v12af1c1;
assign v1668d80 = hgrant5_p & v1668d7f | !hgrant5_p & v1668d7d;
assign d2fd3e = hbusreq2 & d2fd3c | !hbusreq2 & d2fd3d;
assign v1216a9b = hmaster0_p & v1216a95 | !hmaster0_p & v1216a9a;
assign v1215ffe = hbusreq1 & v1215ffd | !hbusreq1 & v845542;
assign a65adb = hgrant2_p & v845542 | !hgrant2_p & a65ada;
assign v12ae83d = jx2_p & v12aee5f | !jx2_p & v12ae83c;
assign v121572f = hbusreq5_p & v121572d | !hbusreq5_p & !v121572e;
assign v1215be0 = hbusreq5_p & v1215bde | !hbusreq5_p & v1215bdf;
assign d2fc56 = hgrant1_p & d2fbcb | !hgrant1_p & d2fc55;
assign f2f392 = hbusreq0 & f2f387 | !hbusreq0 & f2f391;
assign d3071d = hbusreq1_p & d3071c | !hbusreq1_p & v845542;
assign v16a1c00 = hmaster1_p & v16a1bfc | !hmaster1_p & v16a1bff;
assign v12ad569 = hmaster0_p & v12ad565 | !hmaster0_p & v12ad52d;
assign v1216791 = hmaster1_p & v1216790 | !hmaster1_p & v1216a9b;
assign v12ae1f9 = hbusreq4_p & v12ae1f8 | !hbusreq4_p & v12afe60;
assign v12ad612 = hbusreq0 & v12ad611 | !hbusreq0 & !v12afe63;
assign v1446706 = hmaster1_p & v1446705 | !hmaster1_p & v1446436;
assign v134d3bf = hbusreq0_p & v134d1e8 | !hbusreq0_p & v845542;
assign d301b7 = hbusreq5 & d30197 | !hbusreq5 & d301b6;
assign v1445f06 = hbusreq5_p & v1445e6e | !hbusreq5_p & v1445f05;
assign d2fcb4 = hbusreq0 & d305fc | !hbusreq0 & d30604;
assign v12ae209 = decide_p & v12ae201 | !decide_p & v12afe76;
assign v14461bd = hmaster1_p & v144617c | !hmaster1_p & v1445ffc;
assign v16a1d67 = hbusreq3 & v16a1d66 | !hbusreq3 & v16a209f;
assign v14058a6 = hlock4_p & v140583f | !hlock4_p & v1405854;
assign v1405920 = hmaster0_p & v14058bb | !hmaster0_p & v1405896;
assign d80754 = hburst1_p & v845542 | !hburst1_p & d80753;
assign v16a1ce7 = hbusreq5 & v16a1cdb | !hbusreq5 & v16a1ce6;
assign v16a197c = hbusreq0 & v16a209a | !hbusreq0 & v16a197b;
assign v1445b32 = hmaster1_p & v1445b31 | !hmaster1_p & v14458fd;
assign v15533ad = hgrant4_p & v845542 | !hgrant4_p & v15533ac;
assign v14453e9 = hbusreq3 & v14453e7 | !hbusreq3 & v14453e8;
assign v1445459 = hlock2 & v1445446 | !hlock2 & v1445458;
assign v1215c7b = hbusreq5 & v1215c52 | !hbusreq5 & v1215c7a;
assign v14058aa = hbusreq0_p & v1405854 | !hbusreq0_p & v140589a;
assign v1216238 = hmaster1_p & v1216237 | !hmaster1_p & v1216224;
assign v1446419 = hlock0 & v1446418 | !hlock0 & v1446414;
assign v1445ba4 = hbusreq3 & v1445ba3 | !hbusreq3 & v1445b86;
assign v1668d8d = hgrant2_p & v1668d1f | !hgrant2_p & v1668d8c;
assign v15533a3 = hmaster2_p & v155339f | !hmaster2_p & v15533a2;
assign v140591a = hready_p & v1405910 | !hready_p & v1405919;
assign v1214c99 = hgrant2_p & v121536e | !hgrant2_p & v1214c98;
assign v1445a4c = hbusreq1 & v14459b6 | !hbusreq1 & v14459b7;
assign v1405918 = hbusreq2_p & v1405879 | !hbusreq2_p & v1405917;
assign v10d4012 = decide_p & v10d4009 | !decide_p & v10d4011;
assign v16a1e01 = hbusreq2 & v16a1dff | !hbusreq2 & v16a1e00;
assign v12af98c = hbusreq0 & v12af987 | !hbusreq0 & v12af98b;
assign v134ce5e = hmaster2_p & v134ce52 | !hmaster2_p & v845542;
assign v14463f9 = hbusreq2_p & v14463f0 | !hbusreq2_p & v14463f8;
assign v151570e = hready_p & v1515646 | !hready_p & v151570d;
assign v144628d = hbusreq5_p & v1446411 | !hbusreq5_p & v144628c;
assign v1214fb8 = hlock4_p & v1215765 | !hlock4_p & v1214fb7;
assign v155305a = hbusreq1 & v1553058 | !hbusreq1 & v1553059;
assign v1216a96 = hbusreq4_p & v16a1bc6 | !hbusreq4_p & v845570;
assign v1405895 = hlock5_p & v1405893 | !hlock5_p & v1405894;
assign v12ad5cf = hbusreq0 & v12ad5ce | !hbusreq0 & v12afe63;
assign v134d515 = hgrant2_p & v134d364 | !hgrant2_p & v134d514;
assign v1215465 = hbusreq4 & v12164cf | !hbusreq4 & v845542;
assign v1215b7a = hlock4_p & v1215b78 | !hlock4_p & v1215b79;
assign v138a3e9 = hgrant5_p & v845570 | !hgrant5_p & !v1515837;
assign v10d40d9 = hgrant2_p & v10d40d7 | !hgrant2_p & v10d40d8;
assign v16a1aea = hgrant2_p & v845542 | !hgrant2_p & !v16a1ae9;
assign v1215457 = hmaster1_p & v121543b | !hmaster1_p & v121540f;
assign v1445ff9 = hbusreq5_p & v1445fcb | !hbusreq5_p & v1445ff8;
assign v1515844 = hbusreq5_p & v1515842 | !hbusreq5_p & !v1515843;
assign v12af223 = hgrant1_p & d30690 | !hgrant1_p & v12af222;
assign a65af1 = hmaster0_p & a65ae9 | !hmaster0_p & a65af0;
assign f2f372 = hbusreq1 & v1668d58 | !hbusreq1 & v845542;
assign d30883 = hmaster1_p & d30882 | !hmaster1_p & d307f4;
assign v1446125 = hbusreq2_p & v1446122 | !hbusreq2_p & v1446124;
assign v14458e8 = hbusreq1 & v14458db | !hbusreq1 & v14458e7;
assign d2fb33 = decide_p & d2fb32 | !decide_p & v845570;
assign v1446286 = hbusreq2_p & v144627f | !hbusreq2_p & v1446285;
assign d30864 = hmaster2_p & d30863 | !hmaster2_p & d30654;
assign v12aec4f = decide_p & v12aec4e | !decide_p & v12afe76;
assign v1214d7a = hmaster1_p & v1214c7b | !hmaster1_p & v1214c74;
assign v1445b39 = hgrant2_p & v1445b37 | !hgrant2_p & v1445b38;
assign d302d9 = hmaster0_p & d302d7 | !hmaster0_p & d302d8;
assign v138a361 = hlock2_p & v138a35e | !hlock2_p & v138a360;
assign v1445bac = decide_p & v1445bab | !decide_p & v144639b;
assign v12160a8 = hmaster0_p & v121605f | !hmaster0_p & v121606b;
assign d306e3 = hmaster2_p & d306dd | !hmaster2_p & d306e2;
assign v1216a71 = hmaster0_p & v1216a70 | !hmaster0_p & v1216a6c;
assign v14459a9 = hlock4 & v144639c | !hlock4 & v14459a8;
assign v1445a10 = hbusreq0_p & v1445a0f | !hbusreq0_p & v144639e;
assign v12aead3 = decide_p & v12af1c2 | !decide_p & v12afe76;
assign v1214eed = hmaster1_p & v1214ed8 | !hmaster1_p & v1214eec;
assign v1445bc6 = hmaster0_p & v845542 | !hmaster0_p & v14464a5;
assign v1668dbf = hbusreq5_p & v1668dbd | !hbusreq5_p & !v1668dbe;
assign d8075a = busreq_p & d80758 | !busreq_p & !d80759;
assign v144541b = hgrant2_p & v1445418 | !hgrant2_p & v144541a;
assign f2f222 = hmaster0_p & f2f221 | !hmaster0_p & v845542;
assign v1215441 = hbusreq3 & v1215417 | !hbusreq3 & v1215440;
assign v1216a65 = stateA1_p & v845542 | !stateA1_p & v1216a64;
assign d2f996 = hmaster1_p & d2fef8 | !hmaster1_p & d2f995;
assign v1668da9 = hmaster1_p & v1668da8 | !hmaster1_p & v845570;
assign v1445479 = hmaster0_p & v1445473 | !hmaster0_p & v1446404;
assign v16a1e6a = hbusreq2_p & v16a1dc0 | !hbusreq2_p & v16a1e69;
assign d30135 = hlock5_p & d30133 | !hlock5_p & d30134;
assign v1515ae6 = hlock4_p & v1515ae4 | !hlock4_p & !v1515ae5;
assign v140584a = hbusreq0_p & v14463b1 | !hbusreq0_p & v1405844;
assign v1214cc0 = hgrant5_p & v121537d | !hgrant5_p & v1214cbf;
assign v1445f13 = hgrant2_p & v1445ef7 | !hgrant2_p & v1445f12;
assign v1405894 = hgrant5_p & v1405856 | !hgrant5_p & v1405892;
assign v1214cf0 = hmaster2_p & v1214c2a | !hmaster2_p & v1214c31;
assign v144631d = hmaster0_p & v14462e6 | !hmaster0_p & v144631c;
assign v134ce54 = hbusreq0 & v134ce53 | !hbusreq0 & v134d274;
assign v10d4287 = hmastlock_p & v10d4286 | !hmastlock_p & v845580;
assign v12ad012 = hgrant1_p & v12ad5d2 | !hgrant1_p & v12ad011;
assign bf1f79 = hgrant1_p & bf1f52 | !hgrant1_p & bf1f78;
assign v121654d = hlock5_p & v121654c | !hlock5_p & v1216547;
assign v1445bae = stateG10_5_p & v1445f89 | !stateG10_5_p & !v14463a6;
assign v14466a2 = hgrant5_p & v1446426 | !hgrant5_p & v14466a1;
assign v14459a4 = hmaster2_p & v144639c | !hmaster2_p & v14458e5;
assign v10d4068 = hbusreq1_p & v10d4061 | !hbusreq1_p & v10d4067;
assign v14461d5 = hbusreq2_p & v14461c4 | !hbusreq2_p & v14461d4;
assign v12160db = hbusreq1 & v12164dc | !hbusreq1 & v845542;
assign v14459ed = hmaster2_p & v14459ec | !hmaster2_p & v14459e7;
assign v14058d3 = hgrant0_p & v14058d2 | !hgrant0_p & v140584b;
assign v12ad034 = hbusreq2 & v12ad030 | !hbusreq2 & v12ad033;
assign v14465bd = hlock4 & v144639c | !hlock4 & v14465bc;
assign v1445f4e = hlock2 & v1445f4b | !hlock2 & v1445f4d;
assign v134d4fb = hbusreq4_p & v134d273 | !hbusreq4_p & v134d36d;
assign v138a31a = hlock5_p & v151563f | !hlock5_p & v845542;
assign v1405b64 = hready_p & v1405b5a | !hready_p & v1405b63;
assign v11e596a = hgrant5_p & v845542 | !hgrant5_p & v11e5969;
assign v12162dd = hbusreq2 & v12162d2 | !hbusreq2 & v12162dc;
assign v16a19d0 = hbusreq4_p & v16a183f | !hbusreq4_p & !v845542;
assign f2f3c2 = hgrant5_p & f2f3c1 | !hgrant5_p & f2f36a;
assign v140589f = hmaster2_p & v1405854 | !hmaster2_p & v1405845;
assign v12ad56b = hmaster0_p & v12ad565 | !hmaster0_p & v12ad531;
assign v121628d = hgrant2_p & v1216187 | !hgrant2_p & v1216286;
assign v12acfe5 = hmaster1_p & v12acfcb | !hmaster1_p & v12acfdb;
assign v1446176 = hgrant2_p & v1446173 | !hgrant2_p & v1446175;
assign v14058b3 = hgrant2_p & v1405887 | !hgrant2_p & v14058b2;
assign d30821 = hlock5_p & d3081f | !hlock5_p & !d30820;
assign v1445b7a = hmaster0_p & v1445b79 | !hmaster0_p & v1446340;
assign v151560e = hbusreq1_p & a65851 | !hbusreq1_p & v151560d;
assign v1552d83 = hbusreq5_p & v1552d80 | !hbusreq5_p & v1552d82;
assign v144579c = hbusreq0 & v144579b | !hbusreq0 & v1445776;
assign v12162e8 = hmaster2_p & v1216048 | !hmaster2_p & v845542;
assign v121571f = hbusreq4_p & v121571e | !hbusreq4_p & v845542;
assign f2e4e3 = jx2_p & f2e4c9 | !jx2_p & f2e4e2;
assign v144611c = hbusreq2_p & v1446119 | !hbusreq2_p & v144611b;
assign v144626a = hmaster0_p & v1446267 | !hmaster0_p & v1446269;
assign v1668ddc = hbusreq5_p & v1668dda | !hbusreq5_p & !v1668ddb;
assign v155343a = hbusreq4_p & v1553220 | !hbusreq4_p & v1553439;
assign v1552d4e = hgrant2_p & v1553380 | !hgrant2_p & v1552d4d;
assign v1214c30 = hbusreq0_p & v12164cf | !hbusreq0_p & v845542;
assign v12150f6 = hbusreq2_p & v12150f5 | !hbusreq2_p & v12150f1;
assign d3078d = locked_p & d3078c | !locked_p & !v845542;
assign v12aeb1a = hmaster0_p & v845542 | !hmaster0_p & v12aeb19;
assign v1445e2a = hmaster1_p & v1445e0d | !hmaster1_p & v1445e28;
assign v1445a2c = hbusreq1 & v1445a2a | !hbusreq1 & v1445a2b;
assign v134d1f7 = hlock1_p & v134d1f6 | !hlock1_p & v845542;
assign v144576c = hlock2 & v1445769 | !hlock2 & v144576b;
assign v1214f6a = hbusreq2 & v1214f69 | !hbusreq2 & v845542;
assign v138a344 = hbusreq5_p & v138a343 | !hbusreq5_p & !v845542;
assign d302f4 = decide_p & d302f3 | !decide_p & v845570;
assign v16a13d1 = hbusreq2 & v16a13d0 | !hbusreq2 & v16a1f98;
assign v134cd44 = jx2_p & v134d4c7 | !jx2_p & v134d541;
assign v12166e5 = hready & v12166e4 | !hready & !v845542;
assign v14465da = hbusreq1_p & v14465b2 | !hbusreq1_p & v14465d7;
assign v1214ccf = hgrant5_p & v1214ccd | !hgrant5_p & !v1214cce;
assign f2f3e6 = hmaster0_p & f2f396 | !hmaster0_p & f2f350;
assign v15534f4 = hlock2 & v15534dd | !hlock2 & v15534f3;
assign v1446214 = hbusreq5_p & v144639c | !hbusreq5_p & v1446213;
assign v12164e4 = hmaster0_p & v12164d5 | !hmaster0_p & v12164e3;
assign v144633e = hlock0 & v144633d | !hlock0 & v144633c;
assign v15157bc = hgrant4_p & v15157bb | !hgrant4_p & v845570;
assign f2f2e8 = hmaster2_p & f2f2c9 | !hmaster2_p & !f2f2e7;
assign v1446211 = hmaster2_p & v14463b1 | !hmaster2_p & !v144639c;
assign v144537a = hmaster1_p & v1445b33 | !hmaster1_p & v1445a82;
assign v121670a = hgrant2_p & v12166c2 | !hgrant2_p & v1216709;
assign hmaster1 = v143fd7d;
assign v1405931 = hmaster1_p & v1405930 | !hmaster1_p & v14058b1;
assign v15156bb = hgrant1_p & v15156ba | !hgrant1_p & v1515654;
assign v1216013 = hmastlock_p & v1515618 | !hmastlock_p & v845542;
assign a65403 = hmaster0_p & a6538f | !hmaster0_p & a65401;
assign v1405886 = hmaster1_p & v1405885 | !hmaster1_p & v140584d;
assign v14458a3 = hbusreq0 & v14458a1 | !hbusreq0 & v14458a2;
assign v14466ab = hgrant2_p & v14465ab | !hgrant2_p & v14466aa;
assign v16a207e = hgrant1_p & v84554d | !hgrant1_p & v16a207d;
assign v1445eb7 = hmaster2_p & v144639c | !hmaster2_p & v1445e80;
assign f2f36e = hgrant5_p & f2f363 | !hgrant5_p & f2f36a;
assign v16a1ad7 = hready_p & v845555 | !hready_p & !v16a1ad6;
assign v121622b = hgrant5_p & v12160e2 | !hgrant5_p & v121622a;
assign v1216109 = hlock1_p & v1216106 | !hlock1_p & v1216108;
assign d2fae4 = hgrant5_p & d2f973 | !hgrant5_p & !d2fae3;
assign v1445e8b = hgrant4_p & v1445e89 | !hgrant4_p & v1445e8a;
assign v12ad502 = hbusreq0 & v12ad501 | !hbusreq0 & v845542;
assign v1445ee2 = hgrant2_p & v1445ee1 | !hgrant2_p & v1445ece;
assign v1215450 = hbusreq2_p & v121544f | !hbusreq2_p & v121544e;
assign v1553442 = hgrant2_p & v845542 | !hgrant2_p & v1553441;
assign v16a1db2 = hmaster1_p & v16a1db1 | !hmaster1_p & v16a1d53;
assign v16a1e57 = decide_p & v16a1dda | !decide_p & !v16a1e56;
assign v1215dad = hbusreq5 & v1215d95 | !hbusreq5 & v1215dac;
assign v1668c1c = locked_p & v1668c1b | !locked_p & v845542;
assign v155341d = hmaster1_p & v1553385 | !hmaster1_p & v155341c;
assign v1215d9d = hgrant2_p & v1215d69 | !hgrant2_p & v1215d9c;
assign v1215710 = hbusreq4 & v1216528 | !hbusreq4 & !v845547;
assign v1445432 = hbusreq3 & v1445430 | !hbusreq3 & v1445431;
assign v144544f = hbusreq2 & v1445445 | !hbusreq2 & v144544e;
assign v14454ec = hmaster2_p & v1445412 | !hmaster2_p & v1446645;
assign d2f97a = hbusreq1_p & d2fea1 | !hbusreq1_p & d2f979;
assign v1446082 = hmaster0_p & v144603f | !hmaster0_p & v1446081;
assign v134d378 = hmaster2_p & v845542 | !hmaster2_p & v134d377;
assign v1668c66 = hmaster2_p & a658c6 | !hmaster2_p & !v1668c64;
assign v14463ad = hbusreq1 & v14463ab | !hbusreq1 & v14463ac;
assign v121652d = hgrant4_p & v1216524 | !hgrant4_p & v121652c;
assign d305e3 = hmaster1_p & d305e2 | !hmaster1_p & d305db;
assign v138a357 = hbusreq2_p & v138a352 | !hbusreq2_p & v138a356;
assign a65b09 = hmaster0_p & a66287 | !hmaster0_p & a6629b;
assign v1215bc2 = hmaster0_p & v1215bc1 | !hmaster0_p & !v12163a8;
assign f2f232 = hgrant5_p & v845542 | !hgrant5_p & !f2f231;
assign f2f444 = hgrant2_p & f2f417 | !hgrant2_p & f2f443;
assign v140592f = hgrant5_p & v1405859 | !hgrant5_p & v140592e;
assign d3077a = hlock3_p & d30766 | !hlock3_p & d30779;
assign v1214c59 = hbusreq1 & v1215364 | !hbusreq1 & v845547;
assign v16a196a = hgrant2_p & v845542 | !hgrant2_p & !v16a1969;
assign v1389f98 = hbusreq2_p & v1389f8f | !hbusreq2_p & v1389f97;
assign v16a1963 = hgrant5_p & v845542 | !hgrant5_p & !v16a194c;
assign v1215fe5 = hready_p & v12167ac | !hready_p & v1215fe4;
assign d2f984 = hmaster1_p & d2f980 | !hmaster1_p & d2f983;
assign v12153d9 = hbusreq4_p & v12153d8 | !hbusreq4_p & v845542;
assign v1214c1c = hmaster1_p & v1214c07 | !hmaster1_p & v1214bcf;
assign v1446326 = hbusreq2_p & v1446301 | !hbusreq2_p & v1446325;
assign v1553219 = hmaster0_p & v1553218 | !hmaster0_p & v845542;
assign v15530a0 = hbusreq2 & v155309e | !hbusreq2 & v155309f;
assign v12ad5c0 = hbusreq4_p & v12ad5be | !hbusreq4_p & !v12ad5bf;
assign v14466ef = hbusreq5 & v14466d7 | !hbusreq5 & v14466ee;
assign v1445bb4 = hbusreq2_p & v1445bb2 | !hbusreq2_p & v1445bb3;
assign v1668d3d = hmaster2_p & v1668d2f | !hmaster2_p & v1668d3c;
assign v12acfef = decide_p & v12acfee | !decide_p & !v845542;
assign v1445ffb = hlock0 & v1445ffa | !hlock0 & v1445ff9;
assign d2fce9 = hmaster0_p & d2fce8 | !hmaster0_p & v16693aa;
assign v16a1cd7 = hbusreq2_p & v16a1b02 | !hbusreq2_p & v16a1cd6;
assign v16a188b = hbusreq2 & v16a1889 | !hbusreq2 & v16a188a;
assign d2fc27 = hmaster0_p & d2fc23 | !hmaster0_p & d2fc26;
assign v16a1e71 = hmaster1_p & v16a1e64 | !hmaster1_p & !v16a1f96;
assign v10d3fec = hmaster0_p & v10d3fda | !hmaster0_p & v10d3feb;
assign v1214e63 = hmaster1_p & v1214e62 | !hmaster1_p & !v12163a9;
assign v16a1da6 = hmaster1_p & v16a1acc | !hmaster1_p & v16a2672;
assign v16a140d = hmaster0_p & v16a1d91 | !hmaster0_p & v16a1d8c;
assign v1216088 = hmaster1_p & v121606c | !hmaster1_p & v1216082;
assign v16693ac = hmaster2_p & v845542 | !hmaster2_p & v16693ab;
assign v1446696 = hlock4 & v14465bc | !hlock4 & v14465bb;
assign v1445a63 = hgrant2_p & v1445a60 | !hgrant2_p & v1445a62;
assign v144619b = hbusreq3 & v1446199 | !hbusreq3 & v144619a;
assign a658b0 = hbusreq4_p & a658ad | !hbusreq4_p & v845542;
assign v16a13fd = hbusreq5 & v16a13ea | !hbusreq5 & v16a13fc;
assign v1552da1 = hbusreq3_p & v1552d99 | !hbusreq3_p & v1552da0;
assign v1445ae3 = hlock5 & v1445abf | !hlock5 & v1445ae1;
assign v12ad55e = hlock2_p & v12ad55c | !hlock2_p & v12ad55d;
assign v121578a = hbusreq2_p & v1215788 | !hbusreq2_p & v1215789;
assign d2fd12 = hbusreq2 & d2fd11 | !hbusreq2 & d2fcd8;
assign f2f38e = hmaster2_p & f2f38a | !hmaster2_p & f2f38d;
assign v1215c31 = hgrant5_p & v1215be1 | !hgrant5_p & v1215c30;
assign a658b7 = hmaster2_p & a658b0 | !hmaster2_p & a658b6;
assign d3070c = locked_p & v845580 | !locked_p & !v845542;
assign v1553503 = hlock2 & v1553500 | !hlock2 & v1553502;
assign d30166 = hmaster0_p & d30111 | !hmaster0_p & d2fe9b;
assign v10d40dc = hready_p & v10d40d0 | !hready_p & !v10d40db;
assign d308d3 = hbusreq3_p & d30847 | !hbusreq3_p & !d308d2;
assign v12af1bf = hbusreq0 & v12af1bb | !hbusreq0 & v12af1be;
assign v16a1ae8 = hbusreq0 & v16a1ae7 | !hbusreq0 & v16a209b;
assign v1515aec = hgrant2_p & v1515aeb | !hgrant2_p & !v845542;
assign v1214c2f = hmaster0_p & v1214c2c | !hmaster0_p & v1214c2e;
assign v1389e2d = hbusreq5_p & v1389e2c | !hbusreq5_p & !v845542;
assign v10d4053 = hmaster0_p & v10d3ff1 | !hmaster0_p & v10d4052;
assign d3077c = hready_p & d30713 | !hready_p & d3077b;
assign v1405b5d = hmaster0_p & v1405b2d | !hmaster0_p & v1405b16;
assign v1284cbd = hmaster0_p & v1284cb9 | !hmaster0_p & v1284cbc;
assign v1215358 = hmaster1_p & v121534e | !hmaster1_p & v1215357;
assign v1405abb = locked_p & v1405a86 | !locked_p & v1405aa2;
assign v16a1a2d = hbusreq2 & v16a1a2a | !hbusreq2 & v16a1a2c;
assign v1216a89 = stateG3_2_p & v845542 | !stateG3_2_p & v1216a88;
assign v1552f59 = hmaster2_p & v845542 | !hmaster2_p & v1552f58;
assign v1215d6e = hmaster0_p & v1215d6c | !hmaster0_p & v1215d6d;
assign v1446698 = hbusreq4_p & v144639c | !hbusreq4_p & v1446697;
assign a65372 = hgrant1_p & a65362 | !hgrant1_p & !a65371;
assign v1405a88 = locked_p & v1405a87 | !locked_p & !v845542;
assign v14460c0 = hbusreq2_p & v14460b8 | !hbusreq2_p & v14460bf;
assign d2fbf2 = hbusreq0 & d2fbf1 | !hbusreq0 & d302e0;
assign v10d42be = hready_p & v10d42aa | !hready_p & !v10d42bd;
assign d30813 = hbusreq2_p & d30811 | !hbusreq2_p & d30812;
assign v1445b13 = hlock2 & v1445b10 | !hlock2 & v1445b12;
assign v1216571 = hmaster2_p & v121655f | !hmaster2_p & v1216570;
assign v14458ee = hbusreq5_p & v14458ec | !hbusreq5_p & v14458ed;
assign v138953c = hmaster1_p & v845542 | !hmaster1_p & !v138953b;
assign v14463c2 = hmaster0_p & v14463aa | !hmaster0_p & v14463c1;
assign v12acfdb = hmaster0_p & v12acfda | !hmaster0_p & !v12acfb8;
assign v12ad57b = hmaster0_p & v12ad531 | !hmaster0_p & v12ad536;
assign v1445f5a = hmaster0_p & v1446448 | !hmaster0_p & v144667f;
assign v1446462 = hgrant0_p & v845542 | !hgrant0_p & v1446398;
assign d307ff = hmaster2_p & d307a0 | !hmaster2_p & d307bf;
assign d30913 = hmaster2_p & v845542 | !hmaster2_p & !d30911;
assign v1445dfa = hlock0 & v1445df9 | !hlock0 & v1445df4;
assign v15157e4 = hbusreq0 & v15157e0 | !hbusreq0 & v15157e3;
assign v1215096 = hbusreq1 & v1215038 | !hbusreq1 & v1215095;
assign v1668daf = hbusreq2_p & v1668daa | !hbusreq2_p & !v1668dae;
assign v16a1e55 = hbusreq3 & v16a1e4f | !hbusreq3 & v16a1e54;
assign v1214efa = hmaster0_p & v1214ef4 | !hmaster0_p & v1214ef9;
assign a66272 = stateG2_p & v845542 | !stateG2_p & !v156645f;
assign v1216545 = hlock1_p & v1216544 | !hlock1_p & !v845542;
assign v140585d = hlock3_p & v1405852 | !hlock3_p & v140585c;
assign d2fb8c = hbusreq0 & d2fb8b | !hbusreq0 & v845542;
assign d30806 = hmaster1_p & d30805 | !hmaster1_p & d307f4;
assign v134d43c = hbusreq1 & v134d370 | !hbusreq1 & v134d273;
assign v155338a = hready & v1553389 | !hready & v1553217;
assign v12160ba = hmaster1_p & v12160a1 | !hmaster1_p & v1216082;
assign v1553505 = hbusreq2 & v1553503 | !hbusreq2 & v1553504;
assign v14457a9 = hlock2 & v14457a5 | !hlock2 & v14457a8;
assign d307aa = hgrant5_p & v84554e | !hgrant5_p & d307a8;
assign v1445dc1 = hlock2 & v1445db4 | !hlock2 & v1445dbb;
assign v1552d7c = locked_p & v1552d7b | !locked_p & v845542;
assign v14457ae = hmaster1_p & v1445779 | !hmaster1_p & v1445e28;
assign v1215d84 = hbusreq2_p & v1215d7b | !hbusreq2_p & v1215d83;
assign d30842 = hbusreq2_p & d30840 | !hbusreq2_p & d30841;
assign v1445f42 = hbusreq2 & v1445f38 | !hbusreq2 & v1445f41;
assign v121623e = hgrant2_p & v1216202 | !hgrant2_p & v121623d;
assign v1515829 = hbusreq2 & v1515828 | !hbusreq2 & v15167ed;
assign v138a43f = hmaster1_p & v138a43b | !hmaster1_p & v138a43e;
assign d3080e = hmaster0_p & v84554e | !hmaster0_p & d3070e;
assign v12166f6 = hgrant5_p & v845542 | !hgrant5_p & v12166c5;
assign v12ad323 = hbusreq1_p & v12ae1fa | !hbusreq1_p & v12ad322;
assign v1668cae = hbusreq2_p & v1668caa | !hbusreq2_p & v1668cad;
assign d307a7 = hmaster2_p & d306cd | !hmaster2_p & v845542;
assign v16a2072 = hmastlock_p & v16a2667 | !hmastlock_p & !v845542;
assign v14461c0 = hlock2 & v144617b | !hlock2 & v14461bf;
assign v151564f = hmaster2_p & v151564d | !hmaster2_p & !v84556a;
assign f2f282 = hgrant1_p & f2f281 | !hgrant1_p & !v845542;
assign v121577e = hbusreq0 & v1215779 | !hbusreq0 & v121577d;
assign a65473 = hbusreq4_p & a65472 | !hbusreq4_p & !v845542;
assign v12ad5cd = hgrant5_p & v12ad5c7 | !hgrant5_p & !v12ad5cc;
assign v1216527 = locked_p & v1216526 | !locked_p & !v845542;
assign v12153b1 = hbusreq0 & v12153b0 | !hbusreq0 & v845542;
assign v14457bf = hlock2 & v14457bc | !hlock2 & v14457be;
assign v1445ee9 = hmaster2_p & v1445ec0 | !hmaster2_p & v1445def;
assign f2f450 = hbusreq5_p & f2f3c8 | !hbusreq5_p & !f2f44f;
assign v144671d = hlock3 & v1446700 | !hlock3 & v144671c;
assign v12ad517 = hbusreq0 & v12ad516 | !hbusreq0 & !v845542;
assign v1216054 = hbusreq1 & v1216ada | !hbusreq1 & v845542;
assign v134d3b8 = hlock3 & v134d3b5 | !hlock3 & v134d3b7;
assign v144623d = hmaster1_p & v144621d | !hmaster1_p & v1446236;
assign v144544e = hlock2 & v1445446 | !hlock2 & v144544d;
assign v144550e = hlock2 & v14454fa | !hlock2 & v144550d;
assign v134d236 = hlock2 & v134d227 | !hlock2 & v134d235;
assign v15168fc = hlock2_p & v15168fb | !hlock2_p & !v845542;
assign v1405841 = hmaster2_p & v140583d | !hmaster2_p & v14463b1;
assign v1515825 = hbusreq3 & v151581e | !hbusreq3 & v1515824;
assign d307de = hgrant5_p & d30705 | !hgrant5_p & d307dc;
assign v1445df3 = hmaster2_p & v1445df2 | !hmaster2_p & v1445def;
assign d300ef = hgrant5_p & d300d4 | !hgrant5_p & d300ee;
assign v134d3b0 = hgrant2_p & v134d3af | !hgrant2_p & v134d39b;
assign v144603d = hgrant1_p & v144639c | !hgrant1_p & v144603c;
assign v14058fd = hgrant1_p & v1446403 | !hgrant1_p & v14058fc;
assign v1668de6 = hbusreq3 & v1668de5 | !hbusreq3 & v845542;
assign v1515854 = hbusreq3_p & v151580b | !hbusreq3_p & v1515853;
assign v12150fb = hmaster1_p & v121543b | !hmaster1_p & v12150ef;
assign a6545d = hbusreq2_p & a6545a | !hbusreq2_p & a6545c;
assign v12afe67 = hmaster1_p & v12afe47 | !hmaster1_p & v12afe66;
assign v134d454 = hlock2 & v134d451 | !hlock2 & v134d453;
assign v1553100 = hbusreq2 & v15530ff | !hbusreq2 & v155321a;
assign v1516958 = hready_p & v1516900 | !hready_p & !v1516957;
assign v1216280 = hmaster0_p & v121600e | !hmaster0_p & v1215ff0;
assign v16a19b8 = hmaster1_p & v16a19b0 | !hmaster1_p & !v16a2672;
assign v1405872 = hmaster0_p & v1405861 | !hmaster0_p & v1405871;
assign d3084e = hbusreq1_p & d306fe | !hbusreq1_p & !v845542;
assign v16a2061 = hbusreq2 & v16a205f | !hbusreq2 & v16a2060;
assign v1445f27 = hmaster0_p & v1445da9 | !hmaster0_p & v144639c;
assign v1214eee = hgrant5_p & v845542 | !hgrant5_p & v1216531;
assign v1284ce9 = locked_p & v1284c8e | !locked_p & !v1405844;
assign v134d432 = hmaster0_p & v134d379 | !hmaster0_p & v134d431;
assign f2f404 = hmaster1_p & f2f3ef | !hmaster1_p & !f2f330;
assign d2fb11 = hmaster1_p & d2faf1 | !hmaster1_p & d2fb10;
assign v144539b = hlock2 & v1445396 | !hlock2 & v144539a;
assign v144609c = hmaster0_p & v1446404 | !hmaster0_p & v1446077;
assign v1214815 = hbusreq2 & v12147ff | !hbusreq2 & v121671a;
assign v121573f = hgrant5_p & v1215731 | !hgrant5_p & v121573e;
assign a658d4 = hmastlock_p & a658d3 | !hmastlock_p & v845580;
assign v134cdc9 = hbusreq5 & v134cdc7 | !hbusreq5 & v134cdc8;
assign bf1f64 = hlock5_p & bf1f61 | !hlock5_p & bf1f63;
assign v138a363 = hmaster1_p & v138a362 | !hmaster1_p & v138a341;
assign v1553425 = hready_p & v1553306 | !hready_p & v1553424;
assign v134d4a3 = hgrant2_p & v134d4a2 | !hgrant2_p & v134d49b;
assign v1389ff5 = hbusreq3 & v1389fe9 | !hbusreq3 & v1389ff2;
assign v12ad61f = hmaster1_p & v12ad61e | !hmaster1_p & !v12ad617;
assign v16a13dc = hmaster2_p & v16a207e | !hmaster2_p & v16a208a;
assign d2feb4 = hbusreq4_p & d2feb3 | !hbusreq4_p & v845542;
assign v14466e8 = hlock2 & v14466e5 | !hlock2 & v14466e7;
assign v1214ecb = hgrant5_p & v1216a5a | !hgrant5_p & v1216539;
assign v1515c86 = hbusreq2 & v15160fc | !hbusreq2 & v1515c85;
assign v134ce73 = hmaster1_p & v134ce72 | !hmaster1_p & v845542;
assign a65b21 = hready_p & a65b1a | !hready_p & a65b20;
assign v1445f1d = hbusreq5 & v1445f03 | !hbusreq5 & v1445f1c;
assign v144604f = hgrant1_p & v1445fcf | !hgrant1_p & v144604e;
assign v12ad0b8 = hmaster2_p & v845542 | !hmaster2_p & v12ad0b7;
assign v1445bdf = hgrant3_p & v1445bbd | !hgrant3_p & v1445bde;
assign v1669599 = hmaster0_p & v845570 | !hmaster0_p & v1668da6;
assign v14838ba = hgrant1_p & v845558 | !hgrant1_p & v14838b7;
assign v1405afb = hbusreq2_p & v1405af2 | !hbusreq2_p & v1405afa;
assign v1214bc1 = hlock2_p & v1214bbe | !hlock2_p & v1214bc0;
assign v12157ad = hgrant0_p & v845542 | !hgrant0_p & !v845559;
assign v14459ea = hmaster2_p & v144660b | !hmaster2_p & v14458eb;
assign d2fb7e = hbusreq0 & d2fb7d | !hbusreq0 & v845542;
assign v134d39c = hgrant2_p & v134d364 | !hgrant2_p & v134d39b;
assign v114a230 = hgrant4_p & v845542 | !hgrant4_p & !v845572;
assign v15530b4 = hready_p & v1553444 | !hready_p & v15530b3;
assign v15161cf = hbusreq2_p & v15161ce | !hbusreq2_p & !v845542;
assign v1445e87 = hbusreq0_p & v1446403 | !hbusreq0_p & v1445e5d;
assign v1215cc4 = hgrant5_p & v1215c82 | !hgrant5_p & v1215cc3;
assign d30844 = hbusreq5 & d30814 | !hbusreq5 & d30843;
assign v121507d = hgrant2_p & v1215024 | !hgrant2_p & v121507c;
assign v1552d48 = hlock0 & v1552d47 | !hlock0 & v1553392;
assign v16a1374 = hmaster1_p & v16a1329 | !hmaster1_p & v16a1f96;
assign v134d4f4 = hmaster2_p & v134d36d | !hmaster2_p & v845542;
assign v10d42d0 = hmaster0_p & v10d42a5 | !hmaster0_p & v10d428d;
assign v1445e45 = hbusreq4_p & v1446483 | !hbusreq4_p & v144649b;
assign d2fc65 = hbusreq0 & d2fc64 | !hbusreq0 & d302e7;
assign d30140 = hgrant5_p & d3013a | !hgrant5_p & !d300ee;
assign v138936e = hbusreq5_p & v138936d | !hbusreq5_p & v845542;
assign a658ba = stateA1_p & v156645f | !stateA1_p & !v110b6cc;
assign v1214fc2 = hmaster2_p & v12157b1 | !hmaster2_p & v1215750;
assign v1215789 = hgrant2_p & v1215786 | !hgrant2_p & v1215780;
assign v1445e80 = hgrant1_p & v1445dec | !hgrant1_p & v1445e68;
assign bf1f96 = hmaster2_p & bf1f91 | !hmaster2_p & bf1f95;
assign v134d1dd = locked_p & v134d1dc | !locked_p & v845542;
assign v1445791 = hmaster0_p & v144578b | !hmaster0_p & v1445e13;
assign v1214dea = hmaster0_p & v12162e9 | !hmaster0_p & v12162e8;
assign v12af5aa = hgrant1_p & v845542 | !hgrant1_p & v12af5a9;
assign v121632f = hbusreq2_p & v121632c | !hbusreq2_p & v1216326;
assign v1552fce = hbusreq2 & v1552fcc | !hbusreq2 & v1552fcd;
assign d3087b = decide_p & d3087a | !decide_p & v845570;
assign v16a1af0 = decide_p & v16a1aef | !decide_p & v16a20a5;
assign v1215409 = hbusreq2_p & v1215408 | !hbusreq2_p & v12153fc;
assign v1668cfc = hbusreq5_p & v1668cfb | !hbusreq5_p & v1668cc8;
assign v1668dc2 = hmaster2_p & a6588d | !hmaster2_p & v845570;
assign v134cd8e = hready_p & v134d34f | !hready_p & v134cd8d;
assign v1214c52 = hmaster2_p & v1214c4c | !hmaster2_p & v1214c51;
assign v15156d6 = hgrant1_p & v15156d5 | !hgrant1_p & a658bd;
assign v1445b70 = hbusreq2_p & v1445b64 | !hbusreq2_p & v1445b6f;
assign v1215cec = hmaster0_p & v1215ce6 | !hmaster0_p & v1215ceb;
assign v12ad4ff = hmaster0_p & v12ad4fb | !hmaster0_p & v12ad4fe;
assign v10d42a6 = hmaster0_p & v10d428d | !hmaster0_p & v10d42a5;
assign v1215077 = hmaster2_p & v1215060 | !hmaster2_p & !v1215467;
assign v12164c5 = hbusreq2_p & v12164c4 | !hbusreq2_p & v12164c3;
assign v1215c0c = hbusreq1_p & v121652d | !hbusreq1_p & v1216123;
assign d3021b = hmaster2_p & v845580 | !hmaster2_p & !d307ac;
assign d306d2 = hmaster0_p & d306ce | !hmaster0_p & d306d1;
assign v12afdb3 = hbusreq0 & v12afda5 | !hbusreq0 & v12afdb2;
assign v1446043 = hbusreq1_p & v1446634 | !hbusreq1_p & v14465bb;
assign v1214c28 = hbusreq0_p & v12164cf | !hbusreq0_p & v845547;
assign v1668ce7 = hmaster1_p & v1668cd9 | !hmaster1_p & v1668ce6;
assign v1446684 = hlock2 & v1446676 | !hlock2 & v1446683;
assign v1215ddd = hbusreq3_p & v1215db0 | !hbusreq3_p & v1215ddc;
assign v144581a = hlock3 & v1445800 | !hlock3 & v1445819;
assign v1215078 = hmaster2_p & v1214ffe | !hmaster2_p & v121503a;
assign v1668cbf = hmaster0_p & a658ad | !hmaster0_p & v1668cbe;
assign d308dc = hmaster2_p & v845542 | !hmaster2_p & d308db;
assign v14453ac = hbusreq2_p & v14453a6 | !hbusreq2_p & v14453ab;
assign v1214ef2 = hgrant5_p & v845542 | !hgrant5_p & !v1216547;
assign v16a1d9a = hmaster1_p & v16a1d92 | !hmaster1_p & v16a1f96;
assign v138a3ce = hmaster2_p & v845542 | !hmaster2_p & v15157a9;
assign v1215082 = hgrant2_p & v1215063 | !hgrant2_p & v1215081;
assign v1214d64 = hbusreq2 & v1214d61 | !hbusreq2 & v1214d63;
assign v14465d0 = hbusreq1 & v14465cc | !hbusreq1 & v14465cf;
assign v15534dc = hmaster1_p & v1553385 | !hmaster1_p & v15534db;
assign v1553388 = hmastlock_p & v1553387 | !hmastlock_p & v845542;
assign d308c5 = hbusreq5_p & d3082d | !hbusreq5_p & d308c4;
assign v12acfd5 = hbusreq2 & v12acfcd | !hbusreq2 & v12acfd4;
assign v1552d76 = decide_p & v155342e | !decide_p & v155341e;
assign d306ea = stateG3_0_p & v845542 | !stateG3_0_p & !v84556c;
assign v16a1be7 = hbusreq0 & v16a1be5 | !hbusreq0 & v16a1be6;
assign v10d4046 = hbusreq0_p & v10d3fef | !hbusreq0_p & !v10d402b;
assign v14459f2 = hlock1 & v14459ac | !hlock1 & v14459b6;
assign v1216062 = hlock2_p & v121605e | !hlock2_p & v1216061;
assign v1445e4b = hmaster1_p & v1446466 | !hmaster1_p & v1445e4a;
assign v15168f8 = hbusreq1_p & v15168f7 | !hbusreq1_p & v845542;
assign d3079c = hgrant4_p & d30783 | !hgrant4_p & v845542;
assign v1389e32 = hmaster1_p & v1389e27 | !hmaster1_p & v1389e31;
assign v1215383 = hbusreq5_p & v1215381 | !hbusreq5_p & v1215382;
assign v134ce53 = hmaster2_p & v845542 | !hmaster2_p & v134ce52;
assign v1445af4 = hbusreq2 & v1445aed | !hbusreq2 & v1445af3;
assign v1405851 = hmaster1_p & v1405850 | !hmaster1_p & v140584d;
assign v1389809 = hlock5_p & v1389808 | !hlock5_p & !v845542;
assign v1446194 = hmaster1_p & v1446193 | !hmaster1_p & v1445fde;
assign v138a3c3 = hmaster0_p & v138a2fa | !hmaster0_p & v138a2f8;
assign v12ad4cd = hmaster2_p & v12ad4ca | !hmaster2_p & v12ad4cc;
assign d2fba4 = hbusreq2_p & d2fba3 | !hbusreq2_p & d2fb9f;
assign v11e597f = hbusreq2_p & v11e595e | !hbusreq2_p & v11e597e;
assign v144643d = hmaster2_p & v144639c | !hmaster2_p & v1446407;
assign v1553148 = hbusreq4_p & v1553147 | !hbusreq4_p & v845542;
assign v1215b84 = hbusreq5_p & v1215b82 | !hbusreq5_p & v1215b83;
assign v138a44f = hmaster1_p & v138a44e | !hmaster1_p & v138a341;
assign v121506d = hgrant2_p & v1215024 | !hgrant2_p & v121506c;
assign v12147fe = hgrant2_p & v845542 | !hgrant2_p & v12147fd;
assign d3067c = hmaster0_p & d3067a | !hmaster0_p & d3067b;
assign v12ad59d = hlock0_p & v1515714 | !hlock0_p & !v845542;
assign a66290 = hgrant5_p & v845542 | !hgrant5_p & a6628f;
assign v121629b = hbusreq0 & v1216193 | !hbusreq0 & v121629a;
assign v16a1d9f = decide_p & v16a1d2b | !decide_p & !v16a1d9e;
assign v1446331 = hbusreq0 & v1446330 | !hbusreq0 & v14462e7;
assign v1284cd3 = hgrant5_p & v14058a2 | !hgrant5_p & v1284cd2;
assign v134cf42 = hbusreq3_p & v134ced0 | !hbusreq3_p & v134cf41;
assign v1215cd3 = hbusreq5_p & v1215cd1 | !hbusreq5_p & !v1215cd2;
assign v14465c1 = hbusreq4 & v14465bf | !hbusreq4 & v14465c0;
assign d305df = hmaster2_p & v845570 | !hmaster2_p & !d305de;
assign a65ae4 = hgrant1_p & v845542 | !hgrant1_p & !a65ae2;
assign d30873 = hbusreq2 & d30871 | !hbusreq2 & d30872;
assign v1214bca = hmaster2_p & v1215399 | !hmaster2_p & v121539d;
assign v138a347 = hbusreq2_p & v138a342 | !hbusreq2_p & v138a346;
assign v16695ab = hbusreq2_p & v1669596 | !hbusreq2_p & v845570;
assign v1215068 = hgrant2_p & v1215063 | !hgrant2_p & v1215067;
assign v1215d36 = hmaster2_p & v845570 | !hmaster2_p & v1216596;
assign v12acff4 = hmaster1_p & v12acff3 | !hmaster1_p & v12ad5e1;
assign a658de = hbusreq0_p & a658dc | !hbusreq0_p & a658ca;
assign v1214d1e = hmaster0_p & v1214d1d | !hmaster0_p & !v1214d03;
assign v16a1f93 = hbusreq2 & v16a267a | !hbusreq2 & v16a267b;
assign v144642d = hbusreq5_p & v144642c | !hbusreq5_p & v144642a;
assign v138a3dc = hgrant5_p & v845570 | !hgrant5_p & !v1515781;
assign v1214bcf = hmaster0_p & v1214bce | !hmaster0_p & v12153a8;
assign v16a1a8b = hbusreq2 & v16a1a88 | !hbusreq2 & !v16a1a8a;
assign d3014b = hlock5_p & d30149 | !hlock5_p & d3014a;
assign v1445825 = hmaster1_p & v14457e4 | !hmaster1_p & v1445ef0;
assign v10d3ffb = hmaster0_p & v10d3ff6 | !hmaster0_p & v10d3ffa;
assign a65376 = hgrant4_p & v845570 | !hgrant4_p & !a65852;
assign v16a1cdc = hmaster1_p & v16a1ccc | !hmaster1_p & !v16a1f96;
assign v1446338 = hbusreq2 & v1446327 | !hbusreq2 & v1446337;
assign v121657c = hmaster0_p & v845542 | !hmaster0_p & v1216a7f;
assign f2f3de = hgrant2_p & f2f3b4 | !hgrant2_p & !f2f3da;
assign v138a3c8 = hgrant5_p & v845570 | !hgrant5_p & !v151572e;
assign f2f2b1 = decide_p & f2f2b0 | !decide_p & v845542;
assign v1216572 = hlock5_p & v121656e | !hlock5_p & v1216571;
assign v138a336 = hbusreq1 & v1668cbd | !hbusreq1 & !v138a335;
assign v1445b64 = hgrant2_p & v144634f | !hgrant2_p & v1445b60;
assign v121613b = hbusreq4 & v1215fec | !hbusreq4 & v1216014;
assign v121651f = hmaster1_p & v121651e | !hmaster1_p & v845547;
assign v12160a5 = hbusreq2_p & v12160a4 | !hbusreq2_p & v12160a3;
assign v1553140 = hmastlock_p & v155313f | !hmastlock_p & v845542;
assign d306a5 = hgrant4_p & v845558 | !hgrant4_p & d306a4;
assign v16a1dba = decide_p & v16a1db8 | !decide_p & v16a1db9;
assign v134ce3c = hbusreq0_p & v134d37d | !hbusreq0_p & v134d273;
assign v1445893 = hbusreq1 & v1445890 | !hbusreq1 & v1445892;
assign v1552d6a = hlock5 & v155341e | !hlock5 & v1552d5a;
assign v16a1cf9 = hmaster1_p & v16a1cf8 | !hmaster1_p & v16a1be8;
assign v144606b = hmaster2_p & v144605a | !hmaster2_p & v144606a;
assign d307f7 = hmaster2_p & d306fc | !hmaster2_p & !d307ad;
assign d307bc = hbusreq1 & d307bb | !hbusreq1 & v845542;
assign v1445bd3 = hgrant5_p & v14465d5 | !hgrant5_p & v1445bd2;
assign v16a144b = jx0_p & v16a16b7 | !jx0_p & v16a144a;
assign v1214eb4 = hbusreq5 & v1214e67 | !hbusreq5 & v1214eb3;
assign d30833 = hgrant5_p & d306d0 | !hgrant5_p & d307fa;
assign v1445ada = hmaster1_p & v14458aa | !hmaster1_p & v14458c1;
assign d30694 = hbusreq0 & d30692 | !hbusreq0 & d30693;
assign v1445dd0 = hlock0 & v1445dcf | !hlock0 & v1445dce;
assign v144578f = hmaster1_p & v144578e | !hmaster1_p & v1445e07;
assign v16a2076 = hgrant1_p & v84554d | !hgrant1_p & v16a2075;
assign d300ca = hlock4_p & v845542 | !hlock4_p & d300ba;
assign v1215bf4 = hgrant5_p & v121601c | !hgrant5_p & !v1215bf2;
assign a6544c = hgrant2_p & a6540a | !hgrant2_p & a6543a;
assign v15167c1 = hmaster1_p & v15167c0 | !hmaster1_p & v845542;
assign v1214c41 = hready_p & v121538e | !hready_p & v1214c40;
assign v1553415 = hbusreq0 & v1553414 | !hbusreq0 & v1553218;
assign v1445bd8 = hmaster0_p & v144643b | !hmaster0_p & v1446636;
assign f2f33d = hbusreq2_p & f2f33b | !hbusreq2_p & f2f33c;
assign v1445fb9 = hgrant5_p & v1445fb7 | !hgrant5_p & !v1445fb8;
assign f2f3b4 = hmaster1_p & f2f3b3 | !hmaster1_p & ae2496;
assign v121678f = hgrant3_p & v121651a | !hgrant3_p & v121678e;
assign d30705 = hmaster2_p & d30701 | !hmaster2_p & d30704;
assign v138a340 = hbusreq0 & v138a33b | !hbusreq0 & v138a33f;
assign v12ad560 = hbusreq2_p & v12ad55e | !hbusreq2_p & v12ad55f;
assign v13895a0 = hlock5_p & v138959f | !hlock5_p & v845542;
assign d30281 = hbusreq5_p & d30280 | !hbusreq5_p & !d3027f;
assign v1215728 = hbusreq4_p & v1215727 | !hbusreq4_p & v845542;
assign d30617 = hbusreq2_p & d30616 | !hbusreq2_p & d3060e;
assign v16a1ae4 = hbusreq2_p & v16a2098 | !hbusreq2_p & v16a1ae3;
assign d307d4 = hbusreq0_p & v845542 | !hbusreq0_p & d307ac;
assign v16a19bf = hbusreq2 & v16a19b7 | !hbusreq2 & v16a19b9;
assign v1515668 = hgrant1_p & v1515667 | !hgrant1_p & a658e0;
assign v1405900 = hmaster0_p & v14058f8 | !hmaster0_p & !v14058ff;
assign v12ad0cc = hready_p & v845542 | !hready_p & v12ad0cb;
assign v1668dd9 = hbusreq5_p & v1668dd7 | !hbusreq5_p & !v1668dd8;
assign v1668d53 = hbusreq1_p & v1668d51 | !hbusreq1_p & !v1668d52;
assign v1215795 = hbusreq5_p & v1215793 | !hbusreq5_p & v1215794;
assign v1445b91 = hgrant2_p & v1445b65 | !hgrant2_p & v1445b90;
assign f2f429 = hgrant5_p & f2f363 | !hgrant5_p & f2f428;
assign v12153c4 = decide_p & v1215bab | !decide_p & v12153c3;
assign v1215bd7 = hbusreq3 & v845542 | !hbusreq3 & v12164e7;
assign v14466d6 = hlock3 & v14466d3 | !hlock3 & v14466d5;
assign d30788 = stateG2_p & v845542 | !stateG2_p & a66292;
assign v10d407f = hmaster2_p & v10d3fd5 | !hmaster2_p & v10d3fdf;
assign v12afe71 = hmaster1_p & v12afe47 | !hmaster1_p & v12afe70;
assign v14461db = hbusreq2 & v14461d6 | !hbusreq2 & v14461da;
assign v12166ec = hgrant5_p & v845542 | !hgrant5_p & v12166eb;
assign v16a197e = hbusreq0 & v16a209a | !hbusreq0 & v16a197d;
assign v1215364 = hlock0_p & v845547 | !hlock0_p & !v845542;
assign v138959f = hmaster2_p & v15160ff | !hmaster2_p & v845542;
assign v14058b7 = hmaster2_p & v1405891 | !hmaster2_p & v1405844;
assign v1216a69 = hlock5_p & v1216a62 | !hlock5_p & v1216a68;
assign v14457d2 = hlock5 & v1445786 | !hlock5 & v14457d0;
assign v1445a20 = hbusreq0 & v1445a1c | !hbusreq0 & v1445a1f;
assign v1445f5e = hlock2 & v144673f | !hlock2 & v1445f5d;
assign v11e5952 = hlock4_p & v11e593a | !hlock4_p & v845570;
assign v12ad50b = hbusreq3 & v12ad505 | !hbusreq3 & !v12ad50a;
assign v1215384 = hbusreq0 & v1215383 | !hbusreq0 & v845542;
assign v1216184 = hmaster2_p & v845542 | !hmaster2_p & v121601d;
assign v1215cbe = hgrant5_p & v1215c82 | !hgrant5_p & v1215cbd;
assign v1445f0b = hgrant2_p & v1445ee8 | !hgrant2_p & v1445f0a;
assign v1216009 = hlock1_p & v1216005 | !hlock1_p & v1216008;
assign v1553089 = hbusreq1 & v155304d | !hbusreq1 & v155304e;
assign d80777 = hlock5_p & d80775 | !hlock5_p & !d80776;
assign v10d42ca = hmaster2_p & v10d42c9 | !hmaster2_p & v10d403a;
assign v155351c = jx2_p & v1553448 | !jx2_p & v155351b;
assign f2e4f4 = decide_p & f2e4f3 | !decide_p & f2f23c;
assign d3081a = hgrant5_p & v84554e | !hgrant5_p & d307a1;
assign v1446090 = hgrant5_p & v1445fe8 | !hgrant5_p & v144608f;
assign v1445912 = hbusreq2_p & v144590f | !hbusreq2_p & v1445911;
assign v14460fe = hbusreq2 & v14460fc | !hbusreq2 & v14460fd;
assign v1405b19 = hgrant4_p & v1405abf | !hgrant4_p & v1405b18;
assign v16a1cf1 = hgrant2_p & v845542 | !hgrant2_p & v16a1cf0;
assign v1446702 = hbusreq2 & v14466f8 | !hbusreq2 & v1446701;
assign v1284d47 = hgrant2_p & v1284d44 | !hgrant2_p & v1284d46;
assign v1668c46 = hbusreq3 & v1668c3e | !hbusreq3 & v1668c45;
assign v1552f5f = hgrant0_p & v1552f5e | !hgrant0_p & v845542;
assign f2f3be = hbusreq0 & f2f3ba | !hbusreq0 & f2f3bd;
assign v15530a9 = hmaster0_p & v155308b | !hmaster0_p & v845542;
assign v1214de3 = decide_p & v1214dde | !decide_p & v1214de2;
assign f2f457 = hbusreq2_p & f2f444 | !hbusreq2_p & f2f456;
assign a65366 = stateA1_p & v845542 | !stateA1_p & !a65365;
assign f2f353 = hbusreq1 & v1668d2e | !hbusreq1 & v845542;
assign v1215d08 = hgrant2_p & v1215cdc | !hgrant2_p & v1215cfb;
assign v134d277 = decide_p & v134d272 | !decide_p & v134d276;
assign d301d8 = hmaster2_p & d301d7 | !hmaster2_p & v845542;
assign v1446423 = hlock0_p & v1446403 | !hlock0_p & v1446422;
assign v14460c4 = hbusreq2_p & v14460b8 | !hbusreq2_p & v14460c3;
assign v134cd7b = hmaster2_p & v134cd6e | !hmaster2_p & v845542;
assign v134d27e = hgrant1_p & v845542 | !hgrant1_p & v134d27d;
assign v1445a0a = hbusreq4 & v1445a09 | !hbusreq4 & v14459b3;
assign d30780 = hbusreq4 & d306c8 | !hbusreq4 & v845542;
assign v1216ae4 = hmaster2_p & v1216adf | !hmaster2_p & v1216ae3;
assign d30103 = hbusreq5_p & d30102 | !hbusreq5_p & d30101;
assign v1216022 = hlock1_p & v1216021 | !hlock1_p & !v845542;
assign d2fbd7 = hgrant5_p & d2fb4d | !hgrant5_p & d2fbd6;
assign v1446078 = hbusreq0 & v1446076 | !hbusreq0 & v1446077;
assign v16a1d6e = hmaster0_p & v16a1d6c | !hmaster0_p & v16a1d6d;
assign a653ad = hbusreq1 & a653a9 | !hbusreq1 & v845558;
assign v14453fb = hlock2 & v14453f5 | !hlock2 & v14453fa;
assign v1445ac9 = hlock2 & v1445ac6 | !hlock2 & v1445ac8;
assign v1214f03 = hbusreq0 & v1214f01 | !hbusreq0 & v1214f02;
assign f2f2d7 = hbusreq1 & a658e0 | !hbusreq1 & !v845542;
assign v1445af5 = hmaster0_p & v1445a4f | !hmaster0_p & v14458d4;
assign v14058bf = hbusreq2_p & v14058b3 | !hbusreq2_p & v14058be;
assign v1214bd2 = hlock2_p & v1214bd0 | !hlock2_p & v1214bd1;
assign v16a195e = hgrant2_p & v845542 | !hgrant2_p & !v16a195c;
assign v10d426b = hgrant1_p & v10d4019 | !hgrant1_p & v10d426a;
assign d2fee0 = hbusreq2 & d2fedb | !hbusreq2 & d2fedf;
assign v16a1985 = decide_p & v16a196d | !decide_p & v16a1984;
assign v1215cdb = hmaster1_p & v1215cda | !hmaster1_p & v845542;
assign d8076e = hmaster2_p & d8076d | !hmaster2_p & v845542;
assign d3025a = hgrant2_p & d3021d | !hgrant2_p & !d30259;
assign v16a1d73 = hgrant2_p & v845542 | !hgrant2_p & !v16a1d6f;
assign v134d430 = hbusreq0 & v134d42f | !hbusreq0 & v134d429;
assign f2f338 = hmaster1_p & f2f2ed | !hmaster1_p & !f2f330;
assign v12ad5be = hlock0_p & v1515744 | !hlock0_p & d2fbe5;
assign v1668d25 = hbusreq4 & v10d3fd8 | !hbusreq4 & !v845542;
assign d30792 = hbusreq1_p & d30791 | !hbusreq1_p & v845542;
assign v15156e3 = hmaster2_p & v15156c7 | !hmaster2_p & !v1668cc6;
assign v1214f64 = decide_p & v1214ec1 | !decide_p & v1214f63;
assign v14457ed = hmaster0_p & v1445eb6 | !hmaster0_p & v144639c;
assign v1445449 = hbusreq2_p & v1445448 | !hbusreq2_p & v1445bb3;
assign v14058e8 = hgrant0_p & v140587c | !hgrant0_p & v14058e7;
assign v12153f3 = hmaster2_p & v12153ce | !hmaster2_p & v12153d9;
assign v1214fc6 = hmaster1_p & v1214fc5 | !hmaster1_p & v1214fbf;
assign v12ad547 = hbusreq2 & v12ad53f | !hbusreq2 & v12ad546;
assign a6567a = hmaster1_p & a6566b | !hmaster1_p & a65678;
assign v1446047 = hbusreq1_p & v144663e | !hbusreq1_p & v14465d7;
assign v14457a4 = hmaster1_p & v14457a3 | !hmaster1_p & v1445e07;
assign d30126 = hmaster0_p & d2fe80 | !hmaster0_p & d30125;
assign v14458b2 = hmaster1_p & v14458b1 | !hmaster1_p & v14458af;
assign d3071c = hlock1_p & v845542 | !hlock1_p & d305ea;
assign v16a1abe = hmaster1_p & v16a1abd | !hmaster1_p & !v16a2672;
assign v1215d65 = hmaster2_p & v845570 | !hmaster2_p & v12164d9;
assign d306f5 = hlock1_p & d306f4 | !hlock1_p & d305de;
assign v134d4ae = hmaster0_p & v134d4ad | !hmaster0_p & v134d499;
assign v1445a0f = hbusreq4 & v1445a0e | !hbusreq4 & v14459c3;
assign v14463f2 = hbusreq1 & v14463d8 | !hbusreq1 & v14463f1;
assign v134cd67 = hmaster2_p & v134d389 | !hmaster2_p & v134cd66;
assign v1668d19 = hmaster2_p & a65851 | !hmaster2_p & v1668d18;
assign v138945e = hmaster0_p & v1389de1 | !hmaster0_p & v1389ffd;
assign v16a1407 = hbusreq2 & v16a1406 | !hbusreq2 & !v16a209e;
assign v1215c43 = hgrant5_p & v1216029 | !hgrant5_p & !v1215c41;
assign v1446625 = hlock0_p & v144639c | !hlock0_p & v1446624;
assign v1215b93 = hmaster2_p & v845542 | !hmaster2_p & v1215b92;
assign d301e3 = hbusreq5_p & d301e2 | !hbusreq5_p & !d301e1;
assign v1215035 = hbusreq1 & v121502d | !hbusreq1 & v1214ff5;
assign v12afe60 = hgrant0_p & v84554a | !hgrant0_p & !v845542;
assign v144613d = hlock2 & v1446125 | !hlock2 & v144613b;
assign v134d1ec = hbusreq4 & v134d1ea | !hbusreq4 & v134d1eb;
assign d30248 = hgrant5_p & d30242 | !hgrant5_p & !d301fa;
assign d2f98c = hbusreq1_p & d2f98b | !hbusreq1_p & v84555a;
assign v1405b45 = hmaster0_p & v1405a96 | !hmaster0_p & v1405af3;
assign v12af9d3 = hgrant1_p & d30690 | !hgrant1_p & v12af9d2;
assign v1214cfa = hmaster2_p & v1214cf9 | !hmaster2_p & v1214cf5;
assign a653e7 = hmaster0_p & a653c0 | !hmaster0_p & a653e6;
assign v14466dd = hmaster1_p & v14466dc | !hmaster1_p & v14463ef;
assign v1215cb4 = hgrant1_p & f2f285 | !hgrant1_p & v1215cad;
assign v14058c8 = hmaster2_p & v14463b1 | !hmaster2_p & v14058c7;
assign f2e711 = hlock1_p & f2e710 | !hlock1_p & !v845542;
assign v14459d5 = hbusreq0_p & v845542 | !hbusreq0_p & v1446403;
assign d3089f = hgrant1_p & v84554c | !hgrant1_p & d3089e;
assign f2e73c = decide_p & f2e734 | !decide_p & f2f23c;
assign d2fd1e = hbusreq5_p & d2fd1d | !hbusreq5_p & !d2fd1c;
assign v1445edd = hmaster2_p & v144639c | !hmaster2_p & v1445edc;
assign v1215720 = hgrant4_p & v845542 | !hgrant4_p & v121571f;
assign v134d4d9 = hgrant1_p & v845542 | !hgrant1_p & v134d4d8;
assign v121603d = hbusreq1_p & v121603c | !hbusreq1_p & v845542;
assign v12ad4c3 = hmaster0_p & v12af73f | !hmaster0_p & v12ad4c2;
assign d2fd4f = jx0_p & d302f9 | !jx0_p & d2fd4e;
assign v14463dd = hbusreq5_p & v14463dc | !hbusreq5_p & v14463a6;
assign v1445e35 = hbusreq5 & v1445e33 | !hbusreq5 & v1445e34;
assign a653df = hgrant4_p & v845570 | !hgrant4_p & !a653de;
assign v1445d95 = hlock0 & v1445d94 | !hlock0 & v1445d8d;
assign v84555c = hbusreq5_p & v845542 | !hbusreq5_p & !v845542;
assign v1214db5 = hbusreq2 & v1214db0 | !hbusreq2 & v1214db4;
assign v14459b7 = hlock1 & v144660b | !hlock1 & v14459b6;
assign v15168f4 = locked_p & v15168f3 | !locked_p & !v845542;
assign v1445b8a = hbusreq5_p & v14462ea | !hbusreq5_p & v1445b89;
assign v1445aee = hmaster0_p & v1445a36 | !hmaster0_p & v14458d4;
assign v12ad4fb = hbusreq0 & v12ad4fa | !hbusreq0 & v845542;
assign d2fc12 = hmaster1_p & d2fbdb | !hmaster1_p & d2fc11;
assign v166959c = hlock3_p & v166959b | !hlock3_p & !v845542;
assign f2e4fe = hbusreq2_p & f2e4fd | !hbusreq2_p & f2ed99;
assign v138a484 = hmaster1_p & v138a483 | !hmaster1_p & v84555c;
assign v155342f = hmaster0_p & v1553416 | !hmaster0_p & v845542;
assign v12160b6 = hlock2_p & v12160b4 | !hlock2_p & v12160b5;
assign d306fd = hmaster2_p & d306fc | !hmaster2_p & !v84554e;
assign v14453c5 = hready_p & v1445bca | !hready_p & v14453c4;
assign v1552d94 = hgrant2_p & v1552d93 | !hgrant2_p & v1552d8f;
assign v1445b28 = hbusreq3 & v1445b1e | !hbusreq3 & v1445b27;
assign v134d510 = hgrant5_p & v845542 | !hgrant5_p & v134d50f;
assign v16a1bfe = hbusreq0 & v16a209a | !hbusreq0 & v16a1bfd;
assign v1445b4d = hgrant2_p & v1445b46 | !hgrant2_p & v1445b48;
assign v16a16ac = hbusreq2_p & v16a1e0b | !hbusreq2_p & v16a16ab;
assign v138a339 = hlock5_p & v138a333 | !hlock5_p & !v138a338;
assign v1445f56 = hmaster1_p & v1446663 | !hmaster1_p & v1446630;
assign v1445f82 = hready_p & v14465a9 | !hready_p & v1445f81;
assign d2fc78 = hbusreq2_p & d2fc13 | !hbusreq2_p & d2fc77;
assign a6568f = hmaster1_p & a65495 | !hmaster1_p & a658e5;
assign a6627a = hmaster2_p & a66278 | !hmaster2_p & !v845542;
assign v16a1d63 = hmaster1_p & v16a1d5d | !hmaster1_p & v16a1d62;
assign a65381 = hgrant1_p & a65362 | !hgrant1_p & !a65380;
assign d2fd27 = hgrant2_p & v845542 | !hgrant2_p & d2fd26;
assign d80758 = stateG2_p & v845542 | !stateG2_p & !d80757;
assign v1445920 = hbusreq2_p & v144591c | !hbusreq2_p & v144591f;
assign v16a1430 = hbusreq5 & v16a142d | !hbusreq5 & v16a142f;
assign v14461fb = hbusreq2_p & v14461ee | !hbusreq2_p & v14461fa;
assign v138a353 = hmaster2_p & v138a32b | !hmaster2_p & a658ca;
assign v12ad009 = hbusreq1_p & v12ad5af | !hbusreq1_p & v12ad002;
assign v12161b0 = hgrant2_p & v12161a8 | !hgrant2_p & v12161af;
assign v16a141f = hbusreq2_p & v16a13c1 | !hbusreq2_p & v16a1da3;
assign v1668cce = hmastlock_p & v1668ccd | !hmastlock_p & !v845542;
assign d3018e = hmaster0_p & d3090c | !hmaster0_p & d3018d;
assign d8077d = hlock0_p & d80733 | !hlock0_p & !v845542;
assign v1214d65 = hmaster1_p & v1214d55 | !hmaster1_p & v1214d5f;
assign v134d4ec = hgrant5_p & v134d36a | !hgrant5_p & v134d4eb;
assign v14453f5 = hbusreq2_p & v1446272 | !hbusreq2_p & v14453f3;
assign d3090f = hbusreq1 & d305ea | !hbusreq1 & !v16693aa;
assign v1389d71 = hmaster2_p & v15168b0 | !hmaster2_p & v845542;
assign f2f39e = hmaster1_p & f2f397 | !hmaster1_p & f2f39d;
assign d2fad8 = hbusreq1_p & d300b7 | !hbusreq1_p & !d2fad7;
assign v144542d = hgrant2_p & v144542b | !hgrant2_p & v144542c;
assign d3021c = hmaster0_p & v845580 | !hmaster0_p & d3021b;
assign v15168fb = hmaster1_p & v15168fa | !hmaster1_p & v1668c44;
assign v121535e = hlock0_p & v1216a73 | !hlock0_p & v121535d;
assign v16a1af1 = decide_p & v16a1ad5 | !decide_p & v16a1ab9;
assign v1284ca5 = hlock0_p & v1284c8e | !hlock0_p & !v14463ba;
assign d301a2 = hmaster2_p & d3094f | !hmaster2_p & !d30952;
assign v134d215 = hmaster2_p & v134d1e8 | !hmaster2_p & v134d214;
assign v138a313 = hlock5_p & v10d3ffa | !hlock5_p & !v845542;
assign v16a1d1f = hmaster0_p & v16a1d1a | !hmaster0_p & v16a1d1e;
assign v16a205a = hbusreq2 & v16a2058 | !hbusreq2 & v16a2059;
assign d2fc7f = hready_p & d2fc7c | !hready_p & d2fc47;
assign d807b2 = hbusreq2_p & d807ad | !hbusreq2_p & d807b1;
assign v1668d6d = locked_p & v1668d6c | !locked_p & !v845542;
assign v144538b = hlock2 & v1445354 | !hlock2 & v144538a;
assign v1668db4 = hgrant5_p & v845542 | !hgrant5_p & !v1668d29;
assign v1214bb6 = hmaster1_p & v1214bb5 | !hmaster1_p & v12153a9;
assign v134ce7b = hready_p & v134d3be | !hready_p & v134ce7a;
assign v16695ac = hmaster0_p & v1668c1d | !hmaster0_p & v1668da6;
assign v1668db9 = hbusreq0 & v1668db5 | !hbusreq0 & v1668db8;
assign v138a45b = hbusreq2_p & v138a458 | !hbusreq2_p & v138a45a;
assign jx2 = v11f3405;
assign d301a1 = hlock2_p & d3019f | !hlock2_p & d301a0;
assign d30795 = hbusreq1_p & d30794 | !hbusreq1_p & v845542;
assign d2f9d1 = hmaster1_p & d2f99c | !hmaster1_p & d2f9d0;
assign a65674 = hgrant5_p & v949cd9 | !hgrant5_p & a6564d;
assign d2fbc4 = decide_p & d2fbc3 | !decide_p & v845570;
assign v151572b = hgrant0_p & a6537d | !hgrant0_p & a65851;
assign a653b6 = hgrant5_p & a653ab | !hgrant5_p & !a653b5;
assign v1214c60 = hlock5_p & v1214c5e | !hlock5_p & v1214c5f;
assign v1214c67 = hbusreq1 & v121536a | !hbusreq1 & v845542;
assign v1214cc7 = hbusreq0_p & v1214cc6 | !hbusreq0_p & !v845542;
assign a65440 = hgrant5_p & a6587e | !hgrant5_p & a653fd;
assign v14457d3 = hbusreq5 & v14457d1 | !hbusreq5 & v14457d2;
assign d2fbc1 = hbusreq2 & d2fbbd | !hbusreq2 & d2fbc0;
assign v16a206c = hgrant4_p & v845559 | !hgrant4_p & v16a206b;
assign v121611b = hlock5_p & v1216119 | !hlock5_p & v121611a;
assign a65361 = hbusreq1 & a65360 | !hbusreq1 & !v845558;
assign v1553433 = hlock3 & v155321a | !hlock3 & v1553432;
assign v1214c61 = hgrant1_p & v1214c46 | !hgrant1_p & v1214c50;
assign d30723 = hbusreq1_p & d30722 | !hbusreq1_p & v84555a;
assign v1515648 = stateA1_p & a658a7 | !stateA1_p & !v1515647;
assign v10d4093 = hmaster0_p & v10d408c | !hmaster0_p & v10d4092;
assign v134d443 = hgrant2_p & v134d442 | !hgrant2_p & v134d433;
assign v1214d5a = hbusreq2 & v1214d57 | !hbusreq2 & v1214d59;
assign v1214bc2 = hbusreq2_p & v1214bc1 | !hbusreq2_p & v1214bc0;
assign v134d3e5 = decide_p & v134d3e4 | !decide_p & v134d316;
assign v1445df4 = hbusreq5_p & v1445df0 | !hbusreq5_p & v1445df3;
assign d300c4 = hgrant1_p & d300c0 | !hgrant1_p & d300c3;
assign v1215d77 = hgrant5_p & v12164df | !hgrant5_p & v12166eb;
assign v1445f95 = hbusreq1_p & v1445f94 | !hbusreq1_p & v14463bb;
assign v1445e7e = hgrant5_p & v1445e79 | !hgrant5_p & v1445e7d;
assign f2ec22 = hbusreq1_p & f2ec21 | !hbusreq1_p & !v845542;
assign v1215742 = hlock5_p & v121573f | !hlock5_p & v1215741;
assign v14457f7 = hmaster0_p & v14457d7 | !hmaster0_p & v1445edf;
assign d30890 = hbusreq1_p & d307bd | !hbusreq1_p & d306a5;
assign v134d380 = hgrant4_p & v134d273 | !hgrant4_p & v845542;
assign v134d50d = hgrant1_p & v845542 | !hgrant1_p & v134d4fc;
assign a6563f = hbusreq5_p & a653ba | !hbusreq5_p & !a6563e;
assign d2fea8 = hlock4_p & d3070c | !hlock4_p & v845542;
assign v1446139 = hmaster0_p & v14460a5 | !hmaster0_p & v1445fea;
assign a658c6 = hmastlock_p & a658c3 | !hmastlock_p & v845542;
assign v16a1d34 = hbusreq3 & v16a1d33 | !hbusreq3 & v16a2063;
assign v1668e09 = decide_p & v1668e08 | !decide_p & !v845542;
assign v8a9c96 = stateG3_0_p & v845542 | !stateG3_0_p & acd334;
assign v1446097 = hlock2 & v1446085 | !hlock2 & v1446096;
assign v1215337 = hbusreq2 & v1215333 | !hbusreq2 & v1215336;
assign v144611f = hbusreq2_p & v1446119 | !hbusreq2_p & v144611e;
assign v1515645 = hlock3_p & v1515637 | !hlock3_p & v1515644;
assign v12af989 = hbusreq1_p & v84554a | !hbusreq1_p & v12af988;
assign a65452 = hbusreq2 & a6544b | !hbusreq2 & a65451;
assign d302db = hbusreq2_p & d302d6 | !hbusreq2_p & d302da;
assign v1405a9b = hmaster0_p & v1405a8a | !hmaster0_p & v1405a96;
assign v1445e96 = hbusreq0 & v1445e92 | !hbusreq0 & v1445e95;
assign v1215052 = hgrant5_p & v121546e | !hgrant5_p & v1215051;
assign v1446146 = hlock2 & v1446143 | !hlock2 & v1446145;
assign v1215b96 = hbusreq3 & v1215b8d | !hbusreq3 & v1215b95;
assign a654ae = hmaster2_p & a658cb | !hmaster2_p & !a6546d;
assign v1446479 = hgrant1_p & v1446478 | !hgrant1_p & v845542;
assign f2f409 = hbusreq2_p & f2f407 | !hbusreq2_p & f2f408;
assign v1405b12 = hgrant0_p & v1405abb | !hgrant0_p & v1405aa2;
assign d3027e = hgrant5_p & v845570 | !hgrant5_p & d30669;
assign v1445ace = hbusreq3 & v1445acc | !hbusreq3 & v1445acd;
assign v1214ce4 = hbusreq2_p & v1214cda | !hbusreq2_p & v1214ce3;
assign v134d273 = locked_p & v134d1e8 | !locked_p & v845542;
assign v121540f = hmaster0_p & v121540e | !hmaster0_p & v12153eb;
assign v12161fb = hgrant5_p & f2f2a8 | !hgrant5_p & v12161fa;
assign d2fc4f = hgrant1_p & d2fbcb | !hgrant1_p & d2fc4e;
assign v1668c54 = hready_p & v1668c48 | !hready_p & !v1668c53;
assign v134cd78 = hbusreq2 & v134cd76 | !hbusreq2 & v134cd77;
assign v121579f = hmaster0_p & v121579b | !hmaster0_p & v121579e;
assign v1668d5b = hmaster2_p & v1668d3c | !hmaster2_p & v1668d5a;
assign v10d40a7 = hmaster1_p & v10d3ffd | !hmaster1_p & v10d3ffb;
assign d2febe = hbusreq5_p & d2febd | !hbusreq5_p & d2febc;
assign v16a1e4c = hgrant2_p & v16a1d31 | !hgrant2_p & v16a1e4b;
assign v1515630 = locked_p & v151562f | !locked_p & !v845542;
assign v1668c99 = hmaster2_p & a658bd | !hmaster2_p & !v1668c64;
assign v1214dc8 = hready_p & v1214da6 | !hready_p & v1214dc7;
assign v14465f6 = hbusreq0_p & v144639c | !hbusreq0_p & v14465be;
assign d8073c = hlock1_p & d80732 | !hlock1_p & !v845542;
assign a6585c = locked_p & a6585b | !locked_p & v10d3fd8;
assign v121627a = hmaster1_p & v1216279 | !hmaster1_p & v12160e0;
assign v1445f89 = hmaster2_p & v14463b1 | !hmaster2_p & !v14463a5;
assign v1445783 = hmaster1_p & v1445782 | !hmaster1_p & v1445e1b;
assign v1445f4b = hbusreq2_p & v1445f48 | !hbusreq2_p & v1445f4a;
assign v12165a0 = hgrant4_p & v1216a98 | !hgrant4_p & v121659f;
assign v140589b = hbusreq1_p & v1405898 | !hbusreq1_p & v140589a;
assign v1215460 = hbusreq4 & v12164d3 | !hbusreq4 & v845542;
assign v14462ff = hmaster0_p & v14462f5 | !hmaster0_p & v14462fe;
assign d30800 = hgrant5_p & d306e6 | !hgrant5_p & d307ff;
assign v10d4272 = hmaster2_p & v10d426b | !hmaster2_p & v10d403a;
assign d2f9a3 = hbusreq5_p & d2fec1 | !hbusreq5_p & d2f9a2;
assign v12160f3 = hbusreq4_p & v12160f2 | !hbusreq4_p & !v845542;
assign d80760 = locked_p & d8075c | !locked_p & d8075f;
assign d307b9 = hgrant5_p & d307ad | !hgrant5_p & d307b8;
assign v1446562 = hmaster0_p & v144655a | !hmaster0_p & v1446561;
assign v12afdad = hbusreq4_p & v12afdab | !hbusreq4_p & v12afdac;
assign v12153bb = hbusreq0_p & v1215bb0 | !hbusreq0_p & v12160f2;
assign v1215768 = hbusreq4_p & v1215767 | !hbusreq4_p & v845542;
assign v1214fbe = hbusreq0 & v121579c | !hbusreq0 & v1214fbd;
assign v1515ae2 = hgrant2_p & v1515ae1 | !hgrant2_p & !v845542;
assign v1515750 = hgrant1_p & v151574f | !hgrant1_p & v1515747;
assign d307e3 = hlock1_p & d307e2 | !hlock1_p & d30658;
assign v138a307 = hbusreq2_p & v138a302 | !hbusreq2_p & v138a306;
assign v1216312 = hbusreq2_p & v121630f | !hbusreq2_p & v1216307;
assign v1214fb5 = hgrant5_p & v845542 | !hgrant5_p & v1214fb4;
assign v1446555 = hgrant2_p & v14464a8 | !hgrant2_p & v14464a2;
assign a65635 = hbusreq0 & a65626 | !hbusreq0 & a65634;
assign v134d38c = hbusreq5_p & v134d388 | !hbusreq5_p & v134d38b;
assign a658ef = hmaster0_p & a658b7 | !hmaster0_p & a658ee;
assign d2f9a0 = hbusreq4_p & d2febf | !hbusreq4_p & v84554a;
assign v14459dc = hmaster2_p & v14459db | !hmaster2_p & v14459cf;
assign v15157eb = hbusreq5_p & v15157e9 | !hbusreq5_p & !v15157ea;
assign v144634b = hlock2 & v144632f | !hlock2 & v1446349;
assign d301c8 = hbusreq5_p & d301c6 | !hbusreq5_p & d301c7;
assign v11e5944 = hgrant0_p & v845542 | !hgrant0_p & !v11e593a;
assign v1445f9d = hlock0 & v1445f9a | !hlock0 & v1445f9c;
assign v1446713 = hmaster1_p & v1446712 | !hmaster1_p & v1446436;
assign d3022c = hbusreq0 & d30226 | !hbusreq0 & d3022b;
assign a65419 = hgrant5_p & a6587e | !hgrant5_p & a6538a;
assign f2e27b = hready_p & v845542 | !hready_p & f2e27a;
assign v12160f4 = hgrant4_p & v12160f3 | !hgrant4_p & v12afe44;
assign v1445bfe = jx1_p & v144620b | !jx1_p & v1445bfa;
assign v1515723 = hgrant1_p & v1515712 | !hgrant1_p & v1515722;
assign v15532c3 = hgrant5_p & v1553225 | !hgrant5_p & v15532c2;
assign v1445ef8 = hmaster1_p & v1445ecd | !hmaster1_p & v1445ef0;
assign v12af7f6 = hmaster2_p & v12af7f5 | !hmaster2_p & d30690;
assign v10d4279 = hbusreq2_p & v10d4271 | !hbusreq2_p & !v10d4278;
assign v12165b1 = hgrant2_p & v12165ab | !hgrant2_p & v12165b0;
assign d301fe = hgrant1_p & d301f3 | !hgrant1_p & d307bb;
assign v151574d = hbusreq1 & v151560d | !hbusreq1 & v845570;
assign v1445520 = hmaster1_p & v1445506 | !hmaster1_p & v1445b7a;
assign v1515650 = hmaster0_p & v151564e | !hmaster0_p & v151564f;
assign v14459bd = hlock4 & v144639c | !hlock4 & v14459bc;
assign v1552d5e = hbusreq0 & v1552d5d | !hbusreq0 & v1553395;
assign v12ad680 = hmaster2_p & v12ad678 | !hmaster2_p & !v12ad67f;
assign d2fcad = hbusreq1 & d305ea | !hbusreq1 & !d305ef;
assign v1216045 = hbusreq2_p & v1216042 | !hbusreq2_p & v1216044;
assign d3066d = hmaster0_p & d30657 | !hmaster0_p & d3066c;
assign v14465aa = hmaster0_p & v1446404 | !hmaster0_p & v144639c;
assign v121620b = hmaster2_p & v12161d0 | !hmaster2_p & v845542;
assign v12163a7 = hmaster2_p & v12163a5 | !hmaster2_p & !v1216acd;
assign d2fbf9 = hgrant5_p & v84554a | !hgrant5_p & d2fbf7;
assign v1215016 = hmaster0_p & v1215001 | !hmaster0_p & v1215015;
assign v12167a8 = hmaster1_p & v12165ae | !hmaster1_p & v12165a5;
assign v10d402b = locked_p & v10d3fde | !locked_p & v10d3fdf;
assign v1445ba3 = hbusreq2 & v1445b9b | !hbusreq2 & v1445b9e;
assign d2fb03 = hbusreq1_p & d300fd | !hbusreq1_p & d2fb02;
assign v12ad030 = hbusreq2_p & v12ad023 | !hbusreq2_p & v12ad02f;
assign v16a1bed = hbusreq5 & v16a1bdf | !hbusreq5 & v16a1bec;
assign v1446130 = hlock2 & v144612c | !hlock2 & v144612f;
assign v1216abd = hlock1_p & v1216abc | !hlock1_p & v845547;
assign v1284d4b = hbusreq1_p & v1284cc6 | !hbusreq1_p & v1284d4a;
assign d2fb51 = hbusreq0 & d2fb4d | !hbusreq0 & v845542;
assign v134d3dc = hgrant4_p & v845542 | !hgrant4_p & v134d3db;
assign v1216a6b = hlock5_p & v1216a5a | !hlock5_p & v845542;
assign v1668d9e = hgrant5_p & v1668d97 | !hgrant5_p & v1668d9d;
assign a65687 = hmaster0_p & a658e8 | !hmaster0_p & a658ee;
assign v1445787 = hlock2 & v1445786 | !hlock2 & v1445780;
assign v1552fd0 = hbusreq3 & v1552fcf | !hbusreq3 & v155321a;
assign v144578b = hlock0 & v144578a | !hlock0 & v1445789;
assign v134ce7e = hgrant3_p & v134ce7b | !hgrant3_p & v134ce7d;
assign v134cebe = hlock5 & v134d270 | !hlock5 & v134cebd;
assign d3010a = hgrant5_p & d2fea1 | !hgrant5_p & d30108;
assign v138a30f = hlock5_p & v10d3ff1 | !hlock5_p & !v845542;
assign v14466cc = hmaster0_p & v14463c9 | !hmaster0_p & v144639c;
assign a65410 = hbusreq2_p & a6540b | !hbusreq2_p & !a6540f;
assign v1445e1a = hlock2 & v1445e0f | !hlock2 & v1445e19;
assign v1445e76 = stateG10_5_p & v1445e6d | !stateG10_5_p & v1445e75;
assign v1214c29 = hlock0_p & v12164cf | !hlock0_p & v1214c28;
assign v16a19e1 = hmaster1_p & v16a19e0 | !hmaster1_p & v16a2672;
assign v14459e3 = hbusreq5_p & v14459d1 | !hbusreq5_p & v14459e2;
assign v1216042 = hmaster1_p & v1216039 | !hmaster1_p & v1216041;
assign v144610b = hmaster1_p & v14460f7 | !hmaster1_p & v1445fbd;
assign v140588b = hbusreq4_p & v140588a | !hbusreq4_p & v140583c;
assign v121538a = hbusreq0 & d2fbe5 | !hbusreq0 & v845542;
assign d80776 = hgrant5_p & v845542 | !hgrant5_p & d80774;
assign d301e0 = hbusreq5_p & d301df | !hbusreq5_p & !d301de;
assign d2fb92 = hbusreq2_p & d2fb91 | !hbusreq2_p & d2fb90;
assign v1214c2c = hbusreq0 & v1214c2b | !hbusreq0 & v16a2243;
assign d30825 = hbusreq5_p & d30821 | !hbusreq5_p & d30824;
assign d30676 = hlock2_p & d30675 | !hlock2_p & v84555e;
assign v16a207a = hgrant5_p & v845542 | !hgrant5_p & v16a206f;
assign d80739 = busreq_p & d80730 | !busreq_p & !v8b8a8c;
assign bf1f59 = hmaster1_p & bf1f58 | !hmaster1_p & v845542;
assign v1389810 = hbusreq5_p & v138980f | !hbusreq5_p & !v845542;
assign v1445ab1 = hmaster1_p & v1445ab0 | !hmaster1_p & v144589f;
assign v11e5953 = hbusreq4_p & v11e5952 | !hbusreq4_p & v845570;
assign a653e6 = hbusreq0 & a653d6 | !hbusreq0 & a653e5;
assign v1405869 = hgrant5_p & v1405865 | !hgrant5_p & v1405868;
assign v1284d07 = hmaster0_p & v140587e | !hmaster0_p & v1284cb9;
assign v121532d = hbusreq2_p & v121532c | !hbusreq2_p & v1215326;
assign v16a1da3 = hmaster1_p & v16a1ac9 | !hmaster1_p & v16a2672;
assign v9745f6 = hmaster1_p & v9109e4 | !hmaster1_p & v845542;
assign v12162ed = hbusreq1_p & v12162ec | !hbusreq1_p & v845547;
assign v1445a05 = hgrant5_p & v14459d4 | !hgrant5_p & v1445a04;
assign v14460a4 = hbusreq0 & v14460a3 | !hbusreq0 & v1446077;
assign v1446154 = hbusreq2_p & v1446152 | !hbusreq2_p & v1446153;
assign v1284d10 = hgrant1_p & v1284c8f | !hgrant1_p & v14465da;
assign v1215d81 = hmaster0_p & v1215d6c | !hmaster0_p & v1215d80;
assign v1284d3c = hmaster2_p & v1284d3b | !hmaster2_p & v144639e;
assign v134d22d = hmaster1_p & v134d22c | !hmaster1_p & v134d208;
assign v16a1417 = hgrant2_p & v16a1dff | !hgrant2_p & v16a1416;
assign v1216265 = hgrant2_p & v1216229 | !hgrant2_p & v1216264;
assign v1215d29 = hmaster2_p & v845570 | !hmaster2_p & v1216a93;
assign v12161f0 = hbusreq1_p & v12161ef | !hbusreq1_p & v845542;
assign d305d5 = hbusreq5_p & d305d4 | !hbusreq5_p & v845542;
assign v10d408f = hmaster0_p & v10d400b | !hmaster0_p & v10d3ffd;
assign v1389371 = hmaster1_p & v845542 | !hmaster1_p & v1389370;
assign a65620 = hgrant1_p & a65362 | !hgrant1_p & !a6561f;
assign v1552f65 = hmaster2_p & v15533a5 | !hmaster2_p & v1552f64;
assign v16a1dc0 = hmaster1_p & v9337f3 | !hmaster1_p & v16a2672;
assign v1216254 = hbusreq2 & v1216250 | !hbusreq2 & v1216253;
assign v134cd88 = hlock3 & v134d3b5 | !hlock3 & v134cd87;
assign v15161d4 = hgrant2_p & v15161d3 | !hgrant2_p & !v845542;
assign v134cd57 = hlock1 & v134d273 | !hlock1 & v134cd56;
assign v1668dcc = hgrant5_p & v845542 | !hgrant5_p & !v1668d7d;
assign v1216035 = hmaster2_p & f2f2a8 | !hmaster2_p & v1216034;
assign v155339e = hbusreq1 & v155339b | !hbusreq1 & v155339d;
assign v1445a82 = hmaster0_p & v1445a81 | !hmaster0_p & v1445a31;
assign v10d4024 = hgrant1_p & v10d401f | !hgrant1_p & v10d4023;
assign v1553430 = hmaster1_p & v155342f | !hmaster1_p & v845542;
assign v1445a23 = hbusreq0_p & v1445a22 | !hbusreq0_p & v14465bb;
assign v134cd5d = hbusreq0 & v134cd5c | !hbusreq0 & v134d379;
assign v1216276 = hmaster1_p & v1216275 | !hmaster1_p & v1216041;
assign v1515753 = hbusreq5_p & v151574b | !hbusreq5_p & !v1515752;
assign v1216206 = hbusreq1_p & v1216205 | !hbusreq1_p & v845547;
assign v12acffb = hbusreq4_p & v12ad5a6 | !hbusreq4_p & v12acffa;
assign v1445e55 = hbusreq4_p & v14465be | !hbusreq4_p & v14465bb;
assign v121605a = hbusreq1_p & v1216059 | !hbusreq1_p & v845542;
assign v144655c = hgrant1_p & v845542 | !hgrant1_p & v144655b;
assign f2f3ae = hmaster1_p & f2f3ad | !hmaster1_p & f2f2ae;
assign v1216125 = hbusreq1_p & v1216124 | !hbusreq1_p & v845542;
assign d2f979 = hbusreq4_p & d2fea1 | !hbusreq4_p & !v845542;
assign v138a32b = hmastlock_p & v138a328 | !hmastlock_p & !v138a32a;
assign v138a3f7 = hlock5_p & v1668dab | !hlock5_p & v845542;
assign v1515832 = hmaster2_p & v1515609 | !hmaster2_p & v151560d;
assign v1215be7 = hmaster2_p & v845547 | !hmaster2_p & v1215be6;
assign v14466ff = hmaster1_p & v14466fe | !hmaster1_p & v144644d;
assign v134d371 = hlock1 & v134d273 | !hlock1 & v134d370;
assign v1215fb8 = hmaster1_p & v12166f7 | !hmaster1_p & v12166ef;
assign d3063a = hlock2_p & d30639 | !hlock2_p & d30635;
assign v1445fb4 = hbusreq2 & v1445fad | !hbusreq2 & v1445fb3;
assign v16a2064 = hbusreq3 & v16a2061 | !hbusreq3 & v16a2063;
assign v1284d11 = hmaster2_p & v14465b3 | !hmaster2_p & v1284d10;
assign v1216097 = hmaster0_p & v1216096 | !hmaster0_p & v121605c;
assign v16a1dab = hbusreq2 & v16a1daa | !hbusreq2 & v16a205c;
assign v1216a7c = hmaster1_p & v1216a7b | !hmaster1_p & v845542;
assign v1445b47 = hmaster0_p & v1445a3e | !hmaster0_p & v14459a2;
assign v121617b = hgrant5_p & v1216029 | !hgrant5_p & !v1216179;
assign v138a45e = hmaster0_p & v138a354 | !hmaster0_p & v138a34f;
assign v1446656 = hbusreq0 & v1446655 | !hbusreq0 & v1446638;
assign v134d495 = hbusreq0 & v134d376 | !hbusreq0 & v134d379;
assign v16a1bc4 = hbusreq1_p & v16a1bc3 | !hbusreq1_p & v16a2089;
assign v1446072 = hlock0 & v1446067 | !hlock0 & v1446071;
assign v1445fa3 = hmaster0_p & v144639c | !hmaster0_p & v1445fa2;
assign v1405890 = hgrant4_p & v140588b | !hgrant4_p & v140588f;
assign v1214bf5 = hbusreq2_p & v1214bf4 | !hbusreq2_p & v1214bf3;
assign v1445850 = hbusreq2_p & v1445844 | !hbusreq2_p & v144584f;
assign f2f289 = hbusreq5_p & f2f232 | !hbusreq5_p & f2f288;
assign v134d4d0 = hgrant5_p & v134d4cf | !hgrant5_p & v134d4cd;
assign v144552d = hbusreq2_p & v144552c | !hbusreq2_p & v1445bdb;
assign v12af21f = hbusreq5_p & v12af590 | !hbusreq5_p & v12af21e;
assign v1216142 = hbusreq1_p & v1216141 | !hbusreq1_p & v845542;
assign d30756 = hmaster1_p & d3072f | !hmaster1_p & d30754;
assign v14458d2 = hlock0_p & v845542 | !hlock0_p & v144639c;
assign v15156f2 = hmaster0_p & v15156f1 | !hmaster0_p & v151564f;
assign a65663 = hmaster1_p & a65661 | !hmaster1_p & a65439;
assign f2f228 = hgrant1_p & f2f227 | !hgrant1_p & !v845542;
assign v121600b = hmaster2_p & v1216002 | !hmaster2_p & v121600a;
assign d2fb1c = hbusreq5_p & d30153 | !hbusreq5_p & d2fb1b;
assign v1668d6b = hburst0 & a66293 | !hburst0 & v1668d6a;
assign v1445835 = hmaster1_p & v144580e | !hmaster1_p & v1445e28;
assign v14465df = hmaster2_p & v144639c | !hmaster2_p & v1446415;
assign v1214d31 = hbusreq5 & v1214d19 | !hbusreq5 & v1214d30;
assign v1389444 = hbusreq1_p & v15168ad | !hbusreq1_p & v1515c7d;
assign v138a35b = hmaster0_p & v138a34b | !hmaster0_p & v138a344;
assign v16a2674 = hmaster2_p & v16a2668 | !hmaster2_p & v845542;
assign v1215373 = hbusreq3 & v121536f | !hbusreq3 & v1215372;
assign v121503b = hmaster2_p & v121502e | !hmaster2_p & v121503a;
assign v1214bbe = hmaster1_p & v1214bbd | !hmaster1_p & v12153a9;
assign v1445558 = jx0_p & v1445bfe | !jx0_p & v1445557;
assign v1216293 = hgrant2_p & v1216284 | !hgrant2_p & v1216292;
assign v1215c20 = hmaster2_p & v1215c1f | !hmaster2_p & v1215c1a;
assign v1214d6f = hmaster0_p & v1214d08 | !hmaster0_p & v1214c3c;
assign v1215c06 = hmaster0_p & v1215bfb | !hmaster0_p & v1215c05;
assign v144577e = hmaster0_p & v1445778 | !hmaster0_p & v1445e13;
assign v121670c = hmaster1_p & v121670b | !hmaster1_p & v12166ef;
assign a6540e = hmaster1_p & a6540d | !hmaster1_p & a1db63;
assign v1214f6b = decide_p & v1216a82 | !decide_p & v1214f6a;
assign v134d30f = hgrant0_p & v134d1dd | !hgrant0_p & v845542;
assign v15157a1 = hmaster2_p & v1515793 | !hmaster2_p & v845542;
assign v16a1d2a = hbusreq5 & v16a1d25 | !hbusreq5 & v16a1d29;
assign d2feb6 = hlock4_p & d30740 | !hlock4_p & !v16693aa;
assign d2fb43 = hmaster1_p & d2f99c | !hmaster1_p & d2fb42;
assign v12160e6 = decide_p & v12160cf | !decide_p & v12160e5;
assign v1214cd9 = hmaster1_p & v1214cc1 | !hmaster1_p & v1214cd8;
assign v1445a3a = hmaster1_p & v1445a39 | !hmaster1_p & v14458fd;
assign d80740 = hlock5_p & d8073e | !hlock5_p & !d8073f;
assign d2fbec = hgrant4_p & d2fbea | !hgrant4_p & d2fbeb;
assign v1216559 = hgrant1_p & v1216522 | !hgrant1_p & v1216558;
assign v1215bff = hgrant5_p & v1215be4 | !hgrant5_p & !v1215bfd;
assign v12160cd = hbusreq3 & v12160c2 | !hbusreq3 & v12160cc;
assign v15156cc = hbusreq2_p & v15156cb | !hbusreq2_p & v845542;
assign v12150a0 = hbusreq4_p & v121509f | !hbusreq4_p & !v845542;
assign v134d3c1 = hbusreq1_p & v134d1e8 | !hbusreq1_p & v134d3c0;
assign v1405ada = hlock1_p & v1405a88 | !hlock1_p & !v845542;
assign v144615f = decide_p & v1446117 | !decide_p & v144615e;
assign v1668d34 = hbusreq0 & v1668d2d | !hbusreq0 & v1668d33;
assign d308a0 = hbusreq1_p & d307d9 | !hbusreq1_p & d306a5;
assign v12acff5 = hgrant2_p & v12acff2 | !hgrant2_p & v12acff4;
assign d3076a = hlock2_p & d30768 | !hlock2_p & d30769;
assign v1215c5b = hmaster2_p & v1216568 | !hmaster2_p & v845542;
assign v14461d9 = hbusreq2_p & v14461c4 | !hbusreq2_p & v14461d8;
assign v140587d = hmaster2_p & v140587c | !hmaster2_p & v140583f;
assign v134d49b = hmaster1_p & v134d369 | !hmaster1_p & v134d49a;
assign v1445408 = hmaster1_p & v1446466 | !hmaster1_p & v1445407;
assign v12ad615 = hbusreq5_p & v12ad613 | !hbusreq5_p & !v12ad614;
assign v1214c14 = hlock2_p & v1214c12 | !hlock2_p & v1214c13;
assign v1668d8a = hbusreq0 & v1668d81 | !hbusreq0 & v1668d89;
assign v16a1a81 = hbusreq2_p & v16a195e | !hbusreq2_p & v16a1a80;
assign v14460e9 = hmaster1_p & v1445fa2 | !hmaster1_p & v1445f9e;
assign a656d0 = hbusreq2_p & a656c2 | !hbusreq2_p & a656cf;
assign d2fbe9 = hlock4_p & d2fbe6 | !hlock4_p & v84554a;
assign v16a1cc7 = decide_p & v16a1b6b | !decide_p & !v16a1cc6;
assign v16695b9 = hbusreq2_p & v16695a1 | !hbusreq2_p & a7c7c1;
assign v1405af9 = hmaster1_p & v1405af8 | !hmaster1_p & v1405af0;
assign v16a1ad4 = hbusreq3 & v16a1acf | !hbusreq3 & !v16a1ad3;
assign v14466af = hlock0 & v14466ae | !hlock0 & v14466ad;
assign v1446011 = hbusreq1_p & v144647e | !hbusreq1_p & v144648d;
assign bf1f4e = hmaster0_p & bf1f4d | !hmaster0_p & v845542;
assign v134d287 = hgrant5_p & v845542 | !hgrant5_p & v134d285;
assign v1668d66 = hburst0_p & v845542 | !hburst0_p & !v1553930;
assign v14457aa = hlock2 & v1445786 | !hlock2 & v14457a8;
assign v1215435 = hready & v845542 | !hready & a658aa;
assign v10d4033 = hmaster2_p & v10d4024 | !hmaster2_p & !v10d4032;
assign f2f37e = hgrant1_p & v845570 | !hgrant1_p & !f2f37d;
assign v1214ed0 = hgrant5_p & v1214dcc | !hgrant5_p & v1214ecf;
assign hmaster0 = v10a1543;
assign v12ad4dd = hmaster0_p & v12ad4d9 | !hmaster0_p & v12ad4dc;
assign v13897dd = hmaster2_p & v166939b | !hmaster2_p & v845570;
assign a653c6 = hbusreq1 & a653c5 | !hbusreq1 & !v845558;
assign v12af1bb = hbusreq5_p & v12af3a5 | !hbusreq5_p & v12af1ba;
assign d300db = hlock4_p & d307b2 | !hlock4_p & a65382;
assign v1388ce8 = jx1_p & v1389411 | !jx1_p & v1388ce7;
assign d2fedc = hmaster0_p & d2fed5 | !hmaster0_p & d2fecf;
assign v1214c05 = hmaster0_p & v1214bb7 | !hmaster0_p & v1215396;
assign v1445b1b = hlock2 & v1445b18 | !hlock2 & v1445b1a;
assign d3074b = hmaster0_p & d30744 | !hmaster0_p & d30735;
assign v1216178 = hbusreq5_p & v1216176 | !hbusreq5_p & !v1216177;
assign v14453e3 = hbusreq2_p & v144621a | !hbusreq2_p & v14453e2;
assign v1515811 = hbusreq2 & v1515810 | !hbusreq2 & v845542;
assign f2f379 = hbusreq1 & v1668d71 | !hbusreq1 & v845542;
assign v1215b9b = hmaster0_p & v1215b98 | !hmaster0_p & v1215b9a;
assign v16a16a5 = hgrant5_p & v845542 | !hgrant5_p & !v16a1e90;
assign v1668c2c = hmaster1_p & v1668c2b | !hmaster1_p & v845542;
assign v14458c0 = hlock0 & v1445880 | !hlock0 & v14458bf;
assign v1445de9 = hbusreq4_p & v144640a | !hbusreq4_p & v1446406;
assign v1446299 = hlock2 & v1446293 | !hlock2 & v1446298;
assign v134ce63 = hmaster1_p & v134d369 | !hmaster1_p & v134ce62;
assign afe156 = hburst1_p & v906a5a | !hburst1_p & v8af912;
assign v1284cfb = hmaster2_p & v1284cf5 | !hmaster2_p & v1284cfa;
assign v134d20c = hmaster1_p & v134d20b | !hmaster1_p & v134d208;
assign v1216585 = hmaster1_p & v1216584 | !hmaster1_p & v1216a9b;
assign v14465f2 = hgrant4_p & v144639c | !hgrant4_p & v14465f1;
assign d2fc09 = hgrant2_p & d2fc08 | !hgrant2_p & d2fbfe;
assign v11e5980 = decide_p & v11e597f | !decide_p & v11e596d;
assign v1446448 = hlock0 & v1446447 | !hlock0 & v1446446;
assign v1216a76 = hmastlock_p & v1216a75 | !hmastlock_p & v845542;
assign v1445afa = hmaster0_p & v1445a4f | !hmaster0_p & v1445909;
assign v151565a = hmaster2_p & a658c6 | !hmaster2_p & !v1515658;
assign v1668d4d = hmaster2_p & v1668d36 | !hmaster2_p & v1668d4c;
assign v138a49f = decide_p & v138a475 | !decide_p & !v138a406;
assign v138a47d = hmaster0_p & v138a43a | !hmaster0_p & v138a439;
assign v16a1ca2 = hgrant2_p & v16a2059 | !hgrant2_p & v16a1ca1;
assign v134d496 = hlock0 & v134d495 | !hlock0 & v134d376;
assign a653fe = hgrant5_p & a65878 | !hgrant5_p & a653fd;
assign v14058c7 = hgrant1_p & v14058c6 | !hgrant1_p & v1405845;
assign v14460bb = hgrant2_p & v14460b9 | !hgrant2_p & v14460ba;
assign v12ad4d3 = hmaster0_p & v12ad4ce | !hmaster0_p & v12ad4d2;
assign v1389de6 = hlock5_p & v1389de5 | !hlock5_p & !v845542;
assign v1216112 = hmaster2_p & v121610b | !hmaster2_p & v1216111;
assign v15161f9 = hmaster0_p & v1668da6 | !hmaster0_p & d305df;
assign v1215cbf = hgrant5_p & v845542 | !hgrant5_p & !v1215cbd;
assign v1405b3a = decide_p & v1405b39 | !decide_p & v1405a99;
assign v16a1a7d = hmaster1_p & v16a1a7c | !hmaster1_p & v16a195b;
assign v12ad50d = decide_p & v12ad50c | !decide_p & v845542;
assign v14457b2 = hbusreq2_p & v14457ae | !hbusreq2_p & v14457b1;
assign v12166fa = hgrant2_p & v12166f5 | !hgrant2_p & v12166f9;
assign v121510d = hmaster1_p & v121510c | !hmaster1_p & v121546f;
assign v14453b4 = hmaster1_p & v1445366 | !hmaster1_p & v1445a9b;
assign v1446349 = hbusreq2_p & v1446343 | !hbusreq2_p & v1446348;
assign v12ad66b = hmaster0_p & v12ad528 | !hmaster0_p & v12ad517;
assign v1446667 = hbusreq2_p & v1446632 | !hbusreq2_p & v1446666;
assign f2f41e = hgrant1_p & f2f281 | !hgrant1_p & !f2f368;
assign v10d40d0 = decide_p & v10d40c7 | !decide_p & v10d40cf;
assign v1445bec = hmaster1_p & v1445beb | !hmaster1_p & v1446271;
assign v1445ec3 = hlock0 & v1445ec2 | !hlock0 & v1445ec1;
assign v1445531 = hbusreq2_p & v1445530 | !hbusreq2_p & v1445bdb;
assign f2e710 = hbusreq1 & v166939b | !hbusreq1 & !v166939f;
assign v12150dd = hbusreq2_p & v12150d4 | !hbusreq2_p & v12150d3;
assign v1446435 = hlock0 & v144642e | !hlock0 & v1446434;
assign v12afe4d = hgrant0_p & d3065a | !hgrant0_p & !v845542;
assign v1215ffd = hbusreq4_p & v1216a5a | !hbusreq4_p & v1215ff8;
assign v1445fe9 = hbusreq0 & v1445fe8 | !hbusreq0 & v1445fe1;
assign v1668d46 = hbusreq1_p & v1668d44 | !hbusreq1_p & !v1668d45;
assign v144536e = hbusreq2_p & v1445363 | !hbusreq2_p & v144536d;
assign v16a1bbd = hbusreq1_p & v16a1bbc | !hbusreq1_p & v16a206e;
assign v10d40bd = hgrant0_p & v10d401b | !hgrant0_p & !v10d40bc;
assign d307b0 = hbusreq4_p & d307af | !hbusreq4_p & v1668d48;
assign v14454ff = hbusreq2_p & v14454fe | !hbusreq2_p & v1445bdb;
assign f2f53d = hbusreq2_p & f2f52e | !hbusreq2_p & f2f53c;
assign v11e5963 = hgrant5_p & v11e5949 | !hgrant5_p & !v11e5962;
assign v1515839 = hgrant5_p & v10d3ffd | !hgrant5_p & v1515837;
assign v1215cfa = hmaster0_p & v1215cf4 | !hmaster0_p & v1215cf9;
assign v1284c8d = stateA1_p & v146b550 | !stateA1_p & !v85e70d;
assign v12152e5 = hmaster1_p & v12152e4 | !hmaster1_p & v1215b88;
assign v12ad4fa = hbusreq5_p & v12ad4f8 | !hbusreq5_p & !v12ad4f9;
assign d2fc33 = hbusreq5_p & v845542 | !hbusreq5_p & !d2fc32;
assign v12ad1fd = hbusreq2 & v12ad1fc | !hbusreq2 & v12af9b6;
assign v1215028 = hbusreq4_p & v1215027 | !hbusreq4_p & v845547;
assign v1445538 = decide_p & v1445468 | !decide_p & v1445537;
assign v14838be = hready_p & v14838bc | !hready_p & v14838bd;
assign v16a1d8c = hgrant5_p & v845568 | !hgrant5_p & v16a223e;
assign v134d314 = hmaster0_p & v134d30c | !hmaster0_p & v134d313;
assign v1405887 = hlock2_p & v1405884 | !hlock2_p & v1405886;
assign v121576b = hmaster2_p & v845542 | !hmaster2_p & v121576a;
assign v1215c71 = hbusreq0 & v1215c6f | !hbusreq0 & v1215c70;
assign v15157f9 = hmaster0_p & v15157f1 | !hmaster0_p & v15157f8;
assign v1389ff2 = hgrant2_p & v845542 | !hgrant2_p & !v1389de1;
assign d300bb = hlock4_p & d30785 | !hlock4_p & d300ba;
assign f2f2dd = hmaster2_p & f2f2c9 | !hmaster2_p & !f2f2cf;
assign v121629e = hgrant2_p & v12161a7 | !hgrant2_p & v121629d;
assign v1446721 = hlock5 & v1446700 | !hlock5 & v1446720;
assign v134ce74 = hlock2 & v134d276 | !hlock2 & v134ce73;
assign v144553b = hready_p & v144540b | !hready_p & v1445538;
assign v1515639 = hmaster2_p & v10d3fd4 | !hmaster2_p & v845542;
assign v121631a = hbusreq5_p & v1216319 | !hbusreq5_p & v12162ef;
assign v16a1cff = hbusreq5 & v16a1cf5 | !hbusreq5 & v16a1cfe;
assign a658e3 = hbusreq0 & a658d8 | !hbusreq0 & a658e2;
assign v1215771 = hmaster1_p & v1215730 | !hmaster1_p & v1215770;
assign v16a1e8d = hgrant4_p & v845559 | !hgrant4_p & v16a1e8c;
assign v12aeb84 = decide_p & v12aeb83 | !decide_p & v845542;
assign v14453c0 = hlock3 & v1445354 | !hlock3 & v14453be;
assign v1214e5b = hmaster1_p & v1214e5a | !hmaster1_p & v1214e0f;
assign v1515c81 = hmaster2_p & v845542 | !hmaster2_p & v1515c80;
assign f2f3d4 = hbusreq5_p & f2f3d2 | !hbusreq5_p & !f2f3d3;
assign v12160ec = hbusreq4 & v121601c | !hbusreq4 & !v845542;
assign v14462ef = hbusreq5_p & v14462ea | !hbusreq5_p & v14462ee;
assign d302ef = hgrant3_p & d302dd | !hgrant3_p & !d302ee;
assign v1445bc8 = hgrant2_p & v1445bc7 | !hgrant2_p & v1445bc4;
assign v12aeb75 = hmaster2_p & v845542 | !hmaster2_p & v12aeb74;
assign v1445fee = hlock2 & v1445fe6 | !hlock2 & v1445fed;
assign v1445b40 = hmaster0_p & v1445a43 | !hmaster0_p & v1445a5a;
assign v1446289 = hbusreq2 & v1446287 | !hbusreq2 & v1446288;
assign a65627 = hgrant4_p & a662a9 | !hgrant4_p & !a6537f;
assign v1215cff = hgrant5_p & v845542 | !hgrant5_p & v1215c87;
assign v12ad5bd = hbusreq1_p & v12ad5b9 | !hbusreq1_p & !v12ad5bc;
assign v134d20d = hlock2_p & v134d209 | !hlock2_p & v134d20c;
assign d2f97f = hbusreq2_p & d30167 | !hbusreq2_p & d2f97e;
assign v16a1e49 = hbusreq2 & v16a1e2e | !hbusreq2 & v16a1e30;
assign d2fb5c = hmaster1_p & d2fb5b | !hmaster1_p & d2fb55;
assign v12163ab = hmaster1_p & v845542 | !hmaster1_p & !v12163a9;
assign a66284 = hbusreq4_p & a66283 | !hbusreq4_p & !v845542;
assign v1405ae1 = hmaster2_p & d3070c | !hmaster2_p & !v1405a8c;
assign v1446478 = hbusreq1_p & v1446398 | !hbusreq1_p & v1446476;
assign v144599b = hlock1 & v144599a | !hlock1 & v1445999;
assign d3014a = hgrant5_p & v84555a | !hgrant5_p & d30108;
assign v15167ed = hbusreq2_p & v15167ec | !hbusreq2_p & v845542;
assign v12ad8e3 = hbusreq4_p & v12afda1 | !hbusreq4_p & v12af983;
assign v1214bf2 = hmaster0_p & v12153b1 | !hmaster0_p & v1214bf1;
assign v1445ff7 = hbusreq3 & v1445ff5 | !hbusreq3 & v1445ff6;
assign v12acfc0 = hlock2_p & v12acfbd | !hlock2_p & v12acfbf;
assign v16a1bb5 = hburst1 & v16a1bb4 | !hburst1 & v845542;
assign v16a1e77 = hbusreq2_p & v16a1dd7 | !hbusreq2_p & v16a1e76;
assign v16a1331 = hgrant2_p & v16a2059 | !hgrant2_p & v16a1330;
assign v1553058 = hgrant4_p & v1553057 | !hgrant4_p & v845542;
assign v14463b7 = hbusreq1 & v14463b3 | !hbusreq1 & v14463b6;
assign v134d1e4 = hburst0_p & v845584 | !hburst0_p & v134d1e3;
assign v1215048 = hmaster2_p & v845542 | !hmaster2_p & v1215047;
assign v15532c2 = hmaster2_p & v845542 | !hmaster2_p & v15532c1;
assign v1284d21 = hgrant2_p & v1284d08 | !hgrant2_p & v1284d20;
assign f2f418 = hmaster0_p & f2f3a8 | !hmaster0_p & f2f35d;
assign v1216b02 = hlock5_p & v1216b00 | !hlock5_p & !v1216b01;
assign d300b9 = hbusreq4 & d3078d | !hbusreq4 & !d30645;
assign d2fe8b = hmaster2_p & v845542 | !hmaster2_p & d2fe8a;
assign d3083c = hmaster0_p & d3081d | !hmaster0_p & d3083b;
assign v16a1ae9 = hmaster1_p & v16a1ae8 | !hmaster1_p & v16a209c;
assign v16a1389 = hbusreq2 & v16a1385 | !hbusreq2 & v16a1388;
assign d3074a = hbusreq2_p & d30749 | !hbusreq2_p & d30748;
assign v1552d56 = hbusreq2_p & v1552d4e | !hbusreq2_p & v1552d55;
assign v12150b1 = hbusreq5 & v1215076 | !hbusreq5 & v12150b0;
assign v134d28e = hlock0_p & v134d1dd | !hlock0_p & v845542;
assign v1668d88 = hgrant5_p & v1668d7f | !hgrant5_p & v1668d86;
assign v15157ab = hgrant5_p & v15157a6 | !hgrant5_p & v15157aa;
assign v134d264 = hbusreq2_p & v134d263 | !hbusreq2_p & v134d262;
assign v1405a94 = hmaster0_p & v1405a8f | !hmaster0_p & v1405a93;
assign v1216598 = hgrant5_p & v845542 | !hgrant5_p & v1216597;
assign d3025c = hgrant2_p & d30234 | !hgrant2_p & d30251;
assign d305f3 = hbusreq1 & d305ea | !hbusreq1 & !d305f2;
assign d30684 = hbusreq5_p & v84555e | !hbusreq5_p & !v845542;
assign d2fe94 = hmaster2_p & d2fe80 | !hmaster2_p & !d2fe93;
assign d3086a = hbusreq5_p & d30726 | !hbusreq5_p & d30869;
assign a6543a = hmaster1_p & a6541e | !hmaster1_p & a65439;
assign d30219 = hmaster1_p & d301e5 | !hmaster1_p & d30218;
assign v1214df5 = hmaster2_p & v845547 | !hmaster2_p & v1214df3;
assign v1405b32 = decide_p & v1405aba | !decide_p & v1405b31;
assign f2f42f = hgrant1_p & f2f281 | !hgrant1_p & !f2f37a;
assign v12adf63 = hbusreq0 & v12adf5e | !hbusreq0 & v12adf62;
assign v121659a = hbusreq4_p & v1216a8d | !hbusreq4_p & !v1216594;
assign v16a1bc1 = hgrant0_p & v845542 | !hgrant0_p & !v16a1bb9;
assign v1515c7b = hburst1 & v15168a9 | !hburst1 & f2f4ad;
assign v1214cf9 = hgrant1_p & v1214c30 | !hgrant1_p & v1214cf3;
assign a65af7 = hgrant3_p & a662c6 | !hgrant3_p & a65af6;
assign v14457de = hmaster1_p & v14457dd | !hmaster1_p & v1445e07;
assign d30627 = hbusreq3 & d30618 | !hbusreq3 & d30626;
assign v1216539 = hmaster2_p & v1216536 | !hmaster2_p & v1216538;
assign v1515626 = hmastlock_p & v1515625 | !hmastlock_p & !v845542;
assign v1215c47 = hmaster1_p & v1215c46 | !hmaster1_p & v1215c35;
assign v144585a = hbusreq2_p & v1445854 | !hbusreq2_p & v1445859;
assign v1215c2b = hgrant5_p & v1215be1 | !hgrant5_p & v1215c2a;
assign v10d4290 = hbusreq0_p & v10d428f | !hbusreq0_p & v10d3fdf;
assign d300cf = hgrant5_p & d2fe81 | !hgrant5_p & d300ce;
assign v144589c = hmaster2_p & v144589b | !hmaster2_p & v14463bb;
assign v1516218 = decide_p & v1516804 | !decide_p & v845576;
assign d30885 = hmaster0_p & d30850 | !hmaster0_p & d3084d;
assign a6592a = decide_p & a65929 | !decide_p & v845542;
assign v1669591 = decide_p & v16693b0 | !decide_p & v845542;
assign v134cea7 = hbusreq3 & v134cea1 | !hbusreq3 & v134cea6;
assign v12afdae = hgrant4_p & v12afdad | !hgrant4_p & v12afdab;
assign v1445514 = hgrant2_p & v14454e9 | !hgrant2_p & v1445513;
assign v1214da4 = hgrant2_p & v1214da2 | !hgrant2_p & v1214da3;
assign d30255 = hgrant5_p & v845542 | !hgrant5_p & d30221;
assign d2fb49 = hready_p & d2fb33 | !hready_p & d2fb48;
assign v1215d95 = hbusreq3 & v1215d8f | !hbusreq3 & v12164e7;
assign v1445a75 = hmaster2_p & v1445a49 | !hmaster2_p & v14458e5;
assign v16a1afd = hmaster2_p & v16a1afa | !hmaster2_p & !v845542;
assign d30643 = hlock2_p & d30642 | !hlock2_p & v84555e;
assign d2fec5 = hbusreq0 & d2fec1 | !hbusreq0 & d2fec4;
assign a6587b = hbusreq2_p & a65873 | !hbusreq2_p & a6587a;
assign v1215b81 = hbusreq1_p & v1215b7d | !hbusreq1_p & v1215b80;
assign v1216519 = decide_p & v12164ce | !decide_p & v1216518;
assign v1214c6e = hgrant1_p & v1214c68 | !hgrant1_p & v1214c6d;
assign a65672 = hbusreq5_p & a6542f | !hbusreq5_p & a65671;
assign v12ad017 = hmaster0_p & v12ad00e | !hmaster0_p & v12ad016;
assign v138a3cb = hbusreq0 & v138a3c7 | !hbusreq0 & v138a3ca;
assign v1214d43 = hmaster2_p & v845547 | !hmaster2_p & v1214d42;
assign v12161a7 = hmaster1_p & v12161a6 | !hmaster1_p & v845542;
assign d30689 = hbusreq1_p & v845542 | !hbusreq1_p & d30688;
assign v134cf6c = hgrant3_p & v134d3fc | !hgrant3_p & v134cf6b;
assign v1445e28 = hmaster0_p & v1445e27 | !hmaster0_p & v1445e06;
assign v14457f0 = hmaster1_p & v14457ef | !hmaster1_p & v1445ed3;
assign v10d4280 = locked_p & v10d427c | !locked_p & v10d427f;
assign v151583a = hbusreq5_p & v1515838 | !hbusreq5_p & v1515839;
assign v1214edf = hmaster2_p & v1216538 | !hmaster2_p & v121654a;
assign v1668cc8 = hmaster2_p & v845542 | !hmaster2_p & !v1668cc6;
assign v134d3d9 = hbusreq0_p & v134d1dd | !hbusreq0_p & v845542;
assign v12ad8eb = hbusreq0 & v12ad8e6 | !hbusreq0 & v12ad8ea;
assign a65661 = hmaster0_p & a65444 | !hmaster0_p & a6541e;
assign v1215bb7 = hbusreq2_p & v1215bb6 | !hbusreq2_p & v12163ab;
assign v121501c = hmaster2_p & v1214fe6 | !hmaster2_p & v1214ffe;
assign v144663a = hlock0 & v1446639 | !hlock0 & v1446637;
assign v138a3e4 = hmaster0_p & v138a30f | !hmaster0_p & v138a3e3;
assign d2f9b8 = hmaster2_p & d2feb2 | !hmaster2_p & d2f9b7;
assign v1445a9a = hlock0 & v1445a98 | !hlock0 & v1445a99;
assign v16a1bd4 = hbusreq1 & v16a1bd3 | !hbusreq1 & v16a206e;
assign v1445a70 = hlock2 & v1445a69 | !hlock2 & v1445a6f;
assign v144588c = hgrant5_p & v1445889 | !hgrant5_p & !v144588b;
assign v1445868 = decide_p & v1445774 | !decide_p & v1445867;
assign d30700 = hbusreq4_p & v845542 | !hbusreq4_p & a65861;
assign v1553394 = hmaster2_p & v845542 | !hmaster2_p & v1553393;
assign f2e274 = hbusreq1 & v16693a6 | !hbusreq1 & !f2e273;
assign a65b17 = hmaster1_p & a65b14 | !hmaster1_p & a65b09;
assign v134d3d0 = hmaster0_p & v134d3ad | !hmaster0_p & v845542;
assign d30149 = hgrant5_p & d2fe96 | !hgrant5_p & d30108;
assign a6542f = hgrant5_p & a65892 | !hgrant5_p & a653d1;
assign v12ad5e6 = hmaster0_p & v12ad4f4 | !hmaster0_p & v12ad5e5;
assign v1284d1d = hmaster2_p & v1284d19 | !hmaster2_p & v1284d1c;
assign v121537a = hmaster2_p & d2fbe5 | !hmaster2_p & v1215379;
assign v144601c = hmaster1_p & v144601b | !hmaster1_p & v845542;
assign v1446673 = hmaster0_p & v14465b8 | !hmaster0_p & v1446648;
assign bf1fa8 = decide_p & bf1fa7 | !decide_p & v845570;
assign v1445993 = locked_p & v144639c | !locked_p & v1445992;
assign d2fafc = hgrant5_p & d2faf2 | !hgrant5_p & d2fafb;
assign v1445a53 = hgrant1_p & v1445906 | !hgrant1_p & v1445a52;
assign v14461f3 = hgrant2_p & v14461ce | !hgrant2_p & v14461f2;
assign f2f45d = decide_p & f2f45c | !decide_p & f2f23c;
assign v12acfba = hmaster1_p & v12ad67b | !hmaster1_p & !v12acfb9;
assign a6562d = hbusreq1_p & a65387 | !hbusreq1_p & a6562c;
assign v16a1bcb = hgrant1_p & v84554d | !hgrant1_p & v16a1bca;
assign v12153fb = hmaster0_p & v12153f3 | !hmaster0_p & v12153ee;
assign v12162f3 = hbusreq0 & v1216adb | !hbusreq0 & v12162f2;
assign v16a209d = hgrant2_p & v845542 | !hgrant2_p & !v16a209c;
assign d308ea = hgrant2_p & d308e7 | !hgrant2_p & d308de;
assign v1214c0b = hmaster0_p & v1214bb7 | !hmaster0_p & v12153b1;
assign d302d2 = hready_p & d3029e | !hready_p & d301b9;
assign v16a1958 = hmaster2_p & v16a208a | !hmaster2_p & v16a194c;
assign v144623b = hmaster1_p & v144623a | !hmaster1_p & v1446236;
assign v1405a91 = hbusreq0_p & v845542 | !hbusreq0_p & !v1405a87;
assign d2fb50 = hbusreq0 & d2fb4f | !hbusreq0 & v845542;
assign v134d207 = hmaster2_p & v134d205 | !hmaster2_p & v134d206;
assign v1405af8 = hmaster0_p & v1405ad8 | !hmaster0_p & v1405af7;
assign v12ad525 = hmaster0_p & v12ad520 | !hmaster0_p & v12ad524;
assign v1215471 = hmaster2_p & v121545f | !hmaster2_p & v1215466;
assign v155322b = hgrant5_p & v845542 | !hgrant5_p & v1553229;
assign v121606e = hlock2_p & v121606a | !hlock2_p & v121606d;
assign v1445f75 = hbusreq2_p & v1445f71 | !hbusreq2_p & v1445f74;
assign v151580c = hmaster2_p & v10d3fd4 | !hmaster2_p & !v1515741;
assign d306f3 = locked_p & d306f2 | !locked_p & !v845542;
assign v1216aeb = hlock0_p & v1216aea | !hlock0_p & v845547;
assign v1445523 = hlock2 & v14454fa | !hlock2 & v1445522;
assign v12160ab = hbusreq2_p & v12160aa | !hbusreq2_p & v12160a9;
assign d306af = hbusreq1_p & d30661 | !hbusreq1_p & d306ae;
assign v16a1325 = hgrant4_p & v845542 | !hgrant4_p & v16a1324;
assign v121659f = hgrant0_p & v121659e | !hgrant0_p & !v845542;
assign v1215bb0 = hbusreq4 & v16a1bc6 | !hbusreq4 & v845542;
assign v1284cdd = hmaster2_p & v1284cd8 | !hmaster2_p & v1284cdc;
assign v134d44e = hlock0 & v134d44d | !hlock0 & v134d44c;
assign v134ce45 = hbusreq0 & v134ce44 | !hbusreq0 & v134d38b;
assign v1445ed8 = hmaster0_p & v14465b7 | !hmaster0_p & v1445eb8;
assign v144587c = hmaster2_p & v14463b1 | !hmaster2_p & !v1445879;
assign v15168b6 = hbusreq2 & v15168a8 | !hbusreq2 & v15168b5;
assign v16a1e22 = hmaster2_p & v16a1e21 | !hmaster2_p & !v845542;
assign v8b6f6a = jx1_p & v845542 | !jx1_p & !v845542;
assign v1445ebb = hmaster0_p & v14465b7 | !hmaster0_p & v1445eba;
assign v1445e22 = hlock3 & v1445e1f | !hlock3 & v1445e21;
assign v1668c26 = hlock3_p & v1668c25 | !hlock3_p & !v845542;
assign v1445f28 = hmaster1_p & v1445f27 | !hmaster1_p & v1445da4;
assign d308c9 = hgrant2_p & d30886 | !hgrant2_p & !d308c8;
assign v12161b4 = hbusreq2 & v12161a5 | !hbusreq2 & v12161b3;
assign v12153d7 = hbusreq4 & v1216adc | !hbusreq4 & !v845542;
assign v845547 = hready & v845542 | !hready & !v845542;
assign v138a34a = hlock5_p & v138a348 | !hlock5_p & v138a349;
assign v144673a = hgrant2_p & v1446737 | !hgrant2_p & v1446739;
assign v1284cc7 = hgrant1_p & v140583c | !hgrant1_p & v1284cc6;
assign v12161d9 = hmaster2_p & v12161d8 | !hmaster2_p & !v845542;
assign v134cede = hmaster0_p & v134d4a0 | !hmaster0_p & v845542;
assign v12ad53c = hmaster1_p & v12ad53b | !hmaster1_p & !v12ad525;
assign v1445b79 = hlock0 & v1445b78 | !hlock0 & v1445b77;
assign d308e1 = hmastlock_p & d308e0 | !hmastlock_p & v845542;
assign v1668d94 = hmaster1_p & v1668d8f | !hmaster1_p & v1668d93;
assign v12ad5ee = hmaster1_p & v12ad5ed | !hmaster1_p & v12ad5e1;
assign v140590f = hbusreq2_p & v140590c | !hbusreq2_p & v140590e;
assign v12ad5b2 = hgrant5_p & v12ad4d1 | !hgrant5_p & v12ad5b1;
assign d302d7 = hbusreq5_p & d308f4 | !hbusreq5_p & !d3068c;
assign v12ad623 = hgrant2_p & v12ad5fa | !hgrant2_p & !v12ad61f;
assign v16a13e4 = hbusreq0 & v16a2078 | !hbusreq0 & v16a13e3;
assign d30156 = hgrant5_p & v84555a | !hgrant5_p & d30119;
assign v1405b4a = hgrant0_p & v1405a86 | !hgrant0_p & v1405b49;
assign d2fbe2 = hgrant5_p & d2fbdc | !hgrant5_p & d2fbe1;
assign hmaster2 = !v114a3bf;
assign d3020d = hgrant5_p & d301c9 | !hgrant5_p & d3020b;
assign v134ced9 = hbusreq2 & v134ced8 | !hbusreq2 & v134d3ce;
assign f2f236 = hgrant5_p & v845542 | !hgrant5_p & !f2f235;
assign v12ad13d = hgrant2_p & v845542 | !hgrant2_p & v12ad13c;
assign v16a1e2e = hgrant2_p & v16a1dec | !hgrant2_p & v16a1e2d;
assign v121679d = hbusreq2_p & v121679a | !hbusreq2_p & v121679c;
assign v14457cd = hlock2 & v1445786 | !hlock2 & v14457c7;
assign d306c3 = hbusreq5 & d306bb | !hbusreq5 & d306c2;
assign v1516100 = hmaster2_p & v845542 | !hmaster2_p & v15160ff;
assign v1214c9b = hmaster0_p & v845542 | !hmaster0_p & v1215370;
assign v14461cf = hmaster1_p & v1446092 | !hmaster1_p & v14460b6;
assign v10d4019 = hbusreq1_p & v10d3fd5 | !hbusreq1_p & !v10d3fd4;
assign v1215c1d = hgrant5_p & v1215be7 | !hgrant5_p & v1215c1b;
assign v1515815 = hbusreq2_p & v1515814 | !hbusreq2_p & !v845542;
assign v15534ff = hmaster1_p & v1553385 | !hmaster1_p & v15534fe;
assign v144605a = hgrant1_p & v1446057 | !hgrant1_p & v1446059;
assign v16693a4 = hlock3_p & v16693a3 | !hlock3_p & !v845542;
assign d2fcfb = hmaster2_p & v1668c2d | !hmaster2_p & !d2fcaf;
assign v134ced0 = hgrant3_p & v134cec2 | !hgrant3_p & v134cecf;
assign v12ad5da = hgrant4_p & v12ad5d8 | !hgrant4_p & !v12ad5d9;
assign v1553227 = hbusreq1_p & v1553226 | !hbusreq1_p & v845542;
assign d2fbcf = hlock0_p & v845542 | !hlock0_p & !d30645;
assign v16a1ac5 = hmaster1_p & v16a1ac4 | !hmaster1_p & !v16a2672;
assign v1446120 = hlock2 & v144611c | !hlock2 & v144611f;
assign v12162b2 = hmaster0_p & f2f2a8 | !hmaster0_p & v1216035;
assign v1445f37 = hbusreq2_p & v1445f28 | !hbusreq2_p & v1445f36;
assign v1215c4d = hlock2_p & v1215c4c | !hlock2_p & v121657d;
assign v134d465 = hlock5 & v134d276 | !hlock5 & v134d464;
assign v16a193d = hbusreq4 & v16a1bb9 | !hbusreq4 & !v845542;
assign v1405aa7 = hmaster2_p & v845542 | !hmaster2_p & !v1405aa5;
assign bf1fa1 = hmaster2_p & bf1f9b | !hmaster2_p & bf1fa0;
assign v1446617 = hbusreq5_p & v1446616 | !hbusreq5_p & v1446611;
assign v14463ea = hbusreq5_p & v14463e9 | !hbusreq5_p & v14463bc;
assign v16a1957 = hgrant5_p & v845542 | !hgrant5_p & v16a1956;
assign v12ad56d = hlock2_p & v12ad56a | !hlock2_p & v12ad56c;
assign v12afa11 = decide_p & v12afa10 | !decide_p & v12afe76;
assign v16a1e63 = hbusreq5_p & v845568 | !hbusreq5_p & v16a1e62;
assign v14460f4 = hbusreq2 & v14460ee | !hbusreq2 & v14460f3;
assign v121504f = hgrant4_p & v845542 | !hgrant4_p & !v121504e;
assign d301ce = hbusreq1 & v845580 | !hbusreq1 & !v845542;
assign v1214d0e = hmaster0_p & v1214cef | !hmaster0_p & v1214d0d;
assign v1405b06 = hgrant1_p & v1405a92 | !hgrant1_p & v1405b05;
assign v15161fc = hgrant2_p & v15161fb | !hgrant2_p & !v845542;
assign v1445a34 = hgrant2_p & v144598f | !hgrant2_p & v1445a33;
assign v1445b83 = hlock2 & v1445b7f | !hlock2 & v1445b82;
assign v144600c = hgrant5_p & v1446467 | !hgrant5_p & v144647a;
assign d302e5 = hmaster1_p & v845542 | !hmaster1_p & d302e4;
assign v1445a47 = hbusreq2_p & v1445a34 | !hbusreq2_p & v1445a46;
assign v1215390 = hmastlock_p & v121538f | !hmastlock_p & v845542;
assign v16a1951 = hbusreq0 & v16a207a | !hbusreq0 & v16a1950;
assign v1405b0b = hgrant2_p & v1405ad1 | !hgrant2_p & v1405b0a;
assign v134d456 = hbusreq2 & v134d454 | !hbusreq2 & v134d455;
assign v1214bbb = hbusreq2_p & v1214bba | !hbusreq2_p & v1214bb9;
assign v134cdcb = hready_p & v134d3be | !hready_p & v134cdca;
assign v1214cf4 = hbusreq1_p & v1214cbb | !hbusreq1_p & v1214cf3;
assign v16a1a86 = hmaster1_p & v16a1a85 | !hmaster1_p & v16a1968;
assign v1446058 = hbusreq1 & v14465f0 | !hbusreq1 & v144669a;
assign v1405b2a = hmaster1_p & v1405b16 | !hmaster1_p & v1405b29;
assign v134ce96 = hbusreq3 & v134d240 | !hbusreq3 & v134ce95;
assign d3078b = hburst0 & d30789 | !hburst0 & d3078a;
assign v1515742 = hbusreq1 & v1515741 | !hbusreq1 & a65396;
assign v134d3c9 = hlock2 & v134d3c7 | !hlock2 & v134d3c8;
assign v1215334 = hmaster1_p & v121532a | !hmaster1_p & !v121507b;
assign v1214c23 = hbusreq2_p & v1214c22 | !hbusreq2_p & v1214c21;
assign d301fc = hgrant5_p & d301c6 | !hgrant5_p & d301fa;
assign v1216794 = hbusreq2_p & v1216791 | !hbusreq2_p & v1216793;
assign v12153b0 = hmaster2_p & v1215392 | !hmaster2_p & v1215399;
assign v14463fc = hlock2 & v14463f9 | !hlock2 & v14463fb;
assign d2fc58 = hgrant5_p & v84554a | !hgrant5_p & d2fc57;
assign f2f407 = hmaster1_p & f2f3f3 | !hmaster1_p & !f2f330;
assign v12af58d = hbusreq1_p & v12afe4e | !hbusreq1_p & v12afe45;
assign v1446000 = hmaster1_p & v1445feb | !hmaster1_p & v1445ffc;
assign v16a1dff = hmaster1_p & v16a1deb | !hmaster1_p & v16a1f96;
assign v12164c3 = hmaster1_p & v1216afb | !hmaster1_p & v1216af8;
assign decide = !v121482e;
assign v16a1cfb = hbusreq2_p & v16a1bea | !hbusreq2_p & v16a1cfa;
assign v1214fbc = hmaster2_p & v845542 | !hmaster2_p & v1214fbb;
assign v1445e85 = hbusreq0 & v1445e78 | !hbusreq0 & v1445e84;
assign v1445dcc = stateG10_5_p & v1445d8a | !stateG10_5_p & !v1445dcb;
assign v1446056 = hbusreq1 & v14465e7 | !hbusreq1 & v144641e;
assign v10d4006 = hmaster1_p & v10d3ff1 | !hmaster1_p & v10d3ffb;
assign f2f449 = hbusreq0 & f2f446 | !hbusreq0 & f2f448;
assign d30849 = hmaster1_p & d30848 | !hmaster1_p & !d30706;
assign v121653f = hlock1_p & v121653e | !hlock1_p & v845547;
assign v1515673 = hburst1 & v151566f | !hburst1 & v1515672;
assign v1446731 = hmaster0_p & v144664a | !hmaster0_p & v1446663;
assign v1215098 = hgrant1_p & v1215034 | !hgrant1_p & v1215097;
assign v13895a2 = hmaster0_p & v13895a1 | !hmaster0_p & v845542;
assign d2ff00 = hbusreq2_p & d2feff | !hbusreq2_p & d2fefa;
assign v1284d5d = hmaster0_p & v1284d23 | !hmaster0_p & v1284d0e;
assign v1214bbd = hmaster0_p & v12153b1 | !hmaster0_p & v1215396;
assign a658c8 = hburst1 & v845542 | !hburst1 & !v10d3fde;
assign v1445f34 = hbusreq2_p & v1445f28 | !hbusreq2_p & v1445f29;
assign v144585b = hlock2 & v1445857 | !hlock2 & v144585a;
assign v1405b5e = hmaster1_p & v1405b5d | !hmaster1_p & v1405b29;
assign a658d2 = hburst1 & v10d3fd6 | !hburst1 & v845542;
assign v1446232 = hbusreq0 & v144622e | !hbusreq0 & v1446214;
assign f2f235 = hmaster2_p & f2f22a | !hmaster2_p & f2f234;
assign v1216a8f = hbusreq5_p & v1216a8e | !hbusreq5_p & v845542;
assign v15530ed = hbusreq2 & v15530ec | !hbusreq2 & v155341e;
assign v1216a97 = hbusreq0_p & v16a1bc6 | !hbusreq0_p & v845570;
assign v12164c1 = hmaster0_p & v1216afb | !hmaster0_p & v1216ab3;
assign v1214bfd = hbusreq2_p & v1214bfc | !hbusreq2_p & v1214bfb;
assign v14458f1 = hlock4 & v14458d7 | !hlock4 & v14458d6;
assign v138944a = hmaster1_p & v845542 | !hmaster1_p & v1389449;
assign v16a1e0d = hbusreq2 & v16a1e0b | !hbusreq2 & !v16a1e0c;
assign v14058a9 = hgrant1_p & v1405849 | !hgrant1_p & v14058a8;
assign v121602a = hmaster0_p & v121601e | !hmaster0_p & v1216029;
assign v1214cf5 = hgrant1_p & v1214cf2 | !hgrant1_p & v1214cf4;
assign v134d368 = hmaster2_p & v134d367 | !hmaster2_p & v845542;
assign d3082d = hlock5_p & d3082b | !hlock5_p & d3082c;
assign v1445db4 = hbusreq2_p & v1445da5 | !hbusreq2_p & v1445db3;
assign v1445808 = hmaster0_p & v1445802 | !hmaster0_p & v1445eb0;
assign v1515736 = hbusreq5_p & v1515734 | !hbusreq5_p & v1515735;
assign d30697 = hbusreq2_p & d30636 | !hbusreq2_p & d30696;
assign d8076c = hgrant4_p & v845542 | !hgrant4_p & d8076b;
assign v16a132c = hmaster2_p & v16a1326 | !hmaster2_p & v845542;
assign d302e4 = hmaster0_p & d302e0 | !hmaster0_p & d302e3;
assign v12ad53e = hmaster1_p & v12ad53d | !hmaster1_p & !v12ad525;
assign v1214ccc = hgrant5_p & v1214cc2 | !hgrant5_p & v1214ccb;
assign v16a1e51 = hgrant2_p & v16a1dff | !hgrant2_p & v16a1e50;
assign v16a1cc6 = hbusreq5 & v16a1cba | !hbusreq5 & v16a1cc5;
assign v121679b = hmaster0_p & v12166f3 | !hmaster0_p & v12164e3;
assign v1215391 = hready & v1215390 | !hready & !v845542;
assign v12ad5c1 = hgrant0_p & a6537d | !hgrant0_p & !v12ad4d4;
assign v1284d08 = hmaster1_p & v1284d07 | !hmaster1_p & !v1445bb7;
assign a653b8 = hgrant1_p & a6539b | !hgrant1_p & !a65387;
assign v12ad5fa = hmaster1_p & v12ad5f9 | !hmaster1_p & v845542;
assign v12acfb7 = hbusreq5_p & v12ad523 | !hbusreq5_p & v12acfb6;
assign v14460d7 = hbusreq2_p & v14460d1 | !hbusreq2_p & v14460d6;
assign v1215ffc = hbusreq5_p & v1215ff4 | !hbusreq5_p & v1215ffb;
assign d30726 = hmaster2_p & d30723 | !hmaster2_p & d30725;
assign v1214fc8 = hbusreq2_p & v1214fc1 | !hbusreq2_p & v1214fc7;
assign v1668cff = hmaster2_p & v1668cdd | !hmaster2_p & !v1668cdf;
assign v1553509 = hlock5 & v155341e | !hlock5 & v15534f8;
assign v134d505 = hlock0_p & v134d273 | !hlock0_p & v134d504;
assign v1215d0a = hbusreq2 & v1215d07 | !hbusreq2 & v1215d09;
assign d302e9 = hmaster0_p & d302e7 | !hmaster0_p & d302e8;
assign v1216541 = hgrant1_p & v1216540 | !hgrant1_p & v121652d;
assign f2f3c5 = hgrant5_p & f2f3c1 | !hgrant5_p & f2f375;
assign v1516104 = hbusreq2_p & v1516103 | !hbusreq2_p & v845542;
assign v1405b1f = hmaster2_p & v1405b1e | !hmaster2_p & !v1405b1b;
assign v1445e58 = hlock1 & v1445e55 | !hlock1 & v1445e57;
assign v1214df3 = hbusreq1_p & v1214df2 | !hbusreq1_p & v845547;
assign v1215cac = hbusreq5_p & v1215ca9 | !hbusreq5_p & !v1215cab;
assign v144622a = hmaster2_p & v14463f2 | !hmaster2_p & v14463db;
assign v1445f48 = hmaster1_p & v1445f47 | !hmaster1_p & v1445da4;
assign bf1f74 = decide_p & bf1f73 | !decide_p & v845570;
assign v1214d81 = hmaster0_p & v1214c96 | !hmaster0_p & v1214c88;
assign v1668cf5 = hbusreq2_p & v1668cf2 | !hbusreq2_p & v1668ceb;
assign v16a1af3 = hgrant3_p & v16a1ad7 | !hgrant3_p & v16a1af2;
assign v12162eb = hbusreq1 & v1216aad | !hbusreq1 & v1216aea;
assign v1445dd2 = hmaster1_p & v144639c | !hmaster1_p & v1445dd1;
assign v12166f1 = hgrant2_p & v12166c2 | !hgrant2_p & v12166f0;
assign d30863 = hbusreq1_p & d3071a | !hbusreq1_p & d30688;
assign v1553421 = hlock3 & v155341e | !hlock3 & v1553420;
assign a6591f = hbusreq2_p & a6591c | !hbusreq2_p & a6591e;
assign v1216060 = hmaster0_p & v121604c | !hmaster0_p & v121605f;
assign f2f43d = hbusreq2_p & f2f41a | !hbusreq2_p & f2f43c;
assign v1215c1b = hmaster2_p & v1216538 | !hmaster2_p & v1215c1a;
assign v1446039 = hmaster1_p & v14465aa | !hmaster1_p & v1445fde;
assign v1446677 = hbusreq1 & v14465c4 | !hbusreq1 & v14465c5;
assign v121578f = hmaster2_p & v1215b92 | !hmaster2_p & v845542;
assign d301c5 = hbusreq1_p & v845542 | !hbusreq1_p & a65861;
assign v1515607 = hgrant3_p & v15155f0 | !hgrant3_p & !v1515606;
assign v1445be0 = hbusreq3_p & v1445ba9 | !hbusreq3_p & v1445bdf;
assign v1446291 = hmaster1_p & v1446405 | !hmaster1_p & v1446290;
assign v1668c3e = hmaster1_p & v1668c3d | !hmaster1_p & v845570;
assign a653c8 = locked_p & a658d3 | !locked_p & v10d3fd8;
assign v14463da = hbusreq1 & v14463d9 | !hbusreq1 & v14463a1;
assign v1284cfa = hgrant1_p & v140584b | !hgrant1_p & v1284cf9;
assign v1446173 = hmaster1_p & v1446172 | !hmaster1_p & v1445fef;
assign v121623a = hbusreq2_p & v1216239 | !hbusreq2_p & v121622e;
assign v1668c7c = hbusreq0 & v1668c6f | !hbusreq0 & v1668c7b;
assign v1215c72 = hmaster0_p & v1215c56 | !hmaster0_p & v1215c71;
assign v1446436 = hmaster0_p & v1446419 | !hmaster0_p & v1446435;
assign v12aead6 = hbusreq3_p & v12aef0b | !hbusreq3_p & v12aead5;
assign v1405b47 = locked_p & v1405aa1 | !locked_p & v1405a86;
assign v1446156 = hbusreq2_p & v1446152 | !hbusreq2_p & v1446155;
assign v1216104 = hbusreq5_p & v1216102 | !hbusreq5_p & !v1216103;
assign v1446246 = hbusreq3 & v1446229 | !hbusreq3 & v1446245;
assign v1553106 = hready_p & v1553427 | !hready_p & v1553105;
assign v14461ce = hmaster1_p & v144618d | !hmaster1_p & v1445ffc;
assign f2f2a3 = hmaster1_p & f2f297 | !hmaster1_p & f2f2a2;
assign v15157ea = hgrant5_p & v1668dc4 | !hgrant5_p & !v1515751;
assign v12acfcb = hmaster0_p & v12acfc4 | !hmaster0_p & v12ad67b;
assign d2fc00 = hgrant2_p & v84554a | !hgrant2_p & d2fbfe;
assign v1446700 = hbusreq2_p & v14466fd | !hbusreq2_p & v14466ff;
assign v14463b9 = hbusreq4_p & v144639c | !hbusreq4_p & v144639e;
assign v1445eb3 = hmaster2_p & v144639c | !hmaster2_p & v1445df2;
assign v1214ffa = hmaster2_p & v1214ff0 | !hmaster2_p & !v12153b7;
assign v16a1ac7 = hbusreq2 & v16a1ac6 | !hbusreq2 & v16a267b;
assign v138a3d3 = hgrant5_p & v845570 | !hgrant5_p & !v138a3d2;
assign v144634c = hbusreq2 & v144634a | !hbusreq2 & v144634b;
assign v1216a92 = hmaster0_p & v1216a8f | !hmaster0_p & v1216a91;
assign d30624 = hlock2_p & d30623 | !hlock2_p & d3061f;
assign a65693 = hmaster1_p & a658f1 | !hmaster1_p & a658e5;
assign v1215074 = hbusreq2_p & v1215073 | !hbusreq2_p & v1215070;
assign v16a1a27 = hbusreq2_p & v16a188a | !hbusreq2_p & v16a1a26;
assign v16a1bd5 = hbusreq1_p & v16a1bd4 | !hbusreq1_p & v16a206e;
assign f2f4a8 = hlock1_p & f2f4a7 | !hlock1_p & !v845542;
assign v1668cbb = hburst1 & v1668cba | !hburst1 & v845542;
assign v1215073 = hgrant2_p & v1215063 | !hgrant2_p & v1215072;
assign v1214ee6 = hgrant5_p & v845547 | !hgrant5_p & v121655a;
assign v1445ab9 = hmaster1_p & v1445ab8 | !hmaster1_p & v144589f;
assign v1668d1d = hmaster2_p & v1668d1c | !hmaster2_p & a6586b;
assign v12afe3f = decide_p & v12afe3e | !decide_p & v845542;
assign v12150f1 = hmaster1_p & v12153ee | !hmaster1_p & v12150ef;
assign v1215cc7 = hbusreq0 & v1215cc0 | !hbusreq0 & v1215cc6;
assign v1552d74 = decide_p & v155342e | !decide_p & v155321a;
assign v14460b5 = hlock0 & v14460b4 | !hlock0 & v14460b3;
assign v15157b9 = locked_p & v15157b8 | !locked_p & !v845542;
assign v1284cde = hgrant5_p & v140584c | !hgrant5_p & v1284cdd;
assign d2fc51 = hlock0_p & v845542 | !hlock0_p & d2fc50;
assign f2f44f = hgrant5_p & v84554c | !hgrant5_p & f2f431;
assign v15157e0 = hbusreq5_p & v15157de | !hbusreq5_p & !v15157df;
assign d3073b = stateG2_p & v845542 | !stateG2_p & d306ed;
assign v1215c54 = hgrant5_p & v845542 | !hgrant5_p & v1215bf2;
assign v12af73f = hbusreq5_p & v845542 | !hbusreq5_p & d30690;
assign v144537d = hmaster1_p & v1445a43 | !hmaster1_p & v1445a82;
assign v10d3fd2 = stateA1_p & v84557e | !stateA1_p & !v88d3e4;
assign d306dd = hbusreq1_p & d306dc | !hbusreq1_p & v845542;
assign v1553420 = hbusreq2 & v155341b | !hbusreq2 & v155341f;
assign v138a03a = decide_p & v138a039 | !decide_p & v138a406;
assign v140590b = hmaster0_p & v14058db | !hmaster0_p & v1405841;
assign v12aec0a = hmaster1_p & v12afe47 | !hmaster1_p & v12aec09;
assign v12ad58e = hmaster1_p & v12ad57b | !hmaster1_p & v12ad54f;
assign v12153d2 = hlock4_p & v12153d0 | !hlock4_p & v12153d1;
assign d2fc85 = hlock2_p & v845542 | !hlock2_p & d2fc84;
assign v12ad61b = hgrant5_p & v845542 | !hgrant5_p & !v12ad5e8;
assign v1215c13 = hbusreq1 & v121601f | !hbusreq1 & v845542;
assign v14453f3 = hmaster1_p & v14453f2 | !hmaster1_p & v1445bb7;
assign v10d4285 = hgrant1_p & v10d3fd5 | !hgrant1_p & v10d4284;
assign v121602f = hmaster0_p & v121602e | !hmaster0_p & v845542;
assign a65ae8 = hgrant5_p & v845542 | !hgrant5_p & a65ae7;
assign d307a2 = hgrant5_p & d306d1 | !hgrant5_p & d307a1;
assign v14461d8 = hgrant2_p & v14461d7 | !hgrant2_p & v14461cf;
assign d2fd19 = decide_p & d2fd18 | !decide_p & v845570;
assign v1214f55 = hmaster1_p & v1214f54 | !hmaster1_p & v1215d79;
assign v121501b = hmaster1_p & v121501a | !hmaster1_p & v12153bf;
assign v1669593 = hgrant3_p & v16693b2 | !hgrant3_p & !v1669592;
assign v134d1da = stateG3_2_p & v845542 | !stateG3_2_p & v134d1d9;
assign v1445801 = hbusreq0 & v1445ec6 | !hbusreq0 & v1445eb6;
assign v10d3fe8 = hmaster2_p & v10d3fe5 | !hmaster2_p & v10d3fe7;
assign v16a1c96 = hbusreq1_p & v16a1c95 | !hbusreq1_p & v845542;
assign v12acfbd = hmaster1_p & v12acfbc | !hmaster1_p & !v12ad525;
assign v1215dc2 = hready_p & v845542 | !hready_p & v1215dc1;
assign v15533a7 = hgrant5_p & v845542 | !hgrant5_p & v15533a6;
assign v11e5976 = hbusreq4_p & v11e5944 | !hbusreq4_p & v11e5975;
assign d2fb18 = hmaster0_p & d30159 | !hmaster0_p & d30137;
assign v138936c = hmaster2_p & v15155e7 | !hmaster2_p & v845542;
assign v1668d32 = hgrant5_p & v1668d2b | !hgrant5_p & v1668d30;
assign d30852 = hmaster2_p & d3084e | !hmaster2_p & !v845542;
assign f2e883 = hready_p & f2e73c | !hready_p & f2e882;
assign v134d3b4 = hmaster1_p & v134d369 | !hmaster1_p & v134d3b3;
assign v1445a74 = hmaster1_p & v144598e | !hmaster1_p & v144591b;
assign v1445869 = hready_p & v1445e52 | !hready_p & v1445868;
assign v12ad62f = hready_p & v12ad627 | !hready_p & !v12ad62e;
assign v1215c0e = hmaster2_p & v121652e | !hmaster2_p & v1215c0d;
assign d2f990 = hbusreq5_p & d2f98f | !hbusreq5_p & d2f98e;
assign v14465e9 = hbusreq1 & v14465e7 | !hbusreq1 & v14465e8;
assign v1216597 = hmaster2_p & v845542 | !hmaster2_p & v1216596;
assign v12153c0 = hmaster1_p & v12153b6 | !hmaster1_p & v12153bf;
assign v14459f3 = hbusreq1 & v14459f2 | !hbusreq1 & v14459b7;
assign v14058a0 = hgrant5_p & v140589f | !hgrant5_p & v140589d;
assign v134d4a0 = hlock0 & v134d49f | !hlock0 & v134d3aa;
assign d3094e = hburst0 & a658a5 | !hburst0 & d3094d;
assign a658b3 = hburst1 & a658b2 | !hburst1 & v845542;
assign v16a13ba = hmaster1_p & v16a13a8 | !hmaster1_p & v16a2672;
assign v134d467 = decide_p & v134d3ce | !decide_p & v134d466;
assign v16a1cd1 = hmaster0_p & v16a1ccc | !hmaster0_p & v16a1cd0;
assign v15156d5 = hbusreq1_p & a658bd | !hbusreq1_p & a65469;
assign v10d42b2 = hgrant1_p & v10d3fd4 | !hgrant1_p & v10d42b1;
assign v12ad661 = hbusreq0 & v845542 | !hbusreq0 & !v12af73f;
assign v14459be = hbusreq4 & v14459bc | !hbusreq4 & v14459bd;
assign v1214c55 = hbusreq5_p & v1214c53 | !hbusreq5_p & v1214c54;
assign v10d4291 = hlock0_p & v10d428f | !hlock0_p & v10d4290;
assign v1405856 = hmaster2_p & v140583c | !hmaster2_p & v14463b1;
assign v1446460 = hmaster0_p & v845542 | !hmaster0_p & v1446399;
assign v1405928 = hlock0_p & v140588e | !hlock0_p & v1405927;
assign v1405afd = hmaster2_p & v845542 | !hmaster2_p & !v1405afc;
assign v1515841 = hbusreq2 & v1515840 | !hbusreq2 & v1516803;
assign v10d4265 = stateA1_p & v84557e | !stateA1_p & v10d4264;
assign v16a1bba = hgrant0_p & v845542 | !hgrant0_p & v16a1bb9;
assign v16a1378 = hbusreq2 & v16a1375 | !hbusreq2 & v16a1377;
assign v151582f = hbusreq5 & v1515825 | !hbusreq5 & v151582e;
assign v1214fc1 = hgrant2_p & v1215787 | !hgrant2_p & v1214fc0;
assign v1445e4f = hmaster1_p & v1445e4e | !hmaster1_p & v845542;
assign v121531c = hbusreq2_p & v1215317 | !hbusreq2_p & v121531b;
assign d30710 = hmaster1_p & d3070f | !hmaster1_p & v84554e;
assign v15168a7 = hlock2_p & v15168a6 | !hlock2_p & v845542;
assign v12adf62 = hmaster2_p & v845542 | !hmaster2_p & v12adf61;
assign v1215354 = hbusreq4_p & v121534b | !hbusreq4_p & v1215345;
assign v1445e4c = hgrant2_p & v1446461 | !hgrant2_p & v1445e4b;
assign v12147e7 = hgrant2_p & v845542 | !hgrant2_p & v12147e6;
assign d2fc69 = hmaster2_p & d2fc68 | !hmaster2_p & d306a7;
assign v1446686 = hlock3 & v1446676 | !hlock3 & v1446685;
assign v14465bf = hready & v144639e | !hready & v14465bb;
assign v10d42a1 = hmaster0_p & v10d429b | !hmaster0_p & !v10d42a0;
assign v1515743 = hbusreq1_p & v1515740 | !hbusreq1_p & !v1515742;
assign v1445b55 = hmaster2_p & v1446653 | !hmaster2_p & v1446410;
assign f2f413 = hbusreq5 & f2f403 | !hbusreq5 & f2f412;
assign v12ad556 = hmaster1_p & v12ad537 | !hmaster1_p & v12ad54f;
assign d30266 = hmaster1_p & d30265 | !hmaster1_p & v845570;
assign d2fcb3 = hbusreq5_p & d2fcb2 | !hbusreq5_p & !d2fcb1;
assign v155392f = stateG3_0_p & v845586 | !stateG3_0_p & !v845586;
assign d2feb5 = hmaster2_p & d2feb2 | !hmaster2_p & d2feb4;
assign v1389539 = hlock5_p & v1389538 | !hlock5_p & !v845542;
assign v16a1bcd = hgrant5_p & v845542 | !hgrant5_p & v16a1bcc;
assign v16a1d9d = hbusreq3 & v16a1d9c | !hbusreq3 & v16a2063;
assign f2f3e2 = decide_p & f2f3e1 | !decide_p & f2f23c;
assign v1668c19 = hmaster0_p & v1668c18 | !hmaster0_p & v845570;
assign v1215ff2 = hmaster2_p & v1215fea | !hmaster2_p & v1215ff1;
assign v1446465 = hmaster2_p & v1446464 | !hmaster2_p & v845542;
assign v15161cc = hmaster1_p & v15161cb | !hmaster1_p & v845570;
assign d2fec2 = hlock4_p & v845542 | !hlock4_p & !d30727;
assign v1215352 = hbusreq5_p & v1215350 | !hbusreq5_p & v1215351;
assign d301f6 = hgrant5_p & d301f1 | !hgrant5_p & d301f5;
assign v14461e2 = hmaster1_p & v1446081 | !hmaster1_p & v14460cf;
assign v15167c4 = hbusreq2 & v15167b9 | !hbusreq2 & v15167c3;
assign v1215ce0 = hbusreq3 & v1215cdf | !hbusreq3 & v845542;
assign d2fc72 = hbusreq2 & d2fc70 | !hbusreq2 & d2fc71;
assign v1446404 = hmaster2_p & v144639c | !hmaster2_p & v1446403;
assign v14461b1 = hmaster1_p & v1446081 | !hmaster1_p & v14460b6;
assign v14466ba = hbusreq2_p & v14466ab | !hbusreq2_p & v14466b9;
assign v151579f = hbusreq5_p & v151579d | !hbusreq5_p & !v151579e;
assign f2f41d = hgrant1_p & f2f281 | !hgrant1_p & !f2f346;
assign d30236 = hgrant2_p & v845542 | !hgrant2_p & d3022e;
assign v134d459 = hlock5 & v134d449 | !hlock5 & v134d458;
assign d30132 = hbusreq5_p & d30131 | !hbusreq5_p & d30130;
assign v138a48d = hbusreq5 & v138a487 | !hbusreq5 & v138a404;
assign v16a1a20 = hmaster1_p & v16a19df | !hmaster1_p & v16a2672;
assign v12152f0 = hbusreq2_p & v12152eb | !hbusreq2_p & !v12152ef;
assign v144632e = hgrant2_p & v1446328 | !hgrant2_p & v144632d;
assign v1446066 = hgrant5_p & v1445fd9 | !hgrant5_p & v1446065;
assign v1668c70 = hmaster2_p & v1668c6e | !hmaster2_p & !a658e0;
assign d308b0 = hbusreq2_p & d30884 | !hbusreq2_p & !d308af;
assign d306d7 = hbusreq1_p & d306d6 | !hbusreq1_p & v845542;
assign v1446114 = hbusreq3 & v1446112 | !hbusreq3 & v1446113;
assign v1405b10 = hmaster0_p & v1405abd | !hmaster0_p & v1405abc;
assign d306c4 = decide_p & d306c3 | !decide_p & v845570;
assign v16a1418 = hbusreq2_p & v16a1417 | !hbusreq2_p & v16a2062;
assign d2f988 = hlock4_p & d308e1 | !hlock4_p & !d3094f;
assign d3082b = hgrant5_p & d306d0 | !hgrant5_p & d307ee;
assign v1216520 = hlock2_p & v121651c | !hlock2_p & v121651f;
assign v845582 = stateG2_p & v845542 | !stateG2_p & !v845542;
assign v12ae1f5 = hgrant0_p & v12ae1f4 | !hgrant0_p & !v845542;
assign v14461c6 = hmaster1_p & v1446189 | !hmaster1_p & v14460b6;
assign v16a1439 = hmaster2_p & v16a1438 | !hmaster2_p & v16a206f;
assign d30916 = hmaster2_p & a66278 | !hmaster2_p & !d30727;
assign v1445e9c = hlock1 & v1445e8d | !hlock1 & v1445e9b;
assign d3071a = hlock1_p & v845542 | !hlock1_p & d30719;
assign v1445ba9 = hgrant3_p & v14462a5 | !hgrant3_p & v1445ba8;
assign v1446745 = hbusreq2 & v1446735 | !hbusreq2 & v1446744;
assign d308e6 = hmaster0_p & d308e5 | !hmaster0_p & v845542;
assign v12ad56e = hmaster0_p & v12ad565 | !hmaster0_p & v12ad536;
assign v1446699 = hgrant4_p & v1446698 | !hgrant4_p & v14465ef;
assign v14058ad = hgrant4_p & v140584b | !hgrant4_p & v14058ac;
assign d2fd42 = decide_p & d2fd41 | !decide_p & v845570;
assign v134ceb9 = hlock2_p & v134d26d | !hlock2_p & v134ceb8;
assign v12ad5f3 = hmaster0_p & v845542 | !hmaster0_p & v12ad508;
assign v14453bc = hbusreq2_p & v14453b3 | !hbusreq2_p & v14453bb;
assign v1445fce = hbusreq5_p & v1445fcb | !hbusreq5_p & v1445fcd;
assign v1215bae = hbusreq4_p & v1215bad | !hbusreq4_p & v845542;
assign v12af9cf = hgrant0_p & v845542 | !hgrant0_p & !v1405a7d;
assign v1553445 = decide_p & v155342e | !decide_p & v1553423;
assign v1405aef = hgrant5_p & v1405a93 | !hgrant5_p & v1405aee;
assign d307ac = locked_p & v88d3e4 | !locked_p & a65861;
assign a66285 = hgrant4_p & a66284 | !hgrant4_p & !v845542;
assign v16a1d8d = hmaster1_p & v16a1d8c | !hmaster1_p & !v16a2672;
assign v1445f87 = hbusreq1_p & v1445f86 | !hbusreq1_p & v144639e;
assign v16a1dda = hbusreq5 & v16a1dd3 | !hbusreq5 & v16a1dd9;
assign v121574f = hlock5_p & v121574d | !hlock5_p & v121574e;
assign v1215c9a = hmaster2_p & v1215c8c | !hmaster2_p & v1215c99;
assign f2f53c = hgrant2_p & v845542 | !hgrant2_p & f2f53b;
assign v16a1d7c = hmaster1_p & v16a1d7b | !hmaster1_p & v16a1d7a;
assign a662a0 = hgrant1_p & v845542 | !hgrant1_p & !v84557a;
assign v1515613 = hbusreq0_p & a65851 | !hbusreq0_p & v151560d;
assign v1216236 = hgrant5_p & v12160d5 | !hgrant5_p & v1216235;
assign v16a208f = hgrant5_p & v845542 | !hgrant5_p & v16a208e;
assign v1216aed = hbusreq4_p & v1216aeb | !hbusreq4_p & v1216aec;
assign v12166dc = hgrant0_p & v12166db | !hgrant0_p & !v845542;
assign v12162f2 = hmaster2_p & v1216ad6 | !hmaster2_p & v1216aeb;
assign v144581d = hmaster1_p & v14457d8 | !hmaster1_p & v1445e28;
assign v140593a = hgrant2_p & v1405938 | !hgrant2_p & v1405939;
assign v144547e = hlock0 & v144547d | !hlock0 & v1446678;
assign d807c0 = hbusreq3_p & d807b5 | !hbusreq3_p & d807bf;
assign a6586b = hlock0_p & a65851 | !hlock0_p & a6586a;
assign v16a19ab = hmaster2_p & v16a19aa | !hmaster2_p & !v845542;
assign v1446620 = hgrant1_p & v1446432 | !hgrant1_p & v144661f;
assign v14453a8 = hgrant2_p & v144537c | !hgrant2_p & v14453a7;
assign v1553414 = hbusreq5_p & v1553413 | !hbusreq5_p & v1553218;
assign v16a1be2 = hbusreq0 & v16a1be0 | !hbusreq0 & v16a1be1;
assign v12af224 = hmaster2_p & v12af221 | !hmaster2_p & v12af223;
assign a65414 = hgrant5_p & a6587e | !hgrant5_p & a65378;
assign v1552f5e = hlock0_p & v1553217 | !hlock0_p & v1552f5d;
assign v12ad588 = hmaster1_p & v12ad572 | !hmaster1_p & v12ad54f;
assign v1214f1a = hbusreq2 & v1214f19 | !hbusreq2 & v845542;
assign v14058ac = hgrant0_p & v14058ab | !hgrant0_p & v140584b;
assign v15155e8 = hmaster2_p & v845542 | !hmaster2_p & v15155e7;
assign v1215fe2 = hbusreq3 & v12164e7 | !hbusreq3 & v121678b;
assign v1445404 = hmaster2_p & v144646e | !hmaster2_p & v845542;
assign v10d4064 = hgrant5_p & v10d3fdc | !hgrant5_p & v10d4063;
assign v1216a9e = hmaster1_p & v1216a9d | !hmaster1_p & v1216a9b;
assign v1445358 = hbusreq2_p & v1445b35 | !hbusreq2_p & v1445357;
assign v1668cbe = hmaster2_p & a658ad | !hmaster2_p & v1668cbd;
assign f2f3b5 = hgrant2_p & f2f3b4 | !hgrant2_p & !f2f3aa;
assign v15168b5 = hbusreq2_p & v15168b4 | !hbusreq2_p & v845542;
assign f2f38b = hbusreq1 & v1668d84 | !hbusreq1 & v845542;
assign d306ef = stateA1_p & v1553934 | !stateA1_p & !v845542;
assign d30662 = hgrant1_p & v845542 | !hgrant1_p & d30661;
assign v14464a2 = hmaster1_p & v1446466 | !hmaster1_p & v14464a1;
assign v16a188c = hmaster1_p & v16a1846 | !hmaster1_p & !v16a1f96;
assign d30740 = hmastlock_p & d3073f | !hmastlock_p & v845542;
assign v151697d = hmaster2_p & v845542 | !hmaster2_p & v15168ad;
assign d300c2 = hbusreq4_p & d300c1 | !hbusreq4_p & v845542;
assign v1215359 = hbusreq0 & v1215345 | !hbusreq0 & v845542;
assign v1446178 = hmaster1_p & v1446177 | !hmaster1_p & v1445fef;
assign v16a1d76 = hbusreq3 & v16a1d74 | !hbusreq3 & v16a1d56;
assign v1214c44 = hlock2_p & v1214c43 | !hlock2_p & v121536c;
assign v14459ee = stateG10_5_p & v14459eb | !stateG10_5_p & v14459ed;
assign v1445f15 = hlock2 & v1445f11 | !hlock2 & v1445f14;
assign d2f981 = hmaster2_p & v845542 | !hmaster2_p & !d3068e;
assign v1445b06 = hmaster0_p & v1445a6b | !hmaster0_p & v1445909;
assign v1214d0c = hgrant5_p & v1214c3b | !hgrant5_p & v1214d0b;
assign f2f22d = hbusreq1 & a66295 | !hbusreq1 & !v1668c1c;
assign v134d511 = hbusreq0 & v134d50c | !hbusreq0 & v134d510;
assign v1446223 = hmaster0_p & v1446214 | !hmaster0_p & v14463be;
assign v1405ab5 = hmaster0_p & v1405ab0 | !hmaster0_p & v1405aa3;
assign v1214f5c = hbusreq2_p & v1214f5b | !hbusreq2_p & v12164e7;
assign v10d40d5 = hgrant2_p & v10d40d2 | !hgrant2_p & v10d40d4;
assign v1553502 = hbusreq2_p & v1553500 | !hbusreq2_p & v1553501;
assign v1215439 = hmaster2_p & v1215438 | !hmaster2_p & v12153d9;
assign v12ad4ea = hmaster0_p & v12ad4e8 | !hmaster0_p & v12ad4e9;
assign a662a3 = decide_p & a6629f | !decide_p & a662a2;
assign v1446560 = hmaster2_p & v144655c | !hmaster2_p & v144655f;
assign v121601d = hlock1_p & v845547 | !hlock1_p & !v845542;
assign v16a19a8 = hbusreq4_p & v16a19a7 | !hbusreq4_p & v845542;
assign f2f227 = hbusreq1_p & f2f226 | !hbusreq1_p & !v845542;
assign v16a1e67 = hbusreq2 & v16a1e61 | !hbusreq2 & v16a1e66;
assign v12af1c3 = decide_p & v12af1c2 | !decide_p & v845542;
assign v1552f56 = hbusreq1 & v1552f55 | !hbusreq1 & v1553217;
assign v144627b = hlock0 & v144627a | !hlock0 & v1446279;
assign v845558 = hbusreq4_p & v845542 | !hbusreq4_p & !v845542;
assign d305f2 = hgrant4_p & d305f1 | !hgrant4_p & d305ef;
assign v14463cd = hmaster0_p & v14463a8 | !hmaster0_p & v14463bf;
assign v138a349 = hmaster2_p & v1515675 | !hmaster2_p & v138a335;
assign a662ad = hgrant5_p & v845542 | !hgrant5_p & a662ac;
assign v14058c0 = hgrant0_p & v140583d | !hgrant0_p & !v140588e;
assign v1445baf = hgrant5_p & v14463a6 | !hgrant5_p & !v1445bae;
assign bf1f6a = hmaster2_p & bf1f67 | !hmaster2_p & bf1f69;
assign v151570f = hmaster2_p & v1515609 | !hmaster2_p & a65851;
assign v1215b89 = hmaster1_p & v1215b7f | !hmaster1_p & v1215b88;
assign v14465d4 = hgrant5_p & v14465ba | !hgrant5_p & v14465d3;
assign bf1f84 = hgrant5_p & bf1f52 | !hgrant5_p & bf1f83;
assign v144591d = hmaster1_p & v1445903 | !hmaster1_p & v144591b;
assign v1214ee0 = hgrant5_p & v1214ed9 | !hgrant5_p & v1214edf;
assign v121531a = hmaster1_p & v121501d | !hmaster1_p & v1215016;
assign v12ad0b5 = hmaster1_p & v845542 | !hmaster1_p & v12ad0b4;
assign v1445448 = hmaster1_p & v1445447 | !hmaster1_p & v1446236;
assign v12164e1 = hmaster0_p & v12164db | !hmaster0_p & v12164e0;
assign d2feca = hmaster1_p & d2fec9 | !hmaster1_p & d2fec6;
assign v12af9be = hbusreq4_p & v12afe44 | !hbusreq4_p & v12af9bd;
assign v121533e = hbusreq2 & v1215333 | !hbusreq2 & v121533d;
assign d30213 = hgrant5_p & d301c0 | !hgrant5_p & d30212;
assign v1445ff0 = hmaster1_p & v1446405 | !hmaster1_p & v1445fef;
assign v15155eb = hmaster1_p & v15155ea | !hmaster1_p & v845542;
assign v1445b36 = hmaster0_p & v1445902 | !hmaster0_p & v1445a38;
assign v151582b = hlock2_p & v151582a | !hlock2_p & !v1515702;
assign v16a2241 = hmaster1_p & v16a2240 | !hmaster1_p & !v16a2672;
assign v155343f = hgrant5_p & v845542 | !hgrant5_p & v155343e;
assign v10d40a9 = hmaster0_p & v10d3ffd | !hmaster0_p & v10d400b;
assign v1214f58 = hbusreq2 & v1214f57 | !hbusreq2 & v12164e7;
assign v121622c = hmaster0_p & v1216209 | !hmaster0_p & v121622b;
assign v12162bf = hmaster0_p & v121622b | !hmaster0_p & v1216209;
assign d30669 = hmaster2_p & d30659 | !hmaster2_p & d30668;
assign v12ad522 = hbusreq4_p & v12ad521 | !hbusreq4_p & !v1668c6d;
assign d3061e = hmaster0_p & d3061b | !hmaster0_p & d3060c;
assign v1215c5a = hmaster0_p & v1215c56 | !hmaster0_p & v1215c59;
assign v1214f6e = hmaster0_p & v12166f2 | !hmaster0_p & v1215d63;
assign v16a1d17 = hburst1 & v16a1d16 | !hburst1 & v845542;
assign v138a35c = hmaster1_p & v138a35b | !hmaster1_p & v138a341;
assign v1445a12 = hgrant0_p & v14459bb | !hgrant0_p & v1445a11;
assign v12ad54e = hbusreq0 & v12ad54d | !hbusreq0 & !v845542;
assign v1445a3d = hmaster2_p & v14459a0 | !hmaster2_p & v14459ec;
assign v1389f92 = hbusreq5_p & v1389f91 | !hbusreq5_p & v845542;
assign v1215091 = hmaster2_p & v121508d | !hmaster2_p & v1214ffe;
assign v12153ed = hmaster1_p & v12153d4 | !hmaster1_p & v12153ec;
assign v1214da9 = hmaster0_p & v1214d0d | !hmaster0_p & v1214cef;
assign v1215453 = hbusreq2_p & v1215452 | !hbusreq2_p & v121544e;
assign v1216199 = hgrant5_p & v845542 | !hgrant5_p & v1216157;
assign v14453ea = hbusreq2_p & v1446254 | !hbusreq2_p & v14453e2;
assign v1553381 = hgrant0_p & v845542 | !hgrant0_p & v1553217;
assign f2f29a = hbusreq1_p & f2f299 | !hbusreq1_p & v845542;
assign v144541f = hbusreq2_p & v144541e | !hbusreq2_p & v144541b;
assign v16a1e6e = hbusreq3 & v16a1e67 | !hbusreq3 & v16a1e6d;
assign f2e273 = hbusreq4_p & f2f4b0 | !hbusreq4_p & !v845542;
assign v1215fbf = hgrant2_p & v1215fbc | !hgrant2_p & v1215fbe;
assign v1445afe = hlock2 & v1445af2 | !hlock2 & v1445afc;
assign v16a1a91 = hbusreq3_p & v16a19cf | !hbusreq3_p & v16a1a90;
assign v134cdc7 = hbusreq3 & v134cdc6 | !hbusreq3 & v134d276;
assign v12ad524 = hbusreq0 & v12ad523 | !hbusreq0 & v12afdb1;
assign v16a1409 = decide_p & v16a13fd | !decide_p & v16a1408;
assign v1216204 = hbusreq1_p & v1216203 | !hbusreq1_p & v845547;
assign v138a3e5 = hmaster1_p & v138a3e4 | !hmaster1_p & v138a314;
assign v12ad4e4 = hlock0_p & v845570 | !hlock0_p & d2fbe5;
assign v1445f80 = hbusreq5 & v1445f62 | !hbusreq5 & v1445f7f;
assign v1215395 = hmaster2_p & v1215392 | !hmaster2_p & v1215394;
assign v15157d3 = hlock2_p & v1515787 | !hlock2_p & v15157d2;
assign d2fb69 = hlock0_p & v845542 | !hlock0_p & !v16693aa;
assign v121613a = hbusreq1 & v1216139 | !hbusreq1 & v845542;
assign v1216010 = hmaster1_p & v121600f | !hmaster1_p & v121600c;
assign d2fe88 = hbusreq5_p & d2fe86 | !hbusreq5_p & d2fe87;
assign v1446121 = hmaster0_p & v1446077 | !hmaster0_p & v1446404;
assign a653c5 = hbusreq4_p & a653c4 | !hbusreq4_p & v845542;
assign a658dc = hmastlock_p & a658db | !hmastlock_p & v845542;
assign v138a342 = hmaster1_p & v138a32d | !hmaster1_p & v138a341;
assign v1214ec7 = hready_p & v1214de3 | !hready_p & v1214ec6;
assign v138a31f = hlock3_p & v138a30d | !hlock3_p & v138a31e;
assign v1216574 = hbusreq0 & v1216564 | !hbusreq0 & v1216573;
assign v1446164 = hmaster1_p & v1446163 | !hmaster1_p & v1446073;
assign v1214c01 = hmaster1_p & v1214c00 | !hmaster1_p & v12153a9;
assign v16a1423 = hbusreq3 & v16a1420 | !hbusreq3 & v16a1422;
assign a6564c = hgrant1_p & a653c7 | !hgrant1_p & !a6564b;
assign v134d4c9 = hmastlock_p & v134d4c8 | !hmastlock_p & v845542;
assign v1215b76 = hbusreq4_p & v12160eb | !hbusreq4_p & v845542;
assign v1445f8f = hbusreq5_p & v1445f85 | !hbusreq5_p & v1445f8e;
assign v14058f5 = hmaster2_p & v14058f4 | !hmaster2_p & !v14058ee;
assign v1215370 = hbusreq0 & v1216a7f | !hbusreq0 & v845542;
assign d305d6 = hlock5_p & v845542 | !hlock5_p & v845570;
assign v16a1dd8 = hbusreq2 & v16a1dd6 | !hbusreq2 & v16a1dd7;
assign v1405b22 = hbusreq4_p & v845542 | !hbusreq4_p & v1405b18;
assign v1405ab4 = hbusreq2_p & v1405ab3 | !hbusreq2_p & v1405aaf;
assign bf1f69 = hgrant1_p & f2f227 | !hgrant1_p & bf1f68;
assign v1214c16 = hmaster1_p & v1214bfe | !hmaster1_p & v1214bcf;
assign v10d40ac = hmaster1_p & v10d40ab | !hmaster1_p & !v10d3fe9;
assign d30128 = hmaster0_p & v84555a | !hmaster0_p & d2fea9;
assign d2fae1 = hbusreq1_p & d300dd | !hbusreq1_p & d2fae0;
assign v14466a5 = hmaster2_p & v144669c | !hmaster2_p & v144662a;
assign v1552f66 = hgrant5_p & v845542 | !hgrant5_p & v1552f65;
assign v134d36f = hlock4 & v134d273 | !hlock4 & v134d36e;
assign v121510a = hbusreq3 & v12150f7 | !hbusreq3 & v1215109;
assign v144607a = hmaster0_p & v1446404 | !hmaster0_p & v1446079;
assign v1214d36 = hmaster1_p & v1214d35 | !hmaster1_p & v121536b;
assign v12afe53 = hlock0_p & v15168f4 | !hlock0_p & !v845542;
assign v10d427c = hmastlock_p & v10d427b | !hmastlock_p & v10d3fd3;
assign v16a1db9 = hbusreq5 & v16a1d56 | !hbusreq5 & v16a209f;
assign v1216321 = hbusreq5_p & v1216320 | !hbusreq5_p & v12162fe;
assign v121619e = hgrant2_p & v12160ea | !hgrant2_p & v121619d;
assign v1405936 = hgrant2_p & v140591c | !hgrant2_p & v1405935;
assign v14458a0 = hmaster1_p & v144639c | !hmaster1_p & v144589f;
assign v144616e = hmaster1_p & v144616d | !hmaster1_p & v1446073;
assign v121606c = hmaster0_p & v121604c | !hmaster0_p & v121606b;
assign v15157c7 = hgrant1_p & f2f281 | !hgrant1_p & v15157c6;
assign v12ad4c1 = hbusreq5_p & v12adf62 | !hbusreq5_p & v12ad4c0;
assign v144603f = hgrant5_p & v1446404 | !hgrant5_p & v144603e;
assign d307c1 = hgrant5_p & d307ad | !hgrant5_p & d307c0;
assign v1216256 = hgrant2_p & v1216202 | !hgrant2_p & v1216255;
assign f2f44e = hbusreq0 & f2f44b | !hbusreq0 & f2f44d;
assign v1446041 = hmaster2_p & v14465b3 | !hmaster2_p & v14465db;
assign v1216aa9 = hready & v1216aa8 | !hready & !v845542;
assign v121619d = hmaster1_p & v121618e | !hmaster1_p & v121619c;
assign a6590f = hbusreq2_p & a65909 | !hbusreq2_p & a6590e;
assign d3079e = hlock1_p & d3079d | !hlock1_p & d30790;
assign d2fae8 = hbusreq1_p & d300cc | !hbusreq1_p & d2fae7;
assign v1445fc2 = hbusreq2_p & v1445fbe | !hbusreq2_p & v1445fc1;
assign v16a1970 = hgrant1_p & v84554d | !hgrant1_p & v16a196f;
assign v144665a = hbusreq1 & v14465cb | !hbusreq1 & v14465cf;
assign v1216137 = hbusreq4_p & v1216552 | !hbusreq4_p & v1216136;
assign v144663b = hmaster0_p & v1446404 | !hmaster0_p & v144663a;
assign v1284cb2 = hmaster1_p & v1284cb1 | !hmaster1_p & v1284ca7;
assign v1214c34 = hbusreq5_p & v1214c32 | !hbusreq5_p & v1214c33;
assign v1446654 = hmaster2_p & v144639c | !hmaster2_p & v1446653;
assign v14465de = hbusreq5_p & v14465d4 | !hbusreq5_p & v14465dd;
assign v140584f = hmaster2_p & v140583d | !hmaster2_p & v1405844;
assign v1445be5 = hgrant2_p & v1445be3 | !hgrant2_p & v144632d;
assign v1446324 = hmaster1_p & v1446323 | !hmaster1_p & v14462ff;
assign v1445b93 = hmaster1_p & v1446323 | !hmaster1_p & v1445b8d;
assign d308db = hbusreq1_p & d308da | !hbusreq1_p & v845542;
assign v1516979 = hmaster0_p & v845542 | !hmaster0_p & v1668c28;
assign v1515729 = hgrant4_p & v1515715 | !hgrant4_p & v1515728;
assign v1216ad6 = hbusreq4_p & v1216ad5 | !hbusreq4_p & v845547;
assign v1284ce7 = hgrant2_p & v14058b6 | !hgrant2_p & v1284ce6;
assign v14459a0 = hgrant1_p & v14458d2 | !hgrant1_p & v144599a;
assign v1445aa2 = hgrant2_p & v1445a89 | !hgrant2_p & v1445aa1;
assign v1405b61 = hgrant2_p & v1405b5c | !hgrant2_p & v1405b60;
assign v1405b68 = jx1_p & v1405a84 | !jx1_p & v1405b67;
assign v138a321 = stateG3_2_p & v845562 | !stateG3_2_p & d3094a;
assign v1446414 = hbusreq5_p & v1446411 | !hbusreq5_p & v1446413;
assign v16a13c0 = hmaster1_p & v16a2669 | !hmaster1_p & !v16a2672;
assign v1214feb = hgrant1_p & v12153b4 | !hgrant1_p & v1214fea;
assign v10d42ba = hmaster1_p & v10d42b9 | !hmaster1_p & v10d407c;
assign v121678d = decide_p & v12164ce | !decide_p & v121678c;
assign v12150ed = hlock5_p & v12150ec | !hlock5_p & v12150c9;
assign v845548 = hbusreq0_p & v845542 | !hbusreq0_p & !v845542;
assign v8af912 = hburst0_p & v893df7 | !hburst0_p & v845542;
assign v86ab0d = hburst1_p & v845542 | !hburst1_p & v8dfa41;
assign a6537e = hgrant0_p & a6537d | !hgrant0_p & a6536d;
assign v10d40dd = hgrant3_p & v10d40af | !hgrant3_p & !v10d40dc;
assign v12162e1 = hready_p & v12162bc | !hready_p & v12162e0;
assign d2fb9f = hmaster1_p & d2fb7f | !hmaster1_p & d2fb9d;
assign v1214bf6 = hbusreq2 & v1214bdc | !hbusreq2 & v1214bf5;
assign v16a1cc5 = hbusreq3 & v16a1cbf | !hbusreq3 & v16a1cc4;
assign v134d46a = hready_p & v134d3e5 | !hready_p & v134d469;
assign v15534f0 = hmaster0_p & v845542 | !hmaster0_p & v15534ef;
assign v1284cea = hbusreq1_p & v1284c8f | !hbusreq1_p & v1284ce9;
assign v1405899 = stateA1_p & v845542 | !stateA1_p & v1405853;
assign f2f3af = hgrant2_p & f2f3ae | !hgrant2_p & f2f394;
assign v1389462 = hgrant2_p & v845542 | !hgrant2_p & !v1389461;
assign v1446482 = hlock0_p & v1446398 | !hlock0_p & v1446481;
assign v1216561 = hgrant1_p & v845542 | !hgrant1_p & v1216560;
assign v1216194 = hgrant5_p & v121618f | !hgrant5_p & v121612a;
assign v1216ab1 = hmaster2_p & v845542 | !hmaster2_p & !v1216ab0;
assign a65678 = hmaster0_p & a65670 | !hmaster0_p & a65677;
assign v1405a8f = hbusreq5_p & v1405a8d | !hbusreq5_p & !v1405a8e;
assign v12153a9 = hmaster0_p & v12153a2 | !hmaster0_p & v12153a8;
assign v1216176 = hgrant5_p & v121600e | !hgrant5_p & v1216175;
assign v144662c = hgrant5_p & v14465ea | !hgrant5_p & v144662b;
assign v134ce6d = hlock5 & v134d3b5 | !hlock5 & v134ce5d;
assign v16a1848 = hmaster1_p & v16a1842 | !hmaster1_p & v16a2672;
assign d305e9 = stateA1_p & v845542 | !stateA1_p & !v156645f;
assign v16a1ace = hbusreq2_p & v16a1f98 | !hbusreq2_p & v16a1acd;
assign v1515670 = busreq_p & v151566d | !busreq_p & !v845542;
assign d2fad4 = hgrant2_p & d2fad1 | !hgrant2_p & d2fad3;
assign v151564b = hburst1 & v1515648 | !hburst1 & v151564a;
assign f2f39a = hbusreq1_p & f2f399 | !hbusreq1_p & !v845542;
assign a65b18 = hgrant2_p & v845542 | !hgrant2_p & a65b17;
assign v15156c7 = hgrant1_p & v15156c6 | !hgrant1_p & v1668cc4;
assign v1214c8b = hgrant5_p & v16a2243 | !hgrant5_p & v1214c5d;
assign v1515656 = hbusreq1 & a658d4 | !hbusreq1 & !a658dc;
assign v1445859 = hgrant2_p & v1445835 | !hgrant2_p & v1445858;
assign v1552d6b = hbusreq5 & v1552d69 | !hbusreq5 & v1552d6a;
assign f2f454 = hmaster0_p & f2f44e | !hmaster0_p & f2f453;
assign d30290 = hgrant5_p & d3028f | !hgrant5_p & !d30275;
assign v14465c6 = hbusreq1 & v14465c2 | !hbusreq1 & v14465c5;
assign v11e5954 = hgrant4_p & v11e5953 | !hgrant4_p & !v845542;
assign v1214c00 = hmaster0_p & v12153ab | !hmaster0_p & v1214bb7;
assign a65b27 = decide_p & a65b26 | !decide_p & v845542;
assign v1216078 = hmaster0_p & v1216068 | !hmaster0_p & v121606b;
assign v15156b8 = hburst0 & f2f4ad | !hburst0 & v15156b7;
assign v134d282 = hlock1_p & v134d1dd | !hlock1_p & v845542;
assign d2fcae = hlock1_p & d2fcad | !hlock1_p & !v845542;
assign d2fc18 = hbusreq2 & d2fc15 | !hbusreq2 & d2fc17;
assign v12afdab = hlock0_p & d305ef | !hlock0_p & v845542;
assign d8076b = hgrant0_p & v845542 | !hgrant0_p & !d8076a;
assign d2fe9d = hbusreq1_p & v84555a | !hbusreq1_p & d2fe9c;
assign v16a2236 = stateG2_p & v845542 | !stateG2_p & !v16a2235;
assign v1668d4f = hbusreq1_p & v10d3fd8 | !hbusreq1_p & !a65861;
assign v12ad632 = hmaster1_p & v12ad631 | !hmaster1_p & v12ad4ff;
assign v1284ccc = hbusreq1_p & v1284ccb | !hbusreq1_p & !v140589a;
assign v140588c = hlock0_p & v140583d | !hlock0_p & v140583c;
assign f2f3c0 = hgrant5_p & f2f3bf | !hgrant5_p & !f2f35f;
assign v1215bc6 = hbusreq2_p & v1215bc5 | !hbusreq2_p & v1215bc4;
assign v16a1d21 = hbusreq2 & v16a1d1b | !hbusreq2 & v16a1d20;
assign d2f99a = hbusreq1_p & d2feb2 | !hbusreq1_p & d2f999;
assign v1214dd5 = hmaster1_p & v1214dd4 | !hmaster1_p & v845542;
assign v1214d79 = hgrant2_p & v1214d76 | !hgrant2_p & v1214d78;
assign v144549e = hlock3 & v144546f | !hlock3 & v144549d;
assign v1215ba9 = hmaster1_p & v1215ba8 | !hmaster1_p & v845542;
assign d3070d = hlock1_p & d3070c | !hlock1_p & v845542;
assign a65468 = hburst0 & v156645f | !hburst0 & a65467;
assign v1215d80 = hgrant5_p & v12164cf | !hgrant5_p & v12166c5;
assign v1214bdb = hlock2_p & v1214bd9 | !hlock2_p & v1214bda;
assign v11e5946 = hgrant1_p & v845542 | !hgrant1_p & v11e5945;
assign v1284d33 = hmaster1_p & v1284d32 | !hmaster1_p & v1284ca7;
assign v845555 = hbusreq3 & v845542 | !hbusreq3 & !v845542;
assign v14459e7 = hgrant1_p & v14459e5 | !hgrant1_p & v14459e6;
assign v14058f9 = hgrant4_p & v140583f | !hgrant4_p & !v14465b1;
assign v144591e = hbusreq2_p & v144591c | !hbusreq2_p & v144591d;
assign f2f2d8 = hbusreq1_p & f2f2d7 | !hbusreq1_p & !v845542;
assign a65b1a = decide_p & a65b19 | !decide_p & a662a2;
assign v138a30e = hlock5_p & v1515638 | !hlock5_p & !v845542;
assign v11e597e = hgrant2_p & bf1f59 | !hgrant2_p & v11e597d;
assign v1445bef = hgrant2_p & v1445bec | !hgrant2_p & v1445bee;
assign d2fc0f = hbusreq5_p & d2fc0e | !hbusreq5_p & d2fbf0;
assign v166959d = decide_p & v166959c | !decide_p & v845542;
assign v134cee2 = hlock3 & v134d276 | !hlock3 & v134cee1;
assign v134d229 = hbusreq5_p & v134d228 | !hbusreq5_p & v134d1e8;
assign f2f3ea = hbusreq2_p & f2f3e7 | !hbusreq2_p & f2f3e9;
assign v16a1ced = hgrant5_p & v845542 | !hgrant5_p & v16a1cec;
assign v1445e65 = hgrant4_p & v1445dea | !hgrant4_p & v1445e64;
assign v10d3fe1 = hbusreq1_p & v10d3fdb | !hbusreq1_p & v10d3fe0;
assign v13891a5 = hmaster1_p & v845542 | !hmaster1_p & v13891a4;
assign v1215ba0 = hlock4_p & v1216147 | !hlock4_p & !v845542;
assign v12ad4f8 = hmaster2_p & v10d3fd8 | !hmaster2_p & v12ad4f7;
assign v1214c3b = hmaster2_p & v1214c29 | !hmaster2_p & v1214c30;
assign v1445bfa = jx2_p & v1445be0 | !jx2_p & v1445bf9;
assign v1214d28 = hmaster1_p & v1214d27 | !hmaster1_p & !v1214d1e;
assign v121610c = hbusreq1 & v1216537 | !hbusreq1 & v845542;
assign v1516802 = hgrant2_p & v845552 | !hgrant2_p & !v845542;
assign d3028c = hbusreq2_p & d3028b | !hbusreq2_p & !d30286;
assign v1445e6d = hmaster2_p & v14465b3 | !hmaster2_p & v1445e6c;
assign v1216568 = hready & v1216a60 | !hready & v1216567;
assign d2fc6c = hbusreq0 & d2fc6b | !hbusreq0 & d306bc;
assign v12ad578 = hmaster1_p & v12ad577 | !hmaster1_p & !v12ad525;
assign v1216a5c = hburst1_p & v134d1d9 | !hburst1_p & v1216a5b;
assign d300f3 = hmaster2_p & d300f2 | !hmaster2_p & d300ed;
assign v14058f0 = hgrant5_p & v14058ed | !hgrant5_p & !v14058ef;
assign d30826 = hbusreq0 & d30823 | !hbusreq0 & d30825;
assign v1552d5b = hmaster2_p & v1553412 | !hmaster2_p & v845542;
assign v134cec7 = hbusreq2_p & v134d4b0 | !hbusreq2_p & v134d3b5;
assign v138a300 = hbusreq5_p & v138a2ff | !hbusreq5_p & v845542;
assign d30893 = hgrant5_p & d3084f | !hgrant5_p & !d30892;
assign d80766 = hready_p & d80738 | !hready_p & !d80765;
assign v151574c = hmaster2_p & v1515741 | !hmaster2_p & !v10d3ff3;
assign v1214c95 = hgrant5_p & v845542 | !hgrant5_p & v1214c77;
assign v121538b = hmaster0_p & v121537b | !hmaster0_p & v121538a;
assign d2fbca = hlock1_p & d2fb4d | !hlock1_p & v84554a;
assign v16a2086 = hmaster2_p & v16a2085 | !hmaster2_p & v16a2080;
assign d2fee1 = hbusreq3 & d2fed4 | !hbusreq3 & d2fee0;
assign v14459ac = hlock0_p & v14459aa | !hlock0_p & v14459ab;
assign a65699 = hbusreq2 & a65690 | !hbusreq2 & a65698;
assign v16a1444 = hgrant2_p & v845542 | !hgrant2_p & v16a1442;
assign v12153b9 = hmaster2_p & v1215bac | !hmaster2_p & v12153b7;
assign v1214e7f = hmaster1_p & v1214e5a | !hmaster1_p & v1214e73;
assign v1445870 = hlock1 & v144586f | !hlock1 & v144586d;
assign v14466ce = hmaster1_p & v14463c9 | !hmaster1_p & v14463c2;
assign v1446647 = hgrant5_p & v144643d | !hgrant5_p & v1446646;
assign v1216084 = hmaster1_p & v1216060 | !hmaster1_p & v1216082;
assign v1215cab = hgrant5_p & v845542 | !hgrant5_p & !v1215caa;
assign d2f9bc = hbusreq2_p & d2f9bb | !hbusreq2_p & d2f9aa;
assign v1214ec2 = hmaster0_p & v12164d4 | !hmaster0_p & v1215d63;
assign v1445fec = hmaster1_p & v1445feb | !hmaster1_p & v1445fde;
assign v1215717 = hgrant1_p & v121570e | !hgrant1_p & v1215716;
assign v134d231 = hbusreq2_p & v134d230 | !hbusreq2_p & v134d22f;
assign v134d50e = hgrant1_p & v845542 | !hgrant1_p & v134d507;
assign a6541b = hgrant5_p & v845558 | !hgrant5_p & !a6538a;
assign d3024d = hgrant5_p & v845542 | !hgrant5_p & d3020b;
assign v1215bdf = hmaster2_p & v1215ff8 | !hmaster2_p & v1215bdd;
assign v14058cc = hgrant5_p & v14058ca | !hgrant5_p & v14058cb;
assign v1516855 = hgrant3_p & v15167f1 | !hgrant3_p & !v1516854;
assign v1215d42 = hmaster0_p & v1215d2f | !hmaster0_p & v1215d41;
assign v1214c94 = hgrant2_p & v1214c44 | !hgrant2_p & v1214c93;
assign v14465ca = hgrant0_p & v144640c | !hgrant0_p & v14463a0;
assign v15161d2 = hmaster1_p & v15161d1 | !hmaster1_p & v845570;
assign v16a1ccc = hbusreq5_p & v16a1afb | !hbusreq5_p & v16a1ccb;
assign d30817 = hlock5_p & d30815 | !hlock5_p & d30816;
assign v12acfc2 = hmaster2_p & v12ad675 | !hmaster2_p & v12acfc1;
assign v138a33e = hmaster2_p & v1668c6e | !hmaster2_p & !v138a33d;
assign a65866 = hmaster2_p & a65852 | !hmaster2_p & a65864;
assign v134d390 = hgrant0_p & v134d38f | !hgrant0_p & v845542;
assign v1214eda = hmaster2_p & v121652e | !hmaster2_p & v1216541;
assign d2fef0 = hlock2_p & d2feee | !hlock2_p & d2feef;
assign v121605c = hbusreq0 & v1216056 | !hbusreq0 & v121605b;
assign v12152ff = hgrant2_p & v1215786 | !hgrant2_p & v12152fe;
assign v1216274 = hmaster1_p & v1216273 | !hmaster1_p & v1216041;
assign v1284cad = hmaster2_p & v140588d | !hmaster2_p & v144639e;
assign v10d4088 = decide_p & v10d405c | !decide_p & v10d4087;
assign v1214f66 = hgrant3_p & v1214ec7 | !hgrant3_p & v1214f65;
assign v14465ed = hbusreq4_p & v144639c | !hbusreq4_p & v14465ec;
assign v1284d57 = hmaster1_p & v1284ce3 | !hmaster1_p & !v1284cfd;
assign v1553153 = hlock2_p & v155314f | !hlock2_p & v1553152;
assign v12ad504 = hmaster1_p & v12ad503 | !hmaster1_p & v12ad4ff;
assign v12acfe8 = hmaster1_p & v12acfd0 | !hmaster1_p & v12ad54f;
assign d2fe89 = hlock4_p & d306df | !hlock4_p & v845570;
assign v134d1ed = hbusreq4_p & v134d1e8 | !hbusreq4_p & v134d1ec;
assign v144620f = hgrant5_p & v144620c | !hgrant5_p & !v144620e;
assign v1445e9b = hgrant4_p & v1445e02 | !hgrant4_p & v1445e9a;
assign v16a1945 = hbusreq4_p & v16a1944 | !hbusreq4_p & v845542;
assign v1445a95 = hlock5 & v1445a73 | !hlock5 & v1445a94;
assign v1668e0c = hready_p & v845542 | !hready_p & v1668e0b;
assign d2fd28 = hbusreq2_p & d2fd27 | !hbusreq2_p & d302e5;
assign a65af2 = hmaster1_p & a65ae6 | !hmaster1_p & a65af1;
assign v14466e2 = hmaster1_p & v14466cc | !hmaster1_p & v14463ef;
assign v16a1d6b = hgrant5_p & v845542 | !hgrant5_p & v16a1d6a;
assign v1389d58 = hmaster2_p & v1668c49 | !hmaster2_p & !v845542;
assign v12ad5af = hgrant4_p & v12ad5ad | !hgrant4_p & !v12ad5ae;
assign v1446263 = hbusreq5_p & v1446261 | !hbusreq5_p & v1446262;
assign v14466e3 = hmaster0_p & v14463c9 | !hmaster0_p & v14463f6;
assign v1515707 = hlock2_p & v1515706 | !hlock2_p & !v1515702;
assign v12ad028 = hbusreq5_p & v12ad60e | !hbusreq5_p & v12ad027;
assign d2fef7 = hbusreq5 & d2fee1 | !hbusreq5 & d2fef6;
assign d3027d = hbusreq5_p & d3027c | !hbusreq5_p & !d3027b;
assign bf1f6c = hgrant5_p & v845542 | !hgrant5_p & !bf1f6a;
assign v1446269 = hlock0 & v1446268 | !hlock0 & v14465ea;
assign v16a1e4d = hmaster1_p & v16a1e28 | !hmaster1_p & v16a1f96;
assign v1389fff = hmaster2_p & v15168f4 | !hmaster2_p & v845570;
assign v1214c7b = hbusreq0 & v1214c7a | !hbusreq0 & v845542;
assign v1214d01 = hmaster2_p & v1214d00 | !hmaster2_p & v845542;
assign v138a476 = decide_p & v138a475 | !decide_p & !v845542;
assign v1445ecf = hgrant2_p & v1445ec5 | !hgrant2_p & v1445ece;
assign v1445413 = hmaster2_p & v1445412 | !hmaster2_p & v14465b3;
assign v1446619 = hbusreq0_p & v144639c | !hbusreq0_p & v14465c1;
assign v1445ed4 = hmaster1_p & v14465b7 | !hmaster1_p & v1445ed3;
assign d2fc40 = hbusreq0 & d2fb9b | !hbusreq0 & d2fc33;
assign v1445dec = hbusreq4_p & v1446407 | !hbusreq4_p & v1446406;
assign a64715 = hbusreq3_p & a6470a | !hbusreq3_p & a64714;
assign v134d4e4 = decide_p & v134d309 | !decide_p & v134d4e3;
assign v1445a35 = hmaster2_p & v14458d2 | !hmaster2_p & v14459d3;
assign v1214d24 = hgrant2_p & v1214d16 | !hgrant2_p & v1214d1f;
assign v12162c4 = hmaster1_p & v121622b | !hmaster1_p & v1216224;
assign a656c2 = hgrant2_p & v845542 | !hgrant2_p & a656c1;
assign v16a131e = hmastlock_p & v16a131d | !hmastlock_p & !v845542;
assign v12153e7 = hlock0_p & v12153d7 | !hlock0_p & v845542;
assign v1215785 = hmaster0_p & v845542 | !hmaster0_p & v1215ba7;
assign v1214d2d = hgrant2_p & v1214d0a | !hgrant2_p & v1214d2c;
assign v12150d2 = hmaster1_p & v1215443 | !hmaster1_p & v12150d1;
assign d300b2 = hmaster0_p & d2fe81 | !hmaster0_p & d2fe7e;
assign v134d387 = hmaster2_p & v134d383 | !hmaster2_p & v134d386;
assign d30747 = hmaster0_p & d30744 | !hmaster0_p & d3072e;
assign v1446228 = hlock2 & v1446224 | !hlock2 & v1446222;
assign v121608b = hbusreq2 & v1216086 | !hbusreq2 & v121608a;
assign a65409 = hmaster0_p & a6587e | !hmaster0_p & a65890;
assign v15157ce = hgrant5_p & v845542 | !hgrant5_p & !v15157cc;
assign v15534ef = hlock0 & v15534ee | !hlock0 & v15534ed;
assign v1515646 = decide_p & v1515645 | !decide_p & v845542;
assign v144554e = hgrant2_p & v1445bec | !hgrant2_p & v144554d;
assign v1445450 = hlock3 & v144544b | !hlock3 & v144544f;
assign v14457c6 = hmaster1_p & v14457a6 | !hmaster1_p & v1445e28;
assign v10d42a0 = hgrant5_p & v10d3fe8 | !hgrant5_p & v10d429f;
assign v1668ce3 = hlock0_p & v1668cdd | !hlock0_p & v845542;
assign v1214d00 = hgrant1_p & v1214c36 | !hgrant1_p & v1214cff;
assign v1552d64 = hbusreq2_p & v1552d62 | !hbusreq2_p & v1552d63;
assign a65377 = hgrant1_p & a65362 | !hgrant1_p & !a65376;
assign v12161ee = hgrant1_p & v845542 | !hgrant1_p & v12161ed;
assign v1214fe5 = hgrant4_p & v845542 | !hgrant4_p & v1214fe4;
assign v1446630 = hmaster0_p & v14465e6 | !hmaster0_p & v144662f;
assign v1445a50 = hmaster0_p & v14458d4 | !hmaster0_p & v1445a4f;
assign d2fc24 = hmaster2_p & v84554a | !hmaster2_p & !v845542;
assign v1553155 = hmaster0_p & v1553150 | !hmaster0_p & v1553140;
assign v1214f18 = hgrant2_p & v845542 | !hgrant2_p & v1214f17;
assign a6588d = locked_p & a6588a | !locked_p & !v845542;
assign a653d6 = hbusreq5_p & a653d3 | !hbusreq5_p & a653d5;
assign v134d51f = hmaster1_p & v134d369 | !hmaster1_p & v134d51e;
assign v1445da2 = hmaster2_p & v14463b9 | !hmaster2_p & v1445da1;
assign v14461ea = hbusreq2_p & v14461e1 | !hbusreq2_p & v14461e9;
assign v10d404d = hgrant5_p & v10d3ffa | !hgrant5_p & !v10d404b;
assign a6569e = hmaster1_p & a658e8 | !hmaster1_p & !a65916;
assign v151562a = hmaster1_p & v1515629 | !hmaster1_p & v845570;
assign v1445a6c = hmaster0_p & v14458d4 | !hmaster0_p & v1445a6b;
assign v1668d40 = hbusreq5_p & v1668d3e | !hbusreq5_p & v1668d3f;
assign v1216b0d = hmaster0_p & v1216b03 | !hmaster0_p & v1216ab3;
assign v1445fd3 = hlock0 & v1445fd2 | !hlock0 & v1445fce;
assign v1445f1a = hlock3 & v1445edb | !hlock3 & v1445f19;
assign v16a1441 = hbusreq0 & v16a1440 | !hbusreq0 & v16a209b;
assign v1515797 = hgrant5_p & v845570 | !hgrant5_p & v1515796;
assign v1214c73 = hbusreq0 & v1214c72 | !hbusreq0 & v845542;
assign v1515aed = hbusreq2_p & v1515aec | !hbusreq2_p & !v845542;
assign bf1f9d = hbusreq4_p & v845570 | !hbusreq4_p & bf1f9c;
assign v1215cef = hlock5_p & v1215cee | !hlock5_p & !v1215ca8;
assign v1214d6a = hbusreq2 & v1214d66 | !hbusreq2 & v1214d69;
assign v1445a90 = hbusreq2_p & v1445a84 | !hbusreq2_p & v1445a8f;
assign v15167f2 = hmaster0_p & v845570 | !hmaster0_p & v1668c18;
assign v144589a = hlock1 & v1445891 | !hlock1 & v1445899;
assign d300d7 = hlock1_p & d300d5 | !hlock1_p & d300d6;
assign f2f291 = hbusreq3_p & f2f280 | !hbusreq3_p & f2f290;
assign v144670c = hmaster1_p & v144670b | !hmaster1_p & v1446436;
assign f2e4df = decide_p & f2e4de | !decide_p & f2f23c;
assign v144668e = hgrant5_p & v1446688 | !hgrant5_p & v144668d;
assign v14457ba = hmaster1_p & v144578c | !hmaster1_p & v1445e28;
assign d2fc45 = hbusreq2 & d2fc43 | !hbusreq2 & d2fc44;
assign v1216167 = hlock1_p & v1216163 | !hlock1_p & v1216166;
assign v121620c = hgrant5_p & v121620a | !hgrant5_p & v121620b;
assign v10d40d2 = hmaster1_p & v10d40d1 | !hmaster1_p & !v10d3fe9;
assign v134d442 = hmaster1_p & v134d441 | !hmaster1_p & v845542;
assign d30638 = hmaster0_p & d3060c | !hmaster0_p & d30613;
assign v1216abc = hbusreq1 & v1216aad | !hbusreq1 & v1216abb;
assign v12ad5d5 = hlock0_p & v1515762 | !hlock0_p & !v845542;
assign f2ed96 = hbusreq5_p & f2f236 | !hbusreq5_p & f2f288;
assign v15157b7 = hburst0 & a66293 | !hburst0 & v15157b6;
assign d30609 = hmaster1_p & d305ed | !hmaster1_p & d30608;
assign v134d3e1 = hbusreq5_p & v134d280 | !hbusreq5_p & v134d3e0;
assign v1445548 = hgrant2_p & v1445be3 | !hgrant2_p & v1445547;
assign v16a1bb3 = hready_p & v845555 | !hready_p & v16a1bb2;
assign d30667 = hgrant4_p & a66284 | !hgrant4_p & !d30666;
assign v10d40c2 = hmaster2_p & v10d40c1 | !hmaster2_p & v10d403a;
assign v10d4031 = hbusreq1_p & v10d4023 | !hbusreq1_p & v10d4030;
assign v15156eb = hmaster1_p & v15156c9 | !hmaster1_p & v15156e5;
assign v1214c1f = hmaster0_p & v1214bf1 | !hmaster0_p & v12153b1;
assign d30868 = hbusreq1_p & d30724 | !hbusreq1_p & d3068f;
assign v134d4cd = hmaster2_p & v845542 | !hmaster2_p & v134d4cc;
assign v1215363 = hbusreq3 & v121535c | !hbusreq3 & v1215362;
assign v12ad021 = hmaster0_p & v12ad61d | !hmaster0_p & v12ad602;
assign v1215c61 = hgrant5_p & v1215c5b | !hgrant5_p & v1215c1b;
assign v15167f5 = hgrant2_p & v15167f4 | !hgrant2_p & !v845542;
assign v138a3f1 = hmaster0_p & v1668c1f | !hmaster0_p & v138a309;
assign d2ff09 = hbusreq2 & d2ff05 | !hbusreq2 & d2ff08;
assign f2f2ca = hbusreq1 & a658b5 | !hbusreq1 & v845542;
assign v1214c3f = hbusreq2_p & v1214c3a | !hbusreq2_p & v1214c3e;
assign v16a13e2 = hmaster2_p & v16a2085 | !hmaster2_p & v16a208a;
assign d305ff = hbusreq5_p & d305fd | !hbusreq5_p & d305fe;
assign v1445fe6 = hbusreq2_p & v1445fdf | !hbusreq2_p & v1445fe5;
assign v12153cd = hbusreq4 & v1216048 | !hbusreq4 & v845547;
assign v12ad554 = hmaster1_p & v12ad532 | !hmaster1_p & v12ad54f;
assign v14466bf = hbusreq3 & v14466bd | !hbusreq3 & v14466be;
assign v16a1427 = hbusreq2 & v16a1426 | !hbusreq2 & !v16a1f9b;
assign v144545b = hlock3 & v1445456 | !hlock3 & v144545a;
assign d2ff0a = hbusreq5 & d2ff01 | !hbusreq5 & d2ff09;
assign v151561d = hmaster2_p & v845570 | !hmaster2_p & v151561c;
assign d2fb98 = hbusreq3 & d2fb8a | !hbusreq3 & d2fb97;
assign a654b5 = hmaster1_p & a6548c | !hmaster1_p & !a654b0;
assign v16a20a3 = hgrant2_p & v845542 | !hgrant2_p & !v16a20a1;
assign v12ad5a4 = hbusreq0_p & v1515790 | !hbusreq0_p & !v845542;
assign v138a2fb = hmaster0_p & v138a2f8 | !hmaster0_p & v138a2fa;
assign v1389389 = hbusreq0 & v1389de1 | !hbusreq0 & v138a403;
assign v15156bd = hmaster0_p & v15156bc | !hmaster0_p & v151564f;
assign v14462a2 = hlock5 & v1446275 | !hlock5 & v14462a0;
assign v1215018 = hgrant2_p & v1214fe2 | !hgrant2_p & v1215017;
assign a654b9 = hbusreq2 & a654b4 | !hbusreq2 & a654b8;
assign v12afe56 = hgrant1_p & v845542 | !hgrant1_p & v12afe55;
assign v1215bf2 = hmaster2_p & v1215bf1 | !hmaster2_p & v845542;
assign v134ce65 = hgrant2_p & v134ce56 | !hgrant2_p & v134ce63;
assign v1553090 = hlock2 & v1553061 | !hlock2 & v155308f;
assign v1216153 = hbusreq1 & v1216152 | !hbusreq1 & v845542;
assign a65645 = hgrant1_p & a653c7 | !hgrant1_p & !a65644;
assign v15534d6 = hgrant1_p & v845542 | !hgrant1_p & v15534d5;
assign v1668ca5 = hmaster1_p & v1668c75 | !hmaster1_p & !v1668c9c;
assign v1215c85 = hlock2_p & v1215c84 | !hlock2_p & !v845542;
assign v1446144 = hmaster1_p & v144611d | !hmaster1_p & v1445ffc;
assign v144588e = hbusreq0 & v1445878 | !hbusreq0 & v144588d;
assign v1284c90 = hmaster2_p & v140583c | !hmaster2_p & !v1284c8f;
assign v12aec4d = hbusreq3 & v12aec4a | !hbusreq3 & v12afe72;
assign a654bb = hmaster1_p & a65495 | !hmaster1_p & !a654b0;
assign v1216717 = hmaster2_p & v1216716 | !hmaster2_p & v845542;
assign v1284c9f = hmaster2_p & v1405844 | !hmaster2_p & !v1284c9a;
assign v16a12f8 = hbusreq5 & v16a12f1 | !hbusreq5 & v16a12f7;
assign v1446282 = hmaster0_p & v144639c | !hmaster0_p & v1446281;
assign d2fd4e = jx1_p & d2fc82 | !jx1_p & d2fd4d;
assign v144543e = hgrant3_p & v1445403 | !hgrant3_p & v144543d;
assign d2fb3a = hbusreq5_p & d2fec4 | !hbusreq5_p & d2fb39;
assign v1214cbd = hgrant4_p & v121537c | !hgrant4_p & v845572;
assign d2fb30 = hbusreq2_p & d2fb2e | !hbusreq2_p & d2fb2f;
assign f2f386 = hgrant5_p & f2f385 | !hgrant5_p & !f2f37f;
assign v12af227 = hbusreq0 & v12af21f | !hbusreq0 & v12af226;
assign v12af9d9 = hgrant2_p & v12af73f | !hgrant2_p & v12af9d8;
assign v1445f55 = hmaster1_p & v1445f54 | !hmaster1_p & v1446436;
assign v1445f4a = hmaster1_p & v1445f49 | !hmaster1_p & v1445da4;
assign v1668c4a = hmaster2_p & v845542 | !hmaster2_p & !v1668c49;
assign v1445833 = hgrant2_p & v1445831 | !hgrant2_p & v1445832;
assign v10d42da = hmaster1_p & v10d42b8 | !hmaster1_p & v10d407c;
assign v12160ff = hbusreq1_p & v12160fe | !hbusreq1_p & v845542;
assign v134d53c = hready_p & v134d530 | !hready_p & v134d53b;
assign d2fb37 = hbusreq4_p & d2fec2 | !hbusreq4_p & v84554a;
assign v1445401 = hbusreq5 & v14453ff | !hbusreq5 & v1445400;
assign v144672b = hmaster1_p & v144672a | !hmaster1_p & v1446436;
assign v16a1ca5 = hmaster1_p & v16a1ca4 | !hmaster1_p & !v16a2672;
assign v15534d2 = hgrant5_p & v845542 | !hgrant5_p & v15534d1;
assign v1215d0c = hbusreq5 & v1215ce0 | !hbusreq5 & v1215d0b;
assign jx1 = v1284d69;
assign v16a13f7 = hmaster0_p & v16a13f4 | !hmaster0_p & v16a13f6;
assign v1445917 = hmaster2_p & v1445906 | !hmaster2_p & v14458e5;
assign v151567f = hmaster0_p & v151567e | !hmaster0_p & v1515675;
assign v12af9b7 = hbusreq5 & v12af98f | !hbusreq5 & v12af9b6;
assign v16a12c5 = hbusreq2 & v16a12c3 | !hbusreq2 & v16a12c4;
assign v1284cb5 = hmaster0_p & v1284ca9 | !hmaster0_p & v1284cad;
assign v12165b0 = hmaster1_p & v12165af | !hmaster1_p & v12165a5;
assign d30286 = hgrant2_p & v845542 | !hgrant2_p & !d30284;
assign d307eb = hlock1_p & d307ea | !hlock1_p & d30667;
assign v15530e8 = hbusreq2_p & v1552d4e | !hbusreq2_p & v155341e;
assign v1446014 = hgrant1_p & v845542 | !hgrant1_p & v1446013;
assign d30271 = hlock5_p & d3026f | !hlock5_p & !d30270;
assign v14458d0 = hlock5 & v14458b3 | !hlock5 & v14458ce;
assign d80778 = hbusreq5_p & d80777 | !hbusreq5_p & !d80776;
assign v16a1d68 = hbusreq5 & v16a1d57 | !hbusreq5 & v16a1d67;
assign v1214c37 = hmaster2_p & v1214c36 | !hmaster2_p & v845542;
assign v1214d05 = hmaster1_p & v1214cef | !hmaster1_p & v1214d04;
assign d3026c = hlock5_p & d3026a | !hlock5_p & !d3026b;
assign v1553051 = hgrant1_p & v1553050 | !hgrant1_p & v845542;
assign v16a1afe = hmaster0_p & v16a1afb | !hmaster0_p & v16a1afd;
assign v14459b6 = hlock0_p & v14459b4 | !hlock0_p & v14459b5;
assign a65915 = hbusreq5_p & a65912 | !hbusreq5_p & a65913;
assign v12ad515 = hbusreq0_p & a658b5 | !hbusreq0_p & v845542;
assign d2fbb7 = hlock2_p & d2fbb6 | !hlock2_p & d2fbb2;
assign v138a436 = hgrant3_p & v138a3c2 | !hgrant3_p & v138a435;
assign v1284d66 = hbusreq3_p & v1284d2a | !hbusreq3_p & v1284d65;
assign v14463d4 = hlock3 & v14463d1 | !hlock3 & v14463d3;
assign v134d266 = hmaster1_p & v134d265 | !hmaster1_p & v134d208;
assign d2fb77 = hlock4_p & d2fb76 | !hlock4_p & v84554a;
assign v1405ad1 = hmaster1_p & v1405ad0 | !hmaster1_p & !v1405a94;
assign v121639e = hmaster2_p & v845542 | !hmaster2_p & !v1216ac7;
assign v16a1f98 = hmaster1_p & v845564 | !hmaster1_p & !v16a1f96;
assign v138a2ff = hlock5_p & v1515615 | !hlock5_p & v845570;
assign v144541e = hgrant2_p & v1445be3 | !hgrant2_p & v144541d;
assign d30119 = hmaster2_p & d300cd | !hmaster2_p & d300f2;
assign v14453b3 = hgrant2_p & v144538d | !hgrant2_p & v14453b2;
assign d2fb23 = hbusreq5_p & d30141 | !hbusreq5_p & d2fb22;
assign v1215755 = hbusreq1 & v1215b86 | !hbusreq1 & v845542;
assign d30660 = hbusreq4_p & v84555a | !hbusreq4_p & !v845542;
assign v1215735 = hbusreq1 & v1215734 | !hbusreq1 & v1215b97;
assign v10d42cb = hgrant5_p & v10d3ffd | !hgrant5_p & !v10d42ca;
assign v1445541 = hready_p & v144639b | !hready_p & v1445540;
assign v1214f38 = hmaster0_p & v1215d30 | !hmaster0_p & v1215d2f;
assign v14458e2 = hlock0_p & v1446407 | !hlock0_p & v14458e1;
assign v12ad671 = hmastlock_p & v12ad670 | !hmastlock_p & v845542;
assign bf1f91 = hgrant1_p & f2f227 | !hgrant1_p & bf1f90;
assign v1215c8a = hgrant5_p & v845542 | !hgrant5_p & !v1215c88;
assign v1214bb7 = hmaster2_p & v1215392 | !hmaster2_p & v1215364;
assign v144640a = hbusreq4 & v1446408 | !hbusreq4 & v1446409;
assign v1405940 = hbusreq3_p & v1405905 | !hbusreq3_p & v140593f;
assign v12160c4 = hmaster1_p & v12160af | !hmaster1_p & v1216082;
assign f2f3f8 = hbusreq2 & f2f3f2 | !hbusreq2 & f2f3f7;
assign bf1f93 = hgrant5_p & v845542 | !hgrant5_p & !bf1f92;
assign v16a194b = hgrant4_p & v845559 | !hgrant4_p & !v16a194a;
assign v1668c6a = hburst0 & a66272 | !hburst0 & v1668c69;
assign v16a1b62 = hbusreq2 & v16a1b02 | !hbusreq2 & v16a1b03;
assign d30110 = hgrant2_p & d300b4 | !hgrant2_p & d3010f;
assign v134d1e6 = stateG3_2_p & v845542 | !stateG3_2_p & !v134d1e5;
assign v1445bd4 = hbusreq5_p & v1446042 | !hbusreq5_p & v1445bd3;
assign d30224 = hgrant5_p & d30223 | !hgrant5_p & !d30221;
assign v1405ac2 = hmaster2_p & v1405abf | !hmaster2_p & v1405ac0;
assign v10d40b6 = hmaster1_p & v10d40b5 | !hmaster1_p & !v10d404f;
assign d2fd49 = decide_p & d2fd48 | !decide_p & v845570;
assign d300b7 = hlock1_p & d300b5 | !hlock1_p & !d300b6;
assign v16a1d01 = decide_p & v16a1ce7 | !decide_p & !v16a1cc6;
assign d30709 = hmaster0_p & d306fd | !hmaster0_p & d30708;
assign v151699c = hbusreq2_p & v151699b | !hbusreq2_p & v845542;
assign v121630c = hmaster2_p & v1216048 | !hmaster2_p & v1216aea;
assign a662b8 = hmaster1_p & a662ae | !hmaster1_p & a662b7;
assign v16a1dd3 = hbusreq3 & v16a1dbf | !hbusreq3 & v16a1dd2;
assign v1445d92 = hgrant5_p & v1445d8f | !hgrant5_p & !v1445d91;
assign a656a1 = hmaster1_p & a65687 | !hmaster1_p & !a65916;
assign v12ad51c = hbusreq1_p & v12ad51b | !hbusreq1_p & !v1668c63;
assign v1445ad4 = hlock2 & v1445ad1 | !hlock2 & v1445ad3;
assign v1214db8 = hmaster1_p & v1214d0d | !hmaster1_p & !v1214d1e;
assign d302f9 = jx1_p & d308d4 | !jx1_p & d302f8;
assign v1446294 = hmaster1_p & v144626e | !hmaster1_p & v1446290;
assign v138a3ea = hlock5_p & v138a3e9 | !hlock5_p & !v151579c;
assign a65666 = hgrant5_p & v845558 | !hgrant5_p & !a65624;
assign f2e4f8 = decide_p & f2e4e7 | !decide_p & f2f23c;
assign v12153f2 = hbusreq2_p & v12153f1 | !hbusreq2_p & v12153f0;
assign v12add4a = hbusreq0 & v12adf5e | !hbusreq0 & v12add49;
assign d2fd2e = hbusreq2 & d2fd2d | !hbusreq2 & d302f3;
assign v138a34d = hmaster1_p & v138a34c | !hmaster1_p & v138a341;
assign d3075d = hmaster1_p & d30745 | !hmaster1_p & d30754;
assign v1214d4c = hmaster1_p & v12153ab | !hmaster1_p & v1214d4b;
assign f2f298 = hmaster2_p & f2f293 | !hmaster2_p & v845542;
assign v1405b40 = hmaster1_p & v1405b3f | !hmaster1_p & !v1405a94;
assign f2f33c = hmaster1_p & f2f328 | !hmaster1_p & !f2f330;
assign v1216246 = hbusreq2 & v1216242 | !hbusreq2 & v1216245;
assign v16a1e7a = hbusreq5 & v16a1e6e | !hbusreq5 & v16a1e79;
assign v1446085 = hbusreq2_p & v1446075 | !hbusreq2_p & v1446084;
assign v16a1396 = hbusreq2 & v16a1395 | !hbusreq2 & v16a12c4;
assign d302df = hlock5_p & d302de | !hlock5_p & d30656;
assign v16a1dbc = hgrant3_p & v16a1daf | !hgrant3_p & v16a1dbb;
assign v1445507 = hmaster1_p & v1445506 | !hmaster1_p & v14462ff;
assign v1405882 = hready_p & v140585e | !hready_p & v1405881;
assign v144632f = hbusreq2_p & v144632b | !hbusreq2_p & v144632e;
assign v12ad036 = decide_p & v12ad035 | !decide_p & v12afe76;
assign v1553438 = hbusreq0_p & v1553138 | !hbusreq0_p & v845542;
assign v1445e02 = hbusreq4_p & v1446430 | !hbusreq4_p & v1446429;
assign v16a1400 = hgrant2_p & v845542 | !hgrant2_p & v16a13ff;
assign v16a2246 = hbusreq5_p & v16a2245 | !hbusreq5_p & v845542;
assign v12ae1fa = hgrant4_p & v845542 | !hgrant4_p & !v12ae1f9;
assign f2eda4 = jx2_p & f2ed9f | !jx2_p & f2eda3;
assign v1215d04 = hmaster0_p & v1215ce6 | !hmaster0_p & v1215d03;
assign v144615e = hbusreq5 & v144615c | !hbusreq5 & v144615d;
assign v14463f0 = hmaster1_p & v144639c | !hmaster1_p & v14463ef;
assign a662c6 = hready_p & v845542 | !hready_p & a662c5;
assign v1552f6f = hlock0 & v1552f6e | !hlock0 & v1552f6d;
assign v12ad645 = hbusreq5_p & v12ad4fd | !hbusreq5_p & v12ad644;
assign v134cecd = hbusreq5 & v134cecb | !hbusreq5 & v134cecc;
assign a65426 = hgrant5_p & a65424 | !hgrant5_p & !a653b5;
assign v12ad5de = hgrant5_p & v12ad4fd | !hgrant5_p & v12ad5dc;
assign v1284d3d = hbusreq5_p & v1284cad | !hbusreq5_p & v1284d3c;
assign v1215385 = hbusreq4_p & v121537c | !hbusreq4_p & d2fbe5;
assign v121570a = hmaster1_p & v1215709 | !hmaster1_p & !v1215ba1;
assign v1446303 = hbusreq0 & v1446302 | !hbusreq0 & v14462e7;
assign d3069a = hbusreq5_p & v845542 | !hbusreq5_p & d3068a;
assign v1445840 = hlock3 & v14457f6 | !hlock3 & v144583e;
assign v1445fab = hmaster1_p & v1445faa | !hmaster1_p & v1445f9e;
assign f2f367 = hbusreq1 & v1668d4a | !hbusreq1 & v845542;
assign d2ff0c = decide_p & d2ff0b | !decide_p & v845570;
assign v16a1e91 = hgrant5_p & v845542 | !hgrant5_p & v16a1e90;
assign v121624e = hmaster1_p & v121622c | !hmaster1_p & !v121624b;
assign v16a2079 = hlock5_p & v16a2071 | !hlock5_p & v16a2078;
assign d306bd = hbusreq5_p & v845542 | !hbusreq5_p & !d306ac;
assign v10d42d1 = hmaster1_p & v10d42d0 | !hmaster1_p & !v10d42a1;
assign d2fec7 = hmaster1_p & d2feb5 | !hmaster1_p & d2fec6;
assign v1446019 = hgrant2_p & v1446461 | !hgrant2_p & v1446018;
assign v1445ec5 = hmaster1_p & v1445ec4 | !hmaster1_p & v1445e07;
assign v1445fd8 = hbusreq1_p & v1446423 | !hbusreq1_p & v1446429;
assign a653ba = hgrant5_p & a65390 | !hgrant5_p & a653b9;
assign v1216a85 = stateG3_0_p & v845586 | !stateG3_0_p & !v84556c;
assign v121505f = hbusreq2_p & v1215056 | !hbusreq2_p & v121505e;
assign v1668da2 = hmaster0_p & v1668d34 | !hmaster0_p & v1668da1;
assign v1405ad0 = hmaster0_p & v1405a8a | !hmaster0_p & v1405a89;
assign v1216262 = hgrant5_p & v12160e2 | !hgrant5_p & v1216261;
assign d30736 = hmaster0_p & d3071e | !hmaster0_p & d30735;
assign v1445dcf = hbusreq0 & v1445dce | !hbusreq0 & v1445d93;
assign v1445fc7 = hbusreq3 & v1445fc5 | !hbusreq3 & v1445fc6;
assign v14464a1 = hmaster0_p & v144647c | !hmaster0_p & v14464a0;
assign v14458ea = hbusreq5_p & v14458e6 | !hbusreq5_p & v14458e9;
assign v12ad03b = hgrant3_p & v12acff0 | !hgrant3_p & v12ad03a;
assign v140587e = hmaster2_p & v140587c | !hmaster2_p & !v1446403;
assign v134d377 = hgrant1_p & v134d273 | !hgrant1_p & v845542;
assign v134cea2 = hmaster1_p & v134ce84 | !hmaster1_p & v134ce9d;
assign d2fc62 = stateG10_5_p & d2fc60 | !stateG10_5_p & d2fc61;
assign d2febf = hlock4_p & v845542 | !hlock4_p & d305fb;
assign d30778 = hbusreq2 & d30774 | !hbusreq2 & d30777;
assign v1515820 = hmaster0_p & v151581f | !hmaster0_p & v151564f;
assign d306df = hlock0_p & v845542 | !hlock0_p & d306de;
assign v14459d0 = hmaster2_p & v14465b3 | !hmaster2_p & v14459cf;
assign v1515774 = hgrant1_p & v151576a | !hgrant1_p & v1515773;
assign v134d4ed = hmaster2_p & v134d4e8 | !hmaster2_p & v845542;
assign v1284cf2 = hbusreq5_p & v1284ced | !hbusreq5_p & v1284cf0;
assign v1445815 = hmaster1_p & v1445814 | !hmaster1_p & v1445e07;
assign d30160 = hbusreq2_p & d3015e | !hbusreq2_p & d3015f;
assign v14463e1 = hbusreq4 & v14463e0 | !hbusreq4 & v144639f;
assign a6542d = hbusreq5_p & a65429 | !hbusreq5_p & !a6542b;
assign v12ad5e8 = hmaster2_p & v12ad5a8 | !hmaster2_p & v12ad5cb;
assign v1215315 = hmaster0_p & v121501d | !hmaster0_p & v1214fed;
assign v138a3d8 = hbusreq0 & v138a3d1 | !hbusreq0 & v138a3d7;
assign v14058cd = hbusreq5_p & v14058c9 | !hbusreq5_p & v14058cc;
assign v12afe73 = hbusreq5 & v12afe68 | !hbusreq5 & v12afe72;
assign v155313b = hmaster1_p & v155313a | !hmaster1_p & v845542;
assign v14454f7 = hmaster0_p & v14454ed | !hmaster0_p & v1445414;
assign d30955 = hlock5_p & d30953 | !hlock5_p & !d30954;
assign v16a2676 = hmaster0_p & v16a266a | !hmaster0_p & v16a2675;
assign v134d221 = hbusreq5_p & v134d220 | !hbusreq5_p & v134d1e8;
assign f2f4af = hburst0 & a658a5 | !hburst0 & f2f4ae;
assign d2fd23 = hbusreq5_p & d2fd22 | !hbusreq5_p & !d2fd21;
assign d2fb41 = hbusreq5_p & d2fee3 | !hbusreq5_p & d2fb35;
assign v1446710 = hbusreq2 & v144670e | !hbusreq2 & v144670f;
assign v1216530 = hgrant5_p & v845542 | !hgrant5_p & v121652f;
assign d2f992 = hbusreq4_p & d2f991 | !hbusreq4_p & v845542;
assign v1405b2f = hmaster1_p & v1405b2e | !hmaster1_p & v1405b29;
assign v1445fa4 = hmaster1_p & v1445fa3 | !hmaster1_p & v1445f9e;
assign f2f381 = hbusreq1 & v1668d63 | !hbusreq1 & v845542;
assign d2fed4 = hbusreq2 & d2fecc | !hbusreq2 & d2fed3;
assign d80798 = hgrant4_p & v845542 | !hgrant4_p & !d80797;
assign v12167a7 = hmaster1_p & v12167a6 | !hmaster1_p & v1216a9b;
assign d30876 = hmaster1_p & d30865 | !hmaster1_p & d30875;
assign d2f9d8 = decide_p & d2f9d7 | !decide_p & v845570;
assign v16a12c1 = hmaster1_p & v16a1a98 | !hmaster1_p & v16a1f96;
assign v1214f0d = hbusreq0 & v1214f08 | !hbusreq0 & v1214f0c;
assign v1445ee7 = hbusreq3 & v1445ee5 | !hbusreq3 & v1445ee6;
assign v1214da0 = hgrant2_p & v1214d9d | !hgrant2_p & v1214d9f;
assign f2f4b5 = hmaster0_p & f2f4b4 | !hmaster0_p & v845542;
assign v10d4071 = hbusreq4_p & v10d3fd9 | !hbusreq4_p & !v10d3fdf;
assign a653a7 = hmaster2_p & a65377 | !hmaster2_p & a653a3;
assign v16a1e72 = hbusreq2_p & v16a1dd4 | !hbusreq2_p & v16a1e71;
assign v12166cb = stateA1_p & d30714 | !stateA1_p & !v845542;
assign v144544c = hmaster1_p & v1445443 | !hmaster1_p & v1446236;
assign a65ad7 = hmaster0_p & a662cd | !hmaster0_p & a65ad6;
assign d30687 = decide_p & d30686 | !decide_p & v845570;
assign v151576e = hlock0_p & v1668d25 | !hlock0_p & v151576d;
assign v1445b68 = hbusreq2_p & v1445b64 | !hbusreq2_p & v1445b67;
assign v1215be1 = hmaster2_p & v1215ffd | !hmaster2_p & v1216004;
assign v1445e31 = hlock3 & v1445e1f | !hlock3 & v1445e30;
assign d308bc = hbusreq0 & d308b9 | !hbusreq0 & d308bb;
assign a6587f = hburst0_p & v845542 | !hburst0_p & !v155392f;
assign v1284ca1 = hgrant5_p & v1284c9e | !hgrant5_p & !v1284ca0;
assign v1446255 = hmaster1_p & v144623a | !hmaster1_p & v1446250;
assign f2e4d9 = hgrant5_p & v845542 | !hgrant5_p & !f2e4d8;
assign v15530fe = hmaster1_p & v15530fd | !hmaster1_p & v845542;
assign v1668cc5 = hbusreq1 & v1668cbd | !hbusreq1 & !v1668cc4;
assign v1216713 = hbusreq3 & v1216707 | !hbusreq3 & v1216712;
assign v1445aca = hlock2 & v1445abf | !hlock2 & v1445ac8;
assign v10d3ff3 = hbusreq1_p & v10d3fd8 | !hbusreq1_p & !v10d3fdf;
assign v1552d87 = hbusreq0_p & v1553138 | !hbusreq0_p & v1552d7c;
assign v15530f3 = decide_p & v1553216 | !decide_p & v15530f2;
assign v1446301 = hgrant2_p & v14462e9 | !hgrant2_p & v1446300;
assign f2f45a = hbusreq2_p & f2f458 | !hbusreq2_p & !f2f459;
assign f2f462 = jx2_p & f2f291 | !jx2_p & f2f461;
assign v1215326 = hgrant2_p & v1215324 | !hgrant2_p & v1215325;
assign a6548a = hbusreq2_p & a65478 | !hbusreq2_p & a65479;
assign v121576c = hgrant5_p & v1215b87 | !hgrant5_p & v121576b;
assign v1215013 = hgrant1_p & v12153bd | !hgrant1_p & v1215012;
assign v1405b4c = hgrant4_p & v1405a86 | !hgrant4_p & v1405b4b;
assign v12ad5d2 = hbusreq1_p & v12ad5d0 | !hbusreq1_p & v12ad5d1;
assign v1215cc2 = hgrant1_p & v1215cbb | !hgrant1_p & v1216165;
assign v16a1889 = hmaster1_p & v16a1840 | !hmaster1_p & !v16a1f96;
assign v16a1bfa = hbusreq2 & v16a1bf8 | !hbusreq2 & !v16a1bf9;
assign v16a2669 = hmaster2_p & v16a2668 | !hmaster2_p & !v845542;
assign v134d292 = hmaster2_p & v134d28d | !hmaster2_p & v134d291;
assign v1215dae = decide_p & v1215bd5 | !decide_p & v1215dad;
assign v10d4058 = hbusreq5_p & v10d4056 | !hbusreq5_p & !v10d4057;
assign v16a1d30 = hbusreq3 & v16a1d2f | !hbusreq3 & v16a205d;
assign v12acfd4 = hbusreq2_p & v12acfd2 | !hbusreq2_p & v12acfd3;
assign v1445fe2 = hbusreq0 & v1445fe0 | !hbusreq0 & v1445fe1;
assign v12ad5d9 = hbusreq4_p & v12ad5ae | !hbusreq4_p & v12ad5c1;
assign v1445f6d = hlock2 & v1445f68 | !hlock2 & v1445f6c;
assign v12acfc3 = hbusreq5_p & v12ad535 | !hbusreq5_p & v12acfc2;
assign d2faf9 = hbusreq5_p & d300e3 | !hbusreq5_p & d2faf8;
assign v16a1335 = hgrant2_p & v16a205b | !hgrant2_p & v16a1334;
assign v144589e = hlock0 & v1445896 | !hlock0 & v144589d;
assign v144545a = hbusreq2 & v1445445 | !hbusreq2 & v1445459;
assign d2fc30 = hbusreq5_p & d2fb7d | !hbusreq5_p & d2fc2f;
assign d30145 = hgrant5_p & d2fe96 | !hgrant5_p & d300ff;
assign d308c7 = hmaster0_p & d308c1 | !hmaster0_p & d308c6;
assign v1216278 = decide_p & v1216272 | !decide_p & !v1216277;
assign v14466f4 = hbusreq2_p & v14466f1 | !hbusreq2_p & v14466f3;
assign v1446738 = hmaster0_p & v1446648 | !hmaster0_p & v14465b8;
assign v15157cb = hgrant1_p & f2f281 | !hgrant1_p & v15157ca;
assign v1445865 = hbusreq3 & v1445863 | !hbusreq3 & v1445864;
assign v134cf6f = jx1_p & v134ce80 | !jx1_p & v134cf6e;
assign d30810 = hlock2_p & d3080d | !hlock2_p & d3080f;
assign v121657f = hgrant2_p & v121657e | !hgrant2_p & v1216576;
assign v12afa0a = hbusreq5_p & v12afe63 | !hbusreq5_p & v12af9d4;
assign v16a1e8a = hready_p & v845555 | !hready_p & v16a1e89;
assign v121543b = hmaster2_p & v1215438 | !hmaster2_p & v1215b97;
assign v1552d61 = hmaster1_p & v1553385 | !hmaster1_p & v1552d60;
assign v1215cb8 = hbusreq0 & v1215cac | !hbusreq0 & v1215cb7;
assign v16a1d3e = hgrant5_p & v845542 | !hgrant5_p & v16a1d3d;
assign d3074f = hbusreq2 & d3074a | !hbusreq2 & d3074e;
assign a6536d = locked_p & a65369 | !locked_p & !v845542;
assign v12161a2 = hmaster0_p & v121618e | !hmaster0_p & v12161a1;
assign v144551a = hlock2 & v14454fa | !hlock2 & v1445519;
assign v16a19b9 = hgrant2_p & v16a205c | !hgrant2_p & v16a19b8;
assign v10d408d = hmaster1_p & v10d408c | !hmaster1_p & v10d407c;
assign v134d527 = hlock3 & v134d524 | !hlock3 & v134d526;
assign v1553390 = hgrant1_p & v155338f | !hgrant1_p & v845542;
assign v15155fe = hmaster0_p & v15155f7 | !hmaster0_p & v15155fd;
assign v121537e = hbusreq0 & v121537d | !hbusreq0 & v845542;
assign v1216004 = hlock0_p & v1216a5a | !hlock0_p & v1216003;
assign d2fe97 = hmaster0_p & d2fe80 | !hmaster0_p & d2fe96;
assign f2f4c3 = decide_p & f2f4c2 | !decide_p & v845542;
assign v10d4027 = hgrant5_p & v10d3ff1 | !hgrant5_p & !v10d4025;
assign v14461e6 = hgrant2_p & v14461b8 | !hgrant2_p & v14461e5;
assign a65621 = hgrant4_p & a662a9 | !hgrant4_p & !a65863;
assign v12aef09 = decide_p & v12af3ac | !decide_p & v12afe76;
assign a658cf = hmaster2_p & a658b6 | !hmaster2_p & a658ce;
assign v1445b1d = hbusreq2 & v1445b1b | !hbusreq2 & v1445b1c;
assign v1445dff = hmaster2_p & v1446427 | !hmaster2_p & v1445dfe;
assign v1214cfd = hbusreq0 & v1214cfc | !hbusreq0 & v845542;
assign v1405b1c = hmaster2_p & v845542 | !hmaster2_p & !v1405b1b;
assign v1552f72 = hgrant2_p & v1552f71 | !hgrant2_p & v1552f6a;
assign v1515752 = hgrant5_p & v151574c | !hgrant5_p & !v1515751;
assign a658e0 = hlock0_p & a658bd | !hlock0_p & a658de;
assign v1446006 = hbusreq3 & v1446004 | !hbusreq3 & v1446005;
assign a653fa = hgrant5_p & a653f9 | !hgrant5_p & a653f5;
assign d301d4 = hgrant5_p & v845580 | !hgrant5_p & !d301d2;
assign v16a13cc = hbusreq3 & v16a13c3 | !hbusreq3 & v16a13cb;
assign f2f431 = hmaster2_p & f2f42f | !hmaster2_p & f2f430;
assign v1445518 = hgrant2_p & v1445516 | !hgrant2_p & v1445517;
assign v1215d99 = hgrant5_p & v1215d97 | !hgrant5_p & !v1215d98;
assign v1284d25 = hmaster1_p & v1284d24 | !hmaster1_p & !v1284d1f;
assign v15532c6 = hgrant0_p & v1553138 | !hgrant0_p & v845542;
assign v138a43b = hmaster0_p & v138a439 | !hmaster0_p & v138a43a;
assign d2fcfc = hlock5_p & d2fcfb | !hlock5_p & d2fcb1;
assign v144640e = hlock1 & v1446407 | !hlock1 & v144640c;
assign v16a1434 = hgrant3_p & v16a142b | !hgrant3_p & v16a1433;
assign v1215045 = hbusreq4_p & v1215044 | !hbusreq4_p & v845542;
assign d308a3 = hgrant5_p & d30856 | !hgrant5_p & d308a2;
assign v1668d97 = hmaster2_p & a65851 | !hmaster2_p & a65862;
assign v14466c8 = hgrant3_p & v144645f | !hgrant3_p & v14466c7;
assign v14457ce = hbusreq2 & v14457c8 | !hbusreq2 & v14457cd;
assign v1214cdd = hmaster0_p & v121537e | !hmaster0_p & v1214cdc;
assign v1552d90 = hgrant2_p & v155321e | !hgrant2_p & v1552d8f;
assign d308ac = hbusreq0 & d308a4 | !hbusreq0 & d308ab;
assign v14460f1 = hmaster1_p & v1445f85 | !hmaster1_p & v1445fae;
assign d80730 = stateG2_p & v845542 | !stateG2_p & !v936735;
assign d2fd39 = hbusreq2_p & v845552 | !hbusreq2_p & !v845542;
assign v13897e0 = hbusreq5_p & v13897df | !hbusreq5_p & !v845542;
assign v15157bd = hgrant1_p & f2f281 | !hgrant1_p & v15157bc;
assign v1214d30 = hbusreq3 & v1214d26 | !hbusreq3 & v1214d2f;
assign v10d4042 = hgrant4_p & v10d4040 | !hgrant4_p & !v10d4041;
assign v10d3fd5 = locked_p & v845542 | !locked_p & !v10d3fd4;
assign v16a1d82 = decide_p & v16a1d68 | !decide_p & v16a1d81;
assign v1446601 = hlock1 & v1446600 | !hlock1 & v14465fa;
assign d308b5 = hmaster0_p & d3083b | !hmaster0_p & d3081d;
assign d2fb45 = hbusreq2_p & d2ff07 | !hbusreq2_p & d2fb43;
assign v10d429c = hbusreq4_p & v10d4289 | !hbusreq4_p & v10d4292;
assign d2fbb0 = hmaster0_p & d2fb7e | !hmaster0_p & d2fb6c;
assign v10d40a3 = hbusreq2_p & v10d40a0 | !hbusreq2_p & v10d40a2;
assign d2fb8e = hmaster1_p & d2fb8d | !hmaster1_p & d2fb7b;
assign v1445515 = hbusreq2_p & v1445514 | !hbusreq2_p & v1445bdb;
assign v1405b08 = hgrant5_p & v1405a93 | !hgrant5_p & v1405b07;
assign a65af8 = hbusreq3_p & a65ae1 | !hbusreq3_p & a65af7;
assign v14466ad = hbusreq5_p & v14466ac | !hbusreq5_p & v1446643;
assign v1284d43 = hmaster1_p & v1284d42 | !hmaster1_p & v140584d;
assign v1445f72 = hmaster0_p & v1446663 | !hmaster0_p & v14466af;
assign d3074e = hbusreq2_p & d3074d | !hbusreq2_p & d30748;
assign d2fd0d = hbusreq3 & d2fd08 | !hbusreq3 & d2fd0c;
assign v1215c2e = hgrant1_p & v1215c25 | !hgrant1_p & v121615b;
assign v1446334 = hmaster1_p & v1446333 | !hmaster1_p & v144627e;
assign v1445bdb = hgrant2_p & v1445bd9 | !hgrant2_p & v1445bda;
assign v134d43d = hbusreq1_p & v134d43c | !hbusreq1_p & v134d273;
assign v1214e41 = hlock2_p & v1214e10 | !hlock2_p & !v1214e40;
assign d2fadc = hgrant1_p & d2fad8 | !hgrant1_p & d2fadb;
assign v1445ae7 = hmaster0_p & v1445a38 | !hmaster0_p & v1445902;
assign a65632 = hgrant5_p & a653f9 | !hgrant5_p & a65630;
assign v1215716 = hgrant4_p & v845542 | !hgrant4_p & v1215715;
assign v121506a = hbusreq2 & v121505f | !hbusreq2 & v1215069;
assign d301e8 = hlock1_p & d301e6 | !hlock1_p & d301e7;
assign v1215cd8 = hbusreq2_p & v1215cca | !hbusreq2_p & !v1215cd7;
assign v12153b7 = hbusreq1_p & v12153b4 | !hbusreq1_p & v1215bac;
assign v1215740 = hmaster2_p & v1215b97 | !hmaster2_p & v1215b9c;
assign v1215b8e = hready & v845542 | !hready & v1216567;
assign v12166f7 = hbusreq5_p & v12166f6 | !hbusreq5_p & v16a2243;
assign v1215046 = hgrant4_p & v845542 | !hgrant4_p & v1215045;
assign v1216b11 = hlock2_p & v1216b0e | !hlock2_p & v1216b10;
assign v1445e3c = hgrant5_p & v1446467 | !hgrant5_p & v1445e3b;
assign v1215348 = hmaster2_p & v1215345 | !hmaster2_p & v1215347;
assign v12add49 = hmaster2_p & v845542 | !hmaster2_p & v12add48;
assign v12162d2 = hbusreq2_p & v12162cf | !hbusreq2_p & v12162d1;
assign v1446725 = hmaster0_p & v1446440 | !hmaster0_p & v144639c;
assign v16a1321 = hready & v16a223a | !hready & v845542;
assign a65639 = hgrant5_p & a653ab | !hgrant5_p & !a65638;
assign v1445a9c = hmaster1_p & v14459a3 | !hmaster1_p & v1445a9b;
assign v1445bb2 = hmaster1_p & v1445bad | !hmaster1_p & v1445bb1;
assign v1552f60 = hbusreq4_p & v1552f5f | !hbusreq4_p & v15533a0;
assign d30632 = hbusreq5 & d30627 | !hbusreq5 & d30631;
assign v12ad013 = hmaster2_p & v12ad012 | !hmaster2_p & v12af9c1;
assign v1215d86 = hmaster1_p & v1215d85 | !hmaster1_p & v1215d68;
assign v144663d = hlock1 & v14465ce | !hlock1 & v14465c9;
assign v10d42c9 = hgrant1_p & v10d4019 | !hgrant1_p & v10d42c8;
assign v151583c = hmaster0_p & v151583b | !hmaster0_p & v151573b;
assign v1445f79 = hlock2 & v1445f75 | !hlock2 & v1445f78;
assign v1553223 = hmaster2_p & v1553222 | !hmaster2_p & v845542;
assign v1216577 = hgrant2_p & v1216520 | !hgrant2_p & v1216576;
assign v1215723 = hgrant5_p & v1215b7e | !hgrant5_p & v1215722;
assign v134d3c4 = hmaster1_p & v134d3c3 | !hmaster1_p & v134d208;
assign v1216b04 = hmaster0_p & v1216ab3 | !hmaster0_p & v1216b03;
assign d305ef = hmastlock_p & d305ee | !hmastlock_p & v845542;
assign v14460a8 = hgrant2_p & v14460a7 | !hgrant2_p & v1446094;
assign v15156fa = hmaster2_p & v151564d | !hmaster2_p & !a658dc;
assign v1405866 = hlock5_p & v1405864 | !hlock5_p & v1405865;
assign v12166d5 = hbusreq5_p & v12166d4 | !hbusreq5_p & v845542;
assign v151583d = hmaster1_p & v151583c | !hmaster1_p & v1515786;
assign v121546a = hbusreq5_p & v1215468 | !hbusreq5_p & v1215469;
assign v121502a = hgrant1_p & v121545f | !hgrant1_p & v1215029;
assign v121504b = hbusreq0_p & v121504a | !hbusreq0_p & v1215032;
assign v1284cc2 = hmaster0_p & v1405856 | !hmaster0_p & v1284c90;
assign v15156b7 = hburst1 & f2f4ad | !hburst1 & v15156b6;
assign v1445fdf = hmaster1_p & v1446405 | !hmaster1_p & v1445fde;
assign v1445a66 = hmaster0_p & v14459a2 | !hmaster0_p & v1445a3e;
assign v1215c58 = hgrant5_p & v845542 | !hgrant5_p & v1215c01;
assign v1216039 = hmaster0_p & v1216035 | !hmaster0_p & v1216038;
assign d30834 = hgrant5_p & v84554e | !hgrant5_p & d307fa;
assign d300b3 = hmaster1_p & d300b2 | !hmaster1_p & d2fe8c;
assign d30808 = hbusreq2_p & d307f6 | !hbusreq2_p & !d30807;
assign d30259 = hmaster1_p & d30258 | !hmaster1_p & d30250;
assign a656ac = hmaster1_p & a65691 | !hmaster1_p & !a65916;
assign v1405acf = hready_p & v1405a9f | !hready_p & v1405ace;
assign v16a1975 = hbusreq0 & v16a207a | !hbusreq0 & v16a1974;
assign v140591b = hmaster0_p & v140584f | !hmaster0_p & v1405840;
assign d2faff = hbusreq1 & d2f979 | !hbusreq1 & d30660;
assign d306aa = hgrant1_p & d30654 | !hgrant1_p & d306a6;
assign v1445a59 = hbusreq0 & v1445a55 | !hbusreq0 & v1445a58;
assign v15156af = hmaster2_p & v1668cd0 | !hmaster2_p & !v15156ae;
assign f2e734 = hgrant2_p & v845542 | !hgrant2_p & f2e733;
assign v12161cd = hmaster1_p & v12161cc | !hmaster1_p & v1216041;
assign v1446113 = hlock3 & v14460f2 | !hlock3 & v1446111;
assign v845578 = hgrant3_p & v845542 | !hgrant3_p & !v845542;
assign v138949a = hgrant3_p & v138945b | !hgrant3_p & v1389499;
assign v1389fbc = hmaster2_p & f2f4b0 | !hmaster2_p & v845542;
assign d2face = hmaster1_p & d2facd | !hmaster1_p & d2fe8c;
assign v1214e0c = hgrant1_p & v1214e0b | !hgrant1_p & v1216aeb;
assign d30672 = hlock5_p & v845542 | !hlock5_p & v1668c1d;
assign v1445f25 = hmaster1_p & v1445f21 | !hmaster1_p & v845542;
assign v134d4b9 = hbusreq5 & v134d4b7 | !hbusreq5 & v134d4b8;
assign v1389d5b = hmaster0_p & v1389d5a | !hmaster0_p & !v845542;
assign v1445a1c = hgrant5_p & v14458f9 | !hgrant5_p & v1445a1b;
assign f2f2f0 = hmaster1_p & f2f2ef | !hmaster1_p & f2f2db;
assign v1445458 = hbusreq2_p & v1445457 | !hbusreq2_p & v1445bb3;
assign v144538d = hmaster1_p & v144535f | !hmaster1_p & v144591b;
assign v12166c3 = hgrant0_p & v12164cf | !hgrant0_p & !v845542;
assign v1552d8c = hmaster2_p & v1552d86 | !hmaster2_p & v1552d8b;
assign v10d4014 = hmaster0_p & v10d3fdc | !hmaster0_p & v10d3fda;
assign v10d42e0 = hbusreq3_p & v10d42bf | !hbusreq3_p & !v10d42df;
assign v1515720 = locked_p & v151571b | !locked_p & v151571f;
assign v1515835 = hgrant5_p & v10d3ffd | !hgrant5_p & v1515833;
assign v949cd9 = hmaster2_p & v845542 | !hmaster2_p & !v845558;
assign a6566a = hbusreq5_p & a65440 | !hbusreq5_p & !a65669;
assign d30764 = hbusreq2 & d30760 | !hbusreq2 & d30763;
assign a65382 = hgrant0_p & a6537d | !hgrant0_p & v845570;
assign v1668c65 = hmaster2_p & a658b5 | !hmaster2_p & v1668c64;
assign v121571d = hlock0_p & v1216523 | !hlock0_p & !v845542;
assign v1553399 = hbusreq4 & v155338b | !hbusreq4 & v1553217;
assign v144547f = hmaster0_p & v144547e | !hmaster0_p & v1446404;
assign v121659b = hgrant4_p & v121659a | !hgrant4_p & v1216a96;
assign v144631c = hlock0 & v144631b | !hlock0 & v144631a;
assign d30751 = hmaster2_p & d30734 | !hmaster2_p & v84554e;
assign v1445f5b = hmaster1_p & v1445f5a | !hmaster1_p & v1446436;
assign v10d42bf = hgrant3_p & v10d4013 | !hgrant3_p & v10d42be;
assign v121573a = hbusreq4_p & v1215739 | !hbusreq4_p & v845542;
assign v1445a2b = hlock1 & v1445a17 | !hlock1 & v1445a2a;
assign v1445753 = hbusreq2 & v1445f4e | !hbusreq2 & v1445f4f;
assign v11e5960 = hbusreq2_p & v11e595e | !hbusreq2_p & v11e595f;
assign d80744 = hlock0_p & d80732 | !hlock0_p & !v845542;
assign v1215fb3 = hmaster0_p & v12166f7 | !hmaster0_p & v12166c8;
assign v12162e3 = hbusreq3_p & v121626c | !hbusreq3_p & !v12162e2;
assign v1405911 = hbusreq0_p & v1405860 | !hbusreq0_p & !v144639c;
assign v138a480 = hgrant2_p & v138a47e | !hgrant2_p & !v138a47f;
assign v138a3cd = hgrant5_p & v845570 | !hgrant5_p & !v138a3cc;
assign v151575c = hgrant5_p & v151574c | !hgrant5_p & !v151575b;
assign v1216080 = hlock5_p & v121607e | !hlock5_p & v121607f;
assign v1216aa2 = busreq_p & v845542 | !busreq_p & v144646d;
assign f2f2a1 = hmaster2_p & f2f29e | !hmaster2_p & f2f2a0;
assign v1445830 = hgrant2_p & v144582e | !hgrant2_p & v144582f;
assign v1215bb5 = hmaster1_p & v1215bb4 | !hmaster1_p & !v12163a9;
assign v1445fb0 = hmaster0_p & v144639c | !hmaster0_p & v1445f85;
assign v12161f4 = hmaster0_p & v12161dd | !hmaster0_p & v12161f3;
assign v138a002 = hbusreq5_p & v138a001 | !hbusreq5_p & !v845542;
assign v1445a27 = hlock0_p & v144641b | !hlock0_p & v1445a26;
assign d307e6 = hbusreq0_p & a653d9 | !hbusreq0_p & v845542;
assign v1668dda = hgrant5_p & v845570 | !hgrant5_p & v1668d9d;
assign v10d40bf = hgrant4_p & v10d401a | !hgrant4_p & v10d40be;
assign v16a1dc1 = hmaster1_p & v845568 | !hmaster1_p & v16a2672;
assign v16a19dd = hbusreq2_p & v16a1841 | !hbusreq2_p & v16a19d4;
assign v16a223c = hgrant4_p & v845542 | !hgrant4_p & v16a223b;
assign v16a1d9b = hgrant2_p & v16a2060 | !hgrant2_p & v16a1d9a;
assign v14058d6 = hmaster2_p & v14058d0 | !hmaster2_p & v14058d5;
assign v1445b7f = hbusreq2_p & v1445b7c | !hbusreq2_p & v1445b7e;
assign d80756 = stateG2_p & v845542 | !stateG2_p & !d80755;
assign v1515baf = hready_p & v1515aef | !hready_p & !v1515bae;
assign v16a1a95 = hmaster1_p & v16a1a94 | !hmaster1_p & !v16a2672;
assign d300d0 = hgrant5_p & d2fe9b | !hgrant5_p & !d300ce;
assign d3088c = hgrant5_p & d3084f | !hgrant5_p & !d3088b;
assign v1668de4 = hbusreq2_p & v1668de2 | !hbusreq2_p & !v1668de3;
assign v1445811 = hgrant2_p & v144580f | !hgrant2_p & v1445810;
assign v134d4ff = hgrant1_p & v845542 | !hgrant1_p & v134d4fe;
assign v1405b29 = hmaster0_p & v1405b21 | !hmaster0_p & !v1405b28;
assign v1215bfd = hmaster2_p & v1215bf1 | !hmaster2_p & v121652e;
assign v16a1ded = hmaster1_p & v16a2243 | !hmaster1_p & !v16a2672;
assign v1515714 = hbusreq4 & v10d3fd4 | !hbusreq4 & !v845542;
assign v140587a = hbusreq2_p & v1405879 | !hbusreq2_p & v1405878;
assign bf1f52 = locked_p & v845542 | !locked_p & !v84556a;
assign v16a2672 = hmaster0_p & v16a266b | !hmaster0_p & v16a2671;
assign d2fe82 = hmaster0_p & d2fe7e | !hmaster0_p & d2fe81;
assign v1405af5 = hmaster1_p & v1405af4 | !hmaster1_p & !v1405a94;
assign v1216266 = hbusreq2_p & v1216260 | !hbusreq2_p & v1216265;
assign v1215d34 = hgrant5_p & v1215d32 | !hgrant5_p & v1215d33;
assign v12161f9 = hmaster1_p & v12161f8 | !hmaster1_p & v1216041;
assign v134d469 = decide_p & v134d3ce | !decide_p & v134d45b;
assign v1445a01 = hbusreq1 & v14459f8 | !hbusreq1 & v1445a00;
assign v1214c45 = hbusreq1 & v1215345 | !hbusreq1 & v845542;
assign v10d407a = hmaster2_p & v10d4074 | !hmaster2_p & v10d4079;
assign v14460c6 = hbusreq2 & v14460c1 | !hbusreq2 & v14460c5;
assign v16a1d2e = hmaster1_p & v16a1d2d | !hmaster1_p & !v16a2672;
assign v16a1d78 = hbusreq0 & v16a209a | !hbusreq0 & v16a1d77;
assign v15157f6 = hgrant5_p & v845542 | !hgrant5_p & !v1515781;
assign v16a1384 = hmaster1_p & v16a1383 | !hmaster1_p & !v16a2672;
assign v1215376 = hmastlock_p & v1215375 | !hmastlock_p & v845542;
assign d3065c = hgrant4_p & a66284 | !hgrant4_p & d3065b;
assign v144579b = hmaster2_p & v1445de5 | !hmaster2_p & v1445edc;
assign d2fee5 = hmaster0_p & d2fee4 | !hmaster0_p & d2fec5;
assign v1446099 = hmaster0_p & v1446053 | !hmaster0_p & v1446066;
assign d3064d = hbusreq5_p & d3064c | !hbusreq5_p & v845542;
assign v1284d16 = hgrant5_p & v1284d0f | !hgrant5_p & v1284d15;
assign v1214ed3 = hmaster2_p & v1216536 | !hmaster2_p & v845542;
assign v12aeb77 = hmaster0_p & v845542 | !hmaster0_p & v12aeb76;
assign d30136 = hbusreq5_p & d30135 | !hbusreq5_p & d30134;
assign v1446663 = hlock0 & v1446662 | !hlock0 & v1446661;
assign d30275 = hmaster2_p & d3064a | !hmaster2_p & d30651;
assign v144577a = hmaster1_p & v1445779 | !hmaster1_p & v1445e07;
assign v1215000 = hgrant5_p & v1214ffa | !hgrant5_p & !v1214fff;
assign d307b5 = hlock1_p & d307b4 | !hlock1_p & d30649;
assign v12150c4 = hbusreq4_p & v12150c3 | !hbusreq4_p & v845542;
assign v1405876 = hmaster0_p & v1405871 | !hmaster0_p & v1405861;
assign v134d433 = hmaster1_p & v134d369 | !hmaster1_p & v134d432;
assign v1445a8e = hmaster1_p & v1445a6c | !hmaster1_p & v144591b;
assign f2f295 = hbusreq1_p & f2f294 | !hbusreq1_p & v845542;
assign v134d4e5 = hlock4 & v134d36d | !hlock4 & v134d273;
assign v14460dc = hbusreq2 & v14460d8 | !hbusreq2 & v14460db;
assign v155339c = hgrant4_p & v1553217 | !hgrant4_p & v845542;
assign v1214eef = hbusreq5_p & v1214eee | !hbusreq5_p & v1216531;
assign v16a13d3 = hmaster1_p & v16a13c7 | !hmaster1_p & v16a1f96;
assign v134d1fd = hmaster2_p & v845542 | !hmaster2_p & v134d1fc;
assign v14457ad = hbusreq3 & v144579a | !hbusreq3 & v14457ac;
assign v14465e2 = hmaster2_p & v14465b3 | !hmaster2_p & v14465e1;
assign v1284c99 = hlock1_p & v1284c8e | !hlock1_p & !v14463b1;
assign d8079c = hmaster0_p & d80791 | !hmaster0_p & !d8079b;
assign d3078f = hgrant4_p & a66284 | !hgrant4_p & d3078e;
assign v144583b = hgrant2_p & v144583a | !hgrant2_p & v1445836;
assign v1215781 = hgrant2_p & v1215775 | !hgrant2_p & !v1215780;
assign d807a3 = hbusreq2_p & d8079e | !hbusreq2_p & d807a2;
assign v144625c = hlock3 & v1446224 | !hlock3 & v144625b;
assign a6566c = hgrant5_p & a65424 | !hgrant5_p & !a65638;
assign v16a1cea = hbusreq1_p & v16a1bbc | !hbusreq1_p & v16a1ad9;
assign v1405b58 = hgrant2_p & v1405b3e | !hgrant2_p & v1405b57;
assign d300f1 = hlock5_p & d300ef | !hlock5_p & d300f0;
assign v134d1f3 = hmaster2_p & v134d1e8 | !hmaster2_p & v134d1f2;
assign v1515819 = hmaster2_p & v151564d | !hmaster2_p & !a658c6;
assign v138a47a = hmaster0_p & v138a3ec | !hmaster0_p & v138a3cb;
assign a65391 = hbusreq1 & a6585d | !hbusreq1 & a6588f;
assign v15157a5 = hmaster0_p & v15157a0 | !hmaster0_p & v15157a4;
assign d30654 = hbusreq1_p & v84554e | !hbusreq1_p & !v845542;
assign a65655 = hgrant2_p & a6561c | !hgrant2_p & a65653;
assign v12150ac = hmaster1_p & v12150ab | !hmaster1_p & !v12150a6;
assign v144661f = hbusreq1 & v144661d | !hbusreq1 & v144661e;
assign v1405af2 = hgrant2_p & v1405ad2 | !hgrant2_p & v1405af1;
assign v121572c = hmaster2_p & v121572a | !hmaster2_p & v121572b;
assign v134d49a = hmaster0_p & v134d496 | !hmaster0_p & v134d499;
assign v1445ea6 = hmaster2_p & v1446609 | !hmaster2_p & v1445ea5;
assign v14466f5 = hmaster0_p & v144663a | !hmaster0_p & v1446448;
assign v16a1cba = hbusreq3 & v16a1ca3 | !hbusreq3 & v16a1cb9;
assign v1445ad5 = hlock2 & v1445abf | !hlock2 & v1445ad3;
assign v138a446 = hbusreq2_p & v138a442 | !hbusreq2_p & v138a445;
assign d807ab = hgrant5_p & d80762 | !hgrant5_p & d807aa;
assign d300df = hgrant1_p & d300da | !hgrant1_p & d300de;
assign v1668d84 = hgrant4_p & v1668d7a | !hgrant4_p & a653dd;
assign v1445389 = hgrant2_p & v1445388 | !hgrant2_p & v1445384;
assign v1445d8c = hgrant5_p & v1445d89 | !hgrant5_p & !v1445d8b;
assign v1446216 = hlock0 & v1446215 | !hlock0 & v1446210;
assign v12164e6 = hbusreq2_p & v12164e2 | !hbusreq2_p & v12164e5;
assign v1216af5 = hlock5_p & v1216aef | !hlock5_p & v1216af4;
assign v121625c = hgrant1_p & v1216204 | !hgrant1_p & v121625b;
assign v1216555 = hgrant1_p & v1216522 | !hgrant1_p & v1216554;
assign v16a1844 = hmaster1_p & v16a1843 | !hmaster1_p & v16a2672;
assign v144551d = hgrant2_p & v14454e9 | !hgrant2_p & v144551c;
assign v1215024 = hmaster1_p & v1215023 | !hmaster1_p & v121546f;
assign v12161da = hgrant1_p & v845542 | !hgrant1_p & f2f2a8;
assign d301da = hgrant5_p & v845580 | !hgrant5_p & !d301d8;
assign v12ad668 = hbusreq2_p & v12ad65f | !hbusreq2_p & v12ad667;
assign d306b0 = hgrant1_p & v84554c | !hgrant1_p & d306af;
assign v10d3fdd = hmaster0_p & v10d3fda | !hmaster0_p & v10d3fdc;
assign v14458c4 = hbusreq2_p & v14458c2 | !hbusreq2_p & v14458c3;
assign v16a1d60 = hgrant5_p & v845542 | !hgrant5_p & !v16a1d48;
assign v1553233 = hgrant0_p & v1553232 | !hgrant0_p & v845542;
assign d2fbce = hbusreq4_p & d2fbcd | !hbusreq4_p & v84554a;
assign v1553226 = hlock1_p & v1553138 | !hlock1_p & v845542;
assign v1405b0d = hgrant2_p & v1405ad1 | !hgrant2_p & v1405b0c;
assign v11e596e = decide_p & v11e5960 | !decide_p & v11e596d;
assign v134d1f6 = hbusreq1 & v134d1e8 | !hbusreq1 & v134d1f5;
assign d2f9aa = hmaster1_p & d2f99c | !hmaster1_p & d2f9a9;
assign v14459a5 = stateA1_p & v845588 | !stateA1_p & !v845542;
assign v1445bf2 = hbusreq2_p & v1445bef | !hbusreq2_p & v1445bf1;
assign v12165a7 = hgrant2_p & v1216585 | !hgrant2_p & v12165a6;
assign v144553d = hbusreq3_p & v144543e | !hbusreq3_p & v144553c;
assign v134d394 = hgrant1_p & v845542 | !hgrant1_p & v134d393;
assign v1552d68 = hbusreq3 & v1552d67 | !hbusreq3 & v155341e;
assign v12160de = hbusreq1_p & v12160dd | !hbusreq1_p & v845542;
assign a656c4 = hready_p & a656c3 | !hready_p & a65b20;
assign v1553440 = hbusreq5_p & v1553224 | !hbusreq5_p & v155343f;
assign v1515759 = hgrant5_p & v151573d | !hgrant5_p & v1515758;
assign v138a453 = hmaster0_p & v138a344 | !hmaster0_p & v138a354;
assign d2fd4a = hready_p & d2fd49 | !hready_p & d2fd42;
assign v12160c7 = hmaster0_p & v1216099 | !hmaster0_p & v1216093;
assign d2fc38 = hmaster2_p & d2fc37 | !hmaster2_p & d30690;
assign v11e594a = hlock1_p & v11e593a | !hlock1_p & v845570;
assign d30645 = locked_p & d30644 | !locked_p & v845542;
assign v1445774 = hbusreq5 & v1445772 | !hbusreq5 & v1445773;
assign v1445ef3 = hmaster1_p & v1445eb1 | !hmaster1_p & v1445e28;
assign v1215c26 = hgrant1_p & v1215c25 | !hgrant1_p & v1216139;
assign v14460f3 = hlock2 & v14460f2 | !hlock2 & v14460ed;
assign v134d4c8 = stateA1_p & v134d1db | !stateA1_p & v134d1da;
assign v121509c = hmaster2_p & v121509b | !hmaster2_p & v1215098;
assign v1445778 = hlock0 & v1445777 | !hlock0 & v1445775;
assign d8077a = hbusreq4_p & d80779 | !hbusreq4_p & !v845542;
assign v144535e = hbusreq2 & v1445b44 | !hbusreq2 & v144535d;
assign v1445f01 = hlock3 & v1445edb | !hlock3 & v1445f00;
assign v14465b7 = hgrant5_p & v1446404 | !hgrant5_p & v14465b6;
assign a656a5 = hmaster1_p & a65493 | !hmaster1_p & !a65916;
assign v1215037 = hbusreq4_p & v1215036 | !hbusreq4_p & v845542;
assign v14458c6 = hbusreq2_p & v14458c2 | !hbusreq2_p & v14458c5;
assign v144584f = hgrant2_p & v1445829 | !hgrant2_p & v1445848;
assign v12ad5b7 = hbusreq1 & v12ad4cc | !hbusreq1 & !v12ad4e6;
assign v14058bb = hbusreq5_p & v14058ba | !hbusreq5_p & v14058b9;
assign v1215c92 = hmaster2_p & v845570 | !hmaster2_p & v1216a5a;
assign v16a224f = hgrant2_p & v16a205c | !hgrant2_p & v16a224e;
assign v16a1e60 = hmaster1_p & v16a1e5f | !hmaster1_p & v16a2672;
assign v16a207f = hgrant4_p & v845559 | !hgrant4_p & !v845572;
assign v144580c = hgrant2_p & v1445809 | !hgrant2_p & v144580b;
assign v1446092 = hlock0 & v1446091 | !hlock0 & v1446090;
assign v13897ef = hmaster0_p & v13897e0 | !hmaster0_p & v1389de1;
assign a65399 = hbusreq4_p & a65396 | !hbusreq4_p & !v845542;
assign v1215ce9 = hgrant5_p & v845542 | !hgrant5_p & v1215c9a;
assign d2fea3 = hmaster1_p & d2fe9b | !hmaster1_p & !d2fea2;
assign d30608 = hmaster0_p & d305f7 | !hmaster0_p & d30607;
assign v16a1d99 = hgrant2_p & v16a205f | !hgrant2_p & v16a1d98;
assign v1515731 = hbusreq5_p & v151572f | !hbusreq5_p & v1515730;
assign v12ad581 = hbusreq2_p & v12ad550 | !hbusreq2_p & v12ad580;
assign v121509d = hgrant5_p & v121503d | !hgrant5_p & !v121509c;
assign v12166ff = hmaster1_p & v12166fe | !hmaster1_p & v12164e1;
assign d3081e = hmaster2_p & d3080a | !hmaster2_p & v845542;
assign v1445eb8 = hgrant5_p & v1445eb6 | !hgrant5_p & v1445eb7;
assign d2fec9 = hmaster0_p & d2feb5 | !hmaster0_p & d2fec8;
assign v1215c68 = hgrant5_p & v845542 | !hgrant5_p & v1215c30;
assign v1284cfc = hgrant5_p & v140584c | !hgrant5_p & v1284cfb;
assign v151581c = hlock2_p & v151581b | !hlock2_p & !v15156f6;
assign v1668cd7 = hmaster1_p & v1668cbf | !hmaster1_p & v1668cd6;
assign v84554a = hlock0_p & v845542 | !hlock0_p & !v845542;
assign v1215776 = hmaster2_p & v1215717 | !hmaster2_p & v1215747;
assign f2e714 = hmaster2_p & f2f228 | !hmaster2_p & f2e713;
assign v1389d76 = hbusreq5 & v1389d5c | !hbusreq5 & v1389d75;
assign v15156f4 = hmaster2_p & v1515675 | !hmaster2_p & v845542;
assign a65623 = hgrant1_p & a653ae | !hgrant1_p & !a65622;
assign v12ad8e8 = hbusreq1_p & v12add48 | !hbusreq1_p & v12ad8e7;
assign v1215c5e = hlock5_p & v1215c5c | !hlock5_p & v1215c5d;
assign v15156ff = hbusreq2 & v15156fe | !hbusreq2 & v15167ed;
assign v1446344 = hmaster1_p & v1446313 | !hmaster1_p & v1446341;
assign v134d310 = hgrant4_p & v845542 | !hgrant4_p & v134d30f;
assign a6470e = hbusreq2_p & a6470d | !hbusreq2_p & a65b2c;
assign v134d313 = hgrant5_p & v845542 | !hgrant5_p & v134d312;
assign v14460b0 = hmaster2_p & v144608e | !hmaster2_p & v14465db;
assign v1515747 = hgrant4_p & v1515746 | !hgrant4_p & v151560d;
assign v1515757 = hgrant1_p & v1515743 | !hgrant1_p & v1515756;
assign v16a1bc7 = hgrant0_p & v845542 | !hgrant0_p & !v16a1bc6;
assign v14463bb = hlock0_p & v144639c | !hlock0_p & !v14463ba;
assign v16a19b6 = hmaster1_p & v16a19b5 | !hmaster1_p & !v16a2672;
assign v1552d8d = hgrant5_p & v845542 | !hgrant5_p & v1552d8c;
assign v144614c = hmaster1_p & v144612d | !hmaster1_p & v1445ffc;
assign v138945a = decide_p & v1389459 | !decide_p & v845542;
assign f2f538 = hmaster2_p & f2f228 | !hmaster2_p & f2f22a;
assign f2f2e5 = hmaster1_p & f2f2e4 | !hmaster1_p & f2f2db;
assign d30297 = hbusreq2_p & d30295 | !hbusreq2_p & !d30296;
assign v1214d9f = hmaster1_p & v1214d9e | !hmaster1_p & v1214cd8;
assign v1216145 = hlock0_p & v1216523 | !hlock0_p & v1216144;
assign v1214d58 = hmaster1_p & v1214d50 | !hmaster1_p & v1214d4b;
assign v134d28c = hgrant4_p & v134d28b | !hgrant4_p & v845542;
assign v85e755 = hbusreq3_p & a7c7c1 | !hbusreq3_p & !v845542;
assign d3014e = hmaster0_p & d30144 | !hmaster0_p & d3014d;
assign v121631d = hmaster1_p & v12162f7 | !hmaster1_p & v121631b;
assign f2f42b = hmaster2_p & f2f423 | !hmaster2_p & f2f286;
assign v16a16b7 = jx1_p & v16a1d05 | !jx1_p & v16a16b6;
assign v12152e9 = hmaster0_p & v121577e | !hmaster0_p & v1215730;
assign v121629a = hbusreq5_p & v12161aa | !hbusreq5_p & v1216299;
assign v16a208b = hgrant5_p & v845542 | !hgrant5_p & v16a208a;
assign d3083f = hbusreq2_p & d30832 | !hbusreq2_p & !d3083e;
assign v16695a6 = decide_p & v16695a3 | !decide_p & v845542;
assign v134d260 = hbusreq2_p & v134d245 | !hbusreq2_p & v134d244;
assign v1214e57 = hbusreq1_p & v1216ab8 | !hbusreq1_p & v1216ab9;
assign d3076b = hbusreq2_p & d3076a | !hbusreq2_p & d30769;
assign v1215056 = hgrant2_p & v1215024 | !hgrant2_p & v1215055;
assign v12ad5e2 = hmaster1_p & v12ad5b5 | !hmaster1_p & v12ad5e1;
assign v144639c = hmastlock_p & v146d169 | !hmastlock_p & v845542;
assign v1215bd4 = hbusreq5 & v1215bbb | !hbusreq5 & v1215bd3;
assign v1216027 = hmaster0_p & v1216020 | !hmaster0_p & v1216026;
assign v1215d74 = hgrant5_p & v1215d72 | !hgrant5_p & !v1215d73;
assign v16a1e03 = hbusreq5 & v16a1dfe | !hbusreq5 & v16a1e02;
assign v1216ad2 = hmastlock_p & v1446395 | !hmastlock_p & v845542;
assign v1214f60 = hbusreq2_p & v1214f5f | !hbusreq2_p & v12164e7;
assign v1214eeb = hbusreq0 & v1214ee7 | !hbusreq0 & v1214eea;
assign v1515641 = hmaster1_p & v1515640 | !hmaster1_p & v845542;
assign d2feba = hbusreq1_p & d2feb9 | !hbusreq1_p & v84555a;
assign v1216594 = hready & v1216590 | !hready & v1216593;
assign v1445dfc = hbusreq4_p & v1446423 | !hbusreq4_p & v1446429;
assign v1214cc2 = hmaster2_p & v1215379 | !hmaster2_p & v1215380;
assign f2f3b1 = hbusreq1_p & f2f3b0 | !hbusreq1_p & !v845542;
assign d3010e = hmaster0_p & d300f6 | !hmaster0_p & d3010d;
assign d2fbc5 = hready_p & d2fb5f | !hready_p & d2fbc4;
assign v1668d2b = hmaster2_p & v10d3fd8 | !hmaster2_p & v845542;
assign v1668c30 = hmaster0_p & v1668c2f | !hmaster0_p & v845542;
assign v134d4a1 = hmaster0_p & v845542 | !hmaster0_p & v134d4a0;
assign d2fb55 = hmaster0_p & d2fb51 | !hmaster0_p & d2fb54;
assign v134d23c = hmaster0_p & v134d23b | !hmaster0_p & v134d207;
assign v14463fd = hlock2 & v14463d1 | !hlock2 & v14463fb;
assign v15157af = hmaster2_p & v151579b | !hmaster2_p & v15157ae;
assign v15157db = hgrant5_p & v845542 | !hgrant5_p & !v151572e;
assign d30201 = hbusreq5_p & d301fd | !hbusreq5_p & d30200;
assign d3072d = hmaster1_p & d3071e | !hmaster1_p & d3072c;
assign v1445f1f = hready_p & v1445e52 | !hready_p & v1445f1e;
assign v1668d61 = hbusreq0 & v1668d57 | !hbusreq0 & v1668d60;
assign v1216a73 = hready & v1216a60 | !hready & !d305dd;
assign d3060f = hlock2_p & d30609 | !hlock2_p & d3060e;
assign v1668c45 = hmaster1_p & v1668c42 | !hmaster1_p & v1668c44;
assign v1214d3b = hmaster0_p & v1214cdc | !hmaster0_p & v121537e;
assign v1284ce3 = hgrant5_p & v1405859 | !hgrant5_p & v1284ce2;
assign v1214eba = hmaster1_p & v1214eb5 | !hmaster1_p & v1214e73;
assign v1445901 = hbusreq0 & v14458ff | !hbusreq0 & v1445900;
assign v12ad65d = hbusreq2_p & v12ad632 | !hbusreq2_p & v12ad65c;
assign v144641b = hbusreq4 & v144641a | !hbusreq4 & v144640b;
assign v134ce3e = hbusreq4_p & v134d273 | !hbusreq4_p & v134ce3d;
assign d2fe7c = hlock4_p & v845542 | !hlock4_p & a66295;
assign v1445500 = hlock2 & v14454fa | !hlock2 & v14454ff;
assign v144548c = hbusreq2 & v1445481 | !hbusreq2 & v1445482;
assign v134cdc3 = hmaster1_p & v134cdc2 | !hmaster1_p & v845542;
assign v1445f92 = hbusreq1 & v14463ab | !hbusreq1 & v14463e3;
assign v1668c1f = hbusreq5_p & v845570 | !hbusreq5_p & v845542;
assign v1445b43 = hbusreq2_p & v1445b35 | !hbusreq2_p & v1445b42;
assign v1446312 = hlock0 & v1446311 | !hlock0 & v144630b;
assign v1214d15 = hmaster0_p & v1214c2e | !hmaster0_p & v1214d14;
assign v1445879 = hbusreq1_p & v144639c | !hbusreq1_p & v144586f;
assign f2f358 = hgrant1_p & v845570 | !hgrant1_p & !f2f357;
assign v1446104 = hbusreq2_p & v1446102 | !hbusreq2_p & v1446103;
assign d2fbc8 = hmaster1_p & d2fbc7 | !hmaster1_p & d2fb55;
assign a646db = decide_p & a646da | !decide_p & v845542;
assign v134d212 = hlock2_p & v134d210 | !hlock2_p & v134d211;
assign v1445899 = hbusreq4_p & v144639c | !hbusreq4_p & v1445898;
assign d80783 = hmaster0_p & d80778 | !hmaster0_p & !d80782;
assign v1216524 = hbusreq4_p & v1216523 | !hbusreq4_p & v16a19a4;
assign d2fbda = hbusreq5_p & d2fbd9 | !hbusreq5_p & d2fbd8;
assign v1445f83 = hgrant3_p & v1446724 | !hgrant3_p & v1445f82;
assign v1668c29 = hmaster2_p & v845542 | !hmaster2_p & !v84556a;
assign v1405a80 = hmaster1_p & v1405a7d | !hmaster1_p & v1405a7f;
assign v9dde65 = hmaster2_p & v84554c | !hmaster2_p & !v845542;
assign v134d3d4 = hlock3 & v134d276 | !hlock3 & v134d3d3;
assign v12add46 = hlock0_p & v1515c7e | !hlock0_p & v845542;
assign v1405a9e = hlock3_p & v1405a99 | !hlock3_p & v1405a9d;
assign v14458a7 = hmaster0_p & v144639c | !hmaster0_p & v14458a6;
assign v1445f4c = hmaster1_p & v1445db8 | !hmaster1_p & v1445da4;
assign v16a13e0 = hmaster1_p & v16a13df | !hmaster1_p & v16a1d6d;
assign a65aed = hmaster2_p & a65aeb | !hmaster2_p & a65ae4;
assign v12ad59f = stateG2_p & v845542 | !stateG2_p & !v10d4264;
assign v12acfdd = hbusreq2_p & v12acfd7 | !hbusreq2_p & v12acfdc;
assign v16a141a = hbusreq3 & v16a1415 | !hbusreq3 & v16a1419;
assign v12ad4c8 = hgrant3_p & v12ad953 | !hgrant3_p & v12ad4c7;
assign v10d42b7 = hmaster2_p & v10d42b2 | !hmaster2_p & !v10d406d;
assign v1214d63 = hbusreq2_p & v1214c18 | !hbusreq2_p & v1214d62;
assign v144667f = hlock0 & v144667e | !hlock0 & v144667d;
assign v12ad602 = hbusreq0 & v12ad601 | !hbusreq0 & v12afe63;
assign v1215c9f = hmaster0_p & v1215c91 | !hmaster0_p & v1215c9e;
assign v16a18dd = decide_p & v16a1890 | !decide_p & !v16a2065;
assign v1216210 = hbusreq1 & v12166c4 | !hbusreq1 & v845542;
assign v1668d02 = hmaster1_p & v1668cd9 | !hmaster1_p & !v1668d01;
assign d2fb74 = hbusreq5_p & d2fb73 | !hbusreq5_p & d2fb72;
assign d80794 = hgrant1_p & v845542 | !hgrant1_p & !d80793;
assign bf1fa4 = hmaster0_p & bf1f98 | !hmaster0_p & bf1fa3;
assign v15155ef = decide_p & v15155ee | !decide_p & v845542;
assign v14457f3 = hmaster1_p & v14457f2 | !hmaster1_p & v1445e1b;
assign v1215412 = hlock2_p & v1215410 | !hlock2_p & v1215411;
assign v1445e09 = hmaster2_p & v1445de5 | !hmaster2_p & v1445df2;
assign v144617b = hbusreq2_p & v1446176 | !hbusreq2_p & v144617a;
assign v144642f = hbusreq0_p & v1446403 | !hbusreq0_p & v144640c;
assign v1215cee = hgrant5_p & v1215ced | !hgrant5_p & v1215ca6;
assign a65365 = stateG2_p & v845542 | !stateG2_p & a65364;
assign v12aeb1f = hmaster1_p & v845542 | !hmaster1_p & v12aeb1e;
assign v1515c88 = hready_p & v845542 | !hready_p & v1515c87;
assign a65634 = hbusreq5_p & a653fe | !hbusreq5_p & a65632;
assign f2f3d7 = hbusreq5_p & f2f3d5 | !hbusreq5_p & !f2f3d6;
assign f2f36a = hmaster2_p & f2f369 | !hmaster2_p & f2f234;
assign v10d42c8 = hbusreq1_p & v10d426a | !hbusreq1_p & v10d42c7;
assign v1446564 = hgrant2_p & v1446461 | !hgrant2_p & v1446563;
assign v138944f = hmaster1_p & v845542 | !hmaster1_p & v138944e;
assign v14460eb = hmaster0_p & v1445fa2 | !hmaster0_p & v1445fa9;
assign v1445ac6 = hbusreq2_p & v1445ac3 | !hbusreq2_p & v1445ac5;
assign v1445b25 = hlock2 & v1445af2 | !hlock2 & v1445b23;
assign f2f40d = hbusreq2_p & f2f40b | !hbusreq2_p & f2f40c;
assign v12ad27a = hready_p & v12ad22e | !hready_p & v12ad279;
assign d2f9a7 = hbusreq5_p & d2f993 | !hbusreq5_p & d2f9a6;
assign v144542a = hbusreq2_p & v1445429 | !hbusreq2_p & v144541b;
assign v1405b15 = hmaster2_p & v1405b14 | !hmaster2_p & !v845542;
assign f2f3da = hmaster1_p & f2f3d9 | !hmaster1_p & f2f3cf;
assign d807b6 = hmaster0_p & d8079f | !hmaster0_p & v845542;
assign v1215063 = hmaster1_p & v1215062 | !hmaster1_p & v121546f;
assign v1445a14 = hgrant4_p & v1445a0d | !hgrant4_p & v1445a13;
assign v121615d = hgrant4_p & v121613d | !hgrant4_p & v845542;
assign v1215cdf = hbusreq2 & v1215cd8 | !hbusreq2 & v1215cde;
assign f2f3d0 = hmaster1_p & f2f3be | !hmaster1_p & f2f3cf;
assign v10d4076 = hlock0_p & v10d3fd9 | !hlock0_p & v10d4075;
assign d2fc82 = jx2_p & d2fb4b | !jx2_p & d2fc81;
assign v12153e0 = hbusreq5_p & v12153df | !hbusreq5_p & v12153de;
assign v1446717 = hmaster0_p & v144667f | !hmaster0_p & v1446448;
assign v14459e2 = hgrant5_p & v14459d4 | !hgrant5_p & v14459e1;
assign v134d52a = hbusreq5 & v134d528 | !hbusreq5 & v134d529;
assign v16a1cdd = hbusreq2_p & v16a1b64 | !hbusreq2_p & v16a1cdc;
assign v1389498 = decide_p & v1389459 | !decide_p & v138a406;
assign v14453ae = hgrant2_p & v1445388 | !hgrant2_p & v14453aa;
assign f2f22c = hbusreq5_p & f2f229 | !hbusreq5_p & f2f22b;
assign v11f33c5 = jx2_p & v85e75f | !jx2_p & !v85e749;
assign v121618e = hbusreq0 & v121618c | !hbusreq0 & v121618d;
assign a65445 = hmaster0_p & a6541e | !hmaster0_p & a65444;
assign v1215748 = hmaster2_p & v1215747 | !hmaster2_p & v121573d;
assign v1515764 = hbusreq4 & v1515741 | !hbusreq4 & a65396;
assign v1216583 = hbusreq5 & v1216582 | !hbusreq5 & v845542;
assign v1445521 = hgrant2_p & v144551f | !hgrant2_p & v1445520;
assign v14461b8 = hmaster1_p & v144616b | !hmaster1_p & v1445ffc;
assign v121655c = hbusreq4 & v1216a67 | !hbusreq4 & v1216a77;
assign f2f397 = hmaster0_p & f2f350 | !hmaster0_p & f2f396;
assign v1668d3c = hgrant1_p & v1668d23 | !hgrant1_p & v1668d3b;
assign v1214d74 = hmaster0_p & v1215359 | !hmaster0_p & v1215349;
assign v14465ec = hbusreq4 & v14465eb | !hbusreq4 & v14465c3;
assign v16a2095 = hmaster0_p & v16a2091 | !hmaster0_p & v16a2094;
assign v1446407 = locked_p & v845542 | !locked_p & v144639c;
assign v1553518 = decide_p & v155342e | !decide_p & v155350a;
assign v144624a = hmaster2_p & v14463a2 | !hmaster2_p & v14463db;
assign a65b07 = hready_p & v845542 | !hready_p & a65b06;
assign v12164d4 = hmaster2_p & v12164cf | !hmaster2_p & v12164d3;
assign v12161d5 = hmaster2_p & v12161d1 | !hmaster2_p & v845542;
assign v12ad01f = hbusreq2_p & v12ad01b | !hbusreq2_p & !v12ad01e;
assign v1445af8 = hmaster1_p & v1445af7 | !hmaster1_p & v14458fd;
assign v12160f7 = hbusreq1_p & v12160f6 | !hbusreq1_p & v845542;
assign v1216ab8 = hready & v1446397 | !hready & !d305ee;
assign v1516999 = hmaster0_p & v845542 | !hmaster0_p & v1516998;
assign v1215c6a = hmaster0_p & v1215c66 | !hmaster0_p & v1215c69;
assign v134d4b6 = hbusreq3 & v134d4b5 | !hbusreq3 & v134d3b5;
assign v1446639 = hbusreq0 & v1446637 | !hbusreq0 & v1446638;
assign v16a1e26 = hmaster2_p & v16a1e21 | !hmaster2_p & v845542;
assign v138a355 = hmaster0_p & v138a32d | !hmaster0_p & v138a354;
assign v1214d3f = hbusreq2_p & v1214d3c | !hbusreq2_p & v1214d3e;
assign v14459c6 = hlock0_p & v14459c4 | !hlock0_p & v14459c5;
assign v11e5977 = hgrant4_p & v845542 | !hgrant4_p & v11e5976;
assign d307c5 = hlock4_p & v845542 | !hlock4_p & d307c4;
assign v1445eca = hgrant5_p & v1445ec6 | !hgrant5_p & v1445ec9;
assign v144649c = hgrant4_p & v845542 | !hgrant4_p & v144649b;
assign v134d26f = hlock2_p & v134d26d | !hlock2_p & v134d26e;
assign v1445b0c = hlock3 & v1445af2 | !hlock3 & v1445b0b;
assign a65922 = hmaster1_p & a658fd | !hmaster1_p & !a65916;
assign v1284d04 = hgrant2_p & v1284d02 | !hgrant2_p & v1284d03;
assign v1284d09 = locked_p & v140588d | !locked_p & v144639c;
assign v12163a0 = hmaster2_p & v1216ac7 | !hmaster2_p & v1216acf;
assign f2f3a4 = hmaster2_p & f2f355 | !hmaster2_p & f2f374;
assign v1445534 = hlock3 & v14454fa | !hlock3 & v1445532;
assign v10d4276 = hmaster0_p & v10d426f | !hmaster0_p & v10d4275;
assign v16a1d18 = hburst0 & v16a1d16 | !hburst0 & v16a1d17;
assign v1216201 = hmaster0_p & v12160d5 | !hmaster0_p & v12160d4;
assign v1668c9a = hmaster2_p & a658ca | !hmaster2_p & !v1668c64;
assign v1668d69 = stateA1_p & v845542 | !stateA1_p & v1668d68;
assign d301d9 = hgrant5_p & d301bb | !hgrant5_p & d301d8;
assign v138a487 = hbusreq2 & v138a481 | !hbusreq2 & v138a486;
assign v12ad00c = hgrant5_p & v12ad5c7 | !hgrant5_p & !v12ad00b;
assign v10d4095 = hgrant2_p & v10d4090 | !hgrant2_p & v10d4094;
assign v121611d = hready & v121611c | !hready & !v845542;
assign v1284d4e = hgrant5_p & v1405859 | !hgrant5_p & v1284d4d;
assign v144606c = hgrant5_p & v1445fdc | !hgrant5_p & v144606b;
assign v1446615 = hmaster2_p & v1446613 | !hmaster2_p & v1446614;
assign d80735 = hmaster0_p & d80734 | !hmaster0_p & v845542;
assign v1445890 = hbusreq4_p & v144639c | !hbusreq4_p & v144586d;
assign v143fd78 = hgrant4_p & v845542 | !hgrant4_p & v845572;
assign v1515769 = hbusreq1 & v10d3ff9 | !hbusreq1 & !v845542;
assign v1214c26 = hbusreq5 & v1214c11 | !hbusreq5 & v1214c25;
assign v12ad4cc = hbusreq0_p & a6585c | !hbusreq0_p & v845542;
assign v1216041 = hmaster0_p & v121603b | !hmaster0_p & v1216040;
assign d301a4 = hbusreq5_p & d301a3 | !hbusreq5_p & d30954;
assign v16a1da0 = hready_p & v16a1d82 | !hready_p & v16a1d9f;
assign v151581f = hmaster2_p & v151564d | !hmaster2_p & !a658ca;
assign v1214c6c = hbusreq4_p & v1214c6b | !hbusreq4_p & v845547;
assign v16a195b = hmaster0_p & v16a1951 | !hmaster0_p & v16a195a;
assign v1214dc5 = hbusreq3 & v1214dbd | !hbusreq3 & v1214dc4;
assign v1389fbe = hbusreq5_p & v1389fbd | !hbusreq5_p & v845542;
assign v1405aaa = hlock4_p & v1405a87 | !hlock4_p & !v845542;
assign v1446237 = hmaster1_p & v144639c | !hmaster1_p & v1446236;
assign v1216115 = hbusreq5_p & v1216113 | !hbusreq5_p & !v1216114;
assign v144610f = hlock2 & v144610c | !hlock2 & v144610e;
assign v1668d9a = hmaster2_p & v10d3fd8 | !hmaster2_p & !a65861;
assign v134d398 = hbusreq0 & v134d397 | !hbusreq0 & v134d38c;
assign v12161ab = hgrant5_p & v1216094 | !hgrant5_p & v1216132;
assign f2f35f = hmaster2_p & f2f34c | !hmaster2_p & f2f234;
assign f2f2cf = hbusreq1_p & f2f2ce | !hbusreq1_p & !v845542;
assign d8075d = stateG2_p & v845542 | !stateG2_p & d80755;
assign d30959 = hbusreq0 & d305fc | !hbusreq0 & d30958;
assign f2e3f9 = hmaster0_p & f2e715 | !hmaster0_p & f2e3f8;
assign v138a3a2 = hmaster1_p & v138a3a1 | !hmaster1_p & v138a341;
assign v14457c3 = hmaster1_p & v144579e | !hmaster1_p & v1445e28;
assign d2f9a4 = hbusreq4_p & d2f991 | !hbusreq4_p & v84554a;
assign v1445a4a = hmaster2_p & v14458d2 | !hmaster2_p & v1445a49;
assign a6629b = hgrant5_p & v845542 | !hgrant5_p & a6629a;
assign d30823 = hbusreq5_p & d30821 | !hbusreq5_p & d30822;
assign v1445be9 = hgrant3_p & v1445be2 | !hgrant3_p & v1445be8;
assign d300c5 = hmaster2_p & d300be | !hmaster2_p & d300c4;
assign d302f7 = hbusreq3_p & d302f6 | !hbusreq3_p & !d302ef;
assign v1445f99 = hmaster2_p & v1445f97 | !hmaster2_p & v1445f98;
assign v1215769 = hgrant4_p & v845542 | !hgrant4_p & v1215768;
assign v12ad5ea = hgrant5_p & v12ad501 | !hgrant5_p & v12ad5e8;
assign d3012d = hbusreq2_p & d3012b | !hbusreq2_p & d3012c;
assign v1668c77 = hbusreq1_p & v1668c76 | !hbusreq1_p & !v1668c63;
assign v1446641 = hgrant5_p & v1446445 | !hgrant5_p & v1446640;
assign d301ec = hgrant1_p & d301ea | !hgrant1_p & d301eb;
assign a66296 = hlock4_p & a66295 | !hlock4_p & !v845542;
assign v10d402e = hlock0_p & v10d3fe0 | !hlock0_p & v10d3fdf;
assign v14466b0 = hmaster0_p & v14465b8 | !hmaster0_p & v14466af;
assign v14058dd = hmaster1_p & v14058dc | !hmaster1_p & v140584d;
assign v16a1abd = hbusreq5_p & v16a2669 | !hbusreq5_p & v845568;
assign v1214ce2 = hmaster1_p & v1214ce1 | !hmaster1_p & v1214cd8;
assign a65499 = hmaster0_p & a658f1 | !hmaster0_p & a6548b;
assign v1284d46 = hmaster1_p & v1284d45 | !hmaster1_p & !v1284cdf;
assign v14058be = hgrant2_p & v14058b6 | !hgrant2_p & v14058bd;
assign v1446134 = hmaster0_p & v14460a5 | !hmaster0_p & v1446404;
assign d3068f = hbusreq4_p & v845542 | !hbusreq4_p & v84554a;
assign v134d3df = hmaster2_p & v134d3de | !hmaster2_p & v845542;
assign v10d4051 = hgrant2_p & v10d4018 | !hgrant2_p & v10d4050;
assign v15157c8 = hlock0_p & v1515630 | !hlock0_p & !v845542;
assign v1445b87 = hbusreq3 & v1445b72 | !hbusreq3 & v1445b86;
assign v12161ff = hbusreq2_p & v12161f6 | !hbusreq2_p & v12161fe;
assign v12152f5 = hmaster0_p & v12157a4 | !hmaster0_p & v121578e;
assign v1668d39 = hgrant5_p & v10d3fd8 | !hgrant5_p & v1668d37;
assign v16a13c2 = hbusreq2_p & v16a13c1 | !hbusreq2_p & v16a1da2;
assign v1216296 = hbusreq2_p & v1216293 | !hbusreq2_p & !v1216295;
assign v12ad4ef = hbusreq3 & v12ad4e3 | !hbusreq3 & v12ad4ee;
assign d2fb08 = hbusreq4_p & d30104 | !hbusreq4_p & d306a3;
assign v10d405d = hgrant0_p & v10d3fd5 | !hgrant0_p & !v10d3fd4;
assign v151566d = stateG2_p & v845542 | !stateG2_p & d3094b;
assign v12acfb3 = hlock0_p & v1668c6d | !hlock0_p & v845542;
assign v1445b75 = stateG10_5_p & v144668d | !stateG10_5_p & v1445b74;
assign v1214d12 = hbusreq0_p & v12166e5 | !hbusreq0_p & !v845542;
assign a658ea = hmaster0_p & a658b7 | !hmaster0_p & a658e8;
assign v11e5959 = hgrant1_p & v845542 | !hgrant1_p & v11e5958;
assign d305db = hmaster0_p & d305da | !hmaster0_p & d305d7;
assign d30229 = hgrant5_p & d30223 | !hgrant5_p & !d30227;
assign v1284cd1 = hlock5_p & v1284ccf | !hlock5_p & !v1284cd0;
assign v1445b15 = hbusreq2 & v1445b13 | !hbusreq2 & v1445b14;
assign v1515842 = hgrant5_p & v845570 | !hgrant5_p & v1515833;
assign v12160bd = hbusreq2_p & v12160bc | !hbusreq2_p & v12160bb;
assign v121616b = hgrant5_p & v121600b | !hgrant5_p & v121616a;
assign v155298f = jx1_p & v15530b7 | !jx1_p & v155298e;
assign v134cebb = hbusreq2 & v134ceba | !hbusreq2 & v134d270;
assign v134cd76 = hlock2 & v134cd6d | !hlock2 & v134cd75;
assign v12162df = hbusreq5 & v12162cd | !hbusreq5 & v12162de;
assign v1214ed7 = hbusreq0 & v1214ed2 | !hbusreq0 & v1214ed6;
assign f2f35b = hgrant5_p & f2f350 | !hgrant5_p & !f2f359;
assign v12ae76a = decide_p & v12afe3d | !decide_p & v12afe76;
assign v138a44a = hmaster0_p & v138a344 | !hmaster0_p & v138a32d;
assign v1216130 = hbusreq1_p & v121612f | !hbusreq1_p & v845542;
assign v1515702 = hmaster1_p & v15156f5 | !hmaster1_p & v15156e5;
assign d2f9ce = hlock2_p & d2f9cc | !hlock2_p & d2f9cd;
assign v138a441 = hmaster0_p & v138a3f7 | !hmaster0_p & v845542;
assign v1552f85 = hbusreq2 & v1552f83 | !hbusreq2 & v1552f84;
assign v1214dbe = hmaster0_p & v1214d2a | !hmaster0_p & v1214d27;
assign v16a1c04 = hbusreq5 & v16a1bfa | !hbusreq5 & v16a1c03;
assign v1214f07 = hlock5_p & v1214f05 | !hlock5_p & v1214f06;
assign v1216a63 = hburst0_p & v845584 | !hburst0_p & v845542;
assign v15532c7 = hgrant4_p & v845542 | !hgrant4_p & v15532c6;
assign v1215388 = hmaster0_p & v1215384 | !hmaster0_p & v1215387;
assign v1446209 = hgrant3_p & v1446160 | !hgrant3_p & v1446208;
assign a65ae1 = hgrant3_p & a662c6 | !hgrant3_p & a65ae0;
assign v10d428b = hgrant1_p & v10d3fdb | !hgrant1_p & v10d428a;
assign d307bf = hgrant1_p & v845542 | !hgrant1_p & d307be;
assign v12150c7 = hbusreq1_p & v12150c6 | !hbusreq1_p & v1215b97;
assign f2f2ec = hbusreq2 & f2f2e0 | !hbusreq2 & f2f2eb;
assign v121651a = hready_p & v1216aa1 | !hready_p & v1216519;
assign v12afda7 = hlock0_p & v1515c7d | !hlock0_p & v845542;
assign v16a1cf4 = hbusreq2_p & v16a1bde | !hbusreq2_p & v16a1cf3;
assign v138a329 = busreq_p & v845562 | !busreq_p & !v845542;
assign v1389dfb = hgrant2_p & v845542 | !hgrant2_p & !v1389dfa;
assign d2fbbb = hmaster1_p & d2fb7e | !hmaster1_p & d2fb9d;
assign v10d4038 = hmaster2_p & v10d402b | !hmaster2_p & !v10d3ff3;
assign f2f330 = hmaster0_p & f2f32f | !hmaster0_p & !f2f2da;
assign v12ad140 = decide_p & v12ad13f | !decide_p & v12afe76;
assign v1445b94 = hgrant2_p & v1445b69 | !hgrant2_p & v1445b93;
assign v134d271 = hbusreq5 & v134d26c | !hbusreq5 & v134d270;
assign v134cd60 = hlock0_p & v134d273 | !hlock0_p & v134cd5f;
assign v1214fe1 = hmaster0_p & v12153b5 | !hmaster0_p & v1215baf;
assign v1214c84 = hgrant2_p & v121657d | !hgrant2_p & v1214c7d;
assign f2f3dd = hgrant2_p & f2f3ae | !hgrant2_p & f2f3d0;
assign v144604b = hgrant5_p & v1446044 | !hgrant5_p & v144604a;
assign a66293 = stateA1_p & v845542 | !stateA1_p & !a66292;
assign v16a19c6 = hmaster1_p & v16a19b5 | !hmaster1_p & v16a1f96;
assign v12162fd = hmaster2_p & v1216aad | !hmaster2_p & v12162fc;
assign a65851 = locked_p & v845542 | !locked_p & v10d3fd8;
assign v16a19cd = decide_p & v16a1890 | !decide_p & !v16a19cc;
assign v16a1e2b = hbusreq2 & v16a1e25 | !hbusreq2 & v16a1e2a;
assign d2feb2 = hbusreq4_p & d2feb1 | !hbusreq4_p & v845542;
assign d2f98e = hmaster2_p & v84555a | !hmaster2_p & d2f98c;
assign d302dc = decide_p & d302db | !decide_p & v845570;
assign v1216005 = hbusreq1 & v1216004 | !hbusreq1 & v845542;
assign f2f371 = hgrant5_p & f2f35e | !hgrant5_p & !f2f370;
assign v1446191 = hbusreq2_p & v1446186 | !hbusreq2_p & v1446190;
assign a6565a = hgrant2_p & a6540e | !hgrant2_p & !a65653;
assign d2fb88 = hlock2_p & d2fb87 | !hlock2_p & d2fb80;
assign v138a076 = hready_p & v845542 | !hready_p & v138a075;
assign v1215cf9 = hbusreq0 & v1215cf6 | !hbusreq0 & v1215cf8;
assign f2f3bc = hgrant5_p & v84554c | !hgrant5_p & f2f359;
assign v14460f8 = hmaster1_p & v14460f7 | !hmaster1_p & v1445f9e;
assign v14460a3 = hmaster2_p & v144639c | !hmaster2_p & v14460a2;
assign d2fae5 = hbusreq5_p & d30117 | !hbusreq5_p & !d2fae4;
assign v134ce9e = hmaster1_p & v134d20b | !hmaster1_p & v134ce9d;
assign v138a3c5 = hgrant5_p & v845570 | !hgrant5_p & !v1515724;
assign v15157d8 = hgrant5_p & v845542 | !hgrant5_p & !v1515724;
assign v14058b9 = hgrant5_p & v1405859 | !hgrant5_p & v14058b7;
assign v1668d38 = hgrant5_p & a65851 | !hgrant5_p & v1668d37;
assign v1668d50 = hmaster2_p & a65394 | !hmaster2_p & !v1668d4f;
assign v10d401c = hgrant0_p & v10d401b | !hgrant0_p & !v10d3fd4;
assign a653aa = hbusreq1_p & a65360 | !hbusreq1_p & !a653a9;
assign v1445ec7 = hbusreq1 & v1445e65 | !hbusreq1 & v1445e69;
assign v1216b17 = hbusreq3 & v1216b08 | !hbusreq3 & v1216b16;
assign v12167a5 = hgrant2_p & v12167a2 | !hgrant2_p & v12167a4;
assign v960a34 = hburst0_p & v845542 | !hburst0_p & v8a9c96;
assign d306fe = hlock1_p & a65861 | !hlock1_p & !v845542;
assign v12161a9 = hgrant5_p & v1216094 | !hgrant5_p & v121612a;
assign v12160f8 = hgrant1_p & v845542 | !hgrant1_p & v12160f7;
assign v134d293 = hgrant5_p & v845542 | !hgrant5_p & v134d292;
assign v12acff8 = hbusreq0_p & v1515790 | !hbusreq0_p & v845542;
assign v12166c6 = hmaster2_p & v12166c5 | !hmaster2_p & v1216588;
assign a6540a = hmaster1_p & a65409 | !hmaster1_p & a65893;
assign d2faeb = hgrant4_p & v845558 | !hgrant4_p & d2faea;
assign v12aef0b = hgrant3_p & v12af3ae | !hgrant3_p & v12aef0a;
assign d307d0 = hbusreq0_p & v845542 | !hbusreq0_p & v1668d48;
assign v16a1a8c = hbusreq5 & v16a1a82 | !hbusreq5 & v16a1a8b;
assign v14458d9 = hbusreq4 & v14458d7 | !hbusreq4 & v14458d8;
assign v14466d0 = hmaster0_p & v14463c7 | !hmaster0_p & v144639c;
assign v14459ce = hbusreq1_p & v14465b2 | !hbusreq1_p & v14459cd;
assign v138a360 = hmaster1_p & v138a35f | !hmaster1_p & v138a341;
assign v121616c = hgrant5_p & v1216026 | !hgrant5_p & v121616a;
assign v14465c8 = hgrant0_p & v144640a | !hgrant0_p & v14463d8;
assign f2f3bb = hgrant5_p & f2f2a8 | !hgrant5_p & !f2f359;
assign v1515779 = hbusreq4_p & v151572b | !hbusreq4_p & v1515754;
assign v1389f91 = hlock5_p & v1389f90 | !hlock5_p & v845542;
assign v12ad611 = hbusreq5_p & v12ad60e | !hbusreq5_p & v12ad610;
assign v1445adf = hlock3 & v1445ad6 | !hlock3 & v1445ade;
assign v1445db3 = hmaster1_p & v1445db2 | !hmaster1_p & v1445da4;
assign v1445766 = hbusreq2 & v1445760 | !hbusreq2 & v1445761;
assign v1446473 = hgrant5_p & v1446467 | !hgrant5_p & v1446472;
assign v1445444 = hmaster1_p & v1445443 | !hmaster1_p & v1446219;
assign v1515762 = hbusreq4 & a653c8 | !hbusreq4 & !v151563e;
assign f2e715 = hgrant5_p & v845542 | !hgrant5_p & !f2e714;
assign d306a9 = hbusreq5_p & d3064c | !hbusreq5_p & !d306a8;
assign v1216090 = hbusreq1 & v1216048 | !hbusreq1 & v845542;
assign d30614 = hmaster0_p & d305ed | !hmaster0_p & d30613;
assign v1668d8e = hmaster2_p & v10d3fd8 | !hmaster2_p & !a65394;
assign a6563a = hbusreq5_p & a653a8 | !hbusreq5_p & !a65639;
assign v14058d1 = hbusreq0_p & v140583f | !hbusreq0_p & v14058c5;
assign v138a314 = hmaster0_p & v138a312 | !hmaster0_p & v138a313;
assign v1215764 = hlock0_p & v1215b8f | !hlock0_p & v845547;
assign v1552960 = decide_p & v155342e | !decide_p & v15530f2;
assign v12ad599 = hbusreq1 & v12ad4f0 | !hbusreq1 & !v845542;
assign a662c7 = hbusreq1_p & a66285 | !hbusreq1_p & a66289;
assign d306ac = hgrant5_p & v845542 | !hgrant5_p & !d306ab;
assign v144611b = hmaster1_p & v144611a | !hmaster1_p & v1445fde;
assign v138938f = hbusreq0 & v1389ffd | !hbusreq0 & v138a403;
assign v12ad32b = hgrant2_p & v12af73f | !hgrant2_p & v12ad32a;
assign d2fd15 = hbusreq2_p & d2fd14 | !hbusreq2_p & d302d6;
assign d80741 = hbusreq5_p & d80740 | !hbusreq5_p & !d8073f;
assign v1445e75 = hmaster2_p & v1445e74 | !hmaster2_p & v1445e6c;
assign v16693ae = hmaster1_p & v16693ad | !hmaster1_p & v845542;
assign v1515624 = hburst1 & v1552d7a | !hburst1 & v1515623;
assign v134ce3a = hgrant5_p & v134d36a | !hgrant5_p & v134ce39;
assign v1445922 = hlock2 & v1445912 | !hlock2 & v1445920;
assign d30107 = hgrant1_p & d300fa | !hgrant1_p & d30106;
assign v16a1d42 = hgrant5_p & v845542 | !hgrant5_p & v16a1d41;
assign v138a405 = hbusreq5 & v138a3fc | !hbusreq5 & v138a404;
assign v138a343 = hmaster2_p & v138a32b | !hmaster2_p & a658c6;
assign v16a1be9 = hmaster1_p & v16a1be2 | !hmaster1_p & v16a1be8;
assign bf1f5c = hgrant5_p & v845542 | !hgrant5_p & !d3064a;
assign v1668cd1 = hlock0_p & v1668cbd | !hlock0_p & !v845542;
assign v12ad4e7 = hmaster2_p & v12ad4e4 | !hmaster2_p & !v12ad4e6;
assign v14466d1 = hmaster1_p & v14466d0 | !hmaster1_p & v14463cd;
assign v16693a7 = hmaster2_p & v845542 | !hmaster2_p & !v16693a6;
assign v12ad541 = hmaster0_p & v12ad52d | !hmaster0_p & v12ad531;
assign v14454fa = hbusreq2_p & v14454f9 | !hbusreq2_p & v1445bdb;
assign v134ce99 = hlock5_p & v134ce98 | !hlock5_p & v134d1fd;
assign v1389814 = hgrant5_p & a65892 | !hgrant5_p & !v845542;
assign v16a19e5 = hmaster1_p & v16a19e4 | !hmaster1_p & v16a2672;
assign v1668daa = hgrant2_p & v1668da9 | !hgrant2_p & v1668d8c;
assign v16a209b = hgrant5_p & v845542 | !hgrant5_p & !v16a208a;
assign v14453b6 = hbusreq2_p & v14453b3 | !hbusreq2_p & v14453b5;
assign d30189 = hbusreq2_p & d3091b | !hbusreq2_p & d30188;
assign f2f423 = hgrant1_p & f2f281 | !hgrant1_p & !f2f373;
assign v1216180 = hgrant2_p & v1216174 | !hgrant2_p & !v121617f;
assign v12ad002 = hgrant4_p & v12ad5c0 | !hgrant4_p & !v12ad001;
assign v10d409b = hmaster1_p & v10d409a | !hmaster1_p & v10d3ffb;
assign v14453a3 = hbusreq3 & v14453a1 | !hbusreq3 & v14453a2;
assign v1445843 = hmaster1_p & v14457da | !hmaster1_p & v1445f09;
assign v134ce35 = hlock1 & v134d273 | !hlock1 & v134ce34;
assign v1445aa4 = hlock2 & v1445aa0 | !hlock2 & v1445aa3;
assign v144643b = hmaster2_p & v144639c | !hmaster2_p & v1446406;
assign f2f2d3 = hbusreq1_p & f2f2d2 | !hbusreq1_p & v845542;
assign v12152e4 = hmaster0_p & v1215b8a | !hmaster0_p & v1215b7c;
assign v1445377 = hlock3 & v1445354 | !hlock3 & v1445375;
assign v1668d6e = hbusreq4 & a6585c | !hbusreq4 & v1668d6d;
assign v12164dc = hbusreq4_p & v845570 | !hbusreq4_p & v12164cf;
assign v1668d5f = hgrant5_p & v1668d50 | !hgrant5_p & !v1668d5e;
assign v16a1414 = hbusreq2_p & v16a1413 | !hbusreq2_p & v16a205f;
assign v12ad571 = hbusreq2 & v12ad568 | !hbusreq2 & v12ad570;
assign f2e277 = hmaster2_p & v845542 | !hmaster2_p & !f2e276;
assign v1552f7e = hmaster0_p & v1552f7d | !hmaster0_p & v1552f68;
assign v144674b = hmaster0_p & v1446448 | !hmaster0_p & v144663a;
assign d30249 = hlock5_p & d30247 | !hlock5_p & !d30248;
assign v1445a08 = hlock0 & v14459f1 | !hlock0 & v1445a07;
assign v1446400 = hbusreq3 & v14463fe | !hbusreq3 & v14463ff;
assign v144590d = hlock2 & v1445905 | !hlock2 & v144590c;
assign v15155ff = hmaster1_p & v15155fc | !hmaster1_p & v15155fe;
assign v1515636 = hbusreq2 & v1515635 | !hbusreq2 & v845542;
assign v1215ccd = hgrant5_p & v845570 | !hgrant5_p & v1215c87;
assign v1389fe8 = hmaster1_p & v1389de1 | !hmaster1_p & v1389fe7;
assign v1214ced = hmaster2_p & v1214cec | !hmaster2_p & v1214cbc;
assign v1405b3e = hmaster1_p & v1405b3d | !hmaster1_p & !v1405a94;
assign v12afe46 = hgrant1_p & v845542 | !hgrant1_p & v12afe45;
assign v1214c4d = hbusreq1 & v121534b | !hbusreq1 & v845542;
assign d2fbd0 = hgrant0_p & v845542 | !hgrant0_p & d2fbcf;
assign v1216132 = hmaster2_p & v1216131 | !hmaster2_p & v845542;
assign v138a403 = hbusreq5_p & v138a402 | !hbusreq5_p & !v845542;
assign v14058e7 = locked_p & v1405860 | !locked_p & !v144639c;
assign v1445f09 = hmaster0_p & v1445f08 | !hmaster0_p & v1445ea9;
assign v1445bf7 = hready_p & v1445bca | !hready_p & v1445bf3;
assign v15157a2 = hgrant5_p & v1668da6 | !hgrant5_p & v15157a1;
assign v1445553 = hready_p & v1446564 | !hready_p & v1445552;
assign v1445426 = hlock3 & v144541f | !hlock3 & v1445425;
assign v16a12ea = hgrant1_p & v84554d | !hgrant1_p & v16a12e9;
assign v1405907 = hmaster1_p & v1405906 | !hmaster1_p & v140584d;
assign v1445997 = hlock0_p & v1445996 | !hlock0_p & v144639c;
assign v14458b8 = hmaster2_p & v1445871 | !hmaster2_p & v1445885;
assign v1552d99 = hgrant3_p & v155321c | !hgrant3_p & v1552d98;
assign v1552d7e = hgrant1_p & v1552d7d | !hgrant1_p & v845542;
assign v1215792 = hgrant5_p & v1215791 | !hgrant5_p & v121573e;
assign v1445394 = hmaster1_p & v1445366 | !hmaster1_p & v1445a82;
assign v1405883 = hmaster0_p & v1405841 | !hmaster0_p & v1405840;
assign v1668d12 = hlock3_p & v1668cb6 | !hlock3_p & v1668d11;
assign v134d447 = hbusreq2 & v134d445 | !hbusreq2 & v134d446;
assign f2e3fa = hmaster1_p & f2f229 | !hmaster1_p & f2e3f9;
assign a6567e = hgrant2_p & a6540e | !hgrant2_p & !a6567a;
assign f2f357 = hbusreq1_p & f2f356 | !hbusreq1_p & v845542;
assign v121540b = hbusreq3 & v12153f8 | !hbusreq3 & v121540a;
assign f2f3b8 = hgrant5_p & f2f2a8 | !hgrant5_p & !f2f34d;
assign v121508c = hgrant4_p & v1215026 | !hgrant4_p & v121508b;
assign d2feac = hbusreq3 & d2fea7 | !hbusreq3 & !d2feab;
assign v151571e = stateA1_p & v84557e | !stateA1_p & !v151571d;
assign v1216162 = hgrant4_p & v1216148 | !hgrant4_p & v121656a;
assign v12157a3 = hgrant5_p & v845542 | !hgrant5_p & v121577a;
assign f2ec23 = hmaster2_p & v845542 | !hmaster2_p & !f2ec22;
assign v1215473 = hmaster1_p & v1215472 | !hmaster1_p & v121546f;
assign v1214c0f = hbusreq2_p & v1214c0e | !hbusreq2_p & v1214c0d;
assign d30718 = hmastlock_p & d30717 | !hmastlock_p & !v845542;
assign d3014f = hmaster1_p & d30137 | !hmaster1_p & d3014e;
assign v134d42d = hgrant1_p & v845542 | !hgrant1_p & v134d42c;
assign v10d4294 = hbusreq1_p & v10d428a | !hbusreq1_p & v10d4293;
assign v1215c40 = hbusreq5_p & v1215c3e | !hbusreq5_p & !v1215c3f;
assign v16a1cd5 = hmaster0_p & v16a1cd0 | !hmaster0_p & v16a1ccc;
assign v1445abf = hbusreq2_p & v1445abd | !hbusreq2_p & v1445abe;
assign d307da = hbusreq1_p & d307d9 | !hbusreq1_p & v845542;
assign v1445af9 = hbusreq2_p & v1445af6 | !hbusreq2_p & v1445af8;
assign v1446410 = hbusreq1_p & v1446403 | !hbusreq1_p & v144640f;
assign f2f52e = hgrant2_p & v845542 | !hgrant2_p & f2f52d;
assign v12af21c = hgrant1_p & d30690 | !hgrant1_p & v12af21b;
assign v138a011 = hbusreq5 & v1389ff5 | !hbusreq5 & v138a010;
assign v15156e8 = hbusreq2_p & v15156e7 | !hbusreq2_p & v845542;
assign v14458b6 = hlock3 & v14458b3 | !hlock3 & v14458b5;
assign a653c0 = hbusreq0 & a653b7 | !hbusreq0 & a653bf;
assign v12160d4 = hmaster2_p & v12160d1 | !hmaster2_p & v12160d3;
assign v14459d9 = hgrant0_p & v1446403 | !hgrant0_p & v14459d8;
assign v1214fb6 = hbusreq0 & v121578c | !hbusreq0 & v1214fb5;
assign stateG10_4 = !v14838bf;
assign a6538b = hgrant5_p & a65852 | !hgrant5_p & a6538a;
assign d3019e = hmaster0_p & d3019d | !hmaster0_p & !d30917;
assign f2f360 = hgrant5_p & f2f35e | !hgrant5_p & !f2f35f;
assign v1553145 = hlock5_p & v1553143 | !hlock5_p & v1553144;
assign v1445dda = hlock2 & v1445dd7 | !hlock2 & v1445dd9;
assign v12ad01d = hmaster1_p & v12ad01c | !hmaster1_p & v12ad666;
assign v14458fc = hlock0 & v14458fb | !hlock0 & v14458f9;
assign v144599f = hgrant5_p & v14458d4 | !hgrant5_p & v144599e;
assign v12ad5ba = hlock0_p & v1515741 | !hlock0_p & v845542;
assign v14463a8 = hbusreq5_p & v144639c | !hbusreq5_p & v14463a6;
assign d2fb0a = hbusreq1_p & d30106 | !hbusreq1_p & d2fb09;
assign v1553216 = hlock3_p & v1553154 | !hlock3_p & v1553215;
assign a658e7 = hmaster1_p & a658b7 | !hmaster1_p & a658e5;
assign v1516214 = hready_p & v1516201 | !hready_p & !v1516213;
assign v151582a = hmaster1_p & v1515820 | !hmaster1_p & !v15156da;
assign d2fe8f = hmaster0_p & d2fe7e | !hmaster0_p & d2fe8e;
assign f2f3f7 = hbusreq2_p & f2f3f4 | !hbusreq2_p & f2f3f6;
assign v16a1a2f = hbusreq5 & v16a1a23 | !hbusreq5 & v16a1a2e;
assign d30783 = hbusreq4_p & d30782 | !hbusreq4_p & !d30781;
assign d2fb2d = hbusreq2_p & d2fb1a | !hbusreq2_p & !d2fb2c;
assign d30150 = hgrant2_p & d300b4 | !hgrant2_p & d3014f;
assign a653da = hbusreq0_p & a653d9 | !hbusreq0_p & a65396;
assign v1445d98 = hbusreq4_p & v1445d97 | !hbusreq4_p & v14463bb;
assign v1215c97 = hgrant5_p & v845542 | !hgrant5_p & !v1215c95;
assign v121574c = hmaster2_p & v121572b | !hmaster2_p & v121574b;
assign v12af983 = hlock0_p & v84556a | !hlock0_p & v845542;
assign v1214d1c = hbusreq5_p & v1214d1b | !hbusreq5_p & v1214cfb;
assign v138a457 = hmaster0_p & v138a354 | !hmaster0_p & v138a32d;
assign v11e595d = hmaster1_p & v11e5948 | !hmaster1_p & !v11e595c;
assign v1552f5a = hgrant5_p & v1553386 | !hgrant5_p & v1552f59;
assign a656ce = hmaster1_p & a66287 | !hmaster1_p & a656cd;
assign v151563e = locked_p & a658db | !locked_p & v845542;
assign d30677 = hgrant2_p & d30676 | !hgrant2_p & d3066e;
assign v1216326 = hgrant2_p & v1216323 | !hgrant2_p & v121631d;
assign v1668d10 = hbusreq3 & v1668d0f | !hbusreq3 & v845542;
assign v14458df = hlock0_p & v14458dd | !hlock0_p & v14458de;
assign v16a1d56 = hbusreq2 & v16a1d54 | !hbusreq2 & !v16a1d55;
assign v1553236 = hmaster2_p & v1553231 | !hmaster2_p & v1553235;
assign f2e4dc = hmaster1_p & f2f229 | !hmaster1_p & f2e4db;
assign v1668ddd = hbusreq0 & v1668dd9 | !hbusreq0 & v1668ddc;
assign d30244 = hlock5_p & d30241 | !hlock5_p & !d30243;
assign v1445f9f = hmaster1_p & v144639c | !hmaster1_p & v1445f9e;
assign v155338e = hbusreq1 & v155338d | !hbusreq1 & v1553217;
assign v10d4020 = hbusreq4_p & v10d3fdb | !hbusreq4_p & !v10d3fd8;
assign v16a2070 = hmaster2_p & v16a206d | !hmaster2_p & v16a206f;
assign v121655a = hmaster2_p & v1216555 | !hmaster2_p & v1216559;
assign v144647d = hbusreq4_p & v1446398 | !hbusreq4_p & v144646e;
assign v16a197b = hgrant5_p & v845542 | !hgrant5_p & !v16a1970;
assign v1445ba5 = hlock5 & v144632f | !hlock5 & v1445ba4;
assign d30666 = hgrant0_p & d30665 | !hgrant0_p & !v845570;
assign v1445909 = hlock0 & v1445908 | !hlock0 & v1445907;
assign v151560d = locked_p & v845542 | !locked_p & !v10d3fdf;
assign v144547a = hmaster1_p & v1445479 | !hmaster1_p & v144627e;
assign v12150bf = hbusreq2_p & v12150bc | !hbusreq2_p & v12150be;
assign v1445a7c = hmaster2_p & v1445a53 | !hmaster2_p & v14459fc;
assign v1668d45 = hbusreq1 & a65394 | !hbusreq1 & a65396;
assign v16a12f4 = hmaster1_p & v16a12f3 | !hmaster1_p & v16a209c;
assign a66289 = hgrant4_p & v845570 | !hgrant4_p & !v845542;
assign v134d383 = hgrant1_p & v845542 | !hgrant1_p & v134d382;
assign v134ce79 = hbusreq5 & v134ce77 | !hbusreq5 & v134ce78;
assign v1445b02 = hmaster1_p & v1445b01 | !hmaster1_p & v14458fd;
assign v144576d = hlock2 & v1445f40 | !hlock2 & v144576b;
assign d2fd46 = hbusreq2_p & d2fd2c | !hbusreq2_p & !d302eb;
assign v15168f2 = hburst0 & a66293 | !hburst0 & v15168f1;
assign v138a352 = hlock2_p & v138a34d | !hlock2_p & v138a351;
assign v138936d = hlock5_p & v138936c | !hlock5_p & v845542;
assign a65adc = decide_p & a65adb | !decide_p & a662a2;
assign v1405abc = hmaster2_p & v1405abb | !hmaster2_p & v1405a88;
assign v12147ee = hmaster1_p & v12147ed | !hmaster1_p & v1215d79;
assign d30805 = hmaster0_p & d307a6 | !hmaster0_p & d30804;
assign v1445797 = hlock2 & v1445790 | !hlock2 & v1445796;
assign v155321b = decide_p & v1553216 | !decide_p & v155321a;
assign v1216237 = hmaster0_p & v1216209 | !hmaster0_p & v1216236;
assign v1215464 = hmaster0_p & v1215462 | !hmaster0_p & v1215463;
assign v14466a1 = hmaster2_p & v144669c | !hmaster2_p & v1446603;
assign v1668d27 = hgrant4_p & v1668d26 | !hgrant4_p & a6536e;
assign v1552990 = jx0_p & v1552da3 | !jx0_p & v155298f;
assign v14058d9 = hmaster1_p & v14058c4 | !hmaster1_p & v14058d8;
assign v151570d = decide_p & v151570c | !decide_p & v845542;
assign v1214fb9 = hbusreq4_p & v1214fb8 | !hbusreq4_p & v845542;
assign a654b0 = hmaster0_p & a654af | !hmaster0_p & a65475;
assign v16a1968 = hmaster0_p & v16a1964 | !hmaster0_p & v16a1967;
assign v151564c = hburst0 & v1515648 | !hburst0 & v151564b;
assign v16a1d66 = hbusreq2 & v16a1d64 | !hbusreq2 & !v16a1d65;
assign v16a13e7 = hlock2_p & v16a13e0 | !hlock2_p & v16a13e6;
assign d30743 = hbusreq1_p & d30742 | !hbusreq1_p & v845542;
assign v1445eaa = hmaster0_p & v1445e86 | !hmaster0_p & v1445ea9;
assign v1668c2b = hmaster0_p & v1668c2a | !hmaster0_p & v845542;
assign v16a19b2 = hmaster1_p & v16a19b1 | !hmaster1_p & !v16a2672;
assign v16a2085 = hgrant1_p & v84554d | !hgrant1_p & v16a2084;
assign v84556c = start_p & v845542 | !start_p & !v845542;
assign v14465e4 = hbusreq5_p & v14465e3 | !hbusreq5_p & v14465dd;
assign v1405b0a = hmaster1_p & v1405ad8 | !hmaster1_p & v1405b09;
assign v1445e5c = hbusreq1_p & v144639c | !hbusreq1_p & v1445e5b;
assign v10d4011 = hbusreq2_p & v10d400d | !hbusreq2_p & v10d4010;
assign a653e5 = hbusreq5_p & a653e3 | !hbusreq5_p & a653e4;
assign d306eb = hburst0_p & v845542 | !hburst0_p & d306ea;
assign d2fb9a = hlock5_p & d2fb99 | !hlock5_p & d2fb72;
assign d302ec = hbusreq2_p & d302e6 | !hbusreq2_p & !d302eb;
assign v134d23b = hbusreq5_p & v134d23a | !hbusreq5_p & v134d1fd;
assign v1215ff6 = hmastlock_p & v1215ff5 | !hmastlock_p & v845542;
assign v12ad5ce = hbusreq5_p & v12ad5c6 | !hbusreq5_p & !v12ad5cd;
assign v144641e = hlock1 & v144641d | !hlock1 & v144641c;
assign v12160e2 = hmaster2_p & v12160d1 | !hmaster2_p & v12160d8;
assign v121613e = hbusreq4_p & v12160fb | !hbusreq4_p & v12afe44;
assign v14058a7 = hbusreq4_p & v14058a6 | !hbusreq4_p & v140589a;
assign d300ff = hmaster2_p & d30662 | !hmaster2_p & d300fe;
assign f2f34c = hgrant1_p & v845570 | !hgrant1_p & !f2f34b;
assign a6537f = hbusreq4_p & a6537e | !hbusreq4_p & v845542;
assign v12acfbe = hmaster0_p & v12ad528 | !hmaster0_p & v12ad531;
assign d2f97e = hmaster1_p & d2f975 | !hmaster1_p & !d2f97d;
assign v12ad4d4 = hlock0_p & v151560d | !hlock0_p & d2fbe5;
assign v14058c4 = hgrant5_p & v1405841 | !hgrant5_p & v14058c3;
assign d80752 = hlock3_p & d8074c | !hlock3_p & d80751;
assign v1215ce4 = hgrant5_p & v845542 | !hgrant5_p & v1215c8d;
assign v1445d81 = hbusreq4_p & v14463a0 | !hbusreq4_p & v144639e;
assign v134d366 = hgrant4_p & v845542 | !hgrant4_p & v134d365;
assign v134d36c = hmastlock_p & v134d36b | !hmastlock_p & v845542;
assign v14460da = hbusreq2_p & v14460d1 | !hbusreq2_p & v14460d9;
assign v1215089 = hbusreq2_p & v1215086 | !hbusreq2_p & v1215088;
assign v121658d = stateG2_p & v845542 | !stateG2_p & v121658c;
assign v1446622 = hgrant5_p & v14465ea | !hgrant5_p & v1446621;
assign v1446681 = hmaster1_p & v1446680 | !hmaster1_p & v1446436;
assign v1216152 = hgrant4_p & v1216150 | !hgrant4_p & v1216151;
assign v1445a22 = hbusreq4 & v1445a21 | !hbusreq4 & v14459b3;
assign v1215797 = hgrant5_p & v1215791 | !hgrant5_p & v121574c;
assign v1445a0d = hbusreq4_p & v144639c | !hbusreq4_p & v1445a0c;
assign d30231 = hmaster2_p & v845542 | !hmaster2_p & !d3070c;
assign d301f2 = hlock1_p & d306d5 | !hlock1_p & v1668d52;
assign v1445ff4 = hlock2 & v1445ff3 | !hlock2 & v1445fed;
assign v1214f50 = hgrant2_p & v845542 | !hgrant2_p & v1214f4f;
assign d3026f = hgrant5_p & v845570 | !hgrant5_p & d3026e;
assign v1215c36 = hmaster1_p & v1215c06 | !hmaster1_p & v1215c35;
assign v12ad587 = hbusreq2 & v12ad581 | !hbusreq2 & v12ad586;
assign v134d3a9 = hbusreq1 & v134d370 | !hbusreq1 & v134d371;
assign v1215bca = hmaster1_p & v1215bb4 | !hmaster1_p & v1215bc2;
assign v144633c = hbusreq5_p & v144668e | !hbusreq5_p & v144633b;
assign v1515c87 = decide_p & v1515c86 | !decide_p & v845542;
assign d3028f = hmaster2_p & v1668c1c | !hmaster2_p & !v845570;
assign v14454ee = hbusreq0 & v14454eb | !hbusreq0 & v14454ed;
assign v1445b8f = hgrant2_p & v144634f | !hgrant2_p & v1445b8e;
assign v1214c98 = hmaster1_p & v1214c97 | !hmaster1_p & v1214c92;
assign v1515805 = hbusreq2_p & v1515804 | !hbusreq2_p & !v845542;
assign v11e5943 = hlock2_p & v11e5942 | !hlock2_p & bf1f59;
assign v1552f76 = hbusreq2 & v1552f74 | !hbusreq2 & v1552f75;
assign v1446666 = hgrant2_p & v1446659 | !hgrant2_p & v1446665;
assign a65418 = hbusreq5_p & a65414 | !hbusreq5_p & !a65416;
assign v121510e = hmaster0_p & v1215057 | !hmaster0_p & v1215471;
assign d2fc15 = hbusreq2_p & d2fc13 | !hbusreq2_p & d2fc14;
assign v14460be = hmaster1_p & v1446093 | !hmaster1_p & v14460b6;
assign v14460d0 = hmaster1_p & v144603f | !hmaster1_p & v14460cf;
assign a6470a = hgrant3_p & a646dc | !hgrant3_p & a64709;
assign v1216232 = hmaster2_p & v12160d1 | !hmaster2_p & !v1216231;
assign d2fb76 = hlock0_p & v845542 | !hlock0_p & a66275;
assign v16a1bc3 = hbusreq1 & v16a1bc2 | !hbusreq1 & v16a2089;
assign d30886 = hmaster1_p & d30885 | !hmaster1_p & !d30858;
assign v12ad538 = hmaster1_p & v12ad537 | !hmaster1_p & !v12ad525;
assign v1216222 = hgrant5_p & v12160df | !hgrant5_p & v1216221;
assign v1216a9a = hbusreq5_p & v1216a99 | !hbusreq5_p & v845542;
assign v12150a8 = hgrant2_p & v1215063 | !hgrant2_p & v12150a7;
assign v14460bf = hgrant2_p & v14460bd | !hgrant2_p & v14460be;
assign v1445b9c = hgrant2_p & v1445b6e | !hgrant2_p & v1445b93;
assign v1445aae = hready_p & v1445bca | !hready_p & v1445aad;
assign v14458d3 = hmaster2_p & v14458d2 | !hmaster2_p & v144639c;
assign v1215fef = hbusreq1_p & v1215fee | !hbusreq1_p & v845542;
assign v10d40d1 = hmaster0_p & v10d400e | !hmaster0_p & v10d400a;
assign v14465b8 = hbusreq5_p & v14465b5 | !hbusreq5_p & v14465b7;
assign v1445e37 = hready_p & v144639b | !hready_p & v1445e36;
assign a662ae = hbusreq5_p & a66287 | !hbusreq5_p & a662ad;
assign v14457d4 = decide_p & v1445774 | !decide_p & v14457d3;
assign v12164e5 = hmaster1_p & v12164e4 | !hmaster1_p & v12164e1;
assign v1215341 = decide_p & v121545c | !decide_p & v1215340;
assign v138a3e1 = hmaster1_p & v138a3cb | !hmaster1_p & v138a3e0;
assign v144617a = hgrant2_p & v1446178 | !hgrant2_p & v1446179;
assign v16a1db1 = hbusreq0 & v16a1db0 | !hbusreq0 & v16a208b;
assign v1216a9d = hmaster0_p & v1216a8f | !hmaster0_p & v1668c1f;
assign f2f2f1 = hbusreq2_p & f2f2ee | !hbusreq2_p & f2f2f0;
assign v1215c05 = hbusreq0 & v1215c00 | !hbusreq0 & v1215c04;
assign v1216799 = hmaster0_p & v12166f3 | !hmaster0_p & v12164d7;
assign v134ce39 = hmaster2_p & v845542 | !hmaster2_p & v134ce38;
assign f2f44a = hgrant5_p & f2f3c1 | !hgrant5_p & f2f428;
assign v15533ae = hlock1 & v15533a1 | !hlock1 & v15533ad;
assign v1668d06 = hgrant2_p & v1668d02 | !hgrant2_p & v1668d05;
assign v1515806 = hbusreq2 & v1515805 | !hbusreq2 & v1516803;
assign v1445a83 = hmaster1_p & v14459a3 | !hmaster1_p & v1445a82;
assign v1445a60 = hmaster1_p & v144598e | !hmaster1_p & v144590e;
assign v14460b9 = hmaster1_p & v144607a | !hmaster1_p & v1445ffc;
assign v121626f = hmaster0_p & v1216172 | !hmaster0_p & v1216029;
assign v15156bc = hmaster2_p & v151564d | !hmaster2_p & !v15156bb;
assign v16a1c9c = hmaster1_p & v16a1c9b | !hmaster1_p & !v16a2672;
assign v12afe76 = hgrant2_p & v845542 | !hgrant2_p & v12afe75;
assign a656d3 = hgrant3_p & a65b07 | !hgrant3_p & a656d2;
assign v12ad67c = hlock0_p & a658ca | !hlock0_p & v845542;
assign v12166e6 = hbusreq0_p & v12166e5 | !hbusreq0_p & v12166ce;
assign v1445a5c = hmaster1_p & v1445a5b | !hmaster1_p & v1445a32;
assign v14466ac = hgrant5_p & v144643a | !hgrant5_p & v1446640;
assign v1215be8 = hmaster2_p & v121601f | !hmaster2_p & v1215be6;
assign v85e749 = hmaster1_p & v84554c | !hmaster1_p & ae2496;
assign d3088e = hbusreq1_p & d3079e | !hbusreq1_p & d306a5;
assign v144671a = hlock2 & v1446716 | !hlock2 & v1446719;
assign v16a207b = hbusreq5_p & v16a2079 | !hbusreq5_p & v16a207a;
assign d300da = hbusreq1_p & d300d7 | !hbusreq1_p & d300d9;
assign v16a2067 = hready_p & v845555 | !hready_p & !v16a2066;
assign d301b9 = decide_p & d301b8 | !decide_p & v845570;
assign v1405910 = decide_p & v140590a | !decide_p & v140590f;
assign v1216014 = hready & v1216a66 | !hready & v1216013;
assign v14459a1 = hmaster2_p & v14459a0 | !hmaster2_p & v14465b3;
assign v16a13d9 = decide_p & v16a13d8 | !decide_p & !v16a2065;
assign v12164c6 = hmaster0_p & v1216afb | !hmaster0_p & v1216b03;
assign v14463ac = hlock1 & v144639c | !hlock1 & v14463ab;
assign v1445491 = hlock2 & v144546f | !hlock2 & v1445490;
assign v134ce88 = hbusreq2 & v134ce87 | !hbusreq2 & v134d240;
assign v1668ccd = hburst0 & a66272 | !hburst0 & v1668ccc;
assign v1668e0f = jx2_p & v1668e04 | !jx2_p & v1668e0e;
assign v134d203 = hlock0 & v134d202 | !hlock0 & v134d1fe;
assign v10d406d = hgrant1_p & v10d3fe0 | !hgrant1_p & v10d4067;
assign v1405932 = hgrant2_p & v1405924 | !hgrant2_p & v1405931;
assign v12160eb = hbusreq4 & v1215fe8 | !hbusreq4 & v845542;
assign v12ad54f = hmaster0_p & v12ad54e | !hmaster0_p & !v12ad524;
assign v1215451 = hmaster1_p & v1215448 | !hmaster1_p & v121540f;
assign v16a188a = hmaster1_p & v16a1843 | !hmaster1_p & !v16a1f96;
assign v131be8e = decide_p & v131be8a | !decide_p & v131be8d;
assign v1515631 = hmaster2_p & v845570 | !hmaster2_p & v1515630;
assign v1216087 = hmaster1_p & v1216069 | !hmaster1_p & v1216082;
assign v1445a29 = hbusreq4_p & v14465b1 | !hbusreq4_p & v1445a28;
assign v1445fed = hbusreq2_p & v1445fdf | !hbusreq2_p & v1445fec;
assign v16a1db4 = hbusreq2_p & v16a1d54 | !hbusreq2_p & v16a1db3;
assign v845562 = hburst1_p & v845542 | !hburst1_p & !v845542;
assign v12ae201 = hgrant2_p & v845542 | !hgrant2_p & v12ae200;
assign v1214bcd = hbusreq5_p & v1214bcc | !hbusreq5_p & v1214bcb;
assign v14453ee = hbusreq3 & v14453ec | !hbusreq3 & v14453ed;
assign v1446100 = hlock3 & v14460f2 | !hlock3 & v14460fe;
assign v134d4ac = hbusreq0 & v134d4ab | !hbusreq0 & v134d379;
assign v138a3eb = hbusreq5_p & v138a3ea | !hbusreq5_p & !v845542;
assign v14458a4 = hmaster2_p & v144639c | !hmaster2_p & v1445888;
assign v134d286 = hgrant5_p & v134d281 | !hgrant5_p & v134d285;
assign v1214fee = hmaster2_p & v1215bae | !hmaster2_p & v12153b7;
assign v1668dbe = hgrant5_p & v845542 | !hgrant5_p & !v1668d3d;
assign v14453e4 = hbusreq2_p & v1446224 | !hbusreq2_p & v14453e2;
assign d2f995 = hmaster0_p & d2f990 | !hmaster0_p & d2f994;
assign d306e4 = hmaster0_p & d306d9 | !hmaster0_p & d306e3;
assign v1388ce7 = jx2_p & v138949a | !jx2_p & v138a092;
assign v1515824 = hbusreq2 & v1515823 | !hbusreq2 & v15167ed;
assign v1405849 = hbusreq4_p & v14463b1 | !hbusreq4_p & v1405844;
assign v138a324 = stateA1_p & v138a323 | !stateA1_p & a658a5;
assign v134d50a = hgrant1_p & v845542 | !hgrant1_p & v134d509;
assign v1668cab = hmaster1_p & v1668c8a | !hmaster1_p & !v1668ca1;
assign f2f3ab = hgrant2_p & f2f39e | !hgrant2_p & f2f3aa;
assign v12ad644 = hmaster2_p & v12ad4fc | !hmaster2_p & d30690;
assign v121605f = hmaster2_p & v1216049 | !hmaster2_p & v845547;
assign v1215440 = hbusreq2 & v121541b | !hbusreq2 & v121543f;
assign v12ad5a8 = hgrant1_p & v12ad59a | !hgrant1_p & v12ad5a7;
assign v10d4059 = hmaster0_p & v10d4028 | !hmaster0_p & v10d4058;
assign v134cd58 = hbusreq1 & v134cd57 | !hbusreq1 & v134d273;
assign v12ad503 = hmaster0_p & v12ad4f2 | !hmaster0_p & v12ad502;
assign v140584b = hlock0_p & v14463b1 | !hlock0_p & v140584a;
assign v121654a = hgrant1_p & v1216540 | !hgrant1_p & v1216537;
assign v134d22c = hmaster0_p & v134d22b | !hmaster0_p & v134d1e8;
assign v16a1e6b = hmaster1_p & v16a1e63 | !hmaster1_p & v16a2672;
assign v1216065 = hbusreq1 & v1216adc | !hbusreq1 & !v845542;
assign v1445f12 = hmaster1_p & v1445ecd | !hmaster1_p & v1445f09;
assign v1445b6d = hlock2 & v1445b68 | !hlock2 & v1445b6c;
assign v1445fb7 = hmaster2_p & v1445fa6 | !hmaster2_p & v14463a5;
assign v134ce9f = hlock2_p & v134d23d | !hlock2_p & v134ce9e;
assign v1389461 = hlock2_p & v138945f | !hlock2_p & v1389460;
assign a65463 = hbusreq3 & a6545d | !hbusreq3 & !a65461;
assign v12af5a7 = hbusreq1 & v12afe5b | !hbusreq1 & v12af5a6;
assign f2f2dc = hmaster1_p & f2f2cc | !hmaster1_p & f2f2db;
assign a6590b = hmaster0_p & a658ee | !hmaster0_p & a658f1;
assign v121653c = hbusreq5_p & v121653b | !hbusreq5_p & v845542;
assign v138a450 = hmaster0_p & v138a344 | !hmaster0_p & v138a34f;
assign a65669 = hgrant5_p & v845558 | !hgrant5_p & !a65630;
assign d301b6 = hbusreq3 & d301b1 | !hbusreq3 & d308f7;
assign a65400 = hbusreq5_p & a653fe | !hbusreq5_p & a653ff;
assign v16a223b = hgrant0_p & v845542 | !hgrant0_p & !v16a223a;
assign v1552d4d = hmaster1_p & v1553385 | !hmaster1_p & v1552d4c;
assign d2fea0 = hbusreq5_p & d2fe9e | !hbusreq5_p & d2fe9f;
assign v12afdaf = hmaster2_p & v845542 | !hmaster2_p & v12afdae;
assign v144589b = hbusreq1 & v1445899 | !hbusreq1 & v144589a;
assign v134ce82 = hgrant1_p & v134ce81 | !hgrant1_p & v134d1e8;
assign v85e70d = stateG3_2_p & v845542 | !stateG3_2_p & v893df7;
assign v1405b65 = hgrant3_p & v1405b3c | !hgrant3_p & v1405b64;
assign v151561a = hburst0 & v1515618 | !hburst0 & v1515619;
assign v121628e = hgrant2_p & v1216186 | !hgrant2_p & v121628a;
assign v12162f8 = hmaster1_p & v12162f7 | !hmaster1_p & v12162f4;
assign v1515726 = hgrant5_p & v10d3ff1 | !hgrant5_p & v1515724;
assign v1216124 = hbusreq1 & v1216123 | !hbusreq1 & v845542;
assign d30269 = hmaster2_p & d30268 | !hmaster2_p & v845542;
assign v15168fd = hgrant2_p & v15168fc | !hgrant2_p & !v845542;
assign v134d1de = hmaster2_p & v845542 | !hmaster2_p & v134d1dd;
assign v1405b2b = hgrant2_p & v1405b11 | !hgrant2_p & v1405b2a;
assign f2f43a = hmaster0_p & f2f42e | !hmaster0_p & f2f439;
assign v134d235 = hbusreq2_p & v134d234 | !hbusreq2_p & v134d22f;
assign v134d3b9 = hbusreq3 & v134d3b7 | !hbusreq3 & v134d3b8;
assign v14466c5 = hbusreq5 & v1446687 | !hbusreq5 & v14466c4;
assign v1214f4e = hmaster0_p & v1215d6d | !hmaster0_p & v1215d6c;
assign v138a3cc = hmaster2_p & v845542 | !hmaster2_p & v1515749;
assign v1216015 = hbusreq1 & v1216014 | !hbusreq1 & v845542;
assign v1405a84 = jx2_p & v85e75b | !jx2_p & v1405a80;
assign v12150a2 = hgrant1_p & v121546d | !hgrant1_p & v12150a1;
assign a65496 = hmaster1_p & a65495 | !hmaster1_p & a65476;
assign v1215759 = hlock0_p & v1215b78 | !hlock0_p & v1215758;
assign v144550f = hbusreq2 & v1445509 | !hbusreq2 & v144550e;
assign v12ad5c8 = hbusreq1 & v12ad4d4 | !hbusreq1 & v12ad4e4;
assign v1446062 = hgrant1_p & v1445fd7 | !hgrant1_p & v1446061;
assign v16a193e = hgrant0_p & v845542 | !hgrant0_p & v16a193d;
assign v14461c5 = hmaster1_p & v1446187 | !hmaster1_p & v1445ffc;
assign v1216702 = hbusreq5_p & v1216701 | !hbusreq5_p & v16a2243;
assign d2fc66 = hgrant4_p & d2fbf4 | !hgrant4_p & d2fc53;
assign v16a137a = hgrant2_p & v16a2062 | !hgrant2_p & v16a1379;
assign d30857 = hbusreq5_p & d30705 | !hbusreq5_p & d30856;
assign d30820 = hgrant5_p & d3070d | !hgrant5_p & !d307a8;
assign a6585e = hmaster2_p & a65852 | !hmaster2_p & a6585d;
assign v1215019 = hmaster2_p & v1215bac | !hmaster2_p & !v1214ff0;
assign v16a1a87 = hgrant2_p & v845542 | !hgrant2_p & !v16a1a86;
assign v1446073 = hmaster0_p & v1446055 | !hmaster0_p & v1446072;
assign d2fbf1 = hbusreq5_p & d2fbe4 | !hbusreq5_p & d2fbf0;
assign v10d40b0 = hmaster0_p & v10d3feb | !hmaster0_p & v10d3fda;
assign v1445822 = hgrant2_p & v1445820 | !hgrant2_p & v1445821;
assign v14463c1 = hlock0 & v14463c0 | !hlock0 & v14463bd;
assign v1215c89 = hgrant5_p & v1668da6 | !hgrant5_p & v1215c88;
assign v1445855 = hmaster1_p & v144580a | !hmaster1_p & v1445f09;
assign v121501f = hmaster1_p & v121501e | !hmaster1_p & v1215016;
assign v1389169 = hready_p & v138981d | !hready_p & v1389168;
assign v16a1ce4 = hbusreq2_p & v16a1b68 | !hbusreq2_p & v16a1ce3;
assign v16a1324 = hgrant0_p & v16a131b | !hgrant0_p & !v16a1323;
assign v14463de = hbusreq0 & v14463dd | !hbusreq0 & v14463a8;
assign v144632a = hmaster1_p & v14465b7 | !hmaster1_p & v1446329;
assign d306d1 = hmaster2_p & d306cb | !hmaster2_p & d306d0;
assign v134d464 = hbusreq3 & v134d463 | !hbusreq3 & v134d276;
assign v134cee1 = hbusreq2 & v134cee0 | !hbusreq2 & v134d276;
assign d30270 = hgrant5_p & v845542 | !hgrant5_p & !d3026e;
assign v134ce95 = hlock3 & v134ce88 | !hlock3 & v134ce94;
assign v1553060 = hmaster1_p & v1553385 | !hmaster1_p & v155305f;
assign v134d45f = hmaster0_p & v134d440 | !hmaster0_p & v845542;
assign v144666a = hmaster0_p & v14465e4 | !hmaster0_p & v1446617;
assign v134d397 = hbusreq5_p & v134d396 | !hbusreq5_p & v134d38b;
assign d302e8 = hbusreq5_p & d302e2 | !hbusreq5_p & !d306b2;
assign d307dd = hgrant5_p & d306e3 | !hgrant5_p & d307dc;
assign v16a1d37 = hready_p & v845555 | !hready_p & v16a1d36;
assign v1515828 = hbusreq2_p & v1515827 | !hbusreq2_p & v845542;
assign v10d4009 = hbusreq2_p & v10d4006 | !hbusreq2_p & v10d4008;
assign v155298b = hready_p & v1553306 | !hready_p & v1552d97;
assign bf1f8c = hready_p & bf1f8b | !hready_p & !bf1f56;
assign v1553050 = hbusreq1_p & v1553217 | !hbusreq1_p & v155304f;
assign v1215d83 = hgrant2_p & v1215d7d | !hgrant2_p & v1215d82;
assign v121577f = hmaster0_p & v1215730 | !hmaster0_p & v121577e;
assign locked = d2fd4f;
assign v1216077 = hmaster1_p & v1216068 | !hmaster1_p & v121605d;
assign v1214c1b = hmaster1_p & v1214c05 | !hmaster1_p & v1214bcf;
assign v1445f38 = hlock2 & v1445f34 | !hlock2 & v1445f37;
assign v134d455 = hlock2 & v134d3b5 | !hlock2 & v134d451;
assign v16a1a24 = hmaster1_p & v16a19d3 | !hmaster1_p & !v16a1f96;
assign v12ad516 = hmaster2_p & v12ad514 | !hmaster2_p & !v12ad515;
assign v121630e = hmaster1_p & v121630d | !hmaster1_p & v12162f4;
assign v12162cc = hbusreq2_p & v12162cb | !hbusreq2_p & v12162c5;
assign v1216055 = hbusreq1_p & v1216054 | !hbusreq1_p & v845542;
assign v14458f9 = hmaster2_p & v14458f8 | !hmaster2_p & v1446429;
assign f2f2e0 = hbusreq2_p & f2f2dc | !hbusreq2_p & f2f2df;
assign v1445e82 = stateG10_5_p & v1445e7d | !stateG10_5_p & v1445e81;
assign d2fce6 = hbusreq1_p & d305ef | !hbusreq1_p & d305f0;
assign v1446432 = hbusreq1 & v1446430 | !hbusreq1 & v1446431;
assign v1446674 = hmaster1_p & v1446673 | !hmaster1_p & v144666a;
assign v11e5942 = hmaster1_p & v11e5941 | !hmaster1_p & v845542;
assign v144603c = hbusreq1_p & v144603b | !hbusreq1_p & v144639c;
assign v16a1e54 = hbusreq2 & v16a1e51 | !hbusreq2 & v16a1e53;
assign v16a1e78 = hbusreq2 & v16a1e75 | !hbusreq2 & v16a1e77;
assign v1668c3a = hbusreq3_p & v1668c38 | !hbusreq3_p & !v1668c39;
assign v151621b = hgrant3_p & v1516217 | !hgrant3_p & !v151621a;
assign v12ad620 = hgrant2_p & v12ad5e7 | !hgrant2_p & v12ad61f;
assign v1515603 = hbusreq2 & v15155f6 | !hbusreq2 & v1515602;
assign v12acfb9 = hmaster0_p & v12acfb2 | !hmaster0_p & v12acfb8;
assign v1215fe6 = hgrant3_p & v12167a0 | !hgrant3_p & v1215fe5;
assign v1214bc9 = hbusreq3 & v1214bbc | !hbusreq3 & v1214bc8;
assign d306b2 = hgrant5_p & v845542 | !hgrant5_p & !d306b1;
assign v11e5967 = hgrant4_p & v845542 | !hgrant4_p & !v11e5966;
assign d305e2 = hmaster0_p & d305e1 | !hmaster0_p & d305d7;
assign f2f519 = hmaster2_p & f2f228 | !hmaster2_p & f2f230;
assign v1668c8c = hmaster1_p & v1668c8a | !hmaster1_p & v1668c72;
assign v12153d6 = hbusreq4 & v1216aea | !hbusreq4 & v12153d5;
assign v10d4002 = decide_p & v10d4001 | !decide_p & v10d3fee;
assign v138a3a1 = hmaster0_p & v138a34f | !hmaster0_p & v138a32d;
assign d302d3 = hgrant3_p & d301ba | !hgrant3_p & d302d2;
assign a658d5 = hbusreq0_p & a658d4 | !hbusreq0_p & !a658c6;
assign v1216a93 = hbusreq1_p & v16a1bc6 | !hbusreq1_p & v845570;
assign v15530b6 = hbusreq3_p & v15530a8 | !hbusreq3_p & v15530b5;
assign a6591b = hbusreq2_p & a65917 | !hbusreq2_p & a65919;
assign bf1f65 = hbusreq5_p & bf1f64 | !hbusreq5_p & bf1f63;
assign v1445ae4 = hbusreq5 & v1445ae2 | !hbusreq5 & v1445ae3;
assign v1214eca = hbusreq5_p & v1214ec8 | !hbusreq5_p & v1214ec9;
assign v1445f78 = hbusreq2_p & v1445f71 | !hbusreq2_p & v1445f77;
assign f2f285 = hbusreq1_p & f2f233 | !hbusreq1_p & !v845542;
assign d3080c = hmaster0_p & d306d0 | !hmaster0_p & d3080b;
assign v1215c3d = hmaster2_p & v1215bf1 | !hmaster2_p & v1215c15;
assign a653ff = hgrant5_p & a653f9 | !hgrant5_p & a653fd;
assign v144633d = hbusreq0 & v144633c | !hbusreq0 & v14462f3;
assign v16a1a2c = hbusreq2_p & v16a188d | !hbusreq2_p & v16a1a2b;
assign v1215408 = hlock2_p & v1215407 | !hlock2_p & v12153fc;
assign v14466ee = hlock5 & v14466d3 | !hlock5 & v14466ed;
assign v10d426a = hgrant4_p & v10d401a | !hgrant4_p & v10d4269;
assign v10d403d = hbusreq5_p & v10d4037 | !hbusreq5_p & !v10d403c;
assign v14466e7 = hbusreq2_p & v14466e2 | !hbusreq2_p & v14466e6;
assign d3085e = hmaster0_p & d3085d | !hmaster0_p & d3085b;
assign d301c9 = hmaster2_p & d30700 | !hmaster2_p & d30703;
assign v1446177 = hmaster0_p & v1445fe1 | !hmaster0_p & v1446077;
assign bf1f87 = hgrant2_p & bf1f76 | !hgrant2_p & bf1f86;
assign v1216534 = hgrant0_p & v845542 | !hgrant0_p & !v1216528;
assign v1446687 = hbusreq3 & v1446685 | !hbusreq3 & v1446686;
assign v1214e0b = hbusreq1_p & v1216aeb | !hbusreq1_p & v1216aec;
assign d302f3 = hbusreq2_p & d302e6 | !hbusreq2_p & d302e5;
assign v12ad0b0 = hbusreq1_p & v12afda6 | !hbusreq1_p & v12afda7;
assign d30859 = hmaster1_p & d30851 | !hmaster1_p & !d30858;
assign v12153dc = hbusreq1_p & v12153db | !hbusreq1_p & v1215b97;
assign v134d501 = hlock0_p & v134d273 | !hlock0_p & v134d500;
assign v1446604 = hmaster2_p & v14465f5 | !hmaster2_p & v1446603;
assign d30628 = hbusreq5_p & v845542 | !hbusreq5_p & v84554e;
assign d30167 = hmaster1_p & d30166 | !hmaster1_p & !d2fea2;
assign v14457dd = hmaster0_p & v14457d7 | !hmaster0_p & v1445eb0;
assign a65638 = hmaster2_p & a65623 | !hmaster2_p & a65637;
assign d2fc06 = hmaster0_p & d2fb51 | !hmaster0_p & d2fc05;
assign d30158 = hbusreq5_p & d30157 | !hbusreq5_p & d30156;
assign v16a13ca = hbusreq2_p & v16a13c9 | !hbusreq2_p & !v16a1d0e;
assign f2f44b = hbusreq5_p & f2f3c0 | !hbusreq5_p & !f2f44a;
assign v121652c = hgrant0_p & v1216525 | !hgrant0_p & v845542;
assign d2fbb1 = hmaster1_p & d2fbb0 | !hmaster1_p & d2fb7b;
assign d2fd21 = hgrant5_p & v845542 | !hgrant5_p & !d2fd1f;
assign d30845 = decide_p & d30844 | !decide_p & v845570;
assign d305ea = hmastlock_p & d305e9 | !hmastlock_p & !v845542;
assign v1446119 = hmaster1_p & v1446118 | !hmaster1_p & v1445fde;
assign a658ad = hmastlock_p & a658ac | !hmastlock_p & !v845542;
assign v121578b = hbusreq2 & v1215782 | !hbusreq2 & v121578a;
assign v14453ab = hgrant2_p & v1445383 | !hgrant2_p & v14453aa;
assign v144620a = hbusreq3_p & v14460e3 | !hbusreq3_p & v1446209;
assign v10d42a7 = hmaster1_p & v10d42a6 | !hmaster1_p & !v10d42a1;
assign v1405aa8 = hlock5_p & v1405aa6 | !hlock5_p & !v1405aa7;
assign v14461e1 = hgrant2_p & v144619c | !hgrant2_p & v14461e0;
assign v1214ee4 = hbusreq0 & v1214ede | !hbusreq0 & v1214ee3;
assign v1405a85 = stateA1_p & v845542 | !stateA1_p & v845582;
assign v1216229 = hmaster1_p & v1216228 | !hmaster1_p & v12160e0;
assign v1215ceb = hbusreq0 & v1215ce8 | !hbusreq0 & v1215cea;
assign v121505e = hgrant2_p & v1215059 | !hgrant2_p & v121505d;
assign v16a1330 = hmaster1_p & v16a132f | !hmaster1_p & !v16a2672;
assign d30693 = hbusreq5_p & d30605 | !hbusreq5_p & d30691;
assign d2fd24 = hmaster0_p & d2fd1e | !hmaster0_p & d2fd23;
assign v16a1c01 = hgrant2_p & v845542 | !hgrant2_p & !v16a1c00;
assign v1405b25 = hgrant4_p & v1405ac6 | !hgrant4_p & !v1405b04;
assign v1214d42 = hbusreq1_p & v121539c | !hbusreq1_p & v1214d41;
assign v1214bd1 = hmaster1_p & v12153ac | !hmaster1_p & v1214bcf;
assign v1215c7e = hbusreq1_p & v1216a5a | !hbusreq1_p & v845570;
assign v1668dae = hgrant2_p & v1668dad | !hgrant2_p & !v1668da3;
assign v151584d = hbusreq2_p & v151584c | !hbusreq2_p & !v845542;
assign v12afe3c = hmaster0_p & v845542 | !hmaster0_p & v12afe3b;
assign v1668ca6 = hgrant2_p & v1668ca2 | !hgrant2_p & v1668ca5;
assign v1445480 = hmaster1_p & v144547f | !hmaster1_p & v144627e;
assign v1668d4b = hbusreq1_p & v1668d35 | !hbusreq1_p & v1668d4a;
assign v14461ee = hgrant2_p & v14461c2 | !hgrant2_p & v14461ed;
assign v10d400c = hmaster0_p & v10d400a | !hmaster0_p & v10d400b;
assign v1214bda = hmaster1_p & v1214bbf | !hmaster1_p & v1214bcf;
assign v1215083 = hbusreq2_p & v1215082 | !hbusreq2_p & v121507f;
assign v134cd8d = decide_p & v134d3fa | !decide_p & v134cd8c;
assign v1668cfb = hmaster2_p & v1668cc4 | !hmaster2_p & !v1668cc6;
assign v14460fb = hbusreq2_p & v14460f6 | !hbusreq2_p & v14460fa;
assign v12afdb4 = hmaster0_p & v845542 | !hmaster0_p & v12afdb3;
assign v1214bba = hlock2_p & v1214bb6 | !hlock2_p & v1214bb9;
assign bf1f6d = hlock5_p & bf1f6b | !hlock5_p & !bf1f6c;
assign v1553103 = hlock5 & v155321a | !hlock5 & v1553102;
assign v1216247 = hbusreq3 & v121623b | !hbusreq3 & v1216246;
assign v1215079 = hgrant5_p & v1215077 | !hgrant5_p & !v1215078;
assign v1215d98 = hmaster2_p & v845570 | !hmaster2_p & v12166d2;
assign v1214c51 = hgrant1_p & v1214c4f | !hgrant1_p & v1214c50;
assign v121537b = hbusreq0 & v121537a | !hbusreq0 & v845542;
assign v12aecda = decide_p & v12aeb83 | !decide_p & v12afe76;
assign v1405aff = hmaster2_p & v1405a87 | !hmaster2_p & v1405afc;
assign f2f417 = hmaster1_p & f2f416 | !hmaster1_p & f2f2a2;
assign d307a6 = hbusreq0 & d3079b | !hbusreq0 & d307a5;
assign v14465ae = locked_p & v14465ad | !locked_p & v144639c;
assign v15157d4 = hgrant2_p & v15167ff | !hgrant2_p & !v15157d3;
assign d30146 = hgrant5_p & v84555a | !hgrant5_p & d300ff;
assign v155342d = hmaster1_p & v155342c | !hmaster1_p & v155314e;
assign v12ad018 = hmaster1_p & v12ad008 | !hmaster1_p & v12ad017;
assign v121602b = hmaster1_p & v121602a | !hmaster1_p & !v1216027;
assign v1405844 = hmastlock_p & v1405843 | !hmastlock_p & !v845542;
assign v1389450 = hlock2_p & v138944a | !hlock2_p & v138944f;
assign v1446461 = hmaster1_p & v1446460 | !hmaster1_p & v845542;
assign v1445a1a = hgrant1_p & v14458f8 | !hgrant1_p & v1445a19;
assign v1553387 = stateA1_p & v155313f | !stateA1_p & v155313e;
assign a65615 = hmaster0_p & a65401 | !hmaster0_p & a6538f;
assign v138a337 = hbusreq1_p & v138a336 | !hbusreq1_p & !v845542;
assign d2fd2f = hbusreq5 & d2fd29 | !hbusreq5 & d2fd2e;
assign v10d4281 = hbusreq0_p & v10d4280 | !hbusreq0_p & v10d3fd4;
assign v1445a1f = hgrant5_p & v14458fa | !hgrant5_p & v1445a1e;
assign v1446051 = stateG10_5_p & v1446041 | !stateG10_5_p & v1446050;
assign v121626e = hmaster1_p & v121626d | !hmaster1_p & !v1216027;
assign d30865 = hbusreq5_p & d3072e | !hbusreq5_p & d30864;
assign v134d27b = hlock2_p & v134d27a | !hlock2_p & v845542;
assign bf1f4d = hmaster2_p & v845542 | !hmaster2_p & !v845570;
assign v12af5af = hmaster1_p & v12afe47 | !hmaster1_p & v12af5ae;
assign f2f445 = hgrant5_p & v84554c | !hgrant5_p & f2f41f;
assign v144539c = hmaster1_p & v1445370 | !hmaster1_p & v144591b;
assign v16a12e4 = decide_p & v16a12c7 | !decide_p & v16a2065;
assign v1214d51 = hmaster0_p & v12153ab | !hmaster0_p & v1214d50;
assign v1445805 = hmaster0_p & v1445ecc | !hmaster0_p & v14465b7;
assign v155313f = stateG2_p & v845542 | !stateG2_p & v155313e;
assign d306c0 = hmaster1_p & d306bc | !hmaster1_p & d306bf;
assign v1389fb4 = hbusreq5 & v1389f87 | !hbusreq5 & v1389fb3;
assign d2fc89 = hmaster1_p & d2fc88 | !hmaster1_p & v845570;
assign v1668e08 = hlock3_p & v1668e07 | !hlock3_p & v845542;
assign d3068b = hbusreq5_p & d3060b | !hbusreq5_p & d3068a;
assign v144655d = hgrant0_p & v1446398 | !hgrant0_p & v845542;
assign v1405871 = hmaster2_p & v1405860 | !hmaster2_p & v14463b1;
assign v131be8a = hbusreq5_p & v845542 | !hbusreq5_p & v84557c;
assign bf1f71 = hgrant2_p & bf1f5a | !hgrant2_p & bf1f70;
assign v1515617 = hmaster1_p & v151560c | !hmaster1_p & v1515616;
assign v1216562 = hmaster2_p & v121655f | !hmaster2_p & v1216561;
assign v144609d = hmaster1_p & v144609c | !hmaster1_p & v1445fef;
assign v1552d80 = hgrant5_p & v1553225 | !hgrant5_p & v1552d7f;
assign f2f403 = hbusreq3 & f2f3f8 | !hbusreq3 & f2f402;
assign v1445df2 = hbusreq1 & v1445de9 | !hbusreq1 & v1445df1;
assign v16a1bd1 = hbusreq0 & v16a207a | !hbusreq0 & v16a1bd0;
assign v12160d9 = hmaster2_p & v12160d8 | !hmaster2_p & v845542;
assign v1445a99 = hbusreq0 & v1445a97 | !hbusreq0 & v1445a7f;
assign d2f9b9 = hmaster0_p & d2fec8 | !hmaster0_p & d2f9b8;
assign v1445f1e = decide_p & v1445de1 | !decide_p & v1445f1d;
assign v14457ea = hgrant2_p & v14457e3 | !hgrant2_p & v14457e9;
assign bf1f78 = hgrant4_p & bf1f52 | !hgrant4_p & bf1f77;
assign v10d4065 = hbusreq1_p & v10d3fd9 | !hbusreq1_p & !v10d3fdf;
assign v1668d89 = hbusreq5_p & v1668d87 | !hbusreq5_p & v1668d88;
assign d3011c = hlock5_p & d3011a | !hlock5_p & !d3011b;
assign v1214d2a = hbusreq0 & v1214d0c | !hbusreq0 & v1216718;
assign v1445b10 = hbusreq2_p & v1445b0e | !hbusreq2_p & v1445b0f;
assign v134d529 = hlock5 & v134d524 | !hlock5 & v134d528;
assign v134d4a4 = hbusreq2_p & v134d49c | !hbusreq2_p & v134d4a3;
assign v16a1d3f = hbusreq0 & v16a1d3b | !hbusreq0 & v16a1d3e;
assign v15157e5 = hmaster0_p & v15157dd | !hmaster0_p & v15157e4;
assign v1215cc3 = hmaster2_p & v1215cc1 | !hmaster2_p & v1215cc2;
assign v14462f8 = hgrant5_p & v1446433 | !hgrant5_p & v1446621;
assign d308e2 = hbusreq1 & v845542 | !hbusreq1 & d308e1;
assign v12150fc = hlock2_p & v12150fa | !hlock2_p & v12150fb;
assign d3089c = hbusreq5_p & d307ab | !hbusreq5_p & d3089b;
assign a65b20 = decide_p & a65aff | !decide_p & a662a2;
assign v12160b3 = hmaster0_p & v121606b | !hmaster0_p & v1216068;
assign v12150b6 = hmaster1_p & v12150b5 | !hmaster1_p & !v1215ba1;
assign v1445f7e = hbusreq3 & v1445f7c | !hbusreq3 & v1445f7d;
assign d3029e = decide_p & d3029d | !decide_p & v845570;
assign v12ad57c = hmaster1_p & v12ad57b | !hmaster1_p & !v12ad525;
assign v155350e = hmaster0_p & v15534ef | !hmaster0_p & v845542;
assign v1446418 = hbusreq0 & v1446414 | !hbusreq0 & v1446417;
assign d8078e = hgrant5_p & d80770 | !hgrant5_p & !d8078d;
assign v16a1dbb = hready_p & v16a1dba | !hready_p & v16a1dae;
assign bf1f97 = hgrant5_p & bf1f62 | !hgrant5_p & bf1f96;
assign f2e4fd = hgrant2_p & v845542 | !hgrant2_p & f2e4fc;
assign v1216a66 = hmastlock_p & v1216a65 | !hmastlock_p & v845542;
assign v1446168 = hmaster1_p & v1446081 | !hmaster1_p & v1446073;
assign v10d42d6 = decide_p & v10d42cf | !decide_p & v10d42d5;
assign d2fbba = hmaster1_p & d2fbb0 | !hmaster1_p & d2fb9d;
assign v10d40c6 = hgrant2_p & v10d40b9 | !hgrant2_p & !v10d40c5;
assign v14465a9 = decide_p & v1446556 | !decide_p & v1446564;
assign v1215446 = hlock2_p & v1215444 | !hlock2_p & v1215445;
assign v1445b5d = hbusreq0 & v1445b5c | !hbusreq0 & v14462f3;
assign v1216189 = hgrant2_p & v1216186 | !hgrant2_p & v121617f;
assign d300cb = hbusreq4_p & d300ca | !hbusreq4_p & v845542;
assign d30733 = hlock1_p & v845542 | !hlock1_p & !v16693aa;
assign v16a2091 = hbusreq0 & v16a207a | !hbusreq0 & v16a2090;
assign d3071b = hbusreq1_p & d3071a | !hbusreq1_p & v845542;
assign v1445d96 = hbusreq0_p & v14463b1 | !hbusreq0_p & !v1445d7f;
assign v1445354 = hbusreq2_p & v1445b4d | !hbusreq2_p & v1445353;
assign v1214d49 = hbusreq5_p & v12153a7 | !hbusreq5_p & v1214d48;
assign v134d427 = hgrant1_p & v845542 | !hgrant1_p & v134d426;
assign a6539a = hbusreq1 & a65395 | !hbusreq1 & a65399;
assign d300e1 = hgrant5_p & d300d4 | !hgrant5_p & d300e0;
assign bf1f9a = hbusreq1_p & bf1f66 | !hbusreq1_p & bf1f99;
assign v1445e72 = hlock1 & v1445e68 | !hlock1 & v1445e60;
assign v1552f6b = hgrant2_p & v1553380 | !hgrant2_p & v1552f6a;
assign v1446472 = hmaster2_p & v845542 | !hmaster2_p & v1446471;
assign d2fd1f = hmaster2_p & d30648 | !hmaster2_p & v845542;
assign v14463a3 = hbusreq1_p & v144639c | !hbusreq1_p & v14463a2;
assign v15157b3 = hbusreq0 & v15157ad | !hbusreq0 & v15157b2;
assign v121535d = hbusreq0_p & v1216a77 | !hbusreq0_p & v845542;
assign d2fbd8 = hgrant5_p & v84554a | !hgrant5_p & d2fbd6;
assign d2fc49 = hbusreq0_p & d30645 | !hbusreq0_p & v845542;
assign v1446018 = hmaster1_p & v1446466 | !hmaster1_p & v1446017;
assign v1216001 = hlock1_p & v1215ffe | !hlock1_p & v1216000;
assign v14460cb = hgrant5_p & v14460ca | !hgrant5_p & v14460b1;
assign v1445add = hlock2 & v1445abf | !hlock2 & v1445adb;
assign v16a2075 = hgrant4_p & v845559 | !hgrant4_p & v16a2074;
assign v15530b5 = hgrant3_p & v15530b2 | !hgrant3_p & v15530b4;
assign v1446186 = hgrant2_p & v1446183 | !hgrant2_p & v1446185;
assign v12150ec = hmaster2_p & v12150c4 | !hmaster2_p & v12150c7;
assign v16a13f3 = hgrant5_p & v845542 | !hgrant5_p & !v16a2086;
assign v121608e = hlock2_p & v121608c | !hlock2_p & v121608d;
assign v1216157 = hmaster2_p & v1216143 | !hmaster2_p & v1216156;
assign v1446208 = hready_p & v1446038 | !hready_p & v1446203;
assign d30282 = hbusreq0 & d3027d | !hbusreq0 & d30281;
assign v1445f59 = hlock2 & v1445f53 | !hlock2 & v1445f58;
assign v14453a0 = hbusreq2 & v144539b | !hbusreq2 & v144539f;
assign v1284cb9 = hmaster2_p & v140587c | !hmaster2_p & !v1284c8f;
assign v1553055 = hbusreq0_p & v1553399 | !hbusreq0_p & v1553217;
assign v16a1afa = hready & v16a1af9 | !hready & v845542;
assign v1214ece = hbusreq0 & v1214eca | !hbusreq0 & v1214ecd;
assign v1445e6e = hgrant5_p & v1445e54 | !hgrant5_p & v1445e6d;
assign a653ea = hmaster2_p & a65360 | !hmaster2_p & !a65395;
assign v1405b44 = hgrant2_p & v1405b41 | !hgrant2_p & v1405b43;
assign v16a1bf0 = hgrant1_p & v84554d | !hgrant1_p & v16a1bef;
assign v12ad511 = hburst1 & v12ad510 | !hburst1 & v138a326;
assign v144545f = hlock5 & v1445446 | !hlock5 & v144545d;
assign v1445aef = hmaster1_p & v1445aee | !hmaster1_p & v144590e;
assign v151577a = hgrant4_p & v1515765 | !hgrant4_p & v1515779;
assign v144612c = hbusreq2_p & v1446129 | !hbusreq2_p & v144612b;
assign v121603c = hbusreq1 & v1216a96 | !hbusreq1 & v845542;
assign v155351b = hbusreq3_p & v155350d | !hbusreq3_p & v155351a;
assign v1552f8d = hgrant3_p & v155321c | !hgrant3_p & v1552f8c;
assign v1215731 = hmaster2_p & v1215b7b | !hmaster2_p & v1215b81;
assign a65911 = hbusreq3 & a658f9 | !hbusreq3 & a65910;
assign v151579b = hgrant1_p & f2f281 | !hgrant1_p & v151579a;
assign v1284d62 = hbusreq2_p & v1284d5f | !hbusreq2_p & v1284d61;
assign d30774 = hbusreq2_p & d30773 | !hbusreq2_p & d30772;
assign v138a43c = hbusreq5_p & v138a312 | !hbusreq5_p & v845542;
assign v1668d0b = hmaster1_p & v1668cf1 | !hmaster1_p & !v1668cfd;
assign d80745 = hmaster2_p & d80743 | !hmaster2_p & d80744;
assign v1405ab0 = hmaster2_p & v1405aa2 | !hmaster2_p & !v845542;
assign v1216150 = hbusreq4_p & v121614f | !hbusreq4_p & !v845542;
assign v144545e = hlock5 & v1445452 | !hlock5 & v144545d;
assign v1215c1c = hgrant5_p & v1215c07 | !hgrant5_p & v1215c1b;
assign v1215751 = hmaster2_p & v1215750 | !hmaster2_p & v121574b;
assign v1214ffe = hgrant1_p & v1215bac | !hgrant1_p & v1214ff5;
assign v16a1d49 = hgrant5_p & v845542 | !hgrant5_p & v16a1d48;
assign v15533b5 = hlock0 & v15533a9 | !hlock0 & v15533b4;
assign v144618a = hmaster1_p & v1446189 | !hmaster1_p & v1446073;
assign v16a1d51 = hbusreq2 & v16a1d4d | !hbusreq2 & !v16a1d50;
assign v1214bf7 = hbusreq3 & v1214bd8 | !hbusreq3 & v1214bf6;
assign f2eda5 = jx1_p & f2f462 | !jx1_p & f2eda4;
assign a65367 = hburst1 & a65366 | !hburst1 & v845542;
assign v12ad0b9 = hbusreq0 & v12afda2 | !hbusreq0 & v12ad0b8;
assign v1215bf7 = hmaster2_p & v1215bf6 | !hmaster2_p & v845542;
assign v1215cde = hbusreq2_p & v1215cdd | !hbusreq2_p & !v1215cd7;
assign d3013e = hbusreq5_p & d3013c | !hbusreq5_p & d3013d;
assign v15155ee = hbusreq2 & v151697c | !hbusreq2 & v15155ed;
assign v1552d9d = hready_p & v1552d9c | !hready_p & v1552d74;
assign v138a366 = hbusreq3 & v138a358 | !hbusreq3 & v138a365;
assign f2f382 = hbusreq1_p & f2f381 | !hbusreq1_p & v845542;
assign v16a1e94 = hbusreq4_p & v845572 | !hbusreq4_p & v16a1e93;
assign v14453af = hbusreq2_p & v14453a6 | !hbusreq2_p & v14453ae;
assign v15530a3 = hlock5 & v1553094 | !hlock5 & v15530a2;
assign v1216aee = hgrant4_p & v1216aed | !hgrant4_p & v1216aeb;
assign d2fadf = hbusreq4_p & d300db | !hbusreq4_p & d306a3;
assign v12153a0 = hlock5_p & v121539e | !hlock5_p & v121539f;
assign v15533b6 = hmaster0_p & v1553398 | !hmaster0_p & v15533b5;
assign v16a1b66 = hbusreq2 & v16a1b64 | !hbusreq2 & v16a1b65;
assign v16a1949 = hgrant0_p & v845542 | !hgrant0_p & !v16a1948;
assign v1446561 = hgrant5_p & v845542 | !hgrant5_p & v1446560;
assign v15167f6 = hbusreq2_p & v15167f5 | !hbusreq2_p & !v845542;
assign v134ce33 = hbusreq0_p & v134d370 | !hbusreq0_p & v134d273;
assign v1445b82 = hbusreq2_p & v1445b7c | !hbusreq2_p & v1445b81;
assign v1214cd6 = hgrant5_p & v1215386 | !hgrant5_p & v1214cd5;
assign a656b2 = hbusreq5 & a6569a | !hbusreq5 & a656b1;
assign v1214d09 = hmaster0_p & v1214c2e | !hmaster0_p & v1214d08;
assign f2f2ea = hmaster1_p & f2f2e9 | !hmaster1_p & f2f2db;
assign f2f38f = hgrant5_p & f2f2a1 | !hgrant5_p & !f2f38e;
assign v134d4a7 = hbusreq2 & v134d4a5 | !hbusreq2 & v134d4a6;
assign v1445366 = hmaster0_p & v1445a5a | !hmaster0_p & v1445a43;
assign d30894 = hbusreq5_p & d30802 | !hbusreq5_p & !d30893;
assign v144642c = hmaster2_p & v144641d | !hmaster2_p & v1446423;
assign v14460c3 = hgrant2_p & v14460c2 | !hgrant2_p & v14460be;
assign v144554a = decide_p & v144553f | !decide_p & v1445549;
assign v144644a = hmaster1_p & v1446449 | !hmaster1_p & v1446436;
assign v134ce36 = hbusreq1 & v134ce35 | !hbusreq1 & v134d273;
assign d30164 = hready_p & d30163 | !hready_p & d2ff0c;
assign v11e5972 = hready_p & v11e5971 | !hready_p & !v845542;
assign v12ad550 = hmaster1_p & v12ad517 | !hmaster1_p & v12ad54f;
assign v134d4e0 = hmaster0_p & v845542 | !hmaster0_p & v134d4df;
assign v1215cb2 = hgrant5_p & v845542 | !hgrant5_p & !v1215cb0;
assign v134ce92 = hlock2_p & v134ce91 | !hlock2_p & v134ce85;
assign a6564f = hbusreq5_p & a653e3 | !hbusreq5_p & a6564e;
assign v15168ed = hlock2_p & v15168ec | !hlock2_p & !v845542;
assign v134d44f = hmaster0_p & v134d44e | !hmaster0_p & v134d431;
assign f2f28f = hready_p & f2f28e | !hready_p & f2f27e;
assign v138938a = hmaster2_p & v15155f9 | !hmaster2_p & !v845570;
assign v1215367 = hmaster2_p & v1215364 | !hmaster2_p & v1215366;
assign v10d428c = hmaster2_p & v10d4285 | !hmaster2_p & v10d428b;
assign v16a195d = hgrant2_p & v845542 | !hgrant2_p & v16a195c;
assign v12150b9 = hbusreq2_p & v12150b6 | !hbusreq2_p & v12150b8;
assign d300ee = hmaster2_p & d300c4 | !hmaster2_p & d300ed;
assign v16a194f = hbusreq0 & v16a1943 | !hbusreq0 & v16a194e;
assign v151699f = decide_p & v151699e | !decide_p & v845542;
assign d2fb7f = hmaster0_p & d2fb6c | !hmaster0_p & d2fb7e;
assign v1215c76 = hgrant2_p & v1215c4d | !hgrant2_p & v1215c6b;
assign v12165af = hmaster0_p & v121658b | !hmaster0_p & v12165ae;
assign v1445ac8 = hbusreq2_p & v1445ac3 | !hbusreq2_p & v1445ac7;
assign v10d40cb = hmaster0_p & v10d3feb | !hmaster0_p & v10d407f;
assign a65b14 = hmaster0_p & a65b13 | !hmaster0_p & a66287;
assign v16a1f94 = hbusreq3 & v16a2678 | !hbusreq3 & v16a1f93;
assign v12af9d4 = hgrant5_p & d30690 | !hgrant5_p & v12af9d3;
assign v1215d66 = hmaster2_p & v12164cf | !hmaster2_p & v12164d9;
assign v12ad5f2 = hmaster1_p & v12ad5f1 | !hmaster1_p & v12ad4ed;
assign v16a1380 = decide_p & v16a12c7 | !decide_p & v16a137f;
assign v1445545 = hmaster1_p & v14465b7 | !hmaster1_p & v1445544;
assign d2feb3 = hlock4_p & v845542 | !hlock4_p & d305ea;
assign v10d3ffc = hmaster1_p & v10d3ff2 | !hmaster1_p & v10d3ffb;
assign a65858 = hburst1 & a65857 | !hburst1 & v845542;
assign v1445bcc = hmaster1_p & v1445bcb | !hmaster1_p & v1445bb7;
assign v16a1e5d = hbusreq1_p & v845542 | !hbusreq1_p & v16a1e5c;
assign v1216252 = hgrant2_p & v1216234 | !hgrant2_p & v1216251;
assign v15534f6 = hbusreq2 & v15534f4 | !hbusreq2 & v15534f5;
assign v12af9b3 = hbusreq0 & v12af9b1 | !hbusreq0 & v12af9b2;
assign v134d226 = hlock2_p & v134d223 | !hlock2_p & v134d225;
assign v1515719 = hburst1 & v1515718 | !hburst1 & v151564a;
assign v1552f86 = hlock3 & v155341e | !hlock3 & v1552f85;
assign v1553434 = hbusreq3 & v1553433 | !hbusreq3 & v155321a;
assign v16a1404 = hmaster1_p & v16a1403 | !hmaster1_p & v16a1d7a;
assign a65434 = hgrant5_p & a65892 | !hgrant5_p & a653e2;
assign v1405ad6 = hgrant1_p & v1405a86 | !hgrant1_p & v1405ad5;
assign d2f96d = hbusreq4_p & d300d8 | !hbusreq4_p & !v845542;
assign v1214da5 = hbusreq2_p & v1214da0 | !hbusreq2_p & v1214da4;
assign d2ff05 = hbusreq2_p & d2ff04 | !hbusreq2_p & d2ff03;
assign a662a7 = hgrant3_p & a66281 | !hgrant3_p & a662a6;
assign v1445e2e = hlock2 & v1445e2b | !hlock2 & v1445e2d;
assign v12ad4df = hmaster2_p & v12ad4ca | !hmaster2_p & v12ad4d4;
assign v144552b = hmaster1_p & v14454f0 | !hmaster1_p & v1445b8d;
assign v144586f = hlock0_p & v144639c | !hlock0_p & v144586e;
assign v121651e = hmaster0_p & v845547 | !hmaster0_p & v121651d;
assign v134ce8e = hbusreq0 & v134ce8d | !hbusreq0 & v134d1e8;
assign d307f4 = hmaster0_p & d307c3 | !hmaster0_p & d307f3;
assign f2f4b9 = hgrant2_p & f2f4b6 | !hgrant2_p & f2f4ac;
assign v1668da6 = hmaster2_p & v845570 | !hmaster2_p & v845542;
assign f2e4cb = hmaster1_p & v845542 | !hmaster1_p & f2e4ca;
assign v138a30a = hmaster0_p & v138a309 | !hmaster0_p & v1668c1f;
assign v1216b14 = hlock2_p & v1216b13 | !hlock2_p & v1216b10;
assign v1446140 = hbusreq3 & v1446133 | !hbusreq3 & v144613f;
assign v1405ac6 = hlock0_p & v845542 | !hlock0_p & v1405ac5;
assign v1445bbb = hbusreq2_p & v1445bb8 | !hbusreq2_p & v1445bba;
assign v1216127 = hmaster2_p & v1216126 | !hmaster2_p & v845542;
assign v16a142c = hbusreq2_p & v16a13e8 | !hbusreq2_p & v16a1db3;
assign v15534d7 = hmaster2_p & v15534d0 | !hmaster2_p & v15534d6;
assign v134cf6b = hready_p & v134d34f | !hready_p & v134cf6a;
assign f2f2b0 = hbusreq3 & f2f2a7 | !hbusreq3 & f2f2af;
assign d30702 = hbusreq0_p & v845542 | !hbusreq0_p & a65861;
assign v144582c = hlock2 & v14457f6 | !hlock2 & v144582b;
assign d2feae = decide_p & d2fead | !decide_p & v845570;
assign v12afe5a = hgrant0_p & v12afe59 | !hgrant0_p & v845542;
assign d2fc21 = hready_p & d2fc1a | !hready_p & d2fbc4;
assign v12ad528 = hbusreq0 & v12ad527 | !hbusreq0 & !v845542;
assign d30829 = hlock5_p & d30827 | !hlock5_p & d30828;
assign v12ad59c = hlock0_p & v1515713 | !hlock0_p & d2fbe5;
assign v12ad5f9 = hmaster0_p & v845542 | !hmaster0_p & v12ad5f8;
assign f2f428 = hmaster2_p & f2f41e | !hmaster2_p & f2f286;
assign v1445e0d = hmaster0_p & v1445de6 | !hmaster0_p & v1445e0c;
assign v16a1bb2 = decide_p & v16a1b6b | !decide_p & !v16a2065;
assign v12160fb = hlock0_p & v1216a5a | !hlock0_p & !v845542;
assign v1389fc0 = hmaster1_p & v845542 | !hmaster1_p & v1389fbf;
assign d306b6 = hmaster0_p & d306ad | !hmaster0_p & d306b5;
assign d30228 = hgrant5_p & d30220 | !hgrant5_p & d30227;
assign v14465d3 = hmaster2_p & v14465b3 | !hmaster2_p & v14465d2;
assign v138a007 = hmaster1_p & v1389ffe | !hmaster1_p & v138a006;
assign v1215463 = hmaster2_p & v121545f | !hmaster2_p & v1215bac;
assign v12152ed = hmaster1_p & v12152ec | !hmaster1_p & !v1215ba1;
assign v1214c76 = hgrant2_p & v1214c44 | !hgrant2_p & v1214c75;
assign f2f412 = hbusreq3 & f2f40a | !hbusreq3 & f2f411;
assign v15168ae = hbusreq1 & v15168ad | !hbusreq1 & !v845542;
assign v1445fa8 = hbusreq0 & v1445fa7 | !hbusreq0 & v1445f85;
assign v134cec0 = hlock3_p & v134cea9 | !hlock3_p & v134cebf;
assign v1216a8b = hmastlock_p & v1216a8a | !hmastlock_p & v845542;
assign v16a1bdc = hmaster1_p & v16a1bce | !hmaster1_p & v16a1bdb;
assign f2f2af = hmaster1_p & f2f2ac | !hmaster1_p & f2f2ae;
assign a662b4 = hbusreq5_p & a6629b | !hbusreq5_p & a662ad;
assign v1216a6d = hmaster0_p & v1216a6a | !hmaster0_p & v1216a6c;
assign v12ad559 = hmaster1_p & v12ad53b | !hmaster1_p & v12ad54f;
assign d30267 = hlock2_p & d30266 | !hlock2_p & !v845542;
assign v1216a81 = hmaster1_p & v1216a80 | !hmaster1_p & v845542;
assign v14459d4 = hmaster2_p & v14459d3 | !hmaster2_p & v14458e5;
assign v138a039 = hlock3_p & v138a011 | !hlock3_p & v138a038;
assign v1214db6 = hmaster1_p & v1214da9 | !hmaster1_p & !v1214d1e;
assign v1516800 = hgrant2_p & v15167ff | !hgrant2_p & !v845542;
assign v134cd86 = hlock2 & v134d3b5 | !hlock2 & v134cd82;
assign v1515669 = hmaster2_p & v1668c6e | !hmaster2_p & !v1515668;
assign d30247 = hgrant5_p & v845542 | !hgrant5_p & d301fa;
assign v134cea6 = hlock3 & v134ce88 | !hlock3 & v134cea5;
assign v166939b = hbusreq4_p & a66295 | !hbusreq4_p & v845570;
assign v16a16b6 = jx2_p & v16a1dbd | !jx2_p & v16a16b5;
assign v134d3ac = hbusreq0 & v134d3ab | !hbusreq0 & v134d274;
assign f2f27e = decide_p & f2f223 | !decide_p & f2f23c;
assign v10d4061 = hgrant4_p & v10d3fdb | !hgrant4_p & v10d4060;
assign v1668c40 = hbusreq1_p & v1668c1c | !hbusreq1_p & !v845542;
assign v1405852 = hbusreq2_p & v140584e | !hbusreq2_p & v1405851;
assign v1445436 = hbusreq2_p & v1445435 | !hbusreq2_p & v144541b;
assign v1515bb0 = hgrant3_p & v1516107 | !hgrant3_p & !v1515baf;
assign v138a460 = hlock2_p & v138a45d | !hlock2_p & v138a45f;
assign d2fb6b = hmaster2_p & d2fb69 | !hmaster2_p & d2fb6a;
assign v1216183 = hmaster1_p & v1216182 | !hmaster1_p & v845542;
assign v1515770 = hbusreq0_p & a653c8 | !hbusreq0_p & !v1515741;
assign v14453c2 = hlock5 & v1445354 | !hlock5 & v14453c1;
assign v1216282 = hmaster0_p & v1216029 | !hmaster0_p & v121601e;
assign v13895a6 = hready_p & v845542 | !hready_p & v13895a5;
assign v1214bf3 = hmaster1_p & v1214bf2 | !hmaster1_p & v1214bcf;
assign v14454f3 = hbusreq2_p & v14454f2 | !hbusreq2_p & v1445bdb;
assign v1214c9e = hgrant2_p & v1214c9d | !hgrant2_p & v1214c93;
assign v15167f9 = hmaster0_p & v1668c1f | !hmaster0_p & v15167f8;
assign v1215067 = hmaster1_p & v1215066 | !hmaster1_p & v1215054;
assign v16a16ad = hgrant2_p & v845542 | !hgrant2_p & v16a16aa;
assign v1445fd4 = hbusreq1_p & v144641f | !hbusreq1_p & v1446427;
assign d30950 = hbusreq1 & d305ea | !hbusreq1 & !d3094f;
assign v14463e7 = hlock1 & v14463b5 | !hlock1 & v14463e6;
assign d2fc2f = hmaster2_p & d2fc2e | !hmaster2_p & v84554a;
assign v1215029 = hgrant4_p & v1215026 | !hgrant4_p & v1215028;
assign a65438 = hbusreq0 & a65433 | !hbusreq0 & a65437;
assign v14463e4 = hbusreq1 & v14463e2 | !hbusreq1 & v14463e3;
assign v1445faf = hmaster1_p & v144639c | !hmaster1_p & v1445fae;
assign v1215411 = hmaster1_p & v12153ef | !hmaster1_p & v121540f;
assign v16a1e21 = hgrant1_p & v845547 | !hgrant1_p & v16a1e20;
assign v134d3fc = hready_p & v134d1e2 | !hready_p & v134d3fb;
assign v1216ace = hbusreq1 & v1216ac7 | !hbusreq1 & !v1216acd;
assign d30872 = hbusreq2_p & d3076e | !hbusreq2_p & d30870;
assign v10d4295 = hgrant1_p & v10d4065 | !hgrant1_p & !v10d4294;
assign v1446332 = hlock0 & v1446331 | !hlock0 & v1446330;
assign v14453fe = hbusreq3 & v14453fc | !hbusreq3 & v14453fd;
assign v143fd7a = hgrant5_p & v845542 | !hgrant5_p & v143fd79;
assign v1215cf3 = hbusreq5_p & v1215cf2 | !hbusreq5_p & !v1215cb6;
assign v16693ad = hmaster0_p & v16693ac | !hmaster0_p & v845542;
assign v14460e3 = hgrant3_p & v144600b | !hgrant3_p & v14460e2;
assign v1284cbe = hmaster1_p & v1284cbd | !hmaster1_p & !v1445bb7;
assign d30287 = hbusreq2_p & d30285 | !hbusreq2_p & !d30286;
assign f2f28d = hbusreq2_p & f2f23a | !hbusreq2_p & f2f28c;
assign v14458aa = hlock0 & v14458a3 | !hlock0 & v14458a1;
assign v12160ef = hgrant0_p & v12160ee | !hgrant0_p & !v1216528;
assign v16a1c03 = hbusreq2 & v16a1c01 | !hbusreq2 & !v16a1c02;
assign v1668d26 = hbusreq4_p & v1668d24 | !hbusreq4_p & v1668d25;
assign v1405ac7 = hmaster2_p & v1405ac4 | !hmaster2_p & v1405ac6;
assign v14453b9 = hbusreq2_p & v14453b3 | !hbusreq2_p & v14453b8;
assign v121570f = hlock0_p & v12160eb | !hlock0_p & !v12160ec;
assign v16a2679 = hmaster0_p & v16a2675 | !hmaster0_p & v16a266a;
assign v1215d02 = hbusreq5_p & v1215d01 | !hbusreq5_p & v1215cd0;
assign d2fad9 = hbusreq4_p & d300bb | !hbusreq4_p & d306a3;
assign v1389fdd = hbusreq5_p & v1389fdc | !hbusreq5_p & !v845542;
assign v14457be = hbusreq2_p & v14457ba | !hbusreq2_p & v14457bd;
assign v12153f6 = hlock2_p & v12153f5 | !hlock2_p & v12153f0;
assign v1214e64 = hlock2_p & v1214e5b | !hlock2_p & !v1214e63;
assign v14463b8 = hmaster2_p & v14463ad | !hmaster2_p & v14463b7;
assign v134d243 = hmaster1_p & v134d242 | !hmaster1_p & v134d208;
assign d2fbe5 = hbusreq0_p & v845570 | !hbusreq0_p & v845542;
assign v12af98d = hmaster0_p & v12af73f | !hmaster0_p & v12af98c;
assign v1445bd9 = hmaster1_p & v1445bd8 | !hmaster1_p & v1445bb7;
assign f2f3aa = hmaster1_p & f2f3a9 | !hmaster1_p & f2f393;
assign v1214fe6 = hgrant1_p & v1215bac | !hgrant1_p & v1214fe5;
assign v1445f81 = decide_p & v14466ef | !decide_p & v1445f80;
assign f2ed91 = hready_p & v845542 | !hready_p & f2ed90;
assign v1445bb6 = hbusreq5_p & v1445fcb | !hbusreq5_p & v1446413;
assign v1215d67 = hbusreq5_p & v1215d65 | !hbusreq5_p & v1215d66;
assign d30722 = hlock1_p & v845542 | !hlock1_p & a66278;
assign v11ac67c = hgrant5_p & v84554c | !hgrant5_p & v11ac602;
assign v15155f0 = hready_p & v845542 | !hready_p & v15155ef;
assign v16a1408 = hbusreq5 & v16a1402 | !hbusreq5 & v16a1407;
assign v16a19a4 = hbusreq4 & v845547 | !hbusreq4 & v845542;
assign v1445da6 = hmaster2_p & v144639c | !hmaster2_p & v1445d88;
assign v12ad508 = hbusreq0 & v12ad507 | !hbusreq0 & !v845542;
assign v14453ef = hlock5 & v14453e9 | !hlock5 & v14453ee;
assign v1216198 = hbusreq0 & v1216193 | !hbusreq0 & v1216197;
assign d300d6 = hbusreq1 & v84555a | !hbusreq1 & !d2fea8;
assign v12153aa = hmaster1_p & v1215396 | !hmaster1_p & v12153a9;
assign v12ad4f5 = hmaster0_p & v12ad4f2 | !hmaster0_p & v12ad4f4;
assign v1668c6f = hmaster2_p & v1668c6e | !hmaster2_p & a658d6;
assign v1515794 = hgrant4_p & a662a9 | !hgrant4_p & v845570;
assign v1552fd1 = hlock5 & v155321a | !hlock5 & v1552fd0;
assign v1668c24 = hmaster1_p & v1668c20 | !hmaster1_p & v1668c23;
assign v1516806 = decide_p & v1516805 | !decide_p & v845576;
assign v151584a = hmaster1_p & v1515849 | !hmaster1_p & v15157f9;
assign v16a1440 = hgrant5_p & v845542 | !hgrant5_p & !v16a1439;
assign v1445416 = hgrant2_p & v1445411 | !hgrant2_p & v1445415;
assign v144626e = hmaster0_p & v144639c | !hmaster0_p & v144626d;
assign d2fc0a = hbusreq2_p & d2fc09 | !hbusreq2_p & d2fc00;
assign v14460d2 = hmaster1_p & v1446082 | !hmaster1_p & v14460cf;
assign v1284d37 = hbusreq0_p & v140588d | !hbusreq0_p & v144639c;
assign v12ad675 = hbusreq1_p & v12ad514 | !hbusreq1_p & v12ad674;
assign v14459c7 = hgrant0_p & v14459bb | !hgrant0_p & v14459c6;
assign v134cee6 = decide_p & v134cedd | !decide_p & v134cee5;
assign d2fb59 = hmaster2_p & d2fb4d | !hmaster2_p & d2fb58;
assign v16a13fc = hbusreq2 & v16a13fb | !hbusreq2 & !v16a209e;
assign d80782 = hgrant5_p & v845542 | !hgrant5_p & d80781;
assign v1215d44 = hgrant2_p & v1215d3e | !hgrant2_p & v1215d43;
assign f2f3ee = decide_p & f2f3ed | !decide_p & v845542;
assign v1214d2f = hbusreq2 & v1214d23 | !hbusreq2 & v1214d2e;
assign v16a1ad8 = hbusreq4_p & v845542 | !hbusreq4_p & v845572;
assign d2fed8 = hmaster0_p & d2fed5 | !hmaster0_p & d2fec8;
assign v144610c = hbusreq2_p & v144610a | !hbusreq2_p & v144610b;
assign v1214ddd = hbusreq3 & v845547 | !hbusreq3 & v1214ddc;
assign d30752 = hlock5_p & d30751 | !hlock5_p & v84554e;
assign d8073f = hmaster2_p & v845542 | !hmaster2_p & !d8073d;
assign v12ad5aa = hbusreq1_p & v12ad5a9 | !hbusreq1_p & v1668d22;
assign v16a1976 = hmaster0_p & v16a1972 | !hmaster0_p & v16a1975;
assign v12ad592 = hbusreq5 & v12ad57f | !hbusreq5 & v12ad591;
assign v121544b = hbusreq2_p & v121544a | !hbusreq2_p & v1215445;
assign d2fb54 = hbusreq0 & d2fb53 | !hbusreq0 & v845542;
assign v1216593 = locked_p & v1216592 | !locked_p & v845542;
assign v121627b = hmaster0_p & v1216227 | !hmaster0_p & v12160e2;
assign v1214d86 = hbusreq2_p & v1214d83 | !hbusreq2_p & v1214d85;
assign v1216719 = hmaster1_p & v1216718 | !hmaster1_p & v845542;
assign v134d3dd = hbusreq1_p & v134d27d | !hbusreq1_p & v134d3dc;
assign v12162b5 = hmaster1_p & v12162b4 | !hmaster1_p & v12161f4;
assign v10d40b1 = hmaster1_p & v10d40b0 | !hmaster1_p & v10d3fe9;
assign v1215338 = hmaster0_p & v12150aa | !hmaster0_p & v1215092;
assign f2f21d = hmaster2_p & v845542 | !hmaster2_p & !f2f21c;
assign v1405868 = stateG10_5_p & v1405867 | !stateG10_5_p & v1405865;
assign v1552f62 = hlock1 & v15533a1 | !hlock1 & v1552f61;
assign v16a1add = hgrant5_p & v845542 | !hgrant5_p & v16a1adc;
assign v138a304 = hbusreq5_p & v138a303 | !hbusreq5_p & v845542;
assign v1445ef5 = hgrant2_p & v1445ef3 | !hgrant2_p & v1445ef4;
assign v1284cd6 = hbusreq4_p & v1284cd5 | !hbusreq4_p & !v140589a;
assign v134cdc6 = hlock3 & v134d276 | !hlock3 & v134cdc5;
assign v16a1e56 = hbusreq5 & v16a1e4a | !hbusreq5 & v16a1e55;
assign v1445e06 = hlock0 & v1445e01 | !hlock0 & v1445e05;
assign v144616b = hmaster0_p & v1445fe3 | !hmaster0_p & v144608a;
assign v12153a6 = hbusreq4_p & v12153a5 | !hbusreq4_p & v1215364;
assign a653b4 = hgrant1_p & a653ae | !hgrant1_p & !a653a1;
assign v1216790 = hmaster0_p & v12165a9 | !hmaster0_p & v1216a91;
assign v144630c = hmaster2_p & v144639c | !hmaster2_p & v1446645;
assign d302f0 = hbusreq3_p & d302d3 | !hbusreq3_p & !d302ef;
assign v1553061 = hgrant2_p & v1553380 | !hgrant2_p & v1553060;
assign d2fc86 = hbusreq2_p & d2fc85 | !hbusreq2_p & v845542;
assign d80759 = stateG2_p & v845542 | !stateG2_p & d80757;
assign v1389392 = hgrant2_p & v845542 | !hgrant2_p & !v1389391;
assign f2f2a7 = hbusreq2_p & f2f2a3 | !hbusreq2_p & f2f2a6;
assign a662d0 = hgrant1_p & v845542 | !hgrant1_p & !a662cf;
assign v13893b5 = decide_p & v1389372 | !decide_p & v138a406;
assign v12160a0 = hbusreq5 & v121607d | !hbusreq5 & v121609f;
assign v1445da1 = hbusreq1 & v1445d9f | !hbusreq1 & v1445da0;
assign v16a1f9b = hmaster1_p & v845542 | !hmaster1_p & v16a1f96;
assign v1446714 = hmaster0_p & v144667f | !hmaster0_p & v1446440;
assign a6541f = hmaster2_p & a6588f | !hmaster2_p & a6587e;
assign v12afa0e = hgrant2_p & v12af73f | !hgrant2_p & v12afa0d;
assign v16a1392 = hbusreq2_p & v16a12c1 | !hbusreq2_p & v16a1391;
assign v1446265 = hbusreq5_p & v1446416 | !hbusreq5_p & v1446264;
assign v1445f63 = hmaster0_p & v14466af | !hmaster0_p & v14465b8;
assign v1445874 = hmaster2_p & v1445871 | !hmaster2_p & v1445872;
assign v1668d57 = hbusreq5_p & v1668d4e | !hbusreq5_p & !v1668d56;
assign f2e731 = hgrant5_p & v845542 | !hgrant5_p & !f2e730;
assign d30803 = hbusreq5_p & d30802 | !hbusreq5_p & !d30801;
assign v1214dd3 = hbusreq2 & v1214dd2 | !hbusreq2 & v845542;
assign v1445e54 = hmaster2_p & v144639c | !hmaster2_p & v1445def;
assign v15534fd = hlock0 & v15534fc | !hlock0 & v15534fb;
assign v12ad02d = hmaster0_p & v12ad029 | !hmaster0_p & !v12ad02c;
assign v1216313 = hbusreq2 & v1216308 | !hbusreq2 & v1216312;
assign a65688 = hmaster1_p & a65687 | !hmaster1_p & a658e5;
assign v12ad4da = hbusreq4_p & v12ad4d0 | !hbusreq4_p & v12ad4d4;
assign v14058ef = hmaster2_p & v14465b3 | !hmaster2_p & !v14058ee;
assign d8076f = hgrant5_p & v845542 | !hgrant5_p & d8076e;
assign v138a31b = hmaster0_p & v138a31a | !hmaster0_p & v845542;
assign v10d405e = hgrant4_p & v10d3fd5 | !hgrant4_p & v10d405d;
assign d300f7 = hbusreq1 & d2fe8a | !hbusreq1 & d2fe80;
assign v1515852 = hready_p & v1515850 | !hready_p & !v1515851;
assign d3022b = hbusreq5_p & d3022a | !hbusreq5_p & !d30229;
assign v1668d7d = hmaster2_p & v1668d72 | !hmaster2_p & v1668d7c;
assign v121505b = hgrant5_p & v1215471 | !hgrant5_p & v121505a;
assign v134d38d = hbusreq0 & v134d38c | !hbusreq0 & v134d38b;
assign v14458f5 = hbusreq4_p & v1446403 | !hbusreq4_p & v14458f4;
assign v1445505 = hlock0 & v1445504 | !hlock0 & v1445503;
assign v1445ecd = hmaster0_p & v14465b7 | !hmaster0_p & v1445ecc;
assign v144536a = hmaster0_p & v1445909 | !hmaster0_p & v1445a4f;
assign v1668c86 = hmaster2_p & a658ad | !hmaster2_p & !a658bd;
assign v1668d5c = hgrant5_p & v1668d43 | !hgrant5_p & v1668d5b;
assign v1405a8d = hmaster2_p & v845542 | !hmaster2_p & v1405a8c;
assign v1515651 = stateA1_p & a658a5 | !stateA1_p & !v110b6cc;
assign d2f9b6 = hlock4_p & v845542 | !hlock4_p & !d3094f;
assign d2fece = hbusreq4_p & d2fecd | !hbusreq4_p & v845542;
assign v12ae1fd = hgrant5_p & v845542 | !hgrant5_p & v12ae1fc;
assign v12162dc = hbusreq2_p & v12162d9 | !hbusreq2_p & v12162db;
assign d2fb1d = hgrant5_p & d3068e | !hgrant5_p & d2faee;
assign v1668c4e = hmaster2_p & v845542 | !hmaster2_p & v1668c4d;
assign d2fbf8 = hgrant5_p & d2fb53 | !hgrant5_p & d2fbf7;
assign v121614f = hlock0_p & v1216523 | !hlock0_p & v121614e;
assign v1446339 = hmaster2_p & v144663f | !hmaster2_p & v144668c;
assign v1445a31 = hlock0 & v1445a20 | !hlock0 & v1445a30;
assign v1445d9a = hlock1 & v1445d99 | !hlock1 & v1445d98;
assign v16695ad = hmaster1_p & v16695ac | !hmaster1_p & v845570;
assign v16a140a = hgrant2_p & v16a1d2c | !hgrant2_p & v16a1d8d;
assign a662bc = hready_p & a662bb | !hready_p & a662a4;
assign v1445e1b = hmaster0_p & v1445df8 | !hmaster0_p & v1445e00;
assign d30115 = hgrant5_p & d2fe8e | !hgrant5_p & d30114;
assign v14466e6 = hmaster1_p & v14463c9 | !hmaster1_p & v14463ef;
assign d30819 = hgrant5_p & d306d0 | !hgrant5_p & d307a1;
assign v1216171 = hgrant2_p & v12160ea | !hgrant2_p & v1216170;
assign d2fe85 = hbusreq1_p & d2fe80 | !hbusreq1_p & d2fe84;
assign f2ed9c = decide_p & f2f4bf | !decide_p & f2f23c;
assign v1214d20 = hgrant2_p & v1214ce7 | !hgrant2_p & v1214d1f;
assign v1515649 = stateG2_p & v88d3e4 | !stateG2_p & v845542;
assign v138a39b = hmaster1_p & v138a39a | !hmaster1_p & v138a341;
assign v15160fd = hbusreq4 & v15168ad | !hbusreq4 & v16693aa;
assign v1445ed0 = hbusreq2_p & v1445eac | !hbusreq2_p & v1445ecf;
assign d807b3 = decide_p & d80752 | !decide_p & d807b2;
assign a6588a = hmastlock_p & a65888 | !hmastlock_p & v845542;
assign v144588a = hmaster2_p & v14463b1 | !hmaster2_p & !v1445885;
assign v12166e3 = hmastlock_p & v12166e2 | !hmastlock_p & !v845542;
assign d2fc55 = hbusreq1_p & d2fbd4 | !hbusreq1_p & d2fc54;
assign v121658b = hbusreq5_p & v121658a | !hbusreq5_p & v845542;
assign v12150f5 = hlock2_p & v12150f4 | !hlock2_p & v12150f1;
assign v1214ef7 = hgrant5_p & v845542 | !hgrant5_p & v1216571;
assign a6563c = hmaster2_p & a6562e | !hmaster2_p & a6563b;
assign v1515c82 = hmaster0_p & v845542 | !hmaster0_p & v1515c81;
assign v12ad660 = hbusreq0 & v12ad5f7 | !hbusreq0 & !v12af73f;
assign v1445913 = hlock2 & v1445912 | !hlock2 & v144590c;
assign v1215051 = hmaster2_p & v845542 | !hmaster2_p & v1215050;
assign v1668d78 = hbusreq0_p & v1668d25 | !hbusreq0_p & !v1668d48;
assign v14458a6 = hlock0 & v14458a3 | !hlock0 & v14458a5;
assign v12ad67d = hbusreq4_p & a658ca | !hbusreq4_p & v12ad67c;
assign v1215da0 = hmaster1_p & v1215d81 | !hmaster1_p & !v1215d9b;
assign v134d3d3 = hbusreq2 & v134d3d1 | !hbusreq2 & v134d3d2;
assign d2f976 = hbusreq1_p & v84555a | !hbusreq1_p & d2f971;
assign d80773 = hgrant1_p & d80772 | !hgrant1_p & !v845542;
assign d3060c = hbusreq5_p & d3060b | !hbusreq5_p & v845542;
assign v1445eac = hgrant2_p & v1445e53 | !hgrant2_p & v1445eab;
assign v1214ff1 = hbusreq1_p & v1215bae | !hbusreq1_p & !v1214ff0;
assign v1216586 = hgrant0_p & v845570 | !hgrant0_p & !v845542;
assign v1389efd = hready_p & v1389e37 | !hready_p & v1389efc;
assign v134d4f7 = hbusreq0 & v134d4ef | !hbusreq0 & v134d4f6;
assign v1215780 = hmaster1_p & v121577f | !hmaster1_p & v1215770;
assign v1445df7 = hmaster2_p & v1445dec | !hmaster2_p & v1445df5;
assign v14454e8 = hmaster0_p & v144626d | !hmaster0_p & v144639c;
assign v14454fc = hmaster1_p & v14454fb | !hmaster1_p & v144627e;
assign v1215d76 = hgrant5_p & v12164df | !hgrant5_p & v12166df;
assign d80731 = stateA1_p & d80730 | !stateA1_p & !v936735;
assign v1668c57 = hgrant3_p & v1668c54 | !hgrant3_p & !v1668c56;
assign v16a12f9 = decide_p & v16a12f8 | !decide_p & v16a1db9;
assign v1445ea9 = hlock0 & v1445e96 | !hlock0 & v1445ea8;
assign v138932d = hbusreq3_p & v138916a | !hbusreq3_p & v138932c;
assign v12afe5f = hlock5_p & v12afe58 | !hlock5_p & v12afe5e;
assign v1668db8 = hbusreq5_p & v1668db6 | !hbusreq5_p & !v1668db7;
assign v134ce6a = hlock3 & v134d3b5 | !hlock3 & v134ce69;
assign v84557e = busreq_p & v845542 | !busreq_p & !v845542;
assign c50efc = decide_p & c50efb | !decide_p & v845550;
assign v121656a = hgrant0_p & v1216569 | !hgrant0_p & v845542;
assign v1214d45 = hbusreq0 & v1214d44 | !hbusreq0 & v845542;
assign v1405afa = hgrant2_p & v1405af5 | !hgrant2_p & v1405af9;
assign v12ad31f = hgrant5_p & d30690 | !hgrant5_p & v12ad31e;
assign f2f345 = hbusreq1 & v1668d27 | !hbusreq1 & v845542;
assign v1214ee7 = hbusreq5_p & v1214ee5 | !hbusreq5_p & v1214ee6;
assign v138a3bf = hbusreq5 & v138a3ae | !hbusreq5 & !v138a391;
assign v1445e8c = hbusreq4_p & v144639c | !hbusreq4_p & v144660d;
assign v12af7f5 = hbusreq1_p & v845542 | !hbusreq1_p & v12af7f4;
assign a65392 = hburst1 & v88d3e4 | !hburst1 & !v845542;
assign v16a129c = hbusreq2 & v16a1a95 | !hbusreq2 & v16a1a99;
assign d2fbb4 = hbusreq2_p & d2fbb3 | !hbusreq2_p & d2fbb2;
assign v16a205b = hmaster1_p & v9109e4 | !hmaster1_p & !v16a2672;
assign v1668dcd = hbusreq5_p & v1668dcb | !hbusreq5_p & !v1668dcc;
assign v1284ce6 = hmaster1_p & v1284ce5 | !hmaster1_p & !v1284cdf;
assign v1515ae8 = hmaster2_p & a6587e | !hmaster2_p & v1515ae7;
assign d30212 = hmaster2_p & d30210 | !hmaster2_p & d30211;
assign v10d4084 = hmaster0_p & v10d4064 | !hmaster0_p & v10d4083;
assign v1216701 = hgrant5_p & v845542 | !hgrant5_p & v1216700;
assign v1216255 = hmaster1_p & v121623c | !hmaster1_p & !v121624b;
assign v14058f8 = hbusreq5_p & v14058f0 | !hbusreq5_p & v14058f7;
assign v1552d47 = hbusreq0 & v1553392 | !hbusreq0 & v1553395;
assign v1446181 = hbusreq2 & v1446171 | !hbusreq2 & v1446180;
assign v134d537 = hlock3 & v134d534 | !hlock3 & v134d536;
assign f2f3e7 = hmaster1_p & f2f3e6 | !hmaster1_p & f2f39d;
assign d2fc03 = hlock0_p & v845542 | !hlock0_p & !v1668c1c;
assign v1284d50 = hmaster1_p & v1284d4f | !hmaster1_p & !v1284cdf;
assign f2f3cb = hgrant5_p & f2f2a8 | !hgrant5_p & !f2f38e;
assign f2ed9b = decide_p & f2ed9a | !decide_p & f2f23c;
assign v1214cd1 = hbusreq0 & v1214cd0 | !hbusreq0 & v845542;
assign v144644e = hmaster1_p & v1446405 | !hmaster1_p & v144644d;
assign v14457e2 = hmaster0_p & v14457d7 | !hmaster0_p & v1445ec3;
assign v144669a = hlock1 & v14465f2 | !hlock1 & v1446699;
assign v1214d04 = hmaster0_p & v1214cfd | !hmaster0_p & v1214d03;
assign v1445883 = hlock1 & v1445882 | !hlock1 & v144586d;
assign v138a310 = hmaster0_p & v138a30e | !hmaster0_p & v138a30f;
assign v1445ebe = hbusreq2_p & v1445eac | !hbusreq2_p & v1445ebd;
assign v1215034 = hbusreq1_p & v1215461 | !hbusreq1_p & !v1215033;
assign a65862 = locked_p & v845542 | !locked_p & !a65861;
assign v1215b85 = hlock4_p & v1216145 | !hlock4_p & v121614f;
assign v134d51b = hmaster1_p & v134d51a | !hmaster1_p & v845542;
assign a65890 = hmaster2_p & a6587e | !hmaster2_p & a6588f;
assign f2f238 = hmaster0_p & f2f237 | !hmaster0_p & f2f22c;
assign v1216564 = hbusreq5_p & v1216563 | !hbusreq5_p & v845542;
assign v1214d68 = hmaster1_p & v1214d67 | !hmaster1_p & v1214d5f;
assign d3013b = hgrant5_p & d3013a | !hgrant5_p & !d300e0;
assign v1215c50 = hbusreq2_p & v1215c4e | !hbusreq2_p & v1215c4f;
assign v144621d = hmaster0_p & v144639c | !hmaster0_p & v144621c;
assign v1668e10 = jx1_p & v1668c59 | !jx1_p & v1668e0f;
assign v15167c0 = hmaster0_p & v845542 | !hmaster0_p & v15167bf;
assign v1284d54 = hgrant2_p & v1284d43 | !hgrant2_p & v1284d53;
assign d2f99e = hmaster2_p & d3068e | !hmaster2_p & d2f99d;
assign d30794 = hlock1_p & v845542 | !hlock1_p & d30649;
assign v1446443 = hbusreq2_p & v1446437 | !hbusreq2_p & v1446442;
assign v143fd79 = hgrant1_p & v845542 | !hgrant1_p & v143fd78;
assign v16a1a7c = hbusreq0 & v16a1a7b | !hbusreq0 & v16a194e;
assign v12ad1fc = hbusreq2_p & v12ad0bc | !hbusreq2_p & v12af9b5;
assign v144577f = hmaster1_p & v144577e | !hmaster1_p & v1445e07;
assign v138a006 = hmaster0_p & v138a002 | !hmaster0_p & v1389de1;
assign v121607a = hlock2_p & v1216077 | !hlock2_p & v1216079;
assign v144543a = hlock5 & v144541f | !hlock5 & v1445439;
assign v144673b = hmaster0_p & v144643e | !hmaster0_p & v1446638;
assign v12160e7 = hready_p & v1216046 | !hready_p & v12160e6;
assign v1284c94 = hmaster1_p & v1284c93 | !hmaster1_p & v140584d;
assign f2f299 = hbusreq1 & a65862 | !hbusreq1 & v845542;
assign d2fbaa = hmaster1_p & d2fb93 | !hmaster1_p & d2fb9d;
assign v1215c01 = hmaster2_p & v1215bf6 | !hmaster2_p & v1216538;
assign v14457ef = hmaster0_p & v1445eb8 | !hmaster0_p & v14465b7;
assign v1445a62 = hmaster1_p & v14459a2 | !hmaster1_p & v1445a61;
assign v12afda4 = hmaster2_p & v845542 | !hmaster2_p & !v12afda3;
assign v11e5964 = hgrant4_p & v11e593a | !hgrant4_p & !v845542;
assign v134d44d = hbusreq0 & v134d44c | !hbusreq0 & v134d379;
assign v144546f = hbusreq2_p & v1446272 | !hbusreq2_p & v1445bba;
assign v10d4298 = hgrant1_p & v10d3fe0 | !hgrant1_p & v10d4293;
assign v1445435 = hgrant2_p & v1445411 | !hgrant2_p & v1445434;
assign v134d45a = hlock5 & v134d3b5 | !hlock5 & v134d449;
assign v134d3c0 = hbusreq4_p & v134d1e8 | !hbusreq4_p & v134d3bf;
assign a6540d = hmaster0_p & v845558 | !hmaster0_p & a6540c;
assign d302e2 = hlock5_p & d302e1 | !hlock5_p & d30663;
assign v1445b71 = hlock2 & v144632f | !hlock2 & v1445b70;
assign v16a1a82 = hbusreq2 & v16a1a7f | !hbusreq2 & !v16a1a81;
assign v12afe4e = hgrant4_p & v845542 | !hgrant4_p & !v12afe4d;
assign v1553443 = hbusreq2_p & v155323a | !hbusreq2_p & v1553442;
assign v144608d = hbusreq1_p & v144665a | !hbusreq1_p & v14465d7;
assign v144626d = hlock0 & v144626c | !hlock0 & v1446445;
assign v15156cb = hlock2_p & v15156be | !hlock2_p & !v15156ca;
assign d30650 = hbusreq1_p & d3064f | !hbusreq1_p & !v845542;
assign v1668d65 = hbusreq1_p & v1668d62 | !hbusreq1_p & v1668d64;
assign v12ad614 = hgrant5_p & v845542 | !hgrant5_p & !v12ad5dc;
assign v1214f0f = hmaster0_p & v1214f0d | !hmaster0_p & v1214f0e;
assign f2f378 = hbusreq0 & f2f36f | !hbusreq0 & f2f377;
assign d2f9ca = hbusreq5_p & d2f9c9 | !hbusreq5_p & d2f98e;
assign v155308c = hmaster0_p & v845542 | !hmaster0_p & v155308b;
assign v14459cd = hbusreq1 & v14459c9 | !hbusreq1 & v14459cc;
assign v1515ae1 = hlock2_p & v1515ae0 | !hlock2_p & !v845542;
assign v1668c5f = hmaster2_p & a658ad | !hmaster2_p & !v84556a;
assign v144616d = hmaster0_p & v1446081 | !hmaster0_p & v1446092;
assign v1515810 = hbusreq2_p & v151580f | !hbusreq2_p & v845542;
assign v14460e6 = decide_p & v14460e5 | !decide_p & v144639b;
assign bf1f56 = decide_p & v84556a | !decide_p & bf1f55;
assign v15157f1 = hbusreq0 & v15157eb | !hbusreq0 & v15157f0;
assign v134d3c8 = hbusreq2_p & v134d267 | !hbusreq2_p & v134d3c4;
assign v155341e = hgrant2_p & v1553380 | !hgrant2_p & v155341d;
assign v16a1422 = hbusreq2 & v16a1421 | !hbusreq2 & !v16a205c;
assign v1446718 = hmaster1_p & v1446717 | !hmaster1_p & v1446436;
assign v1445eb4 = hmaster2_p & v144639c | !hmaster2_p & v1445e74;
assign f2f4b1 = hbusreq1 & a66275 | !hbusreq1 & !f2f4b0;
assign v1215711 = hgrant0_p & v121570f | !hgrant0_p & !v1215710;
assign v1284cd0 = hgrant5_p & v140589f | !hgrant5_p & v1284cce;
assign d2fbe8 = hbusreq1_p & d2fbe7 | !hbusreq1_p & v84554a;
assign v1446081 = hlock0 & v1446080 | !hlock0 & v144607d;
assign v1215d9c = hmaster1_p & v1215d6e | !hmaster1_p & !v1215d9b;
assign v1446672 = hmaster1_p & v1446671 | !hmaster1_p & v144644d;
assign v1215d2b = hmaster0_p & v1215d2a | !hmaster0_p & v1216a99;
assign v10d3fd9 = locked_p & v10d3fd7 | !locked_p & v10d3fd8;
assign v1214ed6 = hbusreq5_p & v1214ed4 | !hbusreq5_p & v1214ed5;
assign v12164d8 = hmaster0_p & v12164d5 | !hmaster0_p & v12164d7;
assign v1214ddc = hbusreq2 & v1216a81 | !hbusreq2 & v845542;
assign f2f2de = hmaster0_p & f2f2cc | !hmaster0_p & f2f2dd;
assign d301c0 = hmaster2_p & d306da | !hmaster2_p & d306df;
assign v1668cd2 = hmaster2_p & v1668cd0 | !hmaster2_p & v1668cd1;
assign v1214d37 = hmaster1_p & v845547 | !hmaster1_p & v121536b;
assign a6535b = hmaster0_p & a65852 | !hmaster0_p & a6585e;
assign v16a2060 = hmaster1_p & v9337f3 | !hmaster1_p & v16a1f96;
assign d8077e = hgrant0_p & d8077d | !hgrant0_p & !v845542;
assign d80748 = hmaster2_p & d8073a | !hmaster2_p & !v845542;
assign v134ce57 = hgrant2_p & v134ce56 | !hgrant2_p & v134ce47;
assign a662c3 = hmaster1_p & v845542 | !hmaster1_p & a662c2;
assign v12ad664 = hbusreq5_p & v845542 | !hbusreq5_p & v12ad663;
assign v121639f = hmaster0_p & v845542 | !hmaster0_p & v121639e;
assign v16a139f = jx2_p & v16a1a91 | !jx2_p & v16a139e;
assign v1668cdf = hbusreq1_p & v1668cde | !hbusreq1_p & !v845542;
assign d2fb58 = hlock0_p & v845542 | !hlock0_p & !d305de;
assign d30772 = hmaster1_p & d3072e | !hmaster1_p & d30754;
assign v1389fcd = decide_p & v1389fcc | !decide_p & v845542;
assign d30279 = hbusreq5_p & d30278 | !hbusreq5_p & !d30277;
assign v1668dc7 = hgrant5_p & v1668dc2 | !hgrant5_p & v1668d5b;
assign v12160a7 = hmaster1_p & v12160a6 | !hmaster1_p & v121605d;
assign v14464a7 = hmaster0_p & v845542 | !hmaster0_p & v14464a6;
assign v1445a2e = hmaster2_p & v1445a2d | !hmaster2_p & v144660f;
assign v1214dba = hbusreq2_p & v1214db7 | !hbusreq2_p & v1214db9;
assign d30640 = hready_p & d305e7 | !hready_p & d3063f;
assign v134d370 = hbusreq4 & v134d36e | !hbusreq4 & v134d36f;
assign v1214f1b = hbusreq5 & v1214eff | !hbusreq5 & v1214f1a;
assign f2e4e9 = hready_p & v845542 | !hready_p & f2e4e8;
assign v1668de5 = hbusreq2 & v1668de1 | !hbusreq2 & v1668de4;
assign v1515831 = hready_p & v1515818 | !hready_p & v1515830;
assign v12acfe4 = hmaster1_p & v12acfc9 | !hmaster1_p & v12ad54f;
assign v1215b9c = hbusreq1_p & v1215b99 | !hbusreq1_p & v121611f;
assign v1553431 = hlock2 & v155321a | !hlock2 & v1553430;
assign v1445834 = hbusreq2_p & v1445830 | !hbusreq2_p & v1445833;
assign v1668c8f = hbusreq2 & v1668c83 | !hbusreq2 & v1668c8e;
assign v134d4d5 = hbusreq0_p & v134d1dd | !hbusreq0_p & v134d4ca;
assign v10d40bc = hlock0_p & v10d3fd4 | !hlock0_p & v10d40bb;
assign v138a45a = hmaster1_p & v138a459 | !hmaster1_p & v138a341;
assign v155309e = hlock2 & v155309b | !hlock2 & v155309d;
assign v12af590 = hgrant5_p & v845542 | !hgrant5_p & v12af58f;
assign v1216190 = hgrant5_p & v121618f | !hgrant5_p & v1216118;
assign v155339f = hgrant1_p & v845542 | !hgrant1_p & v155339e;
assign v1215734 = hlock4_p & v1216136 | !hlock4_p & !v845542;
assign v14058d2 = hlock0_p & v140583f | !hlock0_p & v14058d1;
assign v12167ab = hbusreq5 & v12167aa | !hbusreq5 & v845542;
assign v1446212 = stateG10_5_p & v1446211 | !stateG10_5_p & !v144639c;
assign v1445a85 = hmaster1_p & v1445a39 | !hmaster1_p & v144591b;
assign v1553512 = hlock3 & v155321a | !hlock3 & v1553511;
assign v1445bc5 = hgrant2_p & v1446461 | !hgrant2_p & v1445bc4;
assign v1215767 = hlock4_p & v1215765 | !hlock4_p & v1215766;
assign v144552c = hgrant2_p & v14454e9 | !hgrant2_p & v144552b;
assign v14058f4 = hgrant1_p & v14058f1 | !hgrant1_p & v14058f3;
assign v144536f = hlock2 & v1445369 | !hlock2 & v144536e;
assign v10d4045 = hbusreq4_p & v10d3fe7 | !hbusreq4_p & !v10d3ff9;
assign v1668d48 = hbusreq4 & a65861 | !hbusreq4 & v845542;
assign f2f221 = hbusreq5_p & f2f21d | !hbusreq5_p & f2f220;
assign v12ad031 = hgrant2_p & v12ad5f5 | !hgrant2_p & v12ad022;
assign v1284d12 = hgrant5_p & v1284d0f | !hgrant5_p & v1284d11;
assign v121654e = hbusreq5_p & v121654d | !hbusreq5_p & v845542;
assign v1216094 = hmaster2_p & v121602d | !hmaster2_p & v845542;
assign d3015a = hmaster0_p & d30137 | !hmaster0_p & d30159;
assign v121678b = hbusreq2 & v12164e7 | !hbusreq2 & v121671a;
assign v1515629 = hmaster0_p & v1515628 | !hmaster0_p & v1668da6;
assign v12150c0 = decide_p & v12150ba | !decide_p & !v12150bf;
assign v1445ec2 = hbusreq0 & v1445ec1 | !hbusreq0 & v1445eae;
assign v1215fb7 = hmaster1_p & v1215fb6 | !hmaster1_p & v12164e1;
assign v15157c0 = hgrant4_p & a662a9 | !hgrant4_p & v15157bf;
assign v1214eb7 = hlock2_p & v1214eb6 | !hlock2_p & !v12163ab;
assign v144665f = hmaster2_p & v14465b0 | !hmaster2_p & v144665b;
assign v12ad327 = hbusreq5_p & v12ae1fd | !hbusreq5_p & v12ad326;
assign f2e27a = decide_p & f2e279 | !decide_p & v845542;
assign v1215737 = hlock0_p & v121611e | !hlock0_p & v121611f;
assign v1445501 = hbusreq2 & v14454f3 | !hbusreq2 & v1445500;
assign v134ce8f = hlock0 & v134ce8e | !hlock0 & v134ce8d;
assign v1389d72 = hlock5_p & v1389d71 | !hlock5_p & v845542;
assign f2e4c8 = hgrant3_p & f2e27b | !hgrant3_p & f2e4c7;
assign v15167ee = hbusreq2 & v15167eb | !hbusreq2 & v15167ed;
assign v1446477 = hmaster2_p & v1446476 | !hmaster2_p & v845542;
assign a65628 = hbusreq1_p & a65380 | !hbusreq1_p & a65627;
assign v1668c33 = hlock3_p & v1668c32 | !hlock3_p & v845542;
assign v845586 = stateG3_1_p & v845542 | !stateG3_1_p & !v845542;
assign v14453c1 = hbusreq3 & v14453bf | !hbusreq3 & v14453c0;
assign d300c3 = hgrant4_p & v845542 | !hgrant4_p & d300c2;
assign d2fc34 = hbusreq0 & d2fb74 | !hbusreq0 & d2fc33;
assign v14461be = hgrant2_p & v14461bd | !hgrant2_p & v14461b9;
assign v134d519 = hlock0 & v134d518 | !hlock0 & v134d516;
assign v12ad4e3 = hbusreq2_p & v12ad4de | !hbusreq2_p & v12ad4e2;
assign v12150de = hmaster2_p & v12153ce | !hmaster2_p & v12150c4;
assign v12aeb83 = hlock3_p & v12aeb40 | !hlock3_p & v12aeb82;
assign v155305d = hgrant5_p & v845542 | !hgrant5_p & v155305c;
assign v1445ddd = hlock3 & v1445dc6 | !hlock3 & v1445ddc;
assign v1216528 = hready & v1216527 | !hready & v845542;
assign v12ad561 = hbusreq2 & v12ad55b | !hbusreq2 & v12ad560;
assign v14461c1 = hbusreq2 & v14461bc | !hbusreq2 & v14461c0;
assign v14453e6 = hlock2 & v14453e4 | !hlock2 & v14453e5;
assign v1445b16 = hmaster1_p & v1445af5 | !hmaster1_p & v144591b;
assign v1668c5a = hbusreq3 & v845570 | !hbusreq3 & v845542;
assign v138944d = hbusreq5_p & v138944c | !hbusreq5_p & v845542;
assign v12160da = hbusreq5_p & f2f2ad | !hbusreq5_p & v12160d9;
assign v1215bb8 = hbusreq2 & v12163ad | !hbusreq2 & v1215bb7;
assign v138a3dd = hlock5_p & v138a3dc | !hlock5_p & !v15157cc;
assign v845559 = hbusreq4 & v845542 | !hbusreq4 & !v845542;
assign v1389e2a = hmaster2_p & v15168f8 | !hmaster2_p & v845542;
assign v1445acf = hmaster1_p & v1445ab0 | !hmaster1_p & v14458c1;
assign v16a1e8e = hbusreq1_p & v16a206e | !hbusreq1_p & v16a1e8d;
assign v1668c69 = hburst1 & a66272 | !hburst1 & v1668c68;
assign v134d1f2 = hbusreq1_p & v134d1f1 | !hbusreq1_p & v845542;
assign a656ad = hmaster1_p & a658f1 | !hmaster1_p & !a65916;
assign v1446096 = hbusreq2_p & v1446075 | !hbusreq2_p & v1446095;
assign v1215772 = hgrant2_p & v121570b | !hgrant2_p & v1215771;
assign v1389391 = hmaster1_p & v1389389 | !hmaster1_p & !v1389390;
assign v16a1aee = hbusreq2 & v16a1aeb | !hbusreq2 & !v16a1aed;
assign v1445409 = hgrant2_p & v1446461 | !hgrant2_p & v1445408;
assign v1215741 = hgrant5_p & v1215740 | !hgrant5_p & v121573e;
assign f2f281 = hbusreq1_p & v845570 | !hbusreq1_p & !v845542;
assign v1553428 = hbusreq0_p & v1553140 | !hbusreq0_p & v845542;
assign d2fc5c = hgrant4_p & d2fbea | !hgrant4_p & d2fc5b;
assign v144628e = hbusreq0 & v144628d | !hbusreq0 & v1446265;
assign v134d1fe = hbusreq5_p & v134d1fa | !hbusreq5_p & v134d1fd;
assign v12ad8e4 = hbusreq1_p & v12adf5d | !hbusreq1_p & v12ad8e3;
assign v16a13d7 = hbusreq3 & v16a13d1 | !hbusreq3 & v16a13d6;
assign d30657 = hbusreq5_p & d30653 | !hbusreq5_p & d30656;
assign d30912 = hmaster2_p & d305ea | !hmaster2_p & d30911;
assign f2f37d = hbusreq1_p & f2f37c | !hbusreq1_p & v845542;
assign v1214e71 = hlock5_p & v1214e70 | !hlock5_p & v1214df5;
assign v1214e5a = hmaster0_p & v1214e59 | !hmaster0_p & v12162e8;
assign v1446395 = stateG3_2_p & v845542 | !stateG3_2_p & !v1446394;
assign v1405ae2 = hmaster2_p & v1405a87 | !hmaster2_p & v1405adc;
assign v1214d7d = hgrant2_p & v1214c82 | !hgrant2_p & v1214d78;
assign d30880 = hmaster1_p & d3087f | !hmaster1_p & !d30706;
assign v10d409f = hmaster0_p & v10d407f | !hmaster0_p & v10d3fdc;
assign v121606f = hbusreq2_p & v121606e | !hbusreq2_p & v121606d;
assign v12af9c3 = hbusreq5_p & v12afe47 | !hbusreq5_p & v12af9c2;
assign v1214c06 = hmaster1_p & v1214c05 | !hmaster1_p & v12153a9;
assign d3063d = hbusreq5 & d3063c | !hbusreq5 & d30631;
assign v8dfa41 = hburst0_p & v845542 | !hburst0_p & v87abb5;
assign v14459fe = hgrant5_p & v14459a4 | !hgrant5_p & v14459fd;
assign v1446298 = hbusreq2_p & v1446291 | !hbusreq2_p & v1446294;
assign v144660c = hlock0_p & v14463b1 | !hlock0_p & v14463ba;
assign v1445f05 = hgrant5_p & v1445f04 | !hgrant5_p & v1445eeb;
assign a65449 = hgrant2_p & a653f4 | !hgrant2_p & a65446;
assign v16a1a7b = hbusreq5_p & v16a1943 | !hbusreq5_p & v16a1a7a;
assign v1445ad0 = hmaster1_p & v14458a6 | !hmaster1_p & v14458c1;
assign v16695a7 = hready_p & v845542 | !hready_p & v16695a6;
assign v12acfcd = hbusreq2_p & v12acfca | !hbusreq2_p & v12acfcc;
assign v1215020 = hgrant2_p & v121501b | !hgrant2_p & v121501f;
assign v1515768 = hbusreq1 & v1515614 | !hbusreq1 & v845570;
assign v121579c = hgrant5_p & v845542 | !hgrant5_p & v1215760;
assign v16695a2 = hbusreq3 & v166959f | !hbusreq3 & v16695a1;
assign v1214dcd = hmaster0_p & v1216a62 | !hmaster0_p & v1214dcc;
assign v121626a = decide_p & v12160cf | !decide_p & v1216269;
assign v15156f8 = hbusreq2_p & v15156f7 | !hbusreq2_p & v845542;
assign v134cec2 = hready_p & v134d1e2 | !hready_p & v134cec1;
assign v16a266f = hmaster2_p & v845559 | !hmaster2_p & v845542;
assign v14460f7 = hmaster0_p & v1445fa9 | !hmaster0_p & v1445fa2;
assign v1445de8 = hmaster0_p & v1445de6 | !hmaster0_p & v1445de7;
assign v1216a77 = hready & v1216a66 | !hready & v1216a76;
assign v16a16a6 = hbusreq5_p & v16a209a | !hbusreq5_p & v16a16a5;
assign f2f435 = hgrant1_p & f2f281 | !hgrant1_p & !f2f38c;
assign d2fcea = hmaster1_p & d2fce9 | !hmaster1_p & !d2fcb5;
assign v1445b7b = hmaster1_p & v14465b7 | !hmaster1_p & v1445b7a;
assign v1445fc8 = hlock5 & v1445fb6 | !hlock5 & v1445fc7;
assign v14457b4 = hlock2 & v1445786 | !hlock2 & v14457b2;
assign v138a47e = hmaster1_p & v138a47d | !hmaster1_p & v138a43e;
assign v11e594e = hgrant5_p & v11e5949 | !hgrant5_p & !v11e594d;
assign v1214dd9 = hbusreq2_p & v1214dd8 | !hbusreq2_p & v845542;
assign f2f2e9 = hmaster0_p & f2f2cc | !hmaster0_p & f2f2e8;
assign v1445844 = hgrant2_p & v144581d | !hgrant2_p & v1445843;
assign v16a2243 = hmaster2_p & v845547 | !hmaster2_p & v845542;
assign v16a1cbf = hbusreq2 & v16a1cbc | !hbusreq2 & v16a1cbe;
assign v12af9c1 = hgrant1_p & d30690 | !hgrant1_p & v12af9c0;
assign v1446163 = hmaster0_p & v1446081 | !hmaster0_p & v144603f;
assign d2fe92 = hlock4_p & d306f3 | !hlock4_p & d305de;
assign f2e4e2 = hbusreq3_p & f2e4d6 | !hbusreq3_p & f2e4e1;
assign v10d4094 = hmaster1_p & v10d4093 | !hmaster1_p & v10d407c;
assign d302ea = hmaster1_p & d306bc | !hmaster1_p & d302e9;
assign v1445afb = hmaster1_p & v1445afa | !hmaster1_p & v14458fd;
assign d2fd3d = hbusreq2_p & v845542 | !hbusreq2_p & d302da;
assign v1515838 = hgrant5_p & v1515832 | !hgrant5_p & v1515837;
assign v1216139 = hgrant4_p & v1216137 | !hgrant4_p & v1216138;
assign v14457b3 = hlock2 & v14457b0 | !hlock2 & v14457b2;
assign v1446348 = hgrant2_p & v1446334 | !hgrant2_p & v1446347;
assign v151577f = hgrant4_p & v151576f | !hgrant4_p & v151577e;
assign v1405915 = hmaster2_p & v1405914 | !hmaster2_p & v14463b1;
assign v1215ba4 = hmaster0_p & v1215b98 | !hmaster0_p & v1215ba3;
assign v1216108 = hbusreq1 & v1216107 | !hbusreq1 & v845542;
assign v1445de1 = hbusreq5 & v1445ddf | !hbusreq5 & v1445de0;
assign v15532cc = hmaster1_p & v1553224 | !hmaster1_p & v15532cb;
assign v1445e2d = hbusreq2_p & v1445e29 | !hbusreq2_p & v1445e2c;
assign d3066a = hlock5_p & v845542 | !hlock5_p & d30669;
assign v1216141 = hlock1_p & v121613a | !hlock1_p & v1216140;
assign v1445dd7 = hbusreq2_p & v1445dd2 | !hbusreq2_p & v1445dd3;
assign v1216286 = hmaster1_p & v1216285 | !hmaster1_p & v121616f;
assign v12afe55 = hgrant4_p & v845542 | !hgrant4_p & !v12afe54;
assign v16a1a76 = hgrant4_p & v845559 | !hgrant4_p & v16a1a75;
assign v1216a86 = hburst0_p & v118e18f | !hburst0_p & v1216a85;
assign v12adf5d = hbusreq4_p & v12afda1 | !hbusreq4_p & v12afda3;
assign v1552f71 = hmaster1_p & v1552f70 | !hmaster1_p & v845542;
assign v1215040 = hgrant5_p & v121503d | !hgrant5_p & !v121503f;
assign v144618e = hmaster1_p & v144618d | !hmaster1_p & v1445fde;
assign v1668cf0 = hmaster2_p & a658ad | !hmaster2_p & !v1668cc4;
assign d8074c = hbusreq2_p & d8074b | !hbusreq2_p & d8074a;
assign v16a138d = hbusreq2 & v16a138c | !hbusreq2 & v16a129f;
assign v121600c = hmaster0_p & v1215ffc | !hmaster0_p & v121600b;
assign v1214fc5 = hmaster0_p & v1214fb6 | !hmaster0_p & v1214fc4;
assign d3087a = hbusreq5 & d30873 | !hbusreq5 & d30879;
assign v1446069 = hbusreq1_p & v1446068 | !hbusreq1_p & v144660e;
assign v16a1ac6 = hbusreq2_p & v16a267a | !hbusreq2_p & v16a1ac5;
assign v138a0c6 = jx2_p & v138a093 | !jx2_p & v138a092;
assign v12af1bc = hbusreq1_p & v12af3a7 | !hbusreq1_p & !v12af988;
assign v1284d29 = hready_p & v1284d06 | !hready_p & !v1284d28;
assign v1216546 = hgrant1_p & v1216545 | !hgrant1_p & v845542;
assign a6562c = hgrant4_p & a662a9 | !hgrant4_p & !a65384;
assign v1445482 = hlock2 & v144546f | !hlock2 & v1445481;
assign v1668cc9 = hbusreq5_p & v1668cc7 | !hbusreq5_p & !v1668cc8;
assign d30642 = hmaster1_p & d30641 | !hmaster1_p & d305db;
assign d307d7 = hgrant4_p & d307d3 | !hgrant4_p & d307d6;
assign v1552fcf = hlock3 & v155321a | !hlock3 & v1552fce;
assign v1445860 = hbusreq2_p & v1445854 | !hbusreq2_p & v144585c;
assign v16a1e0a = hmaster1_p & v16a1d78 | !hmaster1_p & v16a209c;
assign v12ad66c = hmaster1_p & v12ad66b | !hmaster1_p & !v12ad525;
assign v1445b2b = hbusreq5 & v1445b29 | !hbusreq5 & v1445b2a;
assign a64708 = decide_p & a646da | !decide_p & a662a2;
assign v16a1956 = hmaster2_p & v16a206f | !hmaster2_p & v16a1955;
assign v1445a77 = stateG10_5_p & v14459dc | !stateG10_5_p & v1445a76;
assign v14457f1 = hgrant2_p & v14457ee | !hgrant2_p & v14457f0;
assign v845574 = hgrant1_p & v845542 | !hgrant1_p & !v845542;
assign v1405add = hmaster2_p & v845542 | !hmaster2_p & !v1405adc;
assign v10d3fe5 = hbusreq4_p & v10d3fdb | !hbusreq4_p & v10d3fe0;
assign v12161a6 = hmaster0_p & v845542 | !hmaster0_p & v121602e;
assign v14458db = hlock0_p & v14458d9 | !hlock0_p & v14458da;
assign v14466f0 = hmaster0_p & v144663a | !hmaster0_p & v1446404;
assign f2f45e = decide_p & f2f413 | !decide_p & f2f23c;
assign v144546c = hmaster0_p & v144546b | !hmaster0_p & v1446404;
assign v121532e = hbusreq2 & v1215327 | !hbusreq2 & v121532d;
assign d2fefc = hbusreq2_p & d2fefb | !hbusreq2_p & d2fefa;
assign v1445fff = hbusreq2_p & v1445ffd | !hbusreq2_p & v1445ffe;
assign f2f339 = hmaster1_p & f2f2ef | !hmaster1_p & !f2f330;
assign v1445454 = hbusreq2_p & v1445453 | !hbusreq2_p & v1445bb3;
assign v144615b = hbusreq3 & v1446151 | !hbusreq3 & v144615a;
assign v14465f3 = hlock1 & v14465f2 | !hlock1 & v14465f0;
assign v16a169c = hgrant5_p & v845542 | !hgrant5_p & v16a1e98;
assign v1284d1c = hgrant1_p & v1446429 | !hgrant1_p & v1284d1b;
assign v15534dd = hgrant2_p & v1553380 | !hgrant2_p & v15534dc;
assign v1445770 = hlock3 & v1445f40 | !hlock3 & v144576e;
assign v1445994 = hready & v1445993 | !hready & v144639c;
assign d308df = hburst1 & d3073c | !hburst1 & v845542;
assign v1553393 = hgrant1_p & v1553217 | !hgrant1_p & v845542;
assign v1445ee3 = hbusreq2_p & v1445eac | !hbusreq2_p & v1445ee2;
assign v138a3a6 = hmaster0_p & v138a34f | !hmaster0_p & v138a34b;
assign d30294 = hmaster1_p & d30273 | !hmaster1_p & !d30293;
assign v1446009 = hbusreq5 & v1446007 | !hbusreq5 & v1446008;
assign d2faf5 = hbusreq1_p & d300c3 | !hbusreq1_p & d2fae0;
assign a656b6 = hready_p & a65682 | !hready_p & a656b4;
assign v16a1cc1 = hgrant2_p & v16a2062 | !hgrant2_p & v16a1cc0;
assign v12150cd = hlock4_p & v12150cc | !hlock4_p & !v12153e7;
assign v10d4023 = hgrant4_p & v10d4020 | !hgrant4_p & v10d4022;
assign v134d524 = hbusreq2_p & v134d520 | !hbusreq2_p & v134d523;
assign d308c6 = hbusreq0 & d308c3 | !hbusreq0 & d308c5;
assign v16a1be8 = hmaster0_p & v16a1be4 | !hmaster0_p & v16a1be7;
assign v1445a91 = hlock2 & v1445a69 | !hlock2 & v1445a90;
assign v1446442 = hmaster1_p & v1446441 | !hmaster1_p & v1446436;
assign a66273 = stateA1_p & a66272 | !stateA1_p & !v156645f;
assign f2f45b = hbusreq2 & f2f457 | !hbusreq2 & f2f45a;
assign v16a2666 = stateG2_p & v845542 | !stateG2_p & !v893df7;
assign a65472 = hlock0_p & a65469 | !hlock0_p & a658de;
assign d306c6 = hgrant3_p & d306a2 | !hgrant3_p & d306c5;
assign v1445e36 = decide_p & v1445de1 | !decide_p & v1445e35;
assign d308a7 = hbusreq1_p & d307eb | !hbusreq1_p & d306a5;
assign v14454eb = hgrant5_p & v144643a | !hgrant5_p & v14454ea;
assign v121617c = hbusreq5_p & v121617a | !hbusreq5_p & !v121617b;
assign d308c3 = hbusreq5_p & d30829 | !hbusreq5_p & d308c2;
assign v138a444 = hmaster0_p & v138a443 | !hmaster0_p & v84555c;
assign v1445856 = hgrant2_p & v1445831 | !hgrant2_p & v1445855;
assign v1668c34 = decide_p & v1668c33 | !decide_p & !v845542;
assign v144627d = hlock0 & v144627c | !hlock0 & v1446433;
assign v16a143a = hgrant5_p & v845542 | !hgrant5_p & v16a1439;
assign v1215bd8 = decide_p & v1215bd5 | !decide_p & v1215bd7;
assign v1668c49 = hbusreq1_p & a66275 | !hbusreq1_p & v84556a;
assign a65aea = hbusreq1_p & a66298 | !hbusreq1_p & a662aa;
assign v1284d22 = hmaster2_p & v1284d0c | !hmaster2_p & !v14465d8;
assign v1214bf8 = hbusreq5 & v1214bc9 | !hbusreq5 & v1214bf7;
assign v12acd05 = jx2_p & v12ad27c | !jx2_p & v12ae83c;
assign v12adf61 = hbusreq4_p & v12adf60 | !hbusreq4_p & !v84554a;
assign f2f2ef = hmaster0_p & f2f2e3 | !hmaster0_p & f2f2dd;
assign v1389dfa = hmaster1_p & v1389de1 | !hmaster1_p & v1389df9;
assign v12afe64 = hbusreq5_p & v12afe5f | !hbusreq5_p & v12afe63;
assign v1445a48 = hlock1 & v144660b | !hlock1 & v14459b1;
assign v134ce70 = hready_p & v134d34f | !hready_p & v134ce6f;
assign d30683 = hgrant3_p & d30640 | !hgrant3_p & d30682;
assign v10d3ff6 = hbusreq5_p & v10d3ff4 | !hbusreq5_p & !v10d3ff5;
assign v134d3d8 = hready_p & v134d3be | !hready_p & v134d3d7;
assign v12af3a6 = hbusreq1 & v12afda6 | !hbusreq1 & !v84554a;
assign v1445f26 = decide_p & v1445f25 | !decide_p & v144639b;
assign d301d0 = hbusreq1_p & d301cf | !hbusreq1_p & !d301ce;
assign v134d4d8 = hgrant4_p & v845542 | !hgrant4_p & v134d4d7;
assign a65b3a = decide_p & a65b29 | !decide_p & a662a2;
assign v1445a94 = hbusreq3 & v1445a92 | !hbusreq3 & v1445a93;
assign v16a1386 = hmaster0_p & v16a1383 | !hmaster0_p & v16a1a97;
assign v1405906 = hmaster0_p & v14058b4 | !hmaster0_p & v1405856;
assign v16a1bb6 = hburst0 & v16a1bb4 | !hburst0 & v16a1bb5;
assign v15532be = hgrant2_p & v845542 | !hgrant2_p & v1553239;
assign v1446128 = hmaster0_p & v144608a | !hmaster0_p & v1446404;
assign v15157cf = hbusreq5_p & v15157cd | !hbusreq5_p & !v15157ce;
assign v11e593a = locked_p & v84556a | !locked_p & !v845542;
assign v134d1e3 = stateG3_0_p & v845542 | !stateG3_0_p & !a81304;
assign d2f9d4 = hlock2_p & d2f9d3 | !hlock2_p & d2f9cd;
assign v1668cc0 = stateG3_2_p & v845542 | !stateG3_2_p & !v9f3194;
assign v1446422 = hbusreq0_p & v1446403 | !hbusreq0_p & v1446407;
assign v144583a = hmaster1_p & v1445814 | !hmaster1_p & v1445e28;
assign a6592b = hready_p & a65898 | !hready_p & a6592a;
assign v134d4f2 = hmaster2_p & v845542 | !hmaster2_p & v134d4f1;
assign v134d28f = hgrant0_p & v134d28e | !hgrant0_p & v845542;
assign v1284c8e = hmastlock_p & v1284c8d | !hmastlock_p & v845542;
assign d2fe93 = hbusreq4_p & d2fe92 | !hbusreq4_p & !v845542;
assign v15530a7 = hready_p & v1553306 | !hready_p & v15530a6;
assign v1180b7b = stateG2_p & v88d3e4 | !stateG2_p & v110b6cc;
assign v1445a38 = hlock0 & v1445a37 | !hlock0 & v1445a35;
assign hgrant2 = !v1515857;
assign v1214df4 = hmaster2_p & v1216aad | !hmaster2_p & v1214df3;
assign v140585c = hbusreq2_p & v1405858 | !hbusreq2_p & v140585b;
assign d2fb0f = hbusreq0 & d2fb07 | !hbusreq0 & d2fb0e;
assign d2feab = hmaster1_p & d2feaa | !hmaster1_p & v84555a;
assign v1405b33 = hready_p & v1405b0f | !hready_p & v1405b32;
assign v15161ce = hgrant2_p & v15161cd | !hgrant2_p & !v845542;
assign v16a1c98 = hbusreq1_p & v16a1c97 | !hbusreq1_p & v845542;
assign v1215049 = hgrant5_p & v121546e | !hgrant5_p & v1215048;
assign v14461d4 = hgrant2_p & v14461ce | !hgrant2_p & v14461cf;
assign v1389f86 = hmaster0_p & v1389f85 | !hmaster0_p & !v845542;
assign v12ad56c = hmaster1_p & v12ad56b | !hmaster1_p & !v12ad525;
assign d30141 = hlock5_p & d3013f | !hlock5_p & !d30140;
assign v1445eed = hbusreq5_p & v1445e6e | !hbusreq5_p & v1445eec;
assign v1215c2a = hmaster2_p & v1215c26 | !hmaster2_p & v1215c29;
assign v1515c7c = hburst0 & v15168a9 | !hburst0 & v1515c7b;
assign v138980e = hgrant5_p & v138980d | !hgrant5_p & !v845542;
assign v1215c32 = hgrant5_p & v1215bea | !hgrant5_p & v1215c30;
assign v12acfd8 = hmaster2_p & v12acfc1 | !hmaster2_p & !v12ad67f;
assign v16a205e = hbusreq3 & v16a205a | !hbusreq3 & v16a205d;
assign v14838bb = hgrant5_p & v845558 | !hgrant5_p & v14838ba;
assign v1445edc = hbusreq1 & v1445e59 | !hbusreq1 & v1445e5a;
assign v1405898 = hlock1_p & v140583f | !hlock1_p & v1405854;
assign v10d4018 = hlock2_p & v10d4015 | !hlock2_p & !v10d4017;
assign v138a456 = hbusreq2 & v138a44d | !hbusreq2 & v138a455;
assign v1215bbb = hbusreq3 & v1215bb8 | !hbusreq3 & !v845542;
assign a65ae7 = hmaster2_p & a65ae4 | !hmaster2_p & a662ac;
assign a65495 = hmaster0_p & a658f1 | !hmaster0_p & a658e8;
assign v1215c0b = hbusreq1_p & v1215c09 | !hbusreq1_p & v1215c0a;
assign v1446234 = hbusreq0 & v14463e9 | !hbusreq0 & v14463be;
assign a65690 = hbusreq2_p & a6568e | !hbusreq2_p & a6568f;
assign v1446735 = hlock2 & v144672e | !hlock2 & v1446734;
assign v16693a3 = hbusreq3 & v166939e | !hbusreq3 & v16693a2;
assign a658cc = hbusreq1 & a658c7 | !hbusreq1 & a658cb;
assign v12afa10 = hbusreq5 & v12af9da | !hbusreq5 & v12afa0f;
assign v1214c9a = hbusreq2_p & v1214c94 | !hbusreq2_p & v1214c99;
assign v12150a1 = hgrant4_p & v845542 | !hgrant4_p & !v12150a0;
assign v1405b03 = hgrant1_p & v1405a90 | !hgrant1_p & !v1405b02;
assign v1216b08 = hbusreq2 & v1216aff | !hbusreq2 & v1216b07;
assign v121575d = hbusreq4_p & v121575c | !hbusreq4_p & v845542;
assign v155338d = hlock1 & v1553217 | !hlock1 & v155338c;
assign v14459d8 = hlock0_p & v845542 | !hlock0_p & v14459d7;
assign v1405a7f = hmaster0_p & v1405a7d | !hmaster0_p & v1405a7e;
assign start = v11e5983;
assign d301dd = hbusreq0 & d301d6 | !hbusreq0 & d301dc;
assign v1445dc7 = hlock2 & v1445dc6 | !hlock2 & v1445dbb;
assign v1668c7d = hmaster0_p & v1668c7a | !hmaster0_p & v1668c7c;
assign v138a3f6 = hgrant2_p & v138a3f5 | !hgrant2_p & !v138a3e1;
assign v12ad00d = hbusreq5_p & v12ad5c6 | !hbusreq5_p & !v12ad00c;
assign d306a4 = hbusreq4_p & v845542 | !hbusreq4_p & d306a3;
assign d307fe = hbusreq5_p & d307fd | !hbusreq5_p & !d307fc;
assign v12af5ab = hmaster2_p & v12af5a3 | !hmaster2_p & v12af5aa;
assign v14838b8 = decide_p & v14838b7 | !decide_p & v845558;
assign v1214cf1 = hbusreq0_p & v12166ce | !hbusreq0_p & !v845542;
assign v10d40ce = hgrant2_p & v10d40cc | !hgrant2_p & v10d40cd;
assign v134d21d = hlock2 & v134d213 | !hlock2 & v134d21c;
assign v1214f4f = hmaster1_p & v1214f4e | !hmaster1_p & v1215d79;
assign v1405ae3 = hgrant5_p & v1405ae1 | !hgrant5_p & v1405ae2;
assign d30610 = hbusreq2_p & d3060f | !hbusreq2_p & d3060e;
assign v1515814 = hlock2_p & v1515813 | !hlock2_p & v845542;
assign d3022f = hgrant2_p & d3021d | !hgrant2_p & !d3022e;
assign d301f7 = hbusreq5_p & d301f0 | !hbusreq5_p & d301f6;
assign v1446341 = hmaster0_p & v144633e | !hmaster0_p & v1446340;
assign v16a1d0e = hmaster1_p & v845564 | !hmaster1_p & !v16a2672;
assign v1405862 = hlock1_p & v140583e | !hlock1_p & v14463b1;
assign v1445db9 = hmaster0_p & v144639c | !hmaster0_p & v1445db8;
assign f2f393 = hmaster0_p & f2f378 | !hmaster0_p & f2f392;
assign f2ed8f = hgrant3_p & f2f4c4 | !hgrant3_p & f2ed8e;
assign v14457a6 = hmaster0_p & v144579d | !hmaster0_p & v1445e13;
assign v1668c73 = hmaster1_p & v1668c61 | !hmaster1_p & v1668c72;
assign v15157ff = hbusreq5_p & v15157fe | !hbusreq5_p & !v15157b1;
assign v121504e = hbusreq4_p & v121504d | !hbusreq4_p & !v845542;
assign v1215d6d = hgrant5_p & v12164d6 | !hgrant5_p & v12166c6;
assign d30830 = hmaster0_p & d30826 | !hmaster0_p & d3082f;
assign v14058fc = hgrant4_p & v1446403 | !hgrant4_p & !v14058fb;
assign v16a1af8 = hburst0 & v16a1af6 | !hburst0 & v16a1af7;
assign d2fb8b = hmaster2_p & d2fb69 | !hmaster2_p & d2fb6d;
assign v121543f = hbusreq2_p & v121543e | !hbusreq2_p & v121543d;
assign v16a1950 = hgrant5_p & v845542 | !hgrant5_p & v16a194c;
assign v12ad8ec = hmaster0_p & v12af73f | !hmaster0_p & v12ad8eb;
assign v16a1e25 = hgrant2_p & v16a1d2c | !hgrant2_p & v16a1e24;
assign v1446109 = hbusreq2 & v1446107 | !hbusreq2 & v1446108;
assign d30769 = hmaster1_p & d3072e | !hmaster1_p & d3072c;
assign v1215470 = hmaster1_p & v1215464 | !hmaster1_p & v121546f;
assign v1215030 = hgrant5_p & v1215463 | !hgrant5_p & v121502f;
assign a656cf = hgrant2_p & v845542 | !hgrant2_p & a656ce;
assign v1553141 = hlock1_p & v1553140 | !hlock1_p & v845542;
assign v12161d1 = hgrant1_p & v845542 | !hgrant1_p & v1216037;
assign v155322c = hlock5_p & v155322a | !hlock5_p & v155322b;
assign v1552d55 = hgrant2_p & v1552d54 | !hgrant2_p & v1552d4d;
assign v12aeb72 = hmaster0_p & v845542 | !hmaster0_p & v12aeb71;
assign v1405a92 = hlock0_p & v845542 | !hlock0_p & v1405a91;
assign v1515671 = stateG2_p & v845542 | !stateG2_p & v1668cc0;
assign v1216aea = hready & v1446397 | !hready & !v15168aa;
assign v16a209e = hgrant2_p & v845542 | !hgrant2_p & v16a209c;
assign v134ce48 = hgrant2_p & v134d364 | !hgrant2_p & v134ce47;
assign v134d3cc = hbusreq3 & v134d3ca | !hbusreq3 & v134d3cb;
assign v12160ac = hbusreq2 & v12160a5 | !hbusreq2 & v12160ab;
assign v121506e = hmaster0_p & v1215065 | !hmaster0_p & v121505b;
assign v144674a = hgrant2_p & v1446747 | !hgrant2_p & v1446749;
assign d2fafb = hmaster2_p & d2faed | !hmaster2_p & d2fafa;
assign v14453c6 = hgrant3_p & v1445b30 | !hgrant3_p & v14453c5;
assign v144587b = hmaster2_p & v144586f | !hmaster2_p & v1445879;
assign v12acfb2 = hbusreq0 & v12ad681 | !hbusreq0 & v12af73f;
assign v134ce44 = hgrant5_p & v845542 | !hgrant5_p & v134ce43;
assign v12166f3 = hbusreq5_p & v12166f2 | !hbusreq5_p & v16a2243;
assign v134d499 = hlock0 & v134d497 | !hlock0 & v134d498;
assign d30157 = hlock5_p & d30155 | !hlock5_p & d30156;
assign v16a1da7 = hbusreq2_p & v16a1da5 | !hbusreq2_p & v16a1da6;
assign v15532c1 = hgrant1_p & v1553138 | !hgrant1_p & v845542;
assign v134cedf = hmaster1_p & v134cede | !hmaster1_p & v845542;
assign v1215cf6 = hbusreq5_p & v1215cf5 | !hbusreq5_p & v1215cbd;
assign v144607f = hgrant5_p & v1445fe1 | !hgrant5_p & v144607e;
assign v16a1e30 = hgrant2_p & v16a1ded | !hgrant2_p & v16a1e2f;
assign v140591f = hlock2_p & v140591c | !hlock2_p & v140591e;
assign d2fc3d = hbusreq2_p & d2fbb3 | !hbusreq2_p & d2fc3c;
assign v1214f3b = hbusreq2_p & v1214f3a | !hbusreq2_p & v845542;
assign v144623e = hbusreq2_p & v1446237 | !hbusreq2_p & v144623d;
assign v1446075 = hgrant2_p & v1446039 | !hgrant2_p & v1446074;
assign v16a1bf4 = hgrant5_p & v845542 | !hgrant5_p & v16a1bf3;
assign v1215709 = hmaster0_p & v1215b9a | !hmaster0_p & v1215b98;
assign v1214fbf = hmaster0_p & v121579b | !hmaster0_p & v1214fbe;
assign v1284cc6 = hgrant4_p & v140583c | !hgrant4_p & v1284cc5;
assign v12ad5f5 = hlock2_p & v12ad5f2 | !hlock2_p & !v12ad5f4;
assign v1216a7d = hbusreq3 & v1216a72 | !hbusreq3 & v1216a7c;
assign v12ad54c = hmaster2_p & a658ca | !hmaster2_p & !v12ad51c;
assign f2f231 = hmaster2_p & f2f22a | !hmaster2_p & f2f230;
assign v16a1cd6 = hmaster1_p & v16a1cd5 | !hmaster1_p & v16a2672;
assign v1553932 = hburst1_p & v1553931 | !hburst1_p & v155392f;
assign v1215777 = hgrant5_p & v1215b8a | !hgrant5_p & v1215776;
assign v1515783 = hgrant5_p & v10d3ffa | !hgrant5_p & v1515781;
assign v1215cd4 = hbusreq0 & v1215ccf | !hbusreq0 & v1215cd3;
assign d3023c = hbusreq3 & d30238 | !hbusreq3 & v845542;
assign v12ad55d = hmaster1_p & v12ad541 | !hmaster1_p & v12ad54f;
assign v10d4054 = hmaster1_p & v10d4053 | !hmaster1_p & v10d3ffb;
assign v1216322 = hmaster0_p & v1216321 | !hmaster0_p & v1216302;
assign v121536d = hmaster0_p & v1215365 | !hmaster0_p & v845547;
assign v144664d = hgrant2_p & v144663c | !hgrant2_p & v144664c;
assign v121540a = hbusreq2 & v12153fe | !hbusreq2 & v1215409;
assign v16a1d3a = hmaster2_p & v16a1d39 | !hmaster2_p & v16a206f;
assign d2fbe1 = hmaster2_p & d2fbd5 | !hmaster2_p & d2fbe0;
assign d3012c = hgrant2_p & v84555a | !hgrant2_p & d30120;
assign v1446270 = hbusreq2_p & v144626b | !hbusreq2_p & v144626f;
assign f2f363 = hmaster2_p & f2f362 | !hmaster2_p & !v845542;
assign v12aee5c = decide_p & v12af9b6 | !decide_p & v12afe76;
assign v144672f = hmaster0_p & v1446440 | !hmaster0_p & v1446657;
assign d3029b = hbusreq3 & d3029a | !hbusreq3 & v845542;
assign v1405b4b = hbusreq4_p & v1405ad4 | !hbusreq4_p & v1405b4a;
assign v121482e = jx0_p & v1215ddf | !jx0_p & v121482d;
assign v1446439 = hbusreq1 & v144640a | !hbusreq1 & v1446438;
assign v1446749 = hmaster1_p & v1446748 | !hmaster1_p & v1446630;
assign v138a333 = hmaster2_p & v84556a | !hmaster2_p & !v138a332;
assign v1445dba = hmaster1_p & v1445db9 | !hmaster1_p & v1445da4;
assign d3025f = hbusreq2 & d3025b | !hbusreq2 & d3025e;
assign v1668ca0 = hbusreq5_p & v1668c9e | !hbusreq5_p & v1668c9f;
assign v10d4074 = hgrant1_p & v10d3fe5 | !hgrant1_p & !v10d4073;
assign v16a1979 = hgrant2_p & v845542 | !hgrant2_p & !v16a1977;
assign v144578e = hmaster0_p & v144578b | !hmaster0_p & v1445e0c;
assign a653de = hbusreq4_p & a653dd | !hbusreq4_p & v845542;
assign v12150b2 = decide_p & v121545d | !decide_p & v12150b1;
assign v16a1843 = hmaster0_p & v16a1840 | !hmaster0_p & v16a1842;
assign a6544b = hbusreq2_p & a6543c | !hbusreq2_p & a65449;
assign v138a3c9 = hlock5_p & v138a3c8 | !hlock5_p & !v151579c;
assign d30635 = hmaster1_p & d3060c | !hmaster1_p & d30608;
assign v1445d8d = hbusreq5_p & v1445d86 | !hbusreq5_p & v1445d8c;
assign v1215c16 = hmaster2_p & v1215c15 | !hmaster2_p & v1215c0d;
assign v12160a4 = hlock2_p & v12160a2 | !hlock2_p & v12160a3;
assign v15157aa = hmaster2_p & v1515795 | !hmaster2_p & v15157a9;
assign f2f375 = hmaster2_p & f2f374 | !hmaster2_p & f2f234;
assign d307bb = hgrant4_p & d307b0 | !hgrant4_p & v845542;
assign v16a19c3 = hmaster1_p & v16a19b1 | !hmaster1_p & v16a1f96;
assign v134ce41 = hbusreq1 & v134ce3f | !hbusreq1 & v134ce40;
assign v1668dbb = hgrant5_p & v845542 | !hgrant5_p & !v1668d37;
assign v1446147 = hlock2 & v1446125 | !hlock2 & v1446145;
assign v121616f = hmaster0_p & v1216135 | !hmaster0_p & v121616e;
assign d2fd11 = hbusreq2_p & d2fd10 | !hbusreq2_p & d302d6;
assign d3077f = hlock2_p & d3077e | !hlock2_p & !d30707;
assign f2e4d3 = decide_p & f2e4d2 | !decide_p & f2f23c;
assign a658bd = hmastlock_p & a658bc | !hmastlock_p & v845542;
assign v134d388 = hgrant5_p & v845542 | !hgrant5_p & v134d387;
assign v1216573 = hbusreq5_p & v1216572 | !hbusreq5_p & v845542;
assign v14458b3 = hbusreq2_p & v14458b0 | !hbusreq2_p & v14458b2;
assign v1216073 = hmaster0_p & v1216068 | !hmaster0_p & v121605f;
assign d2fbf5 = hgrant4_p & d2fbf4 | !hgrant4_p & d2fbd3;
assign v12af228 = hmaster0_p & v12af9c3 | !hmaster0_p & v12af227;
assign v1515857 = jx0_p & v151621e | !jx0_p & v1515856;
assign v1216136 = hbusreq4 & v121611d | !hbusreq4 & v845547;
assign v12153c3 = hbusreq2_p & v12153c0 | !hbusreq2_p & v12153c2;
assign v1215d30 = hgrant5_p & v1216a90 | !hgrant5_p & v1216589;
assign v121573e = hmaster2_p & v1215721 | !hmaster2_p & v121573d;
assign d307cc = hbusreq1_p & d307cb | !hbusreq1_p & d30661;
assign a662c0 = hbusreq1_p & a66278 | !hbusreq1_p & a6627b;
assign v144583f = hlock3 & v144582d | !hlock3 & v144583e;
assign v1216069 = hmaster0_p & v121604c | !hmaster0_p & v1216068;
assign v1215cbd = hmaster2_p & v1215cba | !hmaster2_p & v1215cbc;
assign stateG10_1 = !v11ac6ca;
assign v16a1ae3 = hgrant2_p & v845542 | !hgrant2_p & !v16a1ae0;
assign d30675 = hmaster1_p & d30674 | !hmaster1_p & d305db;
assign f2f334 = hmaster1_p & f2f2e4 | !hmaster1_p & !f2f330;
assign v1445b90 = hmaster1_p & v1446313 | !hmaster1_p & v1445b8d;
assign d2fbbf = hlock2_p & d2fbbe | !hlock2_p & d2fbbb;
assign v1445b0f = hmaster1_p & v1445ae7 | !hmaster1_p & v144591b;
assign v1445fbd = hmaster0_p & v1445fbc | !hmaster0_p & v1445f9d;
assign v14466f1 = hmaster1_p & v14466f0 | !hmaster1_p & v1446436;
assign v1215fc1 = hbusreq2 & v1215fba | !hbusreq2 & v1215fc0;
assign v11e593d = hmaster1_p & v11e593c | !hmaster1_p & v845542;
assign v1214c2d = hmaster2_p & v1214c29 | !hmaster2_p & d2fbe5;
assign v1445fb8 = stateG10_5_p & v1445f89 | !stateG10_5_p & !v1445fb7;
assign v1405ab1 = hmaster0_p & v1405aa3 | !hmaster0_p & v1405ab0;
assign d8078b = hbusreq1_p & d80733 | !hbusreq1_p & !d8078a;
assign v1668ceb = hgrant2_p & v1668ce7 | !hgrant2_p & v1668cea;
assign v1445e9f = hmaster2_p & v1446609 | !hmaster2_p & v1445e9e;
assign v1214e80 = hmaster1_p & v1214e62 | !hmaster1_p & v1215bc2;
assign v1216706 = hbusreq2_p & v1216705 | !hbusreq2_p & v12166fa;
assign f2e503 = hbusreq3_p & f2e4fa | !hbusreq3_p & f2e502;
assign v1445837 = hgrant2_p & v1445835 | !hgrant2_p & v1445836;
assign d2fbad = hbusreq2 & d2fba9 | !hbusreq2 & d2fbac;
assign d30787 = hbusreq1 & d30786 | !hbusreq1 & v845542;
assign v1668d15 = hmaster2_p & a65851 | !hmaster2_p & v845542;
assign v12ad322 = hgrant4_p & d3068f | !hgrant4_p & !v12ad321;
assign v14058b4 = hmaster2_p & v140583c | !hmaster2_p & v140589a;
assign v155314e = hmaster0_p & v1553146 | !hmaster0_p & v155314d;
assign v134d37f = hgrant4_p & v134d37e | !hgrant4_p & v845542;
assign v12ad4ca = hlock0_p & v1515609 | !hlock0_p & d2fbe5;
assign d301bc = hbusreq1_p & v845542 | !hbusreq1_p & d306d4;
assign v15168f3 = hmastlock_p & v15168f2 | !hmastlock_p & v845542;
assign v14461dc = hlock3 & v14461c1 | !hlock3 & v14461db;
assign v16a12c0 = hmaster1_p & v16a1a94 | !hmaster1_p & v16a1f96;
assign v121678e = hready_p & v12165b4 | !hready_p & v121678d;
assign d2fbd3 = hgrant0_p & v845542 | !hgrant0_p & d2fb4d;
assign v1446195 = hgrant2_p & v1446194 | !hgrant2_p & v144618f;
assign v12af7e2 = decide_p & v12af7e1 | !decide_p & v845542;
assign v15155fb = hbusreq0 & v15155fa | !hbusreq0 & v845542;
assign f2f3bf = hmaster2_p & f2f2aa | !hmaster2_p & v845542;
assign a66292 = stateG3_2_p & v845542 | !stateG3_2_p & v1553931;
assign v134ce52 = hbusreq1 & v134ce34 | !hbusreq1 & v134ce35;
assign v14465d8 = hgrant1_p & v1446406 | !hgrant1_p & v14465d7;
assign v1389818 = hmaster1_p & v138980a | !hmaster1_p & v1389817;
assign v1215d07 = hbusreq2_p & v1215cfc | !hbusreq2_p & !v1215d06;
assign d30124 = hbusreq4_p & d30123 | !hbusreq4_p & v845542;
assign v1445926 = hlock5 & v1445916 | !hlock5 & v1445925;
assign v151580d = hmaster0_p & v151580c | !hmaster0_p & v1515639;
assign a65ae5 = hgrant5_p & v845542 | !hgrant5_p & a65ae4;
assign v121545e = hbusreq4 & v12164cf | !hbusreq4 & v845547;
assign v15157a6 = hmaster2_p & v151561c | !hmaster2_p & v845570;
assign v14465d1 = hbusreq1_p & v14465b2 | !hbusreq1_p & v14465d0;
assign v14461fa = hgrant2_p & v14461d7 | !hgrant2_p & v14461f2;
assign v12ad546 = hbusreq2_p & v12ad543 | !hbusreq2_p & v12ad545;
assign v1215d2c = hmaster1_p & v1215d27 | !hmaster1_p & v1215d2b;
assign v12aec48 = hmaster0_p & v12afe47 | !hmaster0_p & v12aec47;
assign v134d4f3 = hgrant5_p & v134d36a | !hgrant5_p & v134d4f2;
assign v16a1b03 = hmaster1_p & v16a1afd | !hmaster1_p & v16a2672;
assign d3084d = hbusreq5_p & d307f7 | !hbusreq5_p & d3084c;
assign v144643c = hbusreq5_p & v144643a | !hbusreq5_p & v144643b;
assign v1284d0a = hgrant0_p & v140587c | !hgrant0_p & !v1284d09;
assign v144543b = hbusreq5 & v1445433 | !hbusreq5 & v144543a;
assign f2f4be = hmaster0_p & f2f220 | !hmaster0_p & v845542;
assign v1668d93 = hmaster0_p & v1668d92 | !hmaster0_p & v1668d7f;
assign v16a1cf8 = hbusreq0 & v16a1cf7 | !hbusreq0 & v16a1be1;
assign d308f3 = hmaster2_p & v845542 | !hmaster2_p & v84554e;
assign v144613c = hlock2 & v1446138 | !hlock2 & v144613b;
assign v155309d = hbusreq2_p & v155309b | !hbusreq2_p & v155309c;
assign v14463a9 = hbusreq0 & v14463a7 | !hbusreq0 & v14463a8;
assign v1446088 = hmaster2_p & v144639c | !hmaster2_p & v1446087;
assign v1215c44 = hbusreq5_p & v1215c42 | !hbusreq5_p & !v1215c43;
assign v1214ca2 = hbusreq5 & v1214c86 | !hbusreq5 & v1214ca1;
assign v12af5a2 = hbusreq1_p & v12afe45 | !hbusreq1_p & v12afe61;
assign v16a12ee = hmaster1_p & v16a12ed | !hmaster1_p & v16a1d53;
assign v134ce60 = hbusreq5_p & v134ce3a | !hbusreq5_p & v134ce5f;
assign v1445373 = hbusreq2_p & v1445363 | !hbusreq2_p & v1445372;
assign v16a1383 = hbusreq0 & v16a1a93 | !hbusreq0 & !v16a1ac9;
assign v151563b = hmaster1_p & v151563a | !hmaster1_p & v10d3ffb;
assign v151578f = hmastlock_p & v151578e | !hmastlock_p & !v845542;
assign d30142 = hgrant5_p & v84555a | !hgrant5_p & d300f3;
assign v12153f0 = hmaster1_p & v12153ef | !hmaster1_p & v12153ec;
assign d2fba3 = hlock2_p & d2fba2 | !hlock2_p & d2fb9f;
assign v16a1e2f = hmaster1_p & v16a1e27 | !hmaster1_p & !v16a2672;
assign v14459eb = hmaster2_p & v14459db | !hmaster2_p & v14459e7;
assign bf1f8a = hgrant3_p & bf1f57 | !hgrant3_p & bf1f89;
assign v1668dcf = hgrant5_p & v845542 | !hgrant5_p & !v1668d86;
assign v138a032 = hmaster0_p & v138a02e | !hmaster0_p & !v1389de1;
assign v14058e9 = hgrant4_p & v140587c | !hgrant4_p & v14058e8;
assign v1445af3 = hlock2 & v1445af2 | !hlock2 & v1445aec;
assign v1215301 = hbusreq2 & v12152fa | !hbusreq2 & v1215300;
assign v12167a2 = hmaster1_p & v12167a1 | !hmaster1_p & v1216a9b;
assign v16a16a2 = hgrant2_p & v845542 | !hgrant2_p & !v16a169f;
assign v1216166 = hbusreq1 & v1216165 | !hbusreq1 & v845542;
assign v1552d7a = stateA1_p & v1553934 | !stateA1_p & v1553933;
assign v16a1438 = hgrant1_p & v84554d | !hgrant1_p & v16a1437;
assign v14459ca = hgrant0_p & v14458e2 | !hgrant0_p & v144586f;
assign v1389f8d = hbusreq5_p & v1389f8c | !hbusreq5_p & v845542;
assign v1445ad1 = hbusreq2_p & v1445acf | !hbusreq2_p & v1445ad0;
assign v12160c1 = hbusreq2_p & v12160c0 | !hbusreq2_p & v12160bf;
assign v151582e = hbusreq3 & v1515829 | !hbusreq3 & v151582d;
assign v1445557 = jx1_p & v14453c8 | !jx1_p & v1445556;
assign v14462a3 = hbusreq5 & v14462a1 | !hbusreq5 & v14462a2;
assign v1284cdb = hgrant4_p & v140584b | !hgrant4_p & !v1284cda;
assign a6546c = hbusreq1 & a658b6 | !hbusreq1 & !a6546a;
assign v14058c9 = hgrant5_p & v1405897 | !hgrant5_p & v14058c8;
assign f2f23c = hgrant2_p & v845542 | !hgrant2_p & f2f23b;
assign v1445fbc = hlock0 & v1445fbb | !hlock0 & v1445fba;
assign a6561f = hbusreq1_p & a65371 | !hbusreq1_p & a6561d;
assign d3069f = hbusreq2_p & d30631 | !hbusreq2_p & d3069e;
assign d2f973 = hmaster2_p & d2f96c | !hmaster2_p & !d2f972;
assign v14466dc = hmaster0_p & v14463f6 | !hmaster0_p & v14463c9;
assign v1389449 = hmaster0_p & v1389448 | !hmaster0_p & v845542;
assign v134d3bc = hready_p & v134d34f | !hready_p & v134d3bb;
assign v12162fa = hbusreq1 & v1216aad | !hbusreq1 & v1216ab9;
assign v1215d3d = hmaster0_p & v1668da6 | !hmaster0_p & v12165a8;
assign a656bd = hmaster2_p & a66299 | !hmaster2_p & a6628b;
assign v144672a = hmaster0_p & v1446440 | !hmaster0_p & v144663a;
assign v16a1cf0 = hmaster1_p & v16a1cef | !hmaster1_p & v16a1bdb;
assign v12ad50c = hlock3_p & v12ad4ef | !hlock3_p & v12ad50b;
assign v138a394 = hbusreq5_p & v138a393 | !hbusreq5_p & !v845542;
assign v138a402 = hlock5_p & v84557c | !hlock5_p & !v845542;
assign v140583e = hmastlock_p & v85e70d | !hmastlock_p & !v845542;
assign d2fec6 = hmaster0_p & d2febe | !hmaster0_p & d2fec5;
assign v1284d2f = hmaster1_p & v1284d2e | !hmaster1_p & v140584d;
assign v16a1abf = hbusreq2_p & v16a2673 | !hbusreq2_p & v16a1abe;
assign v138a3ef = hgrant2_p & v138a3e5 | !hgrant2_p & !v138a3ee;
assign v16a1e64 = hmaster0_p & v16a1e5f | !hmaster0_p & v16a1e63;
assign v16a1984 = hbusreq5 & v16a197a | !hbusreq5 & v16a1983;
assign a653bf = hbusreq5_p & a653ba | !hbusreq5_p & !a653bd;
assign d305ee = stateA1_p & a658a5 | !stateA1_p & a658a3;
assign v16a197d = hgrant5_p & v845542 | !hgrant5_p & !v16a1973;
assign v134d26b = hlock3 & v134d264 | !hlock3 & v134d26a;
assign v1445b8b = hbusreq0 & v1445b8a | !hbusreq0 & v14462f3;
assign v134d37c = hlock0 & v134d37b | !hlock0 & v134d37a;
assign v121623f = hmaster0_p & v1216236 | !hmaster0_p & v121622b;
assign d2fb93 = hmaster0_p & d2fb8c | !hmaster0_p & d2fb85;
assign d3067d = hmaster1_p & v845542 | !hmaster1_p & d3067c;
assign v1552d96 = decide_p & v15532bf | !decide_p & v1552d95;
assign a65387 = hgrant4_p & v845570 | !hgrant4_p & !a65384;
assign v1445fde = hmaster0_p & v1445fd3 | !hmaster0_p & v1445fdd;
assign v138a3c0 = hlock3_p & v138a392 | !hlock3_p & v138a3bf;
assign d2fc11 = hmaster0_p & d2fc10 | !hmaster0_p & d2fbfc;
assign v151621c = hbusreq3_p & v1516215 | !hbusreq3_p & v151621b;
assign v134d450 = hmaster1_p & v134d369 | !hmaster1_p & v134d44f;
assign v12ad4fc = hbusreq4_p & v10d3fd8 | !hbusreq4_p & !v12ad4f6;
assign v12160b7 = hbusreq2_p & v12160b6 | !hbusreq2_p & v12160b5;
assign v14466d4 = hlock2 & v14466d3 | !hlock2 & v14466cf;
assign v12152e8 = hlock2_p & v12152e5 | !hlock2_p & !v12152e7;
assign bf1fa7 = hbusreq2_p & bf1f71 | !hbusreq2_p & !bf1fa6;
assign v1216226 = hgrant2_p & v1216202 | !hgrant2_p & v1216225;
assign v1445b27 = hlock3 & v1445af2 | !hlock3 & v1445b26;
assign v1389fe9 = hgrant2_p & v845542 | !hgrant2_p & !v1389fe8;
assign v1445a04 = stateG10_5_p & v14459ff | !stateG10_5_p & v1445a03;
assign v1552d95 = hbusreq2_p & v1552d90 | !hbusreq2_p & v1552d94;
assign v138a092 = hgrant3_p & v138a076 | !hgrant3_p & v138a091;
assign v155342e = hbusreq2_p & v1553158 | !hbusreq2_p & v155342d;
assign v1215cb3 = hlock5_p & v1215cb1 | !hlock5_p & !v1215cb2;
assign v1215c4e = hgrant2_p & v1215c4d | !hgrant2_p & v1215c36;
assign v1445aba = hbusreq2_p & v1445ab1 | !hbusreq2_p & v1445ab9;
assign v14466d5 = hbusreq2 & v14466cf | !hbusreq2 & v14466d4;
assign v1552d7b = hmastlock_p & v1552d7a | !hmastlock_p & v845542;
assign v16a1329 = hbusreq0 & v16a1328 | !hbusreq0 & v845568;
assign v134d4dd = hmaster1_p & v134d280 | !hmaster1_p & v134d4dc;
assign v16a1daf = hready_p & v845555 | !hready_p & v16a1dae;
assign d30102 = hlock5_p & d30100 | !hlock5_p & d30101;
assign d3083b = hbusreq0 & d30836 | !hbusreq0 & d3083a;
assign v1214de2 = hbusreq2 & v1214de1 | !hbusreq2 & v845542;
assign v16a1d02 = hready_p & v16a1d00 | !hready_p & v16a1d01;
assign v15530a8 = hgrant3_p & v155321c | !hgrant3_p & v15530a7;
assign v134d278 = hready_p & v134d1e2 | !hready_p & v134d277;
assign d3018d = hmaster2_p & d30718 | !hmaster2_p & !v16693aa;
assign a654c6 = hbusreq5 & a654ac | !hbusreq5 & a654c5;
assign v12ad5cc = hmaster2_p & v12ad5cb | !hmaster2_p & v12ad5c4;
assign v121534c = hmaster2_p & v1215345 | !hmaster2_p & v121534b;
assign v14461f2 = hmaster1_p & v1446092 | !hmaster1_p & v14460cf;
assign v1445aa8 = hbusreq2 & v1445aa4 | !hbusreq2 & v1445aa7;
assign d2f96f = hmaster2_p & d2f96c | !hmaster2_p & !d2f96e;
assign d2fad0 = hmaster1_p & d2facf | !hmaster1_p & !d2fea2;
assign v16a20a2 = hgrant2_p & v845542 | !hgrant2_p & v16a20a1;
assign v12acfd9 = hbusreq5_p & v12ad54b | !hbusreq5_p & v12acfd8;
assign v1214e74 = hmaster1_p & v1214dea | !hmaster1_p & v1214e73;
assign v14457a5 = hbusreq2_p & v144579f | !hbusreq2_p & v14457a4;
assign v1668e04 = hbusreq3_p & v1668e03 | !hbusreq3_p & !v1668c39;
assign v14465b0 = hgrant1_p & v144639c | !hgrant1_p & v14465af;
assign v1446705 = hmaster0_p & v1446657 | !hmaster0_p & v1446440;
assign f2f32e = hmaster2_p & f2f2e7 | !hmaster2_p & f2f21f;
assign v134cd7c = hgrant5_p & v134cd7b | !hgrant5_p & v134cd5b;
assign v1215796 = hgrant5_p & v121578f | !hgrant5_p & v121574c;
assign v1216023 = hbusreq0_p & v845547 | !hbusreq0_p & v121601f;
assign v14460ae = hmaster1_p & v14465aa | !hmaster1_p & v1445ffc;
assign v1215322 = hgrant2_p & v121531f | !hgrant2_p & v1215321;
assign v134d27f = hmaster2_p & v134d27e | !hmaster2_p & v845542;
assign d300e6 = hbusreq1 & d2fe9c | !hbusreq1 & v84555a;
assign v144605d = hbusreq1_p & v1446602 | !hbusreq1_p & v144660e;
assign v1445362 = hmaster1_p & v1445361 | !hmaster1_p & v1445a32;
assign v1445990 = busreq_p & v146d169 | !busreq_p & !v845588;
assign v16a16b3 = hready_p & v16a16b1 | !hready_p & v16a16b2;
assign v151571a = hburst0 & v1515718 | !hburst0 & v1515719;
assign v12150bb = hmaster0_p & v1215019 | !hmaster0_p & v12153b5;
assign v1216243 = hmaster1_p & v1216236 | !hmaster1_p & v1216224;
assign v144619a = hlock3 & v144617b | !hlock3 & v1446198;
assign v16a1af9 = hmastlock_p & v16a1af8 | !hmastlock_p & !v845542;
assign v134cebf = hbusreq5 & v134d270 | !hbusreq5 & v134cebe;
assign v1215b7e = hmaster2_p & v1215b76 | !hmaster2_p & v1215b7d;
assign v134d528 = hbusreq3 & v134d526 | !hbusreq3 & v134d527;
assign v10d4034 = hgrant5_p & v10d4029 | !hgrant5_p & !v10d4033;
assign a658fd = hmaster0_p & a658ee | !hmaster0_p & a658e8;
assign v12af22c = decide_p & v12af22b | !decide_p & v12afe76;
assign v16a1bb9 = hready & v16a1bb8 | !hready & v845542;
assign v1446048 = hgrant1_p & v1446046 | !hgrant1_p & v1446047;
assign v10d3fed = hmaster1_p & v10d3fec | !hmaster1_p & v10d3fe9;
assign v14465e1 = hgrant1_p & v144639c | !hgrant1_p & v14465e0;
assign v134d431 = hlock0 & v134d42a | !hlock0 & v134d430;
assign v1389e31 = hmaster0_p & v1389e2d | !hmaster0_p & v1389e27;
assign v1214e6e = hbusreq1_p & v1216aea | !hbusreq1_p & v1216ab9;
assign v12160d0 = hbusreq1 & v12164cf | !hbusreq1 & v845547;
assign v1214f02 = hgrant5_p & v845542 | !hgrant5_p & v1214ed3;
assign v16a1d4a = hbusreq0 & v16a1d49 | !hbusreq0 & v16a1d45;
assign v16a1447 = hready_p & v16a1446 | !hready_p & !v16a2065;
assign a653ae = hbusreq1_p & a653ac | !hbusreq1_p & !a653ad;
assign v16a1d53 = hbusreq0 & v16a207a | !hbusreq0 & v16a208b;
assign v12ad572 = hmaster0_p & v12ad531 | !hmaster0_p & v12ad517;
assign v144617f = hbusreq2_p & v1446165 | !hbusreq2_p & v144617e;
assign v15156e4 = hbusreq5_p & v15156e3 | !hbusreq5_p & v1668cc8;
assign v1405937 = hmaster0_p & v140584f | !hmaster0_p & v14058db;
assign v14458ff = hmaster2_p & v14458d2 | !hmaster2_p & v14458e8;
assign v14463f3 = hmaster2_p & v144639c | !hmaster2_p & v14463f2;
assign v1446657 = hlock0 & v1446656 | !hlock0 & v1446655;
assign v1389e27 = hbusreq5_p & v1389e26 | !hbusreq5_p & !v845542;
assign v1216710 = hgrant2_p & v12166ff | !hgrant2_p & v121670f;
assign v1515775 = hmaster2_p & v1515767 | !hmaster2_p & v1515774;
assign a65441 = hgrant5_p & v845558 | !hgrant5_p & !a653fd;
assign v12afe61 = hgrant4_p & v845542 | !hgrant4_p & !v12afe60;
assign v1214c62 = hmaster2_p & v1214c61 | !hmaster2_p & v1214c5c;
assign v12163ac = hlock2_p & v12163aa | !hlock2_p & v12163ab;
assign v1445a0e = hlock4 & v14459bc | !hlock4 & v14465ad;
assign v1445788 = hbusreq2 & v1445781 | !hbusreq2 & v1445787;
assign v16a1d25 = hbusreq3 & v16a1d21 | !hbusreq3 & !v16a1d0f;
assign v121618a = hbusreq2_p & v1216188 | !hbusreq2_p & v1216189;
assign v1446316 = hbusreq2_p & v1446301 | !hbusreq2_p & v1446315;
assign v1445537 = hbusreq5 & v144552a | !hbusreq5 & v1445536;
assign v1445e93 = hgrant1_p & v1445dfc | !hgrant1_p & v1445e8d;
assign d306f6 = hbusreq1_p & d306f5 | !hbusreq1_p & !v845542;
assign v1445f96 = hmaster2_p & v1445f93 | !hmaster2_p & v1445f95;
assign v1445397 = hmaster1_p & v144536a | !hmaster1_p & v144591b;
assign v16a1ad1 = hmaster1_p & v16a1ad0 | !hmaster1_p & v16a1f96;
assign v1405903 = decide_p & v140587b | !decide_p & v1405902;
assign v144586b = hbusreq3_p & v1445f20 | !hbusreq3_p & v144586a;
assign v14465ba = hmaster2_p & v144639c | !hmaster2_p & v14465b9;
assign d305dc = hmaster1_p & d305d8 | !hmaster1_p & d305db;
assign d307b1 = hlock0_p & d306d4 | !hlock0_p & a65861;
assign v138a319 = hbusreq2_p & v138a315 | !hbusreq2_p & v138a318;
assign v134d230 = hlock2_p & v134d22d | !hlock2_p & v134d22f;
assign f2f3a9 = hmaster0_p & f2f35d | !hmaster0_p & f2f3a8;
assign v12af986 = hmaster2_p & d30690 | !hmaster2_p & !v12af985;
assign v146d169 = stateG2_p & v845542 | !stateG2_p & !v845588;
assign v138a38e = hlock5_p & v845568 | !hlock5_p & !v845542;
assign v1214c68 = hbusreq1_p & v1214c66 | !hbusreq1_p & v1214c67;
assign d2fbc9 = hlock2_p & d2fbc8 | !hlock2_p & v84554a;
assign v1445aeb = hmaster1_p & v1445aea | !hmaster1_p & v14458fd;
assign v1214bc3 = hmaster1_p & v12153b1 | !hmaster1_p & v12153a9;
assign d301d5 = hlock5_p & d301d3 | !hlock5_p & !d301d4;
assign v1214d5b = hbusreq3 & v1214d54 | !hbusreq3 & v1214d5a;
assign v1405a9a = hmaster1_p & v1405a8a | !hmaster1_p & !v1405a94;
assign v1214c69 = hbusreq0_p & v121655c | !hbusreq0_p & v845542;
assign v1553097 = hbusreq5_p & v1553053 | !hbusreq5_p & v1553096;
assign v1215c83 = hmaster0_p & v1215c81 | !hmaster0_p & v1215c82;
assign v16a2081 = hmaster2_p & v16a207e | !hmaster2_p & v16a2080;
assign v1405838 = stateA1_p & v845542 | !stateA1_p & !v146d169;
assign v134d208 = hmaster0_p & v134d203 | !hmaster0_p & v134d207;
assign v1446426 = hmaster2_p & v144641f | !hmaster2_p & v1446425;
assign v16a1d5d = hmaster0_p & v16a1d5a | !hmaster0_p & v16a1d5c;
assign v121545f = hbusreq4_p & v121545e | !hbusreq4_p & v845547;
assign v134ce75 = hbusreq2 & v134ce73 | !hbusreq2 & v134ce74;
assign v16a1d35 = hbusreq5 & v16a1d30 | !hbusreq5 & v16a1d34;
assign v12ad008 = hbusreq0 & v12ad007 | !hbusreq0 & v12afa0a;
assign v1446459 = hlock3 & v1446455 | !hlock3 & v1446457;
assign v1405b11 = hmaster1_p & v1405b10 | !hmaster1_p & !v1405ac8;
assign v134d3e4 = hbusreq2_p & v134d296 | !hbusreq2_p & v134d3e3;
assign v1216ae5 = hlock5_p & v1216adb | !hlock5_p & v1216ae4;
assign v144578a = hbusreq0 & v1445789 | !hbusreq0 & v1445776;
assign v1215fba = hbusreq2_p & v1215fb5 | !hbusreq2_p & v1215fb9;
assign v1515640 = hmaster0_p & v151563f | !hmaster0_p & v845542;
assign d2fbc2 = hbusreq5 & d2fbb9 | !hbusreq5 & d2fbc1;
assign a654ad = hmaster2_p & a6546a | !hmaster2_p & !a6546d;
assign a658a9 = stateG2_p & v845542 | !stateG2_p & a658a8;
assign v1515608 = jx2_p & v15155e5 | !jx2_p & v1515607;
assign v1445905 = hbusreq2_p & v14458fe | !hbusreq2_p & v1445904;
assign v12acffc = hgrant4_p & v12ad59e | !hgrant4_p & !v12acffb;
assign v14463b3 = hlock0_p & v144639c | !hlock0_p & !v14463b2;
assign d2fea9 = hmaster2_p & v84555a | !hmaster2_p & !d2fea8;
assign v1446138 = hbusreq2_p & v1446135 | !hbusreq2_p & v1446137;
assign v1215b99 = hlock4_p & v16a19a4 | !hlock4_p & !v845542;
assign v14463c6 = hbusreq5_p & v14463c4 | !hbusreq5_p & v14463c5;
assign d30715 = stateA1_p & a658a7 | !stateA1_p & !d30714;
assign v14461fd = hbusreq2 & v14461f5 | !hbusreq2 & v14461fc;
assign v1405b1b = hgrant1_p & v1405a88 | !hgrant1_p & !v1405b1a;
assign v1214cc6 = hready & v1214cc5 | !hready & v1216593;
assign v12ad60d = hgrant5_p & v12ad60c | !hgrant5_p & !v12ad5c5;
assign v1214f71 = hbusreq2 & v1214f70 | !hbusreq2 & v12164e7;
assign v1445ac2 = hmaster0_p & v14458aa | !hmaster0_p & v144639c;
assign v1215d37 = hgrant5_p & v1215d35 | !hgrant5_p & !v1215d36;
assign d2fb7b = hmaster0_p & d2fb75 | !hmaster0_p & d2fb7a;
assign d30814 = hbusreq2 & d30808 | !hbusreq2 & d30813;
assign v14462ee = hgrant5_p & v14462eb | !hgrant5_p & v14462ed;
assign d300ec = hbusreq5_p & d300e3 | !hbusreq5_p & d300eb;
assign v1445530 = hgrant2_p & v14454e9 | !hgrant2_p & v144552f;
assign v151562b = stateG3_2_p & v845542 | !stateG3_2_p & !a65883;
assign v1215468 = hmaster2_p & v1215bac | !hmaster2_p & v1215467;
assign d2fc79 = hbusreq2_p & d2fc16 | !hbusreq2_p & d2fc77;
assign d2f9d9 = hready_p & d2f987 | !hready_p & !d2f9d8;
assign v15157df = hgrant5_p & v845542 | !hgrant5_p & !v1515733;
assign v1216000 = hbusreq1 & v1215fff | !hbusreq1 & v845542;
assign v1215bec = hmaster1_p & v1215be5 | !hmaster1_p & !v1215beb;
assign v1215d31 = hmaster0_p & v1215d2f | !hmaster0_p & v1215d30;
assign v1668d2c = hgrant5_p & v1668d2b | !hgrant5_p & v1668d29;
assign v1445bee = hmaster1_p & v1445bed | !hmaster1_p & v1446329;
assign v16a1bff = hmaster0_p & v16a1bfe | !hmaster0_p & v16a1bfc;
assign d308a2 = hmaster2_p & d3089f | !hmaster2_p & d308a1;
assign v14459e6 = hbusreq1_p & v14465b2 | !hbusreq1_p & v14459cb;
assign v1284d42 = hmaster0_p & v1405859 | !hmaster0_p & v1284c90;
assign v1445a26 = hbusreq0_p & v144641b | !hbusreq0_p & v1446406;
assign v12ad4c4 = hmaster1_p & v12af7f7 | !hmaster1_p & v12ad4c3;
assign d2fbdf = hbusreq1_p & d2fbde | !hbusreq1_p & v84554a;
assign v134d52e = hmaster0_p & v134d4df | !hmaster0_p & v845542;
assign v16a1d26 = hmaster1_p & v16a1d1a | !hmaster1_p & !v16a1f96;
assign v12161b1 = hmaster1_p & v12161a2 | !hmaster1_p & v12161ae;
assign v1668c1e = hbusreq5_p & v1668c1d | !hbusreq5_p & v845542;
assign v1445552 = decide_p & v144553f | !decide_p & v1445551;
assign v1214c48 = hbusreq4_p & v1214c47 | !hbusreq4_p & v16a19a4;
assign v1284d49 = hbusreq4_p & v1284cc5 | !hbusreq4_p & v1284d48;
assign v1445a18 = hlock1 & v1445a17 | !hlock1 & v1445a14;
assign d3021d = hmaster1_p & d3021c | !hmaster1_p & !d301ca;
assign v1445ef2 = hgrant2_p & v1445ee8 | !hgrant2_p & v1445ef1;
assign v134d216 = hbusreq5_p & v134d215 | !hbusreq5_p & v134d1e8;
assign v1445f7c = hlock3 & v1445f6f | !hlock3 & v1445f7b;
assign v14457ff = hlock2 & v14457f6 | !hlock2 & v14457fe;
assign v1216214 = hgrant5_p & v121620f | !hgrant5_p & !v1216213;
assign v1445b21 = hbusreq2_p & v1445b1f | !hbusreq2_p & v1445b20;
assign v1216111 = hgrant1_p & v845542 | !hgrant1_p & v1216110;
assign v15168fa = hmaster0_p & v1668c3f | !hmaster0_p & v15168f9;
assign v12162c7 = hmaster0_p & v12160e2 | !hmaster0_p & v1216232;
assign a6538f = hbusreq0 & a6537b | !hbusreq0 & a6538e;
assign v134ce7c = decide_p & v134d3ce | !decide_p & v134ce6e;
assign v1668d72 = hgrant1_p & v1668d65 | !hgrant1_p & v1668d71;
assign v12aeb1b = hmaster1_p & v845542 | !hmaster1_p & v12aeb1a;
assign v16a141e = hgrant3_p & v16a13da | !hgrant3_p & v16a141d;
assign d301a0 = hmaster1_p & d3090c | !hmaster1_p & !d3019e;
assign v1668d4c = hgrant1_p & v1668d46 | !hgrant1_p & v1668d4b;
assign v144542e = hbusreq2_p & v144542d | !hbusreq2_p & v144541b;
assign v144538a = hbusreq2_p & v144537b | !hbusreq2_p & v1445389;
assign v1214bd4 = hmaster1_p & v1214bb5 | !hmaster1_p & v1214bcf;
assign v12aeb7c = hbusreq2_p & v12aeb73 | !hbusreq2_p & v12aeb7b;
assign v1284ca6 = hmaster2_p & v1284ca4 | !hmaster2_p & v1284ca5;
assign v1216213 = hmaster2_p & v1216212 | !hmaster2_p & v845542;
assign v121543e = hlock2_p & v121543a | !hlock2_p & v121543d;
assign v1405aaf = hmaster1_p & v1405aa3 | !hmaster1_p & v1405aae;
assign v12161af = hmaster1_p & v121618e | !hmaster1_p & v12161ae;
assign v134cd6c = hmaster1_p & v134d369 | !hmaster1_p & v134cd6b;
assign jx0 = v1405b69;
assign v15530f0 = hlock5 & v15530eb | !hlock5 & v15530ef;
assign v12161f8 = hmaster0_p & v1216038 | !hmaster0_p & v12161f7;
assign a65926 = hbusreq2_p & a65924 | !hbusreq2_p & a65925;
assign v121657b = hmaster1_p & v121657a | !hmaster1_p & v845542;
assign v1446273 = hmaster0_p & v144639c | !hmaster0_p & v144643d;
assign v12af3ac = hmaster1_p & v845542 | !hmaster1_p & v12af3ab;
assign v134ce7d = hready_p & v134d3e5 | !hready_p & v134ce7c;
assign d2fb00 = hbusreq1_p & d300f9 | !hbusreq1_p & d2faff;
assign d305e6 = hlock3_p & d305e5 | !hlock3_p & v84555e;
assign v16a1da4 = hbusreq2_p & v16a1da2 | !hbusreq2_p & v16a1da3;
assign v1215345 = hlock0_p & v1216a5a | !hlock0_p & v845542;
assign v1214c87 = hgrant5_p & v845542 | !hgrant5_p & v1214c52;
assign v1216303 = hmaster0_p & v1216300 | !hmaster0_p & v1216302;
assign a6568d = hbusreq2 & a65686 | !hbusreq2 & a6568b;
assign v15156f3 = hmaster1_p & v15156f2 | !hmaster1_p & v151566b;
assign d2fb04 = hgrant1_p & d2fb00 | !hgrant1_p & d2fb03;
assign d30258 = hmaster0_p & d30240 | !hmaster0_p & d30257;
assign v1216aaf = stateG2_p & v845542 | !stateG2_p & !v1446394;
assign v138a483 = hmaster0_p & v84555c | !hmaster0_p & v138a443;
assign v16a1bea = hgrant2_p & v845542 | !hgrant2_p & !v16a1be9;
assign v1216044 = hmaster1_p & v1216043 | !hmaster1_p & v1216041;
assign v12147ff = hbusreq2_p & v12147fe | !hbusreq2_p & v12164e7;
assign v144668a = hbusreq1 & v1446689 | !hbusreq1 & v14465c5;
assign v134d4b2 = hbusreq2_p & v134d4b0 | !hbusreq2_p & v134d4b1;
assign v121631b = hmaster0_p & v121631a | !hmaster0_p & v12162f3;
assign v15156fe = hbusreq2_p & v15156fd | !hbusreq2_p & v845542;
assign d2fb28 = hbusreq5_p & d3014b | !hbusreq5_p & !d2fb27;
assign v151573a = hbusreq5_p & v1515738 | !hbusreq5_p & v1515739;
assign v1405b54 = hbusreq2_p & v1405b44 | !hbusreq2_p & v1405b53;
assign v1215ca6 = hmaster2_p & v1215c94 | !hmaster2_p & v1215ca5;
assign v144579f = hmaster1_p & v144579e | !hmaster1_p & v1445e07;
assign v1284cf7 = hlock0_p & v1284c8f | !hlock0_p & v1284cf6;
assign v1405aa5 = hbusreq1_p & v1405aa4 | !hbusreq1_p & v1405a87;
assign v1446287 = hlock2 & v1446284 | !hlock2 & v1446286;
assign d30721 = hbusreq5_p & d30720 | !hbusreq5_p & v84554e;
assign v1445b19 = hmaster1_p & v1445afa | !hmaster1_p & v144591b;
assign d2f98b = hlock1_p & d2f98a | !hlock1_p & v84555a;
assign v1284d4a = hgrant4_p & v140583c | !hgrant4_p & v1284d49;
assign d301e1 = hgrant5_p & d301c3 | !hgrant5_p & !d301d8;
assign v138a395 = hmaster0_p & v138a394 | !hmaster0_p & v138a344;
assign v1215416 = hbusreq2_p & v1215415 | !hbusreq2_p & v1215411;
assign f2f3fd = hbusreq2_p & f2f3fa | !hbusreq2_p & f2f3fc;
assign d2fb70 = hbusreq1_p & d2fb6f | !hbusreq1_p & v84554a;
assign v1214c8e = hbusreq5_p & v1214c8c | !hbusreq5_p & v1214c8d;
assign v12162ee = hmaster2_p & v1216aad | !hmaster2_p & v12162ed;
assign v1446609 = hgrant1_p & v1446427 | !hgrant1_p & v1446608;
assign v134cd70 = hbusreq0 & v134cd6f | !hbusreq0 & v134d274;
assign v121604e = hlock5_p & v121604d | !hlock5_p & v16a2243;
assign v138a2f9 = hlock5_p & v151570f | !hlock5_p & v845570;
assign v12161aa = hlock5_p & v1216194 | !hlock5_p & v12161a9;
assign d2fb5b = hmaster0_p & d2fb5a | !hmaster0_p & d2fb51;
assign d301a9 = hgrant2_p & d301a6 | !hgrant2_p & d301a0;
assign v134cd64 = hlock1 & v134d385 | !hlock1 & v134cd63;
assign v1445784 = hmaster0_p & v1445776 | !hmaster0_p & v1445e0a;
assign v1216271 = hbusreq2_p & v121626e | !hbusreq2_p & v1216270;
assign v1215708 = hmaster1_p & v1215707 | !hmaster1_p & v1215b88;
assign v15155f9 = hlock0_p & v1668c1c | !hlock0_p & v15155f8;
assign v1446153 = hmaster1_p & v1446136 | !hmaster1_p & v1445ffc;
assign d2fd0a = hlock2_p & v845542 | !hlock2_p & !d2fd09;
assign v1214d34 = hgrant3_p & v1214c41 | !hgrant3_p & v1214d33;
assign v14459c2 = hgrant4_p & v14458db | !hgrant4_p & v14459c1;
assign v10d40a8 = hbusreq2_p & v10d40a6 | !hbusreq2_p & v10d40a7;
assign v144587f = hbusreq5_p & v144587a | !hbusreq5_p & v144587e;
assign v1445f5f = hbusreq2 & v1445f59 | !hbusreq2 & v1445f5e;
assign a65467 = hburst1 & v156645f | !hburst1 & a65466;
assign v1668e0b = decide_p & v1668e08 | !decide_p & v845542;
assign d300bd = hgrant4_p & v845542 | !hgrant4_p & d300bc;
assign v134d274 = hmaster2_p & v845542 | !hmaster2_p & v134d273;
assign v140586c = hbusreq4_p & v140586b | !hbusreq4_p & v14463b1;
assign v140589a = locked_p & v1405899 | !locked_p & v1405844;
assign d301af = hlock2_p & d301ae | !hlock2_p & d301a0;
assign v1214ce7 = hmaster1_p & v1214ce6 | !hmaster1_p & v1214c39;
assign v134cd77 = hlock2 & v134d3b5 | !hlock2 & v134cd6d;
assign d306cc = hlock1_p & v845542 | !hlock1_p & a66295;
assign a6585d = hbusreq4_p & a6585c | !hbusreq4_p & v845542;
assign v1445a43 = hlock0 & v1445a3f | !hlock0 & v1445a42;
assign v12153ba = hbusreq5_p & v12153b8 | !hbusreq5_p & v12153b9;
assign v12ad4eb = hmaster2_p & v12ad4e4 | !hmaster2_p & v845542;
assign v1668db1 = hbusreq3 & v1668db0 | !hbusreq3 & v845542;
assign d30206 = hgrant1_p & d30205 | !hgrant1_p & d307c9;
assign d307b6 = hbusreq1_p & d307b5 | !hbusreq1_p & v845542;
assign v16a206b = hgrant0_p & v845542 | !hgrant0_p & v16a206a;
assign v15156d9 = hbusreq5_p & v15156d7 | !hbusreq5_p & v15156d8;
assign d307f0 = hgrant5_p & d30705 | !hgrant5_p & d307ee;
assign d307e2 = hbusreq1 & d307e1 | !hbusreq1 & v845542;
assign v16695bb = hlock3_p & v16695ba | !hlock3_p & v845542;
assign v1445887 = hlock1 & v144586f | !hlock1 & v1445882;
assign v138a33c = hbusreq4_p & a658e0 | !hbusreq4_p & a65472;
assign v12ad001 = hbusreq4_p & v12ad5c1 | !hbusreq4_p & v12ad000;
assign a658ee = hmaster2_p & a658b0 | !hmaster2_p & !a658be;
assign v1215727 = hlock4_p & v1215726 | !hlock4_p & v845572;
assign d307c9 = hgrant4_p & d307c7 | !hgrant4_p & d307c8;
assign v1446611 = hgrant5_p & v144642a | !hgrant5_p & v1446610;
assign d3081b = hlock5_p & d30819 | !hlock5_p & d3081a;
assign v1446556 = hbusreq2_p & v14464a3 | !hbusreq2_p & v1446555;
assign d80787 = hbusreq2_p & d80785 | !hbusreq2_p & d80786;
assign v12ad625 = hbusreq2 & v12ad621 | !hbusreq2 & v12ad624;
assign v1215d70 = hmaster2_p & v1216588 | !hmaster2_p & v12166d2;
assign f2f39d = hmaster0_p & f2f39c | !hmaster0_p & f2f385;
assign v1216292 = hmaster1_p & v1216291 | !hmaster1_p & v121619c;
assign v12160f2 = hbusreq4 & v845570 | !hbusreq4 & v845542;
assign v12153b6 = hmaster0_p & v1215baf | !hmaster0_p & v12153b5;
assign v16a1dac = hbusreq3 & v16a1da8 | !hbusreq3 & !v16a1dab;
assign v1445be6 = hbusreq2_p & v1445be4 | !hbusreq2_p & v1445be5;
assign v1445e79 = hmaster2_p & v144639c | !hmaster2_p & v1445df5;
assign v16a1e07 = hgrant2_p & v845542 | !hgrant2_p & v16a1e06;
assign d30757 = hlock2_p & d30755 | !hlock2_p & d30756;
assign d80786 = hgrant2_p & v845542 | !hgrant2_p & d80784;
assign v1445f9c = hmaster2_p & v1445f93 | !hmaster2_p & v1445f9b;
assign v1515846 = hgrant5_p & v845542 | !hgrant5_p & !v1515837;
assign v1214ff6 = hbusreq1_p & v1214fea | !hbusreq1_p & v1214ff5;
assign a65471 = hbusreq5_p & a6546f | !hbusreq5_p & !a65470;
assign v14058ba = hlock5_p & v14058b8 | !hlock5_p & v14058b9;
assign v16a13c6 = hmaster1_p & v16a13c5 | !hmaster1_p & v16a2672;
assign v1445894 = hmaster2_p & v1445893 | !hmaster2_p & v14463bb;
assign v1446635 = hmaster2_p & v144639c | !hmaster2_p & v1446634;
assign v121609c = hlock2_p & v1216098 | !hlock2_p & v121609b;
assign v12161fa = hmaster2_p & v12161d0 | !hmaster2_p & v12161da;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hbusreq2_p = 0;
  hlock2_p = 0;
  hbusreq3_p = 0;
  hlock3_p = 0;
  hbusreq4_p = 0;
  hlock4_p = 0;
  hbusreq5_p = 0;
  hlock5_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmaster1_p = 0;
  hmaster2_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  hgrant2_p = 0;
  hgrant3_p = 0;
  hgrant4_p = 0;
  hgrant5_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  stateG10_2_p = 0;
  stateG10_3_p = 0;
  stateG10_4_p = 0;
  stateG10_5_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hbusreq2_p = hbusreq2;
  hlock2_p = hlock2;
  hbusreq3_p = hbusreq3;
  hlock3_p = hlock3;
  hbusreq4_p = hbusreq4;
  hlock4_p = hlock4;
  hbusreq5_p = hbusreq5;
  hlock5_p = hlock5;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmaster1_p = hmaster1;
  hmaster2_p = hmaster2;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  hgrant2_p = hgrant2;
  hgrant3_p = hgrant3;
  hgrant4_p = hgrant4;
  hgrant5_p = hgrant5;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  stateG10_2_p = stateG10_2;
  stateG10_3_p = stateG10_3;
  stateG10_4_p = stateG10_4;
  stateG10_5_p = stateG10_5;
  jx0_p = jx0;
  jx1_p = jx1;
  jx2_p = jx2;
    end
endmodule

