module main(clock, StoB_REQ0_n, StoB_REQ1_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, jx0_n, jx1_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844fa7;
  wire v85d449;
  wire v84ff94;
  wire v85d456;
  wire v844f9b;
  wire v85a6f2;
  wire v85a9de;
  wire v85d584;
  wire v85d507;
  wire v85a87f;
  wire v85b457;
  wire v858ca9;
  wire v858cc1;
  wire v859ee0;
  wire v844f99;
  wire v84f639;
  wire v844fab;
  wire v85a33b;
  wire v84f61b;
  wire v85a854;
  wire v85d4b0;
  wire v85d44e;
  wire v85d4c8;
  wire v85d445;
  wire v85d444;
  wire v85add3;
  wire v85d42d;
  wire v85d4f7;
  wire v85d463;
  wire v85d440;
  wire v85d43d;
  wire v85a260;
  wire v85d45c;
  wire v844faf;
  wire v844f9f;
  wire v85a68e;
  wire v85d4cf;
  wire v85d4d0;
  wire v85a8c6;
  wire v85d4ff;
  wire v85d44c;
  wire v85d45d;
  wire v85d4ed;
  wire v85d485;
  wire v85d4c6;
  wire v84f5b2;
  wire v85d593;
  wire v85a6f5;
  wire v85a9ac;
  wire v84f724;
  wire v85a797;
  wire v85a82c;
  wire v85d490;
  wire v85a78d;
  wire v85d479;
  wire v85a8fa;
  wire v84f6ed;
  wire v85a70b;
  wire v85d610;
  wire v84f6cb;
  wire v858cc2;
  wire v85a6c5;
  wire v85d42a;
  wire v85d4c7;
  wire v85a770;
  wire v85a815;
  wire v84edb2;
  wire v85d4d7;
  wire v85a646;
  wire v85a705;
  wire v85a757;
  wire v84ed3f;
  wire v85d466;
  wire v859ec3;
  wire v85a245;
  wire v85a7d9;
  wire v85a914;
  wire v85a331;
  wire v85a235;
  wire v85d4d5;
  wire v859ebe;
  wire v85d43c;
  wire v84ecfb;
  wire v85a8c1;
  wire v85a776;
  wire v85a96d;
  wire v84faa7;
  wire v85046f;
  wire v85d4cd;
  wire v85d457;
  wire v85d514;
  wire v85a941;
  wire v85a833;
  wire v85d534;
  wire v85b465;
  wire v844f95;
  wire v844f9d;
  wire v8544ec;
  wire v85b456;
  wire v85a8d5;
  wire v85d4a7;
  wire v85bdde;
  wire v85d4fe;
  wire v85d45e;
  wire v85d429;
  wire v85d44b;
  wire v85a894;
  wire v85a779;
  wire v85d47a;
  wire v85d4af;
  wire v85cfa5;
  wire v85d566;
  wire v85d508;
  wire v85d505;
  wire v85bd9c;
  wire v85d5a2;
  wire v85a9aa;
  wire v85d426;
  wire v85ae01;
  wire v84f197;
  wire v85a975;
  wire v85d439;
  wire v85bf72;
  wire v85a6bc;
  wire v85a32f;
  wire v85adcc;
  wire v85d486;
  wire v84fe9e;
  wire v85a259;
  wire v85a718;
  wire v844f97;
  wire v85d4d4;
  wire v85d4ee;
  wire v85d46e;
  wire v85d48f;
  wire v85d434;
  wire v85a792;
  wire v85d49b;
  wire v850262;
  wire v85a2fd;
  wire v85cfa7;
  wire v85ae0d;
  wire v84f976;
  wire v85d452;
  wire v84f975;
  wire v85d5b7;
  wire v85c725;
  wire v85042c;
  wire v844fb1;
  wire v85aa1a;
  wire v85ae0f;
  wire v85bf68;
  wire v85ade5;
  wire v85d4ef;
  wire v85d47b;
  wire v85a820;
  wire v85a924;
  wire v85a30d;
  wire v85d586;
  wire v85d58a;
  wire v855693;
  wire v85d4ea;
  wire v84d668;
  wire v85a737;
  wire v85d4fd;
  wire v85d601;
  wire v85a9b1;
  wire v85a298;
  wire v85b414;
  wire v84ffcf;
  wire v85a8ec;
  wire v85adc8;
  wire v85d467;
  wire v85d503;
  wire v85cfa6;
  wire v85d482;
  wire v85bdd5;
  wire v85d4c4;
  wire v85aa06;
  wire v8504a5;
  wire v84f229;
  wire v85d425;
  wire v85569b;
  wire v85adee;
  wire v85d464;
  wire v85a9eb;
  wire v858c4d;
  wire v85a7be;
  wire v85d4ce;
  wire v85a653;
  wire v858c78;
  wire v85a7c2;
  wire v85a8cd;
  wire v85d450;
  wire v85d460;
  wire v85a256;
  wire v85d59b;
  wire v85a808;
  wire v85a8f2;
  wire v85d496;
  wire v85bde6;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  wire SLC0_n;
  wire ENQ_n;

assign v85cfa6 = DEQ_p & v844f91 | !DEQ_p & v85d503;
assign BtoS_ACK0_n = v85bf72;
assign v85042c = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v84f976;
assign v85a331 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85a914;
assign v85d426 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v85a9aa;
assign v85d429 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85d45e;
assign v85a6f5 = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v85d593;
assign v85ade5 = BtoR_REQ1_p & v85aa1a | !BtoR_REQ1_p & v844fb1;
assign v85bdde = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v85d4a7;
assign DEQ_n = !v859ee0;
assign v85a2fd = BtoS_ACK0_p & v85d434 | !BtoS_ACK0_p & !v850262;
assign v85a87f = BtoS_ACK1_p & v85d456 | !BtoS_ACK1_p & v85d584;
assign v84f976 = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & !v844f97;
assign v84f639 = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v844f91;
assign v85d586 = RtoB_ACK0_p & v844fb1 | !RtoB_ACK0_p & v85ae0f;
assign v859ec3 = BtoS_ACK0_p & v84edb2 | !BtoS_ACK0_p & v85d466;
assign BtoR_REQ1_n = !v85b465;
assign v85a33b = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v844fab;
assign v85a705 = StoB_REQ1_p & v85a770 | !StoB_REQ1_p & v85a646;
assign v85a9de = BtoR_REQ0_p & v85a6f2 | !BtoR_REQ0_p & !v84ff94;
assign v85a833 = BtoS_ACK0_p & v85d457 | !BtoS_ACK0_p & v85a941;
assign v85a9aa = BtoR_REQ0_p & v85d566 | !BtoR_REQ0_p & v85d5a2;
assign v84ff94 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v85d449;
assign v85d425 = BtoS_ACK1_p & v85d467 | !BtoS_ACK1_p & v84f229;
assign v844fb1 = stateG12_p & v844f91 | !stateG12_p & !v844f91;
assign v858cc1 = BtoS_ACK0_p & v85d584 | !BtoS_ACK0_p & v85b457;
assign v85d4ce = stateG7_1_p & v844fb1 | !stateG7_1_p & v844f91;
assign v84f6cb = jx1_p & v85a82c | !jx1_p & v85d610;
assign v85adc8 = BtoR_REQ0_p & v85bf68 | !BtoR_REQ0_p & v85a8ec;
assign v844f9d = FULL_p & v844f91 | !FULL_p & !v844f91;
assign v85a235 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v85a331;
assign v85bd9c = RtoB_ACK1_p & v85d508 | !RtoB_ACK1_p & v85d505;
assign v85d4ef = RtoB_ACK1_p & v85ade5 | !RtoB_ACK1_p & v85aa1a;
assign v84faa7 = BtoS_ACK1_p & v85a776 | !BtoS_ACK1_p & v85a96d;
assign v85d440 = BtoS_ACK0_p & v85d4c8 | !BtoS_ACK0_p & v85d463;
assign v84f197 = StoB_REQ0_p & v85ae01 | !StoB_REQ0_p & v844f91;
assign v85b456 = RtoB_ACK0_p & v8544ec | !RtoB_ACK0_p & !v844f91;
assign v84ed3f = BtoS_ACK1_p & v85d4c7 | !BtoS_ACK1_p & v85a815;
assign v85bf68 = RtoB_ACK0_p & v85aa1a | !RtoB_ACK0_p & v85ae0f;
assign v85a894 = BtoS_ACK0_p & v844f95 | !BtoS_ACK0_p & !v85d44b;
assign v85d4f7 = BtoS_ACK1_p & v84f639 | !BtoS_ACK1_p & v85d44e;
assign v85a32f = BtoR_REQ1_p & v844faf | !BtoR_REQ1_p & v844f91;
assign v85d4c4 = BtoR_REQ1_p & v85cfa6 | !BtoR_REQ1_p & v844fb1;
assign v85d4a7 = RtoB_ACK1_p & v85a8d5 | !RtoB_ACK1_p & !v844f91;
assign v84ffcf = RtoB_ACK1_p & v85ade5 | !RtoB_ACK1_p & v85b414;
assign v85d44c = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85d4ff;
assign v85a9b1 = StoB_REQ1_p & v85d58a | !StoB_REQ1_p & v85d601;
assign v85d59b = BtoS_ACK1_p & v85a7be | !BtoS_ACK1_p & v85a256;
assign v85a7d9 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v85a245;
assign v85a8c6 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v85d4d0;
assign v85d4c8 = StoB_REQ0_p & v84f639 | !StoB_REQ0_p & v85d44e;
assign v85a298 = StoB_REQ0_p & v85a30d | !StoB_REQ0_p & v85a9b1;
assign v85d4d5 = StoB_REQ1_p & v85a770 | !StoB_REQ1_p & v85a235;
assign v85aa06 = RtoB_ACK1_p & v85d4c4 | !RtoB_ACK1_p & v85cfa6;
assign v85d505 = BtoR_REQ1_p & v8544ec | !BtoR_REQ1_p & !v844f91;
assign v85d47b = RtoB_ACK0_p & v844fb1 | !RtoB_ACK0_p & v85d4ef;
assign v85d479 = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v85a78d;
assign v85a854 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v84f61b;
assign v85d45d = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v85d44c;
assign v85d4fd = RtoB_ACK0_p & v844fb1 | !RtoB_ACK0_p & v85a737;
assign v85a8cd = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v85a7c2;
assign v85a776 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v85a8c1;
assign v858c4d = RtoB_ACK0_p & v844fb1 | !RtoB_ACK0_p & v85a9eb;
assign v844fa7 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v844f91;
assign v84f6ed = BtoS_ACK1_p & v85a8fa | !BtoS_ACK1_p & v85d4b0;
assign v84f229 = BtoR_REQ0_p & v85bdd5 | !BtoR_REQ0_p & v8504a5;
assign v85d42a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85a6c5;
assign v85d4ee = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & v85d4d4;
assign v844f91 = 1;
assign v85ae01 = BtoS_ACK1_p & v85d426 | !BtoS_ACK1_p & !v85a9aa;
assign v85d4cd = BtoS_ACK0_p & v85d4d5 | !BtoS_ACK0_p & v85046f;
assign v85d4ed = StoB_REQ1_p & v85d45c | !StoB_REQ1_p & v85d45d;
assign v85d5b7 = jx1_p & v844f91 | !jx1_p & !v84f975;
assign v85d456 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v84ff94;
assign v84f5b2 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v85d4c6;
assign v85d464 = BtoR_REQ1_p & v85aa1a | !BtoR_REQ1_p & v85adee;
assign v85a792 = BtoS_ACK1_p & v844f97 | !BtoS_ACK1_p & !v844f91;
assign v85b414 = BtoR_REQ1_p & v85aa1a | !BtoR_REQ1_p & v844faf;
assign v85aa1a = DEQ_p & v844f91 | !DEQ_p & v844fb1;
assign v85a8d5 = BtoR_REQ1_p & v8544ec | !BtoR_REQ1_p & !v844f9d;
assign v85a256 = StoB_REQ1_p & v84f229 | !StoB_REQ1_p & v85d460;
assign v85d58a = BtoR_REQ0_p & v85d586 | !BtoR_REQ0_p & v844fb1;
assign v85d508 = BtoR_REQ1_p & v8544ec | !BtoR_REQ1_p & v844f91;
assign v85a770 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v85a78d;
assign v85bf72 = jx0_p & v85a894 | !jx0_p & v85d439;
assign v85a914 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v85a7d9;
assign v85d486 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85adcc;
assign v85d5a2 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85bd9c;
assign v85a96d = StoB_REQ1_p & v85a770 | !StoB_REQ1_p & v85a776;
assign v85a7be = BtoR_REQ0_p & v85aa1a | !BtoR_REQ0_p & v858c4d;
assign v85d434 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v85d48f;
assign v85d460 = BtoR_REQ0_p & v85d4ce | !BtoR_REQ0_p & v85d450;
assign v84f724 = BtoS_ACK1_p & v85a6f5 | !BtoS_ACK1_p & v85a9ac;
assign BtoS_ACK1_n = !v85cfa7;
assign v85d496 = jx1_p & v85a8f2 | !jx1_p & !v844f91;
assign v855693 = stateG12_p & v844f9f | !stateG12_p & v844f91;
assign v85b465 = jx0_p & v859ec3 | !jx0_p & v85d534;
assign v85d534 = jx1_p & v85d4cd | !jx1_p & v85a833;
assign v85a646 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v85d4d7;
assign v85add3 = StoB_REQ1_p & v85d444 | !StoB_REQ1_p & v84f639;
assign v844faf = DEQ_p & v844f91 | !DEQ_p & !v844f91;
assign v85a6c5 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844fa7;
assign v85d43d = RtoB_ACK1_p & v844fa7 | !RtoB_ACK1_p & v85a33b;
assign v85d45c = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v85a260;
assign v85d445 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85a33b;
assign v85d4c6 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v85d485;
assign v85d482 = RtoB_ACK1_p & v844fb1 | !RtoB_ACK1_p & v85cfa6;
assign v85d514 = BtoS_ACK1_p & v85d4c7 | !BtoS_ACK1_p & v85d457;
assign v85d507 = StoB_REQ0_p & v85d456 | !StoB_REQ0_p & v85d584;
assign v844f9b = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844f91;
assign v85d4ea = DEQ_p & v844fb1 | !DEQ_p & !v855693;
assign v85d439 = jx1_p & v85d4af | !jx1_p & v85a975;
assign v85a9ac = StoB_REQ1_p & v85d45c | !StoB_REQ1_p & v85a6f5;
assign v85d4cf = ENQ_p & v844faf | !ENQ_p & v85a68e;
assign v85d450 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85a8cd;
assign v858ca9 = BtoS_ACK0_p & v85d507 | !BtoS_ACK0_p & v85b457;
assign v85d444 = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v85d445;
assign v85a820 = BtoR_REQ0_p & v85bf68 | !BtoR_REQ0_p & v85d47b;
assign v85d4fe = BtoR_REQ0_p & v85b456 | !BtoR_REQ0_p & !v85bdde;
assign v85bde6 = jx0_p & v85042c | !jx0_p & !v85d496;
assign v85a757 = BtoS_ACK1_p & v85a646 | !BtoS_ACK1_p & v85a705;
assign v85d485 = stateG7_1_p & v85a68e | !stateG7_1_p & v844f91;
assign v858cc2 = jx0_p & v85d440 | !jx0_p & v84f6cb;
assign v85a259 = StoB_REQ1_p & v84fe9e | !StoB_REQ1_p & !v844f91;
assign v85d566 = RtoB_ACK0_p & v8544ec | !RtoB_ACK0_p & v85cfa5;
assign v859ebe = stateG7_1_p & v844f91 | !stateG7_1_p & v85a68e;
assign v85d4d7 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v85a6c5;
assign v8504a5 = RtoB_ACK0_p & v844fb1 | !RtoB_ACK0_p & v85aa06;
assign v85a6bc = RtoB_ACK0_p & v844faf | !RtoB_ACK0_p & v85cfa5;
assign v84f61b = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v85a33b;
assign v85a68e = DEQ_p & v844f91 | !DEQ_p & v844f9f;
assign v85a70b = StoB_REQ0_p & v84f6ed | !StoB_REQ0_p & v84f639;
assign v85a30d = StoB_REQ1_p & v85a820 | !StoB_REQ1_p & v85a924;
assign v85d46e = BtoS_ACK0_p & v85a718 | !BtoS_ACK0_p & !v85d4ee;
assign v85569b = DEQ_p & v844fb1 | !DEQ_p & !v844f91;
assign v85a808 = StoB_REQ0_p & v85d425 | !StoB_REQ0_p & v85d59b;
assign v85c725 = jx0_p & v85d452 | !jx0_p & v85d5b7;
assign v85a260 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85d43d;
assign jx1_n = !v85bde6;
assign BtoR_REQ0_n = !v858cc2;
assign v85a815 = StoB_REQ1_p & v85a770 | !StoB_REQ1_p & v85d4c7;
assign v85ae0f = RtoB_ACK1_p & v844fb1 | !RtoB_ACK1_p & v85aa1a;
assign v85d601 = BtoR_REQ0_p & v844fb1 | !BtoR_REQ0_p & v85d4fd;
assign v85a6f2 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f9b;
assign v85d490 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v85a33b;
assign v85d44e = StoB_REQ1_p & v85d4b0 | !StoB_REQ1_p & v84f639;
assign v85d467 = StoB_REQ1_p & v85adc8 | !StoB_REQ1_p & v85d58a;
assign v85a941 = StoB_REQ0_p & v85a770 | !StoB_REQ0_p & v85d514;
assign v85ae0d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f97;
assign v85d47a = StoB_REQ0_p & v85a779 | !StoB_REQ0_p & v844f91;
assign v85bdd5 = RtoB_ACK0_p & v85cfa6 | !RtoB_ACK0_p & v85d482;
assign v85cfa7 = jx0_p & v85d46e | !jx0_p & v85a2fd;
assign v85d42d = BtoS_ACK1_p & v84f639 | !BtoS_ACK1_p & v85add3;
assign v844f99 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v85d610 = BtoS_ACK0_p & v84f639 | !BtoS_ACK0_p & v85a70b;
assign v85d584 = StoB_REQ1_p & v85a9de | !StoB_REQ1_p & v85d456;
assign v85d4b0 = BtoR_REQ0_p & v844f99 | !BtoR_REQ0_p & v85a854;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v85a8f2 = BtoS_ACK0_p & v85a298 | !BtoS_ACK0_p & v85a808;
assign v85a8c1 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v84ecfb;
assign v85d452 = BtoS_ACK0_p & v85ae0d | !BtoS_ACK0_p & v84f976;
assign v844f9f = EMPTY_p & v844f91 | !EMPTY_p & !v844f91;
assign v85b457 = StoB_REQ0_p & v85a9de | !StoB_REQ0_p & v85a87f;
assign v85d457 = StoB_REQ1_p & v85a646 | !StoB_REQ1_p & v85d4c7;
assign v85d4d4 = StoB_REQ1_p & v85a9aa | !StoB_REQ1_p & !v844f91;
assign v85a7c2 = BtoR_REQ1_p & v85a653 | !BtoR_REQ1_p & v858c78;
assign v84f975 = BtoS_ACK0_p & v844f95 | !BtoS_ACK0_p & !v844f95;
assign v85a82c = BtoS_ACK0_p & v85d4ed | !BtoS_ACK0_p & v85a797;
assign v85d466 = StoB_REQ0_p & v85a757 | !StoB_REQ0_p & v84ed3f;
assign v85d45e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v85d4fe;
assign v85a78d = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v85d490;
assign v85d4af = BtoS_ACK0_p & v844f95 | !BtoS_ACK0_p & !v85d47a;
assign v85a797 = StoB_REQ0_p & v85d45c | !StoB_REQ0_p & v84f724;
assign v85a653 = stateG7_1_p & v844f91 | !stateG7_1_p & v844fb1;
assign v85a975 = BtoS_ACK0_p & v844f95 | !BtoS_ACK0_p & !v84f197;
assign v85a718 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v85a259;
assign v859ee0 = jx0_p & v858ca9 | !jx0_p & v858cc1;
assign v85a245 = stateG7_1_p & v844f91 | !stateG7_1_p & v85d4cf;
assign v85d44b = StoB_REQ0_p & v85d429 | !StoB_REQ0_p & v844f91;
assign v84edb2 = StoB_REQ0_p & v85d4c7 | !StoB_REQ0_p & v85a815;
assign v85adcc = RtoB_ACK1_p & v85a32f | !RtoB_ACK1_p & v85d505;
assign v85adee = ENQ_p & v85569b | !ENQ_p & v85d4ea;
assign v84fe9e = BtoR_REQ0_p & v85a6bc | !BtoR_REQ0_p & v85d486;
assign v85d48f = StoB_REQ1_p & v85d4fe | !StoB_REQ1_p & !v844f91;
assign v85046f = StoB_REQ0_p & v85a770 | !StoB_REQ0_p & v84faa7;
assign v844fab = stateG7_1_p & v844f91 | !stateG7_1_p & !v844f91;
assign v85d503 = stateG12_p & v844f91 | !stateG12_p & v844f9d;
assign v85d449 = RtoB_ACK1_p & v844fa7 | !RtoB_ACK1_p & v844f91;
assign v84d668 = BtoR_REQ1_p & v844fb1 | !BtoR_REQ1_p & v85d4ea;
assign v850262 = StoB_REQ0_p & v85a792 | !StoB_REQ0_p & v85d49b;
assign v85d49b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85d48f;
assign v85a8fa = StoB_REQ1_p & v85d479 | !StoB_REQ1_p & v85d4b0;
assign v85d4ff = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v85a8c6;
assign v85cfa5 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8544ec;
assign v85d43c = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v859ebe;
assign v85a9eb = RtoB_ACK1_p & v85ade5 | !RtoB_ACK1_p & v85d464;
assign v85a924 = BtoR_REQ0_p & v85aa1a | !BtoR_REQ0_p & v85d47b;
assign v85d593 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v84f5b2;
assign v8544ec = DEQ_p & v844f91 | !DEQ_p & !v844f9d;
assign v85d463 = StoB_REQ0_p & v85d42d | !StoB_REQ0_p & v85d4f7;
assign v85a779 = BtoS_ACK1_p & v85d45e | !BtoS_ACK1_p & !v85d4fe;
assign v84ecfb = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v85d43c;
assign v85a737 = RtoB_ACK1_p & v844fb1 | !RtoB_ACK1_p & v84d668;
assign v85a8ec = RtoB_ACK0_p & v844fb1 | !RtoB_ACK0_p & v84ffcf;
assign jx0_n = !v85c725;
assign v858c78 = DEQ_p & v844f91 | !DEQ_p & !v855693;
assign v85d4d0 = stateG7_1_p & v85d4cf | !stateG7_1_p & v844f91;
assign v85d4c7 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v85d42a;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign SLC0_n = (!BtoS_ACK0_n & ((StoB_REQ1_n & ((BtoS_ACK1_n)))));
assign ENQ_n = (BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((SLC0_n)));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  jx0_p = 0;
  jx1_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
