module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, StoB_REQ4_n, StoB_REQ5_n, StoB_REQ6_n, StoB_REQ7_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoS_ACK4_n, BtoS_ACK5_n, BtoS_ACK6_n, BtoS_ACK7_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, SLC2_n, jx0_n, jx1_n, jx2_n, jx3_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844fb9;
  wire v8af02f;
  wire v844fa1;
  wire v8af916;
  wire v8b25a2;
  wire v912554;
  wire v8ae9c2;
  wire v8c66bb;
  wire v912724;
  wire v873367;
  wire v91180b;
  wire v844f9f;
  wire v8aef02;
  wire v8b33a8;
  wire v911787;
  wire v8afe4c;
  wire v8dd6a6;
  wire v8ae4e9;
  wire v91129a;
  wire v8b06bb;
  wire v8b04d6;
  wire v8ae487;
  wire v8c0457;
  wire v8aeed6;
  wire v912312;
  wire v8af9cf;
  wire v8aeecd;
  wire v8b76f4;
  wire v8b4c61;
  wire v9125e2;
  wire v8c4cc9;
  wire v8b11c5;
  wire v911218;
  wire v844f9d;
  wire v8ae516;
  wire v8b07c0;
  wire v8b0a55;
  wire v8b2019;
  wire v8b0cbb;
  wire v8b6d87;
  wire v8b0eab;
  wire v8b267f;
  wire v8aed8c;
  wire v91159f;
  wire v9116c2;
  wire v8afcd6;
  wire v8e9852;
  wire v8b3227;
  wire v844f9b;
  wire v8b034f;
  wire v91244d;
  wire v8b03cf;
  wire v8b10cf;
  wire v9114dc;
  wire v890bdc;
  wire v9125cc;
  wire v8b208f;
  wire v8afe2c;
  wire v9124ad;
  wire v8af564;
  wire v844f99;
  wire v8b7804;
  wire v912518;
  wire v9124fd;
  wire v8c0b90;
  wire v8b27a6;
  wire v887bda;
  wire v8ae0b9;
  wire v8c39e2;
  wire v867e4e;
  wire v911914;
  wire v911be0;
  wire v8af5ee;
  wire v844f97;
  wire v8c5845;
  wire v91257d;
  wire v9112ad;
  wire v9125eb;
  wire v911fe4;
  wire v9124c0;
  wire v9114e5;
  wire v8b2197;
  wire v8b3d1f;
  wire v912644;
  wire v8b336e;
  wire v8af68d;
  wire v911610;
  wire v91157d;
  wire v88c831;
  wire v91272c;
  wire v85f776;
  wire v9125e5;
  wire v8c53cf;
  wire v8af753;
  wire v8f958b;
  wire v8b0086;
  wire v8b21eb;
  wire v885339;
  wire v912561;
  wire v8c704b;
  wire v91263f;
  wire v911053;
  wire v8816a0;
  wire v8c702a;
  wire v8b2aa2;
  wire v8b52fa;
  wire v911289;
  wire v8cc108;
  wire v8c3d7b;
  wire v8b0ebf;
  wire v8b2f92;
  wire v9110fc;
  wire v911fd5;
  wire v8b0fe0;
  wire v911a56;
  wire v8909b7;
  wire v8af03f;
  wire v91127a;
  wire v8afc92;
  wire v8b3013;
  wire v8b09ce;
  wire v8af334;
  wire v912651;
  wire v912769;
  wire v9124bc;
  wire v8b1e91;
  wire v8714a5;
  wire v8c0508;
  wire v8afe22;
  wire v91272f;
  wire v91239a;
  wire v8b029e;
  wire v8b2815;
  wire v85e7ac;
  wire v8af748;
  wire v91250a;
  wire v8ae7a9;
  wire v911b4f;
  wire v912650;
  wire v8b2f95;
  wire v9124c9;
  wire v912424;
  wire v91177a;
  wire v8c57ef;
  wire v911539;
  wire v890930;
  wire v9110fb;
  wire v8d6cda;
  wire v8b246f;
  wire v8b1d12;
  wire v8bb768;
  wire v910ca3;
  wire v911692;
  wire v9123da;
  wire v912186;
  wire v8ae562;
  wire v8b085b;
  wire v8fed43;
  wire v8b2f8c;
  wire v9125e0;
  wire v8b1ff0;
  wire v894072;
  wire v8b2d81;
  wire v89409b;
  wire v912649;
  wire v911c45;
  wire v912430;
  wire v89288a;
  wire v892501;
  wire v8c65f8;
  wire v8fed90;
  wire v8af7b2;
  wire v8ae169;
  wire v9124e9;
  wire v9123a2;
  wire v8b2073;
  wire v9124be;
  wire v869876;
  wire v9125b2;
  wire v912648;
  wire v8b0062;
  wire v8b2590;
  wire v8b2ee4;
  wire v87cf4c;
  wire v9125ea;
  wire v8aeb91;
  wire v911d4b;
  wire v8af049;
  wire v91185f;
  wire v8b2920;
  wire v8b2e22;
  wire v910884;
  wire v91253b;
  wire v911c9a;
  wire v8aef67;
  wire v8af066;
  wire v911411;
  wire v911a59;
  wire v912578;
  wire v9110bd;
  wire v8b0b83;
  wire v8803b6;
  wire v912569;
  wire v8b22c1;
  wire v912746;
  wire v8b77ef;
  wire v912481;
  wire v9123e9;
  wire v911d50;
  wire v8b2e7b;
  wire v8b2639;
  wire v911eb1;
  wire v8c6e13;
  wire v844fa7;
  wire v887acc;
  wire v844fa5;
  wire v8b039c;
  wire v8b0339;
  wire v856df0;
  wire v8af65e;
  wire v890b14;
  wire v87cf6f;
  wire v8a8ba5;
  wire v844fa3;
  wire v8ae4b3;
  wire v8ae6f0;
  wire v8c3fe8;
  wire v8f956e;
  wire v8b263d;
  wire v8b52f8;
  wire v890ae8;
  wire v87d270;
  wire v8c3def;
  wire v8b0774;
  wire v8afbd6;
  wire v8ae6e0;
  wire v890a25;
  wire v8b0485;
  wire v8ae6f2;
  wire v8b1166;
  wire v8aec57;
  wire v85ed5d;
  wire v911917;
  wire v9124de;
  wire v8b2657;
  wire v8c23d8;
  wire v911fd9;
  wire v912623;
  wire v8afaa7;
  wire v912777;
  wire v86f676;
  wire v8afaed;
  wire v8af372;
  wire v8c48a1;
  wire v9114f1;
  wire v8b1fd2;
  wire v912617;
  wire v8b2bee;
  wire v912456;
  wire v910db7;
  wire v912581;
  wire v910e12;
  wire v8b32c2;
  wire v8b0764;
  wire v89085d;
  wire v8cc153;
  wire v8940a8;
  wire v8af095;
  wire v8b77fb;
  wire v8c3b67;
  wire v912682;
  wire v892ea3;
  wire v9126fc;
  wire v8b13b1;
  wire v8b1276;
  wire v8b032e;
  wire v8dd691;
  wire v8ae0da;
  wire v911174;
  wire v8ae104;
  wire v882eb7;
  wire v8af7c1;
  wire v8fed36;
  wire v91259e;
  wire v8b4ffd;
  wire v869205;
  wire v8b1d6c;
  wire v9117c1;
  wire v8b1fc9;
  wire v8dd654;
  wire v8af92f;
  wire v8aea38;
  wire v844fa0;
  wire v8b327a;
  wire v8aeab1;
  wire v8b6e0a;
  wire v8b12eb;
  wire v91273c;
  wire v8c0bf1;
  wire v912780;
  wire v912668;
  wire v844f9e;
  wire v8aff01;
  wire v9126c4;
  wire v912745;
  wire v911fdd;
  wire v8b279b;
  wire v91116d;
  wire v91258f;
  wire v911cf2;
  wire v8ae7ea;
  wire v912709;
  wire v8af452;
  wire v8b2fd3;
  wire v9123eb;
  wire v8924fb;
  wire v8c7054;
  wire v9114a2;
  wire v8b2878;
  wire v844f95;
  wire v8a8ba3;
  wire v8c6bfa;
  wire v8b1e7d;
  wire v9125d2;
  wire v911f72;
  wire v9123fe;
  wire v8c0435;
  wire v8b0e8e;
  wire v8b004e;
  wire v91187a;
  wire v8b0823;
  wire v8b21ba;
  wire v8c3050;
  wire v8b2bd9;
  wire v9126d5;
  wire v9113da;
  wire v8b0945;
  wire v9112bc;
  wire v9121d1;
  wire v8b1161;
  wire v8b0a12;
  wire v8af82e;
  wire v9124c4;
  wire v9124e1;
  wire v8b32c1;
  wire v8e9855;
  wire v8c049b;
  wire v8af53c;
  wire v8b2464;
  wire v8e98d2;
  wire v8ae162;
  wire v892893;
  wire v844faf;
  wire v912548;
  wire v912711;
  wire v912698;
  wire v8b33d3;
  wire v911075;
  wire v8b1eff;
  wire v8ae6ab;
  wire v911219;
  wire v8ae925;
  wire v8b3c24;
  wire v9110f5;
  wire v91271d;
  wire v88709f;
  wire v912520;
  wire v8d6d04;
  wire v912609;
  wire v8aefe5;
  wire v8b2789;
  wire v8b293f;
  wire v8b2ddd;
  wire v8c568f;
  wire v8b1e7b;
  wire v890ac7;
  wire v8c5c8c;
  wire v9124c3;
  wire v9125a0;
  wire v91118f;
  wire v8b12af;
  wire v9126de;
  wire v8b27f9;
  wire v8c4a3e;
  wire v8af808;
  wire v9126a1;
  wire v8b2c79;
  wire v91130e;
  wire v912408;
  wire v91267e;
  wire v8b2e24;
  wire v8db217;
  wire v8af4ee;
  wire v9125d7;
  wire v8c23d2;
  wire v91245f;
  wire v8b0753;
  wire v8b2c5d;
  wire v8b2b2d;
  wire v8ae714;
  wire v8ae88e;
  wire v8ae151;
  wire v8af894;
  wire v8fed5e;
  wire v892858;
  wire v911fbe;
  wire v9123ba;
  wire v8af275;
  wire v85a510;
  wire v912593;
  wire v8c3e7e;
  wire v8c49c6;
  wire v89098b;
  wire v912507;
  wire v8af192;
  wire v8b21c9;
  wire v912122;
  wire v8aff68;
  wire v8aea95;
  wire v844fb7;
  wire v8afea6;
  wire v9123ef;
  wire v8afdde;
  wire v8c6bef;
  wire v9125ad;
  wire v8b251f;
  wire v8aee6c;
  wire v91263c;
  wire v8b1195;
  wire v910efa;
  wire v8c0443;
  wire v912474;
  wire v8b2445;
  wire v911e75;
  wire v8ae6ee;
  wire v8b1385;
  wire v8c6cd3;
  wire v8cc202;
  wire v91275f;
  wire v912080;
  wire v8b2ae9;
  wire v8c6a96;
  wire v8fed23;
  wire v8c43ba;
  wire v8af9f2;
  wire v8c4c96;
  wire v8afdec;
  wire v8b23d4;
  wire v8c3cff;
  wire v8b4fb2;
  wire v882969;
  wire v9115c6;
  wire v8b5a58;
  wire v8d6d16;
  wire v8b10c6;
  wire v912765;
  wire v8b2ab3;
  wire v9126d9;
  wire v8c6dff;
  wire v8fed7c;
  wire v8afb03;
  wire v8c72da;
  wire v8cc1e2;
  wire v89407e;
  wire v91274f;
  wire v910c69;
  wire v9110c2;
  wire v91270f;
  wire v8b12b1;
  wire v8e9859;
  wire v910bbe;
  wire v8b788f;
  wire v8b12be;
  wire v8b2792;
  wire v8b24cc;
  wire v8c5cc7;
  wire v8ae81f;
  wire v8af8f5;
  wire v8b2a2e;
  wire v9123e0;
  wire v8894e7;
  wire v88abf5;
  wire v87d0f8;
  wire v91266e;
  wire v9126bc;
  wire v890b4a;
  wire v91157e;
  wire v9123c6;
  wire v8b2e70;
  wire v8c09e5;
  wire v9112aa;
  wire v8c5e9b;
  wire v8af624;
  wire v8c0bc2;
  wire v91253f;
  wire v8af39f;
  wire v912450;
  wire v87d059;
  wire v91270b;
  wire v8af0fb;
  wire v912543;
  wire v912631;
  wire v8db203;
  wire v890b41;
  wire v8af004;
  wire v8e9884;
  wire v8b26af;
  wire v8ba4a1;
  wire v912756;
  wire v912657;
  wire v91151f;
  wire v912692;
  wire v8b0e67;
  wire v8c56dd;
  wire v8aef35;
  wire v8aecf5;
  wire v910e34;
  wire v8afe33;
  wire v85c16c;
  wire v9124ab;
  wire v91188e;
  wire v911fd1;
  wire v8c6e2e;
  wire v8d6d00;
  wire v88227e;
  wire v9124e5;
  wire v8ae83c;
  wire v8feced;
  wire v911fcd;
  wire v8b0e1d;
  wire v8e98e4;
  wire v9123f6;
  wire v8c0acd;
  wire v91254d;
  wire v912761;
  wire v875d13;
  wire v8aec34;
  wire v887b94;
  wire v912516;
  wire v8c0b6f;
  wire v912706;
  wire v8f960f;
  wire v911a0d;
  wire v8af159;
  wire v8b2812;
  wire v8c53ab;
  wire v8b0c94;
  wire v8b0b0c;
  wire v8b3237;
  wire v8b029c;
  wire v8c39b8;
  wire v91250d;
  wire v8b02de;
  wire v8b217f;
  wire v88df14;
  wire v9121f2;
  wire v8b26ec;
  wire v9123a3;
  wire v9123dd;
  wire v91265c;
  wire v8b2569;
  wire v8af683;
  wire v8db1b0;
  wire v8afe49;
  wire v912496;
  wire v8b0b7f;
  wire v8af340;
  wire v8b2220;
  wire v9112b6;
  wire v9123c2;
  wire v86bf27;
  wire v8b0446;
  wire v8b7801;
  wire v8af0b0;
  wire v8c534d;
  wire v8c3053;
  wire v8b0f2f;
  wire v8af55a;
  wire v911fc3;
  wire v8b002e;
  wire v911bcd;
  wire v8c6c00;
  wire v8c3f33;
  wire v8bfab7;
  wire v8b2fc4;
  wire v8ae722;
  wire v8b08ac;
  wire v8afce6;
  wire v9124f8;
  wire v8b03fe;
  wire v8fec78;
  wire v8e990d;
  wire v8aeeeb;
  wire v912181;
  wire v8c45e8;
  wire v8aef4e;
  wire v8af84d;
  wire v91153e;
  wire v8d14b5;
  wire v8b0a36;
  wire v884a20;
  wire v8b0693;
  wire v91240f;
  wire v8c36a2;
  wire v87dbe0;
  wire v8aeb12;
  wire v8b0dd3;
  wire v8b021e;
  wire v8b01bd;
  wire v8c50eb;
  wire v9124f2;
  wire v911e65;
  wire v912411;
  wire v9111f5;
  wire v912718;
  wire v8b0dd0;
  wire v8db1c7;
  wire v91241a;
  wire v8b52c1;
  wire v911d25;
  wire v8c47c3;
  wire v8c3d52;
  wire v8b2642;
  wire v863493;
  wire v8c0433;
  wire v8f9724;
  wire v844fb1;
  wire v8b2353;
  wire v8af215;
  wire v9125e3;
  wire v912190;
  wire v9115b8;
  wire v912487;
  wire v912702;
  wire v88b300;
  wire v91215f;
  wire v912683;
  wire v8c4a47;
  wire v8909eb;
  wire v8c7305;
  wire v8afd2b;
  wire v8c5357;
  wire v8b2180;
  wire v879d5b;
  wire v8af431;
  wire v8b11a0;
  wire v911797;
  wire v911fc2;
  wire v8b3d12;
  wire v910ba7;
  wire v912182;
  wire v911d7e;
  wire v887c34;
  wire v9120ec;
  wire v8b0633;
  wire v8c4a25;
  wire v8c6cee;
  wire v8c390a;
  wire v911fd2;
  wire v8ae93f;
  wire v912636;
  wire v8af193;
  wire v8c4072;
  wire v8d540a;
  wire v8aed0c;
  wire v8ae048;
  wire v8ae12e;
  wire v8ae0b8;
  wire v8b7794;
  wire v91265d;
  wire v8b11f0;
  wire v8ae77f;
  wire v8b1a14;
  wire v8b2f6b;
  wire v8ae446;
  wire v9126da;
  wire v8b1130;
  wire v8b1dbd;
  wire v912505;
  wire v887bdb;
  wire v8b222c;
  wire v8af410;
  wire v8c3af9;
  wire v8b23d9;
  wire v91269d;
  wire v88fef2;
  wire v8b1d1f;
  wire v912414;
  wire v8742de;
  wire v8b2fc3;
  wire v88ed6a;
  wire v845125;
  wire v8e98af;
  wire v8b76c6;
  wire v8ae673;
  wire v9125e8;
  wire v8b1e70;
  wire v8c34ba;
  wire v8ae8bf;
  wire v8b114d;
  wire v85c0eb;
  wire v911e3b;
  wire v91238f;
  wire v86ce5c;
  wire v8b0f42;
  wire v8b2e72;
  wire v8b0acf;
  wire v8b1e33;
  wire v8fed5b;
  wire v8c3619;
  wire v8bfa1e;
  wire v911fa7;
  wire v91268f;
  wire v91194c;
  wire v8c420b;
  wire v8b2ba6;
  wire v911e1d;
  wire v8b070e;
  wire v912522;
  wire v911bc6;
  wire v8b0d57;
  wire v8b2ac2;
  wire v8e5d29;
  wire v8ae5e2;
  wire v8aeef8;
  wire v8aee79;
  wire v911173;
  wire v8b265b;
  wire v894810;
  wire v8b0358;
  wire v912628;
  wire v8b085a;
  wire v912201;
  wire v8ae582;
  wire v8c5781;
  wire v8ae7de;
  wire v8af1e9;
  wire v8ae806;
  wire v912154;
  wire v8b1ea2;
  wire v8f96e8;
  wire v91180a;
  wire v9123bf;
  wire v8b25f9;
  wire v890c1b;
  wire v8ae4a3;
  wire v9124a0;
  wire v8b1fc5;
  wire v8b209b;
  wire v9124ef;
  wire v8af3b2;
  wire v8ae765;
  wire v8c42f9;
  wire v91219b;
  wire v9123c7;
  wire v9123b7;
  wire v8c4569;
  wire v8c460a;
  wire v8b0599;
  wire v8dd637;
  wire v8b2fea;
  wire v8b1247;
  wire v8b1003;
  wire v89217c;
  wire v8af6e2;
  wire v8af8b0;
  wire v8aeaf7;
  wire v9124d5;
  wire v8b26cf;
  wire v8ae6c7;
  wire v912428;
  wire v8b2843;
  wire v8cc1a9;
  wire v8b1cbb;
  wire v91278c;
  wire v8f9625;
  wire v8aee21;
  wire v8c71fb;
  wire v9123e2;
  wire v91244b;
  wire v8e98d6;
  wire v911ea9;
  wire v8afcf7;
  wire v91119d;
  wire v8b02ab;
  wire v8b1086;
  wire v912589;
  wire v8b09b0;
  wire v85c141;
  wire v911529;
  wire v911e40;
  wire v912752;
  wire v8b05b0;
  wire v8c7385;
  wire v8940d8;
  wire v8b2c4e;
  wire v8b2c52;
  wire v8af601;
  wire v8c55bf;
  wire v8aea93;
  wire v8b02dd;
  wire v87bd82;
  wire v8c0a9d;
  wire v8b25f8;
  wire v91241f;
  wire v86d734;
  wire v911f49;
  wire v912276;
  wire v8b24e9;
  wire v8fedea;
  wire v890a64;
  wire v8b07d3;
  wire v887bcc;
  wire v8b3383;
  wire v892f3e;
  wire v91273e;
  wire v912690;
  wire v91258e;
  wire v8884e5;
  wire v9125ab;
  wire v8cc1c4;
  wire v9126c3;
  wire v8e990e;
  wire v88ef39;
  wire v8fedc9;
  wire v8b2345;
  wire v8c3e7d;
  wire v8aeabb;
  wire v91177e;
  wire v8afed8;
  wire v8aea7b;
  wire v912739;
  wire v8c4189;
  wire v8fecb7;
  wire v9123c5;
  wire v911631;
  wire v8b244c;
  wire v8c4b6c;
  wire v8b1e9a;
  wire v911f8b;
  wire v8b0d4e;
  wire v8afdfc;
  wire v8b23e9;
  wire v912407;
  wire v88e856;
  wire v8c3fcf;
  wire v9124dd;
  wire v9125c8;
  wire v8af586;
  wire v8c48a8;
  wire v91275d;
  wire v912471;
  wire v912448;
  wire v8b24af;
  wire v8af98a;
  wire v912490;
  wire v912575;
  wire v8afd20;
  wire v912485;
  wire v8b2a9f;
  wire v8af1ad;
  wire v910f9a;
  wire v8c6dfc;
  wire v8af960;
  wire v912420;
  wire v8b01a4;
  wire v8b0963;
  wire v8af2e0;
  wire v8ae8e3;
  wire v911fdf;
  wire v8b12e9;
  wire v8afa40;
  wire v890880;
  wire v8cc139;
  wire v8b0dd9;
  wire v8b9047;
  wire v8b0903;
  wire v8b0b70;
  wire v911733;
  wire v8aeb6d;
  wire v8b2998;
  wire v8b2cc1;
  wire v912768;
  wire v8b2d5a;
  wire v8b0fac;
  wire v8dd5e1;
  wire v8674d8;
  wire v8c04cb;
  wire v8c0b07;
  wire v912679;
  wire v912728;
  wire v912442;
  wire v88abc8;
  wire v8b0113;
  wire v8af478;
  wire v9107fb;
  wire v9124f6;
  wire v8af5b7;
  wire v91220c;
  wire v8ae83f;
  wire v8b0e4c;
  wire v911367;
  wire v8b2aad;
  wire v9124c5;
  wire v8b0e6d;
  wire v8b08c4;
  wire v9123b3;
  wire v8b3321;
  wire v8af3eb;
  wire v9124b0;
  wire v85915c;
  wire v88bebc;
  wire v8b00a9;
  wire v91256e;
  wire v8c6cae;
  wire v91247b;
  wire v8afedf;
  wire v8b1e10;
  wire v8b2a7e;
  wire v8afcaa;
  wire v8aee3c;
  wire v8b1ec4;
  wire v9123cc;
  wire v912515;
  wire v8b016d;
  wire v8af2ab;
  wire v8b284f;
  wire v911eb5;
  wire v911fbd;
  wire v91100d;
  wire v8ae4cd;
  wire v8b1248;
  wire v87cf78;
  wire v8b2bc5;
  wire v912198;
  wire v89097b;
  wire v8af430;
  wire v8b05e2;
  wire v8908a2;
  wire v8b0b9e;
  wire v8b330f;
  wire v8b2c68;
  wire v912790;
  wire v912699;
  wire v8b2484;
  wire v8ae668;
  wire v912666;
  wire v8b0e72;
  wire v91259f;
  wire v8b0fee;
  wire v8dd687;
  wire v912283;
  wire v8ae041;
  wire v8ae713;
  wire v91255d;
  wire v912525;
  wire v8b0f67;
  wire v8b0211;
  wire v8c575b;
  wire v8afc36;
  wire v9123c1;
  wire v8ae8d3;
  wire v912716;
  wire v8b016c;
  wire v8c3c40;
  wire v8b068b;
  wire v9122e7;
  wire v887bcf;
  wire v8c5239;
  wire v8ae46b;
  wire v8ae9f4;
  wire v8afd31;
  wire v9125dd;
  wire v87cd98;
  wire v8d6d2c;
  wire v8afa70;
  wire v894826;
  wire v910c73;
  wire v912717;
  wire v911e94;
  wire v8b2d68;
  wire v9111c2;
  wire v8c0aba;
  wire v911fd6;
  wire v8d6d0f;
  wire v8e5d84;
  wire v8c043b;
  wire v85c148;
  wire v8af986;
  wire v890992;
  wire v8afa3c;
  wire v8ae887;
  wire v911dbb;
  wire v8af305;
  wire v88b266;
  wire v88f72f;
  wire v870559;
  wire v8b20fa;
  wire v8b101c;
  wire v8b2929;
  wire v8b77ed;
  wire v8afaa6;
  wire v8aeb4c;
  wire v8afea2;
  wire v8b091d;
  wire v8afb96;
  wire v8b2c29;
  wire v9123cd;
  wire v8b28d5;
  wire v8af811;
  wire v912723;
  wire v9125b6;
  wire v8b7bb3;
  wire v8af618;
  wire v911fae;
  wire v912695;
  wire v8c500e;
  wire v9118c2;
  wire v8b276b;
  wire v8b2633;
  wire v8940f1;
  wire v844fbb;
  wire v9123d1;
  wire v8c557b;
  wire v8b2a71;
  wire v8c715a;
  wire v912796;
  wire v8b3382;
  wire v9115ca;
  wire v8afb09;
  wire v8af240;
  wire v91250e;
  wire v8b073b;
  wire v911d44;
  wire v8b0463;
  wire v910df3;
  wire v9123c8;
  wire v91174f;
  wire v8af168;
  wire v8b0dd4;
  wire v8940eb;
  wire v8b2e23;
  wire v912691;
  wire v8ae461;
  wire v8b0569;
  wire v864291;
  wire v8909ff;
  wire v8b0c7c;
  wire v8b290b;
  wire v8b1c79;
  wire v8b2d4a;
  wire v8af382;
  wire v8b120b;
  wire v9126ae;
  wire v8b2df8;
  wire v9124c8;
  wire v8e984d;
  wire v8b6d7e;
  wire v85d9b6;
  wire v910cab;
  wire v912656;
  wire v912632;
  wire v8ae696;
  wire v8c4667;
  wire v8b25a8;
  wire v8b03c8;
  wire v8c6c2f;
  wire v8ae7e5;
  wire v9125da;
  wire v887b47;
  wire v8cc182;
  wire v911fa4;
  wire v9126c6;
  wire v8b2610;
  wire v912499;
  wire v9123ab;
  wire v912550;
  wire v9123ee;
  wire v9123a9;
  wire v8b252f;
  wire v8b210b;
  wire v91259a;
  wire v9125f8;
  wire v8b2080;
  wire v87c076;
  wire v912652;
  wire v8b0611;
  wire v9123f5;
  wire v91161f;
  wire v8b2275;
  wire v911742;
  wire v8af651;
  wire v912750;
  wire v88b998;
  wire v8c5d1b;
  wire v9114e1;
  wire v8fece1;
  wire v8b2b44;
  wire v8b28c6;
  wire v91104c;
  wire v869f57;
  wire v8c3541;
  wire v8b3403;
  wire v89342c;
  wire v8c0429;
  wire v8afb9b;
  wire v8b1129;
  wire v8c6c93;
  wire v8afa37;
  wire v9113a8;
  wire v8e9842;
  wire v8b2252;
  wire v912627;
  wire v91256c;
  wire v8b0d58;
  wire v8b07ff;
  wire v9126cc;
  wire v8b296a;
  wire v8aea07;
  wire v8b1ec0;
  wire v8b3d0c;
  wire v91271f;
  wire v912236;
  wire v8b6d47;
  wire v8b2559;
  wire v9125b0;
  wire v8c3efe;
  wire v8b280c;
  wire v890c16;
  wire v9110bb;
  wire v8b3357;
  wire v8b2cf0;
  wire v8ae854;
  wire v8af052;
  wire v8b2885;
  wire v91115b;
  wire v8ae074;
  wire v8784da;
  wire v912685;
  wire v9124f9;
  wire v8c55e1;
  wire v8b2420;
  wire v882fb4;
  wire v8c049e;
  wire v8c6e8e;
  wire v911d0e;
  wire v892ea4;
  wire v8c7026;
  wire v912592;
  wire v911fe3;
  wire v8b77f9;
  wire v8ae731;
  wire v8924ff;
  wire v8b3399;
  wire v8b0494;
  wire v9115c7;
  wire v911538;
  wire v8cc0f1;
  wire v8b2a14;
  wire v91261a;
  wire v9125ec;
  wire v87ab76;
  wire v8c466d;
  wire v9125a9;
  wire v8b2bc3;
  wire v8b2c0d;
  wire v87ed24;
  wire v8af4fa;
  wire v863839;
  wire v8b0681;
  wire v8b2a8d;
  wire v8b10bf;
  wire v9125af;
  wire v8b2e42;
  wire v85aa58;
  wire v8b2a63;
  wire v912466;
  wire v8ae6e2;
  wire v87bd1c;
  wire v8af7cb;
  wire v8b0584;
  wire v8b109a;
  wire v890ab8;
  wire v8aeccb;
  wire v8afdb9;
  wire v911e03;
  wire v85c182;
  wire v844fad;
  wire v8e988e;
  wire v890ac0;
  wire v8b0260;
  wire v8b016b;
  wire v8ae5a8;
  wire v8f9632;
  wire v87a52a;
  wire v8b2e60;
  wire v8c6c4a;
  wire v8db1b1;
  wire v8c5058;
  wire v8ae825;
  wire v8b22a7;
  wire v85db55;
  wire v8af0e3;
  wire v8c0ae6;
  wire v91256f;
  wire v8c6ccc;
  wire v85a47c;
  wire v8b021d;
  wire v912432;
  wire v8b0496;
  wire v8db139;
  wire v8b22ef;
  wire v8af9be;
  wire v8af36f;
  wire v912568;
  wire v8af949;
  wire v89223a;
  wire v911e6a;
  wire v8b140a;
  wire v9126b0;
  wire v91247e;
  wire v8af06b;
  wire v911d4f;
  wire v912784;
  wire v912291;
  wire v8b2553;
  wire v8e983b;
  wire v8b2e92;
  wire v8b2a5b;
  wire v8b02d7;
  wire v8b1d1e;
  wire v8b10fd;
  wire v8dd5d4;
  wire v8b0808;
  wire v9123d4;
  wire v8b2c06;
  wire v8affb3;
  wire v863629;
  wire v8890ee;
  wire v890ba5;
  wire v8b1de3;
  wire v91268b;
  wire v9125d8;
  wire v912732;
  wire v8b0d9e;
  wire v9126e7;
  wire v8b21a3;
  wire v8b2ca9;
  wire v8b244a;
  wire v8c498b;
  wire v9123b1;
  wire v8c4d16;
  wire v912074;
  wire v8aea9f;
  wire v87cf71;
  wire v8b1083;
  wire v912514;
  wire v9124e0;
  wire v8aed6c;
  wire v8b1ec1;
  wire v8b2173;
  wire v8aec65;
  wire v888766;
  wire v8b266b;
  wire v8b066c;
  wire v8c09de;
  wire v8b11ef;
  wire v8b2df3;
  wire v8dd6bd;
  wire v8b24b0;
  wire v8c3e60;
  wire v8ae02f;
  wire v8ae740;
  wire v8b04f8;
  wire v8c3e1b;
  wire v8b28a7;
  wire v8b261e;
  wire v8bfa5d;
  wire v8b0223;
  wire v8b2262;
  wire v8aedac;
  wire v8b25ff;
  wire v9126f9;
  wire v8b76f2;
  wire v8b12ad;
  wire v8af0b5;
  wire v912600;
  wire v8c23d1;
  wire v8b1cf2;
  wire v9126c2;
  wire v9125c5;
  wire v8b2c39;
  wire v8e9954;
  wire v8afde2;
  wire v911ef0;
  wire v8af83a;
  wire v912529;
  wire v8af34a;
  wire v8aedc6;
  wire v8b1ca6;
  wire v8b1245;
  wire v91259b;
  wire v9123c4;
  wire v8aea76;
  wire v912102;
  wire v91264b;
  wire v91230d;
  wire v9126ff;
  wire v8b0b63;
  wire v8ae805;
  wire v8b0554;
  wire v91093d;
  wire v912584;
  wire v8c70dc;
  wire v911940;
  wire v9124ea;
  wire v911b07;
  wire v8bfaf2;
  wire v8c4d14;
  wire v8b068c;
  wire v8b2fc8;
  wire v8ae46d;
  wire v9123c9;
  wire v8c5bc3;
  wire v8b2267;
  wire v912558;
  wire v8b2088;
  wire v890246;
  wire v8f953d;
  wire v8827a3;
  wire v8b2bbf;
  wire v8b1ddc;
  wire v8ae06b;
  wire v8affe3;
  wire v911fb3;
  wire v8db22c;
  wire v8af03b;
  wire v91155b;
  wire v89209f;
  wire v8c57aa;
  wire v911c80;
  wire v912635;
  wire v8b1d03;
  wire v8aeead;
  wire v8c40de;
  wire v9126a9;
  wire v8ae8e5;
  wire v912556;
  wire v91266f;
  wire v91251c;
  wire v91171d;
  wire v8b1410;
  wire v8b3320;
  wire v8b321d;
  wire v8af0e8;
  wire v8b102a;
  wire v8618ae;
  wire v8c23c8;
  wire v8fec8f;
  wire v8aff15;
  wire v91263e;
  wire v8ae4ee;
  wire v8dd5ff;
  wire v912743;
  wire v9123a8;
  wire v91245a;
  wire v8b028f;
  wire v8c706b;
  wire v8b3416;
  wire v8b0a19;
  wire v912598;
  wire v8b04fc;
  wire v8c7153;
  wire v8e98f8;
  wire v859e1d;
  wire v8b1e11;
  wire v912604;
  wire v91276f;
  wire v91258c;
  wire v8bfab2;
  wire v911e68;
  wire v8b8e79;
  wire v8ae8e8;
  wire v911714;
  wire v912326;
  wire v911de3;
  wire v890a73;
  wire v8b1c7b;
  wire v8b257f;
  wire v911bf3;
  wire v8fed1e;
  wire v912547;
  wire v870c3a;
  wire v85c135;
  wire v9125cb;
  wire v8612be;
  wire v8dd5d9;
  wire v8b2f44;
  wire v887ae1;
  wire v8b33af;
  wire v91243d;
  wire v8b340b;
  wire v8b03d4;
  wire v911f9c;
  wire v9126db;
  wire v912729;
  wire v91144e;
  wire v912423;
  wire v911e5a;
  wire v8b0cbf;
  wire v8b1ddf;
  wire v88ac88;
  wire v8b013b;
  wire v8aff37;
  wire v8af767;
  wire v8af71d;
  wire v8c3d77;
  wire v8af1de;
  wire v8af5f1;
  wire v91180c;
  wire v8dd6ad;
  wire v91269c;
  wire v85c13e;
  wire v8b25d9;
  wire v890bcb;
  wire v8c3926;
  wire v8ae160;
  wire v8fec67;
  wire v9123b6;
  wire v911a08;
  wire v8dd6de;
  wire v9123f4;
  wire v8ae934;
  wire v91243a;
  wire v8af640;
  wire v8b2d73;
  wire v89097f;
  wire v91255f;
  wire v8b1eeb;
  wire v8b1d83;
  wire v8cfeeb;
  wire v910ea7;
  wire v8b2e31;
  wire v87de99;
  wire v8b1f58;
  wire v8b01dd;
  wire v8db28c;
  wire v910e18;
  wire v8af6d0;
  wire v8b0283;
  wire v8b28e6;
  wire v89092e;
  wire v912451;
  wire v88acc3;
  wire v8af634;
  wire v8b229e;
  wire v9123df;
  wire v8ae878;
  wire v8b0661;
  wire v9124f0;
  wire v8b0151;
  wire v8dd5cf;
  wire v859212;
  wire v8b0dc3;
  wire v8b2911;
  wire v87ebfd;
  wire v9126eb;
  wire v8b2a3e;
  wire v8f9614;
  wire v8af27d;
  wire v8dd65f;
  wire v8ae578;
  wire v8b2a92;
  wire v8b3212;
  wire v8af62a;
  wire v8b52f7;
  wire v91260b;
  wire v8c71b4;
  wire v890a66;
  wire v8b101e;
  wire v8ae9bd;
  wire v8c54b4;
  wire v87a09b;
  wire v8c5404;
  wire v875f27;
  wire v8aea72;
  wire v912391;
  wire v8aeec4;
  wire v8b05a5;
  wire v9123cb;
  wire v8af886;
  wire v8af102;
  wire v8b0fb5;
  wire v8b8bdf;
  wire v8c43e6;
  wire v8ae0ee;
  wire v87b5cf;
  wire v8b12f9;
  wire v8b20b7;
  wire v8b22d1;
  wire v8af9bd;
  wire v8b0219;
  wire v8b27ec;
  wire v91264a;
  wire v85c157;
  wire v8af72b;
  wire v8b64b8;
  wire v8afb82;
  wire v8b2bd8;
  wire v8aec42;
  wire v8af89d;
  wire v910947;
  wire v9123cf;
  wire v8b05b7;
  wire v911ad5;
  wire v912565;
  wire v8af9ff;
  wire v8af2f5;
  wire v8af77e;
  wire v8aebed;
  wire v8b131b;
  wire v9123d3;
  wire v8b1dbe;
  wire v91259d;
  wire v8afab8;
  wire v8aeb67;
  wire v8ae768;
  wire v8b2688;
  wire v8c369a;
  wire v890c50;
  wire v9124ff;
  wire v8ae97e;
  wire v8b4fca;
  wire v8b241a;
  wire v8afd1f;
  wire v8af763;
  wire v912409;
  wire v911792;
  wire v9124d8;
  wire v911ae3;
  wire v844fb5;
  wire v8b2e66;
  wire v9112e0;
  wire v8af864;
  wire v8afd4d;
  wire v9114ce;
  wire v8af214;
  wire v8c458b;
  wire v8f965b;
  wire v8afb18;
  wire v910fe2;
  wire v8b2aeb;
  wire v8b0a03;
  wire v844fb3;
  wire v91272d;
  wire v911e9b;
  wire v911695;
  wire v912783;
  wire v9126c1;
  wire v91276a;
  wire v8b11c4;
  wire v911382;
  wire v912733;
  wire v88331f;
  wire v8596e1;
  wire v911978;
  wire v8b0f51;
  wire v8c59a9;
  wire v8b1014;
  wire v87cf74;
  wire v8af1d7;
  wire v8dd5d8;
  wire v8db20a;
  wire v8b0207;
  wire v911e0c;
  wire v912401;
  wire v911ee4;
  wire v8b13ca;
  wire v8b0ae4;
  wire v887b30;
  wire v9124cf;
  wire v8bfa4c;
  wire v8afcf5;
  wire v8aebc7;
  wire v9123fa;
  wire v9125a6;
  wire v912749;
  wire v8b0c81;
  wire v9126aa;
  wire v8b32b6;
  wire v8af2b1;
  wire v9124a9;
  wire v8b051c;
  wire v8b19b1;
  wire v912470;
  wire v911ff4;
  wire v8b0107;
  wire v8b051e;
  wire v8b08fa;
  wire v912753;
  wire v8af563;
  wire v8b8be1;
  wire v8bfa76;
  wire v8d6ceb;
  wire v8bfa26;
  wire v912465;
  wire v8b71c1;
  wire v8af5fe;
  wire v9123aa;
  wire v912462;
  wire v8b1e8a;
  wire v910cda;
  wire v8af1d2;
  wire v8ae47c;
  wire v91248b;
  wire v8c0a23;
  wire v912669;
  wire v8b2a8f;
  wire v8d6cde;
  wire v9125a5;
  wire v8b0626;
  wire v8bb97f;
  wire v8c6caf;
  wire v8b2049;
  wire v8b2ad6;
  wire v9123e6;
  wire v8b21bb;
  wire v8af036;
  wire v9126f0;
  wire v912508;
  wire v8afe97;
  wire v8c7159;
  wire v8b2aaa;
  wire v8b055a;
  wire v8fecf0;
  wire v910d0e;
  wire v8c4c30;
  wire v911484;
  wire v912786;
  wire v8b0d89;
  wire v8b23de;
  wire v8689df;
  wire v8cc104;
  wire v8b2f4e;
  wire v8aff75;
  wire v8b2c35;
  wire v8ae4b6;
  wire v8af40b;
  wire v911fb2;
  wire v8afabd;
  wire v912681;
  wire v8b13f6;
  wire v89286e;
  wire v8ae803;
  wire v88bb7a;
  wire v8e9903;
  wire v8c4c08;
  wire v876670;
  wire v892555;
  wire v8ae5c0;
  wire v8af78e;
  wire v8b2eb4;
  wire v91277d;
  wire v8b0877;
  wire v8b2ba1;
  wire v8afed5;
  wire v912114;
  wire v911304;
  wire v8b0d99;
  wire v911fb6;
  wire v8b2021;
  wire v88fa8c;
  wire v8e9896;
  wire v8b01d5;
  wire v8b0449;
  wire v8b233e;
  wire v8b2eed;
  wire v8b32e2;
  wire v8ae07b;
  wire v86b11f;
  wire v9125d3;
  wire v8b1dfe;
  wire v8b65a2;
  wire v8b1cd7;
  wire v8aec17;
  wire v8b11df;
  wire v912591;
  wire v8fecd9;
  wire v8aed7b;
  wire v9113d6;
  wire v912542;
  wire v8af52b;
  wire v8c56de;
  wire v9126d4;
  wire v91255a;
  wire v912555;
  wire v8af0e6;
  wire v8b22fd;
  wire v8c41af;
  wire v8c6cb4;
  wire v890be4;
  wire v91268d;
  wire v8aef55;
  wire v8b04ba;
  wire v8af524;
  wire v9125ae;
  wire v8c47de;
  wire v912402;
  wire v8b29e2;
  wire v91254a;
  wire v85c0e8;
  wire v9125f2;
  wire v8b113b;
  wire v9123ce;
  wire v8b1e15;
  wire v8dd5ec;
  wire v91264e;
  wire v9126d8;
  wire v911fac;
  wire v8b0648;
  wire v9116e0;
  wire v9123d7;
  wire v8b0cd4;
  wire v911a8d;
  wire v8b07bc;
  wire v8b05f1;
  wire v8b07b6;
  wire v8ae031;
  wire v8dd632;
  wire v9124db;
  wire v8b2df5;
  wire v9121ee;
  wire v91240a;
  wire v8b648c;
  wire v8c44cf;
  wire v8ae4ce;
  wire v911cec;
  wire v911441;
  wire v9114d3;
  wire v890b86;
  wire v8c45bc;
  wire v8c0aef;
  wire v9124e7;
  wire v8afa41;
  wire v8af1ef;
  wire v8aeabf;
  wire v8c3925;
  wire v8af2e3;
  wire v8b0942;
  wire v9124df;
  wire v8b2460;
  wire v8fee03;
  wire v8b07a1;
  wire v8af9e8;
  wire v8b23c7;
  wire v91240c;
  wire v912549;
  wire v9121e7;
  wire v91276d;
  wire v8c45be;
  wire v91265a;
  wire v8af2f9;
  wire v8c3bd5;
  wire v8b0d88;
  wire v91277e;
  wire v8af3b6;
  wire v91239b;
  wire v8c50c4;
  wire v91247c;
  wire v9123ff;
  wire v8af9f6;
  wire v8b2c4c;
  wire v91257a;
  wire v912747;
  wire v8c50c5;
  wire v8c64bf;
  wire v8771a0;
  wire v912517;
  wire v8c38b4;
  wire v8aefa4;
  wire v8b0d78;
  wire v9126f4;
  wire v91277b;
  wire v9113eb;
  wire v8c6aa0;
  wire v9123af;
  wire v8c44a1;
  wire v8c0a48;
  wire v8cffee;
  wire v8c6c56;
  wire v911f38;
  wire v8b085c;
  wire v8b232f;
  wire v8b2c21;
  wire v8b1f47;
  wire v8c4ac3;
  wire v8c71b3;
  wire v887bcd;
  wire v9125e6;
  wire v9125f0;
  wire v890c07;
  wire v8b2b17;
  wire v8c704a;
  wire v911959;
  wire v912501;
  wire v9126cb;
  wire v8ae7c9;
  wire v8b339d;
  wire v8f9659;
  wire v8bfae8;
  wire v8ae936;
  wire v888464;
  wire v8b0934;
  wire v8c0456;
  wire v8b1f50;
  wire v9116aa;
  wire v8b0e50;
  wire v8ae556;
  wire v911f9b;
  wire v911c5d;
  wire v893433;
  wire v9126b2;
  wire v9125c7;
  wire v8b25e2;
  wire v890c2c;
  wire v8b7379;
  wire v8ae69b;
  wire v8c0ab9;
  wire v910ff3;
  wire v912492;
  wire v8aed7c;
  wire v8b2576;
  wire v911772;
  wire v88e0ec;
  wire v8b22f0;
  wire v8afc88;
  wire v90c2e3;
  wire v912482;
  wire v8b26f3;
  wire v911c25;
  wire v8b1f2d;
  wire v8c353f;
  wire v910bd1;
  wire v8cf811;
  wire v8c050d;
  wire v87e29c;
  wire v8aeb97;
  wire v8b29d8;
  wire v8fed12;
  wire v8b20ab;
  wire v9122d7;
  wire v8b1154;
  wire v9032d6;
  wire v8f9622;
  wire v8b2b57;
  wire v8aebd0;
  wire v8b094a;
  wire v8c3b8d;
  wire v87b940;
  wire v8af765;
  wire v91260c;
  wire v8b076f;
  wire v911fda;
  wire v8b76c0;
  wire v8c044b;
  wire v8f9721;
  wire v8c23b9;
  wire v85c164;
  wire v8ae0c6;
  wire v87b54c;
  wire v911aa3;
  wire v8b2f6c;
  wire v8b0d32;
  wire v8ae5ca;
  wire v8c77fe;
  wire v912521;
  wire v9126c8;
  wire v8b0b98;
  wire v8b050b;
  wire v912416;
  wire v8ae9bf;
  wire v87f443;
  wire v8b02b9;
  wire v8af74b;
  wire v8c5192;
  wire v8c5d1c;
  wire v91243f;
  wire v8af518;
  wire v8c6979;
  wire v85c0bd;
  wire v91151a;
  wire v912537;
  wire v8924d2;
  wire v8afd76;
  wire v8f9617;
  wire v91222a;
  wire v911149;
  wire v8b0e57;
  wire v8ae5ff;
  wire v8b06bc;
  wire v8aedf2;
  wire v8b29af;
  wire v8ae64c;
  wire v8b0be4;
  wire v912638;
  wire v872c7c;
  wire v8940ac;
  wire v8b1d42;
  wire v8b004c;
  wire v9110d2;
  wire v8db23e;
  wire v8c5356;
  wire v91231e;
  wire v8bfa99;
  wire v8b21fa;
  wire v911017;
  wire v9123bb;
  wire v8c51e1;
  wire v8c4a94;
  wire v9124b7;
  wire v8b0f57;
  wire v8c6e12;
  wire v91257c;
  wire v912413;
  wire v91134e;
  wire v8b077d;
  wire v8b2d17;
  wire v8ae8c2;
  wire v8b0cf9;
  wire v887c3b;
  wire v9124ed;
  wire v91223a;
  wire v85afd4;
  wire v8affdf;
  wire v8af451;
  wire v8c6c7e;
  wire v9116e8;
  wire v861f8d;
  wire v9126df;
  wire v8aede2;
  wire v8affe8;
  wire v9124fe;
  wire v8b282e;
  wire v8b1fcd;
  wire v8aef95;
  wire v912532;
  wire v912776;
  wire v8b129a;
  wire v912755;
  wire v8b1e80;
  wire v8b02cb;
  wire v911f83;
  wire v8af3e7;
  wire v89017d;
  wire v8c7049;
  wire v8b2629;
  wire v9126ab;
  wire v8b77fc;
  wire v8c0b7c;
  wire v8c6964;
  wire v912467;
  wire v8b08e5;
  wire v8db1d7;
  wire v8c40af;
  wire v8b1ef8;
  wire v911543;
  wire v8b1fee;
  wire v8b2655;
  wire v8af9e6;
  wire v911513;
  wire v8b09ea;
  wire v8ae898;
  wire v911220;
  wire v8b0d0e;
  wire v8b00f2;
  wire v9119da;
  wire v8e9920;
  wire v8b1e6a;
  wire v87bbef;
  wire v9124b4;
  wire v912676;
  wire v89217b;
  wire v8c381a;
  wire v91108c;
  wire v8c537f;
  wire v8c77e6;
  wire v8b6d3d;
  wire v8c36bc;
  wire v8809fb;
  wire v912696;
  wire v8af4b1;
  wire v8b02b0;
  wire v912735;
  wire v8b06d3;
  wire v8b0a04;
  wire v8aeab6;
  wire v8b0653;
  wire v912527;
  wire v8ae60e;
  wire v8c557c;
  wire v8b1cd0;
  wire v91251a;
  wire v91274b;
  wire v8b1406;
  wire v912523;
  wire v8b33fa;
  wire v8af7a3;
  wire v8af094;
  wire v8b1c70;
  wire v8b1fe8;
  wire v912075;
  wire v91216a;
  wire v8c0509;
  wire v91275b;
  wire v8c4517;
  wire v91189f;
  wire v8c6c18;
  wire v8b0b2b;
  wire v8afec3;
  wire v8af80a;
  wire v8c3973;
  wire v8dd5d0;
  wire v8aefc1;
  wire v9126c9;
  wire v91254f;
  wire v8af51f;
  wire v912479;
  wire v8ae92f;
  wire v88b60c;
  wire v912771;
  wire v8b2511;
  wire v8afb17;
  wire v8c4353;
  wire v8dd667;
  wire v91141d;
  wire v8ae909;
  wire v8b1e0b;
  wire v8b09b9;
  wire v912763;
  wire v8b6482;
  wire v912788;
  wire v8b139e;
  wire v911664;
  wire v8b0674;
  wire v8aed74;
  wire v8c0bf4;
  wire v8b048e;
  wire v8c6e5a;
  wire v8b0dc4;
  wire v8af7df;
  wire v8af582;
  wire v892e44;
  wire v861315;
  wire v8af399;
  wire v8c6df7;
  wire v8c0b46;
  wire v8b0dc1;
  wire v8b09b4;
  wire v8b25a4;
  wire v8c4a56;
  wire v8c3651;
  wire v912512;
  wire v8591f3;
  wire v9126b8;
  wire v911faa;
  wire v885d39;
  wire v8b076a;
  wire v86f3ae;
  wire v8af119;
  wire v910e98;
  wire v8c6d04;
  wire v8afd55;
  wire v8c3e35;
  wire v8b22a8;
  wire v8ae956;
  wire v91242f;
  wire v9126b4;
  wire v8af79f;
  wire v887ac4;
  wire v88fa49;
  wire v8b02d5;
  wire v8b038f;
  wire v912744;
  wire v8b3286;
  wire v8aeddc;
  wire v8b6f1f;
  wire v8b24b7;
  wire v911158;
  wire v9119a4;
  wire v912626;
  wire v8b26ee;
  wire v91100c;
  wire v8af2c8;
  wire v912472;
  wire v8b0298;
  wire v8940af;
  wire v91263d;
  wire v8909d0;
  wire v8c04c4;
  wire v8cc197;
  wire v8c043d;
  wire v912680;
  wire v8b1110;
  wire v9123d6;
  wire v8b7802;
  wire v8fed49;
  wire v91255c;
  wire v911aa1;
  wire v912705;
  wire v9124d7;
  wire v9124d6;
  wire v911a76;
  wire v8afc85;
  wire v8b0936;
  wire v8b74aa;
  wire v911fa9;
  wire v9125ce;
  wire v8c57d1;
  wire v8c3617;
  wire v8c39e1;
  wire v8b0429;
  wire v910d87;
  wire v8e9961;
  wire v91257f;
  wire v8c4b39;
  wire v912453;
  wire v8b0500;
  wire v8c3728;
  wire v8b0a89;
  wire v8b0e3d;
  wire v9126ad;
  wire v8db288;
  wire v910d59;
  wire v8aed6d;
  wire v8b2b91;
  wire v8b1f0a;
  wire v8c3c57;
  wire v8b29d6;
  wire v86990d;
  wire v912775;
  wire v912461;
  wire v8b0994;
  wire v91183d;
  wire v8c3a82;
  wire v8c46bf;
  wire v892fa2;
  wire v890960;
  wire v8dd6fe;
  wire v912431;
  wire v8ae096;
  wire v911532;
  wire v8b1dd2;
  wire v85f6d2;
  wire v8b107b;
  wire v9126a8;
  wire v884789;
  wire v8b2935;
  wire v8b2c26;
  wire v8afb06;
  wire v9123ad;
  wire v8b0c67;
  wire v890534;
  wire v8c6cdc;
  wire v8af415;
  wire v9124c6;
  wire v8b0264;
  wire v911c2f;
  wire v8b0b29;
  wire v87cfd0;
  wire v8c5fa2;
  wire v8c6bba;
  wire v8579b7;
  wire v8aee49;
  wire v91246a;
  wire v9123f8;
  wire v9115fc;
  wire v8b2d92;
  wire v8b1f71;
  wire v9112f7;
  wire v8ae9fc;
  wire v9126b3;
  wire v8c5e4c;
  wire v8b2b5c;
  wire v8b3d17;
  wire v8b07f3;
  wire v8b2e7a;
  wire v8af025;
  wire v912737;
  wire v91261d;
  wire v8ae9f2;
  wire v8c70fc;
  wire v8b3d0e;
  wire v912026;
  wire v91271e;
  wire v8b1367;
  wire v8b03e8;
  wire v8af780;
  wire v8c7263;
  wire v8b062d;
  wire v91278f;
  wire v8b2e07;
  wire v911f9d;
  wire v8b00a7;
  wire v8b267a;
  wire v8c3b68;
  wire v8d6d1f;
  wire v91253d;
  wire v91278b;
  wire v91207b;
  wire v8c41aa;
  wire v8b028a;
  wire v871da5;
  wire v9123e7;
  wire v8b2479;
  wire v8c4a78;
  wire v8afe01;
  wire v8b0119;
  wire v8b7791;
  wire v8aeada;
  wire v8858cb;
  wire v8c3731;
  wire v8c4398;
  wire v8ae437;
  wire v912625;
  wire v8b05ce;
  wire v8b0ef5;
  wire v8ae5c6;
  wire v8c387f;
  wire v8b0762;
  wire v8b1fb5;
  wire v911c88;
  wire v8b8e74;
  wire v9125b1;
  wire v8afc68;
  wire v8f9587;
  wire v8b22be;
  wire v8fece4;
  wire v91267c;
  wire v912764;
  wire v8af7b5;
  wire v912588;
  wire v912797;
  wire v8ae519;
  wire v8b2e27;
  wire v8af698;
  wire v8b22c9;
  wire v8c510a;
  wire v8af899;
  wire v892e12;
  wire v91268a;
  wire v9114cd;
  wire v8b085e;
  wire v9125b9;
  wire v912722;
  wire v9124e2;
  wire v8fedd4;
  wire v912793;
  wire v9124fb;
  wire v9116c4;
  wire v89098c;
  wire v912660;
  wire v9126b9;
  wire v85e943;
  wire v912714;
  wire v8b1150;
  wire v8af05a;
  wire v8b4d42;
  wire v8b7669;
  wire v8af0ef;
  wire v912509;
  wire v8b0436;
  wire v9125df;
  wire v8afa7c;
  wire v9124f5;
  wire v912425;
  wire v8b2493;
  wire v8b0738;
  wire v8b0b24;
  wire v87139e;
  wire v8ae14c;
  wire v8b1178;
  wire v8af463;
  wire v8b26bb;
  wire v91271c;
  wire v912513;
  wire v8b2c07;
  wire v87e9d4;
  wire v9115e4;
  wire v8afaec;
  wire v8cc129;
  wire v910c25;
  wire v8b0d2f;
  wire v8b0eea;
  wire v8b0112;
  wire v912557;
  wire v8b7892;
  wire v91269a;
  wire v8ae02e;
  wire v8bfa79;
  wire v8b099d;
  wire v911a5d;
  wire v8b2e17;
  wire v8ae118;
  wire v8f95dd;
  wire v8fecad;
  wire v8f9631;
  wire v8afa8e;
  wire v8af6c8;
  wire v9126b1;
  wire v8b0b7a;
  wire v8e989e;
  wire v911b46;
  wire v911d0d;
  wire v8c3d99;
  wire v87d240;
  wire v8b0b9c;
  wire v8b2592;
  wire v91240d;
  wire v890964;
  wire v9125d9;
  wire v8b0eb6;
  wire v8cc0fb;
  wire v8aec59;
  wire v8af717;
  wire v8b2868;
  wire v8c6167;
  wire v88704a;
  wire v9125bc;
  wire v910ff6;
  wire v8c4a57;
  wire v8c0b9e;
  wire v8ae03c;
  wire v88b1d7;
  wire v8c5d7e;
  wire v911196;
  wire v911bdc;
  wire v85c126;
  wire v85f3d2;
  wire v8b2838;
  wire v88340e;
  wire v8db195;
  wire v8afb51;
  wire v9123a4;
  wire v8aeb57;
  wire v8b09e6;
  wire v8b0a78;
  wire v8ae588;
  wire v8618ff;
  wire v8afc39;
  wire v8bfa98;
  wire v8c7247;
  wire v8cda2f;
  wire v8afb8e;
  wire v912693;
  wire v912672;
  wire v91116e;
  wire v910c72;
  wire v8b29c1;
  wire v8af253;
  wire v9126e1;
  wire v911d22;
  wire v8af756;
  wire v8dd6ff;
  wire v89287e;
  wire v912331;
  wire v8ae756;
  wire v91243e;
  wire v91248d;
  wire v8b0467;
  wire v8b02e9;
  wire v8b09e5;
  wire v8b33ed;
  wire v8aedb1;
  wire v912616;
  wire v91261f;
  wire v8b4fda;
  wire v9123e3;
  wire v8c3ea2;
  wire v8afa56;
  wire v8aee85;
  wire v9124ce;
  wire v8b297c;
  wire v881e63;
  wire v8b1068;
  wire v8aed2e;
  wire v8b28d4;
  wire v86cbb8;
  wire v912394;
  wire v8aedc9;
  wire v911ffb;
  wire v8b33aa;
  wire v8b289a;
  wire v8b12fb;
  wire v912493;
  wire v91250c;
  wire v8b2c5c;
  wire v8b3402;
  wire v8b2f46;
  wire v91257b;
  wire v8b03ed;
  wire v8b01f5;
  wire v8c6c8b;
  wire v8b2b4a;
  wire v892551;
  wire v8b1d71;
  wire v911a2a;
  wire v87dc9f;
  wire v91134b;
  wire v8ae670;
  wire v912643;
  wire v8c48c7;
  wire v91262d;
  wire v8afe84;
  wire v911ed2;
  wire v8b0a17;
  wire v8c3d4b;
  wire v85d63e;
  wire v912477;
  wire v85f4b2;
  wire v8b134f;
  wire v8af366;
  wire v87b84a;
  wire v8af687;
  wire v91275a;
  wire v9124e6;
  wire v9116ad;
  wire v8c715c;
  wire v8839ea;
  wire v8c3027;
  wire v8cc220;
  wire v911d2c;
  wire v911fad;
  wire v8dd5e6;
  wire v912742;
  wire v8b0fab;
  wire v8dd6ae;
  wire v912502;
  wire v887bd4;
  wire v91183a;
  wire v9126d1;
  wire v911fab;
  wire v911ebd;
  wire v8aef7a;
  wire v912605;
  wire v8af918;
  wire v8c426f;
  wire v8b050c;
  wire v8b340c;
  wire v911fc4;
  wire v8af5df;
  wire v8ae147;
  wire v8aea10;
  wire v8b2f6d;
  wire v8b0a2d;
  wire v91230e;
  wire v86c179;
  wire v8afe06;
  wire v8b12d5;
  wire v91271b;
  wire v8bfa65;
  wire v9123d2;
  wire v8b3350;
  wire v887b1c;
  wire v8b236d;
  wire v9124a4;
  wire v8b2b08;
  wire v8af85c;
  wire v912068;
  wire v912694;
  wire v8692ec;
  wire v912400;
  wire v8af2bd;
  wire v911052;
  wire v8ae561;
  wire v8d6d2e;
  wire v8b1fc7;
  wire v8aec85;
  wire v8aefce;
  wire v912166;
  wire v8c47bf;
  wire v91211a;
  wire v8afc08;
  wire v912563;
  wire v91272e;
  wire v8b7bb1;
  wire v8b0817;
  wire v890ba9;
  wire v8af23b;
  wire v8b28fe;
  wire v911fea;
  wire v8b1d80;
  wire v8b2d82;
  wire v85c0b1;
  wire v912792;
  wire v8b1350;
  wire v8aed35;
  wire v91242d;
  wire v9114aa;
  wire v912658;
  wire v887b53;
  wire v8b65a3;
  wire v8b2a34;
  wire v8c70fd;
  wire v9124b5;
  wire v8af0c8;
  wire v8b27ab;
  wire v8b29ed;
  wire v912480;
  wire v8b6e6f;
  wire v9126dd;
  wire v912785;
  wire v8c3afa;
  wire v8aed37;
  wire v8f9630;
  wire v8c3bb7;
  wire v912046;
  wire v9125fc;
  wire v8b0ae9;
  wire v8b29d9;
  wire v8aecbf;
  wire v8b2fbc;
  wire v9123de;
  wire v91101e;
  wire v9114e3;
  wire v8c0b95;
  wire v8b76ff;
  wire v8b1f1b;
  wire v8b2162;
  wire v910e1f;
  wire v8b274c;
  wire v8d6d2f;
  wire v9125c3;
  wire v911a5e;
  wire v8b09fb;
  wire v912642;
  wire v8b1e0f;
  wire v8b2741;
  wire v9119bc;
  wire v912280;
  wire v91268e;
  wire v911466;
  wire v8d50bc;
  wire v8ae7b3;
  wire v8b0fa3;
  wire v8ae64a;
  wire v8b238a;
  wire v911c7e;
  wire v8b2a8c;
  wire v8b1e22;
  wire v8b0df4;
  wire v8bfa8b;
  wire v8577c2;
  wire v8b2c6b;
  wire v9126f5;
  wire v8c3c0d;
  wire v8c5350;
  wire v9122c8;
  wire v8b09a9;
  wire v8b76f1;
  wire v8b320b;
  wire v8c0b8f;
  wire v911bad;
  wire v8b02a9;
  wire v911f54;
  wire v8c568d;
  wire v912576;
  wire v8bfa61;
  wire v8e990a;
  wire v912403;
  wire v912464;
  wire v88b254;
  wire v91246d;
  wire v8e992f;
  wire v8dd5e2;
  wire v8c0b04;
  wire v881ef0;
  wire v864227;
  wire v910c58;
  wire v8bfa12;
  wire v88ffd6;
  wire v911197;
  wire v88d6cf;
  wire v912766;
  wire v8b1199;
  wire v8b0b6b;
  wire v911633;
  wire v890b35;
  wire v8ae033;
  wire v8b0750;
  wire v8c4a4e;
  wire v8b0e9d;
  wire v8c4cc3;
  wire v8af1a2;
  wire v8c4410;
  wire v8c51d8;
  wire v890a9a;
  wire v8af5bd;
  wire v8c43c1;
  wire v8b29c9;
  wire v912390;
  wire v8f96fd;
  wire v8c4b37;
  wire v8c5e54;
  wire v8aec46;
  wire v8b0642;
  wire v8b216f;
  wire v88413b;
  wire v8ae4a5;
  wire v910c1b;
  wire v8af78a;
  wire v91242c;
  wire v887afb;
  wire v86bd18;
  wire v8c723e;
  wire v8f9597;
  wire v8b0a5f;
  wire v9111d2;
  wire v8b2cb0;
  wire v912748;
  wire v890adc;
  wire v86995b;
  wire v88f796;
  wire v8b082d;
  wire v912664;
  wire v8b2000;
  wire v911bd2;
  wire v911632;
  wire v9124a5;
  wire v8b0ce2;
  wire v8ae789;
  wire v8aeb29;
  wire v8b06b8;
  wire v8db180;
  wire v88547b;
  wire v91269f;
  wire v8b236f;
  wire v910bd3;
  wire v8ae86c;
  wire v8b00fe;
  wire v9124c2;
  wire v8cc164;
  wire v8c34da;
  wire v9123b9;
  wire v8b09f9;
  wire v9126d2;
  wire v912417;
  wire v8b0c90;
  wire v8b76f3;
  wire v8b33f2;
  wire v8b1e43;
  wire v911fa0;
  wire v8cc0f3;
  wire v8c7100;
  wire v8b0cf7;
  wire v8af015;
  wire v9112d7;
  wire v8b09a3;
  wire v8ae8b7;
  wire v8b0bd2;
  wire v8b2a31;
  wire v8b31f9;
  wire v912264;
  wire v8b7443;
  wire v8b2c37;
  wire v8ae75b;
  wire v8f96c9;
  wire v8fecf2;
  wire v890940;
  wire v8b02ed;
  wire v87ba6d;
  wire v911f1c;
  wire v911ef8;
  wire v8e994b;
  wire v8ae51a;
  wire v9123be;
  wire v8b31b3;
  wire v8b04f4;
  wire v911fb1;
  wire v8aec8e;
  wire v9124d4;
  wire v8b0cfd;
  wire v8af2cd;
  wire v911765;
  wire v9124bd;
  wire v8b2876;
  wire v890b15;
  wire v91248a;
  wire v912662;
  wire v8aea88;
  wire v8af7f1;
  wire v894087;
  wire v8b0705;
  wire v87d0a9;
  wire v8c3a0b;
  wire v8b23bf;
  wire v8c5419;
  wire v8dd643;
  wire v8aedf0;
  wire v8b25e8;
  wire v8b0bd4;
  wire v892511;
  wire v8dd5ca;
  wire v9126f7;
  wire v8af155;
  wire v8b01e2;
  wire v8af26f;
  wire v9125d4;
  wire v8ae584;
  wire v8b26ed;
  wire v8af73a;
  wire v91244f;
  wire v8b1ffd;
  wire v883aaa;
  wire v91230c;
  wire v8ae728;
  wire v8b065b;
  wire v91176c;
  wire v8c4740;
  wire v911395;
  wire v871abf;
  wire v8b3d09;
  wire v8b2b80;
  wire v85c0ac;
  wire v8b11b0;
  wire v8b08ff;
  wire v8b22c6;
  wire v8b0fb9;
  wire v8c458d;
  wire v8c3a85;
  wire v9123f7;
  wire v8872e8;
  wire v8c37c9;
  wire v8c426e;
  wire v8fed10;
  wire v911a6a;
  wire v8b1ff8;
  wire v91251b;
  wire v911b49;
  wire v911291;
  wire v866ac1;
  wire v912634;
  wire v9125a8;
  wire v85c0ba;
  wire v86ff66;
  wire v8c520c;
  wire v8b0e17;
  wire v910c9d;
  wire v8af205;
  wire v8b038e;
  wire v8b1159;
  wire v912415;
  wire v9123bd;
  wire v8aebc5;
  wire v8b21e7;
  wire v8b3401;
  wire v890aa5;
  wire v912647;
  wire v9126e3;
  wire v8b04b6;
  wire v8afa71;
  wire v8b03fc;
  wire v911ed4;
  wire v8ae745;
  wire v8c0bb8;
  wire v91251d;
  wire v8b2cb5;
  wire v911795;
  wire v8aeeaa;
  wire v9124f3;
  wire v912730;
  wire v8c41ae;
  wire v8b08b3;
  wire v91272b;
  wire v8de9ca;
  wire v9121a4;
  wire v91204e;
  wire v8b2afc;
  wire v8dd5d6;
  wire v9113cc;
  wire v912444;
  wire v8afbaa;
  wire v911dbd;
  wire v912511;
  wire v9123ca;
  wire v910fe3;
  wire v8bfa6b;
  wire v8b0c14;
  wire v8c0a62;
  wire v8b02ce;
  wire v8b128f;
  wire v9123ec;
  wire v91249b;
  wire v8c52db;
  wire v8b0109;
  wire v88ee77;
  wire v8602f3;
  wire v911ed6;
  wire v8af318;
  wire v8b0c98;
  wire v8aebc4;
  wire v911704;
  wire v9118e7;
  wire v9125b3;
  wire v8b27a2;
  wire v8aebc8;
  wire v8b1f9c;
  wire v8b116b;
  wire v912678;
  wire v8afd22;
  wire v8ae0a2;
  wire v8b218f;
  wire v8aee08;
  wire v911fe2;
  wire v9125b4;
  wire v91246b;
  wire v8f96e9;
  wire v8c57f0;
  wire v9123f0;
  wire v911913;
  wire v911f4a;
  wire v8afe6f;
  wire v8cc22c;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg StoB_REQ4_p;
  input StoB_REQ4_n;
  reg StoB_REQ5_p;
  input StoB_REQ5_n;
  reg StoB_REQ6_p;
  input StoB_REQ6_n;
  reg StoB_REQ7_p;
  input StoB_REQ7_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoS_ACK4_p;
  output BtoS_ACK4_n;
  reg BtoS_ACK5_p;
  output BtoS_ACK5_n;
  reg BtoS_ACK6_p;
  output BtoS_ACK6_n;
  reg BtoS_ACK7_p;
  output BtoS_ACK7_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg SLC2_p;
  output SLC2_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  reg jx3_p;
  output jx3_n;
  wire ENQ_n;
  wire SLC0_n;
  wire SLC2_n;
  wire SLC1_n;

assign v8aeddc = StoB_REQ0_p & v911664 | !StoB_REQ0_p & v8b3286;
assign v8b22fd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af0e6;
assign v8d6cde = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b2a8f;
assign v8affb3 = StoB_REQ7_p & v8b0808 | !StoB_REQ7_p & v8b2c06;
assign v912764 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v91267c;
assign v8b1154 = StoB_REQ3_p & v8c44a1 | !StoB_REQ3_p & v8b2a3e;
assign v8b0acf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b2e72;
assign v9125a9 = RtoB_ACK1_p & v8909ff | !RtoB_ACK1_p & v844f91;
assign v8b2ae9 = BtoS_ACK7_p & v8af894 | !BtoS_ACK7_p & v9123ba;
assign v8b2885 = StoB_REQ7_p & v8af052 | !StoB_REQ7_p & v844f91;
assign v8b0cf7 = jx1_p & v8b2a8c | !jx1_p & v8c7100;
assign v890246 = StoB_REQ7_p & v8b2267 | !StoB_REQ7_p & v8b2088;
assign v8b109a = BtoR_REQ1_p & v8b0584 | !BtoR_REQ1_p & v9125af;
assign v8b03d4 = jx1_p & v8b2e60 | !jx1_p & v8b340b;
assign v9125da = BtoR_REQ1_p & v8ae7e5 | !BtoR_REQ1_p & v844f91;
assign v912542 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9113d6;
assign v892f3e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v912683;
assign v8afdec = jx3_p & v9110f5 | !jx3_p & !v8c4c96;
assign v87e29c = BtoS_ACK3_p & v8c050d | !BtoS_ACK3_p & v8c44a1;
assign v8c050d = StoB_REQ3_p & v8c44a1 | !StoB_REQ3_p & v844f9f;
assign v8aee85 = BtoS_ACK7_p & v911149 | !BtoS_ACK7_p & v8afa56;
assign v85e943 = BtoS_ACK1_p & v8ae516 | !BtoS_ACK1_p & v8b0a55;
assign v8ae878 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9123df;
assign v911ef0 = RtoB_ACK1_p & v8afde2 | !RtoB_ACK1_p & v890ac0;
assign v8b0260 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f95;
assign v844fad = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v8aea93 = RtoB_ACK0_p & v8c55bf | !RtoB_ACK0_p & v8b23d9;
assign v9114d3 = BtoR_REQ1_p & v8b05f1 | !BtoR_REQ1_p & v911441;
assign v85afd4 = BtoS_ACK3_p & v8c38b4 | !BtoS_ACK3_p & v91223a;
assign v8b0fe0 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & v8b06bb;
assign v8b0ce2 = ENQ_p & v8b2a8c | !ENQ_p & v9124a5;
assign v8dd6ae = jx0_p & v9126c9 | !jx0_p & v844f91;
assign v9124f5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8afa7c;
assign v912627 = BtoS_ACK4_p & v8b2252 | !BtoS_ACK4_p & v8afea6;
assign v9126f4 = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v8b0d78;
assign v8affe3 = BtoS_ACK6_p & v8b10fd | !BtoS_ACK6_p & v8ae06b;
assign v8af780 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v8b03e8;
assign v911eb5 = stateG7_1_p & v8b284f | !stateG7_1_p & v844f91;
assign v911c88 = BtoS_ACK3_p & v8b1fb5 | !BtoS_ACK3_p & v8b0762;
assign v8b0119 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8afe01;
assign v912074 = jx0_p & v8c4d16 | !jx0_p & !v87a52a;
assign v8b2420 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c55e1;
assign v8b21fa = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8bfa99;
assign v8c3926 = RtoB_ACK1_p & v890bcb | !RtoB_ACK1_p & v844f91;
assign v8b24e9 = BtoS_ACK6_p & v8af431 | !BtoS_ACK6_p & v912276;
assign v885339 = jx2_p & v8b21eb | !jx2_p & v8af02f;
assign v8c77e6 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8c537f;
assign v8c41af = BtoS_ACK7_p & v8b0661 | !BtoS_ACK7_p & v8b22fd;
assign v8ae461 = jx0_p & v8940eb | !jx0_p & v912691;
assign v85c126 = stateG7_1_p & v911bdc | !stateG7_1_p & v8c387f;
assign v8af563 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v912753;
assign v8b1014 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c59a9;
assign v91246d = StoB_REQ6_p & v912576 | !StoB_REQ6_p & v88b254;
assign v911c2f = StoB_REQ7_p & v8c3728 | !StoB_REQ7_p & v8b0264;
assign v8b0774 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8c3def;
assign v912785 = stateG7_1_p & v8afe84 | !stateG7_1_p & v9126dd;
assign v8f9587 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8afc68;
assign v8af478 = jx2_p & v8b0113 | !jx2_p & !v9123fe;
assign v8b0994 = jx2_p & v86990d | !jx2_p & v912461;
assign v863493 = EMPTY_p & v884a20 | !EMPTY_p & v8b2642;
assign v8afc92 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v91127a;
assign v8aeb97 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v87e29c;
assign v8b2345 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fedc9;
assign v844fb3 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v8dd687 = StoB_REQ4_p & v844f9f | !StoB_REQ4_p & !v844f91;
assign v911fbd = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v911eb5;
assign v8e5d84 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8d6d0f;
assign v890ac0 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e988e;
assign v8b1e80 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v912755;
assign v9126b0 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b140a;
assign v8fed5e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ae151;
assign v8afd4d = StoB_REQ2_p & v8b0283 | !StoB_REQ2_p & v8af864;
assign v8ae670 = RtoB_ACK1_p & v91257b | !RtoB_ACK1_p & v91134b;
assign v8b055a = BtoS_ACK6_p & v8ae578 | !BtoS_ACK6_p & v8b2aaa;
assign v91134b = jx2_p & v87dc9f | !jx2_p & v8aed2e;
assign v8af06b = jx1_p & v8b2e60 | !jx1_p & v91247e;
assign v8afcd6 = BtoS_ACK7_p & v8b0cbb | !BtoS_ACK7_p & v9116c2;
assign v912403 = BtoS_ACK1_p & v8c0b8f | !BtoS_ACK1_p & v8e990a;
assign v911b07 = BtoS_ACK6_p & v912432 | !BtoS_ACK6_p & v9124ea;
assign v912777 = jx2_p & v8b1166 | !jx2_p & !v8afaa7;
assign v8d6cda = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9110fb;
assign v8af811 = RtoB_ACK1_p & v8b28d5 | !RtoB_ACK1_p & !v844f91;
assign v892893 = DEQ_p & v8b0823 | !DEQ_p & v8ae162;
assign v91254f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8c0ab9;
assign v91259d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b1dbe;
assign v8afc88 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & v8b22f0;
assign v912690 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91273e;
assign v8b3d0e = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v890b4a;
assign v912716 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ae8d3;
assign v8c0456 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8b0934;
assign v8afedf = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8f956e;
assign v8c09e5 = BtoS_ACK0_p & v8b12af | !BtoS_ACK0_p & v8b2e70;
assign v8b29d8 = StoB_REQ2_p & v87e29c | !StoB_REQ2_p & v8aeb97;
assign v912481 = stateG7_1_p & v8b77ef | !stateG7_1_p & v8c66bb;
assign v8c6a96 = jx0_p & v912080 | !jx0_p & v8b2ae9;
assign v8b1195 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91263c;
assign v8d6d00 = BtoS_ACK0_p & v8d6d04 | !BtoS_ACK0_p & v8c6e2e;
assign v8ae7b3 = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & !v844f91;
assign v9126c8 = StoB_REQ6_p & v8b20ab | !StoB_REQ6_p & v912521;
assign v8b77f9 = StoB_REQ2_p & v912592 | !StoB_REQ2_p & v911fe3;
assign v8ae0b8 = jx1_p & v8b2180 | !jx1_p & v8ae12e;
assign v912166 = BtoS_ACK0_p & v8af918 | !BtoS_ACK0_p & v8aefce;
assign v8b3212 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8b2a92;
assign v8c7054 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v9112ad;
assign v8b297c = jx1_p & v8ae6f2 | !jx1_p & !v9124ce;
assign v8b09ce = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b3013;
assign v8dd6a6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8afe4c;
assign v9125f0 = StoB_REQ1_p & v9126f4 | !StoB_REQ1_p & v9125e6;
assign v8af214 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v9114ce;
assign v91268b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8b1de3;
assign v8b1fc9 = stateG7_1_p & v844f91 | !stateG7_1_p & !v9117c1;
assign v91268f = jx1_p & v8b2180 | !jx1_p & v911fa7;
assign v910e12 = StoB_REQ2_p & v8aec57 | !StoB_REQ2_p & !v912581;
assign v8b1cf2 = ENQ_p & v890ac0 | !ENQ_p & v8c23d1;
assign v8b7bb3 = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v9125b6;
assign v8b7804 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v844f99;
assign v8b113b = jx0_p & v9125f2 | !jx0_p & !v8bfa76;
assign v8b0500 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v912453;
assign v8fee03 = DEQ_p & v911ae3 | !DEQ_p & v8b2460;
assign v8b1ec4 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v8aee3c;
assign v911792 = BtoR_REQ1_p & v912409 | !BtoR_REQ1_p & v844f91;
assign v8ae768 = jx1_p & v9126eb | !jx1_p & v8aeb67;
assign v9119a4 = StoB_REQ7_p & v8aed74 | !StoB_REQ7_p & v911158;
assign v8fed7c = stateG7_1_p & v8c6dff | !stateG7_1_p & v9126d9;
assign v911411 = RtoB_ACK1_p & v8c66bb | !RtoB_ACK1_p & v844f91;
assign v8b04b6 = jx1_p & v9123bd | !jx1_p & !v9126e3;
assign v8c55e1 = StoB_REQ7_p & v9124f9 | !StoB_REQ7_p & v844f91;
assign v912797 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & !v912588;
assign v87b940 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8c3b8d;
assign v8b2ddd = StoB_REQ1_p & v8b293f | !StoB_REQ1_p & v844f91;
assign v911fdd = BtoS_ACK1_p & v844f9e | !BtoS_ACK1_p & v912745;
assign v8aef02 = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v844f9f;
assign v911b46 = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v8e989e;
assign v91260c = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8af765;
assign v9123bf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v91180a;
assign v8b099d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8bfa79;
assign v8c43e6 = StoB_REQ4_p & v8afea6 | !StoB_REQ4_p & !v844f91;
assign v8b10fd = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v844f91;
assign v8c6167 = BtoS_ACK1_p & v912557 | !BtoS_ACK1_p & v8b2868;
assign v8c71b3 = BtoS_ACK3_p & v8b2c21 | !BtoS_ACK3_p & v8c4ac3;
assign v8b0d89 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v912786;
assign v8b25a8 = stateG7_1_p & v8909ff | !stateG7_1_p & v8c4667;
assign v8fed90 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b06bb;
assign v8612be = StoB_REQ0_p & v9125cb | !StoB_REQ0_p & v844f91;
assign v8c3a0b = BtoS_ACK7_p & v911bad | !BtoS_ACK7_p & v87d0a9;
assign v8b2021 = jx1_p & v91277d | !jx1_p & v911fb6;
assign v911bf3 = jx2_p & v911714 | !jx2_p & !v8b257f;
assign v8b2073 = BtoS_ACK1_p & v911787 | !BtoS_ACK1_p & v9123a2;
assign v8b0446 = jx0_p & v86bf27 | !jx0_p & v8c6cd3;
assign v8ae69b = jx1_p & v8771a0 | !jx1_p & v8b7379;
assign v8b76c6 = BtoS_ACK6_p & v8c390a | !BtoS_ACK6_p & v8af193;
assign v8c6ccc = BtoS_ACK6_p & v8c6c4a | !BtoS_ACK6_p & v91256f;
assign v8ae14c = RtoB_ACK0_p & v87139e | !RtoB_ACK0_p & v8b0994;
assign v8b2c39 = jx0_p & v9125c5 | !jx0_p & v890ac0;
assign v8b085b = jx0_p & v8b246f | !jx0_p & v8ae562;
assign v873367 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912724;
assign v911219 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v8ae6ab;
assign v912394 = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v86cbb8;
assign v8b05ce = jx0_p & v912625 | !jx0_p & v8c3c57;
assign v910c73 = jx2_p & v8908a2 | !jx2_p & !v894826;
assign v8b1245 = jx3_p & v8e988e | !jx3_p & v890ac0;
assign v8cc182 = ENQ_p & v844fbb | !ENQ_p & !v887b47;
assign v911ff4 = BtoR_REQ0_p & v887b30 | !BtoR_REQ0_p & v912470;
assign v8ae160 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8c5058;
assign v8c52db = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91249b;
assign v8c09de = BtoS_ACK7_p & v911d4f | !BtoS_ACK7_p & v912291;
assign v8af1a2 = jx2_p & v8ae033 | !jx2_p & !v8c4cc3;
assign v8af4b1 = BtoS_ACK3_p & v91108c | !BtoS_ACK3_p & v912696;
assign v8f9659 = StoB_REQ3_p & v8b339d | !StoB_REQ3_p & v844f9d;
assign v8c3651 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8c4a56;
assign v8b2592 = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v8b0b9c;
assign v85c148 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8c043b;
assign BtoS_ACK7_n = v85c182;
assign v8c6d04 = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v910e98;
assign v9123c5 = jx1_p & v8b2180 | !jx1_p & v8fecb7;
assign v8ae83c = BtoS_ACK7_p & v912609 | !BtoS_ACK7_p & v9124e5;
assign v8b0764 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8b32c2;
assign v8b050c = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v8c426f;
assign v8c3bd5 = StoB_REQ2_p & v8af2f9 | !StoB_REQ2_p & !v91265a;
assign v8b02ed = BtoS_ACK0_p & v8b0df4 | !BtoS_ACK0_p & v890940;
assign v8c534d = BtoS_ACK6_p & v8af894 | !BtoS_ACK6_p & v8af0b0;
assign v8f956e = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9b;
assign v8aed2e = jx1_p & v912623 | !jx1_p & !v8b1068;
assign v8b094a = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8aebd0;
assign v8ae47c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af1d2;
assign v8b1f47 = StoB_REQ4_p & v912517 | !StoB_REQ4_p & v844f91;
assign v8591f3 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v912512;
assign v8c66bb = jx2_p & v8ae9c2 | !jx2_p & v844f91;
assign BtoS_ACK0_n = !v8db28c;
assign v9126d4 = jx1_p & v8aed7b | !jx1_p & v8c56de;
assign v8b1cd7 = BtoS_ACK0_p & v91244d | !BtoS_ACK0_p & v8b65a2;
assign v8b1e7d = BtoS_ACK7_p & v844f95 | !BtoS_ACK7_p & v8c6bfa;
assign v8b2b91 = jx0_p & v844f91 | !jx0_p & v8aed6d;
assign v8c64bf = BtoS_ACK7_p & v844fa1 | !BtoS_ACK7_p & v8c50c5;
assign v890aa5 = BtoS_ACK7_p & v8577c2 | !BtoS_ACK7_p & v8b3401;
assign v87f443 = jx1_p & v8771a0 | !jx1_p & v8ae9bf;
assign v9124ab = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85c16c;
assign v9125b2 = StoB_REQ6_p & v869876 | !StoB_REQ6_p & v844f91;
assign v85f3d2 = BtoR_REQ1_p & v85c126 | !BtoR_REQ1_p & v844f91;
assign v91264b = BtoR_REQ1_p & v8af34a | !BtoR_REQ1_p & v912102;
assign v8b0dd3 = jx3_p & v844f91 | !jx3_p & !v8aeb12;
assign v9111d2 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c43c1;
assign v912466 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8b0681;
assign v8aeb29 = StoB_REQ1_p & v8b0fa3 | !StoB_REQ1_p & v8ae789;
assign v8b0219 = StoB_REQ2_p & v8ae0ee | !StoB_REQ2_p & v8af9bd;
assign v8b2e70 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9123c6;
assign v8cc129 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8afaec;
assign v8aeabf = stateG7_1_p & v8afa41 | !stateG7_1_p & v8af1ef;
assign v91272d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844fb3;
assign v911ed4 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8b03fc;
assign v912581 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8aec57;
assign v8b1d6c = jx1_p & v844f91 | !jx1_p & !v869205;
assign v912501 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v911959;
assign v8e9920 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v9119da;
assign v8b2657 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v9124de;
assign v9114cd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91268a;
assign v8c723e = jx2_p & v91242c | !jx2_p & !v86bd18;
assign v8c7247 = BtoR_REQ0_p & v8db195 | !BtoR_REQ0_p & v8bfa98;
assign v8c5239 = jx3_p & v844f91 | !jx3_p & v8c3c40;
assign v912722 = jx1_p & v8c3a82 | !jx1_p & !v9125b9;
assign v8b1248 = BtoS_ACK3_p & v8ae4cd | !BtoS_ACK3_p & !v8af3eb;
assign v88ed6a = BtoS_ACK6_p & v8af431 | !BtoS_ACK6_p & v8b2fc3;
assign v890534 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b0c67;
assign v8aebc5 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v9126f5;
assign v87139e = jx2_p & v912722 | !jx2_p & v8b0b24;
assign v8b76f4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8aeecd;
assign v9116ad = StoB_REQ6_p & v9116e8 | !StoB_REQ6_p & v8b4fda;
assign v9123aa = BtoS_ACK1_p & v8b229e | !BtoS_ACK1_p & v8af5fe;
assign v9124ff = BtoS_ACK6_p & v8ae578 | !BtoS_ACK6_p & v890c50;
assign v912635 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v911c80;
assign v8c7263 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af780;
assign v911631 = jx2_p & v9123c5 | !jx2_p & v8af8b0;
assign v8af7b2 = BtoS_ACK3_p & v8b33a8 | !BtoS_ACK3_p & v8fed90;
assign v8c3027 = BtoS_ACK7_p & v911149 | !BtoS_ACK7_p & v8839ea;
assign v8b076a = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v885d39;
assign v912561 = RtoB_ACK1_p & v885339 | !RtoB_ACK1_p & v8af02f;
assign v8c65f8 = jx0_p & v892501 | !jx0_p & !v8b25a2;
assign v8afab8 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91259d;
assign v91177e = BtoS_ACK0_p & v879d5b | !BtoS_ACK0_p & v8aeabb;
assign v91157e = StoB_REQ1_p & v890b4a | !StoB_REQ1_p & v844f91;
assign v912746 = stateG7_1_p & v8c66bb | !stateG7_1_p & v8b22c1;
assign v912448 = jx0_p & v912471 | !jx0_p & !v844f99;
assign v8b0485 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v844fa3;
assign v8b004e = BtoR_REQ1_p & v887acc | !BtoR_REQ1_p & v8b0e8e;
assign v91247e = jx0_p & v8b021d | !jx0_p & v9126b0;
assign v912181 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8aeeeb;
assign v8ae582 = RtoB_ACK1_p & v9115b8 | !RtoB_ACK1_p & v912201;
assign v8c426e = BtoS_ACK7_p & v911bad | !BtoS_ACK7_p & v8c37c9;
assign v8b28e6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b0283;
assign v8b2f6b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b1a14;
assign v8b1fb5 = StoB_REQ3_p & v8b0762 | !StoB_REQ3_p & !v844f9f;
assign v911fac = jx2_p & v9126d8 | !jx2_p & v8afe97;
assign v88b254 = BtoS_ACK0_p & v8c0b8f | !BtoS_ACK0_p & v912464;
assign v8b28fe = StoB_REQ2_p & v8b6482 | !StoB_REQ2_p & v8af23b;
assign v911fd5 = EMPTY_p & v8c702a | !EMPTY_p & v9110fc;
assign v91100c = jx1_p & v8771a0 | !jx1_p & v8b26ee;
assign v8e9884 = StoB_REQ7_p & v8db203 | !StoB_REQ7_p & v8af004;
assign v912660 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v89098c;
assign v8809fb = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8c36bc;
assign v8b051c = RtoB_ACK1_p & v9124a9 | !RtoB_ACK1_p & v88acc3;
assign v8618ff = RtoB_ACK0_p & v8b0a78 | !RtoB_ACK0_p & v844f91;
assign v912280 = EMPTY_p & v8b2741 | !EMPTY_p & v9119bc;
assign v9123d3 = StoB_REQ6_p & v911ad5 | !StoB_REQ6_p & v8b131b;
assign v912664 = jx2_p & v8b082d | !jx2_p & !v8c4cc3;
assign v8af410 = jx3_p & v844f91 | !jx3_p & v8b222c;
assign v8afc39 = stateG7_1_p & v8ae588 | !stateG7_1_p & v8618ff;
assign v91108c = StoB_REQ3_p & v8c381a | !StoB_REQ3_p & v844f9f;
assign v9125c8 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9124dd;
assign v8ae4b3 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844fa3;
assign v911ee4 = jx1_p & v911382 | !jx1_p & v912401;
assign v91118f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9125a0;
assign v912515 = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v9123cc;
assign v911664 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b139e;
assign v9115c7 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0494;
assign v912780 = BtoS_ACK6_p & v8b327a | !BtoS_ACK6_p & v8c0bf1;
assign v8b26ee = jx0_p & v912626 | !jx0_p & !v8c0b7c;
assign v8b22a7 = StoB_REQ2_p & v8aefe5 | !StoB_REQ2_p & v8ae825;
assign v911196 = jx2_p & v8c5d7e | !jx2_p & v8ae5c6;
assign v8b24b0 = jx0_p & v8dd6bd | !jx0_p & !v8b1e7d;
assign v8b65a2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b1dfe;
assign v890880 = BtoR_REQ0_p & v8af2e0 | !BtoR_REQ0_p & v8afa40;
assign v85ed5d = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v8aec57;
assign v8b76c0 = jx0_p & v911fda | !jx0_p & !v890c2c;
assign v912549 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v91240c;
assign v8af9e8 = BtoS_ACK3_p & v8b0e4c | !BtoS_ACK3_p & !v844f91;
assign v8fecd9 = BtoS_ACK7_p & v8b2eed | !BtoS_ACK7_p & v912591;
assign v8c3cff = jx2_p & v91275f | !jx2_p & v8b23d4;
assign v8fed23 = BtoS_ACK6_p & v8b33d3 | !BtoS_ACK6_p & !v8ae6ab;
assign v8b2812 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & !v8af159;
assign v8c6bba = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & v8c5fa2;
assign v8b26cf = BtoS_ACK1_p & v879d5b | !BtoS_ACK1_p & v9124d5;
assign v8b0109 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v911197;
assign v8b062d = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c7263;
assign v8b0a17 = BtoR_REQ0_p & v8b01f5 | !BtoR_REQ0_p & v911ed2;
assign v912508 = jx3_p & v844f91 | !jx3_p & v9126f0;
assign v8c0443 = BtoS_ACK0_p & v8d6d04 | !BtoS_ACK0_p & v910efa;
assign v8b0e9d = jx3_p & v844f91 | !jx3_p & v8b0750;
assign v887b53 = jx2_p & v912658 | !jx2_p & v912742;
assign v8c5e9b = BtoS_ACK6_p & v9126de | !BtoS_ACK6_p & v9112aa;
assign v8af094 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8af7a3;
assign v8af1e9 = BtoR_REQ0_p & v8aee79 | !BtoR_REQ0_p & v8ae7de;
assign v8af2f5 = StoB_REQ1_p & v87b5cf | !StoB_REQ1_p & v8af9ff;
assign v8b2a8f = BtoS_ACK0_p & v9123df | !BtoS_ACK0_p & v912669;
assign v8c704a = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8b2b17;
assign v911742 = BtoS_ACK1_p & v8b034f | !BtoS_ACK1_p & v8b2275;
assign v8b33f2 = BtoR_REQ0_p & v9126d2 | !BtoR_REQ0_p & v8b76f3;
assign v9124c4 = jx0_p & v8af82e | !jx0_p & v8b1e7d;
assign v890b35 = jx0_p & v8c0b04 | !jx0_p & v911633;
assign v8afc68 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & !v9125b1;
assign v887c34 = StoB_REQ6_p & v8b3d12 | !StoB_REQ6_p & v911d7e;
assign v8c3617 = BtoR_REQ0_p & v8c57d1 | !BtoR_REQ0_p & v8b0936;
assign v912680 = BtoR_REQ0_p & v8b09b9 | !BtoR_REQ0_p & v8c043d;
assign v8b0dc4 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8c6e5a;
assign v911e9b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91272d;
assign v8b1f2d = jx0_p & v90c2e3 | !jx0_p & !v911c25;
assign v8af5b7 = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v9124f6;
assign v8b08ac = StoB_REQ1_p & v8ae722 | !StoB_REQ1_p & v844f91;
assign v8af916 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844fa1;
assign v8bfa5d = StoB_REQ6_p & v8b261e | !StoB_REQ6_p & v912514;
assign v8b33a8 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8aef02;
assign v8c369a = RtoB_ACK1_p & v910947 | !RtoB_ACK1_p & v8b2688;
assign v9125d3 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86b11f;
assign v8b0223 = BtoS_ACK6_p & v8c6c4a | !BtoS_ACK6_p & v8bfa5d;
assign v911765 = jx2_p & v8ae033 | !jx2_p & !v8af2cd;
assign v8b134f = RtoB_ACK1_p & v85f4b2 | !RtoB_ACK1_p & v8b02e9;
assign v91272e = jx0_p & v912563 | !jx0_p & v844f91;
assign v8c0a9d = BtoS_ACK7_p & v912702 | !BtoS_ACK7_p & v87bd82;
assign v8afce6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b08ac;
assign v8b3383 = jx0_p & v8ae8bf | !jx0_p & !v8c4569;
assign v845125 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88ed6a;
assign v912593 = StoB_REQ7_p & v9123ba | !StoB_REQ7_p & v85a510;
assign v8b282e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v9124fe;
assign v9126df = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v861f8d;
assign v8b2197 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9114e5;
assign v85c0b1 = BtoS_ACK0_p & v8f9617 | !BtoS_ACK0_p & v8b2d82;
assign v8c4b39 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v91257f;
assign v912527 = StoB_REQ6_p & v8809fb | !StoB_REQ6_p & v8b0653;
assign v912649 = jx2_p & v912650 | !jx2_p & v89409b;
assign v9124c2 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b00fe;
assign v8c5192 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v9122d7;
assign v8b265b = stateG7_1_p & v9115b8 | !stateG7_1_p & v911173;
assign v9114e1 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c5d1b;
assign v912753 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b08fa;
assign v8bb97f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0626;
assign v8b2ca9 = jx0_p & v8b21a3 | !jx0_p & !v8b1e7d;
assign v8b233e = BtoS_ACK7_p & v8ae878 | !BtoS_ACK7_p & v8b0449;
assign v9112e0 = StoB_REQ3_p & v910e18 | !StoB_REQ3_p & v844fb5;
assign v8afa7c = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v9125df;
assign v9125e5 = BtoR_REQ0_p & v91157d | !BtoR_REQ0_p & v85f776;
assign v8cc220 = jx0_p & v8c3027 | !jx0_p & v844f91;
assign v8c715a = StoB_REQ7_p & v844f9f | !StoB_REQ7_p & v844f91;
assign v8c3af9 = jx1_p & v887bdb | !jx1_p & v8af410;
assign v91250c = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v912493;
assign v91130e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b2c79;
assign v8c3e35 = jx3_p & v844f91 | !jx3_p & !v8afd55;
assign v8aea72 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v875f27;
assign v8aed37 = jx1_p & v8ae6f2 | !jx1_p & !v8c3afa;
assign v91243f = jx0_p & v8c5192 | !jx0_p & !v8c5d1c;
assign v8b2fc8 = jx1_p & v8b2e60 | !jx1_p & v8b068c;
assign v8b2843 = BtoS_ACK6_p & v8af431 | !BtoS_ACK6_p & v912428;
assign v8b039c = stateG7_1_p & v844f91 | !stateG7_1_p & !v844fa5;
assign v8b3d09 = BtoS_ACK7_p & v8bfa8b | !BtoS_ACK7_p & v871abf;
assign v8ae033 = jx1_p & v8b320b | !jx1_p & v890b35;
assign v8fece4 = StoB_REQ3_p & v8b0762 | !StoB_REQ3_p & !v8b2a3e;
assign v912451 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v89092e;
assign v9126dd = RtoB_ACK0_p & v8b28d4 | !RtoB_ACK0_p & v8afe84;
assign v8c0433 = ENQ_p & v87d0f8 | !ENQ_p & v863493;
assign v91251b = StoB_REQ1_p & v881ef0 | !StoB_REQ1_p & v910c58;
assign v8b2633 = ENQ_p & v8c0aba | !ENQ_p & v8b276b;
assign v8b2a92 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8b2a3e;
assign v8af6d0 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v910e18;
assign v8f9632 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v8ae5a8;
assign v91256f = StoB_REQ6_p & v8c5058 | !StoB_REQ6_p & v8c0ae6;
assign v9110fb = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v890930;
assign v912651 = StoB_REQ6_p & v8af334 | !StoB_REQ6_p & v844f91;
assign v8b0642 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8aec46;
assign v8c537f = BtoS_ACK3_p & v91108c | !BtoS_ACK3_p & v8c381a;
assign v8b03cf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v91244d;
assign v9112b6 = BtoS_ACK6_p & v912609 | !BtoS_ACK6_p & v8b2220;
assign v8dd691 = jx1_p & v8b032e | !jx1_p & v844f91;
assign v9126e7 = StoB_REQ7_p & v9125d8 | !StoB_REQ7_p & v8b0d9e;
assign v892e12 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b2815;
assign v861315 = StoB_REQ0_p & v911664 | !StoB_REQ0_p & v892e44;
assign v9125df = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b0436;
assign v8b1d42 = StoB_REQ7_p & v91276d | !StoB_REQ7_p & v8940ac;
assign v8f9614 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b2a3e;
assign v8ae756 = jx0_p & v912790 | !jx0_p & v844f91;
assign v8b1129 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8afb9b;
assign v8b2553 = StoB_REQ0_p & v8b1a14 | !StoB_REQ0_p & v844f91;
assign v8ae8e3 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8af98a;
assign v91245a = BtoS_ACK6_p & v8b10fd | !BtoS_ACK6_p & v9123a8;
assign v91183d = BtoS_ACK7_p & v8b2019 | !BtoS_ACK7_p & v910d59;
assign v8b08b3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c41ae;
assign v8af0b5 = stateG7_1_p & v8b12ad | !stateG7_1_p & !v8b76f2;
assign v91271d = jx0_p & v844f91 | !jx0_p & v9110f5;
assign v912616 = BtoS_ACK1_p & v8afd76 | !BtoS_ACK1_p & v8aedb1;
assign v8b2df5 = RtoB_ACK1_p & v9124db | !RtoB_ACK1_p & v844f91;
assign v8b0681 = jx2_p & v863839 | !jx2_p & v844f91;
assign v8c0b8f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8aef7a;
assign v9124a9 = jx2_p & v8af2b1 | !jx2_p & v88acc3;
assign v8b21bb = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9123e6;
assign v9126a8 = BtoS_ACK3_p & v9110d2 | !BtoS_ACK3_p & v844fb5;
assign v91257a = jx1_p & v9123ff | !jx1_p & !v8b2c4c;
assign v86f676 = ENQ_p & v890a25 | !ENQ_p & !v912777;
assign v8c044b = jx1_p & v8771a0 | !jx1_p & v8b76c0;
assign v8c049e = jx3_p & v8ae4b3 | !jx3_p & v882fb4;
assign v911797 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b11a0;
assign v8afea6 = StoB_REQ5_p & v844fb7 | !StoB_REQ5_p & v844f91;
assign v912331 = jx1_p & v8ae6f0 | !jx1_p & v89287e;
assign v87cf74 = StoB_REQ6_p & v89092e | !StoB_REQ6_p & v8b1014;
assign v9123ee = BtoR_REQ0_p & v844fbb | !BtoR_REQ0_p & v912550;
assign v8b2fd3 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8af452;
assign v912792 = StoB_REQ6_p & v8b0674 | !StoB_REQ6_p & v85c0b1;
assign v8b28d4 = jx2_p & v8b297c | !jx2_p & v8aed2e;
assign v867e4e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c39e2;
assign v8ae64a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b0fa3;
assign v8b257f = jx1_p & v8b2df3 | !jx1_p & v8b1c7b;
assign v8b0a55 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b07c0;
assign v8c4a94 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8c51e1;
assign v8b0d2f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v910c25;
assign v8ae93f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911fd2;
assign v8afe4c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v911787;
assign v8afe97 = jx1_p & v8c6caf | !jx1_p & v912508;
assign v8b2878 = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v9114a2;
assign v8af687 = stateG7_1_p & v8b02e9 | !stateG7_1_p & v87b84a;
assign v8b2353 = StoB_REQ2_p & v844fb1 | !StoB_REQ2_p & !v844f91;
assign v8b238a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ae64a;
assign v912771 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v88e0ec;
assign v8b2d5a = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v912768;
assign v8ae578 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8dd65f;
assign v911f8b = BtoR_REQ0_p & v8b02dd | !BtoR_REQ0_p & v8b1e9a;
assign v8af240 = jx1_p & v8b2a71 | !jx1_p & v8afb09;
assign v9125b1 = StoB_REQ2_p & v911c88 | !StoB_REQ2_p & !v8b8e74;
assign v911174 = RtoB_ACK1_p & v8ae0da | !RtoB_ACK1_p & v910db7;
assign v8c0a23 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v9123df;
assign v86b11f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8ae07b;
assign v8c44a1 = BtoS_ACK4_p & v9123af | !BtoS_ACK4_p & v912517;
assign v8b2088 = BtoS_ACK6_p & v911d4f | !BtoS_ACK6_p & v912558;
assign v9121d1 = stateG12_p & v9112bc | !stateG12_p & v9126d5;
assign v8909b7 = BtoS_ACK3_p & v8b33a8 | !BtoS_ACK3_p & v911a56;
assign v912623 = jx0_p & v911fd9 | !jx0_p & v844f91;
assign v892fa2 = jx1_p & v8c3a82 | !jx1_p & !v8c46bf;
assign v8afe49 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8db1b0;
assign v911cf2 = jx0_p & v912668 | !jx0_p & v91258f;
assign v8afcaa = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8b2a7e;
assign v9124e1 = jx3_p & v844f91 | !jx3_p & !v9124c4;
assign v8b244a = jx3_p & v844f91 | !jx3_p & v8b2ca9;
assign v8b0e72 = jx0_p & v912790 | !jx0_p & v912666;
assign v8dd637 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b0599;
assign v912557 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9d;
assign v9125bc = BtoS_ACK0_p & v8b7892 | !BtoS_ACK0_p & v88704a;
assign v8b25f9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9123bf;
assign v8c420b = RtoB_ACK1_p & v911e3b | !RtoB_ACK1_p & v91194c;
assign v8b2080 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v9125f8;
assign v871da5 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b0a55;
assign v9123b6 = jx0_p & v8fec67 | !jx0_p & v8af71d;
assign v8b1dfe = BtoS_ACK1_p & v8b034f | !BtoS_ACK1_p & v9125d3;
assign v8940d8 = BtoS_ACK7_p & v88b300 | !BtoS_ACK7_p & v8c7385;
assign v8b1a14 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b7794;
assign v887b94 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8aec34;
assign v9125e2 = StoB_REQ6_p & v8b4c61 | !StoB_REQ6_p & v844f91;
assign v8bfa65 = jx0_p & v91271b | !jx0_p & v844f91;
assign v8b2afc = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91204e;
assign v912465 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8af634;
assign v8b2aaa = StoB_REQ6_p & v8af72b | !StoB_REQ6_p & v8b131b;
assign v8b77ed = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b2929;
assign v86ff66 = BtoS_ACK7_p & v8b1ff8 | !BtoS_ACK7_p & v85c0ba;
assign v8ae713 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v912283;
assign v887acc = stateG7_1_p & v844fa7 | !stateG7_1_p & !v844f91;
assign v8ae6e2 = stateG7_1_p & v8b2a63 | !stateG7_1_p & v912466;
assign v91253b = RtoB_ACK1_p & v910884 | !RtoB_ACK1_p & v8c66bb;
assign v8b2f46 = jx1_p & v8ae6f2 | !jx1_p & !v8b3402;
assign v8b1e0b = RtoB_ACK0_p & v8ae909 | !RtoB_ACK0_p & v8cf811;
assign v8b2cf0 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & !v8b3357;
assign v8af7a3 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8b33fa;
assign v9123de = stateG7_1_p & v8aecbf | !stateG7_1_p & v8b2fbc;
assign v8aeb4c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8afaa6;
assign v8af275 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v911fbe;
assign v8afaed = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8aec57;
assign v912102 = stateG7_1_p & v8aea76 | !stateG7_1_p & v890ac0;
assign v9123b1 = jx2_p & v8af06b | !jx2_p & v8c498b;
assign v912505 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b1dbd;
assign v8cc104 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8689df;
assign v9125d4 = BtoS_ACK7_p & v8577c2 | !BtoS_ACK7_p & v8af26f;
assign v8c6c2f = RtoB_ACK1_p & v8ae696 | !RtoB_ACK1_p & v8b03c8;
assign v8b22c1 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8c66bb;
assign v8b1fe8 = StoB_REQ1_p & v912523 | !StoB_REQ1_p & v8b1c70;
assign v91263d = jx1_p & v8771a0 | !jx1_p & v8940af;
assign v8b0211 = BtoS_ACK1_p & v911787 | !BtoS_ACK1_p & v8b0f67;
assign v91269d = BtoS_ACK7_p & v912702 | !BtoS_ACK7_p & v8afd2b;
assign v8b6d87 = BtoS_ACK1_p & v8b07c0 | !BtoS_ACK1_p & v8b0a55;
assign v8b2e31 = BtoR_REQ0_p & v91255f | !BtoR_REQ0_p & v910ea7;
assign v8c23c8 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & !v8b2f95;
assign v8b52f8 = StoB_REQ2_p & v8b263d | !StoB_REQ2_p & v8f956e;
assign v8db288 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v9126ad;
assign v8b33ed = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v8b09e5;
assign v912472 = stateG7_1_p & v887ac4 | !stateG7_1_p & v8af2c8;
assign v8b1d83 = RtoB_ACK0_p & v9123b1 | !RtoB_ACK0_p & v890bcb;
assign v910ea7 = BtoR_REQ1_p & v8cfeeb | !BtoR_REQ1_p & v8ae934;
assign v87cf71 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8aea9f;
assign v8b7794 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v8afaa7 = jx1_p & v912623 | !jx1_p & v844f91;
assign v912589 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v8b1086;
assign v8b327a = StoB_REQ4_n & v844f91 | !StoB_REQ4_n & v844fa0;
assign v8fed36 = EMPTY_p & v8af7c1 | !EMPTY_p & v912777;
assign v8aff75 = jx1_p & v8b8bdf | !jx1_p & v8b2f4e;
assign v912683 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v91215f;
assign v8c6c7e = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8af451;
assign v911cec = RtoB_ACK0_p & v8ae4ce | !RtoB_ACK0_p & v844f91;
assign v8b9047 = ENQ_p & v912154 | !ENQ_p & v8b0dd9;
assign v8b33af = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v887ae1;
assign v8b1f0a = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8af052;
assign v8d6d0f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v911fd6;
assign v8b2688 = jx2_p & v8ae768 | !jx2_p & v8af886;
assign v9123ad = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8afb06;
assign v9126e1 = FULL_p & v8c7247 | !FULL_p & v8af253;
assign v8b0112 = jx0_p & v8b26bb | !jx0_p & v8b0eea;
assign v8b1ff8 = StoB_REQ6_p & v864227 | !StoB_REQ6_p & v911a6a;
assign v8c6cd3 = BtoS_ACK7_p & v9126de | !BtoS_ACK7_p & v8b1385;
assign v912745 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v9126c4;
assign v911e1d = BtoR_REQ1_p & v8b2ba6 | !BtoR_REQ1_p & v844f91;
assign v8b0283 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8af6d0;
assign v8ae7de = BtoR_REQ1_p & v8b265b | !BtoR_REQ1_p & v8c5781;
assign v8db22c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v911fb3;
assign v9125a5 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v8d6cde;
assign v8b236d = jx1_p & v8b2bee | !jx1_p & !v887b1c;
assign v8b3320 = BtoS_ACK6_p & v912432 | !BtoS_ACK6_p & v8b1410;
assign v8b1ec0 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8aea07;
assign v8b1199 = BtoS_ACK6_p & v864227 | !BtoS_ACK6_p & v912766;
assign v8940ac = BtoS_ACK6_p & v91222a | !BtoS_ACK6_p & v872c7c;
assign v8c43c1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8af5bd;
assign v8feced = StoB_REQ1_p & v8afe22 | !StoB_REQ1_p & v844f91;
assign v910c58 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8db139;
assign v91259a = StoB_REQ2_p & v8b1ea2 | !StoB_REQ2_p & v8b210b;
assign v8cc22c = DEQ_p & v8b0ce2 | !DEQ_p & v8afe6f;
assign v91270b = StoB_REQ1_p & v87d059 | !StoB_REQ1_p & v844f91;
assign v8c56de = jx0_p & v8af52b | !jx0_p & !v8bfa76;
assign v911f54 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8b02a9;
assign v9123f8 = StoB_REQ0_p & v912453 | !StoB_REQ0_p & v91246a;
assign v9126f7 = BtoS_ACK0_p & v8b0df4 | !BtoS_ACK0_p & v8dd5ca;
assign v8b0a03 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b2aeb;
assign v911d2c = jx1_p & v8ae6f2 | !jx1_p & !v8cc220;
assign v8b6d3d = StoB_REQ2_p & v8c537f | !StoB_REQ2_p & v8c77e6;
assign v912425 = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v9124f5;
assign v8b340b = jx0_p & v91243d | !jx0_p & v8c4d14;
assign v91257f = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844fb5;
assign v8b6482 = BtoS_ACK3_p & v912763 | !BtoS_ACK3_p & v9124ed;
assign v8b00fe = StoB_REQ7_p & v911c7e | !StoB_REQ7_p & v8b236f;
assign v8ae936 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8bfae8;
assign v859212 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8dd5cf;
assign v890ab8 = BtoR_REQ0_p & v8ae6e2 | !BtoR_REQ0_p & v8b109a;
assign v8c6e8e = jx1_p & v912685 | !jx1_p & v8c049e;
assign v912431 = stateG7_1_p & v8b0994 | !stateG7_1_p & v8dd6fe;
assign v88ac88 = stateG7_1_p & v844f91 | !stateG7_1_p & v8b1ddf;
assign v8ae9c2 = jx1_p & v912554 | !jx1_p & v844f91;
assign v8c0429 = BtoS_ACK6_p & v8c5845 | !BtoS_ACK6_p & v89342c;
assign v91274b = BtoS_ACK3_p & v91251a | !BtoS_ACK3_p & v8b339d;
assign v8af2ab = jx1_p & v8b016d | !jx1_p & !v9124e1;
assign v8b07ff = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v8b0d58;
assign v8b0496 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v844f91;
assign v8c5c8c = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v890ac7;
assign v91151f = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v912657;
assign v911913 = FULL_p & v8ae0a2 | !FULL_p & v9123f0;
assign v9124bd = StoB_REQ3_p & v8aecf5 | !StoB_REQ3_p & v844f91;
assign v8b076f = StoB_REQ7_p & v9122d7 | !StoB_REQ7_p & v91260c;
assign v8dd5d8 = StoB_REQ7_p & v912451 | !StoB_REQ7_p & v8af1d7;
assign v8c4740 = RtoB_ACK0_p & v91176c | !RtoB_ACK0_p & v8af1a2;
assign v9126c2 = StoB_REQ7_p & v844fad | !StoB_REQ7_p & !v8e988e;
assign v91261f = StoB_REQ0_p & v91277b | !StoB_REQ0_p & v912616;
assign v8b29c1 = BtoR_REQ1_p & v910c72 | !BtoR_REQ1_p & v8afc39;
assign v8827a3 = StoB_REQ0_p & v91219b | !StoB_REQ0_p & v844f91;
assign v91242d = BtoS_ACK7_p & v911149 | !BtoS_ACK7_p & v8aed35;
assign v911a2a = jx0_p & v8b1d71 | !jx0_p & v844f91;
assign v8b2d68 = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v911e94;
assign v8b2220 = BtoS_ACK0_p & v8d6d04 | !BtoS_ACK0_p & v8af340;
assign v8aedc6 = BtoR_REQ1_p & v8af34a | !BtoR_REQ1_p & v890ac0;
assign v91265c = jx0_p & v9123dd | !jx0_p & v9110f5;
assign v8b068b = jx3_p & v8b016c | !jx3_p & v8c3c40;
assign v88abf5 = stateG12_p & v8894e7 | !stateG12_p & v8b2792;
assign v8c4a25 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0633;
assign v8b13ca = jx2_p & v911ee4 | !jx2_p & v911e0c;
assign v8b2b2d = BtoS_ACK6_p & v8af4ee | !BtoS_ACK6_p & v8b2c5d;
assign v888464 = StoB_REQ2_p & v8bfae8 | !StoB_REQ2_p & v8ae936;
assign v9123ce = jx1_p & v8b29e2 | !jx1_p & v8b113b;
assign v9123ec = stateG7_1_p & v844f91 | !stateG7_1_p & v8b128f;
assign v8af9ff = StoB_REQ2_p & v8ae0ee | !StoB_REQ2_p & v912565;
assign v8c4189 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912739;
assign v8af8f5 = RtoB_ACK1_p & v912698 | !RtoB_ACK1_p & v8ae81f;
assign v8afa8e = jx1_p & v8b0112 | !jx1_p & !v8f9631;
assign v8bfa4c = stateG7_1_p & v88acc3 | !stateG7_1_p & v9124cf;
assign v912578 = RtoB_ACK0_p & v8c66bb | !RtoB_ACK0_p & v844f91;
assign v8fed12 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b29d8;
assign v8b28a7 = StoB_REQ0_p & v8b0f42 | !StoB_REQ0_p & v844f91;
assign v911ae3 = ENQ_p & v88acc3 | !ENQ_p & v9124d8;
assign v9124c9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8b2f95;
assign v8b0753 = BtoS_ACK6_p & v8af4ee | !BtoS_ACK6_p & v91245f;
assign v8b7379 = jx0_p & v8ae7c9 | !jx0_p & !v890c2c;
assign v8af2cd = jx1_p & v8ae51a | !jx1_p & !v8b0cfd;
assign v8b09a3 = stateG7_1_p & v9112d7 | !stateG7_1_p & v8b2a8c;
assign v8b2a5b = BtoS_ACK6_p & v911d4f | !BtoS_ACK6_p & v8b2e92;
assign v8bfa6b = BtoR_REQ1_p & v910fe3 | !BtoR_REQ1_p & v844f91;
assign v910ff6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v9125bc;
assign v8c3c57 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v910d59;
assign v8d14b5 = stateG7_1_p & v91153e | !stateG7_1_p & v8af84d;
assign v890a73 = jx0_p & v911de3 | !jx0_p & !v8b1e7d;
assign v912201 = jx2_p & v9115b8 | !jx2_p & v8b085a;
assign v8b20fa = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v870559;
assign v8b2c07 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v912513;
assign v8ae83f = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v844f91;
assign v9124de = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v911917;
assign v8b0f51 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v911978;
assign v911fb3 = StoB_REQ7_p & v8b1ddc | !StoB_REQ7_p & v8affe3;
assign v911aa3 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v87b54c;
assign v8b2fc4 = BtoS_ACK2_p & v88709f | !BtoS_ACK2_p & v8bfab7;
assign v8b27f9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b12af;
assign v8b2c68 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8b330f;
assign v8ae765 = jx0_p & v8c4a25 | !jx0_p & v8af3b2;
assign v8ae516 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9d;
assign v8b0c90 = stateG7_1_p & v8b2a8c | !stateG7_1_p & v912417;
assign v911fd1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91188e;
assign v8b2e17 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v911a5d;
assign v8b0d4e = RtoB_ACK1_p & v8b23d9 | !RtoB_ACK1_p & v844f91;
assign v91211a = BtoS_ACK6_p & v8c426f | !BtoS_ACK6_p & v8c47bf;
assign v8bfa98 = BtoR_REQ1_p & v9123a4 | !BtoR_REQ1_p & v8afc39;
assign v8e98d2 = EMPTY_p & v8b2464 | !EMPTY_p & v9121d1;
assign v8e9859 = stateG7_1_p & v8b12b1 | !stateG7_1_p & v912698;
assign v8af382 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v8b2d4a;
assign v9124f2 = RtoB_ACK0_p & v8b01bd | !RtoB_ACK0_p & v844f91;
assign v9124d6 = jx2_p & v9124d7 | !jx2_p & v910bd1;
assign v9123c9 = StoB_REQ0_p & v8ae46d | !StoB_REQ0_p & v844f91;
assign v8b22ef = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v8db139;
assign v8aee6c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b251f;
assign v912511 = jx1_p & v8b320b | !jx1_p & v911dbd;
assign v8b0d32 = StoB_REQ1_p & v8b29d8 | !StoB_REQ1_p & v8b2f6c;
assign v8af85c = StoB_REQ3_p & v8b2b08 | !StoB_REQ3_p & v844f9f;
assign v8aec46 = BtoS_ACK6_p & v911bad | !BtoS_ACK6_p & v8c5e54;
assign v8c0508 = BtoS_ACK2_p & v8ae516 | !BtoS_ACK2_p & v8714a5;
assign v8c39e1 = FULL_p & v8b74aa | !FULL_p & v8c3617;
assign v911733 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8b0b70;
assign v8c6cee = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v844f91;
assign v91255f = stateG7_1_p & v8b2d73 | !stateG7_1_p & v89097f;
assign v85c157 = StoB_REQ0_p & v8b12f9 | !StoB_REQ0_p & v91264a;
assign v88e856 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b0acf;
assign v8bfa61 = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v8b02a9;
assign v9124b7 = StoB_REQ7_p & v8af3b6 | !StoB_REQ7_p & v8c4a94;
assign v871abf = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c5350;
assign v892511 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8b0df4;
assign v9123e6 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v8b2ad6;
assign v8b2935 = StoB_REQ1_p & v8c4b39 | !StoB_REQ1_p & v884789;
assign v8b336e = jx1_p & v911be0 | !jx1_p & !v912644;
assign v9125d7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8db217;
assign v8aea76 = RtoB_ACK1_p & v890ac0 | !RtoB_ACK1_p & v9123c4;
assign v8ae8e8 = jx0_p & v8b8e79 | !jx0_p & v888766;
assign v912462 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9123aa;
assign v8c57ef = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v91177a;
assign v8b27a2 = jx0_p & v9125b3 | !jx0_p & v88ee77;
assign v8af886 = jx1_p & v8b05a5 | !jx1_p & v9123cb;
assign v91180a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8f96e8;
assign v8aee79 = stateG7_1_p & v8aeef8 | !stateG7_1_p & v9115b8;
assign v8afb9b = StoB_REQ7_p & v8c0429 | !StoB_REQ7_p & v844f91;
assign v8ae9bd = StoB_REQ0_p & v8af62a | !StoB_REQ0_p & v8b101e;
assign v91239b = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8af3b6;
assign v9121f2 = RtoB_ACK0_p & v88df14 | !RtoB_ACK0_p & v912122;
assign v8af5bd = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v890a9a;
assign v9114e5 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9124c0;
assign v912669 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c0a23;
assign v8c0bf4 = StoB_REQ3_p & v9124ed | !StoB_REQ3_p & v844f91;
assign v8afcf5 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v910e18;
assign v8b0a12 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & !v9112ad;
assign v8fed10 = StoB_REQ1_p & v881ef0 | !StoB_REQ1_p & v844f91;
assign v8b3d12 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v911fc2;
assign v8909eb = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8c4a47;
assign v8afa70 = jx3_p & v844f91 | !jx3_p & !v8c3c40;
assign v91254a = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v911ad5;
assign v8c702a = BtoR_REQ0_p & v8c704b | !BtoR_REQ0_p & v8816a0;
assign v8b3402 = jx0_p & v8b2c5c | !jx0_p & v844f91;
assign v8c5fa2 = StoB_REQ3_p & v844fb5 | !StoB_REQ3_p & !v844f91;
assign v910e1f = EMPTY_p & v8b29ed | !EMPTY_p & v8b2162;
assign v8aedac = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b2262;
assign v912565 = BtoS_ACK2_p & v8f9614 | !BtoS_ACK2_p & !v8b20b7;
assign v912769 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912651;
assign v8f9721 = jx2_p & v8c044b | !jx2_p & v910bd1;
assign v8c0a48 = StoB_REQ3_p & v912517 | !StoB_REQ3_p & v8c44a1;
assign v8aedb1 = StoB_REQ1_p & v9126f4 | !StoB_REQ1_p & v8b33ed;
assign v8b3237 = BtoS_ACK6_p & v8b33d3 | !BtoS_ACK6_p & v8b0b0c;
assign v8af0e3 = StoB_REQ0_p & v85db55 | !StoB_REQ0_p & v844f91;
assign v8b07c0 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8ae516;
assign v8858cb = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b0eab;
assign v9110bd = stateG7_1_p & v844f91 | !stateG7_1_p & v912578;
assign v911513 = jx0_p & v8af9e6 | !jx0_p & !v911c25;
assign v9126f9 = jx1_p & v8b2e60 | !jx1_p & v8b25ff;
assign v911dbb = stateG7_1_p & v8ae887 | !stateG7_1_p & v844f91;
assign v8b1ea2 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9d;
assign v8b091d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8afea2;
assign v9124f6 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v9107fb;
assign v8af7b5 = StoB_REQ2_p & v911c88 | !StoB_REQ2_p & !v912764;
assign v8b2c29 = jx3_p & v8afb96 | !jx3_p & !v844f91;
assign v8cc0fb = jx0_p & v844f91 | !jx0_p & v8b0eea;
assign v8dd65f = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8af27d;
assign v8c557c = StoB_REQ7_p & v912676 | !StoB_REQ7_p & v8ae60e;
assign v8b114d = jx0_p & v8ae8bf | !jx0_p & !v844f99;
assign v884a20 = BtoR_REQ0_p & v8b26ec | !BtoR_REQ0_p & v8b0a36;
assign v9120ec = BtoS_ACK6_p & v8af431 | !BtoS_ACK6_p & v887c34;
assign v9123da = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v911692;
assign v8b2e7b = FULL_p & v912569 | !FULL_p & v911d50;
assign v8f958b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8af753;
assign v8c6979 = jx2_p & v8af518 | !jx2_p & v910bd1;
assign v8c4667 = RtoB_ACK0_p & v8ae696 | !RtoB_ACK0_p & v8909ff;
assign v8803b6 = BtoR_REQ1_p & v9110bd | !BtoR_REQ1_p & v8b0b83;
assign v8c50c5 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v844fa1;
assign v8afb82 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b64b8;
assign v8af004 = BtoS_ACK6_p & v8af4ee | !BtoS_ACK6_p & v890b41;
assign v8af05a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b1150;
assign v8fedd4 = BtoS_ACK1_p & v8b07c0 | !BtoS_ACK1_p & v9124e2;
assign v8c3053 = BtoS_ACK7_p & v8af894 | !BtoS_ACK7_p & v8c534d;
assign v8b296a = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & !v9126cc;
assign v8ae9fc = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9112f7;
assign v8b29d6 = jx0_p & v8b1f0a | !jx0_p & !v8c3c57;
assign v8aeabb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c3e7d;
assign v8e990a = StoB_REQ2_p & v8b02a9 | !StoB_REQ2_p & v8bfa61;
assign v8cc164 = jx0_p & v8ae86c | !jx0_p & v9124c2;
assign v8af80a = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v912581;
assign v8b128f = RtoB_ACK0_p & v8af1a2 | !RtoB_ACK0_p & v844f91;
assign v8afb06 = StoB_REQ0_p & v912453 | !StoB_REQ0_p & v8b2c26;
assign v911fa9 = RtoB_ACK1_p & v8cf811 | !RtoB_ACK1_p & v9124d6;
assign v890c2c = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8b25e2;
assign v8af1ef = RtoB_ACK0_p & v8af102 | !RtoB_ACK0_p & v9124db;
assign v8b03e8 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b1367;
assign v8af986 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v85c148;
assign v8b2bc3 = stateG7_1_p & v9125a9 | !stateG7_1_p & v844f91;
assign v8bfa26 = jx1_p & v9126eb | !jx1_p & v8d6ceb;
assign v8ae151 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v8c3e7e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912593;
assign v8b02a9 = StoB_REQ3_p & v8aef02 | !StoB_REQ3_p & v844f91;
assign v91176c = jx2_p & v8c5419 | !jx2_p & !v8b065b;
assign v8c44cf = jx1_p & v844f91 | !jx1_p & v8b648c;
assign v8b0bd2 = BtoR_REQ0_p & v9126d2 | !BtoR_REQ0_p & v8ae8b7;
assign v8aea38 = jx0_p & v8ae4b3 | !jx0_p & !v8b25a2;
assign v9125ad = BtoS_ACK3_p & v88709f | !BtoS_ACK3_p & v8c6bef;
assign v9124e2 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8c04cb;
assign v89085d = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8b0764;
assign BtoS_ACK4_n = !v8fee03;
assign v875f27 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c5404;
assign v9123c4 = jx2_p & v890ac0 | !jx2_p & v91259b;
assign v8e983b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b2553;
assign v8b2792 = BtoR_REQ0_p & v8e9859 | !BtoR_REQ0_p & v8b12be;
assign v8c6e5a = BtoS_ACK3_p & v8c0bf4 | !BtoS_ACK3_p & v8b048e;
assign v91116d = BtoS_ACK6_p & v844f9e | !BtoS_ACK6_p & v8b279b;
assign v8c0ae6 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8af0e3;
assign BtoR_REQ1_n = !v892893;
assign v8c71b4 = StoB_REQ2_p & v8b2a92 | !StoB_REQ2_p & v91260b;
assign v8cc1c4 = jx1_p & v8b3383 | !jx1_p & v9125ab;
assign v8c36a2 = RtoB_ACK0_p & v912122 | !RtoB_ACK0_p & v844f91;
assign v912482 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v844f95;
assign v88bebc = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v85915c;
assign BtoS_ACK2_n = !v8b0903;
assign v8b085c = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v911f38;
assign v87d270 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v890ae8;
assign v9124d4 = jx0_p & v8aec8e | !jx0_p & v8b0750;
assign v890992 = jx0_p & v8af986 | !jx0_p & v912442;
assign v8b1e0f = ENQ_p & v9125c3 | !ENQ_p & !v912642;
assign v8c53ab = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v8b2812;
assign v8b1c70 = StoB_REQ2_p & v91274b | !StoB_REQ2_p & v9116aa;
assign v91177a = BtoS_ACK1_p & v8b034f | !BtoS_ACK1_p & v912424;
assign v8b13b1 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v9126fc;
assign v8816a0 = BtoR_REQ1_p & v911053 | !BtoR_REQ1_p & v8af02f;
assign v912796 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c715a;
assign v8c5419 = jx1_p & v8c51d8 | !jx1_p & v8b23bf;
assign v912656 = jx3_p & v8ae4b3 | !jx3_p & v8ae461;
assign v87bd82 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8909eb;
assign v8af3b6 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v91277e;
assign v91272f = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8afe22;
assign v8aea7b = BtoS_ACK6_p & v8af431 | !BtoS_ACK6_p & v8afed8;
assign v8b267f = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v8b0eab;
assign v8db203 = BtoS_ACK6_p & v8af4ee | !BtoS_ACK6_p & v912631;
assign v912517 = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & v844fb7;
assign v91100d = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v911fbd;
assign v8af84d = jx2_p & v8aef4e | !jx2_p & v8c56dd;
assign v8aeb6d = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v911733;
assign v8b0f42 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b1d1f;
assign v894826 = jx1_p & v8b0e72 | !jx1_p & !v8afa70;
assign v912477 = jx1_p & v8ae6f0 | !jx1_p & v85d63e;
assign v8b0449 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v859212;
assign v8c40de = BtoS_ACK6_p & v8c6c4a | !BtoS_ACK6_p & v8aeead;
assign v911c80 = StoB_REQ2_p & v8afe33 | !StoB_REQ2_p & v8c57aa;
assign v8afc36 = BtoS_ACK0_p & v8afe4c | !BtoS_ACK0_p & v8c575b;
assign v8aed8c = StoB_REQ6_p & v8b267f | !StoB_REQ6_p & v844f91;
assign v9123a4 = stateG7_1_p & v844f91 | !stateG7_1_p & v8afb51;
assign v88227e = BtoS_ACK6_p & v912609 | !BtoS_ACK6_p & v8d6d00;
assign v8aedf2 = StoB_REQ2_p & v8b0e57 | !StoB_REQ2_p & v8b06bc;
assign v8af5ee = BtoS_ACK7_p & v844fa1 | !BtoS_ACK7_p & !v912724;
assign v91268a = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v892e12;
assign v9125e0 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v8b2f8c;
assign v91250d = jx0_p & v8c53ab | !jx0_p & !v8c39b8;
assign v91115b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b2885;
assign v90c2e3 = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v8afc88;
assign v9124e5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88227e;
assign v8b1086 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f99;
assign v912554 = jx0_p & v844f91 | !jx0_p & !v8b25a2;
assign v86ce5c = stateG7_1_p & v8b23d9 | !stateG7_1_p & v91238f;
assign v8c460a = jx0_p & v912505 | !jx0_p & !v8c4569;
assign v91240f = stateG7_1_p & v8b0693 | !stateG7_1_p & v844f91;
assign v87d240 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v8c3d99;
assign v9124f0 = BtoS_ACK1_p & v8b229e | !BtoS_ACK1_p & v9123df;
assign v8c4a47 = BtoS_ACK0_p & v912487 | !BtoS_ACK0_p & v912683;
assign v87a09b = StoB_REQ6_p & v8b52f7 | !StoB_REQ6_p & v8c54b4;
assign v8af564 = BtoS_ACK7_p & v8b10cf | !BtoS_ACK7_p & v9124ad;
assign v9124e9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8ae169;
assign v8af40b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8ae4b6;
assign v912755 = BtoS_ACK3_p & v8b129a | !BtoS_ACK3_p & v8b339d;
assign v8dd5d4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b10fd;
assign v8afe84 = jx2_p & v91262d | !jx2_p & v8aed2e;
assign v8b07d3 = jx0_p & v890a64 | !jx0_p & v9125e8;
assign v8b0934 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v888464;
assign v8b0086 = jx0_p & v8f958b | !jx0_p & v8af02f;
assign v8b1e8a = BtoS_ACK0_p & v9123df | !BtoS_ACK0_p & v912462;
assign v9123b3 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v844f91;
assign v91264a = BtoS_ACK1_p & v8af27d | !BtoS_ACK1_p & v8b27ec;
assign v844fa5 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v8af03b = jx0_p & v8f953d | !jx0_p & v8db22c;
assign v91261a = RtoB_ACK1_p & v911d0e | !RtoB_ACK1_p & v8b2a14;
assign v8b107b = ENQ_p & v8b0a89 | !ENQ_p & v85f6d2;
assign v8b03c8 = jx2_p & v910cab | !jx2_p & v864291;
assign v8c45bc = RtoB_ACK1_p & v8af102 | !RtoB_ACK1_p & v8ae4ce;
assign v8b0e6d = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v9124c5;
assign v8c3c40 = jx0_p & v8c53ab | !jx0_p & v8b1e7d;
assign v9114ce = StoB_REQ1_p & v8b0283 | !StoB_REQ1_p & v8afd4d;
assign v91127a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8af03f;
assign v912114 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8afed5;
assign v8afe6f = ENQ_p & v8b31f9 | !ENQ_p & v911f4a;
assign v8aef95 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b1fcd;
assign v8c4517 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v91275b;
assign v8b0674 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v911664;
assign v912628 = jx3_p & v912190 | !jx3_p & v9115b8;
assign v9126e3 = jx3_p & v8b76f1 | !jx3_p & v912647;
assign v844fb9 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844f91;
assign v8b7802 = RtoB_ACK0_p & v8cf811 | !RtoB_ACK0_p & v8c6979;
assign v8b0b6b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b1199;
assign v8aeab6 = StoB_REQ0_p & v8c36bc | !StoB_REQ0_p & v8b0a04;
assign v8bfaf2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v911b07;
assign v8b021e = jx1_p & v844f91 | !jx1_p & v8b0dd3;
assign v912723 = stateG7_1_p & v8af811 | !stateG7_1_p & v844f91;
assign v9125cb = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v85c135;
assign v8afc08 = StoB_REQ7_p & v911052 | !StoB_REQ7_p & v91211a;
assign v9110d2 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844fb5;
assign v8dd5e1 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8b0fac;
assign v912643 = stateG7_1_p & v8ae670 | !stateG7_1_p & v8b28d4;
assign v8b101e = BtoS_ACK1_p & v8af27d | !BtoS_ACK1_p & v890a66;
assign v8b02b9 = jx2_p & v87f443 | !jx2_p & v910bd1;
assign v91253f = jx0_p & v91118f | !jx0_p & v8c0bc2;
assign v890bcb = jx2_p & v8af1de | !jx2_p & v8b25d9;
assign v8b01bd = jx2_p & v844f91 | !jx2_p & v8b021e;
assign v911a76 = RtoB_ACK0_p & v9124d6 | !RtoB_ACK0_p & v8c6979;
assign v8b08fa = StoB_REQ2_p & v8b0107 | !StoB_REQ2_p & v8b051e;
assign v8c77fe = StoB_REQ0_p & v8fed12 | !StoB_REQ0_p & v8ae5ca;
assign v8c466d = BtoR_REQ0_p & v8c3efe | !BtoR_REQ0_p & v87ab76;
assign v9126ad = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b267f;
assign v912765 = jx0_p & v8b10c6 | !jx0_p & v912408;
assign v912499 = RtoB_ACK1_p & v844fbb | !RtoB_ACK1_p & v8b2610;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v8b02cb = StoB_REQ2_p & v9124fe | !StoB_REQ2_p & v8b1e80;
assign v8c0bb8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ae745;
assign v8af431 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v879d5b;
assign v8aefe5 = BtoS_ACK3_p & v88709f | !BtoS_ACK3_p & v8b33a8;
assign v8894e7 = BtoR_REQ0_p & v8e9859 | !BtoR_REQ0_p & v9123e0;
assign v890ba9 = RtoB_ACK1_p & v9124a4 | !RtoB_ACK1_p & v8b0817;
assign v8b0c81 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912749;
assign v8b0dd9 = EMPTY_p & v911f8b | !EMPTY_p & v8cc139;
assign v8b0dc3 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v859212;
assign v9126b3 = StoB_REQ7_p & v8c3728 | !StoB_REQ7_p & v890534;
assign v8b22a8 = jx1_p & v8af119 | !jx1_p & !v8c3e35;
assign v912676 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v9124b4;
assign v87cf78 = StoB_REQ2_p & v9123b3 | !StoB_REQ2_p & !v8b1248;
assign v8b0c94 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b1eff;
assign v8b7892 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v912557;
assign v8b33aa = StoB_REQ0_p & v91277b | !StoB_REQ0_p & v911ffb;
assign v8b102a = jx0_p & v8ae8e5 | !jx0_p & v8af0e8;
assign v887bcf = jx2_p & v8908a2 | !jx2_p & !v9122e7;
assign v8b0b29 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v911c2f;
assign v91276a = StoB_REQ7_p & v912451 | !StoB_REQ7_p & v9126c1;
assign v8b08c4 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8b0e6d;
assign v91194c = jx2_p & v91268f | !jx2_p & v8c3af9;
assign v890a66 = StoB_REQ1_p & v8b3212 | !StoB_REQ1_p & v8c71b4;
assign v86bf27 = BtoS_ACK7_p & v912609 | !BtoS_ACK7_p & v9123c2;
assign v8b2c5c = BtoS_ACK7_p & v911149 | !BtoS_ACK7_p & v91250c;
assign v911c25 = BtoS_ACK7_p & v844f95 | !BtoS_ACK7_p & v8b26f3;
assign v8b52f7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8af62a;
assign v912784 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v911d4f;
assign v8c7305 = BtoS_ACK6_p & v912702 | !BtoS_ACK6_p & v8909eb;
assign v8f9625 = BtoS_ACK3_p & v91278c | !BtoS_ACK3_p & v844f9d;
assign v8ae731 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b77f9;
assign v91246b = RtoB_ACK0_p & v8af1a2 | !RtoB_ACK0_p & v8aebc4;
assign v8b0107 = BtoS_ACK3_p & v8b0496 | !BtoS_ACK3_p & v844f9d;
assign v8ae5a8 = BtoS_ACK6_p & v844f95 | !BtoS_ACK6_p & !v8b016b;
assign v8b2741 = jx2_p & v8c3fe8 | !jx2_p & !v844f91;
assign v8c50c4 = jx0_p & v8c45be | !jx0_p & !v91239b;
assign v91259e = ENQ_p & v890a25 | !ENQ_p & !v8fed36;
assign v8ae7ea = jx1_p & v8aea38 | !jx1_p & !v911cf2;
assign v8ae8e5 = BtoS_ACK7_p & v8c6c4a | !BtoS_ACK7_p & v9126a9;
assign v9124c5 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8b2aad;
assign v8e990d = BtoS_ACK6_p & v912609 | !BtoS_ACK6_p & v8fec78;
assign v8f95dd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ae118;
assign v8ae096 = RtoB_ACK1_p & v890960 | !RtoB_ACK1_p & v8b0994;
assign v8af463 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9126ad;
assign v91204e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9121a4;
assign v8dd5ff = BtoS_ACK7_p & v911d4f | !BtoS_ACK7_p & v8ae4ee;
assign v912693 = stateG7_1_p & v8cda2f | !stateG7_1_p & v8afb8e;
assign v912402 = jx2_p & v9126d4 | !jx2_p & v8c47de;
assign v8b6e0a = BtoS_ACK2_p & v8b327a | !BtoS_ACK2_p & v8aeab1;
assign v8c3a85 = StoB_REQ0_p & v8b08ff | !StoB_REQ0_p & v8c458d;
assign v8b0653 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8aeab6;
assign v911a59 = stateG7_1_p & v911411 | !stateG7_1_p & v844f91;
assign v911d25 = stateG7_1_p & v91241a | !stateG7_1_p & v8b52c1;
assign v8c5d1b = StoB_REQ7_p & v88b998 | !StoB_REQ7_p & v844f91;
assign v8af618 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v9117c1;
assign v911220 = jx2_p & v912467 | !jx2_p & v8ae898;
assign v8b00a7 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v911f9d;
assign v8b03ed = RtoB_ACK0_p & v91257b | !RtoB_ACK0_p & v8b28d4;
assign v9126f0 = jx0_p & v8af036 | !jx0_p & v8b05a5;
assign v91270f = jx2_p & v9110c2 | !jx2_p & v912698;
assign v88df14 = jx2_p & v875d13 | !jx2_p & v8b217f;
assign v85f6d2 = BtoR_REQ0_p & v912431 | !BtoR_REQ0_p & v8b1dd2;
assign v8674d8 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8ae516;
assign v8af7df = StoB_REQ2_p & v8b6482 | !StoB_REQ2_p & v8b0dc4;
assign v912417 = RtoB_ACK0_p & v9123b9 | !RtoB_ACK0_p & v8b2a8c;
assign v8c6e12 = jx0_p & v8b004c | !jx0_p & !v8b0f57;
assign v8b788f = stateG7_1_p & v912698 | !stateG7_1_p & v910bbe;
assign v9125e6 = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v887bcd;
assign v8b2e7a = RtoB_ACK1_p & v8b07f3 | !RtoB_ACK1_p & v8b0a89;
assign v910db7 = jx2_p & v8b1166 | !jx2_p & !v912456;
assign v8af334 = BtoS_ACK0_p & v8afe4c | !BtoS_ACK0_p & v8b09ce;
assign v8af7cb = RtoB_ACK0_p & v8909ff | !RtoB_ACK0_p & v8b0681;
assign v8b263d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8f956e;
assign v8c353f = jx3_p & v844f91 | !jx3_p & !v8b1f2d;
assign v8b23e9 = RtoB_ACK0_p & v8b23d9 | !RtoB_ACK0_p & v844f91;
assign v911fc4 = BtoS_ACK3_p & v8b340c | !BtoS_ACK3_p & v8b2c21;
assign v912390 = StoB_REQ2_p & v890a9a | !StoB_REQ2_p & v8b29c9;
assign v8b0e3d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b2019;
assign v8b11a0 = StoB_REQ2_p & v8aefe5 | !StoB_REQ2_p & v844f91;
assign v8aefc1 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8dd5d0;
assign v8b05b7 = stateG7_1_p & v8af102 | !stateG7_1_p & v9123cf;
assign v8db1c7 = stateG7_1_p & v912718 | !stateG7_1_p & v8b0dd0;
assign v8c4cc3 = jx1_p & v8c4a4e | !jx1_p & !v8b0e9d;
assign v8ae92f = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v912479;
assign v91268e = EMPTY_p & v8b09fb | !EMPTY_p & v912642;
assign v890c1b = BtoS_ACK1_p & v8c6cee | !BtoS_ACK1_p & v8f96e8;
assign v8b11ef = BtoS_ACK7_p & v8b10fd | !BtoS_ACK7_p & v8b0808;
assign v8b289a = BtoS_ACK0_p & v8f9617 | !BtoS_ACK0_p & v8b33aa;
assign v8c3b68 = BtoS_ACK1_p & v8b07c0 | !BtoS_ACK1_p & v8b267a;
assign v8b20b7 = StoB_REQ3_p & v8c43e6 | !StoB_REQ3_p & !v8b2a3e;
assign v8c37c9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8872e8;
assign v8b028a = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c41aa;
assign v8ae6ab = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v8b1eff;
assign v88ef39 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8e990e;
assign v91251d = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v8b03fc;
assign v8c4d16 = BtoS_ACK7_p & v844f95 | !BtoS_ACK7_p & !v8f9632;
assign v89288a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844fa1;
assign v8b2b17 = StoB_REQ0_p & v91277b | !StoB_REQ0_p & v890c07;
assign v8af192 = jx3_p & v844f91 | !jx3_p & !v912507;
assign v912428 = BtoS_ACK0_p & v879d5b | !BtoS_ACK0_p & v8ae6c7;
assign v8aeef8 = RtoB_ACK1_p & v8ae5e2 | !RtoB_ACK1_p & v9115b8;
assign v91230c = jx0_p & v883aaa | !jx0_p & v8b76f1;
assign v8ae75b = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8b2c37;
assign v89407e = StoB_REQ7_p & v912548 | !StoB_REQ7_p & v912711;
assign v8b12af = StoB_REQ1_p & v8b07c0 | !StoB_REQ1_p & v844f91;
assign v8c575b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b0211;
assign v8f9622 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v9032d6;
assign v8ae147 = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v8af5df;
assign v8aee08 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8b1f9c;
assign v8b2c4e = jx0_p & v8940d8 | !jx0_p & v8c5357;
assign v8db20a = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8dd5d8;
assign v910fe2 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8afb18;
assign v9125f2 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v85c0e8;
assign v8b2e66 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844fb5;
assign v8ae8bf = BtoS_ACK7_p & v91265d | !BtoS_ACK7_p & v8ae77f;
assign v8ae5ca = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b0d32;
assign v8b0705 = BtoS_ACK6_p & v911bad | !BtoS_ACK6_p & v894087;
assign v8c4b37 = StoB_REQ0_p & v8c43c1 | !StoB_REQ0_p & v8f96fd;
assign v8b71c1 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v912465;
assign v9112bc = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8b0945;
assign v88b266 = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v8af305;
assign v8b01d5 = stateG7_1_p & v8c7159 | !stateG7_1_p & v8e9896;
assign v910cda = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b1e8a;
assign v8db139 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8b0496;
assign v8fece1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b7804;
assign v8c47bf = StoB_REQ6_p & v8b0674 | !StoB_REQ6_p & v912166;
assign v864291 = jx1_p & v91174f | !jx1_p & v8b0569;
assign v8b0cfd = jx3_p & v844f91 | !jx3_p & v9124d4;
assign v8b32c2 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v910e12;
assign v8b2445 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v912474;
assign v8b0817 = jx2_p & v8b7bb1 | !jx2_p & v912742;
assign v8c6c56 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8cffee;
assign v9123a9 = stateG12_p & v9123ee | !stateG12_p & v844fbb;
assign v8b0467 = jx1_p & v8ae756 | !jx1_p & !v91248d;
assign v8ae041 = StoB_REQ3_p & v8aef02 | !StoB_REQ3_p & v912283;
assign v912672 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8b0a78;
assign v8b1d1f = StoB_REQ2_p & v9125ad | !StoB_REQ2_p & v844f91;
assign v844faf = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v8afe33 = BtoS_ACK3_p & v88709f | !BtoS_ACK3_p & v910e34;
assign v9124f9 = BtoS_ACK6_p & v8c5845 | !BtoS_ACK6_p & v9125eb;
assign v9126de = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b12af;
assign v8b05e2 = jx0_p & v8b08c4 | !jx0_p & v8af430;
assign v910df3 = StoB_REQ7_p & v8b0463 | !StoB_REQ7_p & v844f91;
assign v8aeb12 = jx0_p & v8b2878 | !jx0_p & !v844f91;
assign v9123ba = BtoS_ACK6_p & v8af894 | !BtoS_ACK6_p & v911fbe;
assign v9123e9 = BtoR_REQ1_p & v912481 | !BtoR_REQ1_p & v8b0b83;
assign v9124c3 = BtoS_ACK6_p & v912609 | !BtoS_ACK6_p & v8c5c8c;
assign v8b25a2 = BtoS_ACK7_p & v844fa1 | !BtoS_ACK7_p & !v8af916;
assign v8b02b0 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8af4b1;
assign v8b0877 = BtoS_ACK0_p & v8b229e | !BtoS_ACK0_p & v8b0151;
assign v8b2911 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b0dc3;
assign v8cc202 = jx0_p & v911e75 | !jx0_p & v8c6cd3;
assign v8af4fa = jx0_p & v8ae4b3 | !jx0_p & v844f91;
assign v9123c2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9112b6;
assign v8b1dd2 = BtoR_REQ1_p & v911532 | !BtoR_REQ1_p & v844f91;
assign v8b3286 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v912744;
assign v8b2f6c = StoB_REQ2_p & v87e29c | !StoB_REQ2_p & v911aa3;
assign v8af0e6 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v912555;
assign v8af2e0 = stateG7_1_p & v8b01a4 | !stateG7_1_p & v8b0963;
assign v910cab = jx1_p & v8b2a71 | !jx1_p & v85d9b6;
assign v8b1247 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b2fea;
assign v912636 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ae93f;
assign v8aeb91 = StoB_REQ6_p & v9125ea | !StoB_REQ6_p & v844f91;
assign v88acc3 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912451;
assign v911382 = jx0_p & v8b0a03 | !jx0_p & v8b11c4;
assign v87ed24 = stateG7_1_p & v844f91 | !stateG7_1_p & v8b2c0d;
assign v91247b = jx1_p & v8aea38 | !jx1_p & !v8c6cae;
assign v8b2929 = BtoS_ACK1_p & v911787 | !BtoS_ACK1_p & v8b101c;
assign v8c70fc = BtoR_REQ0_p & v8af025 | !BtoR_REQ0_p & v8ae9f2;
assign v85c13e = jx3_p & v844f91 | !jx3_p & v91269c;
assign BtoR_REQ0_n = v8940f1;
assign v8aeada = jx0_p & v8b028a | !jx0_p & v8b7791;
assign v911fe3 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v912592;
assign v87c076 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8b2080;
assign v911faa = jx1_p & v8771a0 | !jx1_p & v9126b8;
assign v8c57aa = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8afe33;
assign v911c45 = RtoB_ACK0_p & v912649 | !RtoB_ACK0_p & v8c66bb;
assign v8c3c0d = BtoS_ACK0_p & v8b0df4 | !BtoS_ACK0_p & v9126f5;
assign v8b3013 = BtoS_ACK1_p & v911787 | !BtoS_ACK1_p & v8afc92;
assign v8b2e22 = jx1_p & v8b2920 | !jx1_p & !v8b2d81;
assign v8ae673 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b76c6;
assign v8c3d4b = ENQ_p & v8b02e9 | !ENQ_p & !v8b0a17;
assign v8c4569 = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v9123b7;
assign v911197 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88ffd6;
assign v8aebc4 = jx2_p & v911ed6 | !jx2_p & !v8b0c98;
assign v8db28c = DEQ_p & v8b1cf2 | !DEQ_p & v8b01dd;
assign v91277d = jx0_p & v88bb7a | !jx0_p & v8b2eb4;
assign v8aec57 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9b;
assign v9111c2 = stateG12_p & v8d6d2c | !stateG12_p & v8b2d68;
assign v8b0494 = StoB_REQ7_p & v8b3399 | !StoB_REQ7_p & v844f91;
assign v91258f = BtoS_ACK7_p & v844f9e | !BtoS_ACK7_p & v91116d;
assign v91275b = StoB_REQ6_p & v8af7a3 | !StoB_REQ6_p & v8c0509;
assign v8ae07b = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v8b32e2;
assign v863839 = jx1_p & v8af4fa | !jx1_p & v844f91;
assign v8b32e2 = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & v8af634;
assign v88bb7a = BtoS_ACK7_p & v8b0661 | !BtoS_ACK7_p & v8ae803;
assign v844f9f = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & !v844f91;
assign v91161f = jx1_p & v8b2a71 | !jx1_p & v9123f5;
assign v8b2e92 = StoB_REQ6_p & v8e983b | !StoB_REQ6_p & v912784;
assign v9123d4 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8dd5d4;
assign v8af894 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8ae151;
assign v8c3e1b = stateG7_1_p & v9123b1 | !stateG7_1_p & !v8b04f8;
assign v912744 = StoB_REQ1_p & v8b139e | !StoB_REQ1_p & v8b038f;
assign v89098c = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v9116c4;
assign v8b085a = jx1_p & v9115b8 | !jx1_p & v912628;
assign v8ae4e9 = StoB_REQ6_p & v8dd6a6 | !StoB_REQ6_p & v844f91;
assign v8b2d81 = jx3_p & v8af5ee | !jx3_p & !v894072;
assign v8b2ba1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b0877;
assign v8affe8 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8aede2;
assign v8b339d = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9d;
assign v9123e2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c71fb;
assign v9125f8 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v91259a;
assign v8b2bc5 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v87cf78;
assign v890b86 = BtoR_REQ0_p & v911a8d | !BtoR_REQ0_p & v9114d3;
assign v8b19b1 = stateG7_1_p & v8b051c | !stateG7_1_p & v88acc3;
assign v8ae0b9 = StoB_REQ6_p & v887bda | !StoB_REQ6_p & v844f91;
assign v8e9954 = jx1_p & v8b2c39 | !jx1_p & v890ac0;
assign v8b65a3 = stateG7_1_p & v890ba9 | !stateG7_1_p & v887b53;
assign v8aefa4 = BtoS_ACK3_p & v8c38b4 | !BtoS_ACK3_p & v912517;
assign v8af763 = jx2_p & v8afd1f | !jx2_p & v8af886;
assign v912291 = BtoS_ACK6_p & v911d4f | !BtoS_ACK6_p & v912784;
assign v88abc8 = jx0_p & v8dd5e1 | !jx0_p & v912442;
assign v8b0fa3 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8ae7b3;
assign v8c0b95 = stateG7_1_p & v91101e | !stateG7_1_p & v9114e3;
assign v8afed5 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v8b2ba1;
assign v8aebc8 = jx1_p & v844f91 | !jx1_p & v8b27a2;
assign v911fad = jx0_p & v8af9e6 | !jx0_p & v844f91;
assign v8afd22 = BtoR_REQ1_p & v9123ec | !BtoR_REQ1_p & v912678;
assign v912514 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b1083;
assign v8c53cf = ENQ_p & v8af02f | !ENQ_p & v9125e5;
assign v8aea07 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8b296a;
assign v8b0062 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v912648;
assign v8b276b = EMPTY_p & v88b266 | !EMPTY_p & v9118c2;
assign v8e9852 = jx0_p & v911218 | !jx0_p & v8afcd6;
assign v885d39 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8c0ab9;
assign v9126cb = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v912501;
assign v8af89d = jx1_p & v8b8bdf | !jx1_p & v8aec42;
assign v8b2464 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8af53c;
assign v8b0808 = BtoS_ACK6_p & v8b10fd | !BtoS_ACK6_p & v8dd5d4;
assign v8b0cbb = StoB_REQ6_p & v8b2019 | !StoB_REQ6_p & v844f91;
assign v8b06bc = BtoS_ACK3_p & v8ae5ff | !BtoS_ACK3_p & !v844f91;
assign v8cfeeb = stateG7_1_p & v8b1eeb | !stateG7_1_p & v8b1d83;
assign v8618ae = jx1_p & v912074 | !jx1_p & !v8b102a;
assign v912182 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v910ba7;
assign v912605 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8aef7a;
assign v8b1e70 = jx0_p & v8e98af | !jx0_p & v9125e8;
assign v912548 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844faf;
assign v91220c = ENQ_p & v8aeb6d | !ENQ_p & v8af5b7;
assign v8aed6d = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v910d59;
assign v8b1fc5 = StoB_REQ6_p & v8b25f9 | !StoB_REQ6_p & v9124a0;
assign v8b2c21 = StoB_REQ3_p & v912517 | !StoB_REQ3_p & v8b2a3e;
assign v8b1ec1 = BtoS_ACK7_p & v8c6c4a | !BtoS_ACK7_p & v8aed6c;
assign v8b26af = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e9884;
assign v882fb4 = jx0_p & v8b2420 | !jx0_p & v912691;
assign v8fedc9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v88ef39;
assign v8b1e91 = BtoS_ACK7_p & v8ae4e9 | !BtoS_ACK7_p & v9124bc;
assign v911fc3 = jx3_p & v9110f5 | !jx3_p & !v8af55a;
assign v8b21eb = jx1_p & v8b0086 | !jx1_p & v8af02f;
assign v8aeec4 = jx1_p & v9126eb | !jx1_p & v912391;
assign v8c3fe8 = jx1_p & v8ae6f0 | !jx1_p & !v844f91;
assign v912068 = BtoS_ACK3_p & v8af85c | !BtoS_ACK3_p & v8b2b08;
assign v8c5d1c = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8b1f50;
assign v8b274c = ENQ_p & v9124e6 | !ENQ_p & !v910e1f;
assign v8c71fb = BtoS_ACK1_p & v8c6cee | !BtoS_ACK1_p & v8aee21;
assign v890a25 = jx2_p & v8c3fe8 | !jx2_p & v8ae6e0;
assign v911c7e = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b238a;
assign v911695 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v911e9b;
assign v9123ca = jx2_p & v912511 | !jx2_p & !v8af2cd;
assign v9124ea = StoB_REQ6_p & v912584 | !StoB_REQ6_p & v911940;
assign v892ea4 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v8afea6;
assign v8b0ebf = BtoR_REQ1_p & v911053 | !BtoR_REQ1_p & v8c3d7b;
assign v8c387f = jx2_p & v8b2e07 | !jx2_p & v8ae5c6;
assign v8c3973 = StoB_REQ0_p & v8af80a | !StoB_REQ0_p & v8b32c2;
assign v8b64b8 = BtoS_ACK6_p & v8ae578 | !BtoS_ACK6_p & v8af72b;
assign v8af4ee = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8db217;
assign v910bd3 = StoB_REQ7_p & v8b238a | !StoB_REQ7_p & v8b236f;
assign v912598 = RtoB_ACK0_p & v8b0a19 | !RtoB_ACK0_p & !v9123b1;
assign v8af36f = StoB_REQ0_p & v8af9be | !StoB_REQ0_p & v844f91;
assign v8b2e23 = StoB_REQ7_p & v8c6bfa | !StoB_REQ7_p & v844f91;
assign v911289 = jx2_p & v8af02f | !jx2_p & v8b52fa;
assign v8af305 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v911dbb;
assign v9124e6 = BtoR_REQ0_p & v8af366 | !BtoR_REQ0_p & v91275a;
assign v8940af = jx0_p & v8b0298 | !jx0_p & !v8591f3;
assign v912748 = BtoS_ACK6_p & v911bad | !BtoS_ACK6_p & v8b2cb0;
assign v8b0750 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b09a9;
assign v912485 = jx0_p & v8afd20 | !jx0_p & v9125c8;
assign v91269c = jx0_p & v844f91 | !jx0_p & !v8b1e7d;
assign v8b2a63 = RtoB_ACK1_p & v8909ff | !RtoB_ACK1_p & v8b0681;
assign v8b116b = RtoB_ACK0_p & v8b1f9c | !RtoB_ACK0_p & v844f91;
assign v9123e3 = StoB_REQ6_p & v8b232f | !StoB_REQ6_p & v8b4fda;
assign v8afdb9 = EMPTY_p & v8c466d | !EMPTY_p & v8aeccb;
assign v8ae446 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b2f6b;
assign v8ae4a5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v88413b;
assign v9123dd = BtoS_ACK7_p & v8b33d3 | !BtoS_ACK7_p & v9123a3;
assign v85c0ba = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9125a8;
assign v8c70fd = jx1_p & v8ae6f2 | !jx1_p & !v8b2a34;
assign v8b26f3 = BtoS_ACK6_p & v844f95 | !BtoS_ACK6_p & v912482;
assign v89097f = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8dd6de;
assign v9126ff = stateG12_p & v91230d | !stateG12_p & v8b1ca6;
assign v8b1410 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v91171d;
assign v8b21e7 = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v8aebc5;
assign v8b3321 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9d;
assign v911eb1 = ENQ_p & v911fd5 | !ENQ_p & v8b2639;
assign v8aff01 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9e;
assign v8d6d16 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b5a58;
assign v8c5845 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v844f97;
assign v88ee77 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0109;
assign v8b068c = jx0_p & v8b021d | !jx0_p & v8c4d14;
assign v8b3403 = jx0_p & v9114e1 | !jx0_p & v8c3541;
assign v8af23b = BtoS_ACK2_p & v8924d2 | !BtoS_ACK2_p & v8b048e;
assign v8b0339 = stateG7_1_p & v844fa7 | !stateG7_1_p & v844fa5;
assign v8c557b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v9123d1;
assign v9123ef = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v8afea6;
assign v9125a6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v9123fa;
assign v8b09f9 = RtoB_ACK1_p & v9123b9 | !RtoB_ACK1_p & v8b2a8c;
assign v8b32b6 = jx0_p & v9126aa | !jx0_p & v88acc3;
assign v8b1d03 = StoB_REQ0_p & v912635 | !StoB_REQ0_p & v844f91;
assign v8b21a3 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9126e7;
assign v911c9a = stateG7_1_p & v91253b | !stateG7_1_p & v8c66bb;
assign v85c182 = DEQ_p & v8cc182 | !DEQ_p & v911e03;
assign v9126cc = StoB_REQ2_p & v8b0d58 | !StoB_REQ2_p & !v8b07ff;
assign v912407 = stateG7_1_p & v844f91 | !stateG7_1_p & v8b23e9;
assign v85db55 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b22a7;
assign v9113da = stateG7_1_p & v844f91 | !stateG7_1_p & v844fa5;
assign v8dd5d0 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8c3973;
assign v8c5356 = BtoS_ACK3_p & v9110d2 | !BtoS_ACK3_p & v8db23e;
assign v8b0113 = jx1_p & v8aea38 | !jx1_p & !v88abc8;
assign v8c7026 = StoB_REQ3_p & v892ea4 | !StoB_REQ3_p & v844f9f;
assign v912652 = StoB_REQ7_p & v87c076 | !StoB_REQ7_p & v844f91;
assign v91159f = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8aed8c;
assign v8b23d9 = jx2_p & v8ae0b8 | !jx2_p & v8c3af9;
assign v91271e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v912026;
assign v8b2162 = FULL_p & v8b29d9 | !FULL_p & v8b1f1b;
assign v9124fb = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v912793;
assign v8c3d77 = jx0_p & v8aff37 | !jx0_p & v8af71d;
assign v8b2ba6 = stateG7_1_p & v8c420b | !stateG7_1_p & v91194c;
assign v8c715c = BtoS_ACK6_p & v91222a | !BtoS_ACK6_p & v9116ad;
assign v91267c = BtoS_ACK3_p & v8b1fb5 | !BtoS_ACK3_p & v8fece4;
assign v9117c1 = jx2_p & v844f91 | !jx2_p & v8b1d6c;
assign v8b06b8 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8aeb29;
assign v8ae88e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8ae714;
assign v8fecf0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b055a;
assign v8dd632 = jx1_p & v844f91 | !jx1_p & v8ae031;
assign v8b0b2b = jx0_p & v8b1cd0 | !jx0_p & !v8c6c18;
assign v911075 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b33d3;
assign v8af1ad = jx2_p & v8b2a9f | !jx2_p & v8b24af;
assign v9125ce = RtoB_ACK0_p & v8c6979 | !RtoB_ACK0_p & v9124d6;
assign v8d6d2f = DEQ_p & v8c3d4b | !DEQ_p & v8b274c;
assign v89342c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9125eb;
assign v890ba5 = StoB_REQ0_p & v844f97 | !StoB_REQ0_p & v844f91;
assign v8c48a1 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8af372;
assign v91251c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v91266f;
assign v8a8ba3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v8b2e42 = BtoR_REQ1_p & v87ed24 | !BtoR_REQ1_p & v9125af;
assign v8b4ffd = DEQ_p & v86f676 | !DEQ_p & v91259e;
assign v911e65 = stateG7_1_p & v8c50eb | !stateG7_1_p & v9124f2;
assign v8afbd6 = jx0_p & v8b0774 | !jx0_p & v844f91;
assign v912513 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v91271c;
assign v912391 = jx0_p & v8aea72 | !jx0_p & !v844f9d;
assign v91207b = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v91278b;
assign v910d59 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8db288;
assign v91240c = StoB_REQ2_p & v8b23c7 | !StoB_REQ2_p & v8af9e8;
assign v8b0fab = jx2_p & v911d2c | !jx2_p & v912742;
assign v8f9631 = jx0_p & v8b1f0a | !jx0_p & !v8fecad;
assign v8ae97e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9124ff;
assign v8b1d12 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8b7804;
assign v8b1e15 = jx2_p & v9123ce | !jx2_p & v8afe97;
assign v91273c = BtoS_ACK1_p & v8b327a | !BtoS_ACK1_p & v8b12eb;
assign v8b218f = RtoB_ACK1_p & v8af1a2 | !RtoB_ACK1_p & v8b1f9c;
assign v911f9c = jx2_p & v8b03d4 | !jx2_p & v91155b;
assign v8fec78 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b03fe;
assign v8af155 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v9126f7;
assign v85f776 = BtoR_REQ1_p & v91272c | !BtoR_REQ1_p & v844f91;
assign jx1_n = !v8d6d2f;
assign v912555 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91255a;
assign v8af26f = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b01e2;
assign v85aa58 = BtoR_REQ0_p & v8b2bc3 | !BtoR_REQ0_p & v8b2e42;
assign v8d6d04 = StoB_REQ1_p & v912520 | !StoB_REQ1_p & v844f91;
assign v8b1dbe = BtoS_ACK6_p & v8ae578 | !BtoS_ACK6_p & v9123d3;
assign v8cffee = BtoS_ACK3_p & v8c38b4 | !BtoS_ACK3_p & v8c0a48;
assign v910c25 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v8cc129;
assign v911704 = RtoB_ACK1_p & v8aebc4 | !RtoB_ACK1_p & v844f91;
assign v911529 = jx0_p & v8ae8bf | !jx0_p & !v85c141;
assign v8ae789 = StoB_REQ2_p & v8b0fa3 | !StoB_REQ2_p & !v8ae7b3;
assign v912735 = StoB_REQ2_p & v8c537f | !StoB_REQ2_p & v8b02b0;
assign v8b21ba = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v9117c1;
assign v890b4a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v9126bc;
assign v8b032e = jx0_p & v8b1276 | !jx0_p & v844f91;
assign v9126c4 = BtoS_ACK2_p & v844f9e | !BtoS_ACK2_p & v8aff01;
assign v8b082d = jx1_p & v8b320b | !jx1_p & v88f796;
assign v8b217f = jx1_p & v911a0d | !jx1_p & v8b02de;
assign v8b2000 = RtoB_ACK1_p & v8c723e | !RtoB_ACK1_p & v912664;
assign v912122 = jx2_p & v8b2e24 | !jx2_p & v8b21c9;
assign v8b02de = jx3_p & v9110f5 | !jx3_p & !v91250d;
assign v89209f = jx2_p & v8b2fc8 | !jx2_p & v91155b;
assign v8ae06b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b2bbf;
assign v9125b0 = RtoB_ACK0_p & v8b2559 | !RtoB_ACK0_p & v8909ff;
assign v910884 = jx2_p & v87cf4c | !jx2_p & v8b2e22;
assign v91263c = StoB_REQ1_p & v8aee6c | !StoB_REQ1_p & v844f91;
assign v8aed7b = jx0_p & v8b233e | !jx0_p & v8fecd9;
assign v8c47de = jx1_p & v8c6cb4 | !jx1_p & v9125ae;
assign v9126aa = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0c81;
assign v9126a9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c40de;
assign v91248a = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v9124bd;
assign v9123c8 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v910df3;
assign v912706 = BtoS_ACK6_p & v8af4ee | !BtoS_ACK6_p & v8c0b6f;
assign v8b1d80 = BtoS_ACK1_p & v8afd76 | !BtoS_ACK1_p & v911fea;
assign v8bfa79 = BtoS_ACK1_p & v912557 | !BtoS_ACK1_p & v9124e2;
assign v8af168 = BtoS_ACK6_p & v8c5845 | !BtoS_ACK6_p & v911fe4;
assign v87dbe0 = stateG7_1_p & v844f91 | !stateG7_1_p & v8c36a2;
assign v8c6bfa = BtoS_ACK6_p & v844f95 | !BtoS_ACK6_p & !v8a8ba3;
assign v8b3416 = jx1_p & v8c706b | !jx1_p & v8c3e60;
assign v8ae0a2 = BtoR_REQ0_p & v8b02ce | !BtoR_REQ0_p & v8afd22;
assign v910d0e = BtoS_ACK7_p & v8ae578 | !BtoS_ACK7_p & v8fecf0;
assign v8aeed6 = BtoS_ACK2_p & v8b33a8 | !BtoS_ACK2_p & v8c0457;
assign v912650 = jx1_p & v91180b | !jx1_p & v911b4f;
assign v91250a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af748;
assign v912647 = jx0_p & v890aa5 | !jx0_p & v8b76f1;
assign v8c0509 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v91216a;
assign v8839ea = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v8c715c;
assign v911bc6 = StoB_REQ7_p & v9125e3 | !StoB_REQ7_p & v912190;
assign v912761 = jx0_p & v8ae83c | !jx0_p & v91254d;
assign v8b25f8 = jx0_p & v8c0a9d | !jx0_p & v8c5357;
assign v8b28d5 = jx2_p & v844f91 | !jx2_p & v9123cd;
assign v8b33d3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f97;
assign v912550 = BtoR_REQ1_p & v844fbb | !BtoR_REQ1_p & v9123ab;
assign v8af372 = StoB_REQ2_p & v8aec57 | !StoB_REQ2_p & v8afaed;
assign v890ae8 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8b52f8;
assign v9125c7 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v9126b2;
assign v8c23d8 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8b2657;
assign v8c39e2 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8ae0b9;
assign v9118e7 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912576;
assign v8b2a3e = StoB_REQ4_p & v844f9f | !StoB_REQ4_p & v844f91;
assign v9123b7 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v9123c7;
assign v8b76f1 = BtoS_ACK7_p & v8577c2 | !BtoS_ACK7_p & v8b09a9;
assign v91248d = jx3_p & v844f91 | !jx3_p & v91243e;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v912739 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8aea7b;
assign v844fa1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v844f91;
assign v8af205 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v910c9d;
assign v8b0b9c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v87d240;
assign v911e3b = jx2_p & v8c34ba | !jx2_p & v85c0eb;
assign v91093d = StoB_REQ0_p & v8b0554 | !StoB_REQ0_p & v844f91;
assign v8b2815 = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v8b029e;
assign v8b25e2 = StoB_REQ7_p & v8b1f50 | !StoB_REQ7_p & v9125c7;
assign v8ae81f = jx2_p & v912698 | !jx2_p & v8c5cc7;
assign v8ae6ee = BtoS_ACK6_p & v9126de | !BtoS_ACK6_p & v8af808;
assign v91104c = BtoS_ACK6_p & v912518 | !BtoS_ACK6_p & v8b28c6;
assign v8aea88 = BtoS_ACK1_p & v8c0b8f | !BtoS_ACK1_p & v912662;
assign v911fea = StoB_REQ1_p & v8b139e | !StoB_REQ1_p & v8b28fe;
assign v91153e = RtoB_ACK1_p & v911bcd | !RtoB_ACK1_p & v8af84d;
assign v91262d = jx1_p & v8ae6f2 | !jx1_p & !v8c48c7;
assign v8b77fc = StoB_REQ7_p & v912776 | !StoB_REQ7_p & v9126ab;
assign v912520 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v88709f;
assign v8c6c93 = jx0_p & v8b1129 | !jx0_p & v912691;
assign v911ea9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e98d6;
assign v9125d8 = BtoS_ACK6_p & v890ba5 | !BtoS_ACK6_p & v91268b;
assign v8e988e = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & !v844fad;
assign v8fec67 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8ae160;
assign v912750 = BtoS_ACK0_p & v91244d | !BtoS_ACK0_p & v8af651;
assign v91278f = jx0_p & v8b1f0a | !jx0_p & !v8b062d;
assign v9115e4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87e9d4;
assign v8af3eb = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v8b3321;
assign v8b1385 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ae6ee;
assign v912461 = jx1_p & v8c3c57 | !jx1_p & v912775;
assign v8b2f4e = jx0_p & v910d0e | !jx0_p & !v8cc104;
assign v8ae806 = stateG12_p & v8af1e9 | !stateG12_p & v8b0358;
assign v8b016d = jx0_p & v8afcaa | !jx0_p & v912515;
assign v8b0298 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8c6aa0;
assign v912788 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8b6482;
assign v8b2a7e = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8b1e10;
assign v892e44 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8af582;
assign v8c3e7d = BtoS_ACK1_p & v879d5b | !BtoS_ACK1_p & v8e990e;
assign v9113cc = jx1_p & v8b320b | !jx1_p & v8dd5d6;
assign v911a5e = jx2_p & v8b1166 | !jx2_p & v8b1d6c;
assign v8aeccb = FULL_p & v85aa58 | !FULL_p & v890ab8;
assign v887afb = jx0_p & v844f9b | !jx0_p & !v8b76f1;
assign v8c3b8d = StoB_REQ0_p & v8fed12 | !StoB_REQ0_p & v8b094a;
assign v912668 = BtoS_ACK7_p & v8b327a | !BtoS_ACK7_p & v912780;
assign v8c498b = jx1_p & v8890ee | !jx1_p & v8b244a;
assign v8b2c79 = BtoS_ACK6_p & v9126de | !BtoS_ACK6_p & v9126a1;
assign v8af601 = jx1_p & v911529 | !jx1_p & v8b2c52;
assign v912509 = jx0_p & v9126b9 | !jx0_p & v8af0ef;
assign v8ae956 = jx2_p & v911faa | !jx2_p & v8b22a8;
assign v8b8bdf = jx0_p & v8b0fb5 | !jx0_p & v87ebfd;
assign v912768 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b2cc1;
assign v8ae4b6 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8b2c35;
assign v8e992f = BtoS_ACK6_p & v911bad | !BtoS_ACK6_p & v91246d;
assign v8d6d1f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c3b68;
assign v8b0a89 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c3728;
assign v8c3728 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b0500;
assign v8b2c37 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8b7443;
assign v8b0463 = BtoS_ACK6_p & v912518 | !BtoS_ACK6_p & v887bda;
assign v8b2bd9 = BtoR_REQ1_p & v887acc | !BtoR_REQ1_p & v8c3050;
assign v8c3a82 = jx0_p & v91183d | !jx0_p & v8aed6d;
assign v8b330f = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8b0b9e;
assign v910c72 = stateG7_1_p & v912672 | !stateG7_1_p & v91116e;
assign v912749 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9125a6;
assign v9112f7 = StoB_REQ7_p & v8c3728 | !StoB_REQ7_p & v8b1f71;
assign v911052 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8af2bd;
assign v85f4b2 = jx2_p & v912477 | !jx2_p & !v8b0467;
assign v9125ea = BtoS_ACK0_p & v8b7804 | !BtoS_ACK0_p & v912518;
assign v85c0e8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91254a;
assign v8af0fb = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91270b;
assign v912154 = EMPTY_p & v8b0358 | !EMPTY_p & v8ae806;
assign v8b013b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b261e;
assign v91271f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b3d0c;
assign v8b26ec = stateG7_1_p & v8aef35 | !stateG7_1_p & v9121f2;
assign v8b22c9 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8af698;
assign v91249b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9111d2;
assign v8b7bb1 = jx1_p & v8ae6f2 | !jx1_p & !v91272e;
assign v8af430 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v89097b;
assign v9123f0 = BtoR_REQ0_p & v911fe2 | !BtoR_REQ0_p & v8c57f0;
assign v8fecad = BtoS_ACK7_p & v8ae02e | !BtoS_ACK7_p & v8f95dd;
assign v8b021d = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v85a47c;
assign v91256e = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8b00a9;
assign v91258c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v91276f;
assign v8c34da = jx1_p & v8cc164 | !jx1_p & v9124c2;
assign v912413 = jx2_p & v91257c | !jx2_p & !v91257a;
assign v9124a5 = BtoR_REQ0_p & v8b0a5f | !BtoR_REQ0_p & v911632;
assign v8c55bf = jx2_p & v8b02ab | !jx2_p & v8af601;
assign v8b029c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b3237;
assign v8b0963 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8af1ad;
assign v9110fc = stateG12_p & v8b2f92 | !stateG12_p & v8c702a;
assign v8940eb = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0dd4;
assign v87b5cf = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8ae0ee;
assign v8b03fc = StoB_REQ3_p & v8c6c00 | !StoB_REQ3_p & v844f91;
assign v8b04f4 = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v8b31b3;
assign v912490 = RtoB_ACK1_p & v8af98a | !RtoB_ACK1_p & v844f91;
assign v8aecbf = RtoB_ACK1_p & v8b28d4 | !RtoB_ACK1_p & v8f9630;
assign v8aee3c = StoB_REQ2_p & v844fb1 | !StoB_REQ2_p & v844f91;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v912409 = stateG7_1_p & v8c369a | !stateG7_1_p & v8af763;
assign v8b1e33 = StoB_REQ6_p & v8b0acf | !StoB_REQ6_p & v8b2fc3;
assign v911f49 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86d734;
assign v911bcd = jx2_p & v8b7801 | !jx2_p & v8b002e;
assign v8b0436 = BtoS_ACK0_p & v8b07c0 | !BtoS_ACK0_p & v8b0eab;
assign v8b2a14 = jx2_p & v8cc0f1 | !jx2_p & v9113a8;
assign v91266f = StoB_REQ2_p & v8f9625 | !StoB_REQ2_p & v912556;
assign v91244d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b034f;
assign v8b1068 = jx3_p & v844f91 | !jx3_p & v881e63;
assign v9123f7 = BtoS_ACK0_p & v8c0b8f | !BtoS_ACK0_p & v8c3a85;
assign v91219b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f99;
assign v8b12fb = StoB_REQ6_p & v9113eb | !StoB_REQ6_p & v8b289a;
assign v8afc85 = stateG7_1_p & v8c6979 | !stateG7_1_p & v911a76;
assign v912424 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v9124c9;
assign v8af74b = stateG7_1_p & v8f9721 | !stateG7_1_p & v8b02b9;
assign v8ae854 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8b2cf0;
assign v85c16c = BtoS_ACK2_p & v88709f | !BtoS_ACK2_p & v8afe33;
assign v91265d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b7794;
assign v9124d7 = jx1_p & v8771a0 | !jx1_p & v912705;
assign v8b2460 = ENQ_p & v911ff4 | !ENQ_p & v9124df;
assign v8af7c1 = BtoR_REQ0_p & v912682 | !BtoR_REQ0_p & v882eb7;
assign v8af5df = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v911fc4;
assign v8af960 = BtoR_REQ1_p & v912407 | !BtoR_REQ1_p & v8c6dfc;
assign v8b284f = jx2_p & v91247b | !jx2_p & !v8af2ab;
assign v8af82e = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v8b0a12;
assign v9124dd = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912636;
assign v8afbaa = RtoB_ACK1_p & v8afa71 | !RtoB_ACK1_p & v912444;
assign v8ae4ee = BtoS_ACK6_p & v911d4f | !BtoS_ACK6_p & v91263e;
assign v8bfa12 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v910c58;
assign v8b0fee = BtoS_ACK2_p & v8b33a8 | !BtoS_ACK2_p & v844f91;
assign v912609 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8d6d04;
assign v8b2d73 = RtoB_ACK1_p & v9123b1 | !RtoB_ACK1_p & v8dd6de;
assign v8b1ff0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9125e0;
assign v887bdb = jx0_p & v912505 | !jx0_p & !v844f99;
assign v86bd18 = jx1_p & v887afb | !jx1_p & !v8b76f1;
assign v8b1f1b = BtoR_REQ0_p & v9123de | !BtoR_REQ0_p & v8b76ff;
assign v8b4fca = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8ae97e;
assign v91188e = StoB_REQ1_p & v9124ab | !StoB_REQ1_p & v844f91;
assign v911ffb = BtoS_ACK1_p & v8afd76 | !BtoS_ACK1_p & v8aedc9;
assign v8ae5ff = StoB_REQ3_p & v8b2a3e | !StoB_REQ3_p & !v844f91;
assign v8dd5d9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8612be;
assign v887b30 = stateG7_1_p & v8b0ae4 | !stateG7_1_p & v88acc3;
assign v88709f = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9f;
assign v844fb5 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f91;
assign v912430 = stateG7_1_p & v8c66bb | !stateG7_1_p & v911c45;
assign v8b2262 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b0223;
assign v8c5e4c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9126b3;
assign v8bfab2 = BtoS_ACK6_p & v8c6c4a | !BtoS_ACK6_p & v91258c;
assign v9124f3 = BtoS_ACK0_p & v8c0b8f | !BtoS_ACK0_p & v8aeeaa;
assign v8c5350 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8c3c0d;
assign v912691 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b2e23;
assign v8b293f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b2789;
assign v91144e = BtoR_REQ1_p & v912729 | !BtoR_REQ1_p & !v844f91;
assign v8b2c06 = BtoS_ACK6_p & v8b10fd | !BtoS_ACK6_p & v9123d4;
assign v8c57d1 = stateG7_1_p & v911fa9 | !stateG7_1_p & v9125ce;
assign v8ae031 = jx0_p & v8b07b6 | !jx0_p & !v844f9d;
assign v8b0f67 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v912525;
assign v8c6c8b = StoB_REQ6_p & v8b232f | !StoB_REQ6_p & v8b289a;
assign v8b0d9e = BtoS_ACK6_p & v890ba5 | !BtoS_ACK6_p & v912732;
assign v912730 = StoB_REQ6_p & v8c0bb8 | !StoB_REQ6_p & v9124f3;
assign v9123ab = stateG7_1_p & v912499 | !stateG7_1_p & v844fbb;
assign v8af651 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911742;
assign v8dd654 = BtoR_REQ1_p & v887acc | !BtoR_REQ1_p & v8b1fc9;
assign v8afd76 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8924d2;
assign v8cc197 = jx2_p & v91263d | !jx2_p & v8c04c4;
assign v9124be = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b2073;
assign v8afe06 = BtoS_ACK6_p & v8c426f | !BtoS_ACK6_p & v86c179;
assign v8c0457 = BtoS_ACK3_p & v8b33a8 | !BtoS_ACK3_p & v8ae487;
assign v8af7f1 = StoB_REQ0_p & v890b15 | !StoB_REQ0_p & v8aea88;
assign v9126c1 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912783;
assign v9112aa = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8c09e5;
assign v8c049b = stateG7_1_p & v844f91 | !stateG7_1_p & v8e9855;
assign v8c3e60 = jx3_p & v87a52a | !jx3_p & v8b24b0;
assign v8b6d47 = jx1_p & v8b2a71 | !jx1_p & v912236;
assign v8b24b7 = StoB_REQ6_p & v8b0674 | !StoB_REQ6_p & v8b6f1f;
assign v8b1e10 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8afedf;
assign v8b0fb9 = StoB_REQ2_p & v85c0ac | !StoB_REQ2_p & v8b22c6;
assign v910c1b = BtoS_ACK7_p & v864227 | !BtoS_ACK7_p & v8ae4a5;
assign v8c0bc2 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8af624;
assign v8ae048 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8aed0c;
assign v8b02d7 = StoB_REQ7_p & v912291 | !StoB_REQ7_p & v8b2a5b;
assign v85c164 = stateG7_1_p & v8cf811 | !stateG7_1_p & v8c23b9;
assign v9113a8 = jx1_p & v8b3403 | !jx1_p & v8afa37;
assign v894810 = BtoR_REQ1_p & v8b265b | !BtoR_REQ1_p & v9115b8;
assign v8d6ceb = jx0_p & v8aea72 | !jx0_p & !v8bfa76;
assign v911367 = StoB_REQ2_p & v8ae83f | !StoB_REQ2_p & v8b0e4c;
assign v892551 = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v8b2b4a;
assign v8ae4cd = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b3321;
assign v8c47c3 = BtoR_REQ1_p & v911d25 | !BtoR_REQ1_p & v911e65;
assign v8c36bc = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b6d3d;
assign v8aec17 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b1cd7;
assign v911fb2 = BtoS_ACK1_p & v8b229e | !BtoS_ACK1_p & v8af40b;
assign v8b140a = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v911e6a;
assign v8b2484 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v912699;
assign v8ae9f2 = BtoR_REQ1_p & v91261d | !BtoR_REQ1_p & v8b0a89;
assign v8aeead = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b1d03;
assign v911610 = RtoB_ACK0_p & v8af68d | !RtoB_ACK0_p & v8c66bb;
assign v911ed6 = jx1_p & v844f91 | !jx1_p & v8602f3;
assign v88e0ec = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v8ae745 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v911ed4;
assign v8b028f = BtoS_ACK7_p & v8b10fd | !BtoS_ACK7_p & v91245a;
assign v8afaa6 = BtoS_ACK0_p & v8afe4c | !BtoS_ACK0_p & v8b77ed;
assign v910f9a = RtoB_ACK0_p & v8af1ad | !RtoB_ACK0_p & v844f91;
assign v9123f6 = BtoS_ACK6_p & v9126de | !BtoS_ACK6_p & v8e98e4;
assign v8af253 = BtoR_REQ0_p & v912693 | !BtoR_REQ0_p & v8b29c1;
assign v8b2f6d = BtoS_ACK1_p & v912605 | !BtoS_ACK1_p & v8aea10;
assign v8c59a9 = StoB_REQ0_p & v8b28e6 | !StoB_REQ0_p & v8b0f51;
assign v8b07bc = RtoB_ACK0_p & v8af102 | !RtoB_ACK0_p & v844f91;
assign v8b2789 = BtoS_ACK2_p & v88709f | !BtoS_ACK2_p & v8aefe5;
assign v9126d5 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8b2bd9;
assign v8b1f50 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8c0456;
assign v8ae584 = jx0_p & v8b0bd4 | !jx0_p & !v9125d4;
assign v911fe4 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v9125eb;
assign v8af119 = jx0_p & v912617 | !jx0_p & !v86f3ae;
assign v8afa40 = BtoR_REQ1_p & v8b12e9 | !BtoR_REQ1_p & v8c6dfc;
assign v9123c1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8afc36;
assign v8af102 = jx2_p & v8aeec4 | !jx2_p & v8af886;
assign v8b2e07 = jx1_p & v8b2b91 | !jx1_p & !v91278f;
assign v8940f1 = DEQ_p & v91220c | !DEQ_p & v8b2633;
assign v89097b = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v912198;
assign v8b029e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v91239a;
assign v8aef7a = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v844f91;
assign v8b1f9c = jx2_p & v8aebc8 | !jx2_p & !v8b0c98;
assign v91243d = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b33af;
assign v8b1cbb = BtoS_ACK7_p & v8af431 | !BtoS_ACK7_p & v8cc1a9;
assign v9123f4 = RtoB_ACK0_p & v8dd6de | !RtoB_ACK0_p & v844f91;
assign v8b11b0 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85c0ac;
assign v8dd6de = jx2_p & v911a08 | !jx2_p & v8b25d9;
assign v9124a0 = BtoS_ACK0_p & v8c6cee | !BtoS_ACK0_p & v8ae4a3;
assign v8ae46b = jx1_p & v8b0e72 | !jx1_p & v8c5239;
assign v912186 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9123da;
assign v912543 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8af0fb;
assign v91258e = BtoS_ACK7_p & v88b300 | !BtoS_ACK7_p & v912690;
assign v91101e = RtoB_ACK1_p & v8afe84 | !RtoB_ACK1_p & v8f9630;
assign v912644 = jx3_p & v8af5ee | !jx3_p & !v8b3d1f;
assign v8b2a71 = jx0_p & v8ae4b3 | !jx0_p & v8c557b;
assign v912666 = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v8ae668;
assign v8b2b44 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fece1;
assign v912464 = StoB_REQ0_p & v8c568d | !StoB_REQ0_p & v912403;
assign v8aea95 = jx0_p & v8aff68 | !jx0_p & v9110f5;
assign v911f1c = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v87ba6d;
assign v8c54b4 = BtoS_ACK0_p & v8dd65f | !BtoS_ACK0_p & v8ae9bd;
assign v844f91 = 1;
assign v844fbb = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844f91;
assign v87cf4c = jx1_p & v8c65f8 | !jx1_p & v8b2ee4;
assign v91189f = StoB_REQ7_p & v8af094 | !StoB_REQ7_p & v8c4517;
assign v8b22c6 = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v85c0ac;
assign v8b2ac2 = jx0_p & v8b0d57 | !jx0_p & v9115b8;
assign v912662 = StoB_REQ2_p & v9124bd | !StoB_REQ2_p & v91248a;
assign v8aebc7 = BtoS_ACK3_p & v8afcf5 | !BtoS_ACK3_p & !v910e18;
assign v9126d2 = stateG7_1_p & v8b09f9 | !stateG7_1_p & v8b2a8c;
assign v8b232f = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8b085c;
assign v91180c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8af5f1;
assign v8b0b0c = StoB_REQ6_p & v8b0c94 | !StoB_REQ6_p & !v8ae6ab;
assign v911fab = RtoB_ACK0_p & v9126d1 | !RtoB_ACK0_p & v8b28d4;
assign v8ae898 = jx1_p & v911543 | !jx1_p & !v8b09ea;
assign v8b2d82 = StoB_REQ0_p & v911664 | !StoB_REQ0_p & v8b1d80;
assign v8ae934 = stateG7_1_p & v8c3926 | !stateG7_1_p & v9123f4;
assign v8af524 = jx0_p & v8b04ba | !jx0_p & v87ebfd;
assign v8afed8 = StoB_REQ6_p & v8b2345 | !StoB_REQ6_p & v91177e;
assign v8b02dd = stateG7_1_p & v8aeaf7 | !stateG7_1_p & v8aea93;
assign v911fb1 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b04f4;
assign v8b2ee4 = jx0_p & v8b2590 | !jx0_p & v8afcd6;
assign v9122c8 = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v8c5350;
assign v8c6e13 = DEQ_p & v8c53cf | !DEQ_p & v911eb1;
assign v9124db = jx2_p & v8dd632 | !jx2_p & v844f91;
assign v911fda = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8b076f;
assign BtoS_ACK3_n = !v8cc22c;
assign v88413b = BtoS_ACK6_p & v864227 | !BtoS_ACK6_p & v88d6cf;
assign v911de3 = BtoS_ACK7_p & v890ba5 | !BtoS_ACK7_p & v912326;
assign v8b0b24 = jx1_p & v912509 | !jx1_p & v8b0738;
assign v8b0cd4 = RtoB_ACK1_p & v8af102 | !RtoB_ACK1_p & v844f91;
assign v8b04fc = stateG7_1_p & v89209f | !stateG7_1_p & !v912598;
assign v911a08 = jx1_p & v844f91 | !jx1_p & v9123b6;
assign v8b1fee = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v88e0ec;
assign v91275a = BtoR_REQ1_p & v8af687 | !BtoR_REQ1_p & v8b02e9;
assign v88704a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c6167;
assign v8afabd = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911fb2;
assign v8aef67 = BtoR_REQ1_p & v911c9a | !BtoR_REQ1_p & v844f91;
assign v859e1d = jx0_p & v8e98f8 | !jx0_p & !v87a52a;
assign v911d22 = EMPTY_p & v8b2838 | !EMPTY_p & v9126e1;
assign v8b0151 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9124f0;
assign BtoS_ACK6_n = !v8c6e13;
assign v8b050b = StoB_REQ7_p & v9122d7 | !StoB_REQ7_p & v8b0b98;
assign v9125c3 = jx2_p & v8c3fe8 | !jx2_p & !v8b1d6c;
assign v8afdde = BtoS_ACK4_p & v8aef02 | !BtoS_ACK4_p & v9123ef;
assign v8afd2b = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c7305;
assign v91116e = RtoB_ACK0_p & v8b0994 | !RtoB_ACK0_p & v8b0a78;
assign v8b1003 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b1247;
assign v91183a = jx1_p & v8dd6ae | !jx1_p & !v887bd4;
assign v8b31b3 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v9123be;
assign v8b25d9 = jx1_p & v8dd6ad | !jx1_p & v85c13e;
assign v89223a = StoB_REQ6_p & v912568 | !StoB_REQ6_p & v8af949;
assign v844f9e = StoB_REQ4_n & v844f91 | !StoB_REQ4_n & !v844f91;
assign v911484 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8c4c30;
assign v861f8d = StoB_REQ6_p & v9116e8 | !StoB_REQ6_p & v8c704a;
assign v911291 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911b49;
assign v8c500e = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v912695;
assign v8b0cf9 = BtoR_REQ1_p & v8ae8c2 | !BtoR_REQ1_p & v912747;
assign v8bfa99 = StoB_REQ1_p & v8c3bd5 | !StoB_REQ1_p & v91231e;
assign v8579b7 = StoB_REQ2_p & v8c4b39 | !StoB_REQ2_p & v8c6bba;
assign v9110f5 = BtoS_ACK7_p & v911075 | !BtoS_ACK7_p & v8b3c24;
assign v8ae02e = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91269a;
assign v8c23d1 = BtoR_REQ0_p & v8c3e1b | !BtoR_REQ0_p & !v912600;
assign v9123cf = RtoB_ACK0_p & v910947 | !RtoB_ACK0_p & v8af102;
assign v8c043b = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8e5d84;
assign v9126fc = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v892ea3;
assign v8cda2f = RtoB_ACK1_p & v8b0994 | !RtoB_ACK1_p & v8b0a78;
assign v8dd6ff = DEQ_p & v8b107b | !DEQ_p & v8af756;
assign v88b1d7 = jx0_p & v8b1f0a | !jx0_p & !v8ae03c;
assign v8b8be1 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8af563;
assign v8cc0f3 = jx2_p & v8b2a8c | !jx2_p & v911fa0;
assign v8b2e27 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8ae519;
assign v8b32c1 = jx1_p & v8924fb | !jx1_p & !v9124e1;
assign v8c6bef = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8afdde;
assign v8e9896 = RtoB_ACK0_p & v88fa8c | !RtoB_ACK0_p & v8af102;
assign v876670 = BtoS_ACK0_p & v9123df | !BtoS_ACK0_p & v8c4c08;
assign v8b7791 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0119;
assign v9123ff = jx0_p & v912790 | !jx0_p & !v912666;
assign v88fef2 = jx0_p & v91269d | !jx0_p & v8c5357;
assign v8b1130 = BtoS_ACK6_p & v91265d | !BtoS_ACK6_p & v9126da;
assign v9111f5 = BtoR_REQ0_p & v91240f | !BtoR_REQ0_p & v912411;
assign v8b2267 = BtoS_ACK6_p & v911d4f | !BtoS_ACK6_p & v8c5bc3;
assign v910fe3 = stateG7_1_p & v8afbaa | !stateG7_1_p & v9123ca;
assign v890964 = jx3_p & v8aed6d | !jx3_p & v91240d;
assign v8b2c0d = RtoB_ACK0_p & v8909ff | !RtoB_ACK0_p & v844f91;
assign v912080 = BtoS_ACK7_p & v8af4ee | !BtoS_ACK7_p & v8b0753;
assign v912682 = stateG7_1_p & v910db7 | !stateG7_1_p & v8c3b67;
assign v9125b4 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8aebc4;
assign v88ffd6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8bfa12;
assign v8ae46d = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v912450;
assign v912456 = jx1_p & v8b2bee | !jx1_p & v844f91;
assign v8c510a = StoB_REQ7_p & v8b22be | !StoB_REQ7_p & v8b22c9;
assign v9124d5 = StoB_REQ2_p & v8afe33 | !StoB_REQ2_p & v844f91;
assign v8af83a = stateG7_1_p & v911ef0 | !stateG7_1_p & v890ac0;
assign v8c3619 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8fed5b;
assign v912326 = BtoS_ACK6_p & v890ba5 | !BtoS_ACK6_p & !v8b1de3;
assign v8c70dc = StoB_REQ0_p & v9125f8 | !StoB_REQ0_p & v844f91;
assign v911f83 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b02cb;
assign v8b29c9 = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v890a9a;
assign v911d4b = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8aeb91;
assign v8afe22 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8c0508;
assign v8af049 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v911d4b;
assign v87b54c = BtoS_ACK3_p & v8c050d | !BtoS_ACK3_p & v8ae0c6;
assign v8b02d5 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v88fa49;
assign v8afaec = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9115e4;
assign v8afd1f = jx1_p & v9126eb | !jx1_p & v8b241a;
assign v91250e = BtoS_ACK6_p & v8b03cf | !BtoS_ACK6_p & v9125cc;
assign v8b29af = StoB_REQ1_p & v91240c | !StoB_REQ1_p & v8aedf2;
assign v8c6c00 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v9123ef;
assign v8b0569 = jx3_p & v844f91 | !jx3_p & v8ae461;
assign v8aed35 = StoB_REQ7_p & v911052 | !StoB_REQ7_p & v8b1350;
assign v9110bb = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v890c16;
assign v912604 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b1e11;
assign v8b065b = jx1_p & v8ae584 | !jx1_p & !v8ae728;
assign v8c706b = jx0_p & v8dd5ff | !jx0_p & v8b028f;
assign v8af39f = jx1_p & v91271d | !jx1_p & v91253f;
assign v912714 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e943;
assign v9119bc = stateG12_p & v9125c3 | !stateG12_p & v8b2741;
assign v9114aa = jx0_p & v91242d | !jx0_p & v844f91;
assign v8b2493 = jx0_p & v912425 | !jx0_p & v8aed6d;
assign v8b2876 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v9124bd;
assign BtoS_ACK5_n = !v8dd6ff;
assign v8c4d14 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8bfaf2;
assign v8c23b9 = RtoB_ACK0_p & v8f9721 | !RtoB_ACK0_p & v8cf811;
assign v8c4a78 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b2479;
assign v89287e = jx0_p & v8c45be | !jx0_p & v844f91;
assign v8b0942 = FULL_p & v890b86 | !FULL_p & v8af2e3;
assign v8af1de = jx1_p & v844f91 | !jx1_p & v8c3d77;
assign v881ef0 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b0496;
assign v8b1350 = BtoS_ACK6_p & v91222a | !BtoS_ACK6_p & v912792;
assign v8aed6c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9124e0;
assign v8b2511 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & !v912771;
assign v8f96e9 = stateG7_1_p & v9125b4 | !stateG7_1_p & v91246b;
assign v8c0b46 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8c6df7;
assign v8aedc9 = StoB_REQ1_p & v9126f4 | !StoB_REQ1_p & v912394;
assign v912276 = BtoS_ACK0_p & v879d5b | !BtoS_ACK0_p & v911f49;
assign v8b31f9 = EMPTY_p & v8b33f2 | !EMPTY_p & v8b2a31;
assign v91243a = BtoR_REQ1_p & v88ac88 | !BtoR_REQ1_p & v8ae934;
assign v8b2aa2 = jx3_p & v844fb9 | !jx3_p & !v8af02f;
assign v8b09b4 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8b0dc1;
assign v8c3731 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8858cb;
assign v8af2c8 = jx2_p & v91100c | !jx2_p & v8ae898;
assign v8af9f2 = BtoS_ACK7_p & v8b33d3 | !BtoS_ACK7_p & v8c43ba;
assign v87de99 = FULL_p & v8af640 | !FULL_p & v8b2e31;
assign v8b2559 = jx2_p & v8b6d47 | !jx2_p & v912632;
assign v91174f = jx0_p & v911d44 | !jx0_p & v9123c8;
assign v8af864 = BtoS_ACK3_p & v8b2e66 | !BtoS_ACK3_p & !v9112e0;
assign v91246a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8aee49;
assign v8b11c5 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c4cc9;
assign v87b84a = RtoB_ACK0_p & v85f4b2 | !RtoB_ACK0_p & v8b02e9;
assign v8d50bc = DEQ_p & v8b1e0f | !DEQ_p & v911466;
assign v8c5d7e = jx1_p & v8cc0fb | !jx1_p & !v88b1d7;
assign v8b2f95 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f9b;
assign v8ae9bf = jx0_p & v912416 | !jx0_p & !v890c2c;
assign v87dc9f = jx1_p & v8ae6f2 | !jx1_p & !v911a2a;
assign v8c6aa0 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v9113eb;
assign v911ad5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b12f9;
assign v8b2569 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v9123ef;
assign v8af052 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8ae854;
assign v8ae7e5 = stateG7_1_p & v8c6c2f | !stateG7_1_p & v8b03c8;
assign v912783 = StoB_REQ6_p & v911695 | !StoB_REQ6_p & v8f965b;
assign v8b1ef8 = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v8c40af;
assign v8b2c5d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91245f;
assign v8b09ea = jx3_p & v844f91 | !jx3_p & !v911513;
assign v91244b = BtoS_ACK0_p & v8c6cee | !BtoS_ACK0_p & v9123e2;
assign v9123bd = jx0_p & v8f96c9 | !jx0_p & !v912415;
assign v8af9e6 = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v8b2655;
assign v8884e5 = jx0_p & v91258e | !jx0_p & v8c5357;
assign v912679 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8c0b07;
assign v911940 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c70dc;
assign v8af949 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v912432;
assign v91254d = BtoS_ACK7_p & v9126de | !BtoS_ACK7_p & v8c0acd;
assign v9123a2 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v9124e9;
assign v910ba7 = BtoS_ACK1_p & v879d5b | !BtoS_ACK1_p & v8b11a0;
assign v875d13 = jx1_p & v8aea95 | !jx1_p & v912761;
assign v8fecf2 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b0df4;
assign v8b1fc7 = StoB_REQ1_p & v8b139e | !StoB_REQ1_p & v8d6d2e;
assign v8af03f = BtoS_ACK2_p & v8b33a8 | !BtoS_ACK2_p & v8909b7;
assign v912420 = BtoR_REQ0_p & v8afdfc | !BtoR_REQ0_p & v8af960;
assign v8aed74 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8b0674;
assign v88b300 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v912702;
assign v89098b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b3c24;
assign v8b0d57 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v911bc6;
assign v8b244c = RtoB_ACK1_p & v9126c3 | !RtoB_ACK1_p & v911631;
assign v8b3d0c = StoB_REQ7_p & v8b1ec0 | !StoB_REQ7_p & v844f91;
assign v8b06d3 = StoB_REQ1_p & v8b6d3d | !StoB_REQ1_p & v912735;
assign v8dd5ec = RtoB_ACK1_p & v912402 | !RtoB_ACK1_p & v8b1e15;
assign v8af025 = stateG7_1_p & v8b2e7a | !stateG7_1_p & v8b0a89;
assign v8bfa1e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c3619;
assign v911ebd = stateG7_1_p & v8b0fab | !stateG7_1_p & v911fab;
assign v8c4c30 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9d;
assign v911a6a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fed10;
assign v890adc = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v912748;
assign v8b1166 = jx1_p & v8ae6f2 | !jx1_p & v844f91;
assign v912743 = StoB_REQ0_p & v8b1086 | !StoB_REQ0_p & !v844f91;
assign v8b2868 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8af717;
assign v8b0264 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9124c6;
assign v8b2d4a = BtoS_ACK3_p & v8b1c79 | !BtoS_ACK3_p & v8b290b;
assign v8b1ddf = RtoB_ACK0_p & v9123b1 | !RtoB_ACK0_p & v844f91;
assign v8b0b98 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v9126c8;
assign v91259b = jx1_p & v890ac0 | !jx1_p & v8b1245;
assign v8b2180 = jx0_p & v844f91 | !jx0_p & v8c5357;
assign v8d540a = BtoS_ACK6_p & v8c390a | !BtoS_ACK6_p & v8c4072;
assign v8af3e7 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v911f83;
assign v8b1c7b = jx3_p & v87a52a | !jx3_p & v890a73;
assign v8b21c9 = jx1_p & v8c49c6 | !jx1_p & v8af192;
assign v9126b9 = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v912660;
assign v912474 = BtoS_ACK6_p & v912609 | !BtoS_ACK6_p & v8c0443;
assign v9125b9 = jx0_p & v8af899 | !jx0_p & !v8b085e;
assign v911e94 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v912717;
assign v8fedea = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b24e9;
assign v9121a4 = BtoS_ACK6_p & v911a6a | !BtoS_ACK6_p & v8de9ca;
assign v88c831 = RtoB_ACK1_p & v8af68d | !RtoB_ACK1_p & v8c66bb;
assign v8b051e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8b0107;
assign v8c72da = BtoR_REQ0_p & v882969 | !BtoR_REQ0_p & v8afb03;
assign v8b0b7f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v912496;
assign v912733 = StoB_REQ3_p & v910e18 | !StoB_REQ3_p & !v844f91;
assign v8ba4a1 = jx0_p & v8b26af | !jx0_p & v8c3e7e;
assign v8b1fd2 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v9114f1;
assign v8aeab1 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b327a;
assign v911787 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b33a8;
assign v8b016c = BtoS_ACK7_p & v91259f | !BtoS_ACK7_p & v912716;
assign v8af68d = jx2_p & v8b3227 | !jx2_p & v8b336e;
assign v8aeaf7 = jx2_p & v8c42f9 | !jx2_p & v8af8b0;
assign v8b0611 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912652;
assign v8b2655 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & v8b1fee;
assign v86f3ae = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v8b076a;
assign v8b77ef = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8c66bb;
assign v8af683 = BtoS_ACK3_p & v88709f | !BtoS_ACK3_p & v8b2569;
assign v91263f = RtoB_ACK0_p & v885339 | !RtoB_ACK0_p & v8af02f;
assign v8c4b6c = stateG7_1_p & v8b244c | !stateG7_1_p & v911631;
assign v912416 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8b050b;
assign v8b0f2f = jx0_p & v912080 | !jx0_p & v8c3053;
assign v91278b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91253d;
assign v8b2b57 = StoB_REQ2_p & v87e29c | !StoB_REQ2_p & v8f9622;
assign v9124ed = BtoS_ACK4_p & v8b1f47 | !BtoS_ACK4_p & v912517;
assign v8afcf7 = BtoS_ACK7_p & v8c390a | !BtoS_ACK7_p & v911ea9;
assign v8f96c9 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8ae75b;
assign v9123fa = StoB_REQ2_p & v8b0283 | !StoB_REQ2_p & v8aebc7;
assign v8af98a = jx2_p & v8c48a8 | !jx2_p & v8b24af;
assign v8c5058 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8db1b1;
assign v8b2f44 = StoB_REQ6_p & v912547 | !StoB_REQ6_p & v8dd5d9;
assign v8af1d2 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v910cda;
assign v85a510 = BtoS_ACK6_p & v8af894 | !BtoS_ACK6_p & v8af275;
assign v8af0ef = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v8b7669;
assign v8ae5e2 = jx2_p & v8e5d29 | !jx2_p & v9115b8;
assign v8b2a9f = jx1_p & v844f91 | !jx1_p & v912485;
assign v8b0b83 = stateG7_1_p & v911411 | !stateG7_1_p & v912578;
assign v8b23d4 = jx1_p & v8c6a96 | !jx1_p & v8afdec;
assign v8ae162 = ENQ_p & v8b1161 | !ENQ_p & v8e98d2;
assign v911304 = BtoS_ACK7_p & v8b0661 | !BtoS_ACK7_p & v912114;
assign v8ae588 = RtoB_ACK1_p & v8b0a78 | !RtoB_ACK1_p & v844f91;
assign v9115b8 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912190;
assign v8c4cc9 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9125e2;
assign v8cc153 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v89085d;
assign v8c38b4 = StoB_REQ3_p & v912517 | !StoB_REQ3_p & v844f9f;
assign v8c4a57 = BtoS_ACK6_p & v91269a | !BtoS_ACK6_p & v910ff6;
assign v8aeeeb = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e990d;
assign v8c3bb7 = RtoB_ACK1_p & v8f9630 | !RtoB_ACK1_p & v8afe84;
assign v91255c = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8b232f;
assign v911466 = ENQ_p & v912280 | !ENQ_p & !v91268e;
assign v911fb6 = jx3_p & v87ebfd | !jx3_p & v8b0d99;
assign v8c50eb = RtoB_ACK1_p & v8b01bd | !RtoB_ACK1_p & v844f91;
assign v8cf811 = jx2_p & v8ae69b | !jx2_p & v910bd1;
assign v8b12ad = RtoB_ACK1_p & v8ae740 | !RtoB_ACK1_p & !v8b76f2;
assign v912756 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v9112ad;
assign v9124d8 = BtoR_REQ0_p & v8b05b7 | !BtoR_REQ0_p & v911792;
assign v8c5cc7 = jx1_p & v912698 | !jx1_p & v8b24cc;
assign v9123bb = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v911017;
assign v912518 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b7804;
assign v912591 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b11df;
assign v8b07f3 = jx2_p & v8b3d17 | !jx2_p & v8c5e4c;
assign v912576 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c568d;
assign v8db1b1 = StoB_REQ0_p & v911797 | !StoB_REQ0_p & v844f91;
assign v8afd55 = jx0_p & v8c6d04 | !jx0_p & !v911c25;
assign v8b2bee = jx0_p & v912617 | !jx0_p & v844f91;
assign v8afb51 = RtoB_ACK0_p & v8b0994 | !RtoB_ACK0_p & v844f91;
assign v8db180 = StoB_REQ0_p & v8ae64a | !StoB_REQ0_p & v8b06b8;
assign v9125d2 = jx0_p & v8b2878 | !jx0_p & v8b1e7d;
assign v8b33fa = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v912523;
assign v911d0e = jx2_p & v8784da | !jx2_p & v8c6e8e;
assign v8aea9f = StoB_REQ2_p & v9125ad | !StoB_REQ2_p & v8b2998;
assign v864227 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v881ef0;
assign v912415 = BtoS_ACK7_p & v8577c2 | !BtoS_ACK7_p & v8b1159;
assign v890ac7 = BtoS_ACK0_p & v8d6d04 | !BtoS_ACK0_p & v8b1e7b;
assign v912711 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912548;
assign v8af53c = BtoR_REQ1_p & v887acc | !BtoR_REQ1_p & v8c049b;
assign v8c458d = BtoS_ACK1_p & v8c0b8f | !BtoS_ACK1_p & v8b0fb9;
assign v911543 = jx0_p & v912617 | !jx0_p & !v8b1ef8;
assign v869876 = BtoS_ACK0_p & v8afe4c | !BtoS_ACK0_p & v9124be;
assign DEQ_n = !v8a8ba5;
assign v8af3b2 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9124ef;
assign v8909ff = jx2_p & v8af240 | !jx2_p & v864291;
assign v8b0738 = jx3_p & v8aed6d | !jx3_p & v8b2493;
assign v8c704b = stateG7_1_p & v912561 | !stateG7_1_p & v8af02f;
assign v912728 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v912679;
assign v911d44 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b073b;
assign v91257d = StoB_REQ6_p & v8c5845 | !StoB_REQ6_p & v844f91;
assign v912190 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9125e3;
assign v8b12f9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v87b5cf;
assign v8b2eed = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b03cf;
assign v8e98d6 = BtoS_ACK6_p & v8c390a | !BtoS_ACK6_p & v91244b;
assign v8b3382 = StoB_REQ7_p & v844f9d | !StoB_REQ7_p & v844f91;
assign v8b0945 = BtoR_REQ1_p & v887acc | !BtoR_REQ1_p & v9113da;
assign v8ae825 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8aefe5;
assign v91223a = StoB_REQ3_p & v912517 | !StoB_REQ3_p & v9124ed;
assign v8577c2 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8bfa8b;
assign v8b0dd0 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8b01bd;
assign v8aec8e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v911fb1;
assign v8c48c7 = jx0_p & v8c5192 | !jx0_p & v844f91;
assign v8af2bd = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v912400;
assign v911fa7 = jx0_p & v8bfa1e | !jx0_p & v8ae048;
assign v8b1dbd = StoB_REQ7_p & v8ae77f | !StoB_REQ7_p & v8b1130;
assign v9125a0 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9124c3;
assign v8b0d99 = jx0_p & v911304 | !jx0_p & v87ebfd;
assign v9126ab = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8b2629;
assign v91241f = StoB_REQ2_p & v8af683 | !StoB_REQ2_p & v844f91;
assign v8ae0c6 = StoB_REQ3_p & v8c44a1 | !StoB_REQ3_p & v8b1f47;
assign v8b2cc1 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b2998;
assign v8c568d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v911f54;
assign v8d6d2e = StoB_REQ2_p & v8b6482 | !StoB_REQ2_p & v8ae561;
assign v8e5d29 = jx1_p & v8b2ac2 | !jx1_p & v9115b8;
assign v8b6d7e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8e984d;
assign v8afa56 = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v8c3ea2;
assign v8b2838 = BtoR_REQ0_p & v8b1178 | !BtoR_REQ0_p & v85f3d2;
assign v8b2a8d = RtoB_ACK1_p & v8b0681 | !RtoB_ACK1_p & v844f91;
assign v8aec65 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b2173;
assign v887bda = BtoS_ACK0_p & v8b7804 | !BtoS_ACK0_p & v8b27a6;
assign v912600 = BtoR_REQ1_p & v8af0b5 | !BtoR_REQ1_p & !v844f91;
assign v8b1e6a = StoB_REQ2_p & v9119da | !StoB_REQ2_p & !v8e9920;
assign v91271b = BtoS_ACK7_p & v8b050c | !BtoS_ACK7_p & v8b12d5;
assign v8af02f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v844fb9;
assign v8b0eab = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b6d87;
assign v9123c7 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v91219b;
assign v91231e = StoB_REQ2_p & v8af2f9 | !StoB_REQ2_p & !v8c5356;
assign v9124c6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v9123ad;
assign v8c381a = BtoS_ACK4_p & v89217b | !BtoS_ACK4_p & v912517;
assign v8bfae8 = BtoS_ACK3_p & v8f9659 | !BtoS_ACK3_p & v8b339d;
assign v8b2639 = EMPTY_p & v8af066 | !EMPTY_p & v8b2e7b;
assign v8b0633 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9120ec;
assign v87e9d4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b2c07;
assign v887ac4 = RtoB_ACK1_p & v8ae956 | !RtoB_ACK1_p & v8af79f;
assign v8b2d17 = RtoB_ACK0_p & v912413 | !RtoB_ACK0_p & v912747;
assign v8b0c67 = StoB_REQ6_p & v8b0500 | !StoB_REQ6_p & v9123ad;
assign v9114dc = BtoS_ACK1_p & v8b034f | !BtoS_ACK1_p & v91244d;
assign v912442 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v912728;
assign v911fdf = RtoB_ACK0_p & v8b23d9 | !RtoB_ACK0_p & v8af98a;
assign v8b2bd8 = BtoS_ACK7_p & v8ae578 | !BtoS_ACK7_p & v8afb82;
assign v85915c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v9124b0;
assign v9126db = RtoB_ACK1_p & v911bf3 | !RtoB_ACK1_p & !v911f9c;
assign v86d734 = BtoS_ACK1_p & v879d5b | !BtoS_ACK1_p & v91241f;
assign v8b6f1f = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8aeddc;
assign v8b208f = StoB_REQ6_p & v9125cc | !StoB_REQ6_p & v844f91;
assign v8db23e = StoB_REQ3_p & v8b3321 | !StoB_REQ3_p & v844fb5;
assign v8c7049 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v89017d;
assign v8b12be = BtoR_REQ1_p & v8b788f | !BtoR_REQ1_p & v912698;
assign v912648 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v9125b2;
assign v8c6c4a = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v844f91;
assign v8af634 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f9d;
assign v911632 = BtoR_REQ1_p & v911bd2 | !BtoR_REQ1_p & v844f91;
assign v912547 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8fed1e;
assign v8b6e6f = stateG7_1_p & v912480 | !stateG7_1_p & v8afe84;
assign jx2_n = !v8b4ffd;
assign v8af79f = jx2_p & v9126b4 | !jx2_p & v8ae898;
assign v882eb7 = BtoR_REQ1_p & v8ae104 | !BtoR_REQ1_p & v8ae0da;
assign v8b251f = BtoS_ACK2_p & v88709f | !BtoS_ACK2_p & v9125ad;
assign v8bfa76 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8b8be1;
assign v883aaa = BtoS_ACK7_p & v8577c2 | !BtoS_ACK7_p & v8b1ffd;
assign v8c4a4e = jx0_p & v844f9b | !jx0_p & !v8b0750;
assign v8aeeaa = StoB_REQ0_p & v8ae745 | !StoB_REQ0_p & v911795;
assign v8ae728 = jx3_p & v8b76f1 | !jx3_p & v91230c;
assign v8b3357 = StoB_REQ2_p & v890c16 | !StoB_REQ2_p & !v9110bb;
assign v8c3fcf = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v88e856;
assign v8b09e6 = jx1_p & v844f91 | !jx1_p & !v8aeb57;
assign v9124bc = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v912769;
assign v912493 = BtoS_ACK6_p & v91222a | !BtoS_ACK6_p & v8b12fb;
assign v8b26bb = BtoS_ACK7_p & v8b2019 | !BtoS_ACK7_p & v8af463;
assign v9124c0 = StoB_REQ6_p & v911fe4 | !StoB_REQ6_p & v844f91;
assign v912479 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8af51f;
assign v8af318 = jx0_p & v844f9b | !jx0_p & !v844f91;
assign v8afa71 = jx2_p & v8b0e17 | !jx2_p & !v8b04b6;
assign v91261d = stateG7_1_p & v8b0a89 | !stateG7_1_p & v912737;
assign v8dd6bd = BtoS_ACK7_p & v890ba5 | !BtoS_ACK7_p & v9125d8;
assign v890b14 = EMPTY_p & v844f91 | !EMPTY_p & !v8af65e;
assign v9123a8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v912743;
assign v912563 = BtoS_ACK7_p & v8b050c | !BtoS_ACK7_p & v8afc08;
assign v9123cb = jx3_p & v844f91 | !jx3_p & v8b05a5;
assign v8b27ab = BtoR_REQ1_p & v8b65a3 | !BtoR_REQ1_p & v8af0c8;
assign v8af340 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b0b7f;
assign v856df0 = BtoR_REQ1_p & v8b039c | !BtoR_REQ1_p & !v8b0339;
assign v911e0c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0207;
assign v8cc0f1 = jx1_p & v8b2a71 | !jx1_p & v911538;
assign v8aeecd = BtoS_ACK1_p & v911787 | !BtoS_ACK1_p & v8af9cf;
assign v8c51e1 = StoB_REQ6_p & v91277e | !StoB_REQ6_p & v9123bb;
assign v911ed2 = BtoR_REQ1_p & v912643 | !BtoR_REQ1_p & v8afe84;
assign v8afa41 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v9124db;
assign v844fa0 = StoB_REQ5_n & v844f91 | !StoB_REQ5_n & !v844f91;
assign v8b77fb = jx2_p & v8b1166 | !jx2_p & !v8af095;
assign v8b2aad = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v911367;
assign v91129a = StoB_REQ5_n & v844f9f | !StoB_REQ5_n & !v844f91;
assign v89217c = jx0_p & v8b1003 | !jx0_p & v8b222c;
assign v91157d = stateG7_1_p & v8c66bb | !stateG7_1_p & v911610;
assign v890960 = jx2_p & v892fa2 | !jx2_p & v8aed6d;
assign v91119d = jx0_p & v8b1cbb | !jx0_p & v8afcf7;
assign v8af808 = BtoS_ACK0_p & v8b12af | !BtoS_ACK0_p & v8c4a3e;
assign v8fed43 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v9125eb;
assign v8b2019 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b0a55;
assign v8aec59 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v91266e;
assign v8af72b = BtoS_ACK0_p & v8dd65f | !BtoS_ACK0_p & v85c157;
assign v9124b5 = jx1_p & v8b032e | !jx1_p & !v887b1c;
assign v8afb18 = StoB_REQ6_p & v89092e | !StoB_REQ6_p & v8f965b;
assign v8c3ea2 = BtoS_ACK6_p & v91222a | !BtoS_ACK6_p & v9123e3;
assign v9124f8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8afce6;
assign v8b23de = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8b0d89;
assign v8c3afa = jx0_p & v911aa1 | !jx0_p & v844f91;
assign v8b1fcd = StoB_REQ2_p & v9124fe | !StoB_REQ2_p & v8b282e;
assign v912592 = BtoS_ACK3_p & v8c7026 | !BtoS_ACK3_p & v892ea4;
assign v911053 = stateG7_1_p & v8af02f | !stateG7_1_p & v91263f;
assign v8b0e17 = jx1_p & v8b2b80 | !jx1_p & v8c520c;
assign v890c50 = StoB_REQ6_p & v911ad5 | !StoB_REQ6_p & v8af72b;
assign v8e984d = StoB_REQ7_p & v9124c8 | !StoB_REQ7_p & v844f91;
assign v8b2f92 = BtoR_REQ0_p & v8c704b | !BtoR_REQ0_p & v8b0ebf;
assign v8ae925 = BtoS_ACK6_p & v8b33d3 | !BtoS_ACK6_p & v911219;
assign v8ae6c7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b26cf;
assign v8af9cf = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v912312;
assign v8af0e8 = BtoS_ACK7_p & v912432 | !BtoS_ACK7_p & v8b321d;
assign v9114e3 = RtoB_ACK0_p & v8b28d4 | !RtoB_ACK0_p & v8f9630;
assign v9125b6 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v912723;
assign v8e989e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b0b7a;
assign v8ae8d3 = BtoS_ACK6_p & v8dd6a6 | !BtoS_ACK6_p & v9123c1;
assign v8c3def = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v87d270;
assign v91278c = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & !v844f91;
assign v8b26ed = BtoS_ACK0_p & v8b1e22 | !BtoS_ACK0_p & v9126f5;
assign v911aa1 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v91255c;
assign v8c3efe = stateG7_1_p & v8e9842 | !stateG7_1_p & v9125b0;
assign v8b04ba = BtoS_ACK7_p & v8b0661 | !BtoS_ACK7_p & v8aef55;
assign v89017d = StoB_REQ0_p & v8aef95 | !StoB_REQ0_p & v911f83;
assign v8b2479 = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v9123e7;
assign v9123a3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v911219;
assign v8b24af = jx1_p & v912448 | !jx1_p & v844f91;
assign v8afe01 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v8c4a78;
assign v8c0ab9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844fb1;
assign v8c4353 = jx0_p & v8afb17 | !jx0_p & !v911c25;
assign v8b29e2 = jx0_p & v844f91 | !jx0_p & v8fecd9;
assign v8771a0 = jx0_p & v8b0485 | !jx0_p & !v8c64bf;
assign v91266e = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8ae516;
assign v8b0a78 = jx2_p & v8b09e6 | !jx2_p & v844f91;
assign v9116c4 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v9124fb;
assign v8b2576 = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v8aed7c;
assign v8c4398 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v8c3731;
assign v9125eb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v9112ad;
assign v8e98e4 = BtoS_ACK0_p & v8b12af | !BtoS_ACK0_p & v8b0e1d;
assign v8b2b5c = jx0_p & v8ae9fc | !jx0_p & v8c5e4c;
assign v8b25e8 = BtoS_ACK6_p & v844f9b | !BtoS_ACK6_p & v8aedf0;
assign v8890ee = jx0_p & v8b1d1e | !jx0_p & v863629;
assign v912408 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91130e;
assign v8c0b6f = BtoS_ACK0_p & v8db217 | !BtoS_ACK0_p & v912516;
assign v9124ce = jx0_p & v8aee85 | !jx0_p & v844f91;
assign v87cf6f = ENQ_p & v8af65e | !ENQ_p & !v890b14;
assign v8b0d58 = BtoS_ACK3_p & v91256c | !BtoS_ACK3_p & v912627;
assign v86c179 = StoB_REQ6_p & v9113eb | !StoB_REQ6_p & v91230e;
assign v8c520c = jx0_p & v8c426e | !jx0_p & v86ff66;
assign v8b0fb5 = BtoS_ACK7_p & v8ae878 | !BtoS_ACK7_p & v8b2911;
assign v8af9bd = BtoS_ACK2_p & v8f9614 | !BtoS_ACK2_p & !v8b22d1;
assign v91269f = StoB_REQ6_p & v8b238a | !StoB_REQ6_p & v88547b;
assign v9116c2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91159f;
assign v912705 = jx0_p & v911aa1 | !jx0_p & !v8c5d1c;
assign v8b05f1 = stateG7_1_p & v844f91 | !stateG7_1_p & v8b07bc;
assign v844fb1 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v8ae556 = StoB_REQ1_p & v888464 | !StoB_REQ1_p & v8b0e50;
assign v8b04d6 = BtoS_ACK4_p & v8aef02 | !BtoS_ACK4_p & v8b06bb;
assign v912698 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912711;
assign v8ae64c = BtoS_ACK1_p & v8afd76 | !BtoS_ACK1_p & v8b29af;
assign v8b0f57 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v9124b7;
assign v8b10c6 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8d6d16;
assign v8ae169 = BtoS_ACK2_p & v8b33a8 | !BtoS_ACK2_p & v8af7b2;
assign v8bfa8b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b0df4;
assign v8b2ad6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b2049;
assign v912625 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8ae437;
assign v8b0207 = StoB_REQ7_p & v912451 | !StoB_REQ7_p & v910fe2;
assign v8b1d1e = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b02d7;
assign v8c6964 = jx0_p & v8affe8 | !jx0_p & !v8c0b7c;
assign v887bcc = jx1_p & v8b25f8 | !jx1_p & v8b07d3;
assign v9125ae = jx3_p & v87ebfd | !jx3_p & v8af524;
assign v911795 = BtoS_ACK1_p & v8c0b8f | !BtoS_ACK1_p & v8b2cb5;
assign v8af518 = jx1_p & v8771a0 | !jx1_p & v91243f;
assign v911532 = stateG7_1_p & v8ae096 | !stateG7_1_p & v8b0994;
assign v8b0a36 = BtoR_REQ1_p & v8d14b5 | !BtoR_REQ1_p & v844f91;
assign v8b139e = StoB_REQ2_p & v8b6482 | !StoB_REQ2_p & v912788;
assign v91245f = BtoS_ACK0_p & v8db217 | !BtoS_ACK0_p & v8c23d2;
assign v911a5d = BtoS_ACK0_p & v8b7892 | !BtoS_ACK0_p & v8b099d;
assign v8b1eff = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9112ad;
assign v8b0fac = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8b2d5a;
assign v9126a1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8af808;
assign v8aebd0 = StoB_REQ1_p & v8b29d8 | !StoB_REQ1_p & v8b2b57;
assign v91272b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b08b3;
assign v890be4 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b0151;
assign v91248b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8ae47c;
assign v91275f = jx1_p & v8aea95 | !jx1_p & v8cc202;
assign v8b0358 = BtoR_REQ0_p & v8aee79 | !BtoR_REQ0_p & v894810;
assign v9126b2 = StoB_REQ6_p & v8c0456 | !StoB_REQ6_p & v893433;
assign v88b60c = jx0_p & v9126c9 | !jx0_p & !v8ae92f;
assign v912694 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v912068;
assign v912525 = StoB_REQ2_p & v8b0fee | !StoB_REQ2_p & v91255d;
assign v8b3d17 = jx1_p & v87cfd0 | !jx1_p & v8b2b5c;
assign v89217b = StoB_REQ4_p & v912517 | !StoB_REQ4_p & !v844f91;
assign v8b52c1 = RtoB_ACK0_p & v912122 | !RtoB_ACK0_p & v8b01bd;
assign v87a52a = BtoS_ACK7_p & v8b0260 | !BtoS_ACK7_p & v8f9632;
assign v912532 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8aef95;
assign v8b2d92 = StoB_REQ6_p & v8b0500 | !StoB_REQ6_p & v9115fc;
assign v892555 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v876670;
assign v8ae6f2 = jx0_p & v8b0485 | !jx0_p & v844f91;
assign v8b0d88 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8c3bd5;
assign v8872e8 = BtoS_ACK6_p & v911bad | !BtoS_ACK6_p & v9123f7;
assign v9124fe = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8b339d;
assign v912467 = jx1_p & v8771a0 | !jx1_p & v8c6964;
assign v8dd5e6 = jx3_p & v844f91 | !jx3_p & v911fad;
assign v87d0f8 = EMPTY_p & v8b2792 | !EMPTY_p & v88abf5;
assign v8af92f = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8dd654;
assign v9123d1 = StoB_REQ7_p & v8af916 | !StoB_REQ7_p & !v844f91;
assign v912401 = jx0_p & v8db20a | !jx0_p & v911e0c;
assign v8af2b1 = jx1_p & v88acc3 | !jx1_p & v8b32b6;
assign v8e9842 = jx2_p & v91161f | !jx2_p & v9113a8;
assign v9125d9 = jx1_p & v911d0d | !jx1_p & v890964;
assign v912521 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8c77fe;
assign v8b01a4 = RtoB_ACK1_p & v8b23d9 | !RtoB_ACK1_p & v8af1ad;
assign v9119da = BtoS_ACK3_p & v8b00f2 | !BtoS_ACK3_p & v8b0d0e;
assign v8b216f = BtoS_ACK7_p & v911bad | !BtoS_ACK7_p & v8b0642;
assign v912556 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8f9625;
assign v91242f = jx0_p & v8b09b4 | !jx0_p & !v8c0b7c;
assign v8af27d = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8f9614;
assign v8af6c8 = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v8b2019;
assign v892ea3 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8aec57;
assign v91259f = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8dd6a6;
assign v912692 = jx0_p & v91151f | !jx0_p & !v89098b;
assign v910ca3 = BtoS_ACK0_p & v8b7804 | !BtoS_ACK0_p & v8bb768;
assign v911b4f = jx0_p & v8b1e91 | !jx0_p & v8ae7a9;
assign v912790 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8b2c68;
assign v9126d9 = jx2_p & v8b2ab3 | !jx2_p & v8b21c9;
assign v8ae6e0 = jx1_p & v8afbd6 | !jx1_p & v844f91;
assign v8b0936 = BtoR_REQ1_p & v8fed49 | !BtoR_REQ1_p & v8afc85;
assign v91276f = StoB_REQ0_p & v912604 | !StoB_REQ0_p & v844f91;
assign v9110c2 = jx1_p & v910c69 | !jx1_p & v912698;
assign v863629 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8affb3;
assign v8c5bc3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9123c9;
assign v8b76f2 = jx2_p & v9126f9 | !jx2_p & v8c498b;
assign v91180b = jx0_p & v873367 | !jx0_p & !v8b25a2;
assign v912496 = StoB_REQ1_p & v8afe49 | !StoB_REQ1_p & v844f91;
assign v8af451 = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v8affdf;
assign v912718 = RtoB_ACK1_p & v912122 | !RtoB_ACK1_p & v8b01bd;
assign v887c3b = BtoR_REQ0_p & v8b077d | !BtoR_REQ0_p & v8b0cf9;
assign v8b2590 = BtoS_ACK7_p & v8ae4e9 | !BtoS_ACK7_p & v8b0062;
assign v8cc139 = FULL_p & v912420 | !FULL_p & v890880;
assign v8c0435 = jx2_p & v8ae7ea | !jx2_p & !v9123fe;
assign v8dd6fe = RtoB_ACK0_p & v890960 | !RtoB_ACK0_p & v8b0994;
assign v8fed1e = StoB_REQ0_p & v88ef39 | !StoB_REQ0_p & v844f91;
assign v8c5e54 = BtoS_ACK0_p & v8c0b8f | !BtoS_ACK0_p & v8c4b37;
assign v91151a = BtoR_REQ0_p & v85c164 | !BtoR_REQ0_p & v85c0bd;
assign v8b2a31 = stateG12_p & v8b0bd2 | !stateG12_p & v8b33f2;
assign v8c6dff = RtoB_ACK1_p & v8c3cff | !RtoB_ACK1_p & v9126d9;
assign v8c6caf = jx0_p & v91248b | !jx0_p & v8bb97f;
assign v91268d = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v890be4;
assign v8b2cb5 = StoB_REQ2_p & v8b03fc | !StoB_REQ2_p & v91251d;
assign v91215f = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v912487;
assign v9125fc = stateG7_1_p & v8c3bb7 | !stateG7_1_p & v912046;
assign v8b09b9 = stateG7_1_p & v911220 | !stateG7_1_p & v8b1e0b;
assign v8940a8 = jx0_p & v8cc153 | !jx0_p & v844f91;
assign v8b070e = BtoR_REQ0_p & v86ce5c | !BtoR_REQ0_p & v911e1d;
assign v8cc1a9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b2843;
assign v8596e1 = StoB_REQ2_p & v8b0283 | !StoB_REQ2_p & v88331f;
assign v8c7153 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b016b;
assign v912752 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & !v911e40;
assign v8ae437 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c4398;
assign v8b1083 = StoB_REQ0_p & v87cf71 | !StoB_REQ0_p & v844f91;
assign v912617 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8b1fd2;
assign v912747 = jx2_p & v91247c | !jx2_p & !v91257a;
assign v9124a4 = jx2_p & v9123d2 | !jx2_p & v8b236d;
assign v911fae = stateG7_1_p & v8af618 | !stateG7_1_p & v844f91;
assign v8ae805 = StoB_REQ2_p & v8b1ea2 | !StoB_REQ2_p & v8db139;
assign v9116e0 = BtoR_REQ1_p & v8b0648 | !BtoR_REQ1_p & v844f91;
assign v85e7ac = StoB_REQ6_p & v8b2815 | !StoB_REQ6_p & v844f91;
assign v86995b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v890adc;
assign v8af159 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9112ad;
assign v910c9d = BtoS_ACK0_p & v8b0df4 | !BtoS_ACK0_p & v8bfa8b;
assign v9126f5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b2c6b;
assign v8af55a = jx0_p & v8af82e | !jx0_p & !v8c39b8;
assign v9125cc = BtoS_ACK0_p & v91244d | !BtoS_ACK0_p & v890bdc;
assign v8b04f8 = RtoB_ACK0_p & v8ae740 | !RtoB_ACK0_p & !v9123b1;
assign v8b1eeb = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v890bcb;
assign v8b2610 = jx2_p & v844fbb | !jx2_p & v9126c6;
assign v8af036 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b21bb;
assign v8c3541 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v869f57;
assign v911f72 = jx3_p & v844f91 | !jx3_p & !v9125d2;
assign v8b209b = BtoS_ACK6_p & v8c390a | !BtoS_ACK6_p & v8b1fc5;
assign v8fecb7 = jx0_p & v8c4189 | !jx0_p & v8af3b2;
assign v8aeb67 = jx0_p & v8afab8 | !jx0_p & !v844f9d;
assign v912631 = BtoS_ACK0_p & v8db217 | !BtoS_ACK0_p & v912543;
assign v912568 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8af36f;
assign v89286e = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v8b13f6;
assign v890930 = StoB_REQ6_p & v911539 | !StoB_REQ6_p & v844f91;
assign v8b0ae4 = RtoB_ACK1_p & v8b13ca | !RtoB_ACK1_p & v88acc3;
assign v87d0a9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b0705;
assign v911f9d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8ae516;
assign v9126d8 = jx1_p & v9126eb | !jx1_p & v91264e;
assign v912658 = jx1_p & v8ae6f2 | !jx1_p & !v9114aa;
assign v8c4a3e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b27f9;
assign v91239a = BtoS_ACK1_p & v8b07c0 | !BtoS_ACK1_p & v91272f;
assign v8c426f = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v8af918;
assign v9126c9 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8aefc1;
assign v8b74aa = BtoR_REQ0_p & v9123d6 | !BtoR_REQ0_p & v8b0936;
assign v912470 = BtoR_REQ1_p & v8bfa4c | !BtoR_REQ1_p & v8b19b1;
assign v911bd2 = stateG7_1_p & v8b2000 | !stateG7_1_p & v912664;
assign v8e98f8 = BtoS_ACK7_p & v844f95 | !BtoS_ACK7_p & !v8c7153;
assign v91277b = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v9126f4;
assign v8b0b70 = stateG7_1_p & v9117c1 | !stateG7_1_p & !v844f91;
assign v8af73a = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b26ed;
assign v9125e8 = BtoS_ACK7_p & v8c390a | !BtoS_ACK7_p & v8ae673;
assign v8ae6f0 = jx0_p & v8ae4b3 | !jx0_p & !v844f91;
assign v911a8d = stateG7_1_p & v8b0cd4 | !stateG7_1_p & v844f91;
assign v9123af = StoB_REQ4_p & v912517 | !StoB_REQ4_p & v844f9f;
assign v9122e7 = jx1_p & v8b0e72 | !jx1_p & v8b068b;
assign v8b0ef5 = jx3_p & v844f91 | !jx3_p & v8b05ce;
assign v910e34 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8aecf5;
assign v911bdc = RtoB_ACK1_p & v8b0eb6 | !RtoB_ACK1_p & v911196;
assign v8b2df8 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v9126ae;
assign v9115ca = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b3382;
assign v85c0ac = StoB_REQ3_p & v9123ef | !StoB_REQ3_p & v844f91;
assign v910e18 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & !v844f91;
assign v844f9d = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v844f91;
assign v9113eb = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v91277b;
assign v8c6c18 = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v91189f;
assign v912264 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v912450;
assign v8b2eb4 = BtoS_ACK7_p & v8b0661 | !BtoS_ACK7_p & v8af78e;
assign v8af2f9 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v91265a;
assign v9123be = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9126f5;
assign v8c6cae = jx0_p & v8b08c4 | !jx0_p & v91256e;
assign v8c23d2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9125d7;
assign v911fcd = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8feced;
assign v912423 = BtoR_REQ0_p & v8b04fc | !BtoR_REQ0_p & !v91144e;
assign v8e9855 = jx2_p & v8ae7ea | !jx2_p & !v8b32c1;
assign v88b998 = BtoS_ACK6_p & v8b03cf | !BtoS_ACK6_p & v912750;
assign v888766 = BtoS_ACK7_p & v912432 | !BtoS_ACK7_p & v8aec65;
assign v912702 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v912487;
assign v8ae02f = jx1_p & v8b2df3 | !jx1_p & v8c3e60;
assign v8b2bbf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8827a3;
assign v8b2e24 = jx1_p & v91271d | !jx1_p & v91267e;
assign v8b1161 = EMPTY_p & v9126d5 | !EMPTY_p & v9121d1;
assign v9123fe = jx1_p & v8924fb | !jx1_p & !v911f72;
assign v911158 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8b24b7;
assign v910bbe = RtoB_ACK0_p & v91270f | !RtoB_ACK0_p & v912698;
assign v911fc2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911797;
assign v8b077d = stateG7_1_p & v91134e | !stateG7_1_p & v912747;
assign v8e9961 = DEQ_p & v912537 | !DEQ_p & v910d87;
assign v8afb03 = BtoR_REQ1_p & v8fed7c | !BtoR_REQ1_p & v844f91;
assign v91185f = BtoS_ACK7_p & v9124fd | !BtoS_ACK7_p & v8af049;
assign v8af095 = jx1_p & v8940a8 | !jx1_p & v844f91;
assign v8692ec = StoB_REQ2_p & v912068 | !StoB_REQ2_p & v912694;
assign v8b279b = BtoS_ACK0_p & v844f9e | !BtoS_ACK0_p & v911fdd;
assign v911714 = jx1_p & v859e1d | !jx1_p & !v8ae8e8;
assign v8742de = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v912414;
assign v8b05b0 = BtoS_ACK6_p & v912702 | !BtoS_ACK6_p & v912752;
assign v87ebfd = BtoS_ACK7_p & v8b0661 | !BtoS_ACK7_p & v8b2911;
assign v8c0a62 = RtoB_ACK1_p & v8af1a2 | !RtoB_ACK1_p & v844f91;
assign v8b2629 = StoB_REQ6_p & v8af3e7 | !StoB_REQ6_p & v8c7049;
assign v8b27a6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c0b90;
assign v8b01dd = ENQ_p & v8b0b63 | !ENQ_p & v8b1f58;
assign v8b101c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b20fa;
assign v8af767 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v912568;
assign v91171d = StoB_REQ0_p & v91251c | !StoB_REQ0_p & v844f91;
assign v91230e = BtoS_ACK0_p & v8af918 | !BtoS_ACK0_p & v8b0a2d;
assign v8c45e8 = jx0_p & v912181 | !jx0_p & v8c0bc2;
assign v8aede2 = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v9126df;
assign v8b1de3 = StoB_REQ0_p & v9112ad | !StoB_REQ0_p & !v844f91;
assign v8c40af = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8db1d7;
assign v8b1e22 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v8b09fb = jx2_p & v8b1166 | !jx2_p & v844f91;
assign v8b038f = StoB_REQ2_p & v8b6482 | !StoB_REQ2_p & v8b02d5;
assign v8c6cb4 = jx0_p & v87ebfd | !jx0_p & v8c41af;
assign v8c0bf1 = BtoS_ACK0_p & v8b327a | !BtoS_ACK0_p & v91273c;
assign v910ff3 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v8c0ab9;
assign v887bd4 = jx3_p & v844f91 | !jx3_p & v912502;
assign v881e63 = jx0_p & v90c2e3 | !jx0_p & v844f91;
assign v8af51f = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v91254f;
assign v8b02e9 = jx2_p & v912331 | !jx2_p & !v8b0467;
assign v8b1e9a = BtoR_REQ1_p & v8c4b6c | !BtoR_REQ1_p & v844f91;
assign v8b0b63 = EMPTY_p & v8b1ca6 | !EMPTY_p & v9126ff;
assign v8a8ba5 = DEQ_p & v844f91 | !DEQ_p & !v87cf6f;
assign v8b0e57 = BtoS_ACK2_p & v8924d2 | !BtoS_ACK2_p & v8af9e8;
assign v911e03 = ENQ_p & v8b252f | !ENQ_p & !v8afdb9;
assign v8afb96 = BtoS_ACK7_p & v91259f | !BtoS_ACK7_p & v8b091d;
assign v8c6dfc = stateG7_1_p & v912490 | !stateG7_1_p & v910f9a;
assign v8b0661 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8ae878;
assign v8afdfc = stateG7_1_p & v8b0d4e | !stateG7_1_p & v844f91;
assign v8c390a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c6cee;
assign v8b1406 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v91274b;
assign v911692 = StoB_REQ6_p & v910ca3 | !StoB_REQ6_p & v844f91;
assign v911f38 = StoB_REQ2_p & v8aefa4 | !StoB_REQ2_p & v8c6c56;
assign v8b1d71 = BtoS_ACK7_p & v911149 | !BtoS_ACK7_p & v892551;
assign v8af748 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v85e7ac;
assign v912411 = BtoR_REQ1_p & v87dbe0 | !BtoR_REQ1_p & v911e65;
assign v912681 = BtoS_ACK0_p & v9123df | !BtoS_ACK0_p & v8afabd;
assign v8cc108 = RtoB_ACK1_p & v8af02f | !RtoB_ACK1_p & v911289;
assign v8de9ca = StoB_REQ6_p & v911197 | !StoB_REQ6_p & v866ac1;
assign v9125b3 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9118e7;
assign v912453 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8c4b39;
assign v8b0e1d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911fcd;
assign v8f953d = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v890246;
assign v8b252f = EMPTY_p & v844fbb | !EMPTY_p & v9123a9;
assign v8c7100 = jx3_p & v911c7e | !jx3_p & v8b2a8c;
assign v8afea2 = BtoS_ACK6_p & v8dd6a6 | !BtoS_ACK6_p & v8aeb4c;
assign v91238f = RtoB_ACK0_p & v911e3b | !RtoB_ACK0_p & v8b23d9;
assign v890bdc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v9114dc;
assign v869205 = jx3_p & v844f91 | !jx3_p & !v844f91;
assign v8af77e = BtoS_ACK1_p & v8af27d | !BtoS_ACK1_p & v8af2f5;
assign v91275d = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8ae446;
assign v912638 = BtoS_ACK0_p & v8f9617 | !BtoS_ACK0_p & v8b0be4;
assign v88340e = RtoB_ACK1_p & v8b0994 | !RtoB_ACK1_p & v844f91;
assign v9121e7 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v912549;
assign v9122d7 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8b20ab;
assign v9123f5 = jx0_p & v912796 | !jx0_p & v8b0611;
assign v8b340c = StoB_REQ3_p & v912517 | !StoB_REQ3_p & v844f91;
assign v910efa = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b1195;
assign v8b2fbc = RtoB_ACK0_p & v8afe84 | !RtoB_ACK0_p & v8f9630;
assign v911e40 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v912683;
assign v8dd5e2 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8e992f;
assign v8af586 = jx0_p & v8c3fcf | !jx0_p & v9125c8;
assign v8aec85 = BtoS_ACK1_p & v912605 | !BtoS_ACK1_p & v8b1fc7;
assign v9123d6 = stateG7_1_p & v8b1110 | !stateG7_1_p & v8c6979;
assign v8c0aef = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8ae4ce;
assign v91255d = BtoS_ACK3_p & v8ae041 | !BtoS_ACK3_p & v8ae713;
assign v91243e = jx0_p & v8c53ab | !jx0_p & v844f91;
assign v911fd6 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8af683;
assign v8c4410 = BtoS_ACK7_p & v8bfa8b | !BtoS_ACK7_p & v8b09a9;
assign v911772 = jx0_p & v911fd9 | !jx0_p & !v8b2576;
assign v8fed49 = stateG7_1_p & v8c6979 | !stateG7_1_p & v8b7802;
assign v91271c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v91266e;
assign v912569 = BtoR_REQ0_p & v911a59 | !BtoR_REQ0_p & v8803b6;
assign v8b1e43 = jx3_p & v9124c2 | !jx3_p & v8b2a8c;
assign v8af78e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ae5c0;
assign v9125a8 = BtoS_ACK6_p & v911a6a | !BtoS_ACK6_p & v912634;
assign v912432 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v844f91;
assign v87bd1c = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8b0681;
assign v911959 = StoB_REQ6_p & v8b232f | !StoB_REQ6_p & v8c704a;
assign v8af415 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c6cdc;
assign v8b8e79 = BtoS_ACK7_p & v8c6c4a | !BtoS_ACK7_p & v911e68;
assign v8afb09 = jx0_p & v912796 | !jx0_p & v9115ca;
assign v8ae519 = StoB_REQ0_p & v8afc68 | !StoB_REQ0_p & v912797;
assign v8aed7c = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v912492;
assign v8f9617 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v8afd76;
assign v911fa0 = jx1_p & v8b2a8c | !jx1_p & v8b1e43;
assign v8aee21 = StoB_REQ2_p & v8f9625 | !StoB_REQ2_p & v844f91;
assign v9115c6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8c0443;
assign v91263e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8aff15;
assign v9121ee = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b52f7;
assign v8b0e50 = StoB_REQ2_p & v8bfae8 | !StoB_REQ2_p & v9116aa;
assign v8b05a5 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b2911;
assign v8dd667 = jx3_p & v844f91 | !jx3_p & !v8c4353;
assign v8b3350 = jx0_p & v8c6d04 | !jx0_p & v844f91;
assign v8af5fe = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b71c1;
assign v8afb8e = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8b0a78;
assign v912685 = jx0_p & v911d44 | !jx0_p & v8c3541;
assign v9113d6 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8af72b;
assign v8c3d52 = BtoR_REQ0_p & v8db1c7 | !BtoR_REQ0_p & v8c47c3;
assign v9126d1 = jx2_p & v8b2f46 | !jx2_p & v91183a;
assign v9126b1 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8af6c8;
assign v8ae740 = jx2_p & v8b066c | !jx2_p & !v8ae02f;
assign v8b2e60 = jx0_p & v844f91 | !jx0_p & v87a52a;
assign v8dd5ca = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v892511;
assign v8ae8b7 = BtoR_REQ1_p & v8b0c90 | !BtoR_REQ1_p & v8b09a3;
assign v8affdf = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85afd4;
assign v912742 = jx1_p & v8b2bee | !jx1_p & !v8dd5e6;
assign v8ae722 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b2fc4;
assign v911149 = StoB_REQ6_p & v844f9f | !StoB_REQ6_p & v91222a;
assign v912775 = jx3_p & v844f91 | !jx3_p & v8c3c57;
assign v8b3227 = jx1_p & v91180b | !jx1_p & v8e9852;
assign v911e68 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8bfab2;
assign v8aff68 = BtoS_ACK7_p & v8b33d3 | !BtoS_ACK7_p & v8b3c24;
assign v8b085e = BtoS_ACK7_p & v8b0e3d | !BtoS_ACK7_p & v9114cd;
assign v8b002e = jx1_p & v8b0f2f | !jx1_p & v911fc3;
assign v912529 = RtoB_ACK0_p & v8afde2 | !RtoB_ACK0_p & v890ac0;
assign v91222a = StoB_REQ0_p & v844f9f | !StoB_REQ0_p & v8f9617;
assign v894087 = BtoS_ACK0_p & v8c0b8f | !BtoS_ACK0_p & v8af7f1;
assign v8b0dd4 = StoB_REQ7_p & v8af168 | !StoB_REQ7_p & v844f91;
assign v8b07a1 = jx0_p & v8ae4b3 | !jx0_p & v8b25a2;
assign v86cbb8 = BtoS_ACK2_p & v8924d2 | !BtoS_ACK2_p & v8b2c21;
assign v8ae60e = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v912527;
assign v8c5781 = stateG7_1_p & v8ae582 | !stateG7_1_p & v9115b8;
assign v8b11c4 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91276a;
assign v8af52b = BtoS_ACK7_p & v8ae578 | !BtoS_ACK7_p & v912542;
assign v8ae887 = jx2_p & v8afa3c | !jx2_p & !v8b32c1;
assign v911538 = jx0_p & v9115c7 | !jx0_p & v8b0611;
assign v887ae1 = BtoS_ACK6_p & v8c6c4a | !BtoS_ACK6_p & v8b2f44;
assign v8b7443 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v912264;
assign v8b0648 = stateG7_1_p & v8dd5ec | !stateG7_1_p & v911fac;
assign v8b2df3 = jx0_p & v8c09de | !jx0_p & v8b11ef;
assign v8b0bd4 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8b25e8;
assign v8af215 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8b2353;
assign v8ae074 = jx0_p & v91115b | !jx0_p & v9115ca;
assign v8c5404 = BtoS_ACK6_p & v8ae578 | !BtoS_ACK6_p & v87a09b;
assign v8b648c = jx0_p & v91240a | !jx0_p & !v844f9d;
assign v9123eb = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8b2fd3;
assign v91241a = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & v8b01bd;
assign v890940 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fecf2;
assign v9123e0 = BtoR_REQ1_p & v8b788f | !BtoR_REQ1_p & v8b2a2e;
assign v9032d6 = BtoS_ACK3_p & v8c050d | !BtoS_ACK3_p & v8b1154;
assign v8af71d = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8af767;
assign v8ae561 = BtoS_ACK2_p & v8aef7a | !BtoS_ACK2_p & v8c6e5a;
assign v8ae8c2 = stateG7_1_p & v912747 | !stateG7_1_p & v8b2d17;
assign v8c0b90 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v8b7804;
assign v8b3399 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8924ff;
assign v912575 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b3d12;
assign v8b321d = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b3320;
assign v8afd31 = RtoB_ACK1_p & v887bcf | !RtoB_ACK1_p & v8ae9f4;
assign v8b10bf = RtoB_ACK0_p & v8b0681 | !RtoB_ACK0_p & v844f91;
assign v912776 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v912532;
assign v8dd5d6 = jx0_p & v91272b | !jx0_p & v8b2afc;
assign v8ae487 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b04d6;
assign v8b0626 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9125a5;
assign v911017 = StoB_REQ0_p & v8b0d88 | !StoB_REQ0_p & v8b21fa;
assign v8af765 = StoB_REQ6_p & v8b20ab | !StoB_REQ6_p & v87b940;
assign v8ae118 = BtoS_ACK6_p & v91269a | !BtoS_ACK6_p & v8b2e17;
assign v8b2aeb = StoB_REQ7_p & v89092e | !StoB_REQ7_p & v910fe2;
assign v9125ab = jx3_p & v8c5357 | !jx3_p & v8884e5;
assign v8af399 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v861315;
assign v8c49c6 = jx0_p & v8ae88e | !jx0_p & v8c3e7e;
assign v91260b = BtoS_ACK2_p & v8f9614 | !BtoS_ACK2_p & v8b2a3e;
assign v911dbd = jx0_p & v91272b | !jx0_p & v911633;
assign v8b09a9 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9122c8;
assign v8b22be = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8f9587;
assign v8c4c08 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8e9903;
assign v9123c6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91157e;
assign v8af452 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v912709;
assign v8ae696 = jx2_p & v910cab | !jx2_p & v912632;
assign v912766 = StoB_REQ6_p & v911197 | !StoB_REQ6_p & v88d6cf;
assign v85d63e = jx0_p & v8b004c | !jx0_p & v844f91;
assign v9126b8 = jx0_p & v8b09b4 | !jx0_p & !v8591f3;
assign v91277e = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8b0d88;
assign v8b29ed = BtoR_REQ0_p & v911ebd | !BtoR_REQ0_p & v8b27ab;
assign v8b2b08 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v912517;
assign v911d7e = BtoS_ACK0_p & v879d5b | !BtoS_ACK0_p & v912182;
assign v8b28c6 = BtoS_ACK0_p & v8b7804 | !BtoS_ACK0_p & v8b2b44;
assign v9116aa = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8b339d;
assign v8c568f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b2ddd;
assign v892501 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v89288a;
assign v8b29d9 = BtoR_REQ0_p & v8b6e6f | !BtoR_REQ0_p & v8b0ae9;
assign v9124e7 = stateG7_1_p & v8c45bc | !stateG7_1_p & v8c0aef;
assign v8b0823 = ENQ_p & v8af92f | !ENQ_p & v91187a;
assign v8ae668 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8b2484;
assign v8aecf5 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & v9123ef;
assign v8b246f = BtoS_ACK7_p & v8b10cf | !BtoS_ACK7_p & v8d6cda;
assign v9112ad = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v8d6d2c = BtoR_REQ0_p & v8b039c | !BtoR_REQ0_p & !v87cd98;
assign v8c6e2e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v911fd1;
assign v8b0584 = stateG7_1_p & v87bd1c | !stateG7_1_p & v8af7cb;
assign v8e994b = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v911ef8;
assign v8af899 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8c510a;
assign v8c39b8 = BtoS_ACK7_p & v8b33d3 | !BtoS_ACK7_p & v8b029c;
assign v844fa7 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844f91;
assign v8b02ab = jx1_p & v88fef2 | !jx1_p & v91119d;
assign v911be0 = jx0_p & v8af564 | !jx0_p & v911914;
assign v9125dd = stateG7_1_p & v8afd31 | !stateG7_1_p & v844f91;
assign v8c6df7 = StoB_REQ6_p & v8b0674 | !StoB_REQ6_p & v8af399;
assign v9126c6 = jx1_p & v844fbb | !jx1_p & !v911fa4;
assign v8c0acd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v9123f6;
assign v91253d = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v8d6d1f;
assign v912709 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8b034f;
assign jx3_n = v8d50bc;
assign v912763 = StoB_REQ3_p & v9124ed | !StoB_REQ3_p & v844f9f;
assign v890c16 = BtoS_ACK3_p & v8b280c | !BtoS_ACK3_p & v8afea6;
assign v8c3b67 = RtoB_ACK0_p & v8b77fb | !RtoB_ACK0_p & v912777;
assign v8b22f0 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v88e0ec;
assign v911fbe = BtoS_ACK0_p & v8ae151 | !BtoS_ACK0_p & v892858;
assign v8b1f58 = EMPTY_p & v912423 | !EMPTY_p & v87de99;
assign v8b1ffd = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91244f;
assign v8f960f = BtoS_ACK7_p & v8af4ee | !BtoS_ACK7_p & v912706;
assign v8aff37 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b013b;
assign v910c69 = jx0_p & v91274f | !jx0_p & v912698;
assign v8ae86c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v910bd3;
assign v8b2cb0 = StoB_REQ6_p & v9111d2 | !StoB_REQ6_p & v8c5e54;
assign v890a9a = StoB_REQ3_p & v8afdde | !StoB_REQ3_p & v844f91;
assign v8c3f33 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8c6c00;
assign v911218 = BtoS_ACK7_p & v8ae4e9 | !BtoS_ACK7_p & v8b11c5;
assign v911395 = stateG7_1_p & v911765 | !stateG7_1_p & v8c4740;
assign v88d6cf = BtoS_ACK0_p & v881ef0 | !BtoS_ACK0_p & v864227;
assign v912046 = RtoB_ACK0_p & v8f9630 | !RtoB_ACK0_p & v8afe84;
assign v8f9630 = jx2_p & v8aed37 | !jx2_p & v8aed2e;
assign v8bfab7 = BtoS_ACK3_p & v88709f | !BtoS_ACK3_p & v8c3f33;
assign v8ae03c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8c0b9e;
assign v8af0b0 = BtoS_ACK0_p & v8ae151 | !BtoS_ACK0_p & v8af894;
assign v8dd6ad = jx0_p & v91180c | !jx0_p & v844f91;
assign v91187a = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v8b004e;
assign v8b320b = jx0_p & v844f91 | !jx0_p & v8b76f1;
assign v8c51d8 = jx0_p & v8c4410 | !jx0_p & v8b76f1;
assign v8b004c = BtoS_ACK7_p & v911149 | !BtoS_ACK7_p & v8b1d42;
assign v912026 = BtoS_ACK1_p & v8b07c0 | !BtoS_ACK1_p & v8b3d0e;
assign v8aef55 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91268d;
assign v8924ff = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8ae731;
assign v912502 = jx0_p & v8afb17 | !jx0_p & v844f91;
assign v87cd98 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v9125dd;
assign v88fa8c = jx2_p & v8aff75 | !jx2_p & v8b2021;
assign v8db1d7 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8b08e5;
assign v912444 = jx2_p & v9113cc | !jx2_p & !v8af2cd;
assign v8b0c98 = jx1_p & v8af318 | !jx1_p & !v844f91;
assign v8c04cb = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8674d8;
assign v8b76ff = BtoR_REQ1_p & v8c0b95 | !BtoR_REQ1_p & v9125fc;
assign v8b12e9 = stateG7_1_p & v8ae8e3 | !stateG7_1_p & v911fdf;
assign v911914 = BtoS_ACK7_p & v9124fd | !BtoS_ACK7_p & v867e4e;
assign v91272c = stateG7_1_p & v88c831 | !stateG7_1_p & v8c66bb;
assign v8b0e4c = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & !v844f91;
assign v9115fc = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v9123f8;
assign v8b52fa = jx1_p & v8af02f | !jx1_p & !v8b2aa2;
assign v8b08ff = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b11b0;
assign v911bad = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c0b8f;
assign v8b2c52 = jx3_p & v8c5357 | !jx3_p & v8b2c4e;
assign v8b3401 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b21e7;
assign v8db195 = stateG7_1_p & v88340e | !stateG7_1_p & v844f91;
assign v8b0e67 = jx3_p & v844f91 | !jx3_p & !v912692;
assign v8c41ae = BtoS_ACK6_p & v911bad | !BtoS_ACK6_p & v912730;
assign v8c3d99 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b0eab;
assign v91247c = jx1_p & v8b07a1 | !jx1_p & !v8c50c4;
assign v91274f = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v89407e;
assign v8afec3 = jx1_p & v8771a0 | !jx1_p & v8b0b2b;
assign v8b2920 = jx0_p & v8af564 | !jx0_p & v91185f;
assign v8b1110 = RtoB_ACK1_p & v8cf811 | !RtoB_ACK1_p & v8c6979;
assign v8c3925 = BtoR_REQ1_p & v8aeabf | !BtoR_REQ1_p & v911441;
assign v890c07 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v9125f0;
assign v8c043d = BtoR_REQ1_p & v912472 | !BtoR_REQ1_p & v8cc197;
assign v8dd5cf = BtoS_ACK0_p & v9123df | !BtoS_ACK0_p & v8b0151;
assign v91257b = jx2_p & v8b2f46 | !jx2_p & v8aed2e;
assign v8aebed = StoB_REQ0_p & v8b12f9 | !StoB_REQ0_p & v8af77e;
assign v8b034f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9b;
assign v85d9b6 = jx0_p & v8b6d7e | !jx0_p & v9115ca;
assign v8b02ce = stateG7_1_p & v8c0a62 | !stateG7_1_p & v844f91;
assign v8b4fda = BtoS_ACK0_p & v8f9617 | !BtoS_ACK0_p & v91261f;
assign v8c0b9e = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c4a57;
assign v8ae0ee = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8c43e6;
assign v8b09b0 = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v912589;
assign v8b76f3 = BtoR_REQ1_p & v8b0c90 | !BtoR_REQ1_p & v8b2a8c;
assign v8ae0da = jx2_p & v8b1166 | !jx2_p & !v8dd691;
assign v912516 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v887b94;
assign v884789 = StoB_REQ2_p & v8c4b39 | !StoB_REQ2_p & v9126a8;
assign v911fe2 = stateG7_1_p & v8b218f | !stateG7_1_p & v8aee08;
assign v912558 = StoB_REQ6_p & v8e983b | !StoB_REQ6_p & v8c5bc3;
assign v91276d = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v9121e7;
assign v8b0b7a = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v9126b1;
assign v8af624 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c5e9b;
assign v88547b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8db180;
assign v8c0b07 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8c04cb;
assign v8b0903 = DEQ_p & v912522 | !DEQ_p & v8b9047;
assign v8ae5c0 = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v892555;
assign v8b290b = BtoS_ACK4_p & v8b0c7c | !BtoS_ACK4_p & v8afea6;
assign v89409b = jx1_p & v8b085b | !jx1_p & !v8b2d81;
assign v91134e = RtoB_ACK1_p & v912413 | !RtoB_ACK1_p & v912747;
assign v8b25ff = jx0_p & v8aedac | !jx0_p & v9126b0;
assign v87cfd0 = jx0_p & v8af415 | !jx0_p & v8b0b29;
assign v8fec8f = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8c23c8;
assign v8602f3 = jx0_p & v8c52db | !jx0_p & v88ee77;
assign v8f96fd = BtoS_ACK1_p & v8c0b8f | !BtoS_ACK1_p & v912390;
assign v91273e = BtoS_ACK6_p & v912702 | !BtoS_ACK6_p & v892f3e;
assign v91216a = StoB_REQ0_p & v8b33fa | !StoB_REQ0_p & v912075;
assign v8b0c14 = BtoR_REQ0_p & v911395 | !BtoR_REQ0_p & v8bfa6b;
assign v85a47c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8c6ccc;
assign v890b41 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v912631;
assign v8af2e3 = BtoR_REQ0_p & v9124e7 | !BtoR_REQ0_p & v8c3925;
assign v8b08e5 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8c0ab9;
assign v8b0ae9 = BtoR_REQ1_p & v912785 | !BtoR_REQ1_p & v9125fc;
assign v8b1367 = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v91271e;
assign v9125c5 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & !v9126c2;
assign v8b1c79 = StoB_REQ3_p & v8b290b | !StoB_REQ3_p & !v844f9f;
assign v8aee49 = StoB_REQ1_p & v8c4b39 | !StoB_REQ1_p & v8579b7;
assign v87ba6d = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8b02ed;
assign v9123d2 = jx1_p & v8ae6f2 | !jx1_p & !v8bfa65;
assign v8b24cc = jx3_p & v912711 | !jx3_p & v912698;
assign v890b15 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b2876;
assign v8714a5 = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & v8ae516;
assign v8b280c = StoB_REQ3_p & v8afea6 | !StoB_REQ3_p & !v844f9f;
assign v8dd643 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8b2f95;
assign v8b0eb6 = jx2_p & v8afa8e | !jx2_p & v9125d9;
assign v870c3a = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8bfab7;
assign v8b2ab3 = jx1_p & v91271d | !jx1_p & v912765;
assign v8b2fc3 = BtoS_ACK0_p & v879d5b | !BtoS_ACK0_p & v8742de;
assign v8af698 = StoB_REQ6_p & v8f9587 | !StoB_REQ6_p & v8b2e27;
assign v910e98 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & v88e0ec;
assign v911441 = stateG7_1_p & v8b2df5 | !stateG7_1_p & v911cec;
assign v8f9724 = DEQ_p & v8cc1e2 | !DEQ_p & v8c0433;
assign v912450 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f9b;
assign v8b048e = StoB_REQ3_p & v9124ed | !StoB_REQ3_p & v8b1f47;
assign v8ae714 = StoB_REQ7_p & v8b0753 | !StoB_REQ7_p & v8b2b2d;
assign v8b0429 = EMPTY_p & v912680 | !EMPTY_p & v8c39e1;
assign v893433 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v911c5d;
assign v912523 = StoB_REQ2_p & v91274b | !StoB_REQ2_p & v8b1406;
assign v912537 = ENQ_p & v912747 | !ENQ_p & !v91151a;
assign v8b016b = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v8a8ba3;
assign v87bbef = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & !v8b1e6a;
assign v911a0d = jx0_p & v8f960f | !jx0_p & v8b2ae9;
assign v9118c2 = stateG12_p & v8b7bb3 | !stateG12_p & v8c500e;
assign v844fa3 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844f91;
assign v911fa4 = jx3_p & v844f91 | !jx3_p & !v844fbb;
assign v8b10cf = StoB_REQ6_p & v8b03cf | !StoB_REQ6_p & v844f91;
assign v8b2998 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v9125ad;
assign v86990d = jx1_p & v8b2b91 | !jx1_p & !v8b29d6;
assign v8c0b7c = BtoS_ACK7_p & v844f9d | !BtoS_ACK7_p & v8b77fc;
assign v8c3050 = stateG7_1_p & v844f91 | !stateG7_1_p & v8b21ba;
assign v9124fd = StoB_REQ6_p & v912518 | !StoB_REQ6_p & v844f91;
assign v8b0cbf = stateG7_1_p & v911e5a | !stateG7_1_p & v844f91;
assign v8b1e11 = StoB_REQ2_p & v8af683 | !StoB_REQ2_p & v911fd6;
assign v8b1276 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8b13b1;
assign v8b1e7b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c568f;
assign v910947 = jx2_p & v8af89d | !jx2_p & v87ebfd;
assign v85c0bd = BtoR_REQ1_p & v8af74b | !BtoR_REQ1_p & v8c6979;
assign v8c41aa = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v91207b;
assign v912492 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v910ff3;
assign v8ae562 = BtoS_ACK7_p & v9124fd | !BtoS_ACK7_p & v912186;
assign v8b0a5f = stateG7_1_p & v8af1a2 | !stateG7_1_p & v8f9597;
assign v8afb17 = BtoS_ACK7_p & v844f97 | !BtoS_ACK7_p & v8b2511;
assign v8aefce = StoB_REQ0_p & v911664 | !StoB_REQ0_p & v8aec85;
assign v88fa49 = BtoS_ACK3_p & v912763 | !BtoS_ACK3_p & v8b048e;
assign v9126b4 = jx1_p & v8771a0 | !jx1_p & v91242f;
assign v8aed0c = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8d540a;
assign v8b2049 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b0151;
assign v8b03fe = BtoS_ACK0_p & v8d6d04 | !BtoS_ACK0_p & v9124f8;
assign v911d4f = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v844f91;
assign v8b1ddc = BtoS_ACK6_p & v8b10fd | !BtoS_ACK6_p & v8b2bbf;
assign v912696 = StoB_REQ3_p & v8c381a | !StoB_REQ3_p & v8b2a3e;
assign v9125ec = stateG7_1_p & v91261a | !stateG7_1_p & v8b2a14;
assign v8b2c35 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8af634;
assign v912588 = StoB_REQ1_p & v9125b1 | !StoB_REQ1_p & v8af7b5;
assign v8c4a56 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b25a4;
assign v8b2173 = BtoS_ACK6_p & v912432 | !BtoS_ACK6_p & v8af949;
assign v8af717 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8aec59;
assign v8ae77f = BtoS_ACK6_p & v91265d | !BtoS_ACK6_p & v8b11f0;
assign v8c04c4 = jx1_p & v8909d0 | !jx1_p & !v8c3e35;
assign v85c141 = BtoS_ACK7_p & v844f99 | !BtoS_ACK7_p & v8b09b0;
assign v91256c = StoB_REQ3_p & v912627 | !StoB_REQ3_p & !v844f9f;
assign v9123e7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v871da5;
assign v8b00a9 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v88bebc;
assign v844fb7 = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & !v844f91;
assign v8b038e = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v8af205;
assign v8e990e = StoB_REQ2_p & v8bfab7 | !StoB_REQ2_p & v844f91;
assign v894072 = BtoS_ACK7_p & v91257d | !BtoS_ACK7_p & v8b1ff0;
assign v8af015 = jx2_p & v8b2a8c | !jx2_p & v8b0cf7;
assign v8b0b9e = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8b263d;
assign v8b1cd0 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v8c557c;
assign v8b25a4 = StoB_REQ2_p & v8b339d | !StoB_REQ2_p & v9116aa;
assign v91141d = jx1_p & v88b60c | !jx1_p & !v8dd667;
assign BtoS_ACK1_n = !v8f9724;
assign v8c5357 = BtoS_ACK7_p & v88b300 | !BtoS_ACK7_p & v8afd2b;
assign v912507 = jx0_p & v8b2878 | !jx0_p & !v89098b;
assign v91257c = jx1_p & v8b07a1 | !jx1_p & !v8c6e12;
assign v8aec34 = StoB_REQ1_p & v9124c9 | !StoB_REQ1_p & v844f91;
assign v866ac1 = BtoS_ACK0_p & v8fed10 | !BtoS_ACK0_p & v911291;
assign v8b0554 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ae805;
assign v8ae7c9 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v9126cb;
assign v911917 = StoB_REQ2_p & v8aec57 | !StoB_REQ2_p & v85ed5d;
assign v8b8e74 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & !v911c88;
assign v8aedf0 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8dd643;
assign v8bb768 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8b1d12;
assign v8c7159 = jx2_p & v8bfa26 | !jx2_p & v8afe97;
assign v8b00f2 = StoB_REQ3_p & v8b0d0e | !StoB_REQ3_p & !v844f9f;
assign v8b1150 = BtoS_ACK0_p & v8b0a55 | !BtoS_ACK0_p & v912714;
assign v8b22d1 = BtoS_ACK3_p & v8b20b7 | !BtoS_ACK3_p & v8c43e6;
assign v8af1d7 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v87cf74;
assign v85c135 = StoB_REQ2_p & v8bfab7 | !StoB_REQ2_p & v870c3a;
assign v8b120b = StoB_REQ2_p & v8b2d4a | !StoB_REQ2_p & !v8af382;
assign v9124df = EMPTY_p & v9123d7 | !EMPTY_p & v8b0942;
assign v8b267a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b00a7;
assign v911b49 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v91251b;
assign v8c48a8 = jx1_p & v844f91 | !jx1_p & v8af586;
assign v9124ef = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b209b;
assign v8b13f6 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v912681;
assign v91240d = jx0_p & v8b2592 | !jx0_p & v8aed6d;
assign v8b2c4c = jx3_p & v844f91 | !jx3_p & !v8af9f6;
assign v8b2252 = StoB_REQ4_p & v8afea6 | !StoB_REQ4_p & v844f91;
assign v8b2a8c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v911c7e;
assign v8af918 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v912605;
assign v89092e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b28e6;
assign v8b23c7 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8af9e8;
assign v8af9f6 = jx0_p & v8c53ab | !jx0_p & !v8b1e7d;
assign v8af756 = ENQ_p & v8c70fc | !ENQ_p & v911d22;
assign v9126c3 = jx2_p & v887bcc | !jx2_p & v8cc1c4;
assign v8b12b1 = RtoB_ACK1_p & v91270f | !RtoB_ACK1_p & v912698;
assign v8c57f0 = BtoR_REQ1_p & v8f96e9 | !BtoR_REQ1_p & v912678;
assign v912414 = BtoS_ACK1_p & v879d5b | !BtoS_ACK1_p & v8b1d1f;
assign v8afe2c = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b208f;
assign v8f9597 = RtoB_ACK0_p & v8c723e | !RtoB_ACK0_p & v8af1a2;
assign v85c0eb = jx1_p & v8b114d | !jx1_p & v8c5357;
assign v912512 = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8c3651;
assign v9126da = StoB_REQ6_p & v8ae446 | !StoB_REQ6_p & v8b11f0;
assign v9112d7 = RtoB_ACK1_p & v8cc0f3 | !RtoB_ACK1_p & v8af015;
assign v8af78a = jx0_p & v8b216f | !jx0_p & v910c1b;
assign v8b0e8e = stateG7_1_p & v844f91 | !stateG7_1_p & v8c0435;
assign v911f4a = EMPTY_p & v8b0c14 | !EMPTY_p & v911913;
assign v8b2642 = FULL_p & v9111f5 | !FULL_p & v8c3d52;
assign v911f9b = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8ae556;
assign v911fd2 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8c6cee;
assign v911173 = RtoB_ACK0_p & v8ae5e2 | !RtoB_ACK0_p & v9115b8;
assign v8af066 = BtoR_REQ0_p & v912430 | !BtoR_REQ0_p & v8aef67;
assign v8b066c = jx1_p & v912074 | !jx1_p & !v8b266b;
assign v91155b = jx1_p & v8af03b | !jx1_p & v8b244a;
assign v8c0aba = EMPTY_p & v91100d | !EMPTY_p & v9111c2;
assign v8aeb57 = jx0_p & v8b1f0a | !jx0_p & !v844f91;
assign v8ae5c6 = jx1_p & v8aeada | !jx1_p & v8b0ef5;
assign v8ae803 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v89286e;
assign v9124ad = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8afe2c;
assign v911e5a = RtoB_ACK1_p & v9123b1 | !RtoB_ACK1_p & v844f91;
assign v911633 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0b6b;
assign v88331f = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v912733;
assign v91255a = BtoS_ACK0_p & v9123df | !BtoS_ACK0_p & v8ae878;
assign v912522 = ENQ_p & v9115b8 | !ENQ_p & v8b070e;
assign v8b0a04 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8b06d3;
assign v8c42f9 = jx1_p & v8b2180 | !jx1_p & v8ae765;
assign v912729 = stateG7_1_p & v9126db | !stateG7_1_p & !v911f9c;
assign v8b0be4 = StoB_REQ0_p & v912549 | !StoB_REQ0_p & v8ae64c;
assign v8f96e8 = StoB_REQ2_p & v8b1ea2 | !StoB_REQ2_p & v844f91;
assign v8e9903 = BtoS_ACK1_p & v8af634 | !BtoS_ACK1_p & v9123df;
assign v8b7801 = jx1_p & v91265c | !jx1_p & v8b0446;
assign v8af65e = BtoR_REQ0_p & v887acc | !BtoR_REQ0_p & !v856df0;
assign v8b4fb2 = RtoB_ACK0_p & v8c3cff | !RtoB_ACK0_p & v912122;
assign v912642 = stateG12_p & v911a5e | !stateG12_p & v8b09fb;
assign v91244f = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v8af73a;
assign v8689df = BtoS_ACK6_p & v844f9d | !BtoS_ACK6_p & v8b23de;
assign v8af0c8 = jx2_p & v8c70fd | !jx2_p & v9124b5;
assign v887b1c = jx3_p & v844f91 | !jx3_p & v8b3350;
assign v8b3d1f = BtoS_ACK7_p & v91257d | !BtoS_ACK7_p & v8b2197;
assign v9107fb = stateG7_1_p & v8af478 | !stateG7_1_p & v844f91;
assign v8c43ba = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8fed23;
assign v8b1159 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b038e;
assign v9125e3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8af215;
assign v9124c8 = BtoS_ACK6_p & v844f9f | !BtoS_ACK6_p & v8b2df8;
assign v8c3d7b = stateG7_1_p & v8cc108 | !stateG7_1_p & v8af02f;
assign v912634 = StoB_REQ6_p & v88d6cf | !StoB_REQ6_p & v866ac1;
assign v8b073b = StoB_REQ7_p & v91250e | !StoB_REQ7_p & v844f91;
assign v912312 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8aeed6;
assign v912198 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8b2bc5;
assign v8b2a2e = stateG7_1_p & v8af8f5 | !stateG7_1_p & v912698;
assign v8924d2 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v8b2a3e;
assign jx0_n = !v8e9961;
assign v8ae9f4 = jx2_p & v8908a2 | !jx2_p & !v8ae46b;
assign v8909d0 = jx0_p & v8b1276 | !jx0_p & !v86f3ae;
assign v9123b9 = jx2_p & v8c34da | !jx2_p & v9124c2;
assign v911fd9 = BtoS_ACK7_p & v844f9b | !BtoS_ACK7_p & v8c23d8;
assign v9123cc = BtoS_ACK6_p & v844f99 | !BtoS_ACK6_p & v8b1ec4;
assign v8cc1e2 = ENQ_p & v912698 | !ENQ_p & v8c72da;
assign v8af5f1 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8e983b;
assign v912487 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v87d059 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v912450;
assign v8af366 = stateG7_1_p & v8b134f | !stateG7_1_p & v8b02e9;
assign v8ae104 = stateG7_1_p & v911174 | !stateG7_1_p & v910db7;
assign v8b3c24 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8ae925;
assign v91264e = jx0_p & v8b4fca | !jx0_p & !v8bfa76;
assign v8afd20 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v912575;
assign v912480 = RtoB_ACK1_p & v8b28d4 | !RtoB_ACK1_p & v8afe84;
assign v8b5a58 = BtoS_ACK6_p & v912609 | !BtoS_ACK6_p & v9115c6;
assign v8b23bf = jx0_p & v8c3a0b | !jx0_p & v910c1b;
assign v8c34ba = jx1_p & v88fef2 | !jx1_p & v8b1e70;
assign v8aff15 = StoB_REQ0_p & v8fec8f | !StoB_REQ0_p & v844f91;
assign v8b2e72 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b0f42;
assign v9126ae = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & !v8b120b;
assign v8c4ac3 = StoB_REQ3_p & v912517 | !StoB_REQ3_p & v8b1f47;
assign v8db1b0 = BtoS_ACK2_p & v88709f | !BtoS_ACK2_p & v8af683;
assign v8b01e2 = BtoS_ACK6_p & v8bfa8b | !BtoS_ACK6_p & v8af155;
assign v8b236f = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v91269f;
assign v9124e0 = BtoS_ACK6_p & v8c6c4a | !BtoS_ACK6_p & v912514;
assign v912717 = stateG7_1_p & v910c73 | !stateG7_1_p & v844f91;
assign v8ae4a3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v890c1b;
assign v9114f1 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8c48a1;
assign v8af34a = stateG7_1_p & v890ac0 | !stateG7_1_p & v912529;
assign v8b0693 = RtoB_ACK1_p & v912122 | !RtoB_ACK1_p & v844f91;
assign v8c458b = StoB_REQ0_p & v8b28e6 | !StoB_REQ0_p & v8af214;
assign v8b0d0e = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v912517;
assign v8b0eea = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8b0d2f;
assign v9124b0 = StoB_REQ2_p & v9123b3 | !StoB_REQ2_p & v8af3eb;
assign v879d5b = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v844f91;
assign v8b1ca6 = BtoR_REQ0_p & v8af83a | !BtoR_REQ0_p & v8aedc6;
assign v9123df = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b229e;
assign v8af753 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & !v844fb9;
assign v911d50 = BtoR_REQ0_p & v912746 | !BtoR_REQ0_p & v9123e9;
assign v912657 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & v912756;
assign v8b2c6b = BtoS_ACK1_p & v8b1e22 | !BtoS_ACK1_p & v8b0df4;
assign v912732 = StoB_REQ6_p & v844f91 | !StoB_REQ6_p & v91268b;
assign v911e75 = BtoS_ACK7_p & v912609 | !BtoS_ACK7_p & v8b2445;
assign v8ae909 = jx2_p & v8afec3 | !jx2_p & v91141d;
assign v911ef8 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v911f1c;
assign v8afa37 = jx3_p & v844f91 | !jx3_p & v8c6c93;
assign v912283 = BtoS_ACK4_p & v8dd687 | !BtoS_ACK4_p & v844f9d;
assign v8c6cdc = StoB_REQ7_p & v8b0500 | !StoB_REQ7_p & v890534;
assign v8aef35 = jx2_p & v8af39f | !jx2_p & v8c56dd;
assign v9116e8 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8c6c7e;
assign v8908a2 = jx1_p & v8aea38 | !jx1_p & !v8b05e2;
assign v8aec42 = jx0_p & v8b2bd8 | !jx0_p & !v844f9d;
assign v8b2c26 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b2935;
assign v870559 = BtoS_ACK2_p & v8b33a8 | !BtoS_ACK2_p & v88f72f;
assign v8b261e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b28a7;
assign v8afde2 = jx2_p & v8e9954 | !jx2_p & v890ac0;
assign v910d87 = ENQ_p & v887c3b | !ENQ_p & !v8b0429;
assign v912632 = jx1_p & v91174f | !jx1_p & v912656;
assign v8b0599 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v912683;
assign v911978 = StoB_REQ1_p & v8b0283 | !StoB_REQ1_p & v8596e1;
assign v8b222c = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8afd2b;
assign v911a56 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8b0fe0;
assign v8b2f8c = StoB_REQ6_p & v8fed43 | !StoB_REQ6_p & !v844f91;
assign v911539 = BtoS_ACK0_p & v91244d | !BtoS_ACK0_p & v8c57ef;
assign v8b4c61 = BtoS_ACK0_p & v8afe4c | !BtoS_ACK0_p & v8b76f4;
assign v8b131b = BtoS_ACK0_p & v8dd65f | !BtoS_ACK0_p & v8aebed;
assign v8b7669 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b4d42;
assign v912737 = RtoB_ACK0_p & v8b07f3 | !RtoB_ACK0_p & v8b0a89;
assign v91267e = jx0_p & v91118f | !jx0_p & v912408;
assign v8c0b04 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v8dd5e2;
assign v8c4072 = StoB_REQ6_p & v912636 | !StoB_REQ6_p & v8af193;
assign v9114a2 = BtoS_ACK6_p & v844f97 | !BtoS_ACK6_p & v8c7054;
assign v8b12eb = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8b6e0a;
assign v8ae51a = jx0_p & v8f96c9 | !jx0_p & !v8e994b;
assign v8b241a = jx0_p & v8b4fca | !jx0_p & !v844f9d;
assign v912626 = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v9119a4;
assign v91230d = BtoR_REQ0_p & v8af83a | !BtoR_REQ0_p & v91264b;
assign v8b01f5 = stateG7_1_p & v8b28d4 | !stateG7_1_p & v8b03ed;
assign v8b0a19 = jx2_p & v8618ae | !jx2_p & !v8b3416;
assign v88f796 = jx0_p & v86995b | !jx0_p & v911633;
assign v8b2a34 = jx0_p & v8b0298 | !jx0_p & v844f91;
assign v8af8b0 = jx1_p & v8c460a | !jx1_p & v8af6e2;
assign v8af6e2 = jx3_p & v844f91 | !jx3_p & v89217c;
assign v8b2fea = BtoS_ACK6_p & v912702 | !BtoS_ACK6_p & v8dd637;
assign v911e6a = BtoS_ACK6_p & v912432 | !BtoS_ACK6_p & v89223a;
assign v8af640 = BtoR_REQ0_p & v8b0cbf | !BtoR_REQ0_p & v91243a;
assign v8c46bf = jx0_p & v8b1f0a | !jx0_p & !v8aed6d;
assign v9123cd = jx1_p & v844f91 | !jx1_p & !v8b2c29;
assign v912699 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8aee3c;
assign v8b12d5 = StoB_REQ7_p & v8c6aa0 | !StoB_REQ7_p & v8afe06;
assign v8af9be = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b22ef;
assign v912400 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8692ec;
assign v8c4c96 = jx0_p & v8b2878 | !jx0_p & !v8af9f2;
assign v8b2b4a = BtoS_ACK6_p & v91222a | !BtoS_ACK6_p & v8c6c8b;
assign v8b4d42 = BtoS_ACK6_p & v8b2019 | !BtoS_ACK6_p & v8af05a;
assign v8b0dc1 = StoB_REQ7_p & v8aed74 | !StoB_REQ7_p & v8c0b46;
assign v8db217 = StoB_REQ1_p & v8b034f | !StoB_REQ1_p & v844f91;
assign v912786 = StoB_REQ2_p & v8c4c30 | !StoB_REQ2_p & !v911484;
assign v8aef4e = jx1_p & v91271d | !jx1_p & v8c45e8;
assign v892858 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fed5e;
assign v91240a = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v9121ee;
assign v8b0df4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8b1e22;
assign v8c56dd = jx1_p & v8ba4a1 | !jx1_p & v8b0e67;
assign v8b20ab = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8fed12;
assign v8b0762 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v8afea6;
assign v9126eb = jx0_p & v844f91 | !jx0_p & v87ebfd;
assign v912793 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8fedd4;
assign v8b27ec = StoB_REQ1_p & v87b5cf | !StoB_REQ1_p & v8b0219;
assign v887bcd = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8c71b3;
assign v8afa3c = jx1_p & v8aea38 | !jx1_p & !v890992;
assign v8b0c7c = StoB_REQ4_p & v8afea6 | !StoB_REQ4_p & !v844f9f;
assign v911c5d = StoB_REQ0_p & v8b0934 | !StoB_REQ0_p & v911f9b;
assign v9124b4 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v87bbef;
assign v91269a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b7892;
assign v9125af = stateG7_1_p & v8b2a8d | !stateG7_1_p & v8b10bf;
assign v912471 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91275d;
assign v8b129a = StoB_REQ3_p & v8b339d | !StoB_REQ3_p & v844f91;
assign v8b11f0 = BtoS_ACK0_p & v8b7794 | !BtoS_ACK0_p & v91265d;
assign v912678 = stateG7_1_p & v911704 | !stateG7_1_p & v8b116b;
assign v8b06bb = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v91129a;
assign v882969 = stateG7_1_p & v912122 | !stateG7_1_p & v8b4fb2;
assign v8aea10 = StoB_REQ1_p & v9126f4 | !StoB_REQ1_p & v8ae147;
assign v8924fb = jx0_p & v9123eb | !jx0_p & v844f99;
assign v912695 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v911fae;
assign v912236 = jx0_p & v91271f | !jx0_p & v9115ca;
assign v912075 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8b1fe8;
assign v8b0d78 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8aefa4;
assign v8fed5b = BtoS_ACK6_p & v8af431 | !BtoS_ACK6_p & v8b1e33;
assign v8ae12e = jx0_p & v8c4a25 | !jx0_p & v8ae048;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v8af62a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8b3212;
assign v9124cf = RtoB_ACK0_p & v8b13ca | !RtoB_ACK0_p & v88acc3;
assign v8b266b = jx0_p & v8b1ec1 | !jx0_p & v888766;
assign v87ab76 = BtoR_REQ1_p & v9125ec | !BtoR_REQ1_p & v844f91;
assign v9126bc = BtoS_ACK2_p & v8ae516 | !BtoS_ACK2_p & v91266e;
assign v8b11df = BtoS_ACK6_p & v8ae878 | !BtoS_ACK6_p & v8aec17;
assign v8e98af = BtoS_ACK7_p & v8af431 | !BtoS_ACK7_p & v845125;
assign v8b07b6 = BtoS_ACK7_p & v844f91 | !BtoS_ACK7_p & v91254a;
assign v91242c = jx1_p & v8c51d8 | !jx1_p & v8af78a;
assign v8b2b80 = jx0_p & v8b3d09 | !jx0_p & v8b76f1;
assign v887b47 = BtoR_REQ0_p & v8b25a8 | !BtoR_REQ0_p & v9125da;
assign v8784da = jx1_p & v8b2a71 | !jx1_p & v8ae074;
assign v8c45be = BtoS_ACK7_p & v844f9f | !BtoS_ACK7_p & v91276d;
assign v872c7c = StoB_REQ6_p & v9121e7 | !StoB_REQ6_p & v912638;
assign v91265a = BtoS_ACK3_p & v8ae4cd | !BtoS_ACK3_p & v8b3321;
assign v91251a = StoB_REQ3_p & v8b339d | !StoB_REQ3_p & !v844f91;
assign v8b210b = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8b1ea2;
assign v8b229e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8af634;
assign v8b09e5 = BtoS_ACK2_p & v8924d2 | !BtoS_ACK2_p & v8c4ac3;
assign v8af193 = BtoS_ACK0_p & v8c6cee | !BtoS_ACK0_p & v8c390a;
assign v912724 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8af916;
assign v88f72f = BtoS_ACK3_p & v8b33a8 | !BtoS_ACK3_p & v8c6bef;
assign v910bd1 = jx1_p & v911772 | !jx1_p & !v8c353f;
assign v8af582 = StoB_REQ1_p & v8b139e | !StoB_REQ1_p & v8af7df;
assign v8f965b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c458b;
assign v8b1178 = stateG7_1_p & v8c387f | !stateG7_1_p & v8ae14c;
assign v9123d7 = BtoR_REQ0_p & v8b01d5 | !BtoR_REQ0_p & v9116e0;
assign v912584 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v91093d;
assign v8b1f71 = BtoS_ACK6_p & v844f91 | !BtoS_ACK6_p & v8b2d92;
assign v8ae7a9 = BtoS_ACK7_p & v8b0cbb | !BtoS_ACK7_p & v91250a;
assign v8b0a2d = StoB_REQ0_p & v91277b | !StoB_REQ0_p & v8b2f6d;
assign v890a64 = BtoS_ACK7_p & v8af431 | !BtoS_ACK7_p & v8fedea;
assign v8c7385 = StoB_REQ7_p & v844f91 | !StoB_REQ7_p & v8b05b0;
assign v869f57 = StoB_REQ7_p & v91104c | !StoB_REQ7_p & v844f91;
assign v911d0d = jx0_p & v8aed6d | !jx0_p & v911b46;
assign v8ae4ce = jx2_p & v8c44cf | !jx2_p & v844f91;
assign v8b2275 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v87d059;
assign ENQ_n = (DEQ_n & ((FULL_n & ((stateG12_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))) | (!FULL_n & ((stateG12_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!DEQ_n & ((EMPTY_n & ((stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n) | (!StoB_REQ1_n & ((!jx2_n & ((jx1_n & ((!jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((RtoB_ACK1_n & ((BtoR_REQ0_n) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n))))) | (!RtoB_ACK1_n & ((BtoR_REQ0_n) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n))))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((jx2_n) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n))))))) | (!EMPTY_n & ((!FULL_n & ((stateG12_n & ((stateG7_0_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))) | (!stateG12_n & ((stateG7_0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))))))) | (!StoB_REQ6_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))) | (!StoB_REQ3_n & ((!BtoS_ACK3_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))))))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n) | (!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n))))))) | (!StoB_REQ4_n & ((!BtoS_ACK4_n & ((BtoS_ACK5_n & ((StoB_REQ5_n)))))))))))))))))))))))))))))))))))))))))))))))));
assign SLC0_n = (DEQ_n & ((FULL_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((BtoS_ACK6_n & ((ENQ_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))) | (!BtoS_ACK2_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx3_n))))))))))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))) | (!FULL_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((BtoS_ACK6_n & ((ENQ_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))) | (!BtoS_ACK2_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx3_n))))))))))))))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))) | (!DEQ_n & ((EMPTY_n & ((stateG7_0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((stateG7_0_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((BtoS_ACK6_n & ((ENQ_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))) | (!BtoS_ACK2_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx3_n))))))))))))))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))) | (!stateG12_n & ((stateG7_0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n))))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK4_n))) | (!StoB_REQ3_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((jx3_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx3_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((StoB_REQ3_n & ((!StoB_REQ4_n))) | (!StoB_REQ3_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))))) | (!StoB_REQ7_n & ((!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))) | (!jx0_n & ((SLC1_n))))) | (!jx1_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!jx2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!StoB_REQ0_n & ((ENQ_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx0_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n))))))))))) | (!BtoS_ACK2_n & ((SLC1_n) | (!SLC1_n & ((!BtoS_ACK4_n)))))))))))))))))))))))))))))))))))));
assign SLC2_n = (DEQ_n & ((FULL_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))) | (!BtoS_ACK1_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n) | (!jx1_n & ((!SLC1_n))))) | (!jx3_n))))))))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))))) | (!stateG7_1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))) | (!FULL_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))) | (!BtoS_ACK1_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n) | (!jx1_n & ((!SLC1_n))))) | (!jx3_n))))))))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))))) | (!stateG7_1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))))) | (!DEQ_n & ((EMPTY_n & ((stateG7_0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n))) | (!BtoS_ACK2_n))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n))) | (!BtoS_ACK2_n))))))))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n))))))))))))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((stateG7_0_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n & ((BtoS_ACK1_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))) | (!BtoS_ACK1_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n) | (!jx1_n & ((!SLC1_n))))) | (!jx3_n))))))))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n))) | (!BtoS_ACK2_n))))))))))))))))))) | (!BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n))) | (!BtoS_ACK2_n))))))))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))))))))))) | (!stateG12_n & ((stateG7_0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n))) | (!BtoS_ACK2_n))))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n))) | (!BtoS_ACK2_n))))))))))))))))))) | (!BtoR_REQ1_n & ((SLC0_n & ((BtoS_ACK7_n & ((ENQ_n))) | (!BtoS_ACK7_n & ((StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((jx0_n & ((!SLC1_n))))) | (!jx1_n & ((!SLC1_n))))) | (!jx2_n & ((!SLC1_n))))))))) | (!StoB_REQ6_n & ((ENQ_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))))))) | (!SLC0_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((ENQ_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK0_n & ((ENQ_n & ((BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK2_n))))))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((!jx2_n & ((!jx3_n & ((!jx1_n & ((!jx0_n))))))))))) | (!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((ENQ_n))) | (!BtoS_ACK6_n & ((StoB_REQ6_n & ((!BtoS_ACK0_n & ((ENQ_n & ((!BtoS_ACK2_n))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((ENQ_n & ((!BtoS_ACK2_n))))) | (!StoB_REQ0_n & ((ENQ_n & ((StoB_REQ1_n & ((!BtoS_ACK2_n))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((jx2_n & ((!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n)))))))))))))))))))))))))))))));
assign SLC1_n = (DEQ_n & ((stateG12_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))) | (!stateG7_1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))) | (!DEQ_n & ((EMPTY_n & ((stateG7_0_n & ((stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!StoB_REQ6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((!jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))))) | (!stateG7_0_n & ((stateG7_1_n & ((RtoB_ACK1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))) | (!RtoB_ACK1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n) | (!StoB_REQ6_n & ((jx2_n & ((jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((jx2_n) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!StoB_REQ2_n & ((jx2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx2_n & ((jx3_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx3_n & ((jx1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx2_n & ((jx3_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx3_n & ((jx1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((jx2_n) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n & ((jx2_n) | (!jx2_n & ((jx3_n) | (!jx3_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))))) | (!StoB_REQ2_n & ((jx2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx2_n & ((jx3_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx3_n & ((jx1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))) | (!BtoS_ACK2_n & ((jx2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx2_n & ((jx3_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx3_n & ((jx1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoS_ACK7_n) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((BtoS_ACK0_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK2_n & ((jx2_n & ((jx1_n & ((jx0_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))) | (!jx0_n))) | (!jx1_n))) | (!jx2_n))))))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))))) | (!EMPTY_n & ((!FULL_n & ((stateG12_n & ((stateG7_0_n & ((BtoR_REQ0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ0_n & ((BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))) | (!BtoR_REQ1_n & ((BtoS_ACK7_n & ((StoB_REQ7_n & ((jx2_n) | (!jx2_n & ((jx3_n & ((jx1_n))) | (!jx3_n))))))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))))) | (!stateG7_0_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))))))))) | (!stateG12_n & ((BtoS_ACK7_n & ((StoB_REQ7_n))) | (!BtoS_ACK7_n & ((StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n & ((jx2_n & ((jx1_n & ((!jx0_n))) | (!jx1_n))) | (!jx2_n))))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n))))))))))))) | (!StoB_REQ7_n & ((BtoS_ACK6_n & ((StoB_REQ6_n))) | (!BtoS_ACK6_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK3_n)))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  StoB_REQ4_p = 0;
  StoB_REQ5_p = 0;
  StoB_REQ6_p = 0;
  StoB_REQ7_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoS_ACK4_p = 0;
  BtoS_ACK5_p = 0;
  BtoS_ACK6_p = 0;
  BtoS_ACK7_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  SLC2_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
  jx3_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  StoB_REQ4_p = StoB_REQ4_n;
  StoB_REQ5_p = StoB_REQ5_n;
  StoB_REQ6_p = StoB_REQ6_n;
  StoB_REQ7_p = StoB_REQ7_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoS_ACK4_p = BtoS_ACK4_n;
  BtoS_ACK5_p = BtoS_ACK5_n;
  BtoS_ACK6_p = BtoS_ACK6_n;
  BtoS_ACK7_p = BtoS_ACK7_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  SLC2_p = SLC2_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
  jx3_p = jx3_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
