module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hbusreq2, hlock2, hbusreq3, hlock3, hbusreq4, hlock4, hbusreq5, hlock5, hbusreq6, hlock6, hbusreq7, hlock7, hbusreq8, hlock8, hburst0, hburst1, hmaster0, hmaster1, hmaster2, hmaster3, hmastlock, start, decide, locked, hgrant0, hgrant1, hgrant2, hgrant3, hgrant4, hgrant5, hgrant6, hgrant7, hgrant8, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, stateG10_2, stateG10_3, stateG10_4, stateG10_5, stateG10_6, stateG10_7, stateG10_8, jx0, jx1, jx2, jx3);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v8455ab;
  wire v8455b5;
  wire v8455eb;
  wire v2678bee;
  wire v374a7cd;
  wire v3a5ccfd;
  wire v37286a2;
  wire v377e933;
  wire v3774a95;
  wire v3a59f5a;
  wire v375bb3a;
  wire v3a6d93d;
  wire v377514f;
  wire v3a69f36;
  wire v3a6f717;
  wire v39a4e84;
  wire v3a5bfc8;
  wire v377eea3;
  wire v373499c;
  wire v3a709da;
  wire v3724a10;
  wire v372a3dc;
  wire v3a5f8b2;
  wire v374efeb;
  wire v3772775;
  wire v375ea13;
  wire v3737b1a;
  wire v3a6fceb;
  wire v3732da0;
  wire v2678ca9;
  wire v8455c5;
  wire v376b03a;
  wire v8455dd;
  wire v1e379b9;
  wire v372d9a1;
  wire v3767091;
  wire v3727da5;
  wire v3773881;
  wire v372bc78;
  wire v3a2986b;
  wire v375fb93;
  wire v3a6d2d3;
  wire v3773536;
  wire v3a70a53;
  wire v374b237;
  wire v3a70f5f;
  wire v3737672;
  wire v35d37b1;
  wire v845605;
  wire v3746c8d;
  wire v3776483;
  wire v845601;
  wire v3725f3b;
  wire v3a7111f;
  wire v3738cfc;
  wire v3727fe3;
  wire v3a58cd5;
  wire v3747c3e;
  wire v3a6fe6c;
  wire v376575a;
  wire v374cd37;
  wire v375ad7d;
  wire v375c32d;
  wire v3a6aea2;
  wire v3732b63;
  wire v3a55672;
  wire v3a673d9;
  wire v37547f7;
  wire v377cc72;
  wire v374ac8a;
  wire v375356f;
  wire v3a2a770;
  wire v3a68016;
  wire v35ba2dd;
  wire v3729bf3;
  wire v3a58ddb;
  wire v3775c6e;
  wire v3a6f790;
  wire v3a6da08;
  wire v3777988;
  wire v3a551a4;
  wire v3a5e3d0;
  wire v3a70274;
  wire v3751460;
  wire v3773837;
  wire v373e98b;
  wire v3a71006;
  wire v3748332;
  wire v3730610;
  wire v3a6fd1a;
  wire v373c61e;
  wire v377a865;
  wire v375b659;
  wire v3a7017e;
  wire v3a5db06;
  wire v375b812;
  wire v3a6926b;
  wire v3a6ef8f;
  wire v3a64d96;
  wire v3732cdc;
  wire v372523e;
  wire v373e48c;
  wire v376a454;
  wire v374e20c;
  wire v3a6d70a;
  wire v376c12e;
  wire v3763898;
  wire v3a714bf;
  wire v372abb1;
  wire v376db87;
  wire v37323a5;
  wire v38075aa;
  wire v37717ac;
  wire v374b3af;
  wire a7afd8;
  wire v3722f85;
  wire v3762fcb;
  wire v372320e;
  wire v3729eeb;
  wire v3a6f275;
  wire v3768a1c;
  wire v377b159;
  wire v37533d5;
  wire v3a67370;
  wire v37544fa;
  wire v3a5754b;
  wire v372d7ed;
  wire v376ef46;
  wire v3a714cf;
  wire v37594d4;
  wire v3726a86;
  wire v3a6b19d;
  wire v374cfee;
  wire v37719b4;
  wire v374bc77;
  wire v3753b90;
  wire v3808fc2;
  wire v39a4dd6;
  wire v3a55395;
  wire v3775f25;
  wire v3a54b77;
  wire v3a712a7;
  wire v377afaa;
  wire v3778c9a;
  wire v3a6ec08;
  wire v3a6f337;
  wire v845603;
  wire v3766cf9;
  wire v3a70a28;
  wire v3760a9d;
  wire v20d166d;
  wire v3a70c98;
  wire v3741d83;
  wire v3754afa;
  wire v376bb81;
  wire v3751db0;
  wire v3a66447;
  wire v3a53f4c;
  wire v3a6fbf7;
  wire v3725395;
  wire v3776386;
  wire v3750c50;
  wire v3746487;
  wire v373da59;
  wire v373d8d8;
  wire v3a66335;
  wire v375145d;
  wire v372deb9;
  wire v3727a2b;
  wire v3809da1;
  wire v372a20c;
  wire v3a6a089;
  wire v3a71071;
  wire v373b87c;
  wire v373913e;
  wire v3756cee;
  wire v377d95a;
  wire v377b253;
  wire v376b0fd;
  wire v37484de;
  wire v3a5e9a8;
  wire v374612b;
  wire v377bd5c;
  wire v37395a4;
  wire v37399d0;
  wire v906a66;
  wire v3727d4d;
  wire v3751285;
  wire v3747453;
  wire v3762a54;
  wire v374361e;
  wire v3a63166;
  wire v3776db0;
  wire v3764238;
  wire v3760233;
  wire v37698ab;
  wire c8f3d0;
  wire v3750012;
  wire v3773e52;
  wire v37530cf;
  wire v3728333;
  wire v37753f2;
  wire v3a6e8a4;
  wire v3a6a66f;
  wire v374821f;
  wire v3740212;
  wire v3a70255;
  wire v3a620ef;
  wire v3a6fd50;
  wire v3779f1c;
  wire v373da95;
  wire v3a594ab;
  wire v3a697a5;
  wire v377051a;
  wire v3a6f2f2;
  wire v3746368;
  wire v3a5eb73;
  wire v3730b6d;
  wire v3a5688f;
  wire v3743d8b;
  wire v3739c68;
  wire v3a6af93;
  wire v3a5f413;
  wire v3a70a34;
  wire v377d52e;
  wire v373e32a;
  wire v3a59eb3;
  wire v374cbc0;
  wire v375c278;
  wire v3766de9;
  wire v3768c53;
  wire v3a5e7be;
  wire v3a5858c;
  wire v3729c71;
  wire v3a62615;
  wire v38072fd;
  wire v3a6a19b;
  wire v373790d;
  wire v376ae9f;
  wire v374ceec;
  wire v374aa73;
  wire v3740415;
  wire v3a6f428;
  wire v37748e5;
  wire v3a66e91;
  wire v3a56e5e;
  wire v3770ae6;
  wire v3753b5e;
  wire v377b84e;
  wire v373f7b7;
  wire v3768870;
  wire v3763186;
  wire v3728f3a;
  wire v374a3b8;
  wire v377e9bb;
  wire v3a6f8ae;
  wire v374cbe2;
  wire v3a5ad17;
  wire v3a6f12b;
  wire v374457b;
  wire v373efdf;
  wire v3a5e1b7;
  wire v3763e46;
  wire v3a5f586;
  wire v37684c0;
  wire v373f9ad;
  wire v3765370;
  wire v3769e7f;
  wire v373fd4c;
  wire v3a6bf3c;
  wire v3777517;
  wire v360d00f;
  wire v3741736;
  wire v3a5f546;
  wire v3778f25;
  wire v3739c89;
  wire v373b241;
  wire v3a6f6f8;
  wire v373e491;
  wire v3a6d6b8;
  wire v3a5610f;
  wire v3a63a2a;
  wire v3809de2;
  wire v3a6fa76;
  wire v3a5b4de;
  wire v3a6cb62;
  wire v3a6512b;
  wire v37781a8;
  wire v372e559;
  wire v3771b83;
  wire v3a5b9d6;
  wire v3a5a47b;
  wire v3a6fbc7;
  wire v3a5bc4f;
  wire v376ea88;
  wire v3747917;
  wire v1e37916;
  wire v3773bf5;
  wire v3a5c484;
  wire v372c903;
  wire v3a715ae;
  wire v3a6c1ec;
  wire v37355ce;
  wire v3a703cd;
  wire v372c3b9;
  wire v3a55773;
  wire v3a5c11a;
  wire v374d13d;
  wire v3772021;
  wire v3a6e9b0;
  wire v373f2d2;
  wire v3a705aa;
  wire b30936;
  wire v3741b49;
  wire v376ad73;
  wire v374beb6;
  wire v376a054;
  wire v3a556c2;
  wire v377fc58;
  wire v372954c;
  wire v3a63f9a;
  wire a0a219;
  wire v8637a5;
  wire v3a63699;
  wire v3734fba;
  wire v3a55466;
  wire v374b4c5;
  wire v377ebf3;
  wire v372b721;
  wire v3a58219;
  wire v376f92f;
  wire v3a70acb;
  wire v377576e;
  wire v37680a7;
  wire v3a5cb0e;
  wire v3a6f5ae;
  wire v3a701fe;
  wire v37425a8;
  wire v375f985;
  wire v3a7100a;
  wire v374373c;
  wire v3776691;
  wire v3a708bc;
  wire v3765443;
  wire v3a6f4d6;
  wire v37357d0;
  wire v375e5ed;
  wire v37349e4;
  wire v2092b5f;
  wire v376abcc;
  wire v3a5ee7a;
  wire v377d9fa;
  wire v373121b;
  wire v3776d4b;
  wire v375469c;
  wire v3772bb1;
  wire v37551b2;
  wire v3748d63;
  wire v3769e10;
  wire v3a6165b;
  wire v3767153;
  wire v377ace4;
  wire v377696e;
  wire v377a7ee;
  wire v377e539;
  wire v3728723;
  wire v37283ea;
  wire v3744bac;
  wire v3a70895;
  wire v372b5af;
  wire v3a706a2;
  wire v3777178;
  wire v3771507;
  wire v377d280;
  wire v3a543c5;
  wire v374dbdf;
  wire v3a68183;
  wire v3740052;
  wire v375e22b;
  wire v375a293;
  wire v325c976;
  wire v3a5b614;
  wire v373cf3a;
  wire v3a637e0;
  wire v3732706;
  wire v3765261;
  wire v3773a5b;
  wire v37690ea;
  wire v376e5fe;
  wire v3809ec3;
  wire v3764a07;
  wire v374fc57;
  wire v3a57750;
  wire v3a70e79;
  wire v3761553;
  wire v3a7162a;
  wire a16ae7;
  wire v3a7099b;
  wire v375b18e;
  wire v373031f;
  wire v376a149;
  wire v3a7073b;
  wire v3764601;
  wire v3737647;
  wire v3725b27;
  wire v373dec1;
  wire v2619ada;
  wire v375859f;
  wire v3766e4a;
  wire v377476b;
  wire v3774c77;
  wire v372a939;
  wire v3731230;
  wire v376b5ad;
  wire v3a6d4bf;
  wire v37502ca;
  wire v3726344;
  wire v37778a2;
  wire v3a6fb81;
  wire v38073e8;
  wire v3a5915c;
  wire v3762158;
  wire v3753c73;
  wire v1e37523;
  wire v3a667cf;
  wire v3764dac;
  wire v3a5aa5c;
  wire v3a708d4;
  wire v3745b36;
  wire v3a65c29;
  wire v3746f37;
  wire v3772db0;
  wire v3a5ad13;
  wire v3733cca;
  wire v3a6eefe;
  wire v375d8fb;
  wire v3a70452;
  wire v3a70910;
  wire v3a5f7f3;
  wire v3a6ad59;
  wire v3a6a82a;
  wire v3727703;
  wire v3a703b9;
  wire v37436a8;
  wire v3a7011e;
  wire v373ce84;
  wire v1e37dfd;
  wire v375a166;
  wire v37285eb;
  wire v37264c9;
  wire v1e374ce;
  wire v373c856;
  wire v37442e1;
  wire v37728c2;
  wire v3a6f9e4;
  wire v3a6ef4d;
  wire v3a6f44e;
  wire v375ae91;
  wire v3a70f7a;
  wire v37468e5;
  wire v3a6c5fc;
  wire v37731c3;
  wire v3a58102;
  wire v373bd6c;
  wire v3737bff;
  wire v3756899;
  wire v37566f4;
  wire v3722f58;
  wire v3737f89;
  wire v3a6c2d4;
  wire v3741cd7;
  wire v3741325;
  wire v3a6ff2d;
  wire v377550d;
  wire v3779746;
  wire v376b57f;
  wire v377d6d3;
  wire v376d05f;
  wire v373291e;
  wire v3737909;
  wire v377e825;
  wire v3a713e7;
  wire v376dc6f;
  wire v375d3a2;
  wire v374b0fb;
  wire v376b397;
  wire v3a6eaff;
  wire v3a66ab2;
  wire v3a5e030;
  wire v3a5e618;
  wire v3746da7;
  wire v374294c;
  wire v375ff99;
  wire v3722fb7;
  wire v3a60276;
  wire v372b5c0;
  wire v3739b6a;
  wire v380937f;
  wire v3a7084f;
  wire v3737ceb;
  wire v3758d1e;
  wire v3808f5d;
  wire v3753903;
  wire v380678d;
  wire v373ea10;
  wire v3a6f9ae;
  wire v37393ad;
  wire v3a67cd1;
  wire v3809194;
  wire v372e3ea;
  wire v37791a5;
  wire v3a6f03e;
  wire v37337d2;
  wire v3a6ea3b;
  wire v3754603;
  wire v3a6fe1b;
  wire v3a689e5;
  wire v3729597;
  wire v3a71175;
  wire v377e9d7;
  wire v374998d;
  wire v3778754;
  wire v3a60280;
  wire v377940a;
  wire v3a6620b;
  wire v3a7163f;
  wire v3a70db6;
  wire v37316c9;
  wire v377e241;
  wire v3735539;
  wire v3a6eb5c;
  wire v3767ff6;
  wire v37550bd;
  wire v3a70301;
  wire v374e650;
  wire v3725e9a;
  wire v3a59d6b;
  wire v37716e1;
  wire v3735350;
  wire v3a71545;
  wire v37725c6;
  wire v3a710de;
  wire v3742005;
  wire v3746696;
  wire v375987e;
  wire v3a70e5b;
  wire v374641d;
  wire v3748ba4;
  wire v374ed57;
  wire v37308a9;
  wire v375dcd5;
  wire v3a6fb9d;
  wire v3a702f8;
  wire v376bfc3;
  wire v38074bc;
  wire v3807341;
  wire v3769e3a;
  wire v372cfd2;
  wire v3757c10;
  wire v374b3e2;
  wire v3a70c95;
  wire v3a5bb42;
  wire v3731164;
  wire v373c005;
  wire v3747452;
  wire cd0aed;
  wire v375cc28;
  wire v37486c2;
  wire v37543ae;
  wire v3a6c2ad;
  wire aef673;
  wire v3727807;
  wire v3a65f32;
  wire v372313c;
  wire v3760d16;
  wire v372f759;
  wire v376ab01;
  wire v3a687e0;
  wire v375cda2;
  wire v3a70925;
  wire v3a704de;
  wire v375b3be;
  wire v372cb99;
  wire v37402cd;
  wire v376b0f2;
  wire v3a70f64;
  wire v373d0af;
  wire v3a6a4cf;
  wire v3766e8b;
  wire v3a57f8b;
  wire v376d8c1;
  wire v373e031;
  wire v3a5ab85;
  wire v3a6f4fd;
  wire v376ae41;
  wire v3a56494;
  wire v374503d;
  wire v374c900;
  wire v3a6b8cc;
  wire v375a4ba;
  wire v3a62bcf;
  wire v3a6db7f;
  wire v3723220;
  wire v3a6062e;
  wire v374c9d1;
  wire v3a67d7b;
  wire v3a5e8ac;
  wire v3756ce5;
  wire v375f5f0;
  wire v374ea7d;
  wire v3a64b1e;
  wire v3a6fb14;
  wire v35b779f;
  wire v3a6f338;
  wire v3745b20;
  wire v3762388;
  wire v374aa90;
  wire v3a645b4;
  wire v3a6358e;
  wire v3a651fb;
  wire v37314fc;
  wire v3a5bbc2;
  wire v3a6a236;
  wire v372df43;
  wire v375d10e;
  wire v3a6fbc5;
  wire v376d7c6;
  wire v375bdaf;
  wire v3753d9d;
  wire v376ef4f;
  wire v37520ad;
  wire v3a6dc91;
  wire v3758ff8;
  wire v37576f6;
  wire v3807740;
  wire v910050;
  wire v373c377;
  wire v3a6bada;
  wire v3739635;
  wire v3a7005e;
  wire v3a71566;
  wire v3a6f0f2;
  wire v3a71684;
  wire v360bc71;
  wire v3740404;
  wire v377ecd4;
  wire v3776852;
  wire v3a710dd;
  wire v37617ad;
  wire v3a6a546;
  wire v374283c;
  wire v3a70f43;
  wire v3a57214;
  wire v3807ac3;
  wire v376cf3f;
  wire v3a6f139;
  wire b5f474;
  wire v373bc30;
  wire v3a5524c;
  wire v3a6f907;
  wire v3807670;
  wire afadd1;
  wire v37325ed;
  wire v372c467;
  wire v3772d0e;
  wire v3a71556;
  wire v3735ba1;
  wire v3a6a367;
  wire v3740ff7;
  wire v3776d3e;
  wire v37766d3;
  wire bdbe8b;
  wire v37279df;
  wire v3a71112;
  wire v37315ae;
  wire v3a6f407;
  wire v377133f;
  wire v3809b0a;
  wire v3751e7c;
  wire v377bd76;
  wire v372d691;
  wire v3a68170;
  wire v374c256;
  wire v375cf55;
  wire v3a7019a;
  wire v37522ea;
  wire v376e5d2;
  wire v3778a0a;
  wire v3a70eba;
  wire v3755c19;
  wire v3a6f621;
  wire v373894a;
  wire v374067b;
  wire v376374e;
  wire v3a6be38;
  wire v376f0cd;
  wire v37435b9;
  wire v3a71593;
  wire v38067ba;
  wire v3a6fa18;
  wire v3a59d00;
  wire v3a6430c;
  wire v376a87b;
  wire v37599cb;
  wire v377b27b;
  wire v3a6f77e;
  wire v3734f70;
  wire v3754422;
  wire v377e2ae;
  wire v37237cd;
  wire v37435f7;
  wire v3760353;
  wire v3a64987;
  wire v373dde1;
  wire v3768d6c;
  wire v3a55b5b;
  wire v377c0c3;
  wire v372ce1e;
  wire v3a61820;
  wire v3a6f3c2;
  wire v374544d;
  wire v376fe68;
  wire v376906d;
  wire v3a6ad8b;
  wire v3a6f588;
  wire v3762cc4;
  wire v29256ae;
  wire v3a70e10;
  wire v3a640ab;
  wire v3737e04;
  wire v375ff0d;
  wire v37629b4;
  wire v374284d;
  wire v3a6bc0e;
  wire v3a69758;
  wire v37711ec;
  wire v3734583;
  wire v374be73;
  wire v37243ac;
  wire v3a6f600;
  wire v372cdd4;
  wire v376e7c1;
  wire v3730f97;
  wire v3a5f0f0;
  wire v3a5e65e;
  wire v3a6ffb1;
  wire v3760860;
  wire v3764494;
  wire v3a62229;
  wire v3a6f4ea;
  wire v375571e;
  wire v373a7dc;
  wire v376a59f;
  wire v3761340;
  wire v377e0a4;
  wire v3a66d3e;
  wire v3769325;
  wire v3724547;
  wire v3a608b8;
  wire v3a5def7;
  wire v3a5874e;
  wire v3776c6e;
  wire v37388f6;
  wire v3775709;
  wire v3808e56;
  wire v3a6a720;
  wire v37705be;
  wire v3741cd4;
  wire v3777610;
  wire v3a2986f;
  wire v3a6f851;
  wire v373dc55;
  wire v377dc60;
  wire v372ce4a;
  wire v3744657;
  wire v3a6ccc6;
  wire v3741cc4;
  wire v3764e3f;
  wire v3a70f6d;
  wire v3761f13;
  wire v373ef28;
  wire v1e37ec1;
  wire v3a648f6;
  wire v3a573d2;
  wire v3a71329;
  wire v3a6fc98;
  wire v3725f3e;
  wire v3a62c49;
  wire v3a70c10;
  wire v377bbbd;
  wire v3745b60;
  wire v37396de;
  wire v374a877;
  wire v3a6d81e;
  wire v3a6190f;
  wire v376f0a0;
  wire v3a6ed4c;
  wire v3753073;
  wire v3a706d2;
  wire v373cd0a;
  wire v373f24b;
  wire v3732208;
  wire v372f235;
  wire v372787e;
  wire v377dbd3;
  wire v3761ac7;
  wire v375df95;
  wire v3740bb4;
  wire v3778cdb;
  wire v3747193;
  wire v3727420;
  wire v3a703c5;
  wire v3a6f4bd;
  wire v3a636a7;
  wire v3755ed8;
  wire v3a6fc01;
  wire v376faab;
  wire v373eaf6;
  wire v3a6ad04;
  wire v374cda0;
  wire v3a6de95;
  wire v3a70c55;
  wire v377c3ad;
  wire v3a70e6b;
  wire v372c257;
  wire v373d9b3;
  wire v3736113;
  wire v3a6d686;
  wire v9ca2d6;
  wire v3748ab9;
  wire v3a70bfb;
  wire v3a63f80;
  wire v3735d01;
  wire v3a55076;
  wire v3807174;
  wire v37256c0;
  wire v3a70a3d;
  wire v37676b6;
  wire v3752d7a;
  wire v375b5ca;
  wire v3768e0e;
  wire v3751e62;
  wire v3765008;
  wire v3a6eedf;
  wire v37297f9;
  wire v376af8e;
  wire v38069c0;
  wire v377ccb7;
  wire v37614a9;
  wire v372ed5f;
  wire v3753804;
  wire v3a7038a;
  wire v3a578af;
  wire v23fe343;
  wire v375bf36;
  wire v3734e23;
  wire v3a6fc58;
  wire v37514dd;
  wire v373d238;
  wire v375ae0a;
  wire v3a6f269;
  wire dc6ab1;
  wire v376636b;
  wire v3751dcc;
  wire v375485b;
  wire v3a579d1;
  wire v3a64474;
  wire d284a6;
  wire v3a66538;
  wire v3728346;
  wire v377e087;
  wire v37344a0;
  wire v3733360;
  wire v376b795;
  wire v3a5b885;
  wire v3733716;
  wire v37321c2;
  wire v372d48a;
  wire v3a66f3e;
  wire v3a6c44c;
  wire v372ad5d;
  wire v3a5df87;
  wire v2ff9348;
  wire v374c3d0;
  wire v3a605af;
  wire v3a5f154;
  wire v3a6b18c;
  wire v374f89b;
  wire v3a5fe5e;
  wire v3a615bb;
  wire v37721eb;
  wire v3a5a8c3;
  wire v372fe1b;
  wire v374a096;
  wire v374663d;
  wire v3751c77;
  wire v3a71600;
  wire v3a7045f;
  wire v37748f0;
  wire v3a6ef06;
  wire v3a6ff97;
  wire v3775606;
  wire v3a6624e;
  wire v3a676c6;
  wire v377cdbe;
  wire v3724667;
  wire v3756205;
  wire v3a70b5e;
  wire v3a6fb0c;
  wire v3a70ef2;
  wire v372df47;
  wire v374ec84;
  wire v375899b;
  wire v373d5d6;
  wire v373f622;
  wire v3747569;
  wire v374e43d;
  wire v3a625f8;
  wire v3a648d0;
  wire v3a6f377;
  wire v3723635;
  wire b21e3c;
  wire v377419a;
  wire v3729b48;
  wire v3a6aee6;
  wire v3a6fa78;
  wire v3a6f134;
  wire v37647fc;
  wire v3a6ab14;
  wire v37270dc;
  wire v372d733;
  wire v373d239;
  wire v23fd9cb;
  wire v376b4d4;
  wire v3754445;
  wire v3774372;
  wire v3a59c5e;
  wire v372da0b;
  wire v37250b1;
  wire v376efcf;
  wire v376015e;
  wire v3a6ffa0;
  wire v360d18d;
  wire v3746d07;
  wire v375aeca;
  wire v37305b9;
  wire v3a70414;
  wire v377c214;
  wire v3733690;
  wire v3765f13;
  wire v3a70c2e;
  wire v3754d21;
  wire a012c1;
  wire v372c18e;
  wire v3a5ae1b;
  wire v373fe6f;
  wire v3756c83;
  wire v3754f2e;
  wire v377e87e;
  wire v3a70f32;
  wire v372eaf0;
  wire v3771203;
  wire v3a60ba3;
  wire v3a55aa8;
  wire v3777a66;
  wire v3a70f3d;
  wire v3726054;
  wire v3a6fefc;
  wire v37522e4;
  wire v3760a1c;
  wire v377eee2;
  wire v3a6fc89;
  wire v376a9aa;
  wire v37653bf;
  wire v37737f9;
  wire v37296db;
  wire v3752bcc;
  wire d2819e;
  wire v37773a2;
  wire v3a61f82;
  wire v372ee70;
  wire v3a708a8;
  wire v3a6beb6;
  wire v3768c4c;
  wire v374f5e3;
  wire v3378e07;
  wire v373b92c;
  wire v3764bd6;
  wire v3779f43;
  wire v376e9e9;
  wire v3a6fe09;
  wire v3a62f06;
  wire v3739078;
  wire v3758bbd;
  wire v3a707f2;
  wire v37315d0;
  wire v376e0b6;
  wire v3768858;
  wire v3a6fef0;
  wire v3743156;
  wire v374c28e;
  wire v3a5fbcb;
  wire v3809ab5;
  wire v374952b;
  wire v3a6fb0a;
  wire v37518f0;
  wire v372e49a;
  wire v3763c59;
  wire v3743038;
  wire v373df5c;
  wire v3a7138f;
  wire v3741172;
  wire v374151e;
  wire v3a5d2f1;
  wire v2092c08;
  wire v3726abd;
  wire v37688a5;
  wire v3759020;
  wire v37444d0;
  wire v376faea;
  wire v3739e55;
  wire v2925c39;
  wire v3750d37;
  wire v3a6f441;
  wire v3737a06;
  wire v3737103;
  wire v3a580e3;
  wire v374510a;
  wire v376f032;
  wire v3747bc9;
  wire v37293c3;
  wire v373a58c;
  wire v3a6ef3e;
  wire v377360d;
  wire v374b83f;
  wire v376b164;
  wire v3a6841c;
  wire v3a6e7b3;
  wire v3761785;
  wire v360d016;
  wire v372bffc;
  wire v3a598b7;
  wire v3a6f83c;
  wire v3757772;
  wire v3a6fe18;
  wire v3752ade;
  wire v372d9e8;
  wire v3a706de;
  wire v376fe00;
  wire v3773201;
  wire v3757490;
  wire v37654e1;
  wire v375068c;
  wire v374d42c;
  wire v3a6eb3c;
  wire v374177f;
  wire v39a4ed6;
  wire v3774a77;
  wire v374c5e2;
  wire c61b3c;
  wire v3a709a3;
  wire v3a6eebf;
  wire v37613a8;
  wire v3776b18;
  wire v3a5b90b;
  wire v91a14c;
  wire v37bfc4d;
  wire v3a6fad2;
  wire v3a7031b;
  wire v3a6fcfa;
  wire v3a61fc9;
  wire v3a700da;
  wire v37746d7;
  wire v3722f88;
  wire v3741797;
  wire v1e379e9;
  wire v373ec8e;
  wire v3a6f9f9;
  wire v3764e37;
  wire v3a6f922;
  wire v37579c1;
  wire v372650c;
  wire v3779647;
  wire v37709c5;
  wire v3a71437;
  wire v3a61f3c;
  wire v376ebe6;
  wire v37634d8;
  wire v3741922;
  wire v3a68dab;
  wire v377a57a;
  wire v3a6b72a;
  wire v8ac028;
  wire v325c93a;
  wire v3a6307d;
  wire v3741365;
  wire v376537c;
  wire v37369df;
  wire v3779c7e;
  wire v377d789;
  wire v3a70b2d;
  wire v376f62e;
  wire v374ebac;
  wire v3a67dc7;
  wire v3a62abc;
  wire v3768ec7;
  wire v373da8d;
  wire v3773c36;
  wire v3750ebc;
  wire v3760c3c;
  wire v3a700a8;
  wire v374a296;
  wire v3a70672;
  wire v3a62396;
  wire v3a6f09b;
  wire v372eabb;
  wire v3760d14;
  wire v376cfaa;
  wire v377fbbf;
  wire v374b9e6;
  wire v3a652c7;
  wire v3764818;
  wire v3753f82;
  wire v374cab1;
  wire v375a9d7;
  wire v3a6a63c;
  wire v913004;
  wire v3a704b8;
  wire v3758c4d;
  wire v374dd5f;
  wire v37771cc;
  wire v3a563aa;
  wire v3759ca5;
  wire v3732dc6;
  wire v3765a79;
  wire v373a902;
  wire v3a6f786;
  wire v375e23b;
  wire v376a129;
  wire v3a6f000;
  wire v3a6fdc0;
  wire v3767261;
  wire v3a6fb41;
  wire v3a58792;
  wire v3a6ebc5;
  wire v3a70a54;
  wire v3761b90;
  wire v3a658ad;
  wire v3806e35;
  wire v375798a;
  wire v3768091;
  wire v374d6bd;
  wire v37792d9;
  wire v3a701d8;
  wire v3739be4;
  wire v372b163;
  wire v3a6fb45;
  wire v922f0a;
  wire v3746be0;
  wire v372b2ef;
  wire v3743287;
  wire v375f6f6;
  wire v3763788;
  wire v3a6f133;
  wire v3741c03;
  wire v37462ca;
  wire v3773b2f;
  wire v3746cdc;
  wire v3a6ffe7;
  wire v3a6a580;
  wire v3a6bef4;
  wire v3a6caa5;
  wire v3a5e291;
  wire v3a5f147;
  wire v8b397d;
  wire v3a703a1;
  wire v3751ad8;
  wire v373f1e4;
  wire v1e37762;
  wire v375fd29;
  wire v3734b20;
  wire v3378f5d;
  wire v380732c;
  wire v3a62e20;
  wire v3a6bb4b;
  wire v3a6f77b;
  wire v3a5f5d0;
  wire v377f108;
  wire v3750fea;
  wire v372dee5;
  wire v377f4bb;
  wire v37690db;
  wire v3749e1c;
  wire v37403cf;
  wire v3757568;
  wire v3a6a36d;
  wire v3723a30;
  wire v372e77b;
  wire v3a5e8a1;
  wire v3a5d431;
  wire v3a7142e;
  wire v3779879;
  wire v37544ab;
  wire v374cd43;
  wire v3a6f9a7;
  wire v3a70dfd;
  wire v3770362;
  wire v3a69a06;
  wire v373d0e1;
  wire v3a66151;
  wire v3a6a259;
  wire v3a5bead;
  wire v3a5f4e1;
  wire v37753e0;
  wire v376a2c0;
  wire v1e3773a;
  wire v39ea663;
  wire v3752bbd;
  wire v3a71493;
  wire v373a79f;
  wire v3808904;
  wire v372d0db;
  wire v8455e1;
  wire v37771a2;
  wire v3a70521;
  wire v3808ed2;
  wire v3742322;
  wire v3a5958e;
  wire v3752248;
  wire v3a6b2ea;
  wire v3a70907;
  wire v37744e3;
  wire v3767a42;
  wire v376629b;
  wire v375c7b0;
  wire v375a68d;
  wire v3771fe5;
  wire v292500d;
  wire v8455e7;
  wire v3a58c00;
  wire v373ca17;
  wire v3730a0f;
  wire v3a5fcfc;
  wire v3a7147e;
  wire v376c211;
  wire v373fe5e;
  wire v374176c;
  wire v373f042;
  wire v3739702;
  wire v3a6450a;
  wire v3760e78;
  wire v3a558ce;
  wire v3a6909a;
  wire v3a6eff4;
  wire v3a6fe99;
  wire v3764ca7;
  wire v375e70f;
  wire v9c9282;
  wire v3a6fbc6;
  wire v3a674d5;
  wire v373d825;
  wire v3a6931f;
  wire v3a6fc5a;
  wire v3730f5d;
  wire v373e87e;
  wire v3a70cef;
  wire d99853;
  wire v3a6bddf;
  wire v375b48b;
  wire v374b08d;
  wire v3a71618;
  wire v3767537;
  wire v3a70f05;
  wire v3767d2c;
  wire v376ebc7;
  wire v3775379;
  wire v3a708ff;
  wire v3769bf7;
  wire v3746bdb;
  wire v8455d7;
  wire v3a5a496;
  wire v3745b85;
  wire v39a5381;
  wire v39a537f;
  wire v3a70a83;
  wire v3a67241;
  wire v3a6a939;
  wire v3730dea;
  wire v37566b2;
  wire v373a27c;
  wire v3a69555;
  wire v3a59da9;
  wire v3a6f056;
  wire v3733a6c;
  wire v37643ee;
  wire v3a69ad1;
  wire v3a64235;
  wire v3a6edfa;
  wire v3755019;
  wire v374362e;
  wire v374b204;
  wire v3764437;
  wire v37505e1;
  wire v373db51;
  wire v377f384;
  wire v3732fec;
  wire v3727e80;
  wire v3a555f9;
  wire v3a65a34;
  wire v3a5d74e;
  wire v3a676d6;
  wire v3756954;
  wire v374c120;
  wire v37545b7;
  wire v373aaf0;
  wire v3779cb5;
  wire v375b990;
  wire v3a70a29;
  wire v374cab9;
  wire v3a5d994;
  wire v376a752;
  wire v3a6fbfd;
  wire v3a563ad;
  wire v3758079;
  wire v373bdac;
  wire v37674c1;
  wire v374636c;
  wire v3768695;
  wire v3a70157;
  wire v374db33;
  wire v372c834;
  wire v376d06c;
  wire v3744deb;
  wire v3740171;
  wire v37457fb;
  wire v3733b37;
  wire v3a6f2c9;
  wire v3746b4f;
  wire v373e2c3;
  wire v3a6980b;
  wire v3a663ef;
  wire v3a6f7bf;
  wire v37334c5;
  wire v3760eeb;
  wire v3726464;
  wire v3768ecc;
  wire v3742851;
  wire v376626a;
  wire v3727fcb;
  wire v373930f;
  wire v375a754;
  wire v3a707e7;
  wire v3754f93;
  wire v3a67471;
  wire v3739f49;
  wire v3a6af87;
  wire v375a4a9;
  wire v376b21a;
  wire v372bfcc;
  wire v3730755;
  wire v375a4fa;
  wire v3a6c803;
  wire v3a714cd;
  wire v3751734;
  wire v3a6f3d8;
  wire v374c3f2;
  wire v3a702aa;
  wire v3737d44;
  wire v3777f6e;
  wire v373e70e;
  wire v377027e;
  wire v3764c0d;
  wire v375134f;
  wire v3a71315;
  wire v3734862;
  wire v3730dc1;
  wire v3778a55;
  wire v3a70424;
  wire v3767183;
  wire v3769d3d;
  wire v3a67131;
  wire v3a6299c;
  wire v3a5e687;
  wire v374aa82;
  wire v3755e66;
  wire v3779c8d;
  wire v3a6f731;
  wire v3a54789;
  wire v3779e21;
  wire v374f8b5;
  wire v376c176;
  wire v3a6e584;
  wire v3772c0a;
  wire v37648fb;
  wire v3727a82;
  wire v3771dc9;
  wire v3730766;
  wire v3747cfc;
  wire v3a6fd35;
  wire v3a6e40b;
  wire v372c2da;
  wire v37757cb;
  wire v3747afb;
  wire v3a5b25b;
  wire v3a66db2;
  wire v3727af8;
  wire v3745ab5;
  wire v3747ec9;
  wire v373ba38;
  wire v39a4e19;
  wire v3749f51;
  wire v374b07c;
  wire v372410a;
  wire v3771733;
  wire v38071a9;
  wire v3a605b5;
  wire v3a62329;
  wire v372af67;
  wire v3a5c823;
  wire v374af6a;
  wire v37410d9;
  wire v376f0c1;
  wire v373bd24;
  wire v3a6f4d3;
  wire v3760ef5;
  wire v37481c3;
  wire v373d9e5;
  wire v3a66bdb;
  wire v372cb88;
  wire v3a6f436;
  wire v3a70334;
  wire v3a6e591;
  wire v376498a;
  wire v3a6ec94;
  wire v3a5ae2f;
  wire v375a613;
  wire v37526a0;
  wire v377e582;
  wire v3a6f2a4;
  wire v37773a9;
  wire v3a5c4d5;
  wire v3770bb9;
  wire v3a558c5;
  wire v3a5ab84;
  wire v3763b9e;
  wire v3738253;
  wire v372eafa;
  wire v3731596;
  wire v3744b1b;
  wire v1e374cc;
  wire v3725a56;
  wire v3770c9d;
  wire v3a5e2ee;
  wire v3a704f8;
  wire v3a6c80b;
  wire v376e643;
  wire v377696a;
  wire v3a6251b;
  wire v3a655c2;
  wire v373a66d;
  wire v37362ea;
  wire v3a53877;
  wire v3774c11;
  wire v3a6d922;
  wire v3a6b2ef;
  wire v374a891;
  wire v37300b7;
  wire v3a56338;
  wire v377fc15;
  wire v3736a92;
  wire v3a6900b;
  wire v37349d3;
  wire v3759fb4;
  wire v37323a1;
  wire v3766484;
  wire v376a941;
  wire v377a2e1;
  wire v38092f5;
  wire v373a0f4;
  wire v3735bf3;
  wire v3a61c51;
  wire v3a5e1e4;
  wire v3a706b3;
  wire v372525e;
  wire v3a70cf2;
  wire v377a9e2;
  wire v3778657;
  wire v3a71576;
  wire v373b838;
  wire v37287bd;
  wire v3a62d48;
  wire ca1199;
  wire v3a6fdae;
  wire v3726bff;
  wire v3a67629;
  wire v3728eeb;
  wire v8df61b;
  wire v3726f6c;
  wire v3a6ff7d;
  wire v372d02d;
  wire v3a56ccf;
  wire v37422d8;
  wire v374473f;
  wire v37470eb;
  wire v337904e;
  wire v376f455;
  wire v376e611;
  wire v3726f97;
  wire v3a5f9ad;
  wire v2092b01;
  wire v3734247;
  wire v3753fe0;
  wire v374c4bc;
  wire v3a5b41c;
  wire v3a60aca;
  wire v373d5dc;
  wire v373ad68;
  wire ba83e3;
  wire v3a6ad93;
  wire v377258d;
  wire v372f3fc;
  wire v3a6fb44;
  wire v375df97;
  wire v373436a;
  wire v374ea19;
  wire v23fe353;
  wire v3761287;
  wire v3756f8a;
  wire v292556b;
  wire v377e897;
  wire v3a6810b;
  wire v376539b;
  wire v3747797;
  wire c4d63a;
  wire v3768fc7;
  wire v377c174;
  wire v3a6eb54;
  wire v3a707ab;
  wire v3a64bcf;
  wire v373ac50;
  wire v3734bf8;
  wire v3a708d3;
  wire v3759044;
  wire v372c37f;
  wire v3a57b60;
  wire v3a5a01a;
  wire v3731be6;
  wire v374d542;
  wire v3740140;
  wire v37761b6;
  wire v37579a9;
  wire v3770bd9;
  wire v3a6e516;
  wire v377b779;
  wire v374933f;
  wire v3765b08;
  wire v3753ff9;
  wire v3a6fff9;
  wire v373ab9e;
  wire v3a68c0e;
  wire v375bf96;
  wire v3744104;
  wire v3a65a19;
  wire v3744f86;
  wire v372b96c;
  wire v3a6f09c;
  wire v3a704c2;
  wire v3729214;
  wire v3758fe4;
  wire v374f9c5;
  wire v374b2f7;
  wire v3a5ec91;
  wire v3a6fc21;
  wire v3a578e2;
  wire v37596d5;
  wire v372cbfc;
  wire v373428e;
  wire v37778cf;
  wire v372abc8;
  wire v373c81c;
  wire v377af0a;
  wire v377408e;
  wire v375e7cc;
  wire v3a6fbb4;
  wire v3a59dc4;
  wire v3770c4c;
  wire v3a5bb98;
  wire v3a6f4ef;
  wire v39a53a4;
  wire v37416c8;
  wire v3a685e1;
  wire v3758174;
  wire v3742dfb;
  wire v37618ef;
  wire v3a6fc03;
  wire v372b1e6;
  wire v3734918;
  wire v3a657bf;
  wire v3a71389;
  wire v3a6962d;
  wire v3754871;
  wire v3a70403;
  wire v3741cb9;
  wire v3757663;
  wire v3a55d41;
  wire v39a4d88;
  wire v373c4e4;
  wire v375b2e5;
  wire v3762de1;
  wire v3a60205;
  wire v3a6e9a4;
  wire v3777fc5;
  wire v374a044;
  wire v3a63b90;
  wire v3737416;
  wire v3a6443d;
  wire v3a6eb86;
  wire v3756ebb;
  wire v3a5f41d;
  wire v3738ff9;
  wire v3a70114;
  wire v375199d;
  wire v3a6f255;
  wire v3807a32;
  wire v372d60f;
  wire v374cd18;
  wire v37432d3;
  wire v377eac7;
  wire v3a7165b;
  wire v3758a02;
  wire v37758ad;
  wire v3a6fdd8;
  wire v3a710ba;
  wire v3a6ab8c;
  wire v3a6467a;
  wire v377b4ad;
  wire v374a6fc;
  wire v3734a79;
  wire v3a59d40;
  wire v3a5872a;
  wire v3a70cd5;
  wire v376b4d7;
  wire v3a6f958;
  wire v375de18;
  wire v3a66673;
  wire v3a5d822;
  wire v3757811;
  wire v3a5ca02;
  wire v2acaf23;
  wire v374056e;
  wire ce82b0;
  wire v375ee2a;
  wire v3a66464;
  wire v37624b2;
  wire v3a562a9;
  wire v375d453;
  wire v376969b;
  wire v360d03b;
  wire v3772c89;
  wire v377839d;
  wire v373f2d1;
  wire v377bc9c;
  wire v3a708a9;
  wire v3a70304;
  wire v3a7075b;
  wire v3a68b7b;
  wire v377b416;
  wire v3a6eec3;
  wire v3a64da2;
  wire v373c8db;
  wire v374b0eb;
  wire v3a5cff1;
  wire v3a70681;
  wire v3746cdd;
  wire v3742ffc;
  wire b0c091;
  wire v3735ac3;
  wire v377703d;
  wire v376d007;
  wire v377c3f5;
  wire v37523b5;
  wire v375edd8;
  wire v3a667ea;
  wire v376faf9;
  wire v37294f4;
  wire v374dddd;
  wire v3a6261f;
  wire v23fda46;
  wire v37603af;
  wire v3730383;
  wire v3a5cf0b;
  wire v3a70b47;
  wire v37295fe;
  wire v3757c6f;
  wire v39a5265;
  wire v3a6fc9f;
  wire v360d2c6;
  wire v375214d;
  wire v3a70b19;
  wire v37255a1;
  wire v376f14f;
  wire v3733138;
  wire v3a6eaee;
  wire v37356cc;
  wire v3a6f693;
  wire v3765af5;
  wire v3a70017;
  wire v375ae53;
  wire v3742ecd;
  wire v3a71327;
  wire v3a7140d;
  wire v377ea86;
  wire v2092b0b;
  wire v377e5e1;
  wire v3a5fdc8;
  wire v3808d2f;
  wire v37617d8;
  wire v3a703fc;
  wire v3a6a4e6;
  wire v377a104;
  wire v376d6b9;
  wire v3767902;
  wire v3734397;
  wire v3770891;
  wire v3729f3c;
  wire v3a5e3e2;
  wire v372bda4;
  wire v3759fda;
  wire v374e455;
  wire v3728ac4;
  wire v3730cb5;
  wire v3a70485;
  wire v372dc34;
  wire v3a2a128;
  wire v3a6ffe0;
  wire v376a35c;
  wire v3a715fd;
  wire v37464c8;
  wire v373f4d3;
  wire v2aca977;
  wire v3748529;
  wire v3771ce2;
  wire v374d037;
  wire v374502e;
  wire v3a6f453;
  wire v376de0b;
  wire v3a6446a;
  wire v373a7d4;
  wire v373bf7c;
  wire v372dd8e;
  wire v3a6cfa7;
  wire v37482f8;
  wire v3771b63;
  wire v3a5bb49;
  wire v376c592;
  wire v377f3af;
  wire v37794be;
  wire v37524c6;
  wire v3a71085;
  wire v2092b2f;
  wire v3777a7f;
  wire v3a6fe6a;
  wire v3745b52;
  wire v3a6efc9;
  wire v375f479;
  wire v3775da7;
  wire v3a703df;
  wire v377db8a;
  wire v3a7127f;
  wire v39eb1df;
  wire v373e41c;
  wire v3a6fa63;
  wire v3a5b0b3;
  wire v3a6ab5f;
  wire v377314f;
  wire v3a6f018;
  wire v37407cb;
  wire v3a66645;
  wire v373d223;
  wire v3744037;
  wire a81487;
  wire v3773092;
  wire v3a70b94;
  wire v3740f3d;
  wire v3723118;
  wire v375f030;
  wire v3a5db8a;
  wire v3772c51;
  wire v3a6fcba;
  wire v3745c45;
  wire c7885c;
  wire v3731cc6;
  wire v3726156;
  wire v3a6beff;
  wire v3a5bf56;
  wire v1e38224;
  wire v373ed70;
  wire v37583be;
  wire v3a6eb65;
  wire v374ca8a;
  wire v37682dd;
  wire v3a293c5;
  wire v3740690;
  wire v373ef4b;
  wire v376b4e1;
  wire v374908e;
  wire v3a5f1e8;
  wire v3a6f60c;
  wire v377beee;
  wire v374328c;
  wire v3748b2c;
  wire v372fade;
  wire v3a69c7b;
  wire v376ec1d;
  wire v2aca83b;
  wire v3734b6e;
  wire v373dfbe;
  wire v377b3a8;
  wire v3734e58;
  wire v3751e8d;
  wire v3758f64;
  wire v3775b4d;
  wire v3738877;
  wire v373dad7;
  wire v375640f;
  wire v372df2a;
  wire v37481e4;
  wire v3726609;
  wire v3a68591;
  wire v3a714ff;
  wire v3a6eb52;
  wire v3a6e305;
  wire v375fa71;
  wire v375884e;
  wire v3a705ec;
  wire v3a6f875;
  wire v3778ef8;
  wire v373c3bd;
  wire v39ebac7;
  wire v3a709c6;
  wire v3769cad;
  wire v3768180;
  wire v3a67851;
  wire v3779b03;
  wire v380662a;
  wire v375c196;
  wire v372e6ad;
  wire v3a5bbed;
  wire v377094b;
  wire v377122d;
  wire v3a71422;
  wire v3a708bd;
  wire v3a5f83e;
  wire v3778ac5;
  wire v37446b5;
  wire v3a7107a;
  wire v3a6f17f;
  wire v375c69e;
  wire v3a64ee3;
  wire v3a6eef6;
  wire v3a63abb;
  wire v3734625;
  wire v3734c05;
  wire v3a70131;
  wire v375ecc7;
  wire v375f462;
  wire v3747cf5;
  wire v3a6d30c;
  wire v3a70028;
  wire v23fda38;
  wire v376ef9f;
  wire v3a62c46;
  wire v3a6f1e2;
  wire v3766216;
  wire v3737dc7;
  wire v37349b9;
  wire v3740d4e;
  wire v3a6f45b;
  wire v3758eb3;
  wire d8fb57;
  wire v3725042;
  wire v3a6535f;
  wire v3756465;
  wire v3754aa3;
  wire v377ad9a;
  wire v375aaca;
  wire v3723b0c;
  wire v3a6f6a2;
  wire v37416ea;
  wire v325c960;
  wire v3745014;
  wire v3763668;
  wire v373ac52;
  wire v377167e;
  wire v376b088;
  wire v37422f3;
  wire v3756d28;
  wire v3a70fce;
  wire v375af00;
  wire v3757aa1;
  wire v3a70fbb;
  wire v377b576;
  wire v3a669c2;
  wire v374044c;
  wire v3760750;
  wire v3742e30;
  wire v3762034;
  wire v37291ce;
  wire v3a6f744;
  wire v3760bd6;
  wire v3a68c32;
  wire v3a6fa37;
  wire v37283ff;
  wire v3776f07;
  wire v3768429;
  wire v37579b8;
  wire v372c051;
  wire v3745d14;
  wire v375e217;
  wire v37787ce;
  wire v3a707cc;
  wire v3a662a2;
  wire v3a704eb;
  wire v37496c6;
  wire v3a58261;
  wire v376c208;
  wire v3733168;
  wire v375e5a6;
  wire v373250a;
  wire b3ccfa;
  wire v3a6fb4e;
  wire v372fd11;
  wire v3a5690f;
  wire v3a70385;
  wire v3736539;
  wire v37739ed;
  wire v3769ee7;
  wire v376822d;
  wire v372c79f;
  wire v3a614dd;
  wire v3a607c3;
  wire v377c6b0;
  wire v375f883;
  wire v37606bb;
  wire v37587a6;
  wire v375c6d6;
  wire v8455f7;
  wire v37330d6;
  wire v39a4f35;
  wire v377b311;
  wire v3a7094b;
  wire v3a6ebc6;
  wire v3a6fbc9;
  wire c76b50;
  wire v3778a82;
  wire v375b6fe;
  wire v372d86d;
  wire v3738a50;
  wire v3a672e6;
  wire v374ac6d;
  wire v3725a38;
  wire v37505cd;
  wire v3a6f7a9;
  wire v372c6c4;
  wire v3727d4c;
  wire v3a6f2a8;
  wire v3a53eeb;
  wire v3a6fce6;
  wire v377f09a;
  wire v3738dca;
  wire v3a5f50e;
  wire v3a674ac;
  wire v377dd3b;
  wire v3a57445;
  wire v37570b7;
  wire v3a70056;
  wire ad2d05;
  wire v37598c6;
  wire v35b70e6;
  wire v3a70a05;
  wire v375c845;
  wire v374b8fa;
  wire v3a70cb4;
  wire v377ce66;
  wire v3a58c79;
  wire v3a6f40c;
  wire v3722f12;
  wire v3767d7c;
  wire v3761be0;
  wire v377d67a;
  wire v374ea27;
  wire v374611e;
  wire v3a6f639;
  wire v372ed34;
  wire v3a59c65;
  wire v376afb3;
  wire v375ee68;
  wire v376f942;
  wire v3a5b51d;
  wire v3752a6c;
  wire v3757e71;
  wire v3a5aa64;
  wire v3767dc1;
  wire v373e806;
  wire v3a58980;
  wire d0b9d7;
  wire v377915c;
  wire v374da7f;
  wire v3771a0d;
  wire v3a6a0a6;
  wire v3a56d78;
  wire v377b92f;
  wire v373f785;
  wire v3739bcd;
  wire v3a6feee;
  wire v377972c;
  wire v3772183;
  wire v375ad91;
  wire v376e238;
  wire v3747f5d;
  wire v3a71513;
  wire v3a68dfd;
  wire v376cffc;
  wire v37c033d;
  wire v37361aa;
  wire v375b506;
  wire v3730646;
  wire v3a70cdd;
  wire v3a5b693;
  wire v372626a;
  wire v377a1dd;
  wire v37548b3;
  wire v373562f;
  wire ae13ec;
  wire v2acaf6f;
  wire c98f7c;
  wire v374d7dd;
  wire v3753940;
  wire v3742db5;
  wire v37528d5;
  wire v3776340;
  wire v3736c97;
  wire v3a56aae;
  wire v3772b00;
  wire v3a700fe;
  wire v3a6186a;
  wire v3a70822;
  wire v3a70c9a;
  wire v3759506;
  wire v3752684;
  wire v374f4d4;
  wire v373d79e;
  wire v377c2ba;
  wire v3752648;
  wire v3751c87;
  wire v373a07f;
  wire v37457d1;
  wire v3768428;
  wire v376d3f7;
  wire v3a7052a;
  wire v3a6bf86;
  wire v377baeb;
  wire v376fe88;
  wire v372c219;
  wire v3a5986c;
  wire v377f2a9;
  wire v3749d86;
  wire v3a663c3;
  wire v3a6816a;
  wire v372846c;
  wire v3740473;
  wire v3a552d4;
  wire v3a541ee;
  wire v936e47;
  wire v376a877;
  wire v37659f8;
  wire v37651b4;
  wire v375cdf8;
  wire v3a6fb5a;
  wire v372bef3;
  wire v3a70686;
  wire v3a64c6b;
  wire v3a70fcc;
  wire v3a6c5ed;
  wire v37689aa;
  wire v3770dbf;
  wire v374140e;
  wire v3a6738f;
  wire v375c7b9;
  wire v374e7f2;
  wire v374e409;
  wire v3752fbe;
  wire v376130f;
  wire v38074a8;
  wire v3a5edfe;
  wire v3a70b4c;
  wire v3763cf5;
  wire v37519ed;
  wire v3a635ff;
  wire v377ee58;
  wire v3a65f4c;
  wire v3a6b23f;
  wire v377762d;
  wire v1e37370;
  wire v3a6c933;
  wire v372fa17;
  wire v3772afb;
  wire v3a709f0;
  wire v372cbac;
  wire v3a6e9c0;
  wire v3a6356b;
  wire v3a29dbd;
  wire v3727db5;
  wire v3a60d5e;
  wire v3379070;
  wire v372df82;
  wire v3765722;
  wire v3735554;
  wire v3747585;
  wire v376dd15;
  wire v3a6f222;
  wire v3a70e23;
  wire v377022e;
  wire v37458a3;
  wire v375983d;
  wire v3a6b1d4;
  wire v3a66778;
  wire v374b10b;
  wire v37477d2;
  wire v373bb2d;
  wire v3760c90;
  wire v372f12d;
  wire v372c1a7;
  wire v3728739;
  wire v37265f2;
  wire v373a66b;
  wire v3a58a0d;
  wire v372cd50;
  wire v374d802;
  wire v3a58cb2;
  wire v3a6fa4b;
  wire v2619368;
  wire v8455d2;
  wire v8455ce;
  wire v8455c6;
  wire v8455c2;
  wire v8455ca;
  wire v8455ba;
  wire v8455be;
  wire v8455b6;
  wire v8455ff;
  wire v372fc17;
  wire v376f5fb;
  wire v377ac6f;
  wire v3774b25;
  wire v376e00a;
  wire v3739166;
  wire v37682c6;
  wire v3a7066e;
  wire v373e9a9;
  wire v376a006;
  wire v373fe74;
  wire v373d9aa;
  wire v3a55e7f;
  wire v3a5e0f7;
  wire a0d21b;
  wire v3771609;
  wire v3a6a8c0;
  wire v37447bf;
  wire v37749bf;
  wire v3a5b91d;
  wire v23fdaed;
  wire v374f609;
  wire v3a713e3;
  wire v3776e85;
  wire v3a70d32;
  wire v380919d;
  wire v3769740;
  wire v3729f7b;
  wire v376984f;
  wire v374ed4b;
  wire v3724710;
  wire v372b351;
  wire v3778765;
  wire v377ac7e;
  wire v375dc46;
  wire v37281e7;
  wire c511c2;
  wire v3a6106c;
  wire v3737075;
  wire v3a714be;
  wire v3a6ff08;
  wire be54b2;
  wire v3730a61;
  wire d0e017;
  wire v3775a9f;
  wire v3a66120;
  wire v3a6a7e8;
  wire v3769dcb;
  wire v3a5ce2f;
  wire v375d651;
  wire v377e928;
  wire v3744b38;
  wire v3a6f483;
  wire v3a66dcf;
  wire v3a70b6e;
  wire v3757c91;
  wire v3a632e8;
  wire v3739460;
  wire v375dcf5;
  wire v3a71644;
  wire v376dc58;
  wire v3a53dbf;
  wire v373301d;
  wire v3378f4c;
  wire v3730fb0;
  wire v37375e4;
  wire v3758c32;
  wire v373d737;
  wire v3a57046;
  wire v3a6d7f2;
  wire v3a6fe9a;
  wire v3731aac;
  wire v3a5c816;
  wire v3731b53;
  wire v3a70919;
  wire v3769fe3;
  wire v3a6982f;
  wire v3744999;
  wire v3a711b2;
  wire v3a55dc3;
  wire v3a565a8;
  wire v3735e84;
  wire v3724048;
  wire v3a61344;
  wire v3753001;
  wire v3a703b5;
  wire v375a397;
  wire be0e1a;
  wire v3755aae;
  wire v3724b78;
  wire v375c9a3;
  wire v3740174;
  wire v3a715c1;
  wire v3757100;
  wire v1e37af3;
  wire v3a5b9cd;
  wire v374f526;
  wire v37302fb;
  wire v37335a5;
  wire v3a6f6e1;
  wire v3a6a156;
  wire v375fea8;
  wire v38067ea;
  wire v37587a4;
  wire v3a71654;
  wire a65142;
  wire v3a66f8d;
  wire v3a64718;
  wire v3a68ebe;
  wire v3779d24;
  wire v373025a;
  wire v37401c2;
  wire v3769141;
  wire v360caba;
  wire v3a70122;
  wire v3a64103;
  wire v3776615;
  wire v372b7e5;
  wire v3769d3e;
  wire v375bc08;
  wire v376f7a0;
  wire v3a6fcf9;
  wire v3748d3b;
  wire v3a6f1b2;
  wire v375156a;
  wire v3729511;
  wire v3a71213;
  wire v372e443;
  wire v3a70794;
  wire v3a6f41c;
  wire v3726a2c;
  wire v3a55954;
  wire v3a5d5e7;
  wire v23fe379;
  wire v3728506;
  wire v376d4b7;
  wire v3a6fdf0;
  wire v3a62e01;
  wire v3a6a209;
  wire v3a655e9;
  wire v3750b8c;
  wire v3a6eb7a;
  wire v380755c;
  wire v373d449;
  wire v375a901;
  wire v3a70f03;
  wire v375865a;
  wire v3a2981e;
  wire v37451f8;
  wire v3a70b83;
  wire v372d6e5;
  wire v3a605bd;
  wire v3724002;
  wire v3a6eeff;
  wire v3a662fe;
  wire v37644e0;
  wire v3a71024;
  wire v3770161;
  wire v3757b16;
  wire v3a5c42c;
  wire v23fe217;
  wire v3750c08;
  wire v3a70e76;
  wire v3745614;
  wire v377d521;
  wire v3a554c5;
  wire v3a6f97f;
  wire v372e61a;
  wire v3a6f67e;
  wire v3758fc7;
  wire v3a67de4;
  wire v374d13c;
  wire v377fa89;
  wire v3737d48;
  wire v3a70722;
  wire v3a5fa81;
  wire v373e625;
  wire v3a6fda4;
  wire v3a6ff7c;
  wire v3725fe5;
  wire v3739c81;
  wire v3a700ad;
  wire v3765626;
  wire v37316fd;
  wire v374fa4d;
  wire v376051c;
  wire v37447e9;
  wire v375ec23;
  wire v377eada;
  wire v3730b67;
  wire v3751bdd;
  wire v3a6f98c;
  wire v3a68c19;
  wire v3a6887f;
  wire v3a6f962;
  wire v3a61d5f;
  wire v3a5bf99;
  wire v3a5bda1;
  wire v37578bd;
  wire v375cc11;
  wire v376269a;
  wire v3a6ef5a;
  wire v3747929;
  wire v374d8ea;
  wire v3a71677;
  wire v3a65260;
  wire v373becf;
  wire v37645da;
  wire v3a6b937;
  wire v3a6fefd;
  wire v374a20f;
  wire v374efb9;
  wire v3760091;
  wire bb41ad;
  wire v3a29844;
  wire v376aa3f;
  wire v3a711ee;
  wire v3a55162;
  wire v23fd9fe;
  wire v3a6ae54;
  wire v3739885;
  wire v374c058;
  wire v37317b4;
  wire v3a59fd0;
  wire a1bc5b;
  wire v3a69a9f;
  wire v376b89f;
  wire v3a705d2;
  wire v3777d70;
  wire v3a631f7;
  wire v3757bac;
  wire v3761019;
  wire v375242f;
  wire v3762c4c;
  wire v373ec80;
  wire v3a5ee7e;
  wire v3a6f820;
  wire v37730cd;
  wire v3763ca5;
  wire v3723df5;
  wire v3a6cd1b;
  wire v3a59918;
  wire v3727e15;
  wire v3724744;
  wire v3745509;
  wire v374c862;
  wire v3a63043;
  wire v3a54d59;
  wire v3741e12;
  wire v375104f;
  wire v3745dba;
  wire v374710b;
  wire v3a707f1;
  wire v374b918;
  wire v3a65dc4;
  wire v3755b94;
  wire v3a704d9;
  wire v3a70aa4;
  wire v37463ae;
  wire v3a6f75e;
  wire v374df50;
  wire v373ce86;
  wire v3723430;
  wire v3764834;
  wire v3739d4a;
  wire v3a71287;
  wire v3a70c11;
  wire v3767feb;
  wire v1e38239;
  wire v23fdc13;
  wire v373d434;
  wire v3737a30;
  wire v3a702ec;
  wire v3a6464f;
  wire v3732968;
  wire v3750edc;
  wire v3733e77;
  wire v3a58139;
  wire v3765590;
  wire v3a5bc72;
  wire v37245d9;
  wire v375463f;
  wire v3a6e138;
  wire v3a6f1ae;
  wire v9aea50;
  wire v3779ac2;
  wire v3a68d3f;
  wire v37252d0;
  wire v37654b9;
  wire v3a67ff8;
  wire v37289f0;
  wire v372721d;
  wire v3746877;
  wire v3a55aea;
  wire v3776018;
  wire v37370f1;
  wire v3a5457f;
  wire v3773390;
  wire v374262b;
  wire v377fb00;
  wire v3a6eb33;
  wire v3750d44;
  wire v3a54ba7;
  wire v376c248;
  wire v37494bb;
  wire v3774908;
  wire v3755199;
  wire v372864a;
  wire v3a6a2b5;
  wire v3a581e4;
  wire v3779fd9;
  wire v3a61cd7;
  wire v3a70ba9;
  wire v3a57721;
  wire v3a5f894;
  wire v3737456;
  wire v3738c45;
  wire v373f924;
  wire v376c630;
  wire v373c65b;
  wire v380947a;
  wire v376fca4;
  wire v3a68d0e;
  wire v3a6f617;
  wire v3a7152d;
  wire v375a367;
  wire v37579f1;
  wire v3a53d44;
  wire v3a71094;
  wire v3a691ca;
  wire v3a706ba;
  wire v3775e46;
  wire v37430fb;
  wire v3808865;
  wire b9f306;
  wire v3a70abb;
  wire v3746a87;
  wire v23fd9e7;
  wire v3a70247;
  wire v372ab70;
  wire v37654a9;
  wire v37466a5;
  wire v3a6d48a;
  wire v37445e2;
  wire v3a6fdf9;
  wire v374da33;
  wire v3a69091;
  wire v3777243;
  wire v3735e18;
  wire v374f2d1;
  wire v3a70fc0;
  wire v376b8e9;
  wire v3a29706;
  wire v377c7cf;
  wire v372edf9;
  wire v376db8a;
  wire v3729b37;
  wire v375b7fa;
  wire v3a69d13;
  wire v373ae0a;
  wire v374a1f5;
  wire v3753233;
  wire v374ce92;
  wire v3a5797b;
  wire v373fee1;
  wire v374fb51;
  wire v3a7065a;
  wire v372c06f;
  wire v3723ded;
  wire v3734d12;
  wire v377b4cc;
  wire v3a6fc5e;
  wire v372ba40;
  wire v3739589;
  wire v3752edc;
  wire v37260af;
  wire v3a6ae99;
  wire v3a6e7a7;
  wire v3a6fb84;
  wire v374ed51;
  wire v372869e;
  wire v375ebdd;
  wire v3766315;
  wire v376975e;
  wire v3767b66;
  wire v3a708ef;
  wire v3a65660;
  wire v37764ee;
  wire v9ccd8a;
  wire v374a7b2;
  wire v3762545;
  wire v3775b30;
  wire v373dc68;
  wire v3a6f9f5;
  wire v3a53c18;
  wire v3733bfc;
  wire v39eb565;
  wire v37724b9;
  wire v3740c13;
  wire v3756091;
  wire v377546d;
  wire v375d17d;
  wire v3a57f18;
  wire v375589b;
  wire v3a6fae2;
  wire v3750025;
  wire v3a6b4d7;
  wire v3a6e0f2;
  wire v3a6ffda;
  wire v3a5618d;
  wire v3a5bf28;
  wire v376605a;
  wire v3a6dcb2;
  wire v37749fd;
  wire v373e0ad;
  wire v92141c;
  wire v3a6b62d;
  wire v3a70a81;
  wire v372ba1c;
  wire v23fd7a9;
  wire v376d89f;
  wire v373a438;
  wire v3753f71;
  wire v380989b;
  wire v37788ca;
  wire v3a70888;
  wire v374005b;
  wire v3a6fdf4;
  wire v377d39f;
  wire v373d848;
  wire v3a64f97;
  wire v3774fa6;
  wire v3740625;
  wire v3a655cb;
  wire v3a6cacb;
  wire v375ef27;
  wire v3a701b3;
  wire v377b612;
  wire v3736439;
  wire v3a711c1;
  wire v376d566;
  wire v375a5b6;
  wire v3752c73;
  wire v373ff04;
  wire v3772904;
  wire v3a5d8bb;
  wire v3a6dd1a;
  wire v3a68289;
  wire v3a6f80b;
  wire v373aec3;
  wire v375e3a5;
  wire v375d34f;
  wire v3765d94;
  wire v3a68a46;
  wire v3768196;
  wire v3a6fef2;
  wire v3809d53;
  wire v373cfbd;
  wire v3a61038;
  wire v3732e48;
  wire v3a5c4b0;
  wire v3769a63;
  wire v374bf69;
  wire v3739774;
  wire v372bc0c;
  wire v372f6ec;
  wire v3740a1e;
  wire v8455b0;
  wire v377ed8c;
  wire v3a54bcd;
  wire bef73a;
  wire v37266e1;
  wire v3735fee;
  wire v3a6a867;
  wire v3a6fdd0;
  wire v37686c1;
  wire v375b4a7;
  wire v37627f9;
  wire v373c423;
  wire v3a636fe;
  wire v372ab5a;
  wire v3755e82;
  wire v374e606;
  wire v37257c8;
  wire v3a698c3;
  wire v3a6eb76;
  wire v3746f46;
  wire v376e772;
  wire v3a623ca;
  wire v3a5ddc1;
  wire v3809439;
  wire v9c0027;
  wire v375237c;
  wire v3a590d1;
  wire v3a57fa3;
  wire v3a6fe81;
  wire v3a6fc93;
  wire v3a55cf3;
  wire v37409cd;
  wire v3a708f4;
  wire b3b89e;
  wire v3749535;
  wire v375d512;
  wire v3a5a25a;
  wire v3766809;
  wire v3a62dec;
  wire v372b69c;
  wire v3a7123c;
  wire v3a570c0;
  wire v3749d1d;
  wire v8455fd;
  wire v3749a12;
  wire v376f56d;
  wire v3738b8a;
  wire v374a11d;
  wire v372b164;
  wire v3a70cf1;
  wire v37233e4;
  wire v3777647;
  wire v3a6604e;
  wire v3a715ba;
  wire v3a6ff4b;
  wire v375725f;
  wire v3759c96;
  wire v3a6fd84;
  wire v37412e9;
  wire v3763a12;
  wire v3a6ebf7;
  wire v37682ce;
  wire v373e12b;
  wire v37514f7;
  wire v3a6f9fa;
  wire v3733b9a;
  wire v3a5dbd7;
  wire v360d10b;
  wire v3779fd2;
  wire v3a5ed31;
  wire v37384a9;
  wire v3a5b955;
  wire v3a71118;
  wire v3577324;
  wire v3a70924;
  wire v3a566c1;
  wire v325c957;
  wire v3768e52;
  wire v3a706bd;
  wire v373927b;
  wire v373049b;
  wire v373adea;
  wire v3a560d9;
  wire v3a61e95;
  wire v3a7122f;
  wire v372661f;
  wire v3a635b9;
  wire v376ff3d;
  wire a6c8aa;
  wire v3a626d4;
  wire v375766c;
  wire v377195f;
  wire v374845f;
  wire v372b8a3;
  wire ce8abd;
  wire v3a713f6;
  wire v3757194;
  wire v3763562;
  wire v3a70df5;
  wire v3a7031e;
  wire v374a4c2;
  wire v3763c1f;
  wire v37725ea;
  wire v3a702ee;
  wire v3806f0b;
  wire v3a606b0;
  wire v377b0b0;
  wire v3a6f8c7;
  wire v3779c5d;
  wire v3a67cf0;
  wire v3a68c26;
  wire v37477cb;
  wire v373e4a7;
  wire v375b5d6;
  wire v37351ff;
  wire v37490d7;
  wire v3a67fb5;
  wire v3a6f31f;
  wire v3770b6c;
  wire v8455b2;
  wire v3776b20;
  wire v3760bc2;
  wire v3a64862;
  wire v377559f;
  wire v3764fd7;
  wire v3743677;
  wire v377a468;
  wire v376b1ee;
  wire v376a2e7;
  wire v3a54c8d;
  wire v3775653;
  wire v373df7f;
  wire v3739ab4;
  wire v3779595;
  wire v3a65612;
  wire v3746a67;
  wire v3743017;
  wire v3768274;
  wire v3764d82;
  wire v374aa27;
  wire v3a6836a;
  wire v3757bf1;
  wire v3a70be1;
  wire v376f583;
  wire v3729113;
  wire v38099c8;
  wire v3773650;
  wire v3a65b4a;
  wire v3774db3;
  wire v9e52e0;
  wire v375ed5c;
  wire v3761e97;
  wire v3a620f2;
  wire v3a6402e;
  wire v372a20d;
  wire v376769a;
  wire v373c3ac;
  wire v3a6dbec;
  wire v37c36b9;
  wire v3728a4a;
  wire v3a6844c;
  wire v3a5aa8e;
  wire v373de47;
  wire v377073b;
  wire v3a6f234;
  wire v373e1cc;
  wire v3a5bc0a;
  wire v37532f0;
  wire v3a6fb8f;
  wire v375095e;
  wire v3a71675;
  wire v3a6ff8c;
  wire v376256f;
  wire v377265b;
  wire v2093252;
  wire v3a70aa6;
  wire v3765a2e;
  wire v3723134;
  wire v3a70e0e;
  wire v376f71a;
  wire v3729792;
  wire v3a6f916;
  wire v3a6bb56;
  wire v35b708c;
  wire v3a6a918;
  wire v373553c;
  wire v3a6deec;
  wire v23fda2f;
  wire v3a70df9;
  wire v377fbb9;
  wire v373b58a;
  wire v3a6ff41;
  wire v3755a9f;
  wire v3a66651;
  wire v375646d;
  wire v3a5524f;
  wire v3a541ec;
  wire v3a71338;
  wire v3765e47;
  wire v3732632;
  wire v3a6c892;
  wire v373833b;
  wire v37342cd;
  wire v3a707e5;
  wire v3a6f118;
  wire v3753a28;
  wire v3a703dd;
  wire v3725bdc;
  wire v3a70f44;
  wire v3763dd4;
  wire v3a2a105;
  wire v3756780;
  wire v37744e0;
  wire v377b3ff;
  wire v3a70eea;
  wire v3774859;
  wire v3a6f154;
  wire v3a71039;
  wire v3a6f394;
  wire v3a65100;
  wire v373765a;
  wire v8d9a96;
  wire v3767f58;
  wire v376025f;
  wire v376665a;
  wire v374abee;
  wire v3a674fa;
  wire v3770fdb;
  wire v3a6f4dd;
  wire v3756219;
  wire v3a70b4b;
  wire v374221c;
  wire cd5e35;
  wire v3725be9;
  wire v3a690a6;
  wire v37510d9;
  wire v375ed69;
  wire v373dce8;
  wire v3a67133;
  wire v3728826;
  wire v377f200;
  wire v3a6ef62;
  wire v37697fc;
  wire v374cbe3;
  wire baec07;
  wire v3a5c3d6;
  wire v3774730;
  wire v3766309;
  wire v35b91b9;
  wire v377cd68;
  wire v3a706e1;
  wire v3a70b3b;
  wire v39ebb8a;
  wire v372ad2c;
  wire v375610e;
  wire v3a6f8cf;
  wire v376e587;
  wire v3757765;
  wire v374f0f5;
  wire v3a6de93;
  wire v3a6b931;
  wire v3a70e9e;
  wire v3a5865e;
  wire v3742f25;
  wire v23fdbe3;
  wire v374e51a;
  wire v3a5b8a2;
  wire v3a67095;
  wire v3742a61;
  wire v3a6cc2a;
  wire v37372a1;
  wire v37286f3;
  wire v37612a3;
  wire v3740c94;
  wire v3752f9b;
  wire v3a6fe27;
  wire d390f8;
  wire v3760314;
  wire v2acb110;
  wire dc5778;
  wire v375c6c1;
  wire v376a7da;
  wire v372b61a;
  wire v3723698;
  wire v372a732;
  wire v3748c34;
  wire v374c6b1;
  wire v3729022;
  wire v375af98;
  wire v377b429;
  wire v373016b;
  wire v37540d9;
  wire v3a61094;
  wire v376c505;
  wire v3a6fd9c;
  wire v3778b48;
  wire v3a6f435;
  wire v3a6f518;
  wire c63c1f;
  wire v37482c3;
  wire v3a6fb77;
  wire v3a6a68c;
  wire v3730ae6;
  wire v3750735;
  wire v372eb5b;
  wire v375d113;
  wire v3731800;
  wire v37345a4;
  wire v375ce2d;
  wire c8e1cc;
  wire v375bce2;
  wire v3776fec;
  wire v3768aaa;
  wire v376915a;
  wire v3a714c3;
  wire v377568c;
  wire v375968a;
  wire v375dab2;
  wire v3a5f41b;
  wire v3a6f6bc;
  wire v37354da;
  wire v376efcc;
  wire v3765d2b;
  wire v3745cf8;
  wire v372a2ae;
  wire v3a71372;
  wire v373f4dd;
  wire v372d071;
  wire v3a5646d;
  wire v375089b;
  wire v374113f;
  wire v376a74a;
  wire v2acafdd;
  wire v3a7154d;
  wire v3727171;
  wire v377e962;
  wire v3a70291;
  wire v374cca4;
  wire a61746;
  wire v3a656bd;
  wire v3a622a9;
  wire v37766b2;
  wire v3a5e660;
  wire v3a5f592;
  wire v375076f;
  wire v3a70f2c;
  wire v372ad83;
  wire v3747c9f;
  wire v3739246;
  wire v373ab2b;
  wire v3739cdb;
  wire v35772dd;
  wire v3731fe4;
  wire cea42b;
  wire v373fa33;
  wire v3a70c18;
  wire b1fcb7;
  wire v3723459;
  wire v3a6ffd8;
  wire v3a6ff55;
  wire v3a7058c;
  wire v3a6ef55;
  wire v376e860;
  wire v3a6df62;
  wire v375961b;
  wire v3772d8b;
  wire v3743fee;
  wire v376fb6e;
  wire v376c88f;
  wire v374e06d;
  wire v374158f;
  wire v372d685;
  wire a04f67;
  wire v37fca9f;
  wire v3773343;
  wire v3a66039;
  wire v374c9ab;
  wire v377233c;
  wire v3729360;
  wire v3a607fa;
  wire v3a5f6c3;
  wire v3a6da41;
  wire v373875c;
  wire v3751c12;
  wire v377d8f9;
  wire v3732f31;
  wire v3a703cf;
  wire v377c2e6;
  wire v37562fd;
  wire v3a580a0;
  wire v372e34d;
  wire v372361c;
  wire v3752a7e;
  wire v3a70e9f;
  wire v374b690;
  wire v376bf0a;
  wire v38072f9;
  wire v3a67577;
  wire v3745abb;
  wire v374e033;
  wire v3762ba2;
  wire v3a59746;
  wire v3770f48;
  wire v373ec60;
  wire v3a6f345;
  wire v377faff;
  wire v3a6a56e;
  wire v3a58c07;
  wire v3a6ca54;
  wire v3807074;
  wire v3747454;
  wire v375e6ff;
  wire v3a70a01;
  wire v374ff84;
  wire v3a59314;
  wire v3764678;
  wire v3a7118e;
  wire v374edb8;
  wire v1e378da;
  wire v375c697;
  wire v3a5585e;
  wire v3723ba5;
  wire v373a1b4;
  wire v3a70a42;
  wire v3777763;
  wire v3747b74;
  wire v372cae4;
  wire v373fa04;
  wire v372535d;
  wire v375e074;
  wire v3a5f626;
  wire v3762bdf;
  wire v3734dc5;
  wire v3a60ef2;
  wire v3a60132;
  wire v37765fe;
  wire b4444b;
  wire v3774913;
  wire v37722c6;
  wire v3a6fd15;
  wire v376a65a;
  wire v3a61397;
  wire v37377c8;
  wire v3773b0f;
  wire v3724c46;
  wire v376625e;
  wire v3a6416b;
  wire v3a71036;
  wire v375acae;
  wire v37391e5;
  wire v3a67251;
  wire v3a5d5d3;
  wire v376b307;
  wire v3a6a187;
  wire v377ec9b;
  wire v3a7057b;
  wire v3760d83;
  wire v37533ac;
  wire a29a96;
  wire v377395b;
  wire v3a6b1e4;
  wire v374b8e2;
  wire b12fe4;
  wire v376bd43;
  wire v37270a2;
  wire v3739e36;
  wire v3731499;
  wire v376587d;
  wire v375cc17;
  wire v376ab29;
  wire ad41f9;
  wire v38074aa;
  wire v3a6f144;
  wire v3776311;
  wire v3760317;
  wire v3a570a0;
  wire v37788d7;
  wire v372a0e6;
  wire v373f909;
  wire v3a6ebd8;
  wire v3a70430;
  wire v373f13e;
  wire v372e0b7;
  wire v376e66e;
  wire v3740247;
  wire v3722f50;
  wire v37479ee;
  wire v374f048;
  wire v37366df;
  wire v1e37af7;
  wire v372a2e4;
  wire v3732853;
  wire v376cab5;
  wire v373d8e4;
  wire v3a56aee;
  wire v3a6e0bf;
  wire v3a709f7;
  wire v3772c08;
  wire v3a64ef2;
  wire v3a6f8b2;
  wire v377596e;
  wire v376aa62;
  wire v373ec96;
  wire v3a70b40;
  wire v373c433;
  wire v3723a2c;
  wire b85e8b;
  wire v3a708a2;
  wire a0503f;
  wire v375178f;
  wire v3a65b5d;
  wire v3a6c2df;
  wire v23fe361;
  wire v3730930;
  wire v3a70381;
  wire v374c2e2;
  wire v3a6a9d3;
  wire v377f5db;
  wire v373385b;
  wire v3a6faaa;
  wire v37776c8;
  wire v3a5ca22;
  wire v3a6a42a;
  wire v3728434;
  wire v37367ba;
  wire v3743172;
  wire v3755791;
  wire v375b737;
  wire v3a63057;
  wire v37241fd;
  wire v33790da;
  wire v373291c;
  wire v3757b32;
  wire v3734aef;
  wire v3a5e696;
  wire v373c1a0;
  wire v373519d;
  wire v3a63717;
  wire v37479c3;
  wire v37607af;
  wire v3756813;
  wire v37257cf;
  wire v372b396;
  wire v3751bf3;
  wire v37356d4;
  wire v377a110;
  wire v3a5d7bf;
  wire v376eeac;
  wire v3a6eec2;
  wire v3a65384;
  wire v3760fb0;
  wire v37666f6;
  wire v373f1db;
  wire v3770653;
  wire v3754a0d;
  wire v3736d3a;
  wire v3a6d531;
  wire v375aff8;
  wire v3a70b13;
  wire v3735f30;
  wire v3733e04;
  wire v37410b9;
  wire v37296ca;
  wire v37598e6;
  wire v3a593e0;
  wire v377c17f;
  wire dc6ea3;
  wire v375e5d4;
  wire v3a56dd5;
  wire v38090f4;
  wire v3a5e2a3;
  wire v3742938;
  wire v3756981;
  wire v3752759;
  wire v37679b0;
  wire v3a62f75;
  wire v373d3e5;
  wire v374143e;
  wire v3a6051e;
  wire v3806db2;
  wire v3744f37;
  wire v372e351;
  wire v3a56f2e;
  wire v3a6f233;
  wire v3a6fbb8;
  wire v377b32c;
  wire v3a58546;
  wire v375a94d;
  wire v23fdb05;
  wire v377852a;
  wire v373a4e4;
  wire v3a707ad;
  wire v3a70fb2;
  wire v376d7a5;
  wire v3736b19;
  wire v3a69fe5;
  wire v3a61a3d;
  wire v3a70d99;
  wire v375b445;
  wire v3a705c5;
  wire v3775cb7;
  wire v3762e16;
  wire v37613b3;
  wire v3a6fe92;
  wire v3745158;
  wire v37386f5;
  wire v3a6fbef;
  wire v376641b;
  wire v375f87b;
  wire v37440af;
  wire v374891f;
  wire v8455b9;
  wire v374212c;
  wire v376728e;
  wire v373ea7f;
  wire v3757301;
  wire v37316f3;
  wire v3a701af;
  wire v3735f31;
  wire v3a6f83f;
  wire v373e689;
  wire v376e89b;
  wire v37626d4;
  wire v3768685;
  wire v3766c5c;
  wire v3a71344;
  wire v376b88d;
  wire v3753a06;
  wire v372acd0;
  wire v3762eeb;
  wire v3777412;
  wire v3752e63;
  wire v37428b3;
  wire v375c8e6;
  wire v3a62bce;
  wire v376e25b;
  wire v375f014;
  wire v3a5f711;
  wire v374b116;
  wire v3737ce3;
  wire v37698c3;
  wire v3774eec;
  wire v3728cdc;
  wire v3777c0c;
  wire v3756a20;
  wire v376198e;
  wire v37349cc;
  wire v375ff00;
  wire v3a664e6;
  wire v375dd4c;
  wire v377073f;
  wire v3a6eb2a;
  wire v3a71416;
  wire v3755d64;
  wire v3775bd3;
  wire v3739517;
  wire v372cedb;
  wire v3a6bc65;
  wire v3a7015f;
  wire v3741bce;
  wire v374e4c5;
  wire v3a55e8e;
  wire v3a71453;
  wire v3a6c6ec;
  wire v3737d02;
  wire v3a6ca24;
  wire v374e64f;
  wire v372fba0;
  wire v3770c99;
  wire v372cdd7;
  wire v377300f;
  wire v3779613;
  wire v374dc99;
  wire v37382eb;
  wire v3a6f5d4;
  wire v376cef0;
  wire v3a70cf5;
  wire v374fbb6;
  wire v3751d33;
  wire v374cd15;
  wire v3a70bf9;
  wire v3a6c15d;
  wire v376778a;
  wire v377a5d4;
  wire v3741890;
  wire v3776413;
  wire v37452a4;
  wire v38070c7;
  wire v374c2d6;
  wire v3727651;
  wire v3730878;
  wire v377c0ad;
  wire v3731555;
  wire v3a70df8;
  wire v3729c28;
  wire v377da14;
  wire v376f182;
  wire v3a713d2;
  wire v3a6f622;
  wire v3a71299;
  wire v3a580ca;
  wire v3a5e245;
  wire v3a714ed;
  wire v3a62eaa;
  wire v3a6f863;
  wire v3a59613;
  wire v372f4ea;
  wire v3a71203;
  wire v3a7032b;
  wire v37295e7;
  wire v3746406;
  wire v3755a27;
  wire v377209d;
  wire v377b0f8;
  wire v3a6f3ae;
  wire v3774b71;
  wire v37719a1;
  wire v23fdac1;
  wire v3a5fb90;
  wire v3764378;
  wire v3759628;
  wire v3760e13;
  wire v377f0dc;
  wire v3a6f046;
  wire v37395bc;
  wire v3777ce4;
  wire v3a70f68;
  wire v3a635c3;
  wire v372c84a;
  wire v3770b26;
  wire v3a70baf;
  wire v377cd7f;
  wire v3758472;
  wire v3737acd;
  wire v3a6eff7;
  wire v376871e;
  wire v37355d8;
  wire v377f734;
  wire v374e663;
  wire v375aeb3;
  wire v373dbbb;
  wire v373827a;
  wire v373869b;
  wire v373195f;
  wire v3a7067d;
  wire v375b626;
  wire v3774647;
  wire v3a6d31d;
  wire v3a680cb;
  wire v3a6ef96;
  wire v376dd8b;
  wire v376f01b;
  wire v3807071;
  wire v3753f1a;
  wire v3a703ac;
  wire v3a5d28b;
  wire v374b72f;
  wire v3a6f87f;
  wire v2ff9291;
  wire v3765511;
  wire v37565b0;
  wire v372b9c5;
  wire v3a6f804;
  wire v372874c;
  wire v3745b02;
  wire v377bfc7;
  wire v375a4d0;
  wire v3a56069;
  wire v37312e3;
  wire v3a5b45b;
  wire v375c70a;
  wire v3771088;
  wire v3a6f76d;
  wire v3758fa7;
  wire v374569b;
  wire v373d53f;
  wire v3777955;
  wire bae881;
  wire v3751491;
  wire v376d0ff;
  wire v3a6f0d5;
  wire v35b7169;
  wire v3731826;
  wire v377246f;
  wire v3a68871;
  wire v3a6fc97;
  wire v3772b42;
  wire v37515a6;
  wire a39369;
  wire v3756e20;
  wire v3723ec6;
  wire v3a5f000;
  wire v3a6ec0b;
  wire v3a6eb40;
  wire v1e38301;
  wire v377463a;
  wire v373b779;
  wire v3724596;
  wire v37332fa;
  wire v3a6f2d2;
  wire v3a6765d;
  wire v376b6d8;
  wire ca11a2;
  wire v373dff6;
  wire v3a5e19b;
  wire v372ff75;
  wire v373d746;
  wire v377a893;
  wire v3a70471;
  wire v3727b7f;
  wire v3730389;
  wire v3761f78;
  wire v373e5c8;
  wire v3a71015;
  wire v372fe3c;
  wire v374d9b7;
  wire v372349f;
  wire v3759837;
  wire v3740348;
  wire v376d2b7;
  wire v375a8cf;
  wire v3760658;
  wire v376a040;
  wire v373d2e0;
  wire v37314db;
  wire v3a70b53;
  wire v373cb9c;
  wire v3a6b059;
  wire v3a5e0cc;
  wire v3a5815e;
  wire v3a6affa;
  wire v3a58588;
  wire v372295a;
  wire v3a70a2e;
  wire v3a713b2;
  wire v3a6ef8c;
  wire v3a6f252;
  wire v3748bb1;
  wire v376eb2b;
  wire v3767399;
  wire v3777e08;
  wire v373adae;
  wire v37637d6;
  wire v376c63d;
  wire v3742cde;
  wire v3725786;
  wire v3a6f616;
  wire v3777baa;
  wire v375cade;
  wire v374a70f;
  wire v3a5eaa1;
  wire v375135a;
  wire v3735293;
  wire v377d377;
  wire v3a6b924;
  wire v3752707;
  wire v377d8b3;
  wire v3a592be;
  wire v37456a9;
  wire v373c728;
  wire v3a70283;
  wire v3a6fd71;
  wire v3768c21;
  wire v377e2f1;
  wire v37376c8;
  wire v3759b9a;
  wire v37273c2;
  wire v37403e5;
  wire v3a70394;
  wire v37485ec;
  wire v3a5a0e2;
  wire v37675e2;
  wire v377109d;
  wire v375d774;
  wire v3a70974;
  wire v377c3ea;
  wire v3a67519;
  wire v3763d52;
  wire v3a69444;
  wire v373d107;
  wire v3743e4f;
  wire v3a6f389;
  wire v375dea9;
  wire v3775393;
  wire c7658c;
  wire v3a715ea;
  wire v3731c27;
  wire v377a606;
  wire v3a5dde0;
  wire v3a6f35c;
  wire v3a70cd1;
  wire v3a65562;
  wire v2acaf72;
  wire v360c6f5;
  wire v3a63b56;
  wire v3759c9c;
  wire v377c3fb;
  wire v3a6eb01;
  wire v375d161;
  wire v375ac70;
  wire v3768d79;
  wire c6598e;
  wire v374b5da;
  wire v375c806;
  wire v3a63ff3;
  wire v374610e;
  wire v3a6f0b2;
  wire v375f326;
  wire v3763868;
  wire v3a5f26f;
  wire v3735d9c;
  wire v3a675ad;
  wire v37419df;
  wire v3a6f706;
  wire v37c0282;
  wire v3a70257;
  wire v3744dc6;
  wire v3744aed;
  wire v3a70c02;
  wire v373e7c0;
  wire v375fed9;
  wire v376afc5;
  wire v3761d0c;
  wire v375b7b0;
  wire v3731ca8;
  wire v3a6fe06;
  wire v3761b75;
  wire v373de8a;
  wire v3a6fe8e;
  wire v373b012;
  wire v37649a0;
  wire v375ebe9;
  wire v3764870;
  wire v3a70b80;
  wire v3740d4a;
  wire v377405e;
  wire v3a6fab4;
  wire v3724345;
  wire v3a66c14;
  wire v3a58541;
  wire v3779c40;
  wire v375be25;
  wire v376374b;
  wire v37507d0;
  wire v372eada;
  wire v374978c;
  wire v3a69fbe;
  wire v3751aaa;
  wire v3a7167e;
  wire v3a58b20;
  wire v3a7060a;
  wire v3a60974;
  wire v3a6a093;
  wire v374445b;
  wire v3745cc6;
  wire v3748460;
  wire v3738ca1;
  wire v375e320;
  wire v3a6ef63;
  wire v3a70d92;
  wire v3a5f4ef;
  wire v373e845;
  wire v3a6f448;
  wire v374875f;
  wire v3a59819;
  wire v376702a;
  wire v3754c51;
  wire v3774628;
  wire v3a58615;
  wire v376ca9f;
  wire v3a637a1;
  wire v375f44a;
  wire v3a70144;
  wire v3a7072e;
  wire v373330a;
  wire v3a6c515;
  wire v372f3e0;
  wire v3a707f6;
  wire v377671e;
  wire v377e13b;
  wire v372e92b;
  wire v3a6eab3;
  wire v3732588;
  wire v3a6d219;
  wire v37474c2;
  wire v3757ecc;
  wire v377320c;
  wire v3a7119e;
  wire v3772443;
  wire v3a5cf3d;
  wire v3a62a71;
  wire v3a70062;
  wire b4ac83;
  wire v3778afd;
  wire v376f0ab;
  wire v3777a9a;
  wire v3a6fcf3;
  wire v1e37996;
  wire v372a2f5;
  wire v3a6fb1f;
  wire v3a6f61e;
  wire v372b795;
  wire v3807a8d;
  wire v373228a;
  wire v373e858;
  wire v3a6a1b4;
  wire v3770abd;
  wire v3764015;
  wire v3a700ee;
  wire v35b6a6b;
  wire v375eb56;
  wire v3a702c1;
  wire v375a0a1;
  wire v3a62443;
  wire v374530a;
  wire v37513d1;
  wire v3a5deb7;
  wire v3a71109;
  wire v1e3731f;
  wire v2aca784;
  wire v3a58520;
  wire v3756bb9;
  wire v37312e2;
  wire v374fd45;
  wire v372f1a0;
  wire v3a6f618;
  wire v376fe30;
  wire v3a689eb;
  wire v3a6fc63;
  wire v3a6d364;
  wire v373502e;
  wire v372bfd3;
  wire v375cd4c;
  wire v3a54b63;
  wire v374df63;
  wire v3768076;
  wire v374c0e3;
  wire v376428f;
  wire v3734f7b;
  wire v372ea51;
  wire v3a7120c;
  wire v373fc07;
  wire v3771697;
  wire v3a6867e;
  wire v3a6c6cf;
  wire v37517d2;
  wire v3756a09;
  wire v3755a10;
  wire v3a6fd17;
  wire v3748f48;
  wire v337901e;
  wire v376064b;
  wire v372599c;
  wire v3a58e7f;
  wire v375e6b3;
  wire v3a6c243;
  wire v3a565eb;
  wire v3a63329;
  wire v3a7030f;
  wire v3747178;
  wire v3a66381;
  wire v3a56ca1;
  wire v372f997;
  wire v3a6cc93;
  wire v3722dfe;
  wire v3750ae0;
  wire v3734081;
  wire v3737ba0;
  wire v376d892;
  wire v3a58016;
  wire v3744d2a;
  wire v3725a2e;
  wire v3a70746;
  wire v3a6119e;
  wire v373aaed;
  wire v3a6f96b;
  wire v3a71239;
  wire v3808f3c;
  wire v3761eb6;
  wire v3761d5a;
  wire v3a6fadb;
  wire v3a6f81d;
  wire v1e382a5;
  wire v3726c8d;
  wire v373cf96;
  wire v376f1c0;
  wire v37462e7;
  wire v3a659d0;
  wire v3a544db;
  wire v3a7054a;
  wire v3770ab9;
  wire v37488fe;
  wire v374b05b;
  wire v3725bfb;
  wire v37696fe;
  wire v3a70ad3;
  wire v3a64089;
  wire v3723021;
  wire v3a5d5cc;
  wire v3a6bbeb;
  wire v3741b6c;
  wire v376f345;
  wire v3a6dddb;
  wire v37477ca;
  wire v3808f44;
  wire v3730eae;
  wire v3749ff9;
  wire v374a4d2;
  wire dac328;
  wire v372ec6d;
  wire v3737084;
  wire v3a702f7;
  wire v3754922;
  wire v3732759;
  wire v3728621;
  wire v3a5c6d8;
  wire v3774ee5;
  wire v3a6a680;
  wire v373384b;
  wire v3a69e22;
  wire v375f989;
  wire v9e78af;
  wire v3a6da59;
  wire v380702c;
  wire ac6831;
  wire v3a6f063;
  wire v3755db9;
  wire v3a70dc3;
  wire v374494b;
  wire v3739fc8;
  wire v376be82;
  wire v37485e2;
  wire v37726bf;
  wire v3725a65;
  wire v3752aa3;
  wire v374bba3;
  wire v37470de;
  wire v3763832;
  wire v375259d;
  wire v374d5fa;
  wire v3779d06;
  wire v3756c22;
  wire v37585c9;
  wire v3a582ea;
  wire v3730a7b;
  wire v373287a;
  wire b0ac65;
  wire v373803a;
  wire v37461d8;
  wire v3a6efb1;
  wire v373f0c7;
  wire v3733ac0;
  wire v37466c1;
  wire v3a70f11;
  wire v37536bf;
  wire v3a6aa9e;
  wire v3a6fa6f;
  wire v3a5c6e9;
  wire v372ab8f;
  wire v3a620f1;
  wire v376abd9;
  wire v3743e90;
  wire v3a5a9b3;
  wire v37418f3;
  wire v3733c70;
  wire v3754e8e;
  wire v3731312;
  wire v3775806;
  wire v3740811;
  wire v37390ec;
  wire v376daac;
  wire v3a6a3e5;
  wire v3a585fd;
  wire v372fd5d;
  wire v3763e55;
  wire v3a6d1ea;
  wire v3753592;
  wire v894fb9;
  wire v3a7148c;
  wire v3756524;
  wire v376ea99;
  wire v3a71555;
  wire v3a6fdbd;
  wire v1e373f8;
  wire v374ba57;
  wire v3808eb7;
  wire v3a6fcd8;
  wire v374071d;
  wire v373d0eb;
  wire v37674f2;
  wire v3a7046a;
  wire v372bb4b;
  wire v376f0c3;
  wire v3768ac7;
  wire v3a64f4f;
  wire v37309cf;
  wire v3779b95;
  wire v377f118;
  wire v377c4b8;
  wire v3a6f8e6;
  wire v376ee20;
  wire v37730d2;
  wire v3741a07;
  wire d4044f;
  wire v372c470;
  wire v3731508;
  wire v37546a9;
  wire v376d7d5;
  wire v37304a0;
  wire v377371c;
  wire v3a71523;
  wire v373dff9;
  wire v373d6dd;
  wire v3757188;
  wire v373e674;
  wire v37366eb;
  wire v3747630;
  wire v375c1fd;
  wire v3759b61;
  wire v372ce4b;
  wire v3a6f274;
  wire v372c30a;
  wire v3725eb6;
  wire v373cdef;
  wire v3a5bc70;
  wire v3a577ed;
  wire v3749a98;
  wire v3a70762;
  wire v3776225;
  wire v2acb5a2;
  wire v3a70526;
  wire v3a71652;
  wire v3755cb2;
  wire v209325d;
  wire v376e5b6;
  wire v8c34b7;
  wire v3a6ffe1;
  wire v3a5b404;
  wire v3808d7d;
  wire v372be5d;
  wire v3745249;
  wire v3a66af8;
  wire v3a58519;
  wire v372dc8e;
  wire v3a56aa0;
  wire v372dbb0;
  wire v3a5aa42;
  wire v372cf62;
  wire v373fecd;
  wire v377d219;
  wire v3760d59;
  wire v3a70e3a;
  wire v376a967;
  wire v372fe05;
  wire v376e491;
  wire v3a2a766;
  wire v376acf0;
  wire v377903c;
  wire v376111d;
  wire v377018e;
  wire v372455c;
  wire v3a2ae01;
  wire v3a70e2e;
  wire v3a5d763;
  wire v373a9ef;
  wire v3762452;
  wire v3739443;
  wire v3a7104b;
  wire v376d256;
  wire v3a55033;
  wire v37273b0;
  wire v3724f1d;
  wire v3779075;
  wire v3a70fad;
  wire v373c830;
  wire v374282f;
  wire v374249a;
  wire v3722eee;
  wire v3a6d401;
  wire v3a70e33;
  wire v376fcc3;
  wire v3a59ed6;
  wire v376f9a1;
  wire v375aa07;
  wire v376d9ed;
  wire v3771b2a;
  wire v377d9ab;
  wire v39a535f;
  wire b4f302;
  wire v3748f87;
  wire v3a6419e;
  wire v3762cb2;
  wire v3759cc1;
  wire v3a6eb7f;
  wire v37390ff;
  wire v3a705ac;
  wire v376d79d;
  wire v372a0b0;
  wire v3a58a34;
  wire v3a56582;
  wire v3a6f897;
  wire v3755e23;
  wire v376bae4;
  wire v373ce2b;
  wire v3764d1f;
  wire v3735b3e;
  wire v3a58e93;
  wire v373aef5;
  wire v3a6f2b6;
  wire v3a708c6;
  wire v3772326;
  wire v37311a4;
  wire v37234f5;
  wire cd348d;
  wire v3a61279;
  wire v3a60a32;
  wire v3771e23;
  wire v3779aa8;
  wire v3a60cd0;
  wire v3a5398c;
  wire v37337f1;
  wire v3a57d1f;
  wire v3a713a3;
  wire v37354c1;
  wire v39eb44a;
  wire v372e6d3;
  wire v37702c5;
  wire v3725a39;
  wire v3a6046c;
  wire v325b5ea;
  wire v374ccb7;
  wire v3754202;
  wire v3a6f22c;
  wire v377c9b1;
  wire v3a7119d;
  wire v3a67fd0;
  wire v3774314;
  wire v3747a0d;
  wire v93ca8c;
  wire v3a626bd;
  wire v3a54e42;
  wire v377d0e6;
  wire b5a5ab;
  wire v374b5bc;
  wire v3752535;
  wire v3a6efdf;
  wire v372d417;
  wire v3a56114;
  wire v3a705cf;
  wire v372ee18;
  wire v374e18a;
  wire v377c8c8;
  wire v3773250;
  wire v3751ecb;
  wire v3a593cb;
  wire v3a5ff81;
  wire v37440c3;
  wire v3a6ac2a;
  wire v372ecab;
  wire v376f665;
  wire v37575e7;
  wire v372f012;
  wire v377e05a;
  wire v3a70193;
  wire v373c991;
  wire v37764f7;
  wire v376c30b;
  wire v377ccbf;
  wire v3763474;
  wire v3729430;
  wire v3738321;
  wire v3a60bee;
  wire v3a6f645;
  wire v37488d2;
  wire v377aed3;
  wire v3746559;
  wire v3378ef7;
  wire v3a6f343;
  wire v3754272;
  wire v3a6f742;
  wire v3a70ac2;
  wire v3a6f868;
  wire v3741abc;
  wire v3a6f391;
  wire v3a62f68;
  wire v3a5881c;
  wire v376c010;
  wire v3807b9c;
  wire v3a70ca6;
  wire v376b8e1;
  wire v8455ed;
  wire v3a6f7b2;
  wire v3a69ed4;
  wire v3754c09;
  wire v374f4ae;
  wire v374f0bb;
  wire v2aca396;
  wire v8455ef;
  wire v3a6f457;
  wire v374bda9;
  wire v3a563ed;
  wire v376a966;
  wire v3760198;
  wire v37255d6;
  wire v8455d9;
  wire v37723fb;
  wire v8455db;
  wire v3722e5a;
  wire v190eb62;
  wire v3731e3c;
  wire v375ab35;
  wire v2092f0a;
  wire v3a6fa4f;
  wire aca3c3;
  wire v3775b81;
  wire v3a68b6c;
  wire v3772ab6;
  wire v3a558dc;
  wire v376419b;
  wire v3750382;
  wire v3742f7f;
  wire v377f5e0;
  wire v374a8da;
  wire v33789ca;
  wire v375b15b;
  wire v375a59f;
  wire v373a9db;
  wire v3a6f316;
  wire v37714e6;
  wire v3a66d7b;
  wire v3742370;
  wire v3755167;
  wire v3731724;
  wire v375dfcf;
  wire v3735bbb;
  wire v3724014;
  wire v3762363;
  wire v3738f04;
  wire v377bf0d;
  wire v3a6b297;
  wire v3a70cdf;
  wire v372b0f9;
  wire v3a56094;
  wire v373c99b;
  wire v3758e68;
  wire v3776bb6;
  wire v3a70c1a;
  wire v947c98;
  wire v1e3786e;
  wire v377a1ee;
  wire v373e62a;
  wire v3806fe2;
  wire v3752caa;
  wire v374caa8;
  wire v3809e25;
  wire v3732586;
  wire v3a706ef;
  wire v374ff28;
  wire v37519d9;
  wire v3a70615;
  wire v3750c92;
  wire v3a67ab9;
  wire v376fb18;
  wire v375c0cd;
  wire v3a70dea;
  wire v374036a;
  wire v3a5ba7f;
  wire v3a6b6dc;
  wire v3a6efa4;
  wire v377ec1c;
  wire v3754fb0;
  wire v3769628;
  wire v3a5718e;
  wire v374b4da;
  wire v3a611be;
  wire v373ae1e;
  wire v372e8ff;
  wire v372abd2;
  wire v3742d60;
  wire v373226c;
  wire v3747dd0;
  wire v3a605e8;
  wire v3752b4b;
  wire v376f7ab;
  wire v3a703d9;
  wire v3758c50;
  wire v377040f;
  wire v376b1f6;
  wire v377dd4e;
  wire v3a70ed7;
  wire v3808e0d;
  wire v375c8b0;
  wire v3741d51;
  wire v3747276;
  wire v3758c06;
  wire v37351f5;
  wire v375881d;
  wire v372f7ca;
  wire v3a616cb;
  wire v2acaf12;
  wire v3a70d76;
  wire v3a57646;
  wire v2ff9353;
  wire v3a6b463;
  wire v3a6e78d;
  wire v3a6eb2e;
  wire v2ff9190;
  wire v3a71502;
  wire v3752ab6;
  wire v372fe57;
  wire c5b5f4;
  wire v3a6da9c;
  wire v3766438;
  wire v37508b2;
  wire v37390c4;
  wire v372948c;
  wire v39a53f3;
  wire v376c902;
  wire v3a638fb;
  wire v3a60fa3;
  wire v3756f9b;
  wire v3779a3c;
  wire v376db6d;
  wire v3a6fd90;
  wire v37718d5;
  wire v3722ee2;
  wire v37630f1;
  wire v377b3c4;
  wire v9015e2;
  wire v3757b9b;
  wire v3763344;
  wire v3a6ef89;
  wire v374523d;
  wire v3758c15;
  wire v3a70415;
  wire v373f72a;
  wire v377d766;
  wire v3a7076c;
  wire v3a6ca1f;
  wire v3a7044d;
  wire v372840a;
  wire v89b450;
  wire v3a5ffdd;
  wire v3a6f423;
  wire v3a6a7cb;
  wire v37258e7;
  wire v3a707e8;
  wire v3723a2d;
  wire v376f9be;
  wire v3771319;
  wire v3771724;
  wire v376241e;
  wire v3726c99;
  wire v23fd910;
  wire v3a6f409;
  wire v3a6e708;
  wire v3772470;
  wire v3724b93;
  wire v375add8;
  wire v3768538;
  wire v37494a9;
  wire v3778083;
  wire v3725dce;
  wire v3a6f9e8;
  wire v3749d58;
  wire v3733d71;
  wire v37799f4;
  wire v375eb99;
  wire v3a6f4d7;
  wire v3378a0a;
  wire v3742f38;
  wire v377fabc;
  wire v37533c3;
  wire v3a6de73;
  wire v3a6fa06;
  wire v3a5d156;
  wire v3a6a973;
  wire v3a70ca4;
  wire v39eb4ab;
  wire v3773c57;
  wire v377d6e5;
  wire v3750b85;
  wire v37750c2;
  wire v375995f;
  wire v3806882;
  wire v3a6aac8;
  wire v3a61ce5;
  wire v377dc4a;
  wire v373ac95;
  wire v376b706;
  wire v372fddd;
  wire v3748797;
  wire v3a6fde0;
  wire v3a2a107;
  wire v3737808;
  wire v3a70ad0;
  wire v3a6a539;
  wire v3a7098c;
  wire v374e2a1;
  wire v3727507;
  wire v372e169;
  wire v376d34b;
  wire v3723c0d;
  wire v376144f;
  wire v3733727;
  wire v3729531;
  wire v3750f8f;
  wire v3736b57;
  wire v37233a7;
  wire v3726739;
  wire v372342b;
  wire v376bbcc;
  wire v3a70572;
  wire v3727bc1;
  wire v3a59ce1;
  wire v37668b8;
  wire v373b733;
  wire v3a55bfa;
  wire v376a94b;
  wire v3737143;
  wire v374b589;
  wire v3a5e667;
  wire v3741cfb;
  wire v3a6fffd;
  wire v3a6fa4d;
  wire v37522a0;
  wire v360d195;
  wire v377a91a;
  wire v37798bb;
  wire v3753e3b;
  wire v374cffd;
  wire v3a70719;
  wire v3a652db;
  wire v3762e7a;
  wire v377f037;
  wire v373faf3;
  wire v3a6b560;
  wire v2092f5e;
  wire v3a56608;
  wire v3768d29;
  wire v3769112;
  wire v3a6eb1b;
  wire v3a70960;
  wire v3a71473;
  wire v3753ee0;
  wire v3a61de0;
  wire v376b290;
  wire v377c307;
  wire v3739914;
  wire v373c4a7;
  wire v3a6f83b;
  wire v3741793;
  wire v3a6f6cd;
  wire v376f3ae;
  wire v3a7014f;
  wire v3740839;
  wire v3a6fa7e;
  wire v3742b84;
  wire v3a71197;
  wire v3779008;
  wire dbc26f;
  wire v377d27a;
  wire v3724779;
  wire v3a60f21;
  wire v35b7153;
  wire v37325eb;
  wire v3a70129;
  wire v3a54d25;
  wire v3806df2;
  wire v3758357;
  wire v3a70b85;
  wire v377f253;
  wire v3a6f15a;
  wire v372ecad;
  wire v3756f21;
  wire v3a70133;
  wire v377de7f;
  wire v3734279;
  wire v9f45ca;
  wire v372cf70;
  wire v37786f3;
  wire v3a565a1;
  wire v3726c47;
  wire v377aaa9;
  wire v3a56570;
  wire v37680b5;
  wire v373f28d;
  wire v3766246;
  wire v3a70899;
  wire v374fab7;
  wire v375b563;
  wire v3a6f5bf;
  wire v3771f50;
  wire v3754c4a;
  wire v3757a2b;
  wire v3a5c40e;
  wire v3a544c4;
  wire v37573c5;
  wire v3750da4;
  wire v3a70aa8;
  wire v3806a78;
  wire v376ed63;
  wire v3769069;
  wire v3a70474;
  wire v3a7079c;
  wire v37484b6;
  wire v3a6fbf6;
  wire v375c7a3;
  wire v377ece3;
  wire v3a60628;
  wire v37516ba;
  wire v3755f9d;
  wire v3a70854;
  wire v37725c4;
  wire v3a69e59;
  wire v3748a0a;
  wire v3a6fb4f;
  wire v3a70ab3;
  wire v376ec4f;
  wire v3779d91;
  wire v3a6fee3;
  wire v3774253;
  wire v3a6e2ce;
  wire v3748bb7;
  wire v377c0f5;
  wire v38063c6;
  wire v23fdc46;
  wire v3a572b4;
  wire v37483ff;
  wire v3a665d5;
  wire v375c4f9;
  wire v3735fd1;
  wire v373fe61;
  wire v375478f;
  wire v3a6fad9;
  wire v3a5978c;
  wire v3728cfe;
  wire v3a5f5bb;
  wire v376cc8d;
  wire v3a53356;
  wire v3a714b3;
  wire v377728d;
  wire v3a643d7;
  wire v3a71393;
  wire v3577354;
  wire v3a5f9e6;
  wire v3a7168b;
  wire v374a297;
  wire v377085b;
  wire v3a66f35;
  wire v375411b;
  wire v37615a2;
  wire v3a5cd6c;
  wire v375811e;
  wire v3741338;
  wire v3a5741c;
  wire v372fecf;
  wire v37724db;
  wire v3750f49;
  wire v377640c;
  wire v374297b;
  wire v3764312;
  wire v3a6ec1e;
  wire v3a70cc2;
  wire v3a6687c;
  wire v3742290;
  wire v3742aae;
  wire v3769a1e;
  wire v373abde;
  wire v377723a;
  wire v377db1f;
  wire v376047f;
  wire ac1a2c;
  wire v3a6ce39;
  wire v3a5f43a;
  wire v3776454;
  wire v372414d;
  wire v3a7113c;
  wire v37429a1;
  wire v3a691eb;
  wire v3755b4e;
  wire v3a6ff12;
  wire v3740885;
  wire v3a70856;
  wire v37551f2;
  wire v3769f4a;
  wire v37247e2;
  wire bd3fa8;
  wire v377d5d7;
  wire v373e5fb;
  wire v3753353;
  wire v375cea7;
  wire v372b5b0;
  wire v376ff61;
  wire v3a6da33;
  wire v37300c9;
  wire v3778cdd;
  wire v37430c2;
  wire v3752e71;
  wire v373d4fc;
  wire v391331d;
  wire v3731a3b;
  wire v3a5b841;
  wire v374d28d;
  wire v3a6bf41;
  wire v3778454;
  wire v3a63002;
  wire v3743332;
  wire v372408b;
  wire v3a6f910;
  wire v3a713b8;
  wire v3750c12;
  wire v3a700b7;
  wire v374bce0;
  wire v3a5dd86;
  wire v3a69c98;
  wire v377437a;
  wire v3771e60;
  wire v380730d;
  wire v3a64af7;
  wire v3a6212a;
  wire d70af8;
  wire v376e568;
  wire v39eb4de;
  wire v3a61b7f;
  wire v377b4f2;
  wire v372a960;
  wire v372514f;
  wire v3a6eb8b;
  wire v3733f37;
  wire v3a62465;
  wire v3778787;
  wire v3a7026f;
  wire v376062f;
  wire v376c6a8;
  wire v3a5984d;
  wire v375a3dc;
  wire v373f7a5;
  wire v37560ef;
  wire v3758d56;
  wire v37350f0;
  wire v373d791;
  wire v373e1d0;
  wire v3a70388;
  wire v375b0ad;
  wire v37349f9;
  wire v37697f0;
  wire v3a70d3d;
  wire v373402f;
  wire v3a71693;
  wire v3768734;
  wire v3a62b35;
  wire v37586d1;
  wire v37465d4;
  wire v376aaf5;
  wire v375367c;
  wire v3775e35;
  wire v3743831;
  wire v3777da2;
  wire v37652cb;
  wire v2ff8e9c;
  wire v3772715;
  wire v3755136;
  wire v3776516;
  wire v3a67ecb;
  wire v3738491;
  wire v37342f2;
  wire v928541;
  wire v374525d;
  wire v3a61d77;
  wire v3741906;
  wire v37268cc;
  wire v3a60feb;
  wire v3729dea;
  wire v3a66232;
  wire v3a6e5e8;
  wire v3a7158f;
  wire v377dab6;
  wire v3745bc4;
  wire v3a70fd6;
  wire v3a6f35f;
  wire v3a70488;
  wire v375d924;
  wire v376fd4e;
  wire v3a59ea2;
  wire v372afe7;
  wire v37347b2;
  wire v3a53ce6;
  wire v3a7166a;
  wire v37475f4;
  wire v3738259;
  wire v3a637fd;
  wire v3a61388;
  wire v3a6360c;
  wire v3745ae6;
  wire v3a6b864;
  wire v3764caa;
  wire v3760646;
  wire v3761ff9;
  wire v3a63dbf;
  wire v3739334;
  wire v3a5966b;
  wire v38079dc;
  wire v375d445;
  wire v39eb709;
  wire v3756b8a;
  wire v372976e;
  wire v372e30d;
  wire v37609e7;
  wire v372e6f4;
  wire v37352a5;
  wire v376adaf;
  wire v3762a2a;
  wire v376d2dc;
  wire v3a627b3;
  wire v3a5a93a;
  wire v3a59548;
  wire v3772608;
  wire v3753055;
  wire v3730778;
  wire v3a6a02a;
  wire v3a70e4c;
  wire v3733e88;
  wire v3a55ba9;
  wire v360c6b6;
  wire v3378a03;
  wire v3733334;
  wire v3a6670c;
  wire v375f4e8;
  wire v374b320;
  wire v3a6fa55;
  wire v3a66306;
  wire v37675d5;
  wire v3765eee;
  wire v3a55959;
  wire v373f9df;
  wire v377c023;
  wire v3a5621f;
  wire v376d92b;
  wire v3a6f059;
  wire v376eb1d;
  wire v3740060;
  wire aa3e48;
  wire v373cf8f;
  wire ce378e;
  wire v3759c6c;
  wire v3a5fbb0;
  wire v3a6eba5;
  wire v372bf7f;
  wire v373a5a6;
  wire v3a6f160;
  wire v3a58d67;
  wire v3734d8a;
  wire v3a5bd83;
  wire v3a6f633;
  wire v3732f19;
  wire v37251c9;
  wire v3731725;
  wire v3a6d84a;
  wire v376f7d1;
  wire v374e828;
  wire v3769bb0;
  wire v37682bc;
  wire v376827d;
  wire v3a6107c;
  wire v372b48a;
  wire v377c8ca;
  wire v376dc15;
  wire v37429b9;
  wire v3a6e02d;
  wire v3775a4f;
  wire v3a6f04c;
  wire v374748f;
  wire v3a6d500;
  wire v3a5d2bc;
  wire v3747fa9;
  wire v3a697cc;
  wire v3777301;
  wire v3a71131;
  wire v3a6ee78;
  wire v3a7001d;
  wire v3768eac;
  wire v3a70a8f;
  wire v3755090;
  wire v3745012;
  wire v3771a80;
  wire v375daac;
  wire v3763076;
  wire v3770def;
  wire v376eed8;
  wire cd3c6e;
  wire v3a6d10a;
  wire v3a6f62c;
  wire v3a6abdc;
  wire v3a6f79b;
  wire v372a9a6;
  wire v3751291;
  wire v3a70b06;
  wire d5959b;
  wire v373c612;
  wire v375e9b2;
  wire v375eeb0;
  wire v3726460;
  wire v3749655;
  wire v3746cc0;
  wire v373d219;
  wire v3777d1f;
  wire v3a713f4;
  wire v374de48;
  wire v374fb40;
  wire v375c976;
  wire v3779a88;
  wire v3a7002a;
  wire v3763252;
  wire v3809d8b;
  wire v377baf4;
  wire v3747d30;
  wire v35b9d58;
  wire v375c4b0;
  wire v377a27c;
  wire v3a6c0c1;
  wire v37702e0;
  wire v373b42d;
  wire v3a70426;
  wire v3a715ce;
  wire v376321e;
  wire v3739a9f;
  wire v3728581;
  wire v372ab42;
  wire v374ea10;
  wire v3a6e7ae;
  wire v3744dda;
  wire v3769753;
  wire v376f1d0;
  wire v3777602;
  wire v377f694;
  wire v375c1a7;
  wire v377577b;
  wire v373f408;
  wire v3a5548b;
  wire v372a04c;
  wire v372539e;
  wire v3a700b6;
  wire v372e821;
  wire v377d945;
  wire v35b779e;
  wire v3a6049f;
  wire v3734df5;
  wire v3a5c5e1;
  wire v374c9d9;
  wire v3753404;
  wire v3750559;
  wire v375fecf;
  wire v3747ced;
  wire v3727477;
  wire v374dae3;
  wire v3742f1b;
  wire v3736e1d;
  wire v3a61668;
  wire v3778251;
  wire v377bbbb;
  wire v3a58530;
  wire v37391a1;
  wire v3a6fdb0;
  wire v372fc07;
  wire v9fa0b5;
  wire v3751dd7;
  wire v376c4f9;
  wire v3a71356;
  wire v3740975;
  wire v3740d9a;
  wire v375df5e;
  wire v375fae9;
  wire v23fe209;
  wire v3779cda;
  wire v3755901;
  wire v374fa1e;
  wire v3747b4c;
  wire v373df9c;
  wire v3a6f149;
  wire v374cb4a;
  wire v3a5617a;
  wire v3a5a16b;
  wire v375d05d;
  wire v37326a5;
  wire v3a6e804;
  wire v3a6f2ad;
  wire v3777071;
  wire v3a70ab0;
  wire v376fefa;
  wire v374a7de;
  wire v3a63e9d;
  wire v3775072;
  wire v37730b3;
  wire v37339b7;
  wire v37762ec;
  wire v37c0170;
  wire v37628f3;
  wire v373b647;
  wire v3a54484;
  wire v3a70f7c;
  wire v360cd91;
  wire v37580b6;
  wire v37660f0;
  wire v3727e25;
  wire v376ac10;
  wire v376fb07;
  wire v3740be8;
  wire v37362dc;
  wire v3739769;
  wire v37528b8;
  wire v3a6950d;
  wire v375b96f;
  wire v3777b5f;
  wire v3a7067e;
  wire v37444e7;
  wire v3808e3a;
  wire v3a6fa99;
  wire v373766f;
  wire v3a5f609;
  wire v3729c9a;
  wire v3a7050d;
  wire v3a700d2;
  wire v373d81e;
  wire v3766b6e;
  wire v373d661;
  wire v3a68707;
  wire v3806847;
  wire v375b320;
  wire v3a56855;
  wire v374c297;
  wire v3a6f92d;
  wire v3741863;
  wire v3772dcb;
  wire v3a6d0ae;
  wire v37474c1;
  wire v3771c6a;
  wire v377456d;
  wire v3a636c0;
  wire v3734ca9;
  wire v377bd81;
  wire v374b330;
  wire v373fbc9;
  wire v377cdf0;
  wire v3739a3b;
  wire v3a715a8;
  wire d6eddf;
  wire v3a70a5e;
  wire v37658f9;
  wire v375a202;
  wire v374a3f3;
  wire v3741afa;
  wire v3a5d882;
  wire v3a63a46;
  wire v375ab99;
  wire v3727df1;
  wire v8fac55;
  wire v3a6991b;
  wire v32574c7;
  wire v37499a0;
  wire v376f499;
  wire v3745cea;
  wire v3a6ebfb;
  wire v377ec50;
  wire v3a58cd4;
  wire v3a6218f;
  wire v3747114;
  wire baea86;
  wire b88b06;
  wire v3748560;
  wire v3a6b18b;
  wire v375c75c;
  wire v372e708;
  wire v373096c;
  wire v3a71458;
  wire v375b9a0;
  wire v3a70e60;
  wire v3738c75;
  wire v3a539af;
  wire v377d651;
  wire v3742e6b;
  wire v3a57741;
  wire c81b97;
  wire v377cda9;
  wire v3a65019;
  wire v380705b;
  wire v1e373d9;
  wire v375ac88;
  wire v37355e3;
  wire v373e4ca;
  wire v3a61964;
  wire v373c8a4;
  wire v2092fa9;
  wire v372e775;
  wire v374a7c3;
  wire v376e2bb;
  wire v2ff918d;
  wire v3a701b1;
  wire v372e967;
  wire v3a70b9b;
  wire v377081e;
  wire v37629fc;
  wire d950cb;
  wire v376d23f;
  wire v37531ca;
  wire v3730398;
  wire v37345de;
  wire v372a309;
  wire v376e1fb;
  wire v3a593b0;
  wire v3a67715;
  wire v374d246;
  wire v3a715cb;
  wire v3736779;
  wire v37423c1;
  wire v3a70ad5;
  wire v3a705b0;
  wire v376f98e;
  wire v3a70008;
  wire v3735e52;
  wire v3a56ffa;
  wire v37742d2;
  wire v3a603e0;
  wire v377536e;
  wire v3a5ad94;
  wire v37434f4;
  wire v375a6e6;
  wire v3768130;
  wire v37565be;
  wire v3a7126c;
  wire v31c369c;
  wire v1e37556;
  wire v3729030;
  wire v3727ed2;
  wire v3a6f2d1;
  wire v3761d38;
  wire v377b015;
  wire v374ed0a;
  wire v3809752;
  wire v3775a92;
  wire v3745b0f;
  wire v3723e5d;
  wire v92a03a;
  wire v3a5cb6f;
  wire v377d045;
  wire v3724069;
  wire v377a291;
  wire v3a70734;
  wire v3743dae;
  wire v3a6ebf8;
  wire v376dc16;
  wire v3a70728;
  wire v3a6af67;
  wire v37294db;
  wire v37525c7;
  wire v3755a83;
  wire v377f6ae;
  wire v3a66c9a;
  wire v3a6c905;
  wire d38ecb;
  wire v3a6f9e5;
  wire v3761bb7;
  wire v3a6d6be;
  wire v3a5c58f;
  wire v37428ac;
  wire v372ebaa;
  wire v3759d36;
  wire v377d705;
  wire v3a6f0cc;
  wire v376fc36;
  wire v3a587bc;
  wire v372f6ce;
  wire a17325;
  wire v377123e;
  wire v377c551;
  wire v373a349;
  wire v3a6db1a;
  wire v37233d2;
  wire v3725cc8;
  wire v3763150;
  wire v38063a0;
  wire v3a62aef;
  wire v372b3f6;
  wire ae0bd0;
  wire v3730651;
  wire v377b3b0;
  wire v3a6ff89;
  wire v377661b;
  wire v3a65bb1;
  wire v375c735;
  wire v376f5ed;
  wire v376d3a6;
  wire v377b838;
  wire v3a703f7;
  wire v3a71360;
  wire v372f8d3;
  wire v3a6f2b8;
  wire v3a66e70;
  wire v374b256;
  wire v373193a;
  wire v377028b;
  wire v3a633a7;
  wire v373a5b6;
  wire v3747b3c;
  wire v3a6d558;
  wire v3a6c007;
  wire v3a5a16a;
  wire bb97e8;
  wire v3724703;
  wire v376d4ca;
  wire v37623b8;
  wire v3a6af1d;
  wire v3a7138a;
  wire v3a6f8d7;
  wire v3a61ecf;
  wire v3a69b74;
  wire v3a64f05;
  wire v375afc1;
  wire v377228d;
  wire v374b20c;
  wire v3a6efd2;
  wire v374dffc;
  wire v3724e2a;
  wire v3a7046b;
  wire v374ce71;
  wire v372de3b;
  wire v376f504;
  wire v373794a;
  wire v374b4f8;
  wire v374b7d8;
  wire v3a6f373;
  wire v2619ad3;
  wire v37479b4;
  wire v3744f52;
  wire v3a5c27f;
  wire v380930a;
  wire v375fbe8;
  wire v3a63dcc;
  wire v374fa0d;
  wire v377f611;
  wire v3a571b6;
  wire v3a71540;
  wire v3766727;
  wire v3a5bbeb;
  wire v3a552d2;
  wire v3725e96;
  wire v3a7116a;
  wire v37620eb;
  wire v373dfb4;
  wire v372e7f8;
  wire v373abdd;
  wire v374476d;
  wire v3a60924;
  wire v37389ba;
  wire v3a56200;
  wire v3a60642;
  wire v374a60b;
  wire v377e04e;
  wire v3767be8;
  wire v373de1d;
  wire v37630e2;
  wire v3a55078;
  wire v37354bf;
  wire v374e1f0;
  wire v37393e8;
  wire v3a54a24;
  wire v374ee77;
  wire v3761aa3;
  wire v3744f80;
  wire v377a6c4;
  wire v2ff87db;
  wire v8455b3;
  wire v3a6c2b6;
  wire v3a5eadd;
  wire v1e37cd6;
  wire v376a6f1;
  wire v373ad69;
  wire v3722dd5;
  wire v377f7dd;
  wire v3752ec0;
  wire v3a6eb6b;
  wire v374d2b3;
  wire v377349f;
  wire v3758fa8;
  wire v3724d93;
  wire v3761efb;
  wire v3a703d3;
  wire v37684a8;
  wire v3a6fd72;
  wire v8455e9;
  wire v3742d37;
  wire v3a55349;
  wire v377c31d;
  wire v3749a32;
  wire v3735272;
  wire v1e37b76;
  wire v3761d2f;
  wire v372543f;
  wire v3a5b71a;
  wire v3744710;
  wire v3776a6e;
  wire v3a5903a;
  wire v374ac2c;
  wire c0d46a;
  wire v377c039;
  wire v39eb4a7;
  wire v3a71686;
  wire v3a6a1df;
  wire c35240;
  wire v374bfcf;
  wire v374f318;
  wire v375fabf;
  wire v372f532;
  wire v3a6e5f4;
  wire v372bbb3;
  wire v3a711da;
  wire c7355c;
  wire v375f1ee;
  wire v374950c;
  wire v3770bcd;
  wire v3a6eb3d;
  wire v3735f67;
  wire v377d9b2;
  wire v3a7011b;
  wire v3731a2e;
  wire v3a6aabc;
  wire v372fd00;
  wire v3a6ebb8;
  wire v37665c5;
  wire v37744a3;
  wire v3763086;
  wire v8455c1;
  wire v3a5cc27;
  wire v375ecf8;
  wire v3755082;
  wire v37361a0;
  wire v373270f;
  wire v3807a23;
  wire v372cac5;
  wire v3a5f02e;
  wire v3a713c5;
  wire v37496de;
  wire v3a70276;
  wire d52046;
  wire v3760690;
  wire v373216d;
  wire v3806b0b;
  wire v3a578c3;
  wire v373c30e;
  wire v377047f;
  wire v3a702fd;
  wire v3a62e91;
  wire v373dc1c;
  wire v374d3d7;
  wire v3747d3c;
  wire v3766218;
  wire v374c0e4;
  wire v3738c99;
  wire v37311d6;
  wire v372673b;
  wire v374b1ea;
  wire v3770eb9;
  wire v3746259;
  wire v373bcb6;
  wire v3a58b13;
  wire v373c372;
  wire v3761bac;
  wire v3a713b0;
  wire v3a62f05;
  wire v3a70143;
  wire v3a5ba8a;
  wire v375be2d;
  wire v1e37a30;
  wire v374c154;
  wire v3768f5f;
  wire v3a5b576;
  wire v3768c25;
  wire v3a59de6;
  wire v3a6947c;
  wire v3746fe7;
  wire v376f111;
  wire v38064e5;
  wire c9c058;
  wire v377695e;
  wire v3a5e684;
  wire v3724b74;
  wire v37530c7;
  wire v372bdd9;
  wire v37661db;
  wire v3729e38;
  wire v3a7047c;
  wire db6de7;
  wire v375887e;
  wire v377c28e;
  wire v37793b9;
  wire v37798b9;
  wire v3a61f85;
  wire v374f21c;
  wire v372895b;
  wire v3a6fc61;
  wire v3735a25;
  wire v373ca9e;
  wire v37435e1;
  wire v3a6fddb;
  wire v3774e2b;
  wire v3735b3d;
  wire v3775498;
  wire v376614e;
  wire v377168f;
  wire v3774e9d;
  wire bdb49d;
  wire v375a235;
  wire a8afe1;
  wire v38097db;
  wire v377e31b;
  wire v2ff9287;
  wire v3a606e8;
  wire v3a6f243;
  wire v3725ec4;
  wire v3a656b6;
  wire v373a822;
  wire b5da28;
  wire v3755549;
  wire v8455bd;
  wire v377803f;
  wire v37604b3;
  wire v375248f;
  wire v3742be5;
  wire v3750c0c;
  wire v3809af2;
  wire v37482bb;
  wire v2ff8f1e;
  wire v375d30b;
  wire v376d82f;
  wire v3a6fa28;
  wire v3a6e4de;
  wire v3a64374;
  wire v3767904;
  wire v377affd;
  wire v376f277;
  wire v377ca3b;
  wire v3a64968;
  wire v3a71295;
  wire v3726b10;
  wire v3a63f0c;
  wire v3768495;
  wire v372ec4e;
  wire afdeb4;
  wire v3a55cda;
  wire v3a56a86;
  wire v3a70419;
  wire v37685f1;
  wire v3a5c349;
  wire v376ef20;
  wire v3a6b336;
  wire v372562a;
  wire v3756aa3;
  wire v3a6514f;
  wire v3a5ce6f;
  wire v372cb42;
  wire v3a71188;
  wire v3768589;
  wire v3a66c5c;
  wire v3a5846c;
  wire v37501f3;
  wire v3745241;
  wire v372abac;
  wire v3762dc3;
  wire v3a55290;
  wire v372a1b4;
  wire v372cacb;
  wire v377e345;
  wire v3762651;
  wire v375c573;
  wire v3a71132;
  wire v3729829;
  wire v37668e2;
  wire v37255de;
  wire v3a712d3;
  wire v376799e;
  wire b72b90;
  wire v3a6fa72;
  wire v373b286;
  wire v3745ce8;
  wire v3765576;
  wire v375afe9;
  wire v37388a7;
  wire v3a6ff5b;
  wire v372294a;
  wire v3a659f5;
  wire v3a2aed2;
  wire v3a53977;
  wire v37262ab;
  wire v3a6fba3;
  wire v3742a4d;
  wire v374bb16;
  wire v372f721;
  wire v373c268;
  wire v377435d;
  wire v375fe58;
  wire v375c7cf;
  wire v376f38d;
  wire v375c01d;
  wire v3758a0c;
  wire v3a5a967;
  wire v37435f6;
  wire v3a65a33;
  wire v374c1a9;
  wire v3a7012d;
  wire v3a6f12a;
  wire v37788a6;
  wire v3738ed8;
  wire v376ab39;
  wire v3a6adf2;
  wire v376f516;
  wire v37482c7;
  wire v377ac1e;
  wire v3743a77;
  wire v3a6f974;
  wire v373c5ea;
  wire v3a5d365;
  wire v374490b;
  wire v373f64f;
  wire v3747130;
  wire v3773d27;
  wire v3748fde;
  wire v376a04d;
  wire v3a5b807;
  wire v37560c9;
  wire v374fefc;
  wire v3a706d9;
  wire v37440ff;
  wire v3a62122;
  wire v3760629;
  wire v37571da;
  wire v3a6fc9b;
  wire v3a702de;
  wire v374c23c;
  wire v2619ac3;
  wire v3a7133f;
  wire v3a593bb;
  wire v37411df;
  wire v3a588ef;
  wire v373c4d4;
  wire v37577b7;
  wire v376300a;
  wire v23fdebb;
  wire v372d1f0;
  wire v3a705c7;
  wire v37390f0;
  wire v3727387;
  wire v3a70d23;
  wire v3a6e552;
  wire v3a710c5;
  wire v373647a;
  wire v3a6fd77;
  wire v3748c3f;
  wire v3736257;
  wire v373db92;
  wire v375bbe2;
  wire v377dac2;
  wire v374b24a;
  wire v376a3f7;
  wire v3773137;
  wire bee241;
  wire v3a70362;
  wire v3741833;
  wire v37369eb;
  wire v372e3d8;
  wire v3a7115a;
  wire v37647d8;
  wire v3750b22;
  wire v377de07;
  wire v3761e59;
  wire v37421c0;
  wire v372b6d0;
  wire v3761a8f;
  wire v3a6dd22;
  wire v3762613;
  wire v37541d4;
  wire v374cb0f;
  wire v3748400;
  wire v3a71518;
  wire v3776ae5;
  wire v374de73;
  wire v373c688;
  wire v3a5aaca;
  wire v375f87a;
  wire v37446d8;
  wire v3a60638;
  wire ad7e3b;
  wire v3a6ff58;
  wire v372d816;
  wire v3730b5e;
  wire v375d0cf;
  wire v3742dae;
  wire v3746fd4;
  wire v3a5b57a;
  wire v3a6ebc3;
  wire v3a6866f;
  wire v3745d9c;
  wire v373fe48;
  wire v3729435;
  wire v3a714c5;
  wire v209300b;
  wire v3a6ff07;
  wire v3a65160;
  wire v3a6f662;
  wire v373b130;
  wire v3a5ea57;
  wire v3762396;
  wire v3737c1c;
  wire v372ab1b;
  wire v375c54c;
  wire v374d529;
  wire v3a59b42;
  wire v3a703b8;
  wire v37368d0;
  wire v373b6e4;
  wire v3a60c59;
  wire v3759512;
  wire v375975b;
  wire v375564e;
  wire v375058e;
  wire v372cdde;
  wire v380731d;
  wire v374c885;
  wire v374592e;
  wire v3a708aa;
  wire v3809adf;
  wire v3a648f2;
  wire v3773a3d;
  wire v3a6efc4;
  wire v3748422;
  wire v3745f76;
  wire v373f06b;
  wire v372dccf;
  wire v372f309;
  wire v3a58429;
  wire v3a6a3e6;
  wire v377b460;
  wire v374f5d6;
  wire v3a61e6a;
  wire v3a69487;
  wire v3a5fc34;
  wire v3736679;
  wire v373e114;
  wire v3746b73;
  wire v3770ff9;
  wire v377dc99;
  wire v3a709e8;
  wire v3a70fd5;
  wire v37367a0;
  wire v3a61ab0;
  wire v3735050;
  wire v959f2d;
  wire v37281a4;
  wire v3754b66;
  wire v3743486;
  wire v3a6ffdc;
  wire v3a6f4b5;
  wire v3734200;
  wire v3a6fe90;
  wire v3a67c13;
  wire v3a701e4;
  wire v3730ae3;
  wire v3759749;
  wire v373c3e1;
  wire v3a6ae45;
  wire v376b509;
  wire c61447;
  wire v37484df;
  wire v375d0ed;
  wire v3761ca9;
  wire v377b423;
  wire v1e37d8e;
  wire v3a6d9ca;
  wire v3748229;
  wire v3a631d0;
  wire v375f27b;
  wire v3a5c1a5;
  wire v3761ad0;
  wire v372914b;
  wire v3757559;
  wire v3728d14;
  wire v3742f64;
  wire v37434e1;
  wire v37783ba;
  wire v1e37349;
  wire v373d081;
  wire v374835b;
  wire v376753a;
  wire v372ff79;
  wire v374cf44;
  wire v376d1e2;
  wire v375b2e2;
  wire v37348ee;
  wire v375911a;
  wire v37514c7;
  wire v374de0d;
  wire v374fe1a;
  wire v374b992;
  wire v3a6f496;
  wire v374ac60;
  wire v3a6fd53;
  wire v3750fc9;
  wire v3a5d469;
  wire v374355e;
  wire v372da78;
  wire v377bf71;
  wire v3773506;
  wire v375820e;
  wire v376f4c5;
  wire v3730060;
  wire v3a6c31f;
  wire c46b05;
  wire v377800b;
  wire v3a6f2de;
  wire v377f887;
  wire v3a70555;
  wire v3a6471a;
  wire v376d6ef;
  wire v3a65e9d;
  wire v38092a9;
  wire v3744940;
  wire v375c7cb;
  wire v37294d3;
  wire v376e854;
  wire v3a710e3;
  wire v3a6b8aa;
  wire v3751acf;
  wire v375f847;
  wire v37735b8;
  wire v3739ab6;
  wire v3a710f4;
  wire v3723da9;
  wire v3736be1;
  wire v3a634eb;
  wire v372490a;
  wire v3a6fd7e;
  wire v3a6fc41;
  wire v3a70bbe;
  wire v375790e;
  wire v3a56d3a;
  wire v3a703e4;
  wire v3a63512;
  wire v3a63bbc;
  wire v9181c9;
  wire v372d2ad;
  wire v3729852;
  wire v3a62a13;
  wire v3778e28;
  wire v3729d1a;
  wire v3a5e748;
  wire v3a70006;
  wire v3726ae2;
  wire v23fe339;
  wire v3a6fad6;
  wire v377d86e;
  wire v3751ab7;
  wire v3807a47;
  wire v37510b1;
  wire v374922a;
  wire v374f028;
  wire v376f2a5;
  wire v3725496;
  wire v3a6f335;
  wire v3748266;
  wire v3726845;
  wire v3a59409;
  wire v3746265;
  wire v373a47e;
  wire v3760309;
  wire v2678c97;
  wire v3a5e7dc;
  wire v372f289;
  wire v374da92;
  wire v3a70ce5;
  wire v3a69fcf;
  wire v3a6f5e4;
  wire v3746f4c;
  wire v3777c6d;
  wire d60033;
  wire v37422af;
  wire v377d414;
  wire v3a7039c;
  wire v377f0e7;
  wire v3a576a4;
  wire v3a70356;
  wire v372fb63;
  wire v3a706f0;
  wire v37240c0;
  wire v3a7127c;
  wire v3a5b875;
  wire v3759611;
  wire v3739b37;
  wire v3771171;
  wire v3a680eb;
  wire d692cc;
  wire v3a6f730;
  wire v3a56918;
  wire v3759663;
  wire v374a7f2;
  wire v375be00;
  wire v37597f7;
  wire v3a7031c;
  wire v3378b6c;
  wire v3808d68;
  wire v37721fa;
  wire v3a6eb02;
  wire v373f90a;
  wire v376f2fc;
  wire v377cdf1;
  wire v3736b93;
  wire v375a8db;
  wire v373cba8;
  wire v3740b8c;
  wire v3a6f261;
  wire b539d9;
  wire v3745e54;
  wire v3a67755;
  wire v37666d7;
  wire v374c009;
  wire v37729c7;
  wire v3a711e7;
  wire v376c644;
  wire v3a709af;
  wire db9e30;
  wire v3a5dde7;
  wire v373f911;
  wire v372d060;
  wire v3747079;
  wire v8455c9;
  wire v375e53a;
  wire v3728392;
  wire v3a6fd62;
  wire v3a6a872;
  wire v37278fd;
  wire v375a83f;
  wire v3730d6a;
  wire v3809d6a;
  wire v3723400;
  wire v38097a9;
  wire v3a7076d;
  wire v3a6f541;
  wire v37706dd;
  wire v3a58bb0;
  wire v37613bf;
  wire v3777f01;
  wire v372f89e;
  wire v3a71008;
  wire v37400d8;
  wire v3a592d8;
  wire v3a57b5a;
  wire v3752da9;
  wire v377987e;
  wire v3772616;
  wire v37600ad;
  wire v37331a2;
  wire v3a703e2;
  wire v3a5dfa3;
  wire v3a6f88a;
  wire v37c37ed;
  wire v375e85e;
  wire v373665b;
  wire v37763b2;
  wire v3a6a95e;
  wire v3730b63;
  wire v377433b;
  wire v3a5e90f;
  wire v3a71247;
  wire v3a6603f;
  wire v3746a62;
  wire v373a693;
  wire v3724936;
  wire v372e0fc;
  wire v377ba41;
  wire v373d35d;
  wire v3a70359;
  wire v37331d1;
  wire v3770c2a;
  wire v376d640;
  wire v37514e4;
  wire v3739b7a;
  wire v372e4a7;
  wire v374a369;
  wire v372e4ac;
  wire v3777498;
  wire v3a5b4bd;
  wire v3757d5b;
  wire v3769c43;
  wire v372d238;
  wire v37376f9;
  wire v37354b5;
  wire v3a70a3b;
  wire v3757b58;
  wire v3731fd8;
  wire v376a254;
  wire v375a990;
  wire v3a5b39d;
  wire v376b5c6;
  wire v372ddfa;
  wire v3765396;
  wire v3726810;
  wire v3a711e8;
  wire v37508b9;
  wire v37586bb;
  wire v3769215;
  wire v37674d1;
  wire v3751606;
  wire v3a70015;
  wire v3a6ecb7;
  wire v3776f2c;
  wire v3a2a41f;
  wire v3a54b84;
  wire v3809142;
  wire v3a6f437;
  wire v377ea1b;
  wire v374897d;
  wire v3736d87;
  wire v3769c19;
  wire v3a6f0f7;
  wire v376513f;
  wire v3a66940;
  wire v3a7155b;
  wire v3a5af26;
  wire v3776e33;
  wire v3a70cb3;
  wire v372a94f;
  wire d3ed45;
  wire v3a6f6f1;
  wire v377a571;
  wire v375d966;
  wire v9c8578;
  wire v377d8c8;
  wire v3a6f3fa;
  wire v3765d9e;
  wire v3735055;
  wire b20520;
  wire bfe049;
  wire v372cc01;
  wire v376cda5;
  wire v3a71083;
  wire v377dc20;
  wire v3723583;
  wire v3748126;
  wire v376b744;
  wire v377b209;
  wire v3730e4c;
  wire v3a70029;
  wire v376b036;
  wire v3a6fa2a;
  wire v1e37d3a;
  wire v1e37e29;
  wire v3a62aa3;
  wire v37386af;
  wire v3740ab8;
  wire v3764f06;
  wire v376d559;
  wire v372c064;
  wire v3726eea;
  wire v3a581f1;
  wire v372bdb1;
  wire v23fd869;
  wire v375cb5e;
  wire v3772c9f;
  wire v37269b2;
  wire v3a665ca;
  wire v375e993;
  wire c7ae7d;
  wire v37317da;
  wire v3a6b32d;
  wire v375de73;
  wire v3a62875;
  wire v3a6fc08;
  wire v3a57311;
  wire v376fddd;
  wire v373977e;
  wire v3758cec;
  wire v3a6d6fe;
  wire v3a6fa9f;
  wire v375dbe0;
  wire v3735f02;
  wire v3769981;
  wire v3a6fadc;
  wire v3751b37;
  wire v372a24d;
  wire v3a716a4;
  wire v37368d3;
  wire v3a66b26;
  wire v3768264;
  wire v37305cc;
  wire v3a68b74;
  wire v3a6fd65;
  wire v37548e6;
  wire v3a5bb4f;
  wire v3756516;
  wire v377bf88;
  wire v3744693;
  wire v3771c3a;
  wire v3751364;
  wire v3761f39;
  wire v3a6f119;
  wire v3a70b66;
  wire v3a5c858;
  wire v372998a;
  wire v37666dd;
  wire v376725e;
  wire v3a6abf7;
  wire v375fb9d;
  wire v375c65f;
  wire v37756f8;
  wire v3a53709;
  wire v3722ba9;
  wire v3736421;
  wire v377f785;
  wire v3a7155c;
  wire v3745bbe;
  wire v3767638;
  wire v37263bf;
  wire v37678e2;
  wire v376e029;
  wire v3a660e6;
  wire v377e493;
  wire v373af1f;
  wire v3a66e96;
  wire v377e864;
  wire v375af58;
  wire v3739190;
  wire v375b68b;
  wire v3a55482;
  wire v38064e4;
  wire a875ea;
  wire v3761d4e;
  wire v37283fc;
  wire v3a5e24d;
  wire v3a54bc5;
  wire v3a712e6;
  wire v337947a;
  wire v372c42d;
  wire v373180e;
  wire v3777a07;
  wire v376f978;
  wire v376282b;
  wire v3a7091d;
  wire v37324c0;
  wire v377c47d;
  wire v373a26e;
  wire v3743690;
  wire v3725ef7;
  wire v3735593;
  wire v3a6fc53;
  wire v37728a4;
  wire v3a708ec;
  wire v374063d;
  wire v3a6efd1;
  wire c58ea1;
  wire d4de60;
  wire v3a5def2;
  wire v3a70554;
  wire a747d7;
  wire v377492b;
  wire v373552a;
  wire v3a5dd1a;
  wire v3a70827;
  wire v380a2f5;
  wire v3753bac;
  wire v23fde92;
  wire v90829e;
  wire v375bd1f;
  wire dab321;
  wire v3725310;
  wire v375bc6e;
  wire v3a6613e;
  wire v3a6fc11;
  wire v3a70906;
  wire v374550d;
  wire v3a6890e;
  wire v3768616;
  wire v3a5aa33;
  wire v3a682f7;
  wire v374a510;
  wire v3770690;
  wire v3779233;
  wire v3a6776f;
  wire v3a58589;
  wire v372cdf6;
  wire v3755f9b;
  wire v3752c4d;
  wire v3753429;
  wire v373142a;
  wire v3752304;
  wire v3a6ff9b;
  wire v3a6d349;
  wire v373588a;
  wire v373e12e;
  wire v372475a;
  wire v374fa0a;
  wire v37510ae;
  wire v3a5ee3a;
  wire v3758ff4;
  wire v3a6fdcc;
  wire v376fe6e;
  wire v3a6e96b;
  wire v3752798;
  wire v3a710b3;
  wire v3a6fab3;
  wire v3758532;
  wire v3a6f724;
  wire v3a6f4ca;
  wire v3a5463b;
  wire v3a608c4;
  wire v37322ca;
  wire v3764998;
  wire v374ddcd;
  wire v375b943;
  wire v3a67ffe;
  wire v3808d2e;
  wire v374c523;
  wire v373b303;
  wire v374d6f4;
  wire v3a703d1;
  wire v3771ae3;
  wire v3764463;
  wire v3749c22;
  wire v3806572;
  wire v3751ca5;
  wire v3a60bc8;
  wire c858c6;
  wire v3750f2a;
  wire v3776c9a;
  wire v374f0a4;
  wire v375bb6b;
  wire v3a707c7;
  wire v372b2ba;
  wire v3a5ee7d;
  wire v3778637;
  wire v3768b3d;
  wire v377eda6;
  wire v37bfc35;
  wire v3a5ead4;
  wire v377e3ce;
  wire v3a67142;
  wire v3744934;
  wire v3a67221;
  wire v37780cd;
  wire v3732bc1;
  wire v3725f98;
  wire v376d9d4;
  wire v2acb088;
  wire v3a5e8f6;
  wire v23fe285;
  wire v374047d;
  wire v37381f0;
  wire v3728ca9;
  wire v3a6acab;
  wire v37563fe;
  wire v3a6f557;
  wire v372a4c3;
  wire v372d0de;
  wire v376410a;
  wire v373b671;
  wire v3a5787a;
  wire v3a6908b;
  wire v37799ca;
  wire v39eaa60;
  wire v3743788;
  wire v37518ac;
  wire v376a26b;
  wire v3771ea2;
  wire v3723bf9;
  wire v374a601;
  wire v3a6c9c2;
  wire v373ca4f;
  wire v3768b81;
  wire v3a66668;
  wire v3a5706c;
  wire v372e468;
  wire v3723cff;
  wire v372b74c;
  wire v3753ca0;
  wire v3778962;
  wire v3a6ec03;
  wire v372e669;
  wire v373894d;
  wire v377306c;
  wire v377535e;
  wire v3a6f8c0;
  wire v375f3cf;
  wire v3775928;
  wire v373df1f;
  wire c4d24d;
  wire v3726088;
  wire v372ded7;
  wire v377714d;
  wire v3a627d8;
  wire v374efee;
  wire v373a984;
  wire v3a71098;
  wire v377894b;
  wire v376b576;
  wire v3770e2d;
  wire v3a57f41;
  wire v3a6eb55;
  wire v3a70654;
  wire v3a6d37f;
  wire v373913a;
  wire v374500f;
  wire v376070d;
  wire v3a70f5d;
  wire v3a67588;
  wire v3a68fd3;
  wire v377047a;
  wire v3773ca3;
  wire v3a70a99;
  wire v3734658;
  wire v3a6f593;
  wire v3733664;
  wire v375c999;
  wire v3a5a2a4;
  wire v375b6d4;
  wire v3a65565;
  wire v38094ca;
  wire v3730bd8;
  wire v3755b5c;
  wire v373ca3d;
  wire v3a6eede;
  wire v377f170;
  wire v376967e;
  wire v3729ee6;
  wire v3745b66;
  wire v3768774;
  wire v3a71020;
  wire v3a6f7c7;
  wire v373bfab;
  wire v3a70d01;
  wire v3776c04;
  wire v38093aa;
  wire v3752957;
  wire v37274be;
  wire v3767304;
  wire v3a6fc29;
  wire v3744ca2;
  wire v3a64e91;
  wire v3a6f5f6;
  wire v3749bef;
  wire v3a6bedb;
  wire v3a60a23;
  wire v37425a5;
  wire v37517f4;
  wire v3765053;
  wire v3a708ad;
  wire v3a6f310;
  wire v375e752;
  wire v3a6f9df;
  wire v376e0fa;
  wire v3768ec4;
  wire v377f4e5;
  wire v376acee;
  wire v373fa89;
  wire v3a708f6;
  wire v37536c3;
  wire v3a6708c;
  wire v3749b09;
  wire v3777a52;
  wire v3776d97;
  wire v3a5d555;
  wire v37603a3;
  wire v3a71335;
  wire v3a6f6b6;
  wire v37746ea;
  wire v37652eb;
  wire v3a705a6;
  wire d8c443;
  wire v3a6f11c;
  wire v374648f;
  wire v3a6ef3f;
  wire v372a61c;
  wire v3a70969;
  wire v3726c67;
  wire v374c70d;
  wire v375c705;
  wire v3a702a0;
  wire v376a20e;
  wire v3754076;
  wire v376f178;
  wire v37390ed;
  wire v3741a9b;
  wire v3769010;
  wire v373b88a;
  wire v3728127;
  wire v3778b19;
  wire v39a5380;
  wire v3a53e5b;
  wire v3a71467;
  wire v376079f;
  wire v372b268;
  wire v3755a02;
  wire v375a95b;
  wire v377b6b2;
  wire v8dfd63;
  wire v39eaff9;
  wire v37541b4;
  wire v375548b;
  wire v37451b6;
  wire v376bd2f;
  wire v374f8f6;
  wire v3768918;
  wire v372b3dd;
  wire v3a6f555;
  wire v37774d3;
  wire v376fe45;
  wire v37356aa;
  wire v37446e0;
  wire v3a6738e;
  wire v3a7113b;
  wire v3a55081;
  wire v37400d2;
  wire v3a5b719;
  wire v3a6196d;
  wire v3733641;
  wire v374e3fa;
  wire v3a71527;
  wire v375fd8d;
  wire v3734292;
  wire v37786bb;
  wire v3a53f00;
  wire cc2c2e;
  wire v3a56187;
  wire v374d654;
  wire v37427cf;
  wire v3a6f36e;
  wire v375dcdb;
  wire v3768b07;
  wire v373376b;
  wire v3a605e2;
  wire v374fd8a;
  wire v374c58c;
  wire v373df89;
  wire v375fc0a;
  wire v374e0e9;
  wire v3a6ef2e;
  wire v37307d7;
  wire v374d47d;
  wire v377cd5b;
  wire v374f7b7;
  wire v377f15c;
  wire v3750002;
  wire v3a6c7ef;
  wire v3747800;
  wire v3743851;
  wire v3a70562;
  wire v3a705ef;
  wire v3a6ad1f;
  wire v3774cee;
  wire v373a013;
  wire v380a1a6;
  wire v37691fa;
  wire v3a70624;
  wire v23fe189;
  wire v39eb532;
  wire v37444b2;
  wire v3736e8e;
  wire v3a6d4b7;
  wire v375796c;
  wire v3751b35;
  wire v3767080;
  wire v3a6fdb3;
  wire v375bd37;
  wire v37477aa;
  wire v376fc1c;
  wire v3731383;
  wire v375b142;
  wire v377e39f;
  wire v3a58762;
  wire v3757e0b;
  wire v3a56fcd;
  wire v376d387;
  wire v3a6c088;
  wire v372eaaf;
  wire v3777191;
  wire v39ebb49;
  wire v374de7f;
  wire v3773ca9;
  wire v377395f;
  wire v372af91;
  wire v372f5e7;
  wire v3731e8c;
  wire v3a6fcc5;
  wire v376ca07;
  wire v3a6f95f;
  wire v3a6f342;
  wire v3a7006b;
  wire v3727482;
  wire v3722bc2;
  wire v372570c;
  wire v3a621ea;
  wire v3724368;
  wire v3a5b541;
  wire v375ab02;
  wire v3770c59;
  wire v3748f33;
  wire v376cdf6;
  wire v37311d8;
  wire v3a70d7f;
  wire v3731caa;
  wire v3779a60;
  wire v37627a2;
  wire v3a6f5c6;
  wire v37627a8;
  wire v3a5a75c;
  wire v376c8a4;
  wire v3729eb8;
  wire v37408a1;
  wire v3753f59;
  wire v3a70da8;
  wire v3a7109b;
  wire v3a6c42b;
  wire v373070b;
  wire v3a5ba95;
  wire v3a68f05;
  wire v3a6fd54;
  wire v377efe7;
  wire v3a5c860;
  wire v373c921;
  wire v375b239;
  wire v37377f0;
  wire v375bdd4;
  wire v3a6ebf1;
  wire v3a71617;
  wire v376a0e3;
  wire v3730526;
  wire v3a63559;
  wire v3a55f0d;
  wire v375a2a3;
  wire v37425ab;
  wire v3a63b69;
  wire v3a7079f;
  wire v3a5a801;
  wire v3744f35;
  wire v3a6f549;
  wire v375dbd4;
  wire v3744501;
  wire v3a6157d;
  wire v373c111;
  wire v374a0eb;
  wire v3736058;
  wire v3a6c8e4;
  wire v37542b2;
  wire v3a70ed0;
  wire v375dbb6;
  wire v376aa98;
  wire v3740951;
  wire v374d9c0;
  wire v3725948;
  wire v376aa57;
  wire v3776f5e;
  wire v372a96f;
  wire v3767ee9;
  wire v376e77e;
  wire v3758bbf;
  wire v3a62e3c;
  wire v373617a;
  wire v3748004;
  wire v377e04a;
  wire v3a6fc17;
  wire v3765b09;
  wire v3a5cebb;
  wire v375a5a1;
  wire v3749899;
  wire v3a70195;
  wire v3a6f032;
  wire v37722c4;
  wire v375b045;
  wire v377c6cf;
  wire v374bbc7;
  wire v3a5a6fb;
  wire v3763043;
  wire v37447b4;
  wire v3a6c43c;
  wire v3739768;
  wire v37414cd;
  wire v3726229;
  wire v372b819;
  wire v3a6b6f3;
  wire v375309f;
  wire v377d254;
  wire v3733278;
  wire v377b4c9;
  wire v3767985;
  wire v3726e48;
  wire v375a1fd;
  wire v37798ad;
  wire v3768c16;
  wire v374145d;
  wire v3755793;
  wire v3a64147;
  wire v37523ea;
  wire v3738a63;
  wire v376323b;
  wire v376ce1a;
  wire v376930a;
  wire v37760b8;
  wire v3730d52;
  wire v3759d98;
  wire v374d1b8;
  wire v376ce17;
  wire v375b9cc;
  wire v377432b;
  wire v376cd0a;
  wire v3a70e73;
  wire v377457e;
  wire v37291e4;
  wire v3a64252;
  wire v374f8b1;
  wire v374fa4c;
  wire v3a701c2;
  wire v374be32;
  wire v3a704ae;
  wire v3725036;
  wire v376ad33;
  wire v372760c;
  wire v3743b11;
  wire v3756531;
  wire v374ad24;
  wire v37298b9;
  wire v373c3ba;
  wire v375b019;
  wire v37290ab;
  wire v37250b5;
  wire v3a710cb;
  wire v3742b54;
  wire v373a158;
  wire v3757c5c;
  wire v375210d;
  wire v375ac12;
  wire v3a704d1;
  wire v3762720;
  wire v372b34d;
  wire v3a6aa8d;
  wire v3a700d0;
  wire v3a70abd;
  wire v3a54fb2;
  wire v3a65db0;
  wire v373e5f1;
  wire v3743bc5;
  wire v3a71519;
  wire v3a6f8df;
  wire v3a6f02c;
  wire v3a70f6a;
  wire v3737c2f;
  wire v377766c;
  wire v3a6f586;
  wire v376f569;
  wire v375754a;
  wire v375f0f8;
  wire v375586c;
  wire v3a6f3cf;
  wire v3779801;
  wire v3a6f707;
  wire v374abcc;
  wire v3a6f4ab;
  wire v3a5406b;
  wire v37536ae;
  wire v37334fc;
  wire v376a915;
  wire v3a5f622;
  wire v3767e76;
  wire v3a70bcd;
  wire v3756bde;
  wire v375455d;
  wire v3a6ff88;
  wire v3a5ead2;
  wire v3a6f776;
  wire v373513a;
  wire v3a62a9d;
  wire v3763eaa;
  wire v37618dc;
  wire v377606f;
  wire v3a6f522;
  wire v3a71102;
  wire v2acae91;
  wire v3a6ca53;
  wire v372437c;
  wire v374a8a5;
  wire v3731857;
  wire v3768995;
  wire v3a6469c;
  wire v373fda2;
  wire v3a5be20;
  wire v380a0c2;
  wire v3a7103a;
  wire v3777b2e;
  wire v374e8b4;
  wire v3774449;
  wire v375a4f8;
  wire v3751c54;
  wire v1e37c3e;
  wire v3723efc;
  wire v374fc8e;
  wire v37255d9;
  wire v3808f6f;
  wire v3756f10;
  wire v38071bb;
  wire v3a6d9a6;
  wire v3a5a5c8;
  wire v377b951;
  wire v3a708a1;
  wire v3748e82;
  wire v33790c9;
  wire v37415e4;
  wire v3752c04;
  wire v3727ce4;
  wire v3a69cd8;
  wire v3a694ec;
  wire v375eeb9;
  wire v3771303;
  wire v37467a3;
  wire v372ea9a;
  wire v376e794;
  wire v3a6f6b4;
  wire v3727d1e;
  wire v23fe376;
  wire v372f5bd;
  wire v375be12;
  wire v3a7012e;
  wire v3739c94;
  wire v3809f27;
  wire v37244f4;
  wire v3a5a05d;
  wire v376749b;
  wire v374637b;
  wire v377012f;
  wire v375a4b3;
  wire v37790ef;
  wire v3a7136e;
  wire v3a6d1aa;
  wire v37272ed;
  wire v3a6fdc3;
  wire v3a6b860;
  wire v3a554b9;
  wire v3a6f37f;
  wire v3a66ea9;
  wire v373a3c8;
  wire v3a670fb;
  wire v3a70aa2;
  wire v3751510;
  wire v3a5a28b;
  wire v3a68f16;
  wire v3a71077;
  wire v3764b0a;
  wire v373164a;
  wire v375f664;
  wire v374fad8;
  wire v3a7050e;
  wire v3755a96;
  wire v8d2bbf;
  wire v3732f54;
  wire v3a70936;
  wire v3772327;
  wire v3730d6b;
  wire v375931f;
  wire v3779ac0;
  wire v37639fa;
  wire v37416e1;
  wire v374a00a;
  wire v3733a1a;
  wire v373e8cb;
  wire v377da29;
  wire v372a7c1;
  wire v376dafa;
  wire v372998e;
  wire v3a663dd;
  wire v377181f;
  wire v3a70478;
  wire v3a66f40;
  wire v3768678;
  wire v3a5be8a;
  wire v373b9a9;
  wire v372c0f4;
  wire v374c4e9;
  wire v3a6fabe;
  wire d2dc90;
  wire v374cb97;
  wire v374b824;
  wire v3767cb7;
  wire v3a706e2;
  wire v3758a7b;
  wire v3758a4b;
  wire v3752397;
  wire v37316d9;
  wire v3a5334f;
  wire v3a6f374;
  wire v376c99e;
  wire v377624b;
  wire v377249b;
  wire v376d883;
  wire v35b91b6;
  wire v377bdd6;
  wire v2acae68;
  wire v374c9db;
  wire v375b9e1;
  wire v3764eb2;
  wire v373d2bd;
  wire v3a5a39f;
  wire v3751c8c;
  wire v3a60340;
  wire v3747358;
  wire v37590f4;
  wire v376c5de;
  wire v37261be;
  wire v92c996;
  wire v3a68bdb;
  wire v3a55d78;
  wire v3773712;
  wire v3730f7e;
  wire v377a62e;
  wire v3a574fc;
  wire v3a5b93f;
  wire v373b785;
  wire c39ea5;
  wire v3a65c47;
  wire v374a516;
  wire v39eb1dc;
  wire v3736cd2;
  wire v3764fd5;
  wire v377814d;
  wire v3773661;
  wire v2093068;
  wire v3750295;
  wire v3a6850e;
  wire v3a70cc6;
  wire v374e5eb;
  wire v3a5946d;
  wire v3a6c363;
  wire v3a6cac4;
  wire v3a6c0ab;
  wire v374f9cc;
  wire v37565d3;
  wire v3a709c2;
  wire v372a478;
  wire v3a6b368;
  wire v37361ad;
  wire v8455d1;
  wire v866387;
  wire v8455cd;
  wire v373b287;
  wire v374fa66;
  wire v37702e6;
  wire v375ff1e;
  wire v375e147;
  wire v3751fde;
  wire v35772a5;
  wire v3731d80;
  wire v3a635ea;
  wire v3577306;
  wire v3a6f210;
  wire v35772a6;
  wire v3a6ffae;
  wire v374306c;
  wire v3752b8c;
  wire v865472;
  wire v3728b28;
  wire v35772b3;
  wire v3a5b5d3;
  wire c118e3;
  wire v377975f;
  wire v3734ed6;
  wire v372ccea;
  wire v373e80b;
  wire v3806a74;
  wire v3a658bf;
  wire v374d95a;
  wire v373cd5a;
  wire v375e3fd;
  wire v373c590;
  wire v3739077;
  wire v37350e9;
  wire v3722e5c;
  wire v3a6eb39;
  wire v37582dc;
  wire v3a624da;
  wire v37604e9;
  wire v3764683;
  wire v3775651;
  wire v3770559;
  wire v376df25;
  wire v375ce98;
  wire v372be9b;
  wire v372abd8;
  wire v3774a9c;
  wire v373d5df;
  wire v375da9f;
  wire v374f52f;
  wire v3762145;
  wire v3a713b4;
  wire v374e8c3;
  wire v3762858;
  wire v3778372;
  wire v3a6ec83;
  wire v3a70498;
  wire v37499a4;
  wire v3a68af5;
  wire v3766830;
  wire v3753198;
  wire v376c3c2;
  wire v3748c4c;
  wire v3a6db2d;
  wire v377de29;
  wire v3740a8a;
  wire v376c047;
  wire v3776abb;
  wire v3a70652;
  wire v3a69f2b;
  wire v3a6ece9;
  wire v375b5d3;
  wire v3a70c85;
  wire v3755066;
  wire v374d669;
  wire v377a5cc;
  wire v37470a5;
  wire v3765962;
  wire v3746b7f;
  wire v3a58017;
  wire v3761da5;
  wire v373bdd1;
  wire v3a678de;
  wire v3761916;
  wire v3748da1;
  wire v3756723;
  wire v374bb74;
  wire v3725be8;
  wire v375e1f6;
  wire v3a6feb8;
  wire v374d6de;
  wire v3751ebd;
  wire v37246b5;
  wire v3a70769;
  wire v3a69584;
  wire v3751389;
  wire v8c8903;
  wire v372ffaa;
  wire v37400f8;
  wire v37320bb;
  wire v375db2a;
  wire v372f657;
  wire v3753e6a;
  wire v3a626a1;
  wire v3a6af99;
  wire v3a54427;
  wire v3729480;
  wire v3724b72;
  wire v377b24b;
  wire v3751fa8;
  wire v37286bb;
  wire v3a610e9;
  wire v374fef8;
  wire v37397c3;
  wire v37655d6;
  wire v3a5561b;
  wire v3772e33;
  wire v3768e70;
  wire v3a5fabd;
  wire v37617ef;
  wire v3727b03;
  wire v3a6f4b2;
  wire v3a5c90c;
  wire v3750b04;
  wire v373df0d;
  wire v37665ea;
  wire v3741669;
  wire v373b414;
  wire v3a71571;
  wire v3a6fd6f;
  wire v3737462;
  wire v3a70c38;
  wire v373a181;
  wire v3a70e6f;
  wire v3a5794d;
  wire v3a5f6d5;
  wire v3763b94;
  wire v37612c1;
  wire v3a5b687;
  wire v372bb25;
  wire v3a64931;
  wire v1e379fa;
  wire v3744f6f;
  wire v3766df8;
  wire v3a6f4e3;
  wire v37482da;
  wire v3a704a7;
  wire v3a5a225;
  wire v380775e;
  wire v372dab1;
  wire v372e5d3;
  wire v3a70c66;
  wire v37341bc;
  wire v3a70295;
  wire v3738de9;
  wire v3a70547;
  wire v3a6fff6;
  wire v3a5d0b6;
  wire v3a62654;
  wire v37413d5;
  wire v375bc38;
  wire v3a66ac0;
  wire v372b02f;
  wire v374e079;
  wire v3739fb8;
  wire v3777ee7;
  wire v3775e7e;
  wire v3731684;
  wire v3a713d1;
  wire v3a575a5;
  wire v37494da;
  wire v375fbe1;
  wire v3738aef;
  wire v3a65088;
  wire v3749ba6;
  wire v37565c3;
  wire v372ab0f;
  wire v3a5f2bd;
  wire v375a311;
  wire v3736df1;
  wire v377057c;
  wire v377d01e;
  wire v3a6f9bc;
  wire v374f511;
  wire v3379035;
  wire v37598dc;
  wire v3a682cb;
  wire v3776c43;
  wire v37293b1;
  wire v37566a2;
  wire v3726098;
  wire v372f62a;
  wire v3a64ded;
  wire v3a6fb37;
  wire be0bbd;
  wire v3a6f32d;
  wire v38092b4;
  wire v374eef1;
  wire v3764218;
  wire v3a6aefd;
  wire v374f3a3;
  wire v3a7012f;
  wire v3a6a22c;
  wire v372a347;
  wire v374cb44;
  wire v3a62628;
  wire v3a54108;
  wire v375e7d6;
  wire v3737c6c;
  wire v3a6fd34;
  wire v3a7082d;
  wire v377fad8;
  wire v3a5e0b8;
  wire v3a5c7a8;
  wire v3754b58;
  wire v376aa5e;
  wire v3766b5e;
  wire v372ac3a;
  wire v3a6fbe2;
  wire v376d5a4;
  wire v37506fb;
  wire v3779ea0;
  wire cc9d04;
  wire v376b97b;
  wire v372d593;
  wire v3754c0e;
  wire v377aad8;
  wire v374d4c1;
  wire v3747dfc;
  wire v377a6f2;
  wire v3a625d8;
  wire v3a62a08;
  wire v375d70e;
  wire v373512b;
  wire v3733170;
  wire v374a580;
  wire v376a3fe;
  wire v3a630db;
  wire v3751d73;
  wire v3778b51;
  wire v3755e4e;
  wire v3a6fb2a;
  wire v38095ed;
  wire v3745b4f;
  wire v9f7a48;
  wire v3a713fb;
  wire v3a5d34b;
  wire v360d0a7;
  wire v3751d87;
  wire v37424b5;
  wire v372ad52;
  wire v3a7105c;
  wire v3a563af;
  wire v3774d9a;
  wire v3a6fdb7;
  wire v3744e13;
  wire v375d94c;
  wire v3727187;
  wire v3a6fb4b;
  wire v377b920;
  wire v3739120;
  wire v3a70225;
  wire v373f260;
  wire v9d35e2;
  wire v3a708ee;
  wire v3a5dd10;
  wire v3a66373;
  wire v3769fa2;
  wire v3728085;
  wire v3a704b7;
  wire v375cf46;
  wire v3a6b001;
  wire v3730097;
  wire v37432e1;
  wire v3763f05;
  wire v3775c03;
  wire v377410f;
  wire v3779fbc;
  wire v8bc1c0;
  wire v377cf4f;
  wire v3778ae9;
  wire v3755ab8;
  wire v3753386;
  wire v3768add;
  wire v3746a04;
  wire v375987b;
  wire v372be8e;
  wire v374b27d;
  wire v3761b5e;
  wire v373523c;
  wire v3770331;
  wire v3730145;
  wire v3a5b98b;
  wire v3a5445e;
  wire v3a6a87d;
  wire v3761497;
  wire v3a6fd86;
  wire v37533e3;
  wire v3778b8c;
  wire v372a3de;
  wire v3a5dfad;
  wire v3777bd6;
  wire v377e9a4;
  wire v3a701d7;
  wire v3732931;
  wire v3762c7c;
  wire v3a5b9ba;
  wire v3a642cf;
  wire v9e8a9c;
  wire v372468b;
  wire v3733467;
  wire v375898f;
  wire v3760951;
  wire v376c4ba;
  wire v3728646;
  wire v375b2af;
  wire c2e325;
  wire v3a5cfbb;
  wire v3752781;
  wire v3a650e9;
  wire v376634c;
  wire v37572b6;
  wire v3a70b43;
  wire b8ed55;
  wire v3a62e7b;
  wire v3a69feb;
  wire v38096d8;
  wire v376662b;
  wire v39a4ce0;
  wire v3a700ab;
  wire v377541e;
  wire v37632c6;
  wire v3a5857e;
  wire v377c29b;
  wire v373e2bc;
  wire v374f535;
  wire v3a6f834;
  wire v3722a42;
  wire v3a71125;
  wire v3a56194;
  wire v372d8bd;
  wire v3726277;
  wire v3770d70;
  wire v374db93;
  wire v37614c8;
  wire v375416d;
  wire v374189f;
  wire v37297f4;
  wire v3a7066c;
  wire v372865e;
  wire v372eb43;
  wire v37682a8;
  wire v9d7b97;
  wire v3738d68;
  wire v3767420;
  wire v37259c7;
  wire v37793a4;
  wire v3a5c16e;
  wire v374764e;
  wire v3733d66;
  wire v374c98c;
  wire v3a71340;
  wire v3a54dd4;
  wire v3256555;
  wire v3745e12;
  wire v3a71009;
  wire v373539e;
  wire v376a77a;
  wire v37345f3;
  wire v37483db;
  wire v3735179;
  wire v9ec00e;
  wire v377bb6d;
  wire b62443;
  wire v376fafe;
  wire v3a712b2;
  wire v3737478;
  wire v3a6f842;
  wire v376a822;
  wire v3a680e3;
  wire v376a1dd;
  wire v3a5f76b;
  wire v375dff6;
  wire v3762453;
  wire v375a7bd;
  wire c1a4f5;
  wire v3775abc;
  wire v38063c7;
  wire v3757a13;
  wire v374da36;
  wire v375a697;
  wire v372379e;
  wire v3a5ef3e;
  wire v374c74f;
  wire v3764f8a;
  wire v3a2a2fa;
  wire v376d251;
  wire v3761678;
  wire v3778173;
  wire v3a6f31c;
  wire v372628c;
  wire v3729173;
  wire v375d00d;
  wire v375bacc;
  wire v37462ae;
  wire v376b2f4;
  wire v376b0cc;
  wire v3771533;
  wire v3740ed1;
  wire v3a6fa35;
  wire v3745bee;
  wire v3a573bb;
  wire v3a5c842;
  wire v37386d3;
  wire v373ea50;
  wire v373cc0c;
  wire v373917f;
  wire v376f261;
  wire v373b0f5;
  wire v3767010;
  wire v3760ce0;
  wire v380886b;
  wire v376b03d;
  wire v3a5a2d4;
  wire v3779d09;
  wire v377b6ce;
  wire v3a6fee4;
  wire v3a597d8;
  wire v3a70b5c;
  wire v3a56804;
  wire v377d206;
  wire v3a700a6;
  wire v3774dcd;
  wire v3a5e2fa;
  wire v37750bb;
  wire v3a7159b;
  wire v3a6fd70;
  wire v377d223;
  wire v375811b;
  wire v3758fae;
  wire v372fc51;
  wire v37393f0;
  wire v373217b;
  wire v3740152;
  wire v3747cdb;
  wire ab60dc;
  wire ce419c;
  wire v3a71599;
  wire v3a5a24b;
  wire v377217f;
  wire v37761e4;
  wire v374790d;
  wire v3769157;
  wire v373f4a5;
  wire v3a6c835;
  wire v3a5f3e3;
  wire v2ff8cfd;
  wire v1e37b47;
  wire v372873a;
  wire v37684e6;
  wire v37515e1;
  wire v3769f60;
  wire v3a6437e;
  wire v3a5c2f4;
  wire v377184d;
  wire v372562b;
  wire v3739c14;
  wire v3746905;
  wire v3757727;
  wire v376618c;
  wire v3a71354;
  wire v3759a00;
  wire v3731142;
  wire v3a555b3;
  wire v3a5d327;
  wire v372b445;
  wire v375e232;
  wire v377e158;
  wire v373b600;
  wire v3754b35;
  wire v3753883;
  wire v3a70049;
  wire v373e85a;
  wire v373ff58;
  wire v35b7189;
  wire v37229b8;
  wire v2092eb7;
  wire c04cff;
  wire v3748b0e;
  wire v375d2ee;
  wire v3a70455;
  wire v374c63d;
  wire v3774629;
  wire v374d6b5;
  wire v3a585f5;
  wire v3a68e41;
  wire v3765ded;
  wire v373e02a;
  wire v3a6086a;
  wire v357748a;
  wire v3778ed4;
  wire v3a71635;
  wire v37231c2;
  wire v376c477;
  wire v3a620fd;
  wire v3a6ebda;
  wire v376079e;
  wire v376f49f;
  wire v374d383;
  wire v3a66c34;
  wire v374fddd;
  wire v3739ddd;
  wire v373ee8b;
  wire v3a6e66e;
  wire v3a6eafc;
  wire v377217c;
  wire v3a70dc0;
  wire v37273be;
  wire v37535bd;
  wire v3a6b3d4;
  wire v3735324;
  wire v3a6fbaa;
  wire v372d75d;
  wire v376cdc4;
  wire v3a575d5;
  wire v3a6d8ce;
  wire v3a70b72;
  wire v3a59883;
  wire v37595c8;
  wire v37664ab;
  wire v376fa76;
  wire v377df60;
  wire v3728cd0;
  wire v37240e6;
  wire v3765f60;
  wire v3762d6e;
  wire v373b11a;
  wire v3a697b9;
  wire v3a53986;
  wire v373ea8d;
  wire v375cfe0;
  wire v3726448;
  wire v375bc6f;
  wire v3742de5;
  wire v3a6ef19;
  wire v3a672de;
  wire v3a705a2;
  wire v3773f85;
  wire v3a5a6db;
  wire v3a55aba;
  wire v373c853;
  wire v37532a6;
  wire v3741ef3;
  wire v375f7d1;
  wire v3a6ad22;
  wire v372defe;
  wire v3a5fb15;
  wire v3a634c9;
  wire v3a66d43;
  wire v3739b40;
  wire v3a710f9;
  wire v3755a2f;
  wire v3a7133b;
  wire v37229f0;
  wire v3a54c8b;
  wire v3730a34;
  wire v3766448;
  wire v3768095;
  wire v3a64dbd;
  wire v372da87;
  wire v3737ce6;
  wire v3757651;
  wire v3750b0d;
  wire v377a9a1;
  wire v37617ed;
  wire v376107b;
  wire v3739791;
  wire v377bdc3;
  wire v3749c27;
  wire v1e3757b;
  wire v3751905;
  wire v3a621be;
  wire v372cfbf;
  wire v372c571;
  wire v373bf1d;
  wire v3734caf;
  wire v3a7087c;
  wire v3a6e2ec;
  wire v372b5ed;
  wire v37673a3;
  wire v3742584;
  wire v373ff8d;
  wire v3745d3f;
  wire v374d998;
  wire v373d10a;
  wire v3a71409;
  wire v376bb9f;
  wire v373f200;
  wire v372eff2;
  wire v374c582;
  wire v3a713dd;
  wire v3a53dbb;
  wire v3809399;
  wire v3a6f8cc;
  wire v3768889;
  wire v37559ec;
  wire v37388aa;
  wire v3a6db4b;
  wire v374e4c9;
  wire v37398f3;
  wire v37257f8;
  wire v376e677;
  wire v3a70178;
  wire v375bb15;
  wire v3a5b5ef;
  wire v3a703fa;
  wire v3759ad8;
  wire v3a65532;
  wire v3774346;
  wire v3a6f151;
  wire v37749c3;
  wire v37512c0;
  wire v3a703be;
  wire v3753976;
  wire v376eb57;
  wire v3737e97;
  wire v3763f3f;
  wire v3a5fc64;
  wire v3a70c21;
  wire v372a7c2;
  wire v288971d;
  wire v3a71084;
  wire v3a619c0;
  wire v3a5c945;
  wire v3a66110;
  wire v3a57f59;
  wire v376bd2c;
  wire v3a5bd24;
  wire v3735e39;
  wire v3a6cfc5;
  wire v37297c0;
  wire v360d1cd;
  wire v3766d53;
  wire v374016f;
  wire v37458a2;
  wire v3751e0a;
  wire v376d856;
  wire v3724c9c;
  wire v3a6eaba;
  wire v3725d79;
  wire v3a6f54e;
  wire v373f6f0;
  wire v374f36b;
  wire v3766664;
  wire v3a5bf04;
  wire v3a57867;
  wire v3737bfb;
  wire v377f505;
  wire v374fb02;
  wire v3734c3a;
  wire v3a6f9b6;
  wire v3a70605;
  wire v3a6f443;
  wire v3747816;
  wire v3a6d140;
  wire v37737d2;
  wire v3a58cfc;
  wire v3a5b545;
  wire v374f52a;
  wire v3a582bc;
  wire v3751849;
  wire v373cd8f;
  wire v3a56d30;
  wire v376dd7a;
  wire v3a70c31;
  wire v3772c4d;
  wire v3759032;
  wire v3733e9e;
  wire v37432c6;
  wire v3736104;
  wire v376d285;
  wire v3758166;
  wire v3a61c70;
  wire v3a6ff31;
  wire v376ea4a;
  wire v3732eb2;
  wire v3a53a94;
  wire v372d943;
  wire v3a70272;
  wire v3a658cf;
  wire v37589e1;
  wire v3a6f04e;
  wire v3758b05;
  wire v3a5744d;
  wire v3a69da8;
  wire v37521ed;
  wire v376f70a;
  wire v372c007;
  wire v3a56e63;
  wire v3a56512;
  wire v360d0c7;
  wire v3728e09;
  wire v3767f36;
  wire v3744981;
  wire v3a7011c;
  wire v3a5b68a;
  wire v373a246;
  wire v37365fa;
  wire v3a5408e;
  wire v372b91e;
  wire v376a3f5;
  wire v3a69ec5;
  wire v377bac7;
  wire v3725392;
  wire v373a2f4;
  wire v372eb0f;
  wire v3745714;
  wire v375345f;
  wire v3a70333;
  wire v3a5fcf0;
  wire v3726638;
  wire v3a698e1;
  wire v2ff8e61;
  wire v3a709de;
  wire v3a5a510;
  wire v375f95f;
  wire v3a69028;
  wire v3a71386;
  wire v1e382e7;
  wire v376fce9;
  wire v3a70e25;
  wire v3a70b4f;
  wire v373b90b;
  wire v3764d6b;
  wire v3746ab7;
  wire v37590d5;
  wire v3a656f0;
  wire v3751094;
  wire v3807bf8;
  wire v3a68c1f;
  wire v3a6f92f;
  wire v37502b7;
  wire v39a4dbb;
  wire v3a6f3f5;
  wire v3730c14;
  wire v3a56a0d;
  wire v377adf5;
  wire v376f9a8;
  wire v3736847;
  wire v37635f0;
  wire v3a70eac;
  wire v3774369;
  wire v3a69427;
  wire v3a70c07;
  wire v376d45f;
  wire v3a56cdb;
  wire v37234d1;
  wire v374b879;
  wire v3758ab3;
  wire v3775120;
  wire v3a5a52f;
  wire v3a5891c;
  wire v3768c3c;
  wire v376ef42;
  wire v3a707cd;
  wire v3a5fdd3;
  wire v3a5ade4;
  wire v3a70326;
  wire v3725c63;
  wire v37654c4;
  wire v37702f3;
  wire v376f73c;
  wire v3748609;
  wire v3777467;
  wire v3a7093c;
  wire v3a66d1b;
  wire v3a71528;
  wire v377a9e7;
  wire v3747dd8;
  wire v376cdb7;
  wire v3758f2e;
  wire v37775ce;
  wire v377b8fb;
  wire v3a57eae;
  wire v374c7f4;
  wire v37662dc;
  wire v3a627cc;
  wire v376d550;
  wire v3766bc8;
  wire v38074c2;
  wire v377e004;
  wire v377439e;
  wire v3732e1b;
  wire v3732569;
  wire v37237e8;
  wire v374734d;
  wire v3730343;
  wire v3a71065;
  wire v3747623;
  wire v376ff85;
  wire v37509f2;
  wire v3a6f7c5;
  wire v37796c3;
  wire v3a67e97;
  wire v3a59a60;
  wire v373a1a4;
  wire v377bb57;
  wire v373bbd0;
  wire v376cff4;
  wire v376f5d9;
  wire v3a5e000;
  wire v3747141;
  wire v377a0a1;
  wire v3735fc8;
  wire v3744202;
  wire v3774d13;
  wire v3a70931;
  wire v3761930;
  wire v3a7102a;
  wire c60fa0;
  wire v374d525;
  wire v3760e51;
  wire v3a60836;
  wire v372348f;
  wire v3742dcb;
  wire v377224f;
  wire v3a6fde5;
  wire v3a6f82c;
  wire v3a6f6a8;
  wire v3a6fbaf;
  wire v3726ed7;
  wire v3738b7e;
  wire v3808c89;
  wire v3a703db;
  wire v3730a73;
  wire v372ced7;
  wire v3760e6e;
  wire v3a70071;
  wire v3747465;
  wire v3a70d3a;
  wire v376eed1;
  wire v3a6750f;
  wire v376bc8c;
  wire v3735859;
  wire v3a7068f;
  wire v3a6fd8a;
  wire v37475be;
  wire v372779c;
  wire v376eaf2;
  wire v3773eee;
  wire v377d91c;
  wire v372d149;
  wire v3745a3b;
  wire v3a6eb09;
  wire v3a6f938;
  wire v3744990;
  wire v3a6ad0b;
  wire v3a6b285;
  wire v374f0f1;
  wire v377bcf5;
  wire v3a706c5;
  wire v377478a;
  wire v376fed4;
  wire v3726d0c;
  wire v372de54;
  wire v372d780;
  wire v373a222;
  wire v37357d9;
  wire v374237b;
  wire v3a6f463;
  wire v3778cba;
  wire v3777c7f;
  wire v3761702;
  wire v3a70ca1;
  wire v3a65287;
  wire v3736b3b;
  wire v3759d9c;
  wire v37576ec;
  wire v374b13e;
  wire v374cceb;
  wire v37751bb;
  wire v3754bd4;
  wire v373644e;
  wire v3736d1d;
  wire v3768f71;
  wire v3a65b00;
  wire v373d593;
  wire v3a5ada9;
  wire v3734579;
  wire v3a6d33e;
  wire v3a7115d;
  wire v373580c;
  wire v374727f;
  wire v3a70254;
  wire v373b6dd;
  wire v376f6e4;
  wire v3779883;
  wire v375d46e;
  wire v3a5e1e8;
  wire v37443a2;
  wire v374a37e;
  wire v3756a8f;
  wire v3a65ce5;
  wire v99aa13;
  wire v3a5a1e8;
  wire v380651a;
  wire v373739c;
  wire v3a6fb9b;
  wire v3742360;
  wire v3a6799a;
  wire v375c7c4;
  wire v3727a6b;
  wire v3a649da;
  wire v3a5711b;
  wire v3a694b9;
  wire v3a60026;
  wire v377d596;
  wire v3a7010b;
  wire v3a712a5;
  wire v373a7f7;
  wire v3a6d768;
  wire c03a6a;
  wire v372c335;
  wire v3a6f223;
  wire v3746f18;
  wire v35b7768;
  wire v3a6eaf7;
  wire v3777a8a;
  wire v3726594;
  wire v375d387;
  wire v375e039;
  wire v373cae5;
  wire v3a6fc4a;
  wire v3a58604;
  wire v373ff91;
  wire v377618a;
  wire v3a2a348;
  wire v3754e5a;
  wire v3a70233;
  wire v1e38275;
  wire v3a5e24e;
  wire v376ba47;
  wire v38071c1;
  wire v375cec6;
  wire v373dc2f;
  wire v376a8cf;
  wire v375d7b6;
  wire v3764a16;
  wire v3806e0e;
  wire v3764702;
  wire v3a5c3a0;
  wire v3a6fac2;
  wire v3a645b0;
  wire v3746dd5;
  wire v3770f46;
  wire v3735f56;
  wire v3a70ecf;
  wire v3a64566;
  wire v3a6eb77;
  wire v373e16a;
  wire v3a670a1;
  wire v375825a;
  wire v37705d1;
  wire v3a6a1fd;
  wire v37310be;
  wire v373e474;
  wire v377c15d;
  wire v3732b35;
  wire v3a705bf;
  wire v3740110;
  wire v37434d6;
  wire v375d690;
  wire v3766452;
  wire v377b673;
  wire v3a5d356;
  wire v3a5cc4c;
  wire v37610f8;
  wire v3731f7a;
  wire v375a1ab;
  wire v376d93b;
  wire v376824b;
  wire v3a6497b;
  wire v3778333;
  wire v372b077;
  wire v373c074;
  wire v3776d62;
  wire v375e93c;
  wire v375b6c3;
  wire v3779931;
  wire v376139f;
  wire v3731d75;
  wire v3a5c5fc;
  wire v3725475;
  wire v376e7bc;
  wire v37487ca;
  wire v3770b89;
  wire b27f78;
  wire v374e03d;
  wire v37780f6;
  wire v3808eaa;
  wire v3724fe7;
  wire v37745c3;
  wire v373e5d9;
  wire v3a707e0;
  wire v372e33d;
  wire v3a61a2d;
  wire v372ce29;
  wire v3747210;
  wire v3741759;
  wire v377adc8;
  wire v3a6fc6e;
  wire v374c9c7;
  wire v375bbe9;
  wire v3a5fe1d;
  wire v3a53cc3;
  wire v3744265;
  wire v3772dd1;
  wire v3a7094a;
  wire v37504b9;
  wire d08a74;
  wire v3a709aa;
  wire v3759d5a;
  wire v373c95b;
  wire v375c90b;
  wire v3a66f07;
  wire v3746ab1;
  wire v375607f;
  wire v3758dcb;
  wire v37696c4;
  wire v3a715d9;
  wire v3a6096a;
  wire v3a70d19;
  wire v3a71214;
  wire v3778032;
  wire v3739808;
  wire v377a92d;
  wire v3740f7e;
  wire v3a6a758;
  wire v374e21d;
  wire v3a624ec;
  wire v3a5ceaf;
  wire v3758fc4;
  wire v37350b7;
  wire v377c6d0;
  wire v3a6b60d;
  wire v39eb431;
  wire v376b8c2;
  wire v3771ad8;
  wire v374d726;
  wire v377c49c;
  wire v3a6e005;
  wire v3a650a7;
  wire v377dc72;
  wire v3761c72;
  wire v3774b16;
  wire v3766ed8;
  wire v376d872;
  wire v3a6783b;
  wire v3762929;
  wire v37510e5;
  wire v3723e15;
  wire v39eb520;
  wire v3a70eb0;
  wire v37540e2;
  wire v375ddaf;
  wire v3a709d5;
  wire v3727194;
  wire v3a6bfb5;
  wire v376c7cc;
  wire v3a6fbbd;
  wire v3773336;
  wire v373cedd;
  wire v3a6d9da;
  wire v37539cd;
  wire v37742a4;
  wire v37653ef;
  wire v37548f4;
  wire v3a6491d;
  wire v375eb79;
  wire v373557e;
  wire v3769ed3;
  wire v3a6ebe6;
  wire v37745e0;
  wire v37283a8;
  wire v3725b4f;
  wire v3731b11;
  wire v3a712e3;
  wire v3a6212b;
  wire v37265b8;
  wire v2ff937f;
  wire v3a664b5;
  wire v3777d29;
  wire v376b600;
  wire v376a88b;
  wire v374c801;
  wire v3a5c0ac;
  wire v3a6d21e;
  wire v373ade9;
  wire v3763ff7;
  wire v373de66;
  wire v376defa;
  wire v38068b5;
  wire v3730e5d;
  wire v3768a37;
  wire v2ff8cae;
  wire v375b0e4;
  wire v376aa54;
  wire v37747db;
  wire v377e469;
  wire v3753f17;
  wire v372dcd4;
  wire v3a5880b;
  wire v3a70011;
  wire v3779709;
  wire v3a5ddd4;
  wire v3732e39;
  wire v3a6918e;
  wire v3a684ef;
  wire v3a53f45;
  wire v3741e2a;
  wire v3736ea1;
  wire v372d2dc;
  wire v3729178;
  wire v3a6fc8f;
  wire v3741b92;
  wire v377d821;
  wire v374c107;
  wire v375413c;
  wire v9cc76d;
  wire v376cf8c;
  wire v37712f6;
  wire v374abf3;
  wire v3a70e93;
  wire v376a6d6;
  wire v373e5ad;
  wire v376c2e2;
  wire v37240e8;
  wire v3735a4f;
  wire v88c50b;
  wire v373c07d;
  wire v3764585;
  wire v372e544;
  wire v376eb33;
  wire v374aa1b;
  wire v3a6fcbe;
  wire v3a6f6ca;
  wire v372dc2b;
  wire v3a5b25f;
  wire v373dd3c;
  wire v3a68cb5;
  wire v374a35d;
  wire v3734bd2;
  wire v3754c02;
  wire v3a6973f;
  wire v3a6a64f;
  wire v3750e8a;
  wire v375d41f;
  wire v373e163;
  wire v375e0cb;
  wire v3a547ff;
  wire d1375e;
  wire v3378992;
  wire v3a640fd;
  wire v3a67dd8;
  wire v3758aec;
  wire v37483dd;
  wire v3a6ae68;
  wire v377abd1;
  wire v37402f0;
  wire v380761c;
  wire v3a70d7a;
  wire v374b32b;
  wire v37795d3;
  wire v375ff4e;
  wire v374177d;
  wire v374b199;
  wire v3a7156c;
  wire v3773acc;
  wire v37374d6;
  wire v374925f;
  wire v377d146;
  wire v3a6fd45;
  wire v2093037;
  wire v3a6f3f8;
  wire v375dd84;
  wire v372538e;
  wire v3a71547;
  wire v3772e0a;
  wire v374ebd1;
  wire v3762525;
  wire v3a701e9;
  wire v3a57db8;
  wire v3777b00;
  wire v3757dee;
  wire v3a70f41;
  wire v372601c;
  wire v3759ac1;
  wire v374072b;
  wire v3a70831;
  wire v3a708f8;
  wire v3755b55;
  wire v3a6572c;
  wire v3746d31;
  wire v3809f73;
  wire v373a692;
  wire v3738d19;
  wire v377936c;
  wire v3a6f8e7;
  wire v3a6ffea;
  wire v3773044;
  wire v377cbad;
  wire v376e500;
  wire v375dab1;
  wire v372c11d;
  wire v3a70c73;
  wire v373918a;
  wire v9dc858;
  wire v3770993;
  wire v373c79c;
  wire v3765901;
  wire v37798aa;
  wire v3a5ce1e;
  wire v3a70c9b;
  wire v3a566eb;
  wire v37497dd;
  wire v3775234;
  wire v35b8d36;
  wire v3a6efc6;
  wire v376c03e;
  wire v3a5c5ae;
  wire a38ed7;
  wire v3a6123a;
  wire v3725a06;
  wire v3759fe0;
  wire v3a6ef49;
  wire v37539fc;
  wire v3a70464;
  wire v375043c;
  wire d6db19;
  wire v3a5bcc4;
  wire v374bdfb;
  wire v373c379;
  wire v3761671;
  wire v3a682f9;
  wire v37575fd;
  wire v3a5bccf;
  wire v374ca88;
  wire v3744b27;
  wire v373e37c;
  wire v373cf42;
  wire v1e37d3f;
  wire v37775c4;
  wire v37707eb;
  wire v3772020;
  wire v38076a8;
  wire v375b34f;
  wire v3a60d86;
  wire v375bfdf;
  wire v3a71207;
  wire v37555b4;
  wire v377da41;
  wire v3a6fe1c;
  wire v377e1e8;
  wire v374765b;
  wire v3a70ce6;
  wire v37740ec;
  wire v374ad44;
  wire v372647d;
  wire v373695f;
  wire v374bd2c;
  wire v372de6f;
  wire v3a56323;
  wire v380776b;
  wire v3a70dba;
  wire v3756cea;
  wire v37301f9;
  wire v37474fc;
  wire v37394b7;
  wire v3a6692b;
  wire v3729d0b;
  wire v375c1c5;
  wire v376fd33;
  wire v376f53e;
  wire v37767d7;
  wire v3a63def;
  wire v3752e42;
  wire v376ea13;
  wire v375c0f1;
  wire v3a70e38;
  wire v3769630;
  wire v3807003;
  wire v38072f4;
  wire v3a7150d;
  wire v372e48a;
  wire v3a70eec;
  wire v3745149;
  wire v373ed95;
  wire v37450ff;
  wire v375e6ed;
  wire v377a356;
  wire v374b759;
  wire v3a6425d;
  wire v3a7063c;
  wire v375fac6;
  wire v3760b7a;
  wire v8fc6a0;
  wire v3740187;
  wire v3766d24;
  wire v372d249;
  wire v3738636;
  wire v3a68fc9;
  wire v3731b33;
  wire v39a4e12;
  wire v375f3f0;
  wire v37732c0;
  wire v3a6ebff;
  wire v3a70593;
  wire v3760582;
  wire v3771728;
  wire v374fad3;
  wire v373b8ff;
  wire v377b983;
  wire v373d338;
  wire v372367c;
  wire v374b5c5;
  wire v3a7097c;
  wire v373ec24;
  wire v3762924;
  wire v3752e1b;
  wire v3a61bfd;
  wire v373f159;
  wire v3739761;
  wire v377f812;
  wire v377f76a;
  wire v3732c52;
  wire v376866e;
  wire v374b3e1;
  wire v373b0e5;
  wire v2092f20;
  wire v3746888;
  wire v3776415;
  wire v372ac03;
  wire v37266c6;
  wire v3744c10;
  wire v3733cd1;
  wire v96f7ab;
  wire c0c2de;
  wire v3727d18;
  wire v3a70601;
  wire v375a79d;
  wire v3723780;
  wire v37404c5;
  wire v3a6f051;
  wire v3a67b62;
  wire v372f4ce;
  wire v3765cec;
  wire v375ce8d;
  wire v3762640;
  wire v376ffa7;
  wire v3755596;
  wire v375e7bb;
  wire v3a6f8a2;
  wire v374bdcb;
  wire v3a5b6c8;
  wire v3741b5a;
  wire v3a6f7b8;
  wire v372428a;
  wire v375f2ab;
  wire v374b8fe;
  wire v372d360;
  wire v23fe142;
  wire v3777474;
  wire v3735aa5;
  wire v376ae39;
  wire v372e1bc;
  wire v3a70428;
  wire v3768d8f;
  wire v3a5e2af;
  wire v3a6e31f;
  wire v37565af;
  wire v3753927;
  wire v3769712;
  wire v3a5af94;
  wire v37441fb;
  wire v3808531;
  wire v3749a7c;
  wire v372d6fa;
  wire v3728045;
  wire v37232a3;
  wire v372ac64;
  wire v3a6f973;
  wire v3378b65;
  wire v3746e54;
  wire v372969d;
  wire v3779060;
  wire v372391f;
  wire v3a706f8;
  wire v3a58640;
  wire v373afa4;
  wire v3a6dfb2;
  wire v375e60f;
  wire v37559b4;
  wire v37270ad;
  wire v37519dd;
  wire v377b233;
  wire v3a672c9;
  wire v3a63989;
  wire v376980f;
  wire v374fcfe;
  wire v37609c3;
  wire v3a66593;
  wire v3734967;
  wire v3754b6c;
  wire v37625a8;
  wire v377613b;
  wire v3725ceb;
  wire v3750ac3;
  wire v3a5e357;
  wire v374729b;
  wire v3a6eb66;
  wire v3a5ace5;
  wire v3a6f0c8;
  wire v3761c19;
  wire v3a5a23b;
  wire v3a6eac2;
  wire v96020f;
  wire v3725f77;
  wire v3a5c3d7;
  wire v3a64b57;
  wire v3a695c1;
  wire v3753af9;
  wire v376b1aa;
  wire v3759b2f;
  wire v3a6f43e;
  wire v375641f;
  wire v3a68c94;
  wire v37632f8;
  wire v3734067;
  wire v3a6cf7f;
  wire v37249c7;
  wire v3772b14;
  wire v3a5ee73;
  wire v3a706b0;
  wire v3774c1b;
  wire v37243fe;
  wire v3a55904;
  wire v3727d7e;
  wire v3752977;
  wire v3a70516;
  wire v3733e5a;
  wire v373be25;
  wire v372935c;
  wire v3a6b0c7;
  wire v3a712c8;
  wire v3737860;
  wire v3a68b49;
  wire v372a696;
  wire v3731d87;
  wire v373b0e7;
  wire v372f349;
  wire v3a5cfd9;
  wire v38099c1;
  wire v373e15b;
  wire v374cacb;
  wire v3a70198;
  wire v3a70dab;
  wire v376ca02;
  wire v377bcfc;
  wire v377c56c;
  wire v3808d48;
  wire v3a71194;
  wire v377974f;
  wire v3744af9;
  wire v3a709d1;
  wire v3a5e74c;
  wire v37652d7;
  wire v37380d5;
  wire v376c4fd;
  wire v373fd51;
  wire v3758c0d;
  wire v3a60787;
  wire v37736a6;
  wire v3733d6e;
  wire v3a6a213;
  wire v377851b;
  wire v3a704c7;
  wire v377edba;
  wire v373e267;
  wire v376f979;
  wire v377d74d;
  wire v372493b;
  wire v3a6e065;
  wire v3a707b5;
  wire v37455cd;
  wire v376a8be;
  wire v3742f0b;
  wire v3a6be50;
  wire v377d080;
  wire v3727699;
  wire v37528b0;
  wire v377cfd9;
  wire v37307de;
  wire v372ee7e;
  wire v373e8ad;
  wire v375a3dd;
  wire v3a6f2e1;
  wire v3a5c5f4;
  wire v373cde7;
  wire v376b654;
  wire v373cff4;
  wire v3a6febd;
  wire v373b03b;
  wire v3a60077;
  wire v372ee6a;
  wire v3755e64;
  wire v38087ee;
  wire v372b652;
  wire v3768ae9;
  wire v3a6d5a8;
  wire v3a709cd;
  wire v3a6fe72;
  wire v3a71585;
  wire v376ca61;
  wire v3763863;
  wire v374a9d4;
  wire v377a9b2;
  wire v3747020;
  wire v372a95a;
  wire v374ff02;
  wire v3765298;
  wire v3a713c0;
  wire v3a6f8c5;
  wire v3742e95;
  wire v3a67a78;
  wire v374c4c0;
  wire v3768e1e;
  wire v3a714b7;
  wire v3748984;
  wire v373d09a;
  wire v375d20f;
  wire c8ca6f;
  wire v37738b2;
  wire v377de4d;
  wire v376a0e6;
  wire v37478dd;
  wire v3a70b2a;
  wire v377516c;
  wire v373d4f7;
  wire v3a63cf5;
  wire v3a69df3;
  wire v3a6f74f;
  wire v377c831;
  wire v376d810;
  wire v3a6ef21;
  wire v3a6b5ba;
  wire v3a6f5ff;
  wire v37489a0;
  wire v3779288;
  wire v23fd8b7;
  wire v372a1bd;
  wire v3a6fdce;
  wire v3730876;
  wire v373ad86;
  wire v3740f78;
  wire v3747737;
  wire v37552cb;
  wire v3a5a06e;
  wire v37382ee;
  wire v3726f76;
  wire v375de72;
  wire v3a67d0d;
  wire d7f9ec;
  wire v3a70c80;
  wire v3a65540;
  wire v3a69a50;
  wire v373191d;
  wire v374fc95;
  wire v3a704b3;
  wire v3a70c59;
  wire v377ba7d;
  wire v3a6fc99;
  wire v374fad5;
  wire v372cafb;
  wire v3a66c84;
  wire v374fd12;
  wire v3730828;
  wire v3737846;
  wire v3a6ad46;
  wire v372ffd3;
  wire v3753a9f;
  wire v3731ea5;
  wire v3a6f376;
  wire v8ce84c;
  wire v374c048;
  wire v3775c51;
  wire v37624a5;
  wire v374f5a1;
  wire v372ab63;
  wire v3a53cf1;
  wire v374df3c;
  wire v2acb0b1;
  wire v3a613da;
  wire v3752def;
  wire v3a6f733;
  wire v3777d51;
  wire v3761f2b;
  wire v380946e;
  wire v3772e82;
  wire v3a714b9;
  wire v3734f6d;
  wire v3a6ff71;
  wire v3755c0e;
  wire v3a68377;
  wire v3809e97;
  wire v3770032;
  wire v3a5cd51;
  wire v373e10f;
  wire v3a5ad1d;
  wire v37731ce;
  wire v3a66cd7;
  wire acbf77;
  wire v3a5d97a;
  wire v373bd5e;
  wire v38098bf;
  wire v374943a;
  wire v3a69949;
  wire v3730019;
  wire v3a5f3a1;
  wire v1e374d4;
  wire v3737c88;
  wire v3a710ae;
  wire v3766f2e;
  wire v3a5d841;
  wire v3a5cccf;
  wire v374bfd2;
  wire v3a5373e;
  wire v373fdae;
  wire v373861f;
  wire v372af40;
  wire v3774f07;
  wire v3752f43;
  wire v37389b1;
  wire v3753fe6;
  wire v3a70d48;
  wire v3a70392;
  wire v3a6a9cd;
  wire v3772f09;
  wire v37500e0;
  wire v3a5cb4c;
  wire v377a522;
  wire v372f006;
  wire v377ce5a;
  wire v3a67d49;
  wire v3a5fae4;
  wire v374bc20;
  wire v3736d5e;
  wire v3731866;
  wire d5e2c2;
  wire v3a6fc2b;
  wire v376075c;
  wire v3a6fd5d;
  wire v3a6f5b8;
  wire v372f434;
  wire v376bce3;
  wire v3a54f8a;
  wire v3a58182;
  wire v3726d60;
  wire v3a6fcb6;
  wire v375b342;
  wire v374a50a;
  wire v3772aa4;
  wire v3808943;
  wire v3a692c3;
  wire v3a5943e;
  wire v3778e2d;
  wire v373c5dc;
  wire v38097ae;
  wire v3a6fb3e;
  wire v3764de1;
  wire v3769a62;
  wire v37242f1;
  wire v3a5d94f;
  wire v3a560b8;
  wire v375384f;
  wire v377baf9;
  wire v374f857;
  wire v3731dc1;
  wire v376c322;
  wire v3a54b43;
  wire v3a6d574;
  wire v3a5459f;
  wire v377ed4b;
  wire v377a993;
  wire v3739698;
  wire v3a71215;
  wire v37586cd;
  wire v373b4aa;
  wire v3806fc0;
  wire v37799a0;
  wire v3740766;
  wire v37755ff;
  wire v3a70cb0;
  wire v3767e03;
  wire v1e37e1f;
  wire v373e121;
  wire v3a6f523;
  wire v37266d9;
  wire v373fede;
  wire v8727d2;
  wire v372af6d;
  wire v3a6fbe8;
  wire v3a708b5;
  wire v3806a7b;
  wire v3769b75;
  wire v3766cfc;
  wire v3754e8c;
  wire v376dfc9;
  wire v3769f61;
  wire v377ab1f;
  wire v31c3694;
  wire v373cdbf;
  wire v3a6eeb5;
  wire v374c936;
  wire v3a6665c;
  wire v3a583dc;
  wire v377aede;
  wire v376aedb;
  wire v37432cd;
  wire v3a59505;
  wire v380649c;
  wire v3728eef;
  wire v37243d7;
  wire v3727517;
  wire v3776670;
  wire v3a6f2dd;
  wire v374f1c3;
  wire v3a55630;
  wire v374bf59;
  wire v3777cfc;
  wire v3a624d1;
  wire v3a60a9f;
  wire v3a64fee;
  wire v3a60125;
  wire v3a704af;
  wire v37439a0;
  wire v3a614d5;
  wire v3a5cb95;
  wire v373d11f;
  wire v37571ad;
  wire v3a5a3c7;
  wire v377057a;
  wire v37262fd;
  wire v374288a;
  wire v37455ec;
  wire v37720ca;
  wire v3a7089f;
  wire v3a58db9;
  wire v3a71026;
  wire v3a5e7c4;
  wire v3a5b20c;
  wire v3378c5b;
  wire v3a691ea;
  wire v373b710;
  wire v1e37ca9;
  wire v375b80e;
  wire v39a4dd7;
  wire v3726668;
  wire v37773c1;
  wire v3a6079f;
  wire v377eb7a;
  wire v3773f4e;
  wire v3a5f2c7;
  wire v377a942;
  wire v37320bf;
  wire v3770b73;
  wire v376669c;
  wire a9ca33;
  wire v377af60;
  wire v374a66c;
  wire v3752e82;
  wire v373042a;
  wire v375038a;
  wire v3768de8;
  wire v3a70145;
  wire v99797a;
  wire v3728b31;
  wire v3a70f2d;
  wire v374ef4a;
  wire v374d7a7;
  wire v3763b9b;
  wire v3a6cb16;
  wire v3a71121;
  wire v375917f;
  wire v376dfed;
  wire v3a6f4b6;
  wire v376bf8d;
  wire v375a250;
  wire v3777c39;
  wire v373f704;
  wire v3a701a0;
  wire v374743d;
  wire v3734b97;
  wire v3a70fa7;
  wire v3a70115;
  wire v376b363;
  wire v3a58964;
  wire v37237bc;
  wire v3a71542;
  wire v374578a;
  wire v3a6dd65;
  wire v3742657;
  wire v3a70c3a;
  wire v3a68793;
  wire v372e9ef;
  wire v3723e2f;
  wire v377fb50;
  wire v3a65b10;
  wire v373b956;
  wire v3747aa5;
  wire v3a596df;
  wire v372f55a;
  wire v3768c78;
  wire v37572df;
  wire v37467f7;
  wire v37777a2;
  wire v3a71647;
  wire v3a6fe80;
  wire v3762bf1;
  wire v3754c2d;
  wire v372fb9d;
  wire v3744458;
  wire v3a70393;
  wire v372615f;
  wire v37599eb;
  wire v3733228;
  wire v3767938;
  wire v3763813;
  wire v3a6f8dd;
  wire v3731b88;
  wire v376b23a;
  wire v3809f1c;
  wire v376f938;
  wire v23fe10d;
  wire v3a6bbee;
  wire v373fcae;
  wire v3808c66;
  wire v3a5b7e7;
  wire v372707d;
  wire v373bee7;
  wire v3761ae0;
  wire v3770f17;
  wire v37630ff;
  wire v3764005;
  wire v3a6d88e;
  wire v3738a2a;
  wire v3a6fe7c;
  wire v37504f2;
  wire v3a71541;
  wire v3a62949;
  wire v3a6f7cd;
  wire v375fa16;
  wire v3a70ebc;
  wire v376db9b;
  wire v3a70077;
  wire v3768739;
  wire v3777149;
  wire v37766cf;
  wire v3a5733c;
  wire v3745428;
  wire v377a617;
  wire v3a700ae;
  wire v3774b89;
  wire v3a55a19;
  wire v3a64643;
  wire v372f7c6;
  wire v373ae22;
  wire v3a701a9;
  wire v3756cf0;
  wire v3a5bdd2;
  wire v374006f;
  wire v380949b;
  wire v3a62d18;
  wire v3a71304;
  wire v8ed2d8;
  wire v3a6f1a5;
  wire v3774276;
  wire v3a6efb6;
  wire v3772b34;
  wire v3a63f30;
  wire v3773e41;
  wire v3a660e9;
  wire v3a57c2a;
  wire v3764370;
  wire be166e;
  wire v3740e4c;
  wire v3767b62;
  wire v3a6fc3b;
  wire v3a6814a;
  wire v3749c4b;
  wire v3a6d096;
  wire v3a70446;
  wire v3807a80;
  wire v3a6f454;
  wire a54211;
  wire v37761ae;
  wire v3729880;
  wire v3722eaf;
  wire v3a70bb2;
  wire v3a664b8;
  wire v3a5c904;
  wire v37562f2;
  wire v23fde98;
  wire v373abbb;
  wire v3747400;
  wire v37bfc8b;
  wire v3736411;
  wire v3746d52;
  wire v374c73c;
  wire v3a5591a;
  wire v377586d;
  wire v3724f6b;
  wire abd043;
  wire v37337fd;
  wire v3a6f382;
  wire v3a62fd2;
  wire v3a693b7;
  wire v37327fe;
  wire v3a65e1a;
  wire v377b5dc;
  wire v3a69a00;
  wire v372e44d;
  wire v377f78c;
  wire v377d202;
  wire v3a56243;
  wire v3a5f449;
  wire v37419e7;
  wire v3738bf6;
  wire v38076c9;
  wire v3a63111;
  wire v3a6b6f2;
  wire v3779a66;
  wire v3731003;
  wire v373b3a8;
  wire v3a56d01;
  wire v3a55723;
  wire v373d025;
  wire v3a6f53d;
  wire v3a5e09d;
  wire v3759a88;
  wire v3808881;
  wire v3749c8a;
  wire v3a6039a;
  wire v37233a2;
  wire v376935b;
  wire v3a705de;
  wire v374f557;
  wire v3a61fcc;
  wire v3a70094;
  wire v3a6f54d;
  wire v3a71275;
  wire v37381bb;
  wire v373e782;
  wire v374203a;
  wire v3768a79;
  wire v3a70ece;
  wire v35b7044;
  wire v3761adc;
  wire v3a71420;
  wire v3754892;
  wire v377ea72;
  wire v3a5b89b;
  wire v372479c;
  wire v337948a;
  wire c7f8d6;
  wire v3773069;
  wire v3767527;
  wire v377c4bd;
  wire v3a5cc3c;
  wire v3a6488f;
  wire v3755451;
  wire v3258762;
  wire v377dedb;
  wire v3a6ff80;
  wire v3744ea3;
  wire v376cd2f;
  wire v37247a3;
  wire v2ff9391;
  wire v3767744;
  wire v375b0d4;
  wire v3749cf4;
  wire v23fe052;
  wire v3a5aef6;
  wire v3a69118;
  wire v3a2abf5;
  wire v38064dd;
  wire v3766185;
  wire v375bf12;
  wire v3733c51;
  wire v3a5db7f;
  wire v2ff9397;
  wire v3764c6c;
  wire v39ea2e3;
  wire v372977b;
  wire v3a6fea0;
  wire v3744a2f;
  wire v3a57e21;
  wire v3a6f351;
  wire v3734312;
  wire v3771b20;
  wire v376f30a;
  wire v377d34b;
  wire v3730693;
  wire v375bc5b;
  wire v3a714ac;
  wire v3758988;
  wire v3778151;
  wire v377e172;
  wire v372f5ec;
  wire v3731a49;
  wire v373173b;
  wire v3a550cd;
  wire v37780e2;
  wire v3a7121f;
  wire v3776f93;
  wire v3a66747;
  wire v3768036;
  wire v3758663;
  wire v3a6f543;
  wire v3a70064;
  wire v3a70500;
  wire dc3a01;
  wire v3739c9a;
  wire ce3eb4;
  wire v3744314;
  wire v1e37d71;
  wire v37308ae;
  wire v3752ee5;
  wire v3a5dd60;
  wire v3a70b46;
  wire v373f8c8;
  wire v3a6aada;
  wire v3a53f38;
  wire v3a6f06a;
  wire v373c8c3;
  wire v376fa38;
  wire v3a695fc;
  wire v3746a81;
  wire v3742aff;
  wire v2092ba8;
  wire v38088f5;
  wire v3a6932d;
  wire v37628cd;
  wire v37285fa;
  wire v3a6f814;
  wire v3a58aa5;
  wire v3a59e87;
  wire v3725098;
  wire d23bf8;
  wire v3a70a32;
  wire v3a6eb3f;
  wire v373ad3f;
  wire v3739531;
  wire v3a7114c;
  wire v37626d8;
  wire v3a70ea2;
  wire v3750f60;
  wire v374e168;
  wire v3a66a3a;
  wire v37244f3;
  wire v373418b;
  wire v3a67269;
  wire a792d5;
  wire v3a7064c;
  wire v3a6b07b;
  wire v376480b;
  wire v3755fd4;
  wire v3a688f9;
  wire v373281b;
  wire v3a70069;
  wire v3a6d684;
  wire v3808e82;
  wire v374055c;
  wire v373d07a;
  wire v3a70dd8;
  wire v37733d9;
  wire v3766853;
  wire v3a66ca4;
  wire v37780fd;
  wire v3a694b4;
  wire b6057e;
  wire v37582e6;
  wire v377cbb6;
  wire v3734a96;
  wire v3a644ac;
  wire v3a6f5a6;
  wire v37473c5;
  wire v1e37776;
  wire v37638f9;
  wire v39ea76e;
  wire v3a714d8;
  wire v3a6ff27;
  wire v377a87d;
  wire v3a533d8;
  wire v377ea6c;
  wire v377601b;
  wire v372459b;
  wire v376dae8;
  wire v3a621e6;
  wire v3761f57;
  wire v377866b;
  wire v3779486;
  wire v377e9c1;
  wire v377598a;
  wire v3a6f1bf;
  wire v3a6ed14;
  wire v3a681f5;
  wire d03e23;
  wire v3a70533;
  wire v3724734;
  wire v3a5be0b;
  wire v3a6cbfa;
  wire v9d7045;
  wire v377c490;
  wire v375c67c;
  wire v3a6a893;
  wire v375912e;
  wire v3a6bf00;
  wire v3a6ffde;
  wire v3748d8c;
  wire v3734c60;
  wire v376e41a;
  wire v3a70f19;
  wire v373e748;
  wire v374c53a;
  wire v3a62542;
  wire v3a55b6c;
  wire v3a6ea51;
  wire v374dfd9;
  wire v3766709;
  wire v3757b0e;
  wire v3778567;
  wire v377accc;
  wire v3a70221;
  wire v37606c7;
  wire v373da69;
  wire v3a5e02b;
  wire v3a2981b;
  wire v3a70970;
  wire v372f37d;
  wire v3a6fa93;
  wire v377c8d1;
  wire v3a6fb2f;
  wire v3a672c8;
  wire v3738666;
  wire v3a5c9df;
  wire v37398a1;
  wire v3a708d8;
  wire v3a6f32a;
  wire v3a6f4fc;
  wire v37498be;
  wire v372949c;
  wire v3723ee7;
  wire v37711c5;
  wire v37745a0;
  wire v3a595fe;
  wire v3a5c066;
  wire v3762997;
  wire v372e2cd;
  wire v376ce55;
  wire v3732b3a;
  wire v375abaa;
  wire v3a70ab8;
  wire v3733027;
  wire v3a6ffd3;
  wire v373af55;
  wire v3a6a1d1;
  wire v373fdf0;
  wire v3a70d9b;
  wire ab15ca;
  wire v3a6f7b5;
  wire v3a5ebc8;
  wire v372fc7e;
  wire v3747897;
  wire v3a634b9;
  wire v3a548c2;
  wire v3736471;
  wire v3755096;
  wire v372a264;
  wire v3a5e485;
  wire v3738ce7;
  wire v376454b;
  wire v374b36e;
  wire v372b1c8;
  wire v37380c4;
  wire v377e5ac;
  wire v3748194;
  wire v3a6eeba;
  wire v37545a5;
  wire v3a7137a;
  wire v3a7080a;
  wire v39e9c97;
  wire v372a7ae;
  wire v3735a7c;
  wire v372f100;
  wire v372c1fc;
  wire v3a6ebd2;
  wire v3a70d65;
  wire v3743a2c;
  wire v3737f5f;
  wire v3a59720;
  wire v28896c8;
  wire v3736da4;
  wire v37770d2;
  wire v3a55640;
  wire v373698e;
  wire v372e94f;
  wire v3a5bffe;
  wire v3a70731;
  wire v376460f;
  wire v3a70964;
  wire v3a70070;
  wire v37c014e;
  wire v3a709bf;
  wire v374db9d;
  wire v374b8cb;
  wire v3766345;
  wire v3776ea4;
  wire v380951e;
  wire v37712b7;
  wire v375471b;
  wire v3a711e4;
  wire v3731999;
  wire v374ec57;
  wire v375bb06;
  wire v3a6f5f9;
  wire v3774fee;
  wire v3a70117;
  wire v3a6220e;
  wire v375005c;
  wire v3734de2;
  wire v3a66988;
  wire v375ab04;
  wire v3a71270;
  wire v3a702c6;
  wire v3a6eb4a;
  wire v374c052;
  wire v3a70557;
  wire v373296d;
  wire v3a70adb;
  wire v3776d42;
  wire v3a7167c;
  wire v3737a6e;
  wire v3a6d5e2;
  wire v3740cb5;
  wire v3a703a0;
  wire v3a715c4;
  wire v3726570;
  wire v377baa6;
  wire v3768ce2;
  wire v376d28f;
  wire v375e2d3;
  wire v3775642;
  wire v375c265;
  wire v3378d8f;
  wire v3736610;
  wire v37234e7;
  wire v3728df3;
  wire v3770cd8;
  wire v3747eef;
  wire v3a6f989;
  wire v376a7e8;
  wire v3a64d23;
  wire v3a6e81e;
  wire v2acafcc;
  wire v373f5ab;
  wire v375d9ad;
  wire v3a71043;
  wire v375d351;
  wire v37603f4;
  wire v3762bbe;
  wire v376b3b0;
  wire v376049c;
  wire v3a6f807;
  wire v377d4ab;
  wire v372ef40;
  wire v3a71012;
  wire v3a70957;
  wire v3749846;
  wire v3749a17;
  wire v3728d28;
  wire v374a9fa;
  wire v3779fdf;
  wire v375a26b;
  wire v374910b;
  wire v3a66983;
  wire v3a569e1;
  wire v37474f3;
  wire v3a6f997;
  wire v3a6fa8e;
  wire v374a668;
  wire v3a54c12;
  wire v23fe329;
  wire v3a6937a;
  wire v3770db3;
  wire v3756e39;
  wire v37469db;
  wire v3737fe0;
  wire v3a645f6;
  wire v3a70913;
  wire v373632b;
  wire v3a5d1fb;
  wire v3773b55;
  wire v3a5aa9d;
  wire v3a63d3c;
  wire v374aa71;
  wire v3759279;
  wire v3a71170;
  wire v376c2b7;
  wire v3a5cfed;
  wire v376ad4e;
  wire v373c703;
  wire v39ea273;
  wire v3772c57;
  wire v3739732;
  wire v3739dd4;
  wire v3a632d8;
  wire v372362a;
  wire v3a71459;
  wire v3730a8b;
  wire v3a6fd31;
  wire v373a973;
  wire v374e684;
  wire v377dfbd;
  wire v3724da7;
  wire v3a633bf;
  wire v3733ee4;
  wire v3a612df;
  wire v3a2981d;
  wire v3a6f058;
  wire v373628a;
  wire v375e3a1;
  wire v3a6e733;
  wire v37353be;
  wire v3725688;
  wire v3a5a814;
  wire v3763e6c;
  wire v376e954;
  wire v3736dfd;
  wire v372919e;
  wire v3a70afd;
  wire v38068ec;
  wire v3a67315;
  wire v3a6fc6d;
  wire v9381f3;
  wire v3739d9b;
  wire v3a7132c;
  wire v3a549f5;
  wire v3756bc9;
  wire v375c5a8;
  wire v3749ec6;
  wire v3a695b7;
  wire v3a71041;
  wire v3a6f860;
  wire v3727740;
  wire v2092faa;
  wire v3751861;
  wire v373c642;
  wire v3776eef;
  wire v3740dc8;
  wire v3a6843e;
  wire v37667e4;
  wire v375e91e;
  wire v376a7bf;
  wire v3734965;
  wire v37266bd;
  wire v3730b5a;
  wire v3a68d26;
  wire v375f99c;
  wire v373b9e9;
  wire v3738d54;
  wire v3a5b01c;
  wire v373eeed;
  wire v3a6f227;
  wire v377eed2;
  wire v3a5803d;
  wire v3736fb1;
  wire v3a5c0f8;
  wire v3a54271;
  wire v37358ae;
  wire v37431c0;
  wire v3729f13;
  wire v3732a95;
  wire v3746085;
  wire v376964c;
  wire v373d071;
  wire v3a68931;
  wire dacf90;
  wire v3a60bc1;
  wire v37681ec;
  wire v3a6eef0;
  wire v3737438;
  wire v377815b;
  wire v3a5fae3;
  wire v3726c61;
  wire v3a6f49f;
  wire v377f6c3;
  wire v37476c5;
  wire v3a71193;
  wire v3a5be70;
  wire v373e941;
  wire v3a62e77;
  wire v372647c;
  wire v376b71f;
  wire v3a6f7eb;
  wire v3a5d930;
  wire v374bbca;
  wire v375f3bc;
  wire v3a6202c;
  wire v37348f8;
  wire v372ad5a;
  wire v374f92e;
  wire v3725de9;
  wire v3a6d7a0;
  wire v3a64eb3;
  wire v3747b29;
  wire v37653a2;
  wire v375a30e;
  wire v37247c8;
  wire v3a70657;
  wire v374f7f8;
  wire v3760337;
  wire v3a5de1e;
  wire v3729139;
  wire v3a70ab7;
  wire v3a69adb;
  wire v372fd97;
  wire v3a7152c;
  wire v377c7ce;
  wire v376a31b;
  wire v8a7f7e;
  wire v3a6edb1;
  wire v37790a9;
  wire v3743d58;
  wire v3a6a442;
  wire v3762870;
  wire v376e7f5;
  wire v3753389;
  wire v376596e;
  wire v377adaa;
  wire v3a70bce;
  wire bc7f17;
  wire v3756ca5;
  wire v37609a6;
  wire v37235bd;
  wire v376da22;
  wire v3a715f7;
  wire v377da1e;
  wire v373ebd2;
  wire v3a7089e;
  wire v375c551;
  wire v374ca2d;
  wire v3a6f8a1;
  wire v3a6f04a;
  wire v374c234;
  wire v3a61254;
  wire v3a700a5;
  wire bda6d5;
  wire v3a58836;
  wire v374e0ba;
  wire v3a702ed;
  wire v375b21c;
  wire aef136;
  wire v3763c82;
  wire v3749d74;
  wire v37612f7;
  wire v3a54aa0;
  wire v3a6368a;
  wire v3779324;
  wire v3769039;
  wire v37393cc;
  wire v3a6acbb;
  wire v3749380;
  wire v3a69df1;
  wire v377a551;
  wire v3a6f995;
  wire v3a710f7;
  wire v37229ba;
  wire v3a700e6;
  wire v37523de;
  wire v374648b;
  wire v3729724;
  wire v3732aa6;
  wire v375da3a;
  wire a21c18;
  wire v3a71646;
  wire v37728d3;
  wire v3758700;
  wire v23fdd06;
  wire v3749f86;
  wire v3a61a15;
  wire v377a673;
  wire v373e792;
  wire v3750e4b;
  wire v375452a;
  wire v3a7147c;
  wire v3748544;
  wire v377167d;
  wire v3a6f31d;
  wire v3a67b5e;
  wire v37649ee;
  wire v3771026;
  wire v3745a7b;
  wire v922c1b;
  wire a4764c;
  wire v374774d;
  wire v3a6ef4c;
  wire v37607d2;
  wire v37243dc;
  wire c6a502;
  wire v3771696;
  wire d138a6;
  wire v37551df;
  wire v3a6fc46;
  wire v3a6ef4a;
  wire v3a64bc4;
  wire v376cd0d;
  wire v3757ce3;
  wire v325c9cb;
  wire v3a715f2;
  wire v3a59217;
  wire v37269a2;
  wire v3740083;
  wire v373040e;
  wire v3a714f0;
  wire v3a6494a;
  wire v3a6f6f4;
  wire v377e545;
  wire v3736d03;
  wire v3a7141c;
  wire v3752b8f;
  wire v3a59529;
  wire v3a54e41;
  wire v3a6e986;
  wire v3a60247;
  wire v3a70c17;
  wire v3a70d9e;
  wire v375ed60;
  wire v373c721;
  wire v377a6bf;
  wire v374a849;
  wire v3764f39;
  wire v376beca;
  wire v3a70538;
  wire v3a571d1;
  wire v3738eb0;
  wire v3739239;
  wire v377499f;
  wire v3a6ca1d;
  wire v3776d33;
  wire v3775311;
  wire d27e8c;
  wire v3726605;
  wire v3a6ff15;
  wire v372fb1b;
  wire v3a66584;
  wire v37540df;
  wire v3750b71;
  wire v37516cc;
  wire v376674a;
  wire v3a5d373;
  wire v374ae4a;
  wire v374f329;
  wire v372d42d;
  wire v37593a4;
  wire v373b7f5;
  wire aa6771;
  wire v3777ff7;
  wire v374089e;
  wire v3a630ba;
  wire v3a67dd0;
  wire v3775341;
  wire v374fa94;
  wire v3758c46;
  wire v3759181;
  wire v3744d18;
  wire v3752e24;
  wire v373a629;
  wire v3a6f6ec;
  wire v37585bf;
  wire v37541d3;
  wire v373cd0c;
  wire v373aec4;
  wire v3759bdb;
  wire ca9b68;
  wire v3779e72;
  wire v3a69a1b;
  wire v3734129;
  wire v3777b84;
  wire v3a6bd0f;
  wire v3764f60;
  wire v3a29520;
  wire v375c4c7;
  wire v373c342;
  wire v8f4f53;
  wire v37449e7;
  wire v373627b;
  wire v37493ed;
  wire v3a6efc3;
  wire c8bdc6;
  wire v3763f1d;
  wire v3a70120;
  wire v3754ca0;
  wire v3a70dc1;
  wire v3378a2d;
  wire v3a70a31;
  wire v37c028b;
  wire v3776e2b;
  wire v3745315;
  wire v3763c20;
  wire v3a710d8;
  wire v1e37c79;
  wire v3a704b4;
  wire v374083d;
  wire aeaf7c;
  wire v372542e;
  wire v374fdc9;
  wire v3a61b9d;
  wire v37414be;
  wire v3a649c2;
  wire v3a6f8c9;
  wire v3734b14;
  wire v3807abe;
  wire v3a7156b;
  wire v3735ec7;
  wire v3758c5c;
  wire v3a7121e;
  wire v3a70646;
  wire v376cc0e;
  wire v376f2f4;
  wire v3a70968;
  wire v37662f4;
  wire b66740;
  wire v1e37784;
  wire v9b81ab;
  wire v3a713bb;
  wire v3770093;
  wire v376df3c;
  wire v3a56f2d;
  wire v377a0f2;
  wire v37629ba;
  wire v3a70ee7;
  wire v3a6f312;
  wire v3765466;
  wire v374ad81;
  wire v3a6eaf4;
  wire v37665e1;
  wire v377e7ac;
  wire v373bc28;
  wire v3762807;
  wire v3722caa;
  wire v3a70a82;
  wire v3738a93;
  wire v372fbb1;
  wire v3778e98;
  wire v373485b;
  wire v3808cf7;
  wire v3a61375;
  wire v3a6a82d;
  wire v374e02b;
  wire v3742472;
  wire v373782c;
  wire v3a55ec8;
  wire v373eef7;
  wire v3a7006c;
  wire v3744d60;
  wire v373a7a1;
  wire v3a62541;
  wire v3a6e943;
  wire v375c6f5;
  wire v3768ba9;
  wire v374f34b;
  wire v373afd0;
  wire v376e074;
  wire v3742146;
  wire v37287be;
  wire v3774542;
  wire v375f0f0;
  wire v3a6f665;
  wire v374d0ad;
  wire v3a70cc9;
  wire v3a6f327;
  wire v38068c1;
  wire v37626ab;
  wire v3a6961d;
  wire v3a6aaa4;
  wire v8dc5a6;
  wire v3763590;
  wire v3778f81;
  wire v377f5c9;
  wire v3733b65;
  wire b33e26;
  wire v3a6fcd1;
  wire v3740d36;
  wire c99197;
  wire v3768ab0;
  wire v3577416;
  wire v372dcc2;
  wire v37584c7;
  wire a568f8;
  wire v3a6f415;
  wire v3a6d1a4;
  wire v3758dfe;
  wire v3a6ef23;
  wire v377594d;
  wire v373ad2b;
  wire v375649a;
  wire v3778fab;
  wire v3743e4a;
  wire v3a665b4;
  wire v37485f0;
  wire v3a6eee6;
  wire v377bb21;
  wire v373d72e;
  wire v372e0b0;
  wire v3747586;
  wire v3a6f4ce;
  wire v3768690;
  wire v3745498;
  wire v373b4c8;
  wire v3a6f900;
  wire v377a312;
  wire v376e6ac;
  wire v37431bb;
  wire v373a11f;
  wire v37400f3;
  wire v37650dd;
  wire v3737ac8;
  wire v3744161;
  wire v3754d8a;
  wire v37292df;
  wire v3737c0d;
  wire v374bddc;
  wire v375b98c;
  wire v3727dd4;
  wire v375b3f0;
  wire v372ee98;
  wire v3a5c0de;
  wire v3a6f0e3;
  wire v37317c0;
  wire v3a5db8b;
  wire v3a6fcc3;
  wire v23fe0c9;
  wire v3577484;
  wire v3a53f1a;
  wire v375098f;
  wire v3762244;
  wire v373aa77;
  wire v377d7dd;
  wire v374cc7f;
  wire v3722f3b;
  wire v374affb;
  wire v3a67869;
  wire v37483f9;
  wire v3a695c9;
  wire v3778464;
  wire v3779736;
  wire v375af99;
  wire v3a70382;
  wire v37640de;
  wire v372815e;
  wire v3748929;
  wire v3736c8c;
  wire v373a77b;
  wire v3a6ff1f;
  wire v3748234;
  wire v373d703;
  wire v3735749;
  wire v3a6f925;
  wire v3a7162b;
  wire v3747d69;
  wire v3723d16;
  wire v3a709ce;
  wire v375dcf8;
  wire v3765293;
  wire v3a61c5e;
  wire v374b64d;
  wire v3732aab;
  wire v1e37583;
  wire v3146177;
  wire v377882e;
  wire v3728a9f;
  wire v3a6706d;
  wire v3a644d3;
  wire v3a57b11;
  wire v3a6b475;
  wire v31461d5;
  wire v3a5b6c5;
  wire v375bd0e;
  wire v373f880;
  wire v3736079;
  wire b8cdcc;
  wire v94c82c;
  wire v28e9804;
  wire v3a64792;
  wire v3a6dc83;
  wire v372b88d;
  wire v3759c1f;
  wire v37466b7;
  wire v3735274;
  wire v374a0c4;
  wire v3759886;
  wire v377234d;
  wire v37504eb;
  wire v3773200;
  wire v3743910;
  wire v3759a67;
  wire v375295a;
  wire v3a70e7a;
  wire v375121b;
  wire v377d9aa;
  wire v3740541;
  wire v3772080;
  wire v377a812;
  wire v3a5d94a;
  wire v374da1a;
  wire v374b497;
  wire v3779f92;
  wire v35b7734;
  wire v37480b7;
  wire v3748ac8;
  wire v3a6f42a;
  wire v3a702da;
  wire v360d140;
  wire v3a58803;
  wire v375d3bb;
  wire v37358ab;
  wire v3754a25;
  wire v3a67a6f;
  wire v3a5d7ba;
  wire v373c58c;
  wire v372b006;
  wire v376053b;
  wire v372c09e;
  wire v374ab4c;
  wire v3a6f9be;
  wire v37291f8;
  wire v3734b34;
  wire v375463e;
  wire v3a5f974;
  wire v3755b56;
  wire v3756dd8;
  wire v37519e3;
  wire v3769950;
  wire v377818c;
  wire v3778b60;
  wire v374e6b1;
  wire v3769c6d;
  wire v3730be2;
  wire v3739b4c;
  wire v3a58287;
  wire v376f9eb;
  wire v37579ab;
  wire v3808e2e;
  wire v373859f;
  wire v3a5841e;
  wire v376926f;
  wire v377c9cb;
  wire v375f172;
  wire v37735aa;
  wire v3a70442;
  wire b8f82c;
  wire v3a6fdb6;
  wire v374757c;
  wire v3a53d2b;
  wire v3a6fb65;
  wire v3779071;
  wire v3a6ebfc;
  wire v3759232;
  wire v3a715e6;
  wire v3745a5f;
  wire v3777a00;
  wire v375bb10;
  wire v375c4e6;
  wire v3a70e3d;
  wire v372cdd5;
  wire v3a6870f;
  wire v3744f62;
  wire v3a6b597;
  wire v3a5bea0;
  wire v37744d9;
  wire v37255f6;
  wire v3a6f59d;
  wire v372ae6f;
  wire v3a58e44;
  wire v375ecab;
  wire v3740663;
  wire v37470e2;
  wire v37675f1;
  wire v3743b62;
  wire v374c6c5;
  wire v3775d26;
  wire v3733e30;
  wire v3a66910;
  wire v375fbbb;
  wire v3a6e37c;
  wire v3764132;
  wire v3736db2;
  wire v377ba8a;
  wire v3a69b77;
  wire v3a6f4f9;
  wire v376d86c;
  wire v3a71182;
  wire v377409c;
  wire d6aeaf;
  wire v374cb21;
  wire v3a6f446;
  wire v374350d;
  wire v3a70da2;
  wire v3a66e9f;
  wire v3735a87;
  wire v3a6f76b;
  wire v3a70981;
  wire b4f354;
  wire v3724b94;
  wire v37315fd;
  wire v3763afe;
  wire v3741fea;
  wire v3a6c9aa;
  wire v374db73;
  wire v3779177;
  wire v37bfc8a;
  wire v373a54d;
  wire v37418bf;
  wire v376025c;
  wire v3a59900;
  wire v372589e;
  wire v375bfe5;
  wire v3a6f5cb;
  wire v32587ac;
  wire v3764448;
  wire v3725e4b;
  wire v3725371;
  wire v3766669;
  wire v3726dfd;
  wire v3729949;
  wire v377b7e0;
  wire v3722d8b;
  wire v3a6be9f;
  wire v3a6f72e;
  wire v372e440;
  wire v374c251;
  wire v3a70874;
  wire v372a636;
  wire v376efaa;
  wire v3a6fa8f;
  wire v374dc1b;
  wire v3749975;
  wire v373f75b;
  wire v3a55d4c;
  wire v3758e8d;
  wire v375d76b;
  wire v374156a;
  wire v3a6f259;
  wire v3a56e45;
  wire v372b1e8;
  wire v3a6ce52;
  wire v375a804;
  wire v3a55a58;
  wire v3a65dad;
  wire v3741249;
  wire v374597c;
  wire v2acaec4;
  wire v374c28d;
  wire v373b938;
  wire v3736382;
  wire v3a69dd2;
  wire v375e73a;
  wire v377a68a;
  wire v3773071;
  wire v377d1dc;
  wire v37763d1;
  wire v3a6fd10;
  wire v372cdec;
  wire v1e37b99;
  wire v373b02e;
  wire v373b887;
  wire v3a5cf28;
  wire v3750abf;
  wire v3755f22;
  wire v3a65552;
  wire v3a71435;
  wire v3a55542;
  wire v89fdcf;
  wire v372efcb;
  wire v3762c7f;
  wire v37244f1;
  wire a61f6b;
  wire v375c263;
  wire v3a6e5e1;
  wire v3a65605;
  wire v3752f2e;
  wire v377871a;
  wire v3758d18;
  wire v3755ad5;
  wire v372625f;
  wire v372a5c8;
  wire v3a711d8;
  wire v35b71af;
  wire v372d630;
  wire v3808f45;
  wire v3747d58;
  wire v372b6ec;
  wire v3a6fc7d;
  wire v3772e0c;
  wire v3761300;
  wire v3a5c7a2;
  wire v3a6f796;
  wire v37647de;
  wire v37525c8;
  wire v3754717;
  wire v373d98d;
  wire v377f630;
  wire v33790e7;
  wire v3765739;
  wire v376a943;
  wire v3769e8c;
  wire v374bf55;
  wire v377ad9c;
  wire v3a65fa5;
  wire v3a7106d;
  wire v37297d0;
  wire v374d1dc;
  wire v3736ad7;
  wire v375ab89;
  wire v37510d0;
  wire v373b4dc;
  wire v375a8d6;
  wire v377cef3;
  wire v3a705f1;
  wire v3a7131d;
  wire v3755000;
  wire v3a704a3;
  wire v377d232;
  wire v3731c2f;
  wire v373d42f;
  wire v3a5eb8f;
  wire v3762f5b;
  wire v3a6fbb5;
  wire v3761431;
  wire v3757519;
  wire v3a5b40f;
  wire v98083e;
  wire v37739f4;
  wire v3a576d0;
  wire v3722b92;
  wire v375f486;
  wire v376bca9;
  wire a7394c;
  wire v3a638aa;
  wire v3728685;
  wire v372cde4;
  wire v3a68525;
  wire v37298be;
  wire v37536b8;
  wire v377e871;
  wire v372d1d7;
  wire v3a712dd;
  wire v3a65069;
  wire v3a570ee;
  wire v3a5a162;
  wire v3a6f64d;
  wire v373f1aa;
  wire v3756e63;
  wire v3a6c849;
  wire cc8b5a;
  wire v3a7110e;
  wire v376a84d;
  wire v37673fe;
  wire v3a6ba91;
  wire v377326a;
  wire v375a16a;
  wire v373221a;
  wire v3761c5e;
  wire v377709a;
  wire v377a808;
  wire v3a573c2;
  wire v3a607bd;
  wire v3a71302;
  wire v3769160;
  wire v3764e52;
  wire v39eb4d4;
  wire v3763398;
  wire v37742f1;
  wire v374ebe8;
  wire v372d744;
  wire v374fe54;
  wire v376a63f;
  wire v3a711a4;
  wire v3774000;
  wire v3770bed;
  wire v376a399;
  wire v377d785;
  wire v3775e82;
  wire v3a64ad6;
  wire v3a5af5c;
  wire v3742995;
  wire v375cab0;
  wire v3a6599b;
  wire v3a70b51;
  wire v372567b;
  wire v360d109;
  wire v372cede;
  wire v3a6fd68;
  wire v3a62b11;
  wire v3a6efef;
  wire v3775269;
  wire v3741e54;
  wire v3a67b7f;
  wire v376bb43;
  wire v3a6b2e5;
  wire v372b7cc;
  wire v3733d45;
  wire a8fc27;
  wire v3724273;
  wire v3a56372;
  wire v377876f;
  wire v3a7119f;
  wire v3770027;
  wire v3726458;
  wire v3a702ff;
  wire v373933b;
  wire v375c317;
  wire v374fda4;
  wire a25d5b;
  wire v3a6a6c1;
  wire v3762f76;
  wire v372516b;
  wire v3a6f2d9;
  wire v37481bf;
  wire v3a63628;
  wire v3759aeb;
  wire v3a63e9b;
  wire v3a704d6;
  wire v374eb2d;
  wire v373f8c4;
  wire v37566c9;
  wire v3770a6d;
  wire v3a61532;
  wire v375dc25;
  wire v37520ee;
  wire v37641b8;
  wire v3724aa4;
  wire v1e37eb7;
  wire v3728fee;
  wire v374fd32;
  wire v3a56027;
  wire v377849a;
  wire v377c67b;
  wire v3756a5f;
  wire v3a70ab1;
  wire v3a6fd9f;
  wire v3724718;
  wire v3807686;
  wire v3a6f7ee;
  wire v3a6f130;
  wire v377e002;
  wire v3a70bf3;
  wire v372cd61;
  wire v373e0d0;
  wire v374ccb3;
  wire v3a6fe5c;
  wire v3a6f3e9;
  wire v3a580fb;
  wire v3741ab9;
  wire v3752b5c;
  wire v3724efc;
  wire v3a6652b;
  wire v3a6877a;
  wire v3a70989;
  wire v3806e5b;
  wire v3a70e6e;
  wire v3733cf4;
  wire v3745589;
  wire v375add1;
  wire v377d8d6;
  wire v3a5aca8;
  wire v377ba37;
  wire v3741925;
  wire v3a70fda;
  wire v23fd83c;
  wire v3a6f2ce;
  wire v3723a94;
  wire v3760da6;
  wire v372fa3a;
  wire v376dd48;
  wire v3739112;
  wire v3a585f1;
  wire v374d547;
  wire v376b6ba;
  wire v376beea;
  wire v3723923;
  wire v3777d2e;
  wire v3a6cf6a;
  wire v3757f0d;
  wire v372c8bc;
  wire v375805a;
  wire v37315e2;
  wire v2092ef2;
  wire v3729830;
  wire v97e702;
  wire v37387e6;
  wire v3729308;
  wire v374beee;
  wire v3a5a825;
  wire v372b7b1;
  wire v3a6b22e;
  wire v377c9c3;
  wire v3733955;
  wire v2aca76c;
  wire v375d57e;
  wire v377e89a;
  wire v3a6b478;
  wire v3765222;
  wire v3764257;
  wire v3a592bc;
  wire v3773103;
  wire v3a65ea7;
  wire v3a636d2;
  wire v376f250;
  wire v3808fc8;
  wire v374b6ee;
  wire v372a1f6;
  wire v375c099;
  wire v3a6f2f8;
  wire v373a0dc;
  wire v3769c4c;
  wire v3a704d2;
  wire v374e620;
  wire v3762324;
  wire v3a53a43;
  wire v37563bc;
  wire v37576af;
  wire v37457a8;
  wire v37288c3;
  wire v3742c62;
  wire v3a5b070;
  wire v3753aa5;
  wire v3725bd2;
  wire v3759dc9;
  wire v9c9e05;
  wire v37709d8;
  wire v3743a4d;
  wire v3755608;
  wire v376a246;
  wire v377789d;
  wire v3a67c36;
  wire v3a7097e;
  wire v375d06a;
  wire v376b27a;
  wire v376e1ad;
  wire v3a713a9;
  wire v3755289;
  wire v37235b8;
  wire v3a63d77;
  wire v37348f5;
  wire v3a57b00;
  wire v3740e9c;
  wire v3a70ed8;
  wire v376da8d;
  wire v37383bb;
  wire v37629d2;
  wire v375e34d;
  wire v374db79;
  wire v3a70dae;
  wire v375524f;
  wire v3a70e7b;
  wire v3769921;
  wire v372efcd;
  wire v3a64abe;
  wire v3a70e2d;
  wire v373f1ba;
  wire v3a70d5d;
  wire v3a6fc91;
  wire v3a70b57;
  wire v376b70a;
  wire v3a5f1db;
  wire ac69a2;
  wire v3765dbc;
  wire v374e0b8;
  wire v3a6f1eb;
  wire v3750d6d;
  wire v3a55377;
  wire v3255a0c;
  wire v3a6f728;
  wire v3727c6e;
  wire v37703cb;
  wire v3768e15;
  wire v3747133;
  wire af0958;
  wire v374c9e1;
  wire v3a704e6;
  wire v375df4f;
  wire v3745e63;
  wire v3a6f49b;
  wire v372c3e9;
  wire v3a6fca7;
  wire v3736518;
  wire v3737186;
  wire v37314cc;
  wire v3807aa1;
  wire v37c007b;
  wire v3a5979b;
  wire v3748b83;
  wire v23fde6a;
  wire v3a6fb3f;
  wire v3a5a7c6;
  wire v377c3a1;
  wire v3a6ec04;
  wire v375a67c;
  wire v375dc9b;
  wire v3a6d329;
  wire v3764e55;
  wire v35b7174;
  wire v3752536;
  wire v372b686;
  wire v3a70943;
  wire v3a69910;
  wire v3778cf7;
  wire v3777cb2;
  wire v3a584fd;
  wire v3766dc8;
  wire v3757506;
  wire v375c9f0;
  wire v3a6ef26;
  wire v3a6fb88;
  wire v372ac1d;
  wire v374f26c;
  wire v3a70059;
  wire v374cdc4;
  wire v3a70736;
  wire v37383d3;
  wire v3a70a90;
  wire v372e6d0;
  wire v372d2d2;
  wire v37586e2;
  wire v375f106;
  wire v3a697f1;
  wire v39ebbae;
  wire v3a5fc59;
  wire v3a6f963;
  wire v377278b;
  wire v3766c68;
  wire v37259cc;
  wire v374dce0;
  wire v3759119;
  wire v377f424;
  wire v2ff87d2;
  wire v3a66cad;
  wire v3a6d4f8;
  wire v3a614b1;
  wire v3a68f3d;
  wire v3a60767;
  wire v3746efa;
  wire v3a6f8ef;
  wire v37654ea;
  wire v373361a;
  wire v3769dfe;
  wire v3760700;
  wire v3731b90;
  wire v37232c0;
  wire v375b40c;
  wire v3779283;
  wire v3a5be74;
  wire v372ce8b;
  wire v3a6f7fd;
  wire v3a711b5;
  wire v3750d27;
  wire v373197c;
  wire v3726357;
  wire v3a70ec3;
  wire v376fb50;
  wire v37404bc;
  wire v3a70fec;
  wire v3768953;
  wire v374afa4;
  wire v3764aea;
  wire v3a6f2e7;
  wire v376ce15;
  wire v37601a1;
  wire v3a5dbd1;
  wire v3a70d93;
  wire v374657b;
  wire v3775721;
  wire v3a614d1;
  wire v376bfa7;
  wire v3a5cc77;
  wire v372ca99;
  wire v3750218;
  wire v3a6f5eb;
  wire v3a6f61c;
  wire v3a64641;
  wire v3a5965e;
  wire v377e2a4;
  wire v3a7159a;
  wire v3a628d4;
  wire v3775902;
  wire v38064a3;
  wire v373d64d;
  wire v3736be5;
  wire v374ffd5;
  wire v3757afc;
  wire v372bea3;
  wire v3a6fd19;
  wire v3a71551;
  wire v377dc8f;
  wire v3730289;
  wire v3a6cccd;
  wire v3739b38;
  wire v37526ca;
  wire v3740f9c;
  wire v37276a8;
  wire v373576f;
  wire v3729187;
  wire v3755220;
  wire v37627f6;
  wire v372e1b6;
  wire v37665c9;
  wire v37729bf;
  wire v3a610da;
  wire v3771646;
  wire v376c07e;
  wire v3577344;
  wire v3a5d30d;
  wire v3754e33;
  wire v372814c;
  wire v377a4ef;
  wire v3a5abf4;
  wire v372fbeb;
  wire v373f7ff;
  wire v39a4dac;
  wire v375789b;
  wire v373ccbc;
  wire v37c0339;
  wire v374eb71;
  wire v3756d07;
  wire v375045d;
  wire v3746303;
  wire v3a70f9f;
  wire v374f138;
  wire v372e3b4;
  wire v3753328;
  wire v377b170;
  wire v375b3b9;
  wire v37486d7;
  wire v375b031;
  wire v375d3e2;
  wire v3a65587;
  wire v3a59fbc;
  wire v377ab78;
  wire v376cf03;
  wire v3768d1d;
  wire v3749a29;
  wire v3742c16;
  wire v380761d;
  wire v372d924;
  wire v3779924;
  wire v3a64f5e;
  wire v37794e5;
  wire v3773107;
  wire v2092ff6;
  wire v376db98;
  wire v3a70f40;
  wire v375b776;
  wire v374179c;
  wire v3a70f29;
  wire v3a53e0e;
  wire db86c8;
  wire v3763dd5;
  wire v37577a4;
  wire v3a7049e;
  wire v3a67fee;
  wire v3a5d474;
  wire v3a5657a;
  wire v3724bbf;
  wire v3a6fcd3;
  wire v374c13e;
  wire v380700c;
  wire v3776649;
  wire v3a6a5e6;
  wire v375e431;
  wire v3751440;
  wire v3731c4b;
  wire v3a53cf5;
  wire v377329c;
  wire v372eb00;
  wire v374dcfb;
  wire v374a25d;
  wire v3a6f7db;
  wire v3a5cd0e;
  wire v3a6ef77;
  wire v3740aa8;
  wire v373bafb;
  wire v3a6f3d7;
  wire v373da11;
  wire v37304a2;
  wire v8455f1;
  wire v3749412;
  wire v37274a2;
  wire v376a27b;
  wire v39e9ca4;
  wire v8455f5;
  wire v3727e10;
  wire v3a5a260;
  wire v377b074;
  wire v3769759;
  wire v3a6fb85;
  wire v373eef9;
  wire v3730ab2;
  wire v329f8b7;
  wire v373aaca;
  wire v3a6ff57;
  wire v3778565;
  wire v37405a7;
  wire v3726dfa;
  wire v377eaf2;
  wire v3a6e432;
  wire v37559b2;
  wire v3759569;
  wire v3a71137;
  wire v3a6ac94;
  wire v372a023;
  wire v3778528;
  wire v3a7162d;
  wire v3753a3f;
  wire v3a6c0b3;
  wire v377f149;
  wire a36a2a;
  wire v3a670fe;
  wire v3a6006a;
  wire v375c9ea;
  wire v3a5dd17;
  wire v372f83b;
  wire v3a56d86;
  wire v3a6651d;
  wire v3a603a1;
  wire v3a71282;
  wire v3a712c0;
  wire v3a5c538;
  wire v374e78a;
  wire v3a6add2;
  wire v373d0b2;
  wire v375483e;
  wire v374cc2a;
  wire v3747c93;
  wire v3a5cf53;
  wire v3a6f418;
  wire v3a70fd2;
  wire v3770e30;
  wire v3a704b0;
  wire v373b51b;
  wire v374021a;
  wire v3743adf;
  wire v3a55198;
  wire v3a65e71;
  wire v374b42b;
  wire v3a6225d;
  wire v3a5a615;
  wire v377e81a;
  wire v3a61d1f;
  wire v373c8ac;
  wire v3729d06;
  wire v3725a0b;
  wire v1e37943;
  wire v3a6b58f;
  wire v3779c09;
  wire v3764955;
  wire v3779bde;
  wire v3a63dba;
  wire v3a58673;
  wire v373280e;
  wire v37408b7;
  wire v3a6af5b;
  wire v3734c16;
  wire v376aba9;
  wire v37269de;
  wire v3a58c2f;
  wire v37337b3;
  wire c7d478;
  wire v3a71579;
  wire v3a7136b;
  wire v373cbf9;
  wire v375e133;
  wire v377077a;
  wire v3770322;
  wire v3806b2d;
  wire v3a587a1;
  wire v372d811;
  wire v3a59eab;
  wire v3a5a3d0;
  wire v3a6f55c;
  wire v3738dac;
  wire v3731d76;
  wire v3a70467;
  wire v374a509;
  wire v3771440;
  wire v373e062;
  wire v377df1a;
  wire v3a6a0e4;
  wire v3778676;
  wire v3a6f7a7;
  wire v3742825;
  wire v3767c03;
  wire v374b424;
  wire v377c103;
  wire v377825c;
  wire v374a637;
  wire v374cd48;
  wire v3a60008;
  wire v375a41b;
  wire v377a5a9;
  wire v1e379ef;
  wire v37507dd;
  wire v374b340;
  wire v3766487;
  wire v377b981;
  wire v37496fc;
  wire v3a6f209;
  wire aac06c;
  wire v3779b31;
  wire v3747d0e;
  wire v3a712bc;
  wire v3a6fb20;
  wire v3a715f9;
  wire v373b1c8;
  wire v3742210;
  wire v3757ae7;
  wire v3739743;
  wire v37642a0;
  wire v375534a;
  wire v3a6f567;
  wire v3767c46;
  wire v37232a6;
  wire v3a7156a;
  wire v37433ef;
  wire ba7f1c;
  wire v3a66ca0;
  wire v3728867;
  wire v3747d42;
  wire v373dc53;
  wire v373ec29;
  wire v3a705da;
  wire v3776836;
  wire v3a62e99;
  wire v292555a;
  wire v374c88d;
  wire v3a706da;
  wire v3807a93;
  wire v38074ed;
  wire v3756fee;
  wire v3a70ec4;
  wire v3a70f25;
  wire c10173;
  wire v3742649;
  wire v37249fe;
  wire v3a6f63c;
  wire v376fbe3;
  wire v3763c39;
  wire v37366d5;
  wire v3761dda;
  wire v3767d57;
  wire v3755691;
  wire v3778857;
  wire v3a70423;
  wire v3a6f95a;
  wire v3a60d50;
  wire v373e01f;
  wire v3a705ee;
  wire v974eb9;
  wire v3a62bc6;
  wire v3775b2f;
  wire ca2eb2;
  wire v3750f77;
  wire v375e29b;
  wire v3a70461;
  wire v3754f72;
  wire v3729520;
  wire v373e365;
  wire d893c7;
  wire v3724023;
  wire v372862a;
  wire v37bfc97;
  wire v3775526;
  wire v3a5fa4c;
  wire v375a8a7;
  wire v3a647ce;
  wire v376eb3c;
  wire v377a366;
  wire v3806def;
  wire v376fc09;
  wire v3743ecf;
  wire v3a70879;
  wire v372a6de;
  wire v3741fee;
  wire v3a706a3;
  wire v3747d0a;
  wire v38074c0;
  wire v1e37e04;
  wire v3a6efc1;
  wire v3a6b768;
  wire v37285c9;
  wire v3a5cb2c;
  wire v3a6ae23;
  wire v3a6f467;
  wire v3a70739;
  wire v373a005;
  wire v3766232;
  wire v37681cc;
  wire v373fa48;
  wire v3a713b5;
  wire v372be74;
  wire v374b972;
  wire v37644ee;
  wire v376d258;
  wire v3a5d646;
  wire v3a700ff;
  wire v3a6f04d;
  wire v3a61516;
  wire v3758809;
  wire v373ff40;
  wire v3737c39;
  wire v3a6f078;
  wire v3770648;
  wire v3a5e3d3;
  wire v3725cbf;
  wire v3a558f6;
  wire v373d293;
  wire v3a55641;
  wire v377dacb;
  wire v3a6edbe;
  wire v3a70ae8;
  wire v3a67eb2;
  wire v3a712b5;
  wire v373beae;
  wire v3a60cf8;
  wire v37289d4;
  wire v3731115;
  wire v3a704bd;
  wire v3a6a4d4;
  wire v3a5b474;
  wire v3806ec2;
  wire v375f317;
  wire v372781d;
  wire v3729e5f;
  wire v3775d76;
  wire v3a6a493;
  wire v3a70ad6;
  wire v3725bab;
  wire v373a196;
  wire v373a305;
  wire aa52b8;
  wire v376646f;
  wire v3747931;
  wire v37409f4;
  wire v3773575;
  wire v376d8d1;
  wire v3a6f044;
  wire v374e3a9;
  wire v2092bcb;
  wire v374e085;
  wire v3763e76;
  wire v37771a8;
  wire v375b7b5;
  wire v374f351;
  wire v3a62e1b;
  wire v3a5ee6e;
  wire v375b90a;
  wire v3a62f13;
  wire v3a649fd;
  wire v3a6a934;
  wire v376a3bb;
  wire v376d6b2;
  wire v376be60;
  wire v3777abf;
  wire v37764c0;
  wire v375119e;
  wire v3759aca;
  wire v375d84e;
  wire v3a6f9bd;
  wire v3778bde;
  wire v375352f;
  wire v3762dcf;
  wire v3765bf4;
  wire v975066;
  wire v3727aa3;
  wire v94ea62;
  wire v3a5923c;
  wire v374d8cb;
  wire v375c31a;
  wire v3a6f4bc;
  wire v3759d78;
  wire v3770c66;
  wire v3757f45;
  wire v37657ef;
  wire v3759ee4;
  wire v3a67d4a;
  wire v37443b5;
  wire v3774f24;
  wire v3756a05;
  wire v375d559;
  wire v3807bf7;
  wire v373b78b;
  wire v3a70c7f;
  wire v3758915;
  wire v372f1b9;
  wire v3778546;
  wire v3a6c20e;
  wire v3a6f79e;
  wire v373397b;
  wire v39a4e43;
  wire v3a71064;
  wire v374dc53;
  wire v3755abd;
  wire v3759ef7;
  wire v3747c90;
  wire b96080;
  wire v3754565;
  wire v3a6fae9;
  wire v3726262;
  wire v1e37cba;
  wire v372d643;
  wire v3a5f33d;
  wire v3731d69;
  wire v3731906;
  wire v3a6fddd;
  wire v37562a5;
  wire v3a70e4b;
  wire v28896b4;
  wire v37445b9;
  wire v3a713c8;
  wire v3a712c4;
  wire v23fe159;
  wire v3770735;
  wire v3a6ffcc;
  wire v376112d;
  wire v373d69f;
  wire fc6f92;
  wire v374d451;
  wire v3a6fc6c;
  wire v2619ad0;
  wire v3731dc6;
  wire v3777787;
  wire v3a6772f;
  wire v3756971;
  wire v3a70b73;
  wire v3a5ae6d;
  wire v3a68523;
  wire v3a6ffcf;
  wire v376f3c8;
  wire v3747527;
  wire v377ba5a;
  wire v3a70752;
  wire v374a48c;
  wire v3a6e8d4;
  wire v373f492;
  wire v374af2f;
  wire v20930b8;
  wire v3a2a33d;
  wire v3757009;
  wire v3730052;
  wire v374586b;
  wire v3a6abcc;
  wire v3758d7e;
  wire v374f82e;
  wire v3a70fbf;
  wire v37780cc;
  wire v377190a;
  wire v37787ec;
  wire v377d33e;
  wire v3756261;
  wire v37481f3;
  wire v37231ed;
  wire v3a5d48b;
  wire v3749b84;
  wire v3a6fc64;
  wire v377b073;
  wire v372ae1b;
  wire bf3e2b;
  wire v3a71129;
  wire v3a7014e;
  wire v3a71078;
  wire v376711c;
  wire v3a6ec52;
  wire v95151c;
  wire v372cb44;
  wire v3a620d3;
  wire v37759b5;
  wire v37513bc;
  wire v3777e0e;
  wire v374f9ce;
  wire v3a56122;
  wire v3a6b4e8;
  wire v3770425;
  wire v3a70cee;
  wire v377c7d3;
  wire v3806b0a;
  wire v3a660af;
  wire v3a6f83a;
  wire v37787f5;
  wire v3a6eed9;
  wire v3a6ae0f;
  wire v3728ea6;
  wire v3747398;
  wire v37616e1;
  wire v3a6a7a1;
  wire v3728fb5;
  wire v337907e;
  wire v3806bc8;
  wire v372777c;
  wire v3a5cef4;
  wire v37507da;
  wire v376c4c5;
  wire v372c944;
  wire v3a70a87;
  wire v3a6134b;
  wire v377f70a;
  wire v3a6f8fd;
  wire v3726381;
  wire v373f0e6;
  wire v3806dda;
  wire v373e896;
  wire v8827d7;
  wire v373a18b;
  wire v3a6617b;
  wire v37354f8;
  wire v3a6fc78;
  wire v3a6946d;
  wire v3a66492;
  wire v37735ec;
  wire v3a583f5;
  wire v375a28a;
  wire v372600f;
  wire v37379d7;
  wire v3a702fe;
  wire v37686f6;
  wire v3a6e105;
  wire v1e37972;
  wire v377f73c;
  wire v3775c0b;
  wire v377b7f9;
  wire v377d2ee;
  wire v3757818;
  wire v3a5bd99;
  wire v3a6108b;
  wire v373497f;
  wire v3744a9c;
  wire v372a77f;
  wire v377e124;
  wire v373c059;
  wire v373e8b5;
  wire v3770f51;
  wire v38079d7;
  wire v372f16b;
  wire v375a677;
  wire v377d0fc;
  wire v374650c;
  wire v35b724a;
  wire v3770754;
  wire v3a710b2;
  wire v3724057;
  wire v377c31a;
  wire v373fbc7;
  wire v375d6ba;
  wire v3a6bf89;
  wire v3a5d36a;
  wire v376d312;
  wire v3a707a7;
  wire v3a6f08c;
  wire v3a68116;
  wire v3a69961;
  wire v3770b04;
  wire v3a70519;
  wire v374270c;
  wire v3a71478;
  wire v375f6e3;
  wire v3a69761;
  wire v3723f45;
  wire v375ab8e;
  wire v3735db2;
  wire v375c9bc;
  wire v373bb2f;
  wire v3a68601;
  wire v3378302;
  wire v377261b;
  wire v376ca13;
  wire v37605fb;
  wire v3a56b05;
  wire v3a6c050;
  wire v3a6f8d5;
  wire v377a8e0;
  wire v37445e5;
  wire v3a7020e;
  wire v3a5efb8;
  wire v373ac1c;
  wire v3a63fc5;
  wire v3a58a1b;
  wire v37362b5;
  wire v3a6f56c;
  wire v3737352;
  wire v3767aae;
  wire v3a55cc4;
  wire v3a70927;
  wire v3769a8e;
  wire v37609ab;
  wire v375c044;
  wire v37554a1;
  wire v3a6d3c5;
  wire v372fb48;
  wire v37283fe;
  wire v374e39c;
  wire v3a700c8;
  wire v23fdec8;
  wire v3737b63;
  wire v2acaeda;
  wire v3a5e3be;
  wire v3a57d9e;
  wire v376b8f8;
  wire v3758b89;
  wire v3a62015;
  wire v3a70e3f;
  wire v3744b07;
  wire v3807d59;
  wire v3a6f323;
  wire v37706a7;
  wire v3a6e8a6;
  wire v3a5db97;
  wire v3a70be7;
  wire v3726013;
  wire v3a6f061;
  wire v3a56f67;
  wire v3a71469;
  wire v3a66545;
  wire v3a7085f;
  wire v3a6a1b7;
  wire v37438ca;
  wire v3741d11;
  wire v37377fd;
  wire v37710ad;
  wire v3a6f55d;
  wire v373d5f0;
  wire v37300d3;
  wire v3a6df6c;
  wire v3733173;
  wire v3a70d78;
  wire v2092a89;
  wire v3753942;
  wire v3a62f8e;
  wire a7e544;
  wire v3a5e7e8;
  wire v3747ef9;
  wire v3761950;
  wire v3a633ca;
  wire v3762b55;
  wire v373f03e;
  wire v1e37b3f;
  wire v3742ac7;
  wire v372b5a3;
  wire v3751090;
  wire v3a7151e;
  wire v3a7018a;
  wire v3a6ad38;
  wire v375e2bc;
  wire v372e38f;
  wire v8ef654;
  wire v374bc3e;
  wire v3731cc3;
  wire v377ce51;
  wire v3731c1c;
  wire v376780f;
  wire v372e8cc;
  wire v374617d;
  wire v376a464;
  wire v373cd41;
  wire v3775252;
  wire v3a604bc;
  wire v35b71cf;
  wire v3a6f871;
  wire v372bfd0;
  wire v3777844;
  wire v3a5eaaf;
  wire v377d4de;
  wire v374514e;
  wire v374cf82;
  wire v3727026;
  wire v3739b17;
  wire v37289ee;
  wire v37277c3;
  wire v375d51e;
  wire v37278c8;
  wire v375b93d;
  wire v3752e46;
  wire v376fc98;
  wire v37383c0;
  wire v37470f6;
  wire v3a6fd63;
  wire v3753b3f;
  wire v3729b6a;
  wire v3a6403e;
  wire v373c7db;
  wire v372b858;
  wire v373e76a;
  wire v3809d45;
  wire v3a6f832;
  wire v372301d;
  wire v3730043;
  wire v3808cf1;
  wire v3a6eba3;
  wire v3a6ac66;
  wire v3a6f21c;
  wire v3759b7c;
  wire v3a68bf8;
  wire v3a7078a;
  wire v376b6c9;
  wire v3743eb5;
  wire b755d3;
  wire v375a00a;
  wire v3a6c449;
  wire v3806ec4;
  wire v3a59391;
  wire v3a6d9fa;
  wire v3740f92;
  wire v3a711e2;
  wire v3756eca;
  wire v37752c8;
  wire v372f1b8;
  wire v372aa99;
  wire v3a67284;
  wire v3a64e29;
  wire v37789a0;
  wire v3a644e6;
  wire v376ee03;
  wire v1e37721;
  wire v376c87d;
  wire v3731685;
  wire v23fe175;
  wire v37474dc;
  wire v3a5987a;
  wire v3a54560;
  wire v376d143;
  wire v376a094;
  wire v3809968;
  wire v374ca62;
  wire v3a6facd;
  wire v37528fd;
  wire v3768768;
  wire v372f3e8;
  wire v3a708e0;
  wire v376508b;
  wire v3a6c64d;
  wire v376f2c8;
  wire v3a6fb75;
  wire v3a70f38;
  wire v3a5b0a6;
  wire v3a6b288;
  wire v372cd1f;
  wire v3730f6f;
  wire v372a0cb;
  wire v3a6faf0;
  wire v3a6ac9e;
  wire v3766dfb;
  wire v3775b7e;
  wire v3754328;
  wire v3a6f6c6;
  wire v3758983;
  wire v3742ec5;
  wire v374f528;
  wire v3a5b28d;
  wire v3779c33;
  wire v3736aaa;
  wire v3a70cec;
  wire v3a62e42;
  wire v3a675d9;
  wire v3a533ae;
  wire v3748d17;
  wire v377c41b;
  wire v3a70ff8;
  wire v3775e03;
  wire v377d354;
  wire v3753c2a;
  wire v376693b;
  wire v37753da;
  wire v376b199;
  wire v377fc1f;
  wire v373ac71;
  wire v377d595;
  wire v37770af;
  wire v3a6fee5;
  wire v375fc79;
  wire v3772f37;
  wire v374f273;
  wire v377d45b;
  wire v3737c52;
  wire v372acd3;
  wire v376b1d4;
  wire v3a66349;
  wire v3a70f92;
  wire v373c26c;
  wire v375c924;
  wire v3747c20;
  wire v373e60c;
  wire v3779d96;
  wire v3a70cd7;
  wire v376a383;
  wire v372946a;
  wire v375d2b1;
  wire v377b267;
  wire v3a65130;
  wire v3730b3a;
  wire v374cf79;
  wire v3a56c2e;
  wire v3a6f0e9;
  wire v3730695;
  wire v374e353;
  wire v3759edb;
  wire v37454cc;
  wire v3764825;
  wire v375792f;
  wire v3745790;
  wire v374b6e8;
  wire v3746e10;
  wire v3a6f3a9;
  wire v3778f19;
  wire v373149a;
  wire v374312f;
  wire v3a68c87;
  wire v373f3ac;
  wire c47a78;
  wire v373340d;
  wire v37269f6;
  wire v3741ccb;
  wire v376efb6;
  wire v3a6f9d7;
  wire v3747238;
  wire v3773a00;
  wire v3a6f954;
  wire v3a70712;
  wire v376ed58;
  wire v3768a43;
  wire v3a6fa1d;
  wire v3a6ef07;
  wire v373fcc7;
  wire v377097e;
  wire v373e11e;
  wire v373fa73;
  wire v3735512;
  wire v377d21c;
  wire v374dabe;
  wire v3779810;
  wire v2ff87d7;
  wire v37457c1;
  wire v3738d63;
  wire v37520fc;
  wire v3a7161c;
  wire v3750b64;
  wire v373150d;
  wire v3a704cd;
  wire v3754aa8;
  wire v37451db;
  wire aa5585;
  wire v3a61796;
  wire v3731f35;
  wire v3779749;
  wire v3a70b10;
  wire v37751b4;
  wire v374132e;
  wire v3735ac0;
  wire v376edbb;
  wire v37235fa;
  wire v3743b63;
  wire v3734e70;
  wire v3a6ebee;
  wire v37774b6;
  wire v37484e7;
  wire v3764383;
  wire v3a573ec;
  wire v377d51d;
  wire v3a70207;
  wire v3a70bcb;
  wire v3755113;
  wire v3766746;
  wire v3a68356;
  wire v3762e54;
  wire v3a70c92;
  wire v377a3af;
  wire v3a6b303;
  wire v3728990;
  wire v377c9a1;
  wire v3a61724;
  wire v373d78f;
  wire v375047c;
  wire v372af95;
  wire v375c3c5;
  wire v38079db;
  wire v3a672b6;
  wire v3a6eff6;
  wire v372f744;
  wire v37477d5;
  wire v37500d0;
  wire v3a617ad;
  wire v3760989;
  wire v374fba1;
  wire v3740466;
  wire v3768e14;
  wire v377e071;
  wire v3764869;
  wire v3a6f5a4;
  wire v2092ac1;
  wire v3a6ec01;
  wire v3a715b8;
  wire v376079d;
  wire v3728840;
  wire v3729544;
  wire v3775a8e;
  wire v3766afa;
  wire v3732b92;
  wire v3a6fd4f;
  wire v3725ba5;
  wire v3772e4f;
  wire v3a5b01a;
  wire v372f1a8;
  wire v3748e6a;
  wire v3a6fcf5;
  wire v376cfc9;
  wire v37646ce;
  wire v3a551e2;
  wire v3a6724f;
  wire v3a5971d;
  wire v38064a1;
  wire v37736c4;
  wire v3a595fd;
  wire v3a6f551;
  wire v3743def;
  wire v3a658d5;
  wire v37723b7;
  wire v372790e;
  wire d62aa6;
  wire v3a6b37c;
  wire v375084d;
  wire v3769f84;
  wire v3a64056;
  wire v37591da;
  wire v37771ca;
  wire v3a6f105;
  wire v3a6b51b;
  wire v375aa6b;
  wire v376c2a1;
  wire v3750c27;
  wire v3a6f4df;
  wire v3a5bc77;
  wire v3749674;
  wire v3a66fb3;
  wire v3a5ba1a;
  wire v1e37413;
  wire v3a6f994;
  wire v3a60103;
  wire v377a180;
  wire v3779925;
  wire v3a70e70;
  wire v3754403;
  wire v3770da3;
  wire v3a68904;
  wire v3728c08;
  wire v3a6279b;
  wire v3a5f7c5;
  wire v3741e56;
  wire v373f14d;
  wire v3a6080b;
  wire a374cd;
  wire v3a70b56;
  wire v3768383;
  wire v3a61886;
  wire v3732797;
  wire v2092baa;
  wire v1e37bf6;
  wire v3765784;
  wire v374f7ec;
  wire v3727bcb;
  wire v37711dd;
  wire v372a068;
  wire v3a7106b;
  wire v3742723;
  wire v3a6d1fa;
  wire v3a635f8;
  wire v3776cce;
  wire v3a5fa22;
  wire v373cb58;
  wire v3723404;
  wire v37668cb;
  wire v3755a70;
  wire v3a6adb2;
  wire v3a7164a;
  wire v98381a;
  wire v3a5378e;
  wire v37602cf;
  wire v3730c26;
  wire v376f87a;
  wire v3a603ad;
  wire v1e37a72;
  wire v3a6ebae;
  wire v372452c;
  wire v375a6d3;
  wire v3742bc1;
  wire v374f7cb;
  wire v3a6ffc7;
  wire v377f85a;
  wire v372bf24;
  wire v37385d2;
  wire v3722d9b;
  wire v3a59caa;
  wire v3a5f587;
  wire v377215c;
  wire v3a70fb7;
  wire v3a6f100;
  wire v3a64dbb;
  wire v3a714a6;
  wire v3754107;
  wire v3750cfd;
  wire v37305e3;
  wire v377fbeb;
  wire v3a6a084;
  wire v3a7165e;
  wire v3a5b642;
  wire v3766f30;
  wire v3a7017f;
  wire v3a6feb5;
  wire v1e37b52;
  wire v372c18a;
  wire v372ebc8;
  wire v3a6054b;
  wire v3a6eafe;
  wire v373b1ae;
  wire v375c740;
  wire v3732899;
  wire v3749dc2;
  wire v3a70ffe;
  wire v375f069;
  wire v9bba04;
  wire v3a6f2d5;
  wire v377670f;
  wire v375ed52;
  wire v3a6bfea;
  wire v3a685cd;
  wire v3a6b381;
  wire v3759c90;
  wire v37744f5;
  wire v3745801;
  wire v3a6b4ae;
  wire v373541f;
  wire d9767c;
  wire v3a6f77c;
  wire v3743366;
  wire v376905f;
  wire v373a3dd;
  wire v3a6fdc5;
  wire v3775d56;
  wire v3a5770d;
  wire v3725582;
  wire v3a6f9b9;
  wire v373b6c0;
  wire v377ab46;
  wire v37412c3;
  wire v3723fce;
  wire v37667f7;
  wire v3a5b70a;
  wire v3a67a85;
  wire v3742af4;
  wire v8639e9;
  wire v3778bef;
  wire v3a6f887;
  wire v3760b03;
  wire v3737ace;
  wire v376fe90;
  wire v376f814;
  wire v3a6ecdd;
  wire v374d6ff;
  wire v3a596a5;
  wire v376592c;
  wire v373fb42;
  wire v3a5511c;
  wire v376b44a;
  wire v3a6b4de;
  wire v96ab98;
  wire v3748282;
  wire v377e73f;
  wire v373300a;
  wire v3745e5e;
  wire v3743f11;
  wire v377d7e1;
  wire v3775a7d;
  wire v3a6eee4;
  wire v3746cc5;
  wire v3725589;
  wire v921bc8;
  wire v3a70432;
  wire v374446c;
  wire v37435a0;
  wire v375000b;
  wire v3a70bde;
  wire v376acd5;
  wire v3758395;
  wire v3a58022;
  wire v374d011;
  wire v3a6126c;
  wire v3a70bd2;
  wire v97ecca;
  wire v373da5b;
  wire v3a5f4ff;
  wire v375bd53;
  wire v377a4c1;
  wire v3a57593;
  wire v373d40a;
  wire v37324bb;
  wire v3a6f6eb;
  wire v37739a8;
  wire v3a6ceb0;
  wire v3748cb7;
  wire v377052f;
  wire v3744796;
  wire v376a867;
  wire v3a6bab9;
  wire v376e16e;
  wire v3731415;
  wire v373f0a3;
  wire v375473a;
  wire v376abf6;
  wire v37664d0;
  wire v3a62d56;
  wire v373c2d7;
  wire v3a69169;
  wire v37420b6;
  wire v3a69267;
  wire v3741e82;
  wire v377f190;
  wire v3a65245;
  wire v3a53dff;
  wire v3a6c636;
  wire v357733c;
  wire v373aa3d;
  wire v3770ff4;
  wire v3729031;
  wire v37672af;
  wire v3a70ede;
  wire v373bc2f;
  wire v37314d7;
  wire v3760167;
  wire v3a70406;
  wire v375d98f;
  wire v3a6f650;
  wire v373b4ad;
  wire v3754903;
  wire v37293ea;
  wire v373cc0f;
  wire v3a6f490;
  wire v376ef09;
  wire v373e52d;
  wire v373fef5;
  wire v3a6ef90;
  wire v37606dc;
  wire v374dfd5;
  wire a2aef9;
  wire v3752dbb;
  wire v3a6fbf4;
  wire v3a6fb78;
  wire v3a62d36;
  wire v37535f2;
  wire v3a6fe8a;
  wire v3761031;
  wire v375a03b;
  wire cea55f;
  wire v377f27f;
  wire v377f669;
  wire v377bb56;
  wire v3776ace;
  wire v375c351;
  wire v372529a;
  wire v372e499;
  wire v3739e05;
  wire v360d01e;
  wire v37572eb;
  wire v3756bd2;
  wire v3779b96;
  wire v3767ba9;
  wire v3a70473;
  wire v3749293;
  wire v3a63621;
  wire v37306bb;
  wire v3806507;
  wire v37254c0;
  wire v3a70eb6;
  wire v37548d8;
  wire v373081f;
  wire v3a70bff;
  wire v3743c51;
  wire v3745c75;
  wire v375a38e;
  wire v37600e9;
  wire v3a62caa;
  wire v3737202;
  wire v3a62d5d;
  wire v3a538b3;
  wire v3a6ebb7;
  wire v3a712a3;
  wire v376d327;
  wire v3a70e84;
  wire v372b7b7;
  wire v3a6f613;
  wire v3723e1f;
  wire v3754777;
  wire v375b349;
  wire v3a62197;
  wire v376ffbf;
  wire v3a64e2a;
  wire v37270bc;
  wire v3750ad1;
  wire v3740c5f;
  wire v39372d9;
  wire v3779cf6;
  wire v3736eff;
  wire v37c36bf;
  wire v374c720;
  wire v3a6ff70;
  wire v3752616;
  wire v35b71fc;
  wire v372d3f1;
  wire v3765433;
  wire v374b0d9;
  wire v377e355;
  wire cbfab3;
  wire v374d612;
  wire v3a679fd;
  wire v3a5cf6f;
  wire v3745de0;
  wire v3a6be15;
  wire v376dcca;
  wire v374b274;
  wire v3762037;
  wire v3a708a4;
  wire v375d800;
  wire v37c03ad;
  wire v3a71375;
  wire v372d299;
  wire v3763548;
  wire v3770aee;
  wire v3a70119;
  wire v374f2d2;
  wire v3766f51;
  wire v3a6f1e8;
  wire v376d0b5;
  wire v3a55fe8;
  wire v3746df7;
  wire v376c7d1;
  wire v3732bf9;
  wire v374ad45;
  wire v3a6275e;
  wire v3761cd2;
  wire v3a64200;
  wire v3a5dff7;
  wire v373c7aa;
  wire v375c111;
  wire v3a6c2b2;
  wire v376978a;
  wire v37660d2;
  wire v377c6e8;
  wire v3766b81;
  wire v3a54f85;
  wire v3723903;
  wire v3a625c9;
  wire v376a272;
  wire v3a6f9ac;
  wire v3a70410;
  wire v3751dba;
  wire v3731eff;
  wire v3a6f69f;
  wire v37420e2;
  wire v3741218;
  wire v3a6fe52;
  wire v37495dc;
  wire ce69d1;
  wire v3a70d04;
  wire v3a6ead6;
  wire v3760088;
  wire v3a6f775;
  wire v3a6ffd0;
  wire v3735f79;
  wire v3766160;
  wire v3744f48;
  wire v376d98c;
  wire v3a6f70d;
  wire v372dc5c;
  wire v3a5dcfc;
  wire v375b7e1;
  wire v23fe101;
  wire v3730f35;
  wire v374733b;
  wire v3a6eba0;
  wire v373bd76;
  wire v3a5687e;
  wire v373cd68;
  wire v37775f9;
  wire v3a679e7;
  wire v372a79f;
  wire v3735fdc;
  wire v3741fc9;
  wire v3a6e91d;
  wire v3773b7b;
  wire v37540e7;
  wire v3a539bb;
  wire v3750d46;
  wire v3726505;
  wire v3a7102b;
  wire v372f553;
  wire v37328f1;
  wire v9ae4c2;
  wire v3725bba;
  wire v3a5c3eb;
  wire v3a641d5;
  wire v3a6d499;
  wire v37651c2;
  wire v372348c;
  wire v3a70716;
  wire v377b3df;
  wire v3762ca2;
  wire v3a6830c;
  wire v39a4e5f;
  wire v3a6d9c6;
  wire v374f35a;
  wire v3741694;
  wire v372f76a;
  wire v37551e3;
  wire v374944b;
  wire v3a6ffab;
  wire v377a1d3;
  wire v209300d;
  wire v23fdf30;
  wire v3736d43;
  wire v3a709f2;
  wire v376e5ab;
  wire v3a5b469;
  wire v374bae0;
  wire v3a66b2b;
  wire v3807a92;
  wire v373f0ee;
  wire v376be2c;
  wire v373502a;
  wire v374172f;
  wire v3742905;
  wire v3744877;
  wire v3748de3;
  wire v3a71615;
  wire d5ffe1;
  wire v376a0fc;
  wire v3a6ff2c;
  wire v373dbfe;
  wire v3722a46;
  wire v3a689bb;
  wire v375842f;
  wire v375d417;
  wire v3a650a6;
  wire v375aa47;
  wire a4a7a5;
  wire v37317a9;
  wire v3a710c2;
  wire v3a67aaa;
  wire v374c9f0;
  wire v3756c25;
  wire v3758f1b;
  wire v374d0f9;
  wire v3768723;
  wire v3a5c25e;
  wire v3a7137f;
  wire v3a6f2cb;
  wire v38072bd;
  wire v3775e78;
  wire v377c9cc;
  wire v377abcb;
  wire v377489e;
  wire v3a6fd2a;
  wire v376c8ea;
  wire v3a6fed3;
  wire v3a66051;
  wire v3a55bf6;
  wire v375b044;
  wire v3a69efa;
  wire v377b67d;
  wire v37570db;
  wire v3a612af;
  wire v3a61580;
  wire v3257acb;
  wire v3a6a9d7;
  wire v28896f0;
  wire v375a6e8;
  wire v373e1fb;
  wire v37533b4;
  wire v3a68d2e;
  wire v3a59aa1;
  wire v377744b;
  wire v3a69946;
  wire v376305d;
  wire v37541c6;
  wire v3730c86;
  wire v3731f7f;
  wire v39eb550;
  wire v3a5f602;
  wire v3a6ec0f;
  wire v3a6f7c6;
  wire v3760e1b;
  wire v37667eb;
  wire v1e37a9d;
  wire v376639f;
  wire v3767797;
  wire v3a656be;
  wire v375a86a;
  wire v3770ad8;
  wire v3a5a5a7;
  wire v374871a;
  wire v375bce7;
  wire v374457a;
  wire v3769f23;
  wire v3a5eefd;
  wire v3a6f417;
  wire v372d5e5;
  wire v372d28d;
  wire v377c5de;
  wire v3a6f47a;
  wire v3a60fee;
  wire v375c01e;
  wire v3a538ba;
  wire v3742a4e;
  wire v376c6b3;
  wire v374e8f7;
  wire v372b6b9;
  wire v373e225;
  wire v3a5cb14;
  wire v3738937;
  wire v3a6fb83;
  wire v3a5fefa;
  wire v3a70e98;
  wire v377504a;
  wire v372fff3;
  wire v1e37339;
  wire v374518c;
  wire v375ff94;
  wire v374f707;
  wire v3a70a4d;
  wire v3a70a18;
  wire v3a6603d;
  wire v373ccde;
  wire v3759b63;
  wire v373d076;
  wire v3776bdf;
  wire v3a70172;
  wire v372aec7;
  wire v3a6f501;
  wire v3761175;
  wire v3774e4f;
  wire d7669b;
  wire v3a6f528;
  wire v3a5acb3;
  wire v3a70317;
  wire v37366ed;
  wire v37671eb;
  wire v3742c6c;
  wire v376358f;
  wire v3a63a18;
  wire v3a6fd8f;
  wire v3a70244;
  wire v373dd4a;
  wire v23fd8cb;
  wire v3806ef3;
  wire v375f145;
  wire v374f712;
  wire v37512ca;
  wire v3a712ca;
  wire v37762bd;
  wire v3a5b071;
  wire v37507dc;
  wire v374d7ec;
  wire v3770072;
  wire v3734dd6;
  wire v3a546a2;
  wire v373b203;
  wire v3a6f5a2;
  wire v37437cf;
  wire v376dcbe;
  wire v3a568ee;
  wire v3750ba3;
  wire v37705ec;
  wire v3762ac3;
  wire v3759cb9;
  wire v376a06d;
  wire v3a6f6e8;
  wire v3a5d03e;
  wire v3761f4e;
  wire v3727823;
  wire v3741343;
  wire v3a6caa7;
  wire v3a5c0e1;
  wire v3731720;
  wire v3a5750b;
  wire v37773d6;
  wire v37385d3;
  wire v374c790;
  wire v372f5c5;
  wire v3a5a223;
  wire v3a709fb;
  wire v3a6bbe3;
  wire v3752dc7;
  wire v3a70f63;
  wire v3a64bb1;
  wire v376cba1;
  wire v37669d0;
  wire v377f6a5;
  wire v3a61f33;
  wire v3735d9e;
  wire v3734c26;
  wire v373dcd2;
  wire v3774c4d;
  wire v2889703;
  wire v3a70466;
  wire v3733dd8;
  wire v3752933;
  wire v3773e77;
  wire v3769e70;
  wire v3806f08;
  wire v3a57384;
  wire v3a5e647;
  wire v374518e;
  wire v3758661;
  wire v375aa18;
  wire v377638d;
  wire v3743798;
  wire v375c8db;
  wire v3749ae8;
  wire v3a7117d;
  wire v377aa4d;
  wire v3a70923;
  wire v3a65da2;
  wire v3a5ef89;
  wire db903b;
  wire v376bea3;
  wire v37371b2;
  wire v3a68954;
  wire v3754176;
  wire v377db14;
  wire v372c53a;
  wire v3a58527;
  wire v3a70feb;
  wire v375f9f1;
  wire v37499ac;
  wire v377e31d;
  wire ac8c4a;
  wire v373a36a;
  wire v3771431;
  wire v374868d;
  wire v3746a2b;
  wire v3770075;
  wire v3774df9;
  wire v3777eed;
  wire v3a63da7;
  wire v375a7d3;
  wire v376aa99;
  wire v373ee52;
  wire v3a668da;
  wire v3766acb;
  wire v3a54580;
  wire v3772e85;
  wire v3a7026d;
  wire v3a6f9e6;
  wire v3779593;
  wire v372fdd0;
  wire v3a712f5;
  wire v376e507;
  wire v3773b66;
  wire v3a646fb;
  wire v37649d3;
  wire v376f23f;
  wire v3762656;
  wire v377c079;
  wire v3a67833;
  wire v3a6e6fa;
  wire v372cea0;
  wire v3a6fb7f;
  wire v3a70613;
  wire v3733e1f;
  wire v3a65755;
  wire v37441a3;
  wire v37734d2;
  wire v37712c2;
  wire v3a71227;
  wire v3a6f53e;
  wire v37445f1;
  wire v374ad30;
  wire v373a341;
  wire v3770d41;
  wire v3a7136a;
  wire v374e6e3;
  wire v374ba05;
  wire v372e132;
  wire v3725556;
  wire v3a6efad;
  wire v3a6872e;
  wire v373a6c8;
  wire v373fde6;
  wire v2acaed3;
  wire v3779c2b;
  wire v375c98d;
  wire v3774bdf;
  wire v377e9a5;
  wire v37710a1;
  wire v869938;
  wire v3740bee;
  wire v375c0e8;
  wire v3767a7b;
  wire v3766877;
  wire v3809b31;
  wire v37450b8;
  wire v3a6f4d2;
  wire v375da9c;
  wire v37233e7;
  wire v3a7024c;
  wire v373ff1c;
  wire v3a697e4;
  wire v3758299;
  wire v3a707ce;
  wire v375abab;
  wire v3a5899d;
  wire v37c0158;
  wire v375f370;
  wire v3a59f9b;
  wire v372c134;
  wire v37250a3;
  wire v3773c69;
  wire v3a70d64;
  wire v374dd61;
  wire v37474b8;
  wire v376cc1b;
  wire v3766117;
  wire v373bb2c;
  wire v3a630dc;
  wire b3d3ad;
  wire v375e577;
  wire v3a6f0fd;
  wire v37685ea;
  wire v3736c8d;
  wire v375cdf4;
  wire v375c4ac;
  wire v373bda7;
  wire v377f104;
  wire v3758869;
  wire v3a6fbd1;
  wire v3727c07;
  wire v3a70ef8;
  wire v377b2f3;
  wire v3775687;
  wire v3a59085;
  wire v3a6015c;
  wire v3730789;
  wire v3a71326;
  wire v377f5f2;
  wire v3a66632;
  wire v376b193;
  wire v3a6f9cb;
  wire v377d004;
  wire v3a6c8b0;
  wire v3a6f6fe;
  wire v3a5bed2;
  wire v38065f1;
  wire v3a59ddc;
  wire v3a615c7;
  wire v3746aa9;
  wire v374ace9;
  wire v3a70307;
  wire v37618bf;
  wire v372f0bc;
  wire v3757ad8;
  wire v37790a6;
  wire v3a563cf;
  wire v3a6bedd;
  wire v372f464;
  wire v3a69677;
  wire v374749d;
  wire v3a6087b;
  wire v37553f5;
  wire v3748e09;
  wire v3a6f38b;
  wire v3747fbf;
  wire v23fda4e;
  wire v373eb03;
  wire v3a61132;
  wire v3722b64;
  wire v3751f72;
  wire cf45c3;
  wire v373a493;
  wire v37302c5;
  wire v377d1ab;
  wire v3749008;
  wire v3764c9c;
  wire v3750adf;
  wire v3a6f676;
  wire v3747a0e;
  wire v3727580;
  wire v3a5fc82;
  wire v372eb1a;
  wire v37333bb;
  wire v37393ed;
  wire v3759d41;
  wire v372f07d;
  wire v376d72e;
  wire v372a161;
  wire v373e16b;
  wire v3754a74;
  wire v3a7152f;
  wire v3725380;
  wire v3378a34;
  wire v374a430;
  wire v3a61d2e;
  wire v3a6efea;
  wire v3757254;
  wire v373abae;
  wire v376b2a2;
  wire v3a56cca;
  wire v375a635;
  wire v377ad76;
  wire v360d166;
  wire v3a710eb;
  wire v3757407;
  wire v374aece;
  wire v373b9d6;
  wire v376d4ee;
  wire v3a6ae3e;
  wire v3a6f9a2;
  wire v3755a05;
  wire v3a70186;
  wire v377221f;
  wire v3737681;
  wire v3a58038;
  wire v3a7116e;
  wire v3759536;
  wire v3a710ad;
  wire v3a6afef;
  wire v375c52f;
  wire v3a5784f;
  wire v3775636;
  wire v3a6f8d0;
  wire v374d4d3;
  wire v3768904;
  wire v2093083;
  wire v373d43a;
  wire v3a6ac33;
  wire v37551c4;
  wire cb09e1;
  wire v37559c4;
  wire v375f963;
  wire v3a571fa;
  wire v3a6fb73;
  wire v3724028;
  wire v37440c0;
  wire v374ad17;
  wire v3a5c196;
  wire v374b074;
  wire v3a6fdf5;
  wire v373aa0e;
  wire v3769a6c;
  wire v3a6bba4;
  wire v374ffb8;
  wire v3737265;
  wire v37343f6;
  wire v3749336;
  wire v3a71574;
  wire v3a5d217;
  wire v3764761;
  wire v38095b1;
  wire v376fbfd;
  wire v3737200;
  wire v3a70040;
  wire v376c313;
  wire v372c41f;
  wire v325c90f;
  wire v372668c;
  wire v3a2a911;
  wire v3771428;
  wire v376c8f2;
  wire v376f42c;
  wire v37664b4;
  wire v3a6f625;
  wire v3a66a4f;
  wire b4ede7;
  wire v3776974;
  wire v3728e91;
  wire v3776c6b;
  wire v3a6f9ff;
  wire v373100d;
  wire v3744d54;
  wire v3a6329a;
  wire v3755207;
  wire v3731994;
  wire v374b0a3;
  wire v3a6f474;
  wire v377386a;
  wire v3a555a9;
  wire v3a60223;
  wire v372cb36;
  wire v372a460;
  wire v3a6f86a;
  wire v3a698ab;
  wire v3730402;
  wire v3754cb0;
  wire v3a69fde;
  wire v3a6fb69;
  wire v37560f1;
  wire v37675e9;
  wire v373ba2e;
  wire v374975c;
  wire v3a55491;
  wire v3a6fec6;
  wire v372ce94;
  wire v372b646;
  wire v372f0e0;
  wire v3a67c30;
  wire v3732b1d;
  wire v37563ef;
  wire b9d061;
  wire v3a611d8;
  wire v3774d6e;
  wire v373cb89;
  wire v3a6f4b9;
  wire v3a5ed98;
  wire v37558d3;
  wire v3750375;
  wire v3a299f3;
  wire v3a7016e;
  wire v374c5f6;
  wire v3a6b9d9;
  wire v372a8fd;
  wire v3a6f6e2;
  wire v372c08d;
  wire v3774359;
  wire v3a63c8e;
  wire v3761026;
  wire v372db12;
  wire v37240c8;
  wire v3738a94;
  wire v3772b81;
  wire v360d105;
  wire v3a6678b;
  wire v375c8c8;
  wire v3734868;
  wire v3751fbe;
  wire v3a5b7e3;
  wire v3a648a6;
  wire v3a6f194;
  wire v3779b12;
  wire v3753e28;
  wire v374e5e9;
  wire v372cb77;
  wire v3a58ba8;
  wire v37772db;
  wire v37327ee;
  wire v3746ef3;
  wire v3760464;
  wire v377c6ce;
  wire v3731dfe;
  wire v3764910;
  wire v3a5b912;
  wire v3a6d0af;
  wire v3751261;
  wire v37579f7;
  wire v3727c74;
  wire v3767b5a;
  wire v3779097;
  wire v3773c13;
  wire v3a716a2;
  wire cfe9c3;
  wire v360c1bf;
  wire v376ba89;
  wire v37648cd;
  wire v3736afd;
  wire v3a5e620;
  wire v372c85f;
  wire v3a57c0d;
  wire v3a7138c;
  wire v3776779;
  wire v3a6332f;
  wire v377c798;
  wire v375aa99;
  wire v3736af1;
  wire v3722b6f;
  wire v3807413;
  wire v3a701f7;
  wire v37783d2;
  wire v3754fc6;
  wire v3743522;
  wire v3a63306;
  wire v374dd4c;
  wire v37316cb;
  wire v37410dc;
  wire v3742f76;
  wire v3a66c94;
  wire v3774f1e;
  wire v3736515;
  wire v372f2ed;
  wire v3727363;
  wire v3a7008f;
  wire v3722b21;
  wire v3744c5e;
  wire v373c228;
  wire v3a704fb;
  wire v37281be;
  wire v3a6f58f;
  wire v3a5e7e0;
  wire v3a70175;
  wire v37328fc;
  wire v3734c20;
  wire v3729a1c;
  wire v37445d7;
  wire v3a6f430;
  wire v3a6fa5c;
  wire v3a6a374;
  wire v3739cfb;
  wire v376e02e;
  wire v37504a9;
  wire v3a70480;
  wire v8e6c5f;
  wire v3724715;
  wire v3a54811;
  wire v374af22;
  wire v372efee;
  wire v37548f5;
  wire v3a6de4f;
  wire v3a59649;
  wire v3728903;
  wire v3a5dc67;
  wire v374dbf7;
  wire v37523e9;
  wire v372ff3a;
  wire v37255a7;
  wire v374e9c0;
  wire v3761466;
  wire v2acae4c;
  wire v3a58dce;
  wire v3a710c8;
  wire v375a4eb;
  wire v373029d;
  wire v3743f54;
  wire v3769302;
  wire v3a6898d;
  wire v37688df;
  wire v3732d82;
  wire v3a707ea;
  wire v3a685c7;
  wire v3807513;
  wire v3a70126;
  wire v3a67b48;
  wire v3745a81;
  wire v3764270;
  wire v3a70f28;
  wire v3743fe3;
  wire v3a66316;
  wire v3a5e371;
  wire v373e93e;
  wire v3a60229;
  wire v377ce5e;
  wire v3752321;
  wire v3742a4b;
  wire v3729933;
  wire v375df8e;
  wire v3a707ec;
  wire v3a70da4;
  wire v37404d0;
  wire v3743165;
  wire v3759172;
  wire v3744a91;
  wire v3255b53;
  wire v3a5d3f6;
  wire v3a557d2;
  wire v374bd4a;
  wire v3728870;
  wire v3747598;
  wire v3a579e2;
  wire v3a6f91b;
  wire v3a70510;
  wire v3754164;
  wire v3760644;
  wire v37564d1;
  wire v3767e7f;
  wire v3722b91;
  wire v3757dc4;
  wire v373bbe6;
  wire v3a6abfe;
  wire v3a707e1;
  wire v3808d56;
  wire v3740681;
  wire v3a6fbdb;
  wire v3735c84;
  wire v3724cce;
  wire v3a710ff;
  wire v374159f;
  wire v3a6eef8;
  wire v3766846;
  wire v375e4d9;
  wire v37662d7;
  wire v37645aa;
  wire v3741e9d;
  wire v3730da3;
  wire v3770af1;
  wire v377c6b3;
  wire v37518fa;
  wire v3377af7;
  wire v3a590fb;
  wire v37526d6;
  wire v375d4d9;
  wire v37572f7;
  wire v3a6fba9;
  wire v375add0;
  wire v3744452;
  wire v33789b9;
  wire v3a6fcfd;
  wire v3754379;
  wire v3774d86;
  wire v37759a7;
  wire v372afcc;
  wire ca50c0;
  wire v3a6f750;
  wire v3741b61;
  wire v23fdf14;
  wire v375d5e1;
  wire v3731579;
  wire v3776ce0;
  wire v377b8b9;
  wire v29256bb;
  wire v375b261;
  wire v374d8bb;
  wire v3a6a322;
  wire v3a6eb1e;
  wire v377338f;
  wire v3a70261;
  wire v3a55d3b;
  wire v3a5f8a2;
  wire v3743fba;
  wire v3731d8f;
  wire v360bedd;
  wire v35b73a5;
  wire v3a55ab6;
  wire v3a630bc;
  wire v375f86d;
  wire v3743f9a;
  wire v8b32e5;
  wire v3a70cd2;
  wire v3807c0c;
  wire v37611b7;
  wire v375cf36;
  wire v3726777;
  wire v3a5eafa;
  wire v3773043;
  wire v377d41d;
  wire v37577db;
  wire cb1cc0;
  wire v374a115;
  wire v3a6ff8f;
  wire v373593a;
  wire v3a70321;
  wire v377b292;
  wire v3750866;
  wire v3258db3;
  wire v37719f2;
  wire v374ba04;
  wire v3a59dab;
  wire v3a552f7;
  wire v374a67d;
  wire v377a3ec;
  wire v377ca49;
  wire v3a70761;
  wire v372b794;
  wire v3a67c3b;
  wire v3760bda;
  wire v3a714c8;
  wire v3a56794;
  wire v3734cce;
  wire v373abcf;
  wire v3770f56;
  wire v3a70434;
  wire v3768d56;
  wire v3779cb1;
  wire v3a54eae;
  wire v373d993;
  wire v3742303;
  wire v3a70c69;
  wire v38064d5;
  wire v373edf3;
  wire v35b7033;
  wire v372c492;
  wire v375320f;
  wire v37353d9;
  wire v3734a99;
  wire v3770f7a;
  wire v3762434;
  wire v3a6ff8a;
  wire v372dfbe;
  wire v374e5e4;
  wire v3a60f85;
  wire v37744c1;
  wire v3a6d810;
  wire v3a5a2e2;
  wire v3a68f4d;
  wire v3a702b5;
  wire v3744d36;
  wire d57388;
  wire v3727b4a;
  wire v38099a1;
  wire v3a5bd05;
  wire v3a6f8ee;
  wire v3a5d678;
  wire v374882c;
  wire v377af11;
  wire v3a584d6;
  wire v3736a75;
  wire v373375c;
  wire v3723227;
  wire v3762b32;
  wire v372dd4b;
  wire v3734a80;
  wire v376739e;
  wire v3763105;
  wire v3a6fb6a;
  wire v3770174;
  wire v3a5f451;
  wire v3a7013a;
  wire v3a6f573;
  wire v37702dc;
  wire v3a700ef;
  wire v372a2ff;
  wire v3a6f0f3;
  wire v373867a;
  wire v3a5730e;
  wire v2ff8e3d;
  wire v3a707b4;
  wire v3a6ef1e;
  wire v372d078;
  wire v376e90a;
  wire v374355d;
  wire v372b89e;
  wire v3a68ed1;
  wire v3763d77;
  wire v3a5f83c;
  wire v3a69b93;
  wire v3a5bbec;
  wire v3753258;
  wire v3a5e846;
  wire v377629f;
  wire v374ffb7;
  wire v373785d;
  wire v3a70a4f;
  wire v3a6fab9;
  wire v3a56b4e;
  wire v3a70130;
  wire v376eaca;
  wire v37621ea;
  wire v3760ff4;
  wire v37761cb;
  wire v3a5dc82;
  wire v373f6d5;
  wire v3a70322;
  wire v372b8d7;
  wire v3769c7f;
  wire v3731d67;
  wire v374c6ff;
  wire c86567;
  wire v3769820;
  wire v3a61323;
  wire v3a60755;
  wire v3a68245;
  wire v3a711de;
  wire v373a68a;
  wire v37592ca;
  wire v3752147;
  wire v3a6f1f8;
  wire v3736028;
  wire v3a5b451;
  wire v375b9c1;
  wire v3a6972b;
  wire v23fd923;
  wire v3745039;
  wire v3a7025f;
  wire v3a66773;
  wire v37615aa;
  wire v9762fd;
  wire v3733b4e;
  wire v3a65a24;
  wire v3a590de;
  wire v3a6fbed;
  wire v374732a;
  wire v9c4c8d;
  wire v3755665;
  wire v3a6e21a;
  wire v3a5af1e;
  wire v3a707aa;
  wire v376fc77;
  wire v3a5f580;
  wire v3747ad6;
  wire v3764cea;
  wire v372e58c;
  wire v377d6fc;
  wire v3a6f27d;
  wire v372e5fb;
  wire v373b9ab;
  wire v37596df;
  wire v3a70c6c;
  wire v3a6f4cb;
  wire v372ab06;
  wire v37741f1;
  wire v3a6fa04;
  wire v3754ce8;
  wire v372f885;
  wire v38097c0;
  wire cf8423;
  wire v3a66811;
  wire v375a543;
  wire v372c28d;
  wire v3a6f068;
  wire v37591f2;
  wire v37597fa;
  wire v373c126;
  wire v375967d;
  wire v377167c;
  wire v3724c63;
  wire v372d866;
  wire v3753f1d;
  wire v3a71687;
  wire v375d886;
  wire v3a587dd;
  wire v3a6f0c6;
  wire v3731be2;
  wire v373bb6c;
  wire v376ea5c;
  wire v3731e0e;
  wire v3a6f7b4;
  wire v3731bd7;
  wire v3762712;
  wire v376cd8f;
  wire v3733480;
  wire v3a6f2bb;
  wire v37288b6;
  wire v372e83f;
  wire v372d608;
  wire v372d7a4;
  wire v373e3d5;
  wire v3a61901;
  wire v374e43a;
  wire v1e3799d;
  wire v3a7139e;
  wire v37468ea;
  wire v3740dcd;
  wire v3a6e222;
  wire v8716e3;
  wire v3a5b7b9;
  wire v375ad94;
  wire v3a54455;
  wire v3749e13;
  wire v373df13;
  wire v3a6f60d;
  wire v3764141;
  wire v37696b6;
  wire v3a61c45;
  wire v3a6243f;
  wire v375d8e0;
  wire v3a54919;
  wire v3767892;
  wire v3778430;
  wire bf29af;
  wire v1e37ca4;
  wire v374fe7b;
  wire v375f9df;
  wire v3733132;
  wire v3778390;
  wire v372e618;
  wire v3a6c6f6;
  wire v3746145;
  wire v3770e35;
  wire v3a7144a;
  wire v3a6f709;
  wire v375c3a2;
  wire v3736bcd;
  wire v3767d14;
  wire v3744ff3;
  wire v3735485;
  wire v3a7086d;
  wire v3a71135;
  wire v3727e58;
  wire v375329c;
  wire v375e767;
  wire v37364bd;
  wire v376773a;
  wire v37774c7;
  wire v374e16a;
  wire v3a70c74;
  wire v3a711fb;
  wire v377881b;
  wire v3a70a4c;
  wire v3a6cf19;
  wire v3774209;
  wire v3a5b8e4;
  wire v3a6dd7e;
  wire v376480c;
  wire v3a70dfb;
  wire v37246f1;
  wire v337859c;
  wire v37699f2;
  wire v37711e1;
  wire v37638ee;
  wire v372eeee;
  wire v38097ca;
  wire v3761a96;
  wire v3a70ed9;
  wire v372ce45;
  wire v3764418;
  wire v3a60976;
  wire v3736217;
  wire v377cd7e;
  wire v37715d9;
  wire v3743f3c;
  wire v337902c;
  wire v375138c;
  wire v37390d6;
  wire v942053;
  wire v3a712d4;
  wire v3722a6f;
  wire v3756305;
  wire v3759bf4;
  wire v377982c;
  wire v23fe1ad;
  wire v3a70b63;
  wire v3a6ff16;
  wire v3a5ae05;
  wire v376984d;
  wire v377772d;
  wire v375c9b9;
  wire v37249ff;
  wire v37655bf;
  wire v375523e;
  wire v374d6f6;
  wire v3773a96;
  wire v3758b56;
  wire v3a71492;
  wire v3a6cd48;
  wire v37455ff;
  wire v3771c5f;
  wire v374e6c7;
  wire v1e379c4;
  wire v3a704f0;
  wire v3772b8a;
  wire v377b3a2;
  wire v3730c0b;
  wire v3a66274;
  wire v374674d;
  wire v3a703aa;
  wire v37707db;
  wire v3a6f6bf;
  wire v3a6f791;
  wire v3748299;
  wire v377e547;
  wire v3a5a884;
  wire v374b0e3;
  wire v376959b;
  wire v3a70fb1;
  wire v374b364;
  wire v372b3b6;
  wire v3a5b945;
  wire v373c553;
  wire v3a70b11;
  wire v3a57210;
  wire v373578f;
  wire v373b288;
  wire v3a706c0;
  wire v37722cc;
  wire v37567c7;
  wire v376485c;
  wire v373e296;
  wire aebd68;
  wire v884deb;
  wire v3a6f659;
  wire v376d9aa;
  wire v372a39d;
  wire v372c5da;
  wire v372ff9a;
  wire v3723fcc;
  wire v3725c41;
  wire v3776039;
  wire v3a6d64e;
  wire v377451f;
  wire v377d839;
  wire v3a5ba93;
  wire v3a56687;
  wire v3a5ab7b;
  wire v3a69923;
  wire v3743a4c;
  wire v377d15d;
  wire v37513e6;
  wire v3768737;
  wire v3a70459;
  wire v3a70378;
  wire v3a6f757;
  wire v377ac8a;
  wire v3725c68;
  wire v377542e;
  wire v374956a;
  wire v37559ea;
  wire v373eecc;
  wire v375a92b;
  wire v39eb56c;
  wire v375c728;
  wire v3749437;
  wire v3a70a6e;
  wire v374f3ad;
  wire v3744c08;
  wire v3770db8;
  wire v377857d;
  wire v3a6eecd;
  wire v3751dc9;
  wire v374d480;
  wire v37574d2;
  wire v3729f05;
  wire v3a614cb;
  wire v3a70e97;
  wire v3a68310;
  wire v9a2413;
  wire v373cf9c;
  wire v3a5b87f;
  wire v3a70dcb;
  wire v376aae5;
  wire v3a5b7ad;
  wire v3a70106;
  wire v3723b33;
  wire v33789d0;
  wire v3764461;
  wire v3733294;
  wire v3809964;
  wire v3a6eb69;
  wire v377d428;
  wire v3a6bb47;
  wire v3754295;
  wire v372586f;
  wire v3757e40;
  wire v3777bf4;
  wire v2ff8bbc;
  wire v3a594fe;
  wire v37706ae;
  wire v372e711;
  wire v3a6fb57;
  wire v3a5e783;
  wire v37576e7;
  wire v3806599;
  wire v377f5ca;
  wire v3a71146;
  wire v377c2bc;
  wire v3a70fea;
  wire v373f2fe;
  wire v374178a;
  wire v3a60c49;
  wire v3a70d38;
  wire v37625ef;
  wire v3a6fa4c;
  wire v3755738;
  wire v3a5b86c;
  wire v3a69583;
  wire v3a56e03;
  wire v375d997;
  wire v3a6f7d5;
  wire v3769ce7;
  wire v375bb51;
  wire v3a6f959;
  wire v374a157;
  wire v3a6c044;
  wire v3a714f1;
  wire v374b19b;
  wire v3a5de5f;
  wire v37582e0;
  wire v3731370;
  wire v2092f2c;
  wire v3a6fa10;
  wire v374fef0;
  wire v3747302;
  wire v3743b9e;
  wire v37496fa;
  wire v3a6a195;
  wire v373dd8a;
  wire v37416b5;
  wire v37408a3;
  wire v380693e;
  wire v3a71452;
  wire v3a62fa3;
  wire v3a598a0;
  wire v376e041;
  wire v3a68463;
  wire v3a6f20d;
  wire v372d4de;
  wire v3a68f98;
  wire v3808dd8;
  wire v3a6f9c7;
  wire v373ca1a;
  wire v3a6f4c7;
  wire v3a62965;
  wire v3a67eec;
  wire v37370f8;
  wire v3755a0f;
  wire v3776125;
  wire v377ec08;
  wire v373e521;
  wire v37458dc;
  wire v372310a;
  wire v3726e81;
  wire v3753bb2;
  wire v3a67cff;
  wire v3736cb8;
  wire v37239ed;
  wire v3736e06;
  wire v37692c1;
  wire v3778b8d;
  wire v373c2ec;
  wire v375da82;
  wire v373087b;
  wire v375cfa5;
  wire v1e37e67;
  wire v3778a76;
  wire v377d042;
  wire v3770719;
  wire v373185b;
  wire v3a5e4e5;
  wire v376f0f6;
  wire v3a6f81b;
  wire v374851a;
  wire v3774ab8;
  wire v3a6eb67;
  wire v3748d67;
  wire v377e298;
  wire v373b7c5;
  wire v3725717;
  wire v37458ca;
  wire v37790c8;
  wire v372bd46;
  wire v360d03f;
  wire v375039e;
  wire v375da10;
  wire v3753163;
  wire v376f768;
  wire v3a700b5;
  wire v3a70f74;
  wire v3a6939d;
  wire v3a654c1;
  wire v37577b6;
  wire v3729785;
  wire v3751a86;
  wire v37786a6;
  wire v3776865;
  wire v376f2a7;
  wire v3735ad2;
  wire v3a71582;
  wire v3a5dc35;
  wire v375a8ad;
  wire v376362f;
  wire v3a70c35;
  wire v3a6e985;
  wire v37339f0;
  wire v3a59d9d;
  wire v37276eb;
  wire v3762502;
  wire v3a5cd50;
  wire v375d689;
  wire v3a6ddd4;
  wire v3a6eead;
  wire v376533e;
  wire v3a5408c;
  wire v3744ae4;
  wire v375200e;
  wire v3726c36;
  wire v3a5f265;
  wire v372f8c1;
  wire v3771d77;
  wire v3767cfb;
  wire v3778fec;
  wire v373bf4f;
  wire v37285ad;
  wire v3a71037;
  wire v3a57ac7;
  wire v374d2e5;
  wire v374b6ac;
  wire v3751081;
  wire v3a59bbd;
  wire v3a6eb1c;
  wire v376a44f;
  wire v3a702a2;
  wire d54152;
  wire v3a6e7ed;
  wire v35b85ad;
  wire v37711f0;
  wire v376bb26;
  wire v3a7097d;
  wire v3a5f1d4;
  wire v3a709ef;
  wire v3a5bb64;
  wire v3770cb8;
  wire v3a707b2;
  wire v3757a04;
  wire v377a422;
  wire v337905c;
  wire v3a6fb0e;
  wire v376fc7f;
  wire v377cd41;
  wire v37667d3;
  wire v94b9e7;
  wire v374a89b;
  wire v3753f0d;
  wire v3809a58;
  wire v377b330;
  wire v3a7022c;
  wire v3a7161b;
  wire v3800eea;
  wire v2925d03;
  wire v3a70f09;
  wire v3a6b27d;
  wire v37774ca;
  wire v377e056;
  wire v375d434;
  wire v3753231;
  wire v372f6d3;
  wire v3a6c81d;
  wire v37487a6;
  wire v3770d22;
  wire v373d8ec;
  wire v3774e32;
  wire v3733da4;
  wire v374fe9d;
  wire v3a6fd98;
  wire v3747084;
  wire v377a18b;
  wire v39a4e99;
  wire v3a6f1b9;
  wire v373804d;
  wire v3a670e9;
  wire v3a58d6b;
  wire v3a70213;
  wire v3a6eb7b;
  wire v380909e;
  wire v3a703bf;
  wire v372b4cb;
  wire v3769923;
  wire v372c3c7;
  wire v374db6a;
  wire v38073bb;
  wire v3a70230;
  wire v372f346;
  wire v376132a;
  wire v3a703d7;
  wire v37581cf;
  wire v376a4ec;
  wire v37320ff;
  wire v3735796;
  wire v3a6f138;
  wire v37662e7;
  wire v3a58378;
  wire v37716ca;
  wire v3a66c5b;
  wire v374bd09;
  wire v3767e71;
  wire v3742ca7;
  wire v3739748;
  wire v3a70dbb;
  wire v37330dc;
  wire v28896dc;
  wire v374b23d;
  wire v374f9c6;
  wire v3a6452e;
  wire v3a67b76;
  wire v37385c6;
  wire v374bb76;
  wire v37418dc;
  wire v3775fa5;
  wire v3a65847;
  wire v37558f2;
  wire v3772a57;
  wire v3a6f4da;
  wire v3a63ac4;
  wire v373b0f3;
  wire v376c69d;
  wire v374deba;
  wire v37761dd;
  wire v37435eb;
  wire v3769f4e;
  wire v374bece;
  wire v375e037;
  wire v3748cd9;
  wire v3a6f224;
  wire v3a69329;
  wire v3734ba4;
  wire v372c3c0;
  wire v3a624e7;
  wire v3773633;
  wire v37392e0;
  wire v373b6ee;
  wire v3739f1d;
  wire v373fe0d;
  wire v3a6fdd7;
  wire v376597e;
  wire v3775622;
  wire v37525c5;
  wire v3a7025c;
  wire v3757253;
  wire v3a70a7f;
  wire v2acaffd;
  wire v3a6f03f;
  wire v373698b;
  wire v376992a;
  wire v3743604;
  wire v3759f23;
  wire v3730d34;
  wire v3a5af28;
  wire v23fd9f9;
  wire v3a6f2d8;
  wire v3a64709;
  wire v3730b15;
  wire v374a806;
  wire v3777142;
  wire v3a5f80f;
  wire v373a8a1;
  wire v3a675eb;
  wire v375cfd9;
  wire v376d4d9;
  wire v3a5a3be;
  wire v373128b;
  wire v3757d20;
  wire v3736901;
  wire v3a6224d;
  wire v374d7c1;
  wire cff2df;
  wire v3777daa;
  wire v23fe27f;
  wire v373cdea;
  wire v3770e95;
  wire v3a60ab2;
  wire v3764c7c;
  wire v3806498;
  wire v376dd64;
  wire v374fa18;
  wire v3738087;
  wire v373b667;
  wire v376bb88;
  wire v3740fe0;
  wire v373b11b;
  wire v374376b;
  wire v376beb4;
  wire v3a7165c;
  wire v3738e63;
  wire v37765a3;
  wire v3769ecf;
  wire v3741a71;
  wire v3a6ae14;
  wire v1e3751e;
  wire v375427c;
  wire v3a6a8b4;
  wire v373f6f7;
  wire v374a98e;
  wire v3a6ccfe;
  wire v3a6d665;
  wire v377a6e2;
  wire v3a5e881;
  wire v3765e79;
  wire v3740232;
  wire v3a5f7d7;
  wire v3a61a71;
  wire v375ef49;
  wire v37346e8;
  wire v37356b4;
  wire v37461d9;
  wire v3774385;
  wire v37729e0;
  wire v3a70582;
  wire v3777888;
  wire v3a6279c;
  wire v3a70454;
  wire v374d617;
  wire v3743cf5;
  wire v372a288;
  wire v3a574d7;
  wire v373413c;
  wire v37701cf;
  wire v3a70180;
  wire v3a5f38a;
  wire v37556ec;
  wire v377414c;
  wire v374d80f;
  wire v3749ec0;
  wire v376489b;
  wire v39e9c98;
  wire v3a62819;
  wire v3a61302;
  wire v3728d57;
  wire v3a63688;
  wire v373dd40;
  wire v3a6f9b4;
  wire v3734db5;
  wire v373601e;
  wire v375e12d;
  wire a53cf9;
  wire v3a715a9;
  wire v37629bf;
  wire v376aa76;
  wire v3a70e7d;
  wire v3a62250;
  wire v3a6913c;
  wire v3a5f0a5;
  wire v372f56c;
  wire v37494a7;
  wire v3741572;
  wire v373db82;
  wire v3a7125d;
  wire v37548e7;
  wire v3a70013;
  wire v37645a8;
  wire v3a70b92;
  wire v3806a6f;
  wire v3a70a50;
  wire v376f584;
  wire v3747e8e;
  wire v3a700b0;
  wire v3a65827;
  wire v3a70905;
  wire v3a712ac;
  wire v37283bb;
  wire v3a540a4;
  wire v3756430;
  wire v3a6fbd7;
  wire v3a6f65c;
  wire v373bd77;
  wire v3a6f49e;
  wire v373b687;
  wire v37501ad;
  wire v3730bf9;
  wire v3775144;
  wire v3775831;
  wire v3a70417;
  wire v3a71025;
  wire v3764a7d;
  wire v372b50b;
  wire v3a6adff;
  wire v372a0e3;
  wire v3a6ef17;
  wire v3763571;
  wire v372ca44;
  wire v3779cf9;
  wire v374809d;
  wire v3809788;
  wire v37366fc;
  wire v3a70e75;
  wire v373cdca;
  wire v373059e;
  wire v377e11d;
  wire v3771d4f;
  wire v3a60a6e;
  wire v3a6f3da;
  wire v3738679;
  wire v3a6b393;
  wire v3a6dfc9;
  wire v2aca778;
  wire v375c944;
  wire v3a538bd;
  wire v377bf77;
  wire v373c01b;
  wire v3a5b6de;
  wire v3751c4b;
  wire v3806c41;
  wire v3a58cf7;
  wire v39eb4cb;
  wire v376c80f;
  wire v3754682;
  wire v3735809;
  wire v376e833;
  wire v37639c6;
  wire v376f47f;
  wire v3763fb5;
  wire v3a71054;
  wire v3735051;
  wire v377a50f;
  wire v372b1e3;
  wire v3a7129f;
  wire v37614c1;
  wire v3759263;
  wire v3a7052e;
  wire v3a5b1ea;
  wire v376ff64;
  wire v3a6ff33;
  wire v3758c3d;
  wire v373afe9;
  wire v375491e;
  wire v372e3f5;
  wire v3a7024f;
  wire v37486de;
  wire v375029a;
  wire v38068c8;
  wire v372620f;
  wire v3a57508;
  wire v374217a;
  wire v37438ab;
  wire v3757921;
  wire v3a567ec;
  wire v376fa3e;
  wire v375cf04;
  wire v375aba9;
  wire v3747271;
  wire v374a0ab;
  wire v372c23b;
  wire v3779f1e;
  wire v376f536;
  wire v380909f;
  wire v373c617;
  wire v373a373;
  wire v3a617a6;
  wire v3728493;
  wire v3738c5f;
  wire v374a36b;
  wire v3377aee;
  wire v376d1dd;
  wire v3a713ea;
  wire v3771933;
  wire v37431ce;
  wire v37464e4;
  wire v3a5ebbf;
  wire v37337e7;
  wire v3724bf3;
  wire v375df28;
  wire v3a6022f;
  wire v376366a;
  wire v376d972;
  wire v37795a3;
  wire v3a5bca4;
  wire v3745f9b;
  wire v3a6b90f;
  wire v3809e93;
  wire v373e450;
  wire v37522ff;
  wire v376663a;
  wire v373ae83;
  wire v3a633b9;
  wire v37745b8;
  wire v377bfc0;
  wire v3a5ef6e;
  wire v372fd12;
  wire v3a6ff18;
  wire v373de13;
  wire v3a71267;
  wire v374e436;
  wire v3a70765;
  wire v3770f54;
  wire v37796ce;
  wire v23fe28c;
  wire v3a2a0f4;
  wire v3773666;
  wire v3a6f3cd;
  wire v3a70484;
  wire v3a5b52c;
  wire v3a587be;
  wire v3a710e4;
  wire v3a6f71a;
  wire v3a62fa7;
  wire v3762385;
  wire v37411bc;
  wire v3729fa0;
  wire v3a71166;
  wire v376d1bb;
  wire v374faf5;
  wire v372879a;
  wire v3a701c3;
  wire v374d9b3;
  wire v3a6fe44;
  wire v3734e69;
  wire v377a6dc;
  wire v3a7063e;
  wire v375b42e;
  wire v3a69544;
  wire v1e378b4;
  wire v3a70df4;
  wire v3772404;
  wire v3a6bbf0;
  wire v373bde3;
  wire v376e04c;
  wire v3a70bf1;
  wire v3a6fd6a;
  wire v3769e4c;
  wire v38078e5;
  wire v3a5ffac;
  wire v380946b;
  wire v3759b71;
  wire v3a7026a;
  wire v3a705d1;
  wire v37302c7;
  wire v3a5ff46;
  wire v3a71498;
  wire v3764e69;
  wire v377142b;
  wire v372c0fd;
  wire v3a5aaee;
  wire v37298f1;
  wire v3754df4;
  wire v3771d75;
  wire v3a5be41;
  wire v2093018;
  wire v3a2976c;
  wire v3a6c1f1;
  wire v3a70fc9;
  wire v375370a;
  wire v3a5e909;
  wire v3727943;
  wire v37685c3;
  wire v3756fbd;
  wire v3a6fac1;
  wire v376314e;
  wire v2092ee9;
  wire v8f1dd1;
  wire v3a58723;
  wire v3a6b57d;
  wire v3a5de59;
  wire v375d8f8;
  wire v3748a5d;
  wire v372cd04;
  wire v3727981;
  wire v372984e;
  wire v3a6542a;
  wire v3766b5a;
  wire v8cd321;
  wire v376543b;
  wire v3a5f218;
  wire v3a70bc4;
  wire v372567a;
  wire v373666f;
  wire v37287d2;
  wire v3a640e3;
  wire v37735ba;
  wire v3a5d99f;
  wire v3a702e0;
  wire v3a5df82;
  wire v375ae8d;
  wire v377c47c;
  wire v3a7061f;
  wire a4e409;
  wire v3a57f6c;
  wire v373a09f;
  wire v3a70578;
  wire v374d2d5;
  wire v374d255;
  wire v374b080;
  wire v3a6eaf8;
  wire v372354b;
  wire v372d4eb;
  wire v376a3c2;
  wire v3a5f4c6;
  wire v3746473;
  wire v3a6ff0e;
  wire v37710a4;
  wire v3a6f1d8;
  wire v376e68d;
  wire v39ebaee;
  wire v375e093;
  wire v3741f67;
  wire v3a65e55;
  wire v37261ad;
  wire v3a5f6da;
  wire v372e571;
  wire v375e9ca;
  wire v3755ae2;
  wire v3a70a16;
  wire v37274e6;
  wire v376bf8a;
  wire v37701af;
  wire v3a7022f;
  wire v375c19b;
  wire v3a6d6fb;
  wire v3a6b1bf;
  wire v3772f74;
  wire v3756d6e;
  wire v3a6f6e0;
  wire v3a70b52;
  wire v374efad;
  wire v3756595;
  wire v3769e50;
  wire v3a70a75;
  wire v3a70af0;
  wire v3758b8b;
  wire v3727a6d;
  wire v374bdac;
  wire v376a946;
  wire v3a71032;
  wire v3757a61;
  wire v376f641;
  wire v372ab19;
  wire v373e219;
  wire v373fd94;
  wire v374c6b8;
  wire v3a713d5;
  wire v3a5df66;
  wire v3a6e4ec;
  wire v375ede6;
  wire v3a5cdef;
  wire v37690e7;
  wire v372317f;
  wire v3a70242;
  wire v3772e44;
  wire v3758892;
  wire v3a6a76d;
  wire v3771622;
  wire v3763f20;
  wire v375aff6;
  wire v3759786;
  wire v373ea09;
  wire v37409f6;
  wire v373e873;
  wire v3a6ba08;
  wire v3a70fca;
  wire v3a5ebc2;
  wire v375af91;
  wire v373b2da;
  wire v3758672;
  wire v374f077;
  wire v3734c47;
  wire v3a6f550;
  wire v37583f0;
  wire v3a6f758;
  wire v3771cf7;
  wire v37597f4;
  wire v375372b;
  wire v3a7166f;
  wire v38094b8;
  wire v3a6f8d9;
  wire v3772cab;
  wire v3a58a3b;
  wire v37517f7;
  wire ac4b49;
  wire v3a6dbbf;
  wire v3775ec8;
  wire v37495ed;
  wire v3a69539;
  wire v375049a;
  wire v376bc32;
  wire v3a6a4b9;
  wire v376ae7f;
  wire v377bf7b;
  wire v373c52e;
  wire v3737a8b;
  wire v3a5faf0;
  wire v3a6fa20;
  wire v377113b;
  wire v37345aa;
  wire v3a6f610;
  wire v374d43f;
  wire v374e4fa;
  wire v3a66c12;
  wire v3760276;
  wire v3730252;
  wire v376fdd4;
  wire v3a70676;
  wire v377b058;
  wire v3a7107e;
  wire v3777bcf;
  wire v3a57b57;
  wire v3746746;
  wire v3750f4c;
  wire v37373bb;
  wire v373a4cd;
  wire v9243ac;
  wire v3a6639e;
  wire v3a70c06;
  wire v375f28d;
  wire bd1306;
  wire v37263d2;
  wire v3a6df51;
  wire v3726bb7;
  wire v3a70eee;
  wire v3751a97;
  wire v3a6a6e1;
  wire v3764bf2;
  wire v3a7129c;
  wire v3730fbd;
  wire v3748e0c;
  wire v3763b4d;
  wire v3723d79;
  wire v376769e;
  wire v39eaae9;
  wire v3748059;
  wire v372a683;
  wire v37690da;
  wire v372d773;
  wire v3a5d21b;
  wire v3765203;
  wire v3a6e231;
  wire v3a6f09d;
  wire v377d4dd;
  wire v3a68757;
  wire v3762d09;
  wire v377b0d8;
  wire v3769696;
  wire v3a5584b;
  wire v3a626fe;
  wire v3a61c80;
  wire v373e07e;
  wire v3746f9d;
  wire v377b205;
  wire v3a64f96;
  wire v3726072;
  wire v3745bdc;
  wire v3a5ed86;
  wire v3730722;
  wire v3a68315;
  wire v377cb3d;
  wire v3806465;
  wire v37402a4;
  wire v3a5d62d;
  wire v3a592bb;
  wire v2acb5bc;
  wire v376f51c;
  wire v3a706c9;
  wire v3a6f81c;
  wire v372685c;
  wire v3a710ea;
  wire v3a69b91;
  wire v374a189;
  wire v373f6e7;
  wire v3a6ae19;
  wire v3a715d0;
  wire v377b2e1;
  wire v3a6826a;
  wire v37722a0;
  wire v3a6edb5;
  wire v3763d53;
  wire v3749469;
  wire v9d70f0;
  wire v3734d20;
  wire v376daa7;
  wire v3725673;
  wire v377fc45;
  wire v3751eb6;
  wire v374c522;
  wire v3755bb4;
  wire v372ff54;
  wire v3a70dd3;
  wire v3779a80;
  wire v3a5878e;
  wire v376002d;
  wire v374f272;
  wire v3749fc1;
  wire v374ebbf;
  wire v375d2ff;
  wire v372bce5;
  wire v3740893;
  wire v377b6de;
  wire v2acafac;
  wire v3760a0b;
  wire v3a5b181;
  wire v3a69b19;
  wire v376a06c;
  wire v373168f;
  wire v3a66ea0;
  wire v372c1bb;
  wire v37509c4;
  wire v3751406;
  wire v37392ae;
  wire v3738f30;
  wire v373b4e3;
  wire v3a700af;
  wire v3725c6c;
  wire v375d364;
  wire v375f2e8;
  wire v3a6f1c8;
  wire v3731517;
  wire v372b20b;
  wire v373c8ba;
  wire v377d2bb;
  wire v376e795;
  wire v377b94e;
  wire v3a6f7e9;
  wire v1e377f7;
  wire v3a6b643;
  wire v377caa8;
  wire v3751012;
  wire v373aa47;
  wire v373643b;
  wire v377b7d0;
  wire v3a6f843;
  wire v3773ad7;
  wire v372e83a;
  wire v3a5ac5c;
  wire v3a5905e;
  wire v37386a9;
  wire v3750fc8;
  wire v3a69de7;
  wire v3a64421;
  wire v374a9d0;
  wire v372e8ed;
  wire v3a6fae5;
  wire v372dadb;
  wire v2092ffc;
  wire v37765e1;
  wire v374faa9;
  wire v3726d1f;
  wire v3a70374;
  wire v3a70f66;
  wire v377e328;
  wire v374b285;
  wire v373f6cf;
  wire v3731088;
  wire v3a71055;
  wire v3a6f123;
  wire v37785f8;
  wire v37681a3;
  wire v37497d6;
  wire v372a421;
  wire v376dc21;
  wire v3774fa8;
  wire v3775bf6;
  wire d435c2;
  wire v372dec8;
  wire v3a71345;
  wire v375fbd7;
  wire v372842d;
  wire v3731afc;
  wire v3a6eb0b;
  wire v377c929;
  wire v3a6fefa;
  wire v373a802;
  wire v3764994;
  wire v37650bd;
  wire v3377b1b;
  wire v373af5d;
  wire v37404da;
  wire v2925d19;
  wire v3749bf0;
  wire v373471f;
  wire v37544cb;
  wire v3732086;
  wire v3a5c65e;
  wire v3a6fc7f;
  wire v374581a;
  wire v3755e61;
  wire v3740d3b;
  wire v37297ce;
  wire v37493b4;
  wire v3751383;
  wire v37403b1;
  wire v3a7148d;
  wire v3732b98;
  wire v3a706c7;
  wire v37366d2;
  wire v374b4a4;
  wire v3727db9;
  wire v3a6bb84;
  wire v3a706fe;
  wire v3763da5;
  wire v37512c1;
  wire v38067b3;
  wire v3730038;
  wire v377b4b0;
  wire v3a6f449;
  wire v3727a04;
  wire v3774452;
  wire v3a5b448;
  wire v3a708a6;
  wire v3753278;
  wire v375a842;
  wire v375ac6a;
  wire v3a5a585;
  wire v3a6fbfc;
  wire v3724e67;
  wire v3733ba1;
  wire v3a6440f;
  wire v37524a6;
  wire v3766a98;
  wire v39a5293;
  wire v376999e;
  wire v376572c;
  wire v377d10c;
  wire v3a700e5;
  wire v3a6cc67;
  wire v3a6fd89;
  wire v373506a;
  wire v373d9e0;
  wire v3a6c6ce;
  wire v376e1fd;
  wire v3a62e92;
  wire v3750fee;
  wire v3a707b9;
  wire v3a6f080;
  wire v3a5d25d;
  wire v94335e;
  wire v3a61c73;
  wire v3a712b7;
  wire v37674fb;
  wire b08e51;
  wire aac430;
  wire v375d149;
  wire v23fe0c2;
  wire v3736d47;
  wire v3a6f6a9;
  wire v374de43;
  wire v372c016;
  wire v374f838;
  wire v3a6774e;
  wire v377910a;
  wire v3a572e9;
  wire v376085a;
  wire v37784ad;
  wire v3a70183;
  wire v372af77;
  wire v3747edc;
  wire v9204d4;
  wire v3a58200;
  wire v377ba59;
  wire v3754caa;
  wire v3a5aad8;
  wire v3778c7f;
  wire v374d86e;
  wire v372a704;
  wire v377981a;
  wire v3806ed4;
  wire v375bfc4;
  wire v377c965;
  wire v372a298;
  wire v3727a12;
  wire v3728625;
  wire v37297cb;
  wire v3a6817f;
  wire v3806575;
  wire v375eaea;
  wire v375f0c9;
  wire v3a656c7;
  wire v3779b5b;
  wire v372c00a;
  wire v375c10c;
  wire v3735113;
  wire v3774b58;
  wire v375a455;
  wire v3a603bb;
  wire v3752fb7;
  wire v3a582d6;
  wire v373f953;
  wire v3771ab9;
  wire v374c61d;
  wire v3a71425;
  wire v374faa2;
  wire v3a687a7;
  wire v3725710;
  wire v3768349;
  wire v3a70525;
  wire v3a63331;
  wire v3741bb2;
  wire v37690f3;
  wire v372e9f3;
  wire v375b980;
  wire v3754b2c;
  wire v3a6e793;
  wire v3a6f4af;
  wire v372e873;
  wire v374243d;
  wire v373c3a0;
  wire v3a5e496;
  wire v3747ea2;
  wire v373d955;
  wire v3749e8a;
  wire v377fbd5;
  wire a9f66a;
  wire v3a70dd0;
  wire v37251b9;
  wire v376195f;
  wire v3738d0b;
  wire v3774aa2;
  wire v377e29a;
  wire v373d0d1;
  wire v375c0c4;
  wire v3760b79;
  wire v3759f09;
  wire v3a6f025;
  wire v373b0d2;
  wire v372b8fd;
  wire v8d4314;
  wire v3738e3c;
  wire v377ce3f;
  wire v3a6fa7c;
  wire v377bb38;
  wire v375e1b0;
  wire v3a6eece;
  wire v37397ba;
  wire v377e9b0;
  wire v373308b;
  wire v3a66856;
  wire v377f264;
  wire v372450e;
  wire v3742b31;
  wire v3a7106f;
  wire v3765ce2;
  wire v372b9c6;
  wire v3a64703;
  wire v3a57b0d;
  wire v3a5ab6e;
  wire v3a6c8dc;
  wire v3a54d84;
  wire v39eb3bd;
  wire v3731004;
  wire v373e789;
  wire v3a7103d;
  wire v3747bea;
  wire v3a5e2e1;
  wire v3a57658;
  wire v37346dc;
  wire v3752556;
  wire v372efb4;
  wire v374b526;
  wire v3a69676;
  wire v3a6f914;
  wire v3770bf5;
  wire v3a5a591;
  wire v37789da;
  wire v3a6837d;
  wire v3753d51;
  wire v37406ca;
  wire v374165f;
  wire v3757091;
  wire v3a571fd;
  wire v3a70876;
  wire v3a5ab33;
  wire v3776323;
  wire v375408a;
  wire v37682c0;
  wire v3a62e1e;
  wire v3739f22;
  wire v3a69488;
  wire v372d741;
  wire v23fd967;
  wire v3a67b86;
  wire v37792cf;
  wire v373c7a5;
  wire v3775999;
  wire b04260;
  wire v3751db5;
  wire v3a70b00;
  wire v375e647;
  wire v374b0cb;
  wire v3a6d897;
  wire v375129f;
  wire v375c903;
  wire v3a7160d;
  wire v3a66534;
  wire v3757956;
  wire v3a5992f;
  wire v37577cd;
  wire v3754ba1;
  wire v3734fa9;
  wire v375b3af;
  wire v37275ef;
  wire v3727ffa;
  wire baf7ba;
  wire v3738df9;
  wire v375c439;
  wire v3a70fd1;
  wire v3a67691;
  wire v377af10;
  wire v37652f1;
  wire v3775725;
  wire v3732bd2;
  wire v375f9e9;
  wire v3a614a1;
  wire v3762281;
  wire v372f87b;
  wire v3a70bb7;
  wire v374145b;
  wire v372a13a;
  wire v3741f08;
  wire v376a9ee;
  wire v3749356;
  wire v3a704d0;
  wire v3743425;
  wire v37554c0;
  wire v3a70b76;
  wire v3a70f8d;
  wire v374829e;
  wire v3a6f7ed;
  wire v3730c0a;
  wire v3762e66;
  wire v3a5d08e;
  wire v3a712bf;
  wire v376cd84;
  wire v3a65ce7;
  wire v3a6f4a3;
  wire v37306c6;
  wire v37756ac;
  wire v377002f;
  wire v3a6ed79;
  wire cecaa5;
  wire v3730986;
  wire v373cd03;
  wire v3a60a68;
  wire a72315;
  wire v3a6ef22;
  wire v375166c;
  wire v3a5e6f6;
  wire v3a629a6;
  wire v3a69c57;
  wire v372a85f;
  wire v375bdcc;
  wire v3773eeb;
  wire v375f2a3;
  wire v372ab85;
  wire v3a6f333;
  wire b6b4ea;
  wire v3a709a0;
  wire v3a573e3;
  wire v37407b3;
  wire v3733c39;
  wire v3809b44;
  wire v3a67698;
  wire v3a67603;
  wire v3a6f949;
  wire v3752400;
  wire v372afd2;
  wire v3a703d0;
  wire v3a6f61f;
  wire v3a7118a;
  wire v3a6ffff;
  wire v3762312;
  wire v3a5aacb;
  wire v3a6f0a5;
  wire v3739e7a;
  wire v1e37558;
  wire v373b0d0;
  wire v3764a2d;
  wire v3763b5d;
  wire v3725671;
  wire v375a3a8;
  wire v374523b;
  wire v3a5b1ec;
  wire v3727c62;
  wire v374d33d;
  wire v3a64aa0;
  wire v3778a8b;
  wire v374b3f8;
  wire v373339c;
  wire v3a69b5f;
  wire v3a6ec06;
  wire v3a6f169;
  wire v3760e47;
  wire v3a70bb3;
  wire a22759;
  wire v37427d3;
  wire v3a70ea0;
  wire v3732b81;
  wire v376a34d;
  wire v3a5b2fd;
  wire v3a618b3;
  wire v37398eb;
  wire v376b7db;
  wire v375b2fe;
  wire v3a654af;
  wire v3742b24;
  wire v37266cb;
  wire v3725799;
  wire v37664e7;
  wire v3a67f97;
  wire v376c777;
  wire v3a7081c;
  wire v3a6fe5b;
  wire v374794f;
  wire v3a6abaa;
  wire v377cc23;
  wire v3756398;
  wire v374fd4a;
  wire v3806ff0;
  wire v375abcd;
  wire v3723495;
  wire v3a714d2;
  wire v3a6a051;
  wire v377d9bb;
  wire v377870b;
  wire v3a704e7;
  wire v3a6f326;
  wire v3779264;
  wire d3b3b2;
  wire v3763d3a;
  wire v3751831;
  wire v3749e48;
  wire v3a6e3bb;
  wire v3765c85;
  wire v3760343;
  wire v372dd89;
  wire v374668c;
  wire v3a6fc6a;
  wire v37434ce;
  wire v3732187;
  wire v373f124;
  wire v3a67e53;
  wire v3733ae1;
  wire v3722c80;
  wire v372f59c;
  wire v376e74b;
  wire v3725827;
  wire v2ff8e5c;
  wire v3a63c15;
  wire v3a70c19;
  wire v3758ab0;
  wire v3a6f90c;
  wire v377ee7c;
  wire v3736fb4;
  wire v3766ef9;
  wire v375be5b;
  wire v3728b9d;
  wire v37769ee;
  wire v3a559f0;
  wire v3769605;
  wire ca602f;
  wire v3a6741a;
  wire v3722e4c;
  wire v37259bc;
  wire v3744f0d;
  wire v2093234;
  wire v3a706ed;
  wire v3a5cd72;
  wire v376d29a;
  wire v3a6f08a;
  wire v3a712d1;
  wire v3a5e244;
  wire v3727472;
  wire v3a7026c;
  wire v3767f06;
  wire v377205d;
  wire v372e8d8;
  wire v375624b;
  wire v372bbd2;
  wire v3727d00;
  wire v3777d39;
  wire v3a6f329;
  wire v37584e6;
  wire v3762a76;
  wire v3a7114a;
  wire v375e30b;
  wire v3774d04;
  wire v377ed71;
  wire v372998c;
  wire v3754e7b;
  wire v374abc9;
  wire v377b860;
  wire v3735c9d;
  wire v3722bca;
  wire v3a53a2d;
  wire v3751a9f;
  wire v3a62bae;
  wire v373ead8;
  wire v3a6fdef;
  wire cf4a8f;
  wire v3748cbd;
  wire v3759947;
  wire v3724f7b;
  wire v376dab5;
  wire v372a116;
  wire v3758df6;
  wire v3a700db;
  wire v3a66e6f;
  wire v376d215;
  wire v376e2a4;
  wire v39ea259;
  wire v3723e23;
  wire v3a64b55;
  wire v9c1340;
  wire v3757272;
  wire v3733b02;
  wire v376775d;
  wire v3772a27;
  wire v3377adc;
  wire v373bd70;
  wire v3a5b4d6;
  wire v376ddb6;
  wire v3a7017d;
  wire v3769cc4;
  wire v3809dfb;
  wire v373d943;
  wire v37237f1;
  wire v3a53d04;
  wire v37571c8;
  wire v377aed1;
  wire v373a9fb;
  wire v375e512;
  wire v3731b28;
  wire v3a58f56;
  wire v3a5ef9d;
  wire v373d5b7;
  wire d24921;
  wire v3768fb7;
  wire v3a713ad;
  wire v3a69913;
  wire v376b220;
  wire b0015f;
  wire v3a57037;
  wire v37667f8;
  wire v376cddf;
  wire v377e30e;
  wire v3a6c4bb;
  wire v3a5b89a;
  wire v374b912;
  wire v3a71343;
  wire v3736ae6;
  wire v375c4cb;
  wire v3a642c5;
  wire v3a6d792;
  wire v3739082;
  wire v376256c;
  wire v3a70c33;
  wire v3a6ffc1;
  wire v375c381;
  wire v3726d4a;
  wire v375973d;
  wire v3a63b26;
  wire v3a70f61;
  wire v374d258;
  wire v3740d9e;
  wire v3742725;
  wire v372ab6c;
  wire v3727e69;
  wire v3730370;
  wire v37634d0;
  wire v377ef71;
  wire v373c076;
  wire v3a71427;
  wire v375a28e;
  wire v3742950;
  wire v376a47e;
  wire v3a6fab8;
  wire v3769d4c;
  wire v3a6c922;
  wire v39a4e1f;
  wire v3a70d21;
  wire v3a70f27;
  wire v3778c14;
  wire v3a6c3ac;
  wire v375d1ae;
  wire v3a70a03;
  wire v3a709ec;
  wire v374853c;
  wire v372b8eb;
  wire v373303f;
  wire v3748f03;
  wire v2aca783;
  wire v3739f0e;
  wire v373690a;
  wire v377e889;
  wire v377429c;
  wire v373b50e;
  wire v373a90e;
  wire v3a709d2;
  wire v3a6ff82;
  wire v3a632aa;
  wire v372b906;
  wire v377150c;
  wire v3a6ff10;
  wire v372e790;
  wire v3a6fe33;
  wire v3a6bf22;
  wire v373e154;
  wire v376af98;
  wire v3770f55;
  wire v372febd;
  wire v374db21;
  wire v3a70514;
  wire v3737220;
  wire v3a6f5e1;
  wire v376574a;
  wire v3758e1c;
  wire v3a6efeb;
  wire v3a6e872;
  wire v377653f;
  wire v3750d61;
  wire v3a70e28;
  wire v3748262;
  wire v375f88a;
  wire v3738061;
  wire v37756ab;
  wire v37787c1;
  wire v3a6e318;
  wire v37383da;
  wire v3a5d405;
  wire v3a6deea;
  wire v3768288;
  wire v3759f66;
  wire v3728213;
  wire v3a675f7;
  wire v376af6a;
  wire v3778dd7;
  wire v3746d4a;
  wire v3808fce;
  wire v3724731;
  wire v377d367;
  wire v3a5b7db;
  wire v37760f9;
  wire v3a5715d;
  wire v3808952;
  wire v37318e2;
  wire v357731b;
  wire v3766e55;
  wire v37611a9;
  wire v2ff8e9a;
  wire v3a59d65;
  wire v373a141;
  wire v372e25b;
  wire v3a701a2;
  wire v3a705e6;
  wire v3743f7a;
  wire v373dfb5;
  wire v3a63df4;
  wire v375c432;
  wire v3a6f1fb;
  wire v37449fc;
  wire v948ef2;
  wire v3a6f3f0;
  wire v3759c23;
  wire v3a6ffee;
  wire v3759a4a;
  wire v373ebcf;
  wire v376c89f;
  wire v37245a1;
  wire v3756ead;
  wire v3753298;
  wire v37606f4;
  wire v3a702f6;
  wire v373fb22;
  wire v2acae79;
  wire v3a6fd76;
  wire v3765dbe;
  wire v375c85c;
  wire v3724ced;
  wire v3754c99;
  wire v3736684;
  wire v3a6130e;
  wire v374c576;
  wire v374d31a;
  wire v373432d;
  wire v3a7093f;
  wire v3a62846;
  wire v3a6f59e;
  wire v37288bc;
  wire v376fbb5;
  wire v3a62753;
  wire v375df71;
  wire v372ddbc;
  wire v3737d23;
  wire v3809eb1;
  wire v3a6cf75;
  wire v3723e62;
  wire v3a6a208;
  wire v3728a53;
  wire v3a7076e;
  wire v3a70f62;
  wire v3a56789;
  wire v3778fb5;
  wire v3a5d185;
  wire v373ac84;
  wire v372809b;
  wire v376293b;
  wire v3759b93;
  wire v374f243;
  wire v373f5fc;
  wire v377dadb;
  wire v3a7031f;
  wire v3809a8b;
  wire v3775f4f;
  wire v37793e4;
  wire v3a705d5;
  wire v3748ba9;
  wire v3a6f70b;
  wire v376d542;
  wire v374d59a;
  wire v380704f;
  wire v3a7029b;
  wire v3a5c366;
  wire v3a712b6;
  wire v3724f24;
  wire v37730bf;
  wire v3742cfe;
  wire v3771e8d;
  wire v3754b61;
  wire v372c500;
  wire v372495f;
  wire dc6ded;
  wire v374ad67;
  wire v376c76d;
  wire v3a6fd4b;
  wire v3a66c6c;
  wire v3766d5a;
  wire v3a6b51f;
  wire v374aec2;
  wire v37293e0;
  wire v3a63ece;
  wire v3763a86;
  wire v3774deb;
  wire v3763db6;
  wire v372a1d4;
  wire v3a70d7b;
  wire v3735abc;
  wire v3a6f5aa;
  wire v209306f;
  wire v3733b90;
  wire v3a71512;
  wire v376d36a;
  wire v372c345;
  wire v37251f6;
  wire v23fdf85;
  wire v374d40b;
  wire v3754f5d;
  wire v376d081;
  wire v373fe7b;
  wire v8f559e;
  wire v37659e2;
  wire v3a6b70e;
  wire v3a70336;
  wire v3a70d44;
  wire v3a61a76;
  wire v3a6f998;
  wire v3a70890;
  wire v373f07d;
  wire v3a5aefc;
  wire v37717ee;
  wire v376ecae;
  wire v374ecf9;
  wire v37626b9;
  wire v3a70f35;
  wire v3a647e7;
  wire v3731211;
  wire v373a8d6;
  wire v377538f;
  wire v3772c19;
  wire v337830d;
  wire v3a713be;
  wire v3a5a29e;
  wire v3750f72;
  wire v377704c;
  wire v372673d;
  wire v373a16b;
  wire v37691d1;
  wire v373706e;
  wire v3a5a323;
  wire v3a623dc;
  wire v3a6bab2;
  wire v377cd0d;
  wire v3a658b0;
  wire v373b759;
  wire v3a53bb3;
  wire v3767266;
  wire v3a6767d;
  wire v3777cb9;
  wire v3a55838;
  wire v373f3b5;
  wire v3770fbc;
  wire v3767385;
  wire v37664a1;
  wire v3a296e8;
  wire v377d74c;
  wire v376739f;
  wire v37565a6;
  wire v3753d94;
  wire v376d2c6;
  wire v375ee2e;
  wire v3779a9c;
  wire v38076bb;
  wire v3a5f05e;
  wire v377b8f9;
  wire v3a647e0;
  wire v374a4cc;
  wire v3a60443;
  wire v3a68c27;
  wire v3729a07;
  wire v37406a7;
  wire v376c351;
  wire v3a70125;
  wire v3741dac;
  wire v3a703bb;
  wire v376c30a;
  wire v372cfd5;
  wire v3729b9f;
  wire v3774b98;
  wire v3a6f442;
  wire v3756109;
  wire v377f26e;
  wire v37602e0;
  wire v375e9a9;
  wire v3750087;
  wire v3a70d36;
  wire v3742a8e;
  wire v375f2c7;
  wire v3748494;
  wire v3a61ceb;
  wire v37360c1;
  wire ab0224;
  wire v3a70fc4;
  wire v377b66a;
  wire v3766cfb;
  wire v3a705ae;
  wire v3a614a0;
  wire v3748acd;
  wire a14297;
  wire v3a6c628;
  wire v3a7005b;
  wire v3a6799d;
  wire v3a7128b;
  wire v3808dd0;
  wire v3a62c11;
  wire v372b27e;
  wire v3761d9f;
  wire v373af26;
  wire v3a298b6;
  wire v3a642ab;
  wire v3a6199d;
  wire ac9d0d;
  wire v377f397;
  wire v37621ff;
  wire v372bfbb;
  wire v376b1be;
  wire v376ea51;
  wire v377bf2d;
  wire v3778f6c;
  wire v373d753;
  wire v374cd7e;
  wire v3740de5;
  wire v3a65856;
  wire v372f95b;
  wire v374b310;
  wire v3739e39;
  wire v374e6a5;
  wire v3a6edb9;
  wire v372731e;
  wire v377bb66;
  wire v3a55b61;
  wire v3a65d4e;
  wire v3a6d0a1;
  wire v375a80c;
  wire v3a707a0;
  wire v372d95c;
  wire v3753dd4;
  wire v375cc06;
  wire v3a63884;
  wire v376d86d;
  wire v3746202;
  wire v375f823;
  wire v3733d02;
  wire v375a6be;
  wire v38073be;
  wire v374686d;
  wire v3a5ac38;
  wire v3a6811a;
  wire v3a70933;
  wire v37753dc;
  wire v3762d80;
  wire v3739d22;
  wire v3733dd4;
  wire v3a6c672;
  wire v3745f4a;
  wire v3a6fedb;
  wire v3761909;
  wire v3a5a09c;
  wire v3a6fee9;
  wire v37791a7;
  wire v37425a7;
  wire v3a6bf60;
  wire v3729561;
  wire v375068a;
  wire v376804b;
  wire v3728ea7;
  wire v3759361;
  wire v372c1b0;
  wire v373ace1;
  wire v375e356;
  wire v3768e7e;
  wire v37431ec;
  wire v374184c;
  wire v3a6f751;
  wire v3757695;
  wire v3768304;
  wire v3753b6a;
  wire v372a71e;
  wire v3765021;
  wire v3a6f78a;
  wire v3a6f4ed;
  wire v3a6d09c;
  wire v374dc13;
  wire v375be64;
  wire v373c064;
  wire v360d0db;
  wire v3729115;
  wire v377a43e;
  wire v3749629;
  wire v37366b5;
  wire b516f2;
  wire v3737209;
  wire v376f501;
  wire v372462b;
  wire v3751e5e;
  wire v3a6afe8;
  wire v377d6ba;
  wire v38078ed;
  wire v375431d;
  wire v3a612a4;
  wire v3732715;
  wire v3a6ff3c;
  wire v37389db;
  wire v376e316;
  wire v376b018;
  wire v3a709cf;
  wire v377b4b9;
  wire v3a711fa;
  wire v3a68255;
  wire v380879c;
  wire v3730a93;
  wire v3723d4b;
  wire v3a6b92c;
  wire v3a70b3a;
  wire v37383f6;
  wire v375021b;
  wire v374cb05;
  wire v3a6f30f;
  wire v376f9b5;
  wire v374ed99;
  wire v3a6eddd;
  wire v3729ae9;
  wire v3735c5a;
  wire v377763c;
  wire v376c26e;
  wire v3733440;
  wire v3a669e9;
  wire v3770366;
  wire v377bbd9;
  wire v377e27e;
  wire v3a6ef0e;
  wire v3577421;
  wire v3a6f07d;
  wire v3a70a51;
  wire v375f2f2;
  wire v373c1ff;
  wire v1e379cc;
  wire v375b01e;
  wire v3758ce2;
  wire v376b38c;
  wire v3a5a039;
  wire v375517b;
  wire v3736b4a;
  wire v3a7115e;
  wire v372ebd5;
  wire v3a6f894;
  wire v374bac7;
  wire v3746825;
  wire v3a64e75;
  wire v377e915;
  wire v3a64c14;
  wire a52d64;
  wire v3761847;
  wire v376195b;
  wire v3a54222;
  wire v373f3e4;
  wire v3257687;
  wire v375ae3d;
  wire v377807f;
  wire v376b65a;
  wire v37318e3;
  wire v37287e1;
  wire v377e018;
  wire v37548a5;
  wire v3a6fcdc;
  wire v3a58d5f;
  wire v3a6eb97;
  wire v3a70de3;
  wire v375a33d;
  wire v3776859;
  wire v3740c73;
  wire v88b8eb;
  wire v3766d29;
  wire v373b380;
  wire v3a554f0;
  wire v3a56c60;
  wire v3a6f72f;
  wire v3770e77;
  wire v3749544;
  wire v3746312;
  wire v3a6e33a;
  wire v376f39f;
  wire v3754ee0;
  wire v3a6f6ea;
  wire v3732bff;
  wire v372b5bc;
  wire v377d491;
  wire v3728b10;
  wire v3a6efc7;
  wire v3808e6b;
  wire v3764203;
  wire v3a6fe91;
  wire v375076a;
  wire v377b096;
  wire v3728eca;
  wire v3a6f9ed;
  wire v3a6f9ce;
  wire v3753a1d;
  wire v3745510;
  wire v3745b39;
  wire v3779a9a;
  wire v3769c81;
  wire v377f83c;
  wire v376df02;
  wire v375efc9;
  wire v37796f6;
  wire v3758d37;
  wire v3a55673;
  wire v3771d0f;
  wire v3577376;
  wire v3a680f4;
  wire v377da26;
  wire v376ba2e;
  wire v3770234;
  wire v372dec3;
  wire v3748d1f;
  wire v375d6e8;
  wire v374febd;
  wire v3a5b51a;
  wire v3a5f7b8;
  wire v373d91f;
  wire v377aeba;
  wire v373a333;
  wire v3a6fba1;
  wire v3742521;
  wire v37667b3;
  wire v373557c;
  wire v3a6dae5;
  wire v37512f3;
  wire v372ead6;
  wire v37512dc;
  wire v375dba4;
  wire v373facf;
  wire v39a4c67;
  wire v3a6ddea;
  wire v3a6efa1;
  wire v3a6f3e7;
  wire v3a70030;
  wire v3a71162;
  wire v372f260;
  wire v3a587d6;
  wire v3748972;
  wire v3766799;
  wire v3748755;
  wire v377cece;
  wire v3a6f718;
  wire v3725f9b;
  wire v3749a38;
  wire v3a5d48f;
  wire v3a6f2bf;
  wire v3a551e4;
  wire v3725564;
  wire v3a5de73;
  wire v3737628;
  wire v3725494;
  wire v37763c2;
  wire v374d965;
  wire v3a6f477;
  wire v3a714cc;
  wire v3728963;
  wire v3a55419;
  wire v375c0d6;
  wire v3774f4e;
  wire v3a6f17b;
  wire v37573a3;
  wire v1e37c0d;
  wire v3a70460;
  wire v3a714e1;
  wire v3a6cb4e;
  wire v374c8ec;
  wire v3a714ad;
  wire v3735fca;
  wire v3742f4c;
  wire v3734100;
  wire v3809ee9;
  wire v3a55b93;
  wire v37616e0;
  wire v376d7ee;
  wire v3a6ebcc;
  wire v375fbb7;
  wire v376646a;
  wire v3a627a7;
  wire v374d63f;
  wire v3735444;
  wire v377ae81;
  wire v375df25;
  wire v375e4a0;
  wire v37c00b6;
  wire v376b4a8;
  wire v376bb05;
  wire v3a62589;
  wire v3750ef8;
  wire v37535ae;
  wire v3770ab1;
  wire v3726cc1;
  wire v3a5574a;
  wire v3a709d0;
  wire v374d3b8;
  wire v3a60fd6;
  wire v3a5e10c;
  wire v37263b9;
  wire v3a6b46d;
  wire v3a5e5d0;
  wire v3758ea7;
  wire v375693b;
  wire v3a6fec4;
  wire v377efa7;
  wire v3a70384;
  wire v3731f9a;
  wire v3a70fe9;
  wire v3772310;
  wire v377746e;
  wire v376dc44;
  wire v373931a;
  wire v374f345;
  wire v3a60826;
  wire v3a7115c;
  wire v3756f77;
  wire v37631a9;
  wire v375fdc9;
  wire v373bac6;
  wire v3748966;
  wire v3a64a9a;
  wire v3743ec6;
  wire v3a70e16;
  wire v376a40c;
  wire v3a6eb53;
  wire v3741e9f;
  wire v9e6ddd;
  wire v3a67acf;
  wire v3769b3f;
  wire v37399f7;
  wire v377a89f;
  wire v3a607ba;
  wire v3724d8b;
  wire v377fb55;
  wire v3a6f3be;
  wire v3a6f396;
  wire v3733ba7;
  wire v33789ef;
  wire v3750b02;
  wire bb70de;
  wire v3741bd8;
  wire v376b743;
  wire v3a5bd9c;
  wire v376910a;
  wire v3757f6d;
  wire v3770bca;
  wire v3761351;
  wire v37325b9;
  wire v3a70955;
  wire v373bded;
  wire v3a700a3;
  wire v3a703cb;
  wire v376ec9b;
  wire v3736011;
  wire v3a70b20;
  wire v3a5b960;
  wire v3a5c040;
  wire v3757311;
  wire v3776ff3;
  wire v3751c65;
  wire v3a5eecb;
  wire v3729385;
  wire v3750553;
  wire v3759203;
  wire v3724f05;
  wire v3a6ec29;
  wire v3a6ccc4;
  wire v3a5ad26;
  wire v3a66aa6;
  wire v3763e30;
  wire v374f0ac;
  wire v3734534;
  wire v3a71332;
  wire v374093f;
  wire v3a5b514;
  wire v3724811;
  wire v372f4fe;
  wire v3a7055c;
  wire v37399d4;
  wire v3a713da;
  wire v3a5666f;
  wire v37332eb;
  wire b44720;
  wire v3a70662;
  wire v3a5d2f9;
  wire v377ed18;
  wire v375803d;
  wire v3a5d548;
  wire v373dac4;
  wire v37724fc;
  wire v374e7fa;
  wire v3a6f697;
  wire v37692e3;
  wire v374148a;
  wire v3743f2c;
  wire v377e67a;
  wire v372d1ae;
  wire v376e20f;
  wire v3a60859;
  wire v373b1bb;
  wire v3a70819;
  wire dbf06b;
  wire v3a6fc94;
  wire v3a6ffe2;
  wire v3768c76;
  wire v373bfdd;
  wire v3a5be3f;
  wire v372a4ae;
  wire v3a7104f;
  wire v3806ff5;
  wire v3772f32;
  wire v3a683c6;
  wire d320a7;
  wire v374ca2e;
  wire v3a711c3;
  wire v3726b63;
  wire v37624a9;
  wire v3a66bfa;
  wire v3a2a106;
  wire v372bebe;
  wire v3a6a1d9;
  wire v375e349;
  wire v3a70d7e;
  wire v37242fa;
  wire v375b56c;
  wire v3a5b925;
  wire v37401bb;
  wire v3777c9b;
  wire v3a704ff;
  wire v3748d6c;
  wire v377118b;
  wire v3749f9d;
  wire v375fe15;
  wire v3a6f20f;
  wire v3a6a346;
  wire v3a6f908;
  wire v3752131;
  wire v373b166;
  wire v37650b8;
  wire v376430d;
  wire v3a5e62b;
  wire v375d9df;
  wire v372a39a;
  wire v372f4e6;
  wire v3771633;
  wire v372863f;
  wire v3748d3c;
  wire v3755f23;
  wire v3a706c3;
  wire v3a63eff;
  wire v376ebbf;
  wire v376ee80;
  wire v3735e89;
  wire v37787da;
  wire v37267d6;
  wire d438fc;
  wire v37229e0;
  wire v3a63b7a;
  wire v3a5b109;
  wire v377619b;
  wire v375fda5;
  wire v3a6f911;
  wire v373628e;
  wire v376435f;
  wire v3a5f4b1;
  wire v3a702cb;
  wire v3760881;
  wire v374aacc;
  wire v3a711cb;
  wire v3724b8c;
  wire v377eab7;
  wire v374a79e;
  wire v3a70de5;
  wire v376eeb3;
  wire v3739e4f;
  wire v372552c;
  wire v37277ab;
  wire v3a7026e;
  wire v3779ba9;
  wire v377a525;
  wire v374f252;
  wire v375e0e3;
  wire v3a6f3c6;
  wire v37681ed;
  wire v3a63299;
  wire v373ad16;
  wire v3a65762;
  wire v3745bdf;
  wire v3a61cb2;
  wire v3a6f43a;
  wire v3750fbb;
  wire v376a97b;
  wire v3a5bac7;
  wire v374ed52;
  wire v3a6fb52;
  wire v3a5b310;
  wire v3a66fd9;
  wire v3777536;
  wire v374decf;
  wire v3728793;
  wire v37272ca;
  wire v372e244;
  wire v374d0e3;
  wire v3a64b0f;
  wire v3a7068a;
  wire v3a6002a;
  wire v377d58d;
  wire v3a6628b;
  wire v3a53d12;
  wire v377b946;
  wire v377e85a;
  wire v3754e78;
  wire v3753526;
  wire v3a6eb0a;
  wire v3733b77;
  wire v3745828;
  wire v37413b6;
  wire v3a6eb47;
  wire v3a55f2b;
  wire v3a552c9;
  wire v374852b;
  wire v3749d3f;
  wire v3737d3f;
  wire v3a6efe2;
  wire v3a70168;
  wire v3724fdb;
  wire v3a7090f;
  wire v37572af;
  wire v3a61c1f;
  wire v3a61734;
  wire v3a71202;
  wire v3755731;
  wire v3751ffd;
  wire v3765c49;
  wire v3a70e77;
  wire v37508c2;
  wire v37c3782;
  wire beaea1;
  wire v3758abd;
  wire v375cb51;
  wire v3a57cc8;
  wire v3765f5c;
  wire v3749a6b;
  wire v373e2d3;
  wire v3a70275;
  wire v3a663b9;
  wire v3758a92;
  wire v3a7040e;
  wire v373e891;
  wire v3a6fd9b;
  wire v37745e9;
  wire v3735d84;
  wire v3770edc;
  wire v3a5f6a8;
  wire v3a64539;
  wire v3a70e90;
  wire v376e160;
  wire v3734585;
  wire v3758bc2;
  wire v3a70771;
  wire v1e37405;
  wire v3a6c4c3;
  wire v3a70f0c;
  wire v3774b66;
  wire v3774eed;
  wire v376ad04;
  wire v3a6fbcb;
  wire v3a6d2d7;
  wire v3a64e3e;
  wire v3750ff0;
  wire v3a6209f;
  wire v373b17e;
  wire v3732a04;
  wire v3a5dc5c;
  wire v3a6f931;
  wire v377d831;
  wire v373c15e;
  wire v3779955;
  wire v3a6edab;
  wire v376bade;
  wire v37605bb;
  wire v3752831;
  wire v3a712da;
  wire v374401a;
  wire v3744adf;
  wire v3a70188;
  wire v37671b7;
  wire v3a54dfa;
  wire v374ca4a;
  wire v375e854;
  wire v376a480;
  wire v372713b;
  wire v372a417;
  wire v3806636;
  wire v3757e93;
  wire v3750b29;
  wire v3a702e3;
  wire v3759284;
  wire v3a6fe61;
  wire v3a70e4a;
  wire v3a5d55b;
  wire v3a64994;
  wire v3809093;
  wire v3a5cb68;
  wire v3809516;
  wire v373e7d9;
  wire v376cad6;
  wire v3760d8d;
  wire v3a6ab69;
  wire v3731f08;
  wire v3765219;
  wire v8fffa6;
  wire v376b11e;
  wire v377086b;
  wire v376747e;
  wire v3749840;
  wire v3745eb8;
  wire v37305c2;
  wire v3a71048;
  wire v23fe312;
  wire v37438c9;
  wire v377665f;
  wire v3a55b2d;
  wire v372eae4;
  wire v3768ef1;
  wire v3754ec0;
  wire v374bc27;
  wire v3a5c127;
  wire v37672c8;
  wire v375115e;
  wire v9b03cc;
  wire v3a62245;
  wire v3763f13;
  wire v372494a;
  wire v376c028;
  wire v3a54769;
  wire v373d89b;
  wire v3746b0c;
  wire v3a70cac;
  wire v3a6d434;
  wire v3762d26;
  wire v3a61a7f;
  wire v3741039;
  wire v373a876;
  wire v3737aee;
  wire v373bce7;
  wire v3a70a12;
  wire v3a70c94;
  wire v374197c;
  wire v376d793;
  wire v3a707bb;
  wire v373b0a4;
  wire v3a5a985;
  wire v3744cea;
  wire v37477dd;
  wire v3a67ec4;
  wire v3a5f75a;
  wire v3740a38;
  wire v3730451;
  wire v373d8f2;
  wire v3a710d9;
  wire v377204f;
  wire v37467be;
  wire v377a0d8;
  wire v3a7012b;
  wire v360bc74;
  wire v3a70586;
  wire v374fa11;
  wire v3a70727;
  wire v3749503;
  wire v375fc73;
  wire v377d97d;
  wire v372b4d8;
  wire v3a581bd;
  wire v3a6891e;
  wire v3a6bddd;
  wire v372fe5f;
  wire v3779fec;
  wire v3731399;
  wire v3742d54;
  wire v373e962;
  wire v3a702bc;
  wire v372e798;
  wire v3735d39;
  wire v3a6f88b;
  wire v37510e0;
  wire v357732f;
  wire v380887a;
  wire v3736141;
  wire v3a6ca99;
  wire v376be4c;
  wire v372da76;
  wire v3726d97;
  wire v3a6fa2c;
  wire v3a704f2;
  wire v375f302;
  wire v377dd65;
  wire v37266c2;
  wire v373a9ee;
  wire v37590a2;
  wire v3807b28;
  wire v3a71196;
  wire v3761e45;
  wire v3a65680;
  wire v3774e7b;
  wire v39eaae4;
  wire v3a7051e;
  wire v35b7092;
  wire v37777d5;
  wire v3a7102f;
  wire v372def9;
  wire v375fe83;
  wire v3a6ff9a;
  wire v372c5bc;
  wire v3756ff6;
  wire v37508df;
  wire v372de63;
  wire v37501e6;
  wire v3771232;
  wire v23fe0bb;
  wire v3a6c5ee;
  wire v3a6b8a2;
  wire v3768062;
  wire v3762389;
  wire v373e760;
  wire v3a57959;
  wire v37567d3;
  wire v37565a5;
  wire v3a6b15d;
  wire v3727713;
  wire v3a7056c;
  wire v3a70c7a;
  wire v372e863;
  wire v23fd83f;
  wire v2acb0a5;
  wire v38099e8;
  wire v376f7a7;
  wire v3a6c63e;
  wire v3757ec4;
  wire v380733a;
  wire v3a5fb00;
  wire v943e48;
  wire v37314b5;
  wire v37fc910;
  wire v37413d8;
  wire v3763209;
  wire v375e815;
  wire v373e4db;
  wire v3a63873;
  wire v3747ac9;
  wire v3806e34;
  wire v3a5a7fd;
  wire v373d4ff;
  wire v917087;
  wire v37697ba;
  wire v3a6210a;
  wire v375afc7;
  wire v3761ba8;
  wire v3a5a0d2;
  wire v375d2b3;
  wire v3739ec6;
  wire v374fac7;
  wire v1e37cc1;
  wire v3a6f158;
  wire v3738750;
  wire v376891a;
  wire d2e9f6;
  wire v3a5d6c6;
  wire v3a6f0be;
  wire v3a70cb1;
  wire v3a6e50e;
  wire v3a6ffbd;
  wire v3757cd6;
  wire v3729c45;
  wire v3748481;
  wire v374f76a;
  wire v37538e1;
  wire v3a708c2;
  wire v373184e;
  wire v374212e;
  wire v3a7150e;
  wire v3a710a2;
  wire v3a68f4f;
  wire v372952e;
  wire v3a69a39;
  wire v3a708cf;
  wire v3a648c3;
  wire v375969d;
  wire v3a6fb62;
  wire v3a61cbf;
  wire v3a70715;
  wire ae0781;
  wire v3a6fffc;
  wire v3756057;
  wire v3a711fc;
  wire v3a64cfa;
  wire v377598f;
  wire v374baea;
  wire v372de1e;
  wire v3a5f992;
  wire v374544c;
  wire v3a64a09;
  wire v373026e;
  wire v3731aaf;
  wire v35b77ae;
  wire v375f3ac;
  wire v3a64b90;
  wire v37591f3;
  wire v37476bd;
  wire v372bae3;
  wire v377682b;
  wire v372cec6;
  wire v3756737;
  wire v376a052;
  wire v3a70481;
  wire v3a6e7d8;
  wire v37713fe;
  wire v377c931;
  wire v3a6f1b7;
  wire v972988;
  wire v373547f;
  wire v3a70cc7;
  wire v3a567ea;
  wire v23fd89c;
  wire v375538e;
  wire v3a572e2;
  wire v3a60f1a;
  wire v375ad79;
  wire v3757e32;
  wire v3a70ddd;
  wire v373d66c;
  wire v377a369;
  wire v374c5fc;
  wire v376b72d;
  wire v3778e3f;
  wire v37602c4;
  wire v375da55;
  wire v3a5db58;
  wire v3a65671;
  wire v1e37397;
  wire v374cef4;
  wire v3753a34;
  wire v3736ae5;
  wire v3a6eee7;
  wire v92391b;
  wire v3746444;
  wire v3765734;
  wire v3a593ee;
  wire v377836a;
  wire v375bd8a;
  wire v374d836;
  wire v3746824;
  wire v374a266;
  wire v3a706df;
  wire v3a70a88;
  wire v37560c7;
  wire v8c0e15;
  wire v3a5e9d3;
  wire v372a399;
  wire v3730946;
  wire v376c06f;
  wire v3a6f4ac;
  wire v374acbe;
  wire v373c9b1;
  wire v37672a5;
  wire v37606ba;
  wire v3a70dbe;
  wire v3a713ec;
  wire v374b37d;
  wire v372946e;
  wire v3756304;
  wire v373ac08;
  wire v3a5fcbc;
  wire v375ddb7;
  wire v3a5c700;
  wire v372a6c2;
  wire v3a6f3ad;
  wire v3731ffc;
  wire v3749b37;
  wire v377aa23;
  wire v3775d04;
  wire d305e8;
  wire v376498f;
  wire v374d88f;
  wire v3a6261b;
  wire v37695b1;
  wire v376f0fb;
  wire v3725506;
  wire v3769bcb;
  wire v3a65d01;
  wire v3753456;
  wire v3760a55;
  wire v3a64b83;
  wire v37621eb;
  wire v3742a27;
  wire v3a6a295;
  wire v377cccb;
  wire v372c3d7;
  wire v375cddb;
  wire v377291b;
  wire v376c0c8;
  wire v3a70c4b;
  wire v3a6eb46;
  wire v3740646;
  wire v373ad3c;
  wire v377a63c;
  wire v376f332;
  wire v375588c;
  wire v3735525;
  wire v373dfb8;
  wire v3754877;
  wire v375c946;
  wire v373a568;
  wire v3725360;
  wire v3a55efa;
  wire v377d3b9;
  wire v37729db;
  wire v373fd50;
  wire v37697a3;
  wire v376a297;
  wire v3728d72;
  wire v373e6cf;
  wire v3a70995;
  wire v372ea4b;
  wire v3a6d03c;
  wire v3726979;
  wire v37485ce;
  wire v37429e5;
  wire v376b540;
  wire v3740762;
  wire v3737e2c;
  wire v3768a9c;
  wire v3a7074e;
  wire v3a5395c;
  wire v3a6708d;
  wire v3778138;
  wire v375cb14;
  wire v3807a2e;
  wire v3a6ff99;
  wire v3753a2e;
  wire v3a70961;
  wire v3a6eebd;
  wire v3773838;
  wire v3a674c2;
  wire v375a261;
  wire v3754a42;
  wire v3a53873;
  wire v3723b5b;
  wire v3778d7f;
  wire v374d778;
  wire v374d969;
  wire v374e21e;
  wire v37402b8;
  wire v3773ab1;
  wire v3773ccd;
  wire v37679f0;
  wire v3a5d6f3;
  wire v3a70e54;
  wire v3a651c8;
  wire v3764a6c;
  wire v3770a5a;
  wire v37402d8;
  wire v372a465;
  wire v3a70d2a;
  wire v3a61149;
  wire v37276a0;
  wire v380735e;
  wire v3a701ee;
  wire v376e87e;
  wire v3a6fda1;
  wire v3a5414c;
  wire v37325c5;
  wire v375d95f;
  wire v37515a1;
  wire v3774a4b;
  wire v3a6e29d;
  wire v3757e56;
  wire v3a6f232;
  wire v3a58dfb;
  wire v3751141;
  wire v3a6f212;
  wire v376c0dc;
  wire v3a5ba5b;
  wire v376752b;
  wire v373a57d;
  wire v3a71076;
  wire v37523f8;
  wire v3774cf5;
  wire v37750a5;
  wire v3723025;
  wire v3753fe3;
  wire v3a62dae;
  wire v3774664;
  wire v3a70795;
  wire v3779e9b;
  wire v3732b30;
  wire v3739d2c;
  wire v376d795;
  wire v3753b70;
  wire v3761f69;
  wire v3a6a52c;
  wire v3a64a5d;
  wire v3a57f04;
  wire d3a24d;
  wire v373945c;
  wire v3a6eeb7;
  wire v37610ce;
  wire v3a550e2;
  wire v3a7021a;
  wire v3763e92;
  wire v374eec1;
  wire v3808e88;
  wire a80fe2;
  wire v375c144;
  wire v372aaf8;
  wire v3a6ddc7;
  wire v3a6f6f2;
  wire v3a711be;
  wire v377b481;
  wire v37336b4;
  wire v3a7050f;
  wire v373e2f2;
  wire v376456d;
  wire v37713e8;
  wire v374797c;
  wire v3a70f0d;
  wire v372bcd3;
  wire v37484ac;
  wire v3a63f7b;
  wire v3745d1e;
  wire v3759532;
  wire v3a5f205;
  wire v376956a;
  wire v372d98c;
  wire v3a5565d;
  wire v372b923;
  wire v374333e;
  wire v3728455;
  wire v3a68916;
  wire v3a5d8d3;
  wire v3758bcd;
  wire v3a5d065;
  wire v3733a4c;
  wire v3764684;
  wire v3a6f7b3;
  wire v373124d;
  wire v3734a4f;
  wire v375194a;
  wire v374e873;
  wire v372fcfc;
  wire v3743b2f;
  wire v37741d7;
  wire v3a6cce9;
  wire v375ece3;
  wire v37370c6;
  wire c48c9d;
  wire v3a6e6c2;
  wire v376b374;
  wire v372baf1;
  wire v376a9f7;
  wire v375dd92;
  wire v3776f7d;
  wire v3767b2e;
  wire v376dcf6;
  wire v3a5d4e9;
  wire v37264a3;
  wire v376053f;
  wire v3a5c4c6;
  wire v376c25c;
  wire v37494c3;
  wire v37548e9;
  wire v37359cb;
  wire v3a648c8;
  wire v3766472;
  wire v3772ac1;
  wire v3a6fa69;
  wire v3a7140f;
  wire v3772bda;
  wire v3734914;
  wire v375524c;
  wire v3a62eee;
  wire v376a47b;
  wire v3a6fab1;
  wire v3739eed;
  wire v374752b;
  wire v23fe345;
  wire v3747587;
  wire v3a6e4b8;
  wire v3749e61;
  wire v3733249;
  wire v3a5d153;
  wire v37342ec;
  wire v3776479;
  wire v373fb1a;
  wire v3a6f569;
  wire v3722bb0;
  wire v37741f0;
  wire v377a12e;
  wire v3a6fb06;
  wire v373e587;
  wire v3740953;
  wire v374f359;
  wire v3a6f8a9;
  wire v3a7162f;
  wire v37540dd;
  wire v3757f54;
  wire v3a5eae2;
  wire v3a67f58;
  wire v376158e;
  wire v3728435;
  wire a740cc;
  wire v37372eb;
  wire v375c3b6;
  wire v377817b;
  wire v377e59a;
  wire v3747fda;
  wire v3743fc1;
  wire v3747b97;
  wire v373a0d6;
  wire v3a6e81d;
  wire v1e37c60;
  wire v375652a;
  wire v37630a8;
  wire v3776066;
  wire v3a60509;
  wire v372e741;
  wire v373ec83;
  wire v375075b;
  wire v37758de;
  wire v3a60134;
  wire v3745941;
  wire v3a70e47;
  wire v37300e3;
  wire v37530e8;
  wire v376bfb9;
  wire v3766986;
  wire v377d4e1;
  wire v377bd9b;
  wire v372ff09;
  wire v3761334;
  wire v3744838;
  wire v3750b9d;
  wire v3773cda;
  wire v3766445;
  wire v3a71656;
  wire v3731a95;
  wire v37305e6;
  wire v3a6cd4f;
  wire v3a5e611;
  wire v376957a;
  wire v380910e;
  wire v3756ba5;
  wire v37294a9;
  wire v3764d3e;
  wire v3759c48;
  wire v3739dfa;
  wire v3762dd5;
  wire v3a6fe04;
  wire v3a711cf;
  wire v374407e;
  wire v37776f0;
  wire d193f7;
  wire v372f2ff;
  wire v3a710f8;
  wire v374990a;
  wire v3a69fe0;
  wire v37542a0;
  wire v3729972;
  wire v375fac2;
  wire v3a70577;
  wire v3a6fd41;
  wire v37426ea;
  wire v375970d;
  wire v374caf9;
  wire v3a70ce8;
  wire v3a5f458;
  wire v37557c6;
  wire v3745ee1;
  wire v3a70a46;
  wire v3a6ebdc;
  wire v3a6eb72;
  wire v3758c13;
  wire v3a70859;
  wire v37535fd;
  wire v37712aa;
  wire v3743bde;
  wire v375bcf7;
  wire v37529f6;
  wire v3a638f4;
  wire v3a71264;
  wire v3806c70;
  wire v3a5aa93;
  wire v3a70170;
  wire v374335b;
  wire a56488;
  wire v3a70749;
  wire v3771076;
  wire v375bf61;
  wire v3a6fa2d;
  wire v3762ca6;
  wire v372e374;
  wire v372a027;
  wire v3778d73;
  wire v3a58687;
  wire v3a5a9e6;
  wire v3742c68;
  wire v3a7085c;
  wire v3a58306;
  wire v3752f8e;
  wire v3775903;
  wire v372437d;
  wire v3740a94;
  wire v37503f5;
  wire v3779f68;
  wire v3a70d6d;
  wire v3768070;
  wire v3a56ba2;
  wire v3772318;
  wire v374c9e4;
  wire v3731e55;
  wire v375ceb9;
  wire v3a69391;
  wire v3723db5;
  wire v3a6fb8b;
  wire v372a48e;
  wire v3808ceb;
  wire v3a63777;
  wire v3a709b4;
  wire v3772e8e;
  wire v3a70638;
  wire v3a67eb4;
  wire v3723740;
  wire a50cea;
  wire v3a6f529;
  wire v374e016;
  wire v3a6efb0;
  wire v3a6f5e8;
  wire v376e240;
  wire v3a62d59;
  wire v3a6f0a2;
  wire v3a6fe48;
  wire v3771667;
  wire c2c2bc;
  wire v37447e2;
  wire v373eaee;
  wire v377564e;
  wire v373ac12;
  wire v372e661;
  wire v373855c;
  wire v3a5d079;
  wire v3a5e827;
  wire a19873;
  wire v373a7a5;
  wire v374bfa6;
  wire v376502e;
  wire v373301a;
  wire v37692dc;
  wire v9aa32c;
  wire v3a6f873;
  wire v3773e8d;
  wire v37770df;
  wire v37775c7;
  wire v375f0de;
  wire v37596a6;
  wire v374127d;
  wire v3a60649;
  wire v3745202;
  wire v2ff8e74;
  wire v37476c2;
  wire v375e035;
  wire v3a675bc;
  wire v3a58674;
  wire v37487f7;
  wire v372dde7;
  wire v3a6af0b;
  wire v3733c9e;
  wire v3a6162f;
  wire v3a5f78a;
  wire v3258dc5;
  wire v3a6ebc7;
  wire v3743a8a;
  wire v377cf34;
  wire v3739493;
  wire v3a6f31e;
  wire v3776e45;
  wire v376723e;
  wire v372e9b1;
  wire v3a714fe;
  wire v3a6e8db;
  wire v3779014;
  wire v2aca987;
  wire v3a5dd8a;
  wire v375a251;
  wire v3774247;
  wire v3764306;
  wire v3a6f608;
  wire v374930c;
  wire v377d302;
  wire v37752af;
  wire v37338bb;
  wire v3730688;
  wire v3a62113;
  wire v3a62f50;
  wire v3763478;
  wire v376b044;
  wire v3a65b42;
  wire v376da5f;
  wire v375585a;
  wire v372c97c;
  wire v37657be;
  wire v3726da1;
  wire v372e537;
  wire v37248e4;
  wire v3735fc0;
  wire v37796ee;
  wire v3a705dd;
  wire v372aefc;
  wire v3a63203;
  wire v376a21e;
  wire v37533ea;
  wire v3768751;
  wire v37473ca;
  wire v3a70ff1;
  wire v373d7ea;
  wire v3a6d1b9;
  wire v3a70891;
  wire v3743726;
  wire v375733e;
  wire v374eac6;
  wire v37325cf;
  wire v3a6e3f0;
  wire v373bfea;
  wire v3a555d1;
  wire v3a59264;
  wire v3806f19;
  wire v3752767;
  wire v3a5dd62;
  wire b95629;
  wire v37612d4;
  wire v372d9b0;
  wire v375d059;
  wire v3a5ae95;
  wire v374e843;
  wire v3a71134;
  wire v372883e;
  wire v373ad7b;
  wire v3764ed7;
  wire v376072e;
  wire v377fc51;
  wire v3759be3;
  wire v375cf7d;
  wire v3a651fc;
  wire v3a5836e;
  wire v376d62b;
  wire v377c068;
  wire v3729cbe;
  wire v3774acc;
  wire v380956e;
  wire v375aea6;
  wire v372952d;
  wire v372af57;
  wire v3723dac;
  wire v373d12a;
  wire v3a71526;
  wire v376c5b4;
  wire v3723bac;
  wire v372e88f;
  wire v3724859;
  wire v376819e;
  wire b2eec3;
  wire v3740469;
  wire v3773434;
  wire v372b847;
  wire v2092be1;
  wire v377fada;
  wire v373f1ac;
  wire v3a595ba;
  wire v374fafa;
  wire v3776e8b;
  wire v373ab15;
  wire v3726f2e;
  wire v3a6b53f;
  wire v37674a3;
  wire v37790fb;
  wire v37618ad;
  wire v374875d;
  wire v3a6f10e;
  wire a9c905;
  wire v377f171;
  wire v3a70704;
  wire v3a5a051;
  wire v3742a62;
  wire v3a6bf12;
  wire v3744117;
  wire v376f5b3;
  wire v3a6efb2;
  wire v374b8c5;
  wire v3a616ad;
  wire v3a70c2c;
  wire v3a5e2eb;
  wire v375b880;
  wire v376166b;
  wire v3764552;
  wire v3a61e9a;
  wire v377a002;
  wire bbcc5e;
  wire v3807a26;
  wire v3727b10;
  wire v3727c91;
  wire v37280a3;
  wire v37652d4;
  wire v3766792;
  wire v3763550;
  wire v3728f6d;
  wire v3777d37;
  wire v3729bc6;
  wire v372cb8c;
  wire v37719a0;
  wire v3729988;
  wire v3a5c9d3;
  wire v3a704f5;
  wire v37750e4;
  wire v373ab60;
  wire v3a702fc;
  wire v3a70433;
  wire v3733483;
  wire v3a6673e;
  wire v375d7d2;
  wire v375a0af;
  wire v3a5c2ff;
  wire v3a6e927;
  wire v3772347;
  wire v38072a2;
  wire v3726023;
  wire v3a54466;
  wire v3a64a14;
  wire v375f55e;
  wire v377241f;
  wire v3779b3a;
  wire v3a70220;
  wire v3730094;
  wire v3a6cf88;
  wire v9fecca;
  wire v3a6eca6;
  wire v375d4de;
  wire v3734fc3;
  wire v3a58be6;
  wire v3766298;
  wire v3743057;
  wire v372d2cd;
  wire v37529d6;
  wire v3a5f358;
  wire v377b73b;
  wire v3725c95;
  wire v376baad;
  wire v3808e9f;
  wire v37632c3;
  wire v37311da;
  wire v3a70c75;
  wire v3735b0b;
  wire v37670db;
  wire v3a6d4f3;
  wire v376e1d4;
  wire v372610c;
  wire v3a700be;
  wire v3773f27;
  wire v377375f;
  wire v3732a31;
  wire v374e9d1;
  wire v3a70665;
  wire b8f5a8;
  wire v3771c38;
  wire v3769639;
  wire v3743dce;
  wire v3752215;
  wire v376fddc;
  wire v3a5e0e5;
  wire v376b56b;
  wire v3a2a0f9;
  wire v3a5c3ef;
  wire v37431ac;
  wire v3a702bd;
  wire v3763364;
  wire v3a64608;
  wire v3730c96;
  wire v3a62403;
  wire v3a6de83;
  wire v3a7159f;
  wire v3a671f2;
  wire v3a6f25b;
  wire v374dabc;
  wire v3a615f5;
  wire v375f69e;
  wire v376c5d3;
  wire v3a58bae;
  wire v3761b23;
  wire v3a706ea;
  wire v372c20d;
  wire v3750857;
  wire v376df68;
  wire v3764f2d;
  wire v3a6f5e7;
  wire v3a71368;
  wire v3a6fec1;
  wire v3a71180;
  wire v3771e69;
  wire v3a6094b;
  wire v3a6b8e8;
  wire v374705f;
  wire v3a7071f;
  wire v3762230;
  wire v3a5bc76;
  wire v3807748;
  wire v3742395;
  wire v3740f94;
  wire v373809d;
  wire v3747fdb;
  wire v376784b;
  wire v3735760;
  wire v375a0ad;
  wire v3765998;
  wire v375b801;
  wire v3735a7f;
  wire v3758524;
  wire v3758561;
  wire v3a700d7;
  wire v3752fcb;
  wire v3a5d8e0;
  wire v3756a6a;
  wire v292554f;
  wire v3727960;
  wire v3a57801;
  wire v3a65afd;
  wire v3742676;
  wire v3741418;
  wire v3a6fe07;
  wire v3769870;
  wire v377b5f4;
  wire v374a8db;
  wire v377f1ff;
  wire v376445f;
  wire v3a57ee9;
  wire v3743d5d;
  wire v3a70ccd;
  wire v375caa2;
  wire v3756200;
  wire v377034f;
  wire v373a0f8;
  wire v3a5cf57;
  wire v374e00b;
  wire v372911f;
  wire v3a6ac20;
  wire v3748489;
  wire v374e784;
  wire v3a6fe2d;
  wire v9375a3;
  wire v3772a15;
  wire v3a6f45d;
  wire v372f3a4;
  wire v37369d7;
  wire v3755aca;
  wire v37693a3;
  wire v3a6fe6f;
  wire v3a6094e;
  wire v375316c;
  wire v374e179;
  wire v37380be;
  wire v3726240;
  wire v3757ebc;
  wire v3a6b0eb;
  wire v3744824;
  wire v375521a;
  wire v3726654;
  wire v3770b24;
  wire v3748472;
  wire v374b228;
  wire v3a7113d;
  wire v3a68f22;
  wire v3744f1e;
  wire v3724f54;
  wire v3769510;
  wire v3731304;
  wire v3a6fc0b;
  wire v376ca86;
  wire v37386c6;
  wire v3a68482;
  wire v3a6ec20;
  wire v375eb1b;
  wire v3755f80;
  wire v373f19e;
  wire v3a5b909;
  wire v3a6b4fb;
  wire v3761cec;
  wire v3738397;
  wire v377d8dd;
  wire bdda12;
  wire v3769404;
  wire v37609ac;
  wire v372da4f;
  wire v373c480;
  wire v375b736;
  wire v3a708b9;
  wire v3a676a9;
  wire v373fc8a;
  wire v3a6f0b8;
  wire v37368b3;
  wire v372456c;
  wire v3752cf6;
  wire v3a646ae;
  wire v3a6d840;
  wire v372f76c;
  wire v3a70c72;
  wire v372b881;
  wire v3761d47;
  wire v372cdb0;
  wire v3a61517;
  wire v3732c86;
  wire v380925f;
  wire v37523ef;
  wire v2ff8f33;
  wire v3765b5c;
  wire v3a53392;
  wire v3a63f6b;
  wire v3749f3b;
  wire v373d25a;
  wire v373e0b5;
  wire v374a0f0;
  wire v3a6123e;
  wire v3776b61;
  wire v3736cc7;
  wire v377844d;
  wire v375767e;
  wire v3759ffd;
  wire v3a70b5d;
  wire v3a70ee1;
  wire v3a70ba7;
  wire v372b44a;
  wire v3a6582b;
  wire v3a70753;
  wire v3a70f18;
  wire v3764ced;
  wire v3753030;
  wire v3a70f53;
  wire v375c366;
  wire v3a53ed2;
  wire v3757537;
  wire v37319c5;
  wire v3a70e5e;
  wire v377b647;
  wire v374ef3e;
  wire v3765224;
  wire v3779863;
  wire v3a53cc2;
  wire v376dc2e;
  wire v3774494;
  wire v3a7126a;
  wire v376b269;
  wire v3a66f81;
  wire v373dd9b;
  wire v3a60faf;
  wire v3a538b9;
  wire v375c791;
  wire v373d7e9;
  wire v3753542;
  wire ad187c;
  wire v3771502;
  wire v3a5a647;
  wire v3a714f5;
  wire v3a5ef54;
  wire v3a6d5b3;
  wire d8a75b;
  wire v3732817;
  wire v3741d00;
  wire v3a707de;
  wire v3736c94;
  wire v374059d;
  wire v374ace7;
  wire v375bebd;
  wire v375d84b;
  wire v3726006;
  wire v3769616;
  wire v376ab72;
  wire v3771e95;
  wire v3a6a393;
  wire d9a7db;
  wire v3a7047e;
  wire v37537ef;
  wire v37372c9;
  wire v3759ca7;
  wire v3770cf6;
  wire v3756483;
  wire v38073c9;
  wire v374a4ca;
  wire v3728823;
  wire v3a70eff;
  wire v3a6ebf6;
  wire v3a6500c;
  wire v373c3e4;
  wire v377b4fb;
  wire v372f3f7;
  wire v2092b23;
  wire v376942f;
  wire v3809259;
  wire v3733103;
  wire v3a6ec17;
  wire v372e4de;
  wire v3758a9c;
  wire v3752002;
  wire v3a705e8;
  wire v3a6dcb9;
  wire v3a62968;
  wire v375a4ea;
  wire v3a57ebf;
  wire v375f619;
  wire v3a685db;
  wire v3a55eda;
  wire v372cd65;
  wire v376f09b;
  wire v375822b;
  wire v3730b1c;
  wire v3722b10;
  wire v3a67b58;
  wire v3a6ffe9;
  wire v3776395;
  wire v3772d2f;
  wire v37764b1;
  wire v3a5ce2d;
  wire v3758225;
  wire v375c707;
  wire v37621ee;
  wire v3724c95;
  wire v3758e5f;
  wire v372d880;
  wire v376aa7a;
  wire v3a6f48f;
  wire v37415b2;
  wire v3750547;
  wire v3a6ec6d;
  wire v37440a8;
  wire v3378594;
  wire v3a57b70;
  wire v3a70791;
  wire v377eaa3;
  wire v3a70532;
  wire v3728a76;
  wire b65b94;
  wire a96343;
  wire v3a60b90;
  wire v3a5e9b8;
  wire v3a6febe;
  wire v3754d28;
  wire v377c236;
  wire v3a6a8b2;
  wire b2d8a6;
  wire v3765f12;
  wire v376e663;
  wire v3769e46;
  wire v3a704c3;
  wire v3766101;
  wire v3769023;
  wire v373623d;
  wire v3a707f0;
  wire v3766462;
  wire v3748d2f;
  wire v3728c14;
  wire v3a7107f;
  wire v3a71525;
  wire v3a5d32a;
  wire v3769982;
  wire v3756bd8;
  wire v3a70cc8;
  wire v37604fe;
  wire v3a6fe50;
  wire v375b389;
  wire v3a6c527;
  wire v3729d8d;
  wire v3759f61;
  wire v37522bc;
  wire v3a70376;
  wire v3a6f1c5;
  wire v3a6f02e;
  wire v3a71145;
  wire v3762fc2;
  wire v374cba0;
  wire v35b708f;
  wire v377e26b;
  wire v373abb7;
  wire v3a702a7;
  wire v373120c;
  wire v3763af8;
  wire v375f6ef;
  wire v377e8da;
  wire v3a70d0f;
  wire v376c1e4;
  wire v3729280;
  wire v3733a5f;
  wire v3a53e66;
  wire v376397d;
  wire v37662d3;
  wire v373c219;
  wire v3775293;
  wire v377661c;
  wire v3738602;
  wire v3a5c462;
  wire v3735dae;
  wire v3a6d4f9;
  wire v373d10f;
  wire v3a70511;
  wire v325b5df;
  wire v37648f2;
  wire v3a56d2d;
  wire v37248fd;
  wire v3a66d50;
  wire v377cc27;
  wire b0f188;
  wire v373ed9a;
  wire v374fae5;
  wire v3a7062b;
  wire v3a7134d;
  wire v3a71088;
  wire v37452c7;
  wire v3760e46;
  wire v3748353;
  wire v3754b98;
  wire v3749d78;
  wire v3772567;
  wire v374ba61;
  wire v3a6632a;
  wire v3768af7;
  wire v3726c20;
  wire v3a7114b;
  wire v3a5ddaa;
  wire v373511d;
  wire v3749969;
  wire v3a67d8d;
  wire v375107e;
  wire v3a63d22;
  wire v374ff15;
  wire v372c863;
  wire v3807a4a;
  wire v373f4fb;
  wire v375c3eb;
  wire v373cdd5;
  wire v3739bcb;
  wire v3a702b3;
  wire v3a6f52c;
  wire v373185f;
  wire v377f401;
  wire v3734788;
  wire v3740c75;
  wire v372e474;
  wire v373aa23;
  wire v3a697f2;
  wire v375024d;
  wire v3750e9a;
  wire v3a6f1fd;
  wire v372802c;
  wire v3a6ebf0;
  wire v3742101;
  wire v377ad8f;
  wire v3809865;
  wire cf6441;
  wire v375d009;
  wire v3757955;
  wire v376121f;
  wire v376aeae;
  wire v38090f6;
  wire v375de7f;
  wire v3753923;
  wire v3a6d299;
  wire v374291b;
  wire v37519ea;
  wire v3a709ba;
  wire v3a6fba8;
  wire v3a70b5f;
  wire v3a708fd;
  wire bc9e23;
  wire v37777bf;
  wire v376129a;
  wire v3a6ad19;
  wire v376a7fc;
  wire v3766e5d;
  wire v3752c29;
  wire v3a6d3f3;
  wire v3727615;
  wire v374cd10;
  wire v3a67dbc;
  wire v3729e32;
  wire v3a6f8f7;
  wire v3a70b91;
  wire v373b14a;
  wire v3775e66;
  wire v3a705f7;
  wire v39a5350;
  wire v377b515;
  wire v3a6fac4;
  wire v86d3dc;
  wire v3770855;
  wire v3a638fe;
  wire v3a5dbc7;
  wire v3a63e87;
  wire v3a70b0e;
  wire v372d336;
  wire v3a70e19;
  wire v3a6dc38;
  wire v3a60b96;
  wire v3807113;
  wire v3742f0a;
  wire v3a70caa;
  wire v3a6934e;
  wire v3a630b7;
  wire v3a691f2;
  wire v3a70083;
  wire v373427f;
  wire v3a6567f;
  wire v3a7126e;
  wire v3a6f28a;
  wire v3775508;
  wire v377e692;
  wire v3a70033;
  wire v37606e1;
  wire v3a5a1ef;
  wire v3a70398;
  wire v37444d4;
  wire v3a6ef6f;
  wire v37620b4;
  wire v3a6574d;
  wire v37725b5;
  wire v33790a4;
  wire v23fda78;
  wire v3a6fa02;
  wire v3a5b4ca;
  wire v3a70ed5;
  wire v3732c96;
  wire v37514f1;
  wire v373055b;
  wire v372b7e6;
  wire v3a7066d;
  wire v3769384;
  wire v37688d1;
  wire v376c422;
  wire d73f1d;
  wire v37333de;
  wire v376cd09;
  wire v374b564;
  wire v3725403;
  wire v23fe0ff;
  wire v3740bf7;
  wire v376a252;
  wire v3a6fd20;
  wire v3a6fe10;
  wire v325c974;
  wire v376438f;
  wire v3809542;
  wire cbc7dd;
  wire v37365f8;
  wire v3a669be;
  wire v3a70f4f;
  wire v3763046;
  wire v376fbce;
  wire v3a6dac0;
  wire v377c97f;
  wire v37646a9;
  wire v3725b77;
  wire v3a71679;
  wire v3a60bfb;
  wire v377600d;
  wire v2925cf2;
  wire v375fd99;
  wire v3a695a8;
  wire v375d65c;
  wire v3a692da;
  wire v3a6fd22;
  wire v374eab3;
  wire v3a67965;
  wire v3750eb9;
  wire v3a6ae2f;
  wire v373a6f8;
  wire v3a7138e;
  wire v3a6efb9;
  wire v3759cad;
  wire v3a670d6;
  wire v37577d8;
  wire v3a70544;
  wire v3772a87;
  wire v3a623c7;
  wire v3a6fd48;
  wire v373ea3f;
  wire v3a5e3bb;
  wire v3a6f6e7;
  wire v3757271;
  wire v3758972;
  wire v3a583ee;
  wire v3767429;
  wire v3a6c02f;
  wire v376ab4e;
  wire v3a70bea;
  wire v375c70c;
  wire v3807df0;
  wire v3732355;
  wire bba7f1;
  wire v3a7082a;
  wire v3772596;
  wire v3806388;
  wire v372b373;
  wire v3a6fea8;
  wire v376a2bf;
  wire b4f73f;
  wire v3762c73;
  wire v37372dd;
  wire cc4895;
  wire v3a71569;
  wire v3a57ec9;
  wire v3a70821;
  wire v3a710f3;
  wire v3765740;
  wire v373d5ab;
  wire v376b082;
  wire v3a5b47c;
  wire v37293f6;
  wire v37775eb;
  wire v3a6ba77;
  wire v3a6dbf0;
  wire v3a710f1;
  wire v3a714a2;
  wire v3a6fba6;
  wire v37458d2;
  wire v3a6fc1d;
  wire v3a70b9a;
  wire v3a6984f;
  wire v372f87c;
  wire v3727ff7;
  wire v3765e6a;
  wire v3723f2a;
  wire v3739391;
  wire v376c203;
  wire v377d60e;
  wire v3757863;
  wire v3725f24;
  wire v3a63e9e;
  wire v3751a33;
  wire v374d273;
  wire v3761cbb;
  wire v3778e03;
  wire v372b17b;
  wire v375f71d;
  wire v3a6a116;
  wire v3a5c015;
  wire v377868e;
  wire v3764ca0;
  wire v374e768;
  wire v3a5d06d;
  wire v3a66e41;
  wire v3a6e868;
  wire v3a5e3c0;
  wire v380917f;
  wire v376daf6;
  wire v3a56d0a;
  wire v3723baf;
  wire v3a605f1;
  wire v3a6f722;
  wire v3733bbe;
  wire v39eb452;
  wire v373e4c0;
  wire v3a70dfe;
  wire v3774f35;
  wire v3748b9d;
  wire v376d172;
  wire v3a621e7;
  wire v3760a52;
  wire v3747b15;
  wire v373e38a;
  wire v373a759;
  wire v23fd9e1;
  wire v3a70a89;
  wire v376aaee;
  wire v37416f0;
  wire v375dbeb;
  wire v37521ff;
  wire v3a5e7fd;
  wire v374e06f;
  wire v37233a4;
  wire v373a7a6;
  wire v374c693;
  wire v3738700;
  wire v3753964;
  wire v3a70a45;
  wire v37265b3;
  wire cf3b5d;
  wire v3a65bb5;
  wire v375aae9;
  wire v376c343;
  wire v375b7dc;
  wire v3a69043;
  wire v3a6c7c6;
  wire v3a70688;
  wire v375b0e8;
  wire v377c160;
  wire v37626a4;
  wire v3739da7;
  wire v3a6e6e1;
  wire v3730fc0;
  wire v373f9db;
  wire v373484e;
  wire v3728034;
  wire v376bebb;
  wire v37277c2;
  wire v3735f14;
  wire v37599b1;
  wire a9f810;
  wire v3a55271;
  wire v3a5b563;
  wire v377af64;
  wire v3a6f7c0;
  wire v3723247;
  wire v3a70486;
  wire v37485e0;
  wire v3747704;
  wire v3809958;
  wire v376c883;
  wire v3778fda;
  wire v3a66b88;
  wire v3577338;
  wire v372a94e;
  wire v3772edc;
  wire v3a70405;
  wire v3a7080b;
  wire v377206b;
  wire v3a6fac0;
  wire v3a715b7;
  wire v37590cb;
  wire v3761006;
  wire v376d902;
  wire v374ee8d;
  wire v3747314;
  wire v3779717;
  wire v375af36;
  wire v3a7082c;
  wire v3730a2f;
  wire v3a7108f;
  wire v373187a;
  wire c5fc63;
  wire v372dcf7;
  wire v376c6fb;
  wire v3746540;
  wire v373464d;
  wire v3a71128;
  wire v3a6da6b;
  wire v3a6d71b;
  wire v3a6d407;
  wire v374e5fa;
  wire v3727830;
  wire v3a6d2ed;
  wire v376058c;
  wire v3777362;
  wire v374c8a8;
  wire v3a656a4;
  wire v3731fb9;
  wire v3a706d5;
  wire v3747d33;
  wire v3a55ea1;
  wire v373ed57;
  wire v375a4f6;
  wire v3773a06;
  wire v3a6ffec;
  wire v37472f4;
  wire v3a6dcf3;
  wire v3a71090;
  wire v3779f0a;
  wire v3765442;
  wire v3731455;
  wire v374a543;
  wire v1e378a8;
  wire v3a715e9;
  wire v3a60a84;
  wire v3773078;
  wire v37282f7;
  wire v3a705d4;
  wire v3a6fb43;
  wire v3770733;
  wire v3a6ec88;
  wire v3577487;
  wire v376934b;
  wire v373c334;
  wire v376382f;
  wire v375554d;
  wire v3a70938;
  wire v372838e;
  wire v3a6ed2b;
  wire v376e979;
  wire v377b3bd;
  wire v375e50f;
  wire v3739621;
  wire v375be90;
  wire v3a711b4;
  wire v3a57f7d;
  wire v3a706e6;
  wire v37751c3;
  wire v37352fa;
  wire v376ba2b;
  wire v3a5982a;
  wire v37777d1;
  wire b5394c;
  wire v3a647cd;
  wire v3a5af41;
  wire v3a700e8;
  wire v3743d47;
  wire v377c271;
  wire v37646dc;
  wire v3a70583;
  wire v3765ad4;
  wire v3a69c73;
  wire v3a60ce2;
  wire v3761c4e;
  wire v3730e7d;
  wire v3a5495d;
  wire v3a6f806;
  wire v3a6f15c;
  wire v3774841;
  wire v377cb85;
  wire v375ea58;
  wire v3a62a6d;
  wire v37bfca2;
  wire v37453d7;
  wire v3775782;
  wire v3a6fd2f;
  wire v374c2aa;
  wire v376a65b;
  wire v3751f56;
  wire v377e089;
  wire v3a70fa2;
  wire v372ee9a;
  wire v3774ccf;
  wire v3765a1d;
  wire v374f768;
  wire v3727215;
  wire v3a6be44;
  wire v3a6f6c5;
  wire v3767e47;
  wire v3a6f330;
  wire da0ed3;
  wire v37235f1;
  wire v372bad7;
  wire v37694de;
  wire v377834b;
  wire v3a60395;
  wire v3739021;
  wire v3a6f8de;
  wire v3a68e71;
  wire v37740d0;
  wire v3758d6c;
  wire v3761bd1;
  wire v37591b4;
  wire v3a5a158;
  wire v3775aa7;
  wire v373daa8;
  wire v3742feb;
  wire v3731991;
  wire v3809d9e;
  wire v372a80a;
  wire v3a70630;
  wire v37753b4;
  wire v373c23c;
  wire v373158e;
  wire v373b48c;
  wire v375f906;
  wire v376b3d4;
  wire v3a6f9e9;
  wire v375789e;
  wire v3a57baa;
  wire v3746ed6;
  wire v3a7044e;
  wire v3727f69;
  wire v375a7cd;
  wire v3755dcd;
  wire ce4d7a;
  wire v3750978;
  wire v3729421;
  wire v373c4c2;
  wire v37302f1;
  wire v3775f27;
  wire aed6c7;
  wire v3a70cfb;
  wire v37564e4;
  wire v372ad34;
  wire v374fe8e;
  wire v375400b;
  wire v3a70118;
  wire v3746ea0;
  wire v3807474;
  wire v3a71189;
  wire v3a5c188;
  wire v37350b2;
  wire v37710f3;
  wire v37295a5;
  wire v3a58971;
  wire v375c92f;
  wire v3a6ffd7;
  wire v1e37759;
  wire v3806dc8;
  wire v3770c98;
  wire v377180a;
  wire v37501a3;
  wire v374ef8d;
  wire v3a5c7a3;
  wire v372c483;
  wire v374bbaf;
  wire v37651fe;
  wire v3761fd6;
  wire v377109a;
  wire v3740489;
  wire v3740dcc;
  wire v373635b;
  wire v3a70585;
  wire v3a6fa53;
  wire v37352dc;
  wire v3a56c18;
  wire v372bd5f;
  wire v3a65c31;
  wire v3a6fd36;
  wire v37673e8;
  wire v3a70e53;
  wire v375178a;
  wire v3a6f701;
  wire v3743b64;
  wire v3a71588;
  wire v372a06a;
  wire v37606f0;
  wire v3a5a45e;
  wire v3726a2b;
  wire v9ac541;
  wire v3a6fc3a;
  wire v374fedc;
  wire v375ec51;
  wire v373c6b6;
  wire v39a4df7;
  wire v3a700d4;
  wire v39a4dc7;
  wire v372bee9;
  wire a5d7b0;
  wire v375579f;
  wire v3a707ff;
  wire v3729ffd;
  wire v37244a0;
  wire v375ce35;
  wire v3761719;
  wire v37797ef;
  wire v377efd0;
  wire v374baac;
  wire v3777da6;
  wire v3a5e015;
  wire v3746045;
  wire v35b7299;
  wire v372f72b;
  wire v37433b4;
  wire v3778323;
  wire v3738762;
  wire v3739cda;
  wire v3a640ff;
  wire v3731b41;
  wire v3a5d989;
  wire v3740ad9;
  wire v3777995;
  wire v372648f;
  wire v3730e74;
  wire v3a6ef01;
  wire v3a71254;
  wire v376d3e1;
  wire v373b30b;
  wire v3a6fc68;
  wire v37262ec;
  wire v375fcac;
  wire v375f238;
  wire v3a5fd54;
  wire v38073fd;
  wire v3729b63;
  wire v372d828;
  wire v3a6d621;
  wire v37308b0;
  wire v3751e80;
  wire v3773fc7;
  wire v3a5918c;
  wire v3733d3f;
  wire v3736319;
  wire v3a71558;
  wire v3755420;
  wire v37427e9;
  wire v3766d0a;
  wire v3a6f6c0;
  wire v3a703b0;
  wire v374e8b5;
  wire v3a5d522;
  wire v3a67555;
  wire v3a7047d;
  wire v3726ec0;
  wire v3754227;
  wire v3a63597;
  wire v3a7041e;
  wire v3764bca;
  wire v3773bc6;
  wire v374673a;
  wire v3739f29;
  wire v3a700d8;
  wire v23fdf1a;
  wire v3a70786;
  wire v3a5c57a;
  wire v3a6988c;
  wire v376296b;
  wire v373824d;
  wire v37730ab;
  wire v3a67c9e;
  wire v372e4e3;
  wire v3741be8;
  wire v3a70ce7;
  wire v3734c40;
  wire v373aa96;
  wire v37568c9;
  wire v3a70005;
  wire v3a6cc28;
  wire v3727b18;
  wire v3a681ed;
  wire v373c897;
  wire v377ba8e;
  wire v3a704bf;
  wire v3768a78;
  wire v3778f46;
  wire v3a70499;
  wire v37665f9;
  wire v37441dc;
  wire v3a6aba6;
  wire v3a70287;
  wire v3769c51;
  wire v3745196;
  wire v37691ab;
  wire v3a6f11b;
  wire v3735b5a;
  wire v3755cf7;
  wire v377a8dc;
  wire v3727a10;
  wire v3778b2a;
  wire v3a6762b;
  wire v372ebbf;
  wire v3a70aeb;
  wire d3068c;
  wire v377479e;
  wire v3760e2e;
  wire v3763f48;
  wire v3a6600a;
  wire v3768b99;
  wire v3748ae2;
  wire bd3213;
  wire v3740f70;
  wire v375208a;
  wire v374c6e1;
  wire v3751161;
  wire v3a5f0a7;
  wire v3a6fdf8;
  wire v3a6b710;
  wire v3757b55;
  wire v3a64190;
  wire v377a3bd;
  wire v3a5faba;
  wire v3a6e089;
  wire v3a672e5;
  wire v3a6fbe6;
  wire v3766d1b;
  wire v3727cd0;
  wire v1e37b65;
  wire v373ef30;
  wire v3a6ceb7;
  wire v3a5810a;
  wire v35b7160;
  wire v377bc89;
  wire v376c635;
  wire v373f8b1;
  wire v377b4f7;
  wire v3a70f04;
  wire v3a64b41;
  wire v377e2f7;
  wire v3a6f322;
  wire v3737dad;
  wire v374a08a;
  wire v375ceee;
  wire v3a6a57c;
  wire v374bd1f;
  wire v375a338;
  wire v373946b;
  wire v3a5b615;
  wire v3a7127d;
  wire v3a6b078;
  wire v3729e0b;
  wire v3a70b37;
  wire v3a6f7a1;
  wire v372bf35;
  wire v38094e9;
  wire v374bc10;
  wire v374f860;
  wire v372fbf8;
  wire v375d38f;
  wire v37390ba;
  wire v1e37a69;
  wire v3a6feb9;
  wire v372d5bb;
  wire v3760b17;
  wire v3766996;
  wire v3768933;
  wire v372e88a;
  wire v38095b2;
  wire v3a6ec56;
  wire v3772541;
  wire v3a56b60;
  wire v373d9a2;
  wire v3778419;
  wire v37786f9;
  wire v376b5c0;
  wire v3767cd6;
  wire v37493b9;
  wire v374a8df;
  wire v3a70ac0;
  wire v3a6f102;
  wire v3a6eb5a;
  wire v3a6f4f4;
  wire v3a5c210;
  wire v3758824;
  wire v3a6f0d3;
  wire v3a5b826;
  wire v3a70b7c;
  wire v372ff0a;
  wire v374f432;
  wire v3735c5d;
  wire v3a5927f;
  wire v372b22b;
  wire v3a70e07;
  wire v3730afc;
  wire v3a6f0a9;
  wire v3761fc1;
  wire v3769cd6;
  wire v3764ca8;
  wire v3a6bdd1;
  wire v3774a1e;
  wire v3a7057a;
  wire v375d3cd;
  wire v374ebb6;
  wire v376021d;
  wire v3773d96;
  wire v3809464;
  wire v3a66529;
  wire v376550d;
  wire v3766597;
  wire v3770919;
  wire v3a6fa49;
  wire v3725d7b;
  wire v377e904;
  wire v3a5df33;
  wire v3a61fd3;
  wire v3762be8;
  wire v3807026;
  wire v2925d2c;
  wire v3a6f9d9;
  wire v373561e;
  wire v3757996;
  wire v3a539c3;
  wire v375f97d;
  wire v3a70a5f;
  wire v3752ed7;
  wire v376a799;
  wire v375636e;
  wire v3a6fc19;
  wire v3a6afdd;
  wire v3740bce;
  wire v373703c;
  wire v374ef20;
  wire v372a55a;
  wire v3a5a868;
  wire v37591e8;
  wire v37657e4;
  wire v3a585b7;
  wire v372d75a;
  wire v3779678;
  wire v37429a7;
  wire v3724ab6;
  wire v374df45;
  wire v375fcb7;
  wire v377c94b;
  wire v3731749;
  wire v3733862;
  wire v3a69ae7;
  wire v373530a;
  wire v3a63f3d;
  wire v373e6f1;
  wire v39ebb74;
  wire v3a66999;
  wire v3743bbe;
  wire v373a33d;
  wire v373c8cb;
  wire v3a7049a;
  wire v377f2ea;
  wire v3754237;
  wire v3744cfe;
  wire v3a5b42a;
  wire v3773e09;
  wire v37234e0;
  wire v375e1a2;
  wire v3777692;
  wire v37578b4;
  wire v375cb72;
  wire v3a5b286;
  wire v375c674;
  wire v3a7165d;
  wire v3779e1b;
  wire v373fdfb;
  wire v3770538;
  wire v3a6f6bd;
  wire v3725b75;
  wire v374378e;
  wire v3a70bb8;
  wire v3734abe;
  wire v3a65eba;
  wire v3a6a233;
  wire v23fda6a;
  wire v373dbb0;
  wire v37777d2;
  wire v3a70524;
  wire v3a61298;
  wire v373261a;
  wire v373577f;
  wire v3a65cfb;
  wire v3738b0c;
  wire v3743eda;
  wire v3a56898;
  wire v37718de;
  wire v3756930;
  wire v37364cf;
  wire v3a5950d;
  wire v3a704dc;
  wire v3731de2;
  wire v3a6ff30;
  wire v376a7b2;
  wire v377ba09;
  wire v376daec;
  wire v3729c7e;
  wire v380911c;
  wire v373c23e;
  wire v3742140;
  wire v3a6c7fe;
  wire v37455c2;
  wire v377c5c2;
  wire v3a6c33a;
  wire v372cd45;
  wire v3772ab1;
  wire v3752201;
  wire v37265f6;
  wire v37299fa;
  wire v37684cf;
  wire v3733d5a;
  wire v377005e;
  wire v373374d;
  wire v37436cf;
  wire v372f3f1;
  wire v3a70fdb;
  wire v3a7045e;
  wire v3a70fed;
  wire v3a70fcf;
  wire v3a5b567;
  wire v3a6db03;
  wire v3738aa2;
  wire v374b7ea;
  wire v374ac78;
  wire v37323c5;
  wire v375c62d;
  wire v3a6f6af;
  wire v372bd06;
  wire v372da2f;
  wire v3a6d2eb;
  wire v372fb53;
  wire v39ebb5d;
  wire v37447f7;
  wire v373d1bb;
  wire v3a7035f;
  wire v376f505;
  wire v3a69bbf;
  wire cbb40b;
  wire v3774d12;
  wire v3772ee4;
  wire a6f1de;
  wire v37370b9;
  wire v3a6bdca;
  wire v3724fe8;
  wire v374c425;
  wire v377a511;
  wire v3752222;
  wire v3a711b9;
  wire v3a6ff26;
  wire v3a60723;
  wire v3775ad3;
  wire v375c65a;
  wire v372bc6c;
  wire v2619ad7;
  wire v377a345;
  wire v37275cf;
  wire v3a6b80e;
  wire v3a5faaa;
  wire v376791c;
  wire v37573b9;
  wire v3a713ee;
  wire v3a71219;
  wire v3741020;
  wire v372ecd8;
  wire v37369f2;
  wire v3a71474;
  wire v3a705a8;
  wire v374dd8f;
  wire v37600da;
  wire v3753837;
  wire v380854b;
  wire v3a6b908;
  wire v37471e0;
  wire v3762d3e;
  wire v376d3d1;
  wire v3754f54;
  wire v3730b77;
  wire v373dbc5;
  wire v3a5919f;
  wire v3a70d8a;
  wire v23fd96e;
  wire v376c4a9;
  wire v3a70d85;
  wire v376189d;
  wire v3742a57;
  wire v3759a08;
  wire v37660d9;
  wire v373e284;
  wire v377bf2b;
  wire v3a5d704;
  wire v37611c1;
  wire v3a6e9b8;
  wire v3a66123;
  wire v3a684bb;
  wire v376894a;
  wire v3a6f9a4;
  wire v2619aa7;
  wire v3a70aa3;
  wire v3775729;
  wire v372ead5;
  wire v3749a1d;
  wire v3752b6a;
  wire v372b893;
  wire v8955d0;
  wire v3778091;
  wire v3a65e17;
  wire v3a68b7d;
  wire v3a5a37a;
  wire v3a64fce;
  wire v373127a;
  wire v3765406;
  wire v3a58c95;
  wire v37702e8;
  wire v3a5cf84;
  wire v3a705c0;
  wire v3a6ff06;
  wire v37472b6;
  wire v3735468;
  wire v3751c73;
  wire v3729381;
  wire v375f777;
  wire v3a606d2;
  wire v375ea88;
  wire v3752ebb;
  wire v3a54e0c;
  wire v3746976;
  wire v3733739;
  wire v3a7017b;
  wire v3a68467;
  wire v3a705ea;
  wire v37434eb;
  wire v374a9e4;
  wire v377b732;
  wire v373478e;
  wire v373c1e4;
  wire v374adfa;
  wire v3734c59;
  wire v3809e77;
  wire v375035f;
  wire v37268b6;
  wire v3a701f3;
  wire v377c923;
  wire v37315c8;
  wire v3a29850;
  wire v3a6a5a8;
  wire v3a65f7a;
  wire v3756918;
  wire v3a6fd5e;
  wire v3a71276;
  wire v2ff9229;
  wire v376ea80;
  wire v3743477;
  wire v37392d7;
  wire v375b344;
  wire v2889709;
  wire v3738944;
  wire v3a6f4d5;
  wire v374650b;
  wire v3a68228;
  wire v3777340;
  wire v3a6f5ec;
  wire v372633a;
  wire v372abf1;
  wire v37641ad;
  wire v380a1f3;
  wire v37686ea;
  wire v3a5bf4c;
  wire v3a70f06;
  wire v376740b;
  wire v376bb7b;
  wire v376e0df;
  wire v39ebb64;
  wire v376afdf;
  wire v3742c9b;
  wire v3a70bf8;
  wire v3744081;
  wire v3742b79;
  wire v3738da4;
  wire v377b3d5;
  wire v3a661cd;
  wire v37c03ff;
  wire v37754ac;
  wire v375d758;
  wire v23fdea8;
  wire v3774618;
  wire v3a6f882;
  wire v3728c46;
  wire v373447d;
  wire v3808cee;
  wire v3762c44;
  wire v376ae9c;
  wire v3731cf0;
  wire v3a6bf04;
  wire v374a454;
  wire v3764628;
  wire v374f31c;
  wire v3a7042c;
  wire v3a60a24;
  wire v37523dd;
  wire v3729516;
  wire v376a847;
  wire v3723d1a;
  wire v3a5ef2e;
  wire v37253a5;
  wire v377946d;
  wire v39a4eaa;
  wire v37625a7;
  wire v3a57c47;
  wire v3a669dc;
  wire v3a537c5;
  wire v376f24b;
  wire v3a5b3f9;
  wire v3a6fd1c;
  wire v3a5b78f;
  wire v39eb418;
  wire v372e3db;
  wire v372ad29;
  wire v3a678f9;
  wire v3a6dada;
  wire v3a5e394;
  wire v3a56a52;
  wire v3a5ada2;
  wire v3a6ac81;
  wire v37734ba;
  wire v3772add;
  wire v1e37d82;
  wire v3a57db6;
  wire v2acadfb;
  wire v377957e;
  wire v3763b6c;
  wire v375a64f;
  wire v3a5cdf4;
  wire v3a70360;
  wire v375f046;
  wire v3a5ba6d;
  wire b1ca9b;
  wire v3748caf;
  wire v3757343;
  wire v374c73d;
  wire v375c861;
  wire v374828c;
  wire v3a70a64;
  wire v3a6241d;
  wire v372b1dc;
  wire v3a70c4d;
  wire v37379bb;
  wire v37471f0;
  wire v3a71230;
  wire v3a71119;
  wire v37652b1;
  wire v3736ebd;
  wire v37b6451;
  wire v3a6cb69;
  wire v9da9d2;
  wire v3a703de;
  wire v3722fc0;
  wire v3a5db5f;
  wire v3a710bb;
  wire v372e611;
  wire v373b719;
  wire v3771c59;
  wire v37638de;
  wire v37430f5;
  wire v3739681;
  wire v3a71391;
  wire d1bf3b;
  wire v3a641ea;
  wire v373d029;
  wire v3763ca1;
  wire v37742f4;
  wire v37430db;
  wire v372d1b1;
  wire v3a6f671;
  wire v375b16e;
  wire v3768be2;
  wire v3739ca5;
  wire v3732c24;
  wire v37448f2;
  wire v3a7007b;
  wire v373f2a6;
  wire v3747d5a;
  wire v3753638;
  wire v3730818;
  wire v3774c3f;
  wire v3758e3c;
  wire v3a70823;
  wire v373b5f0;
  wire v3740b82;
  wire v375896e;
  wire v39a4f17;
  wire c9bec3;
  wire v37431b5;
  wire v3762a9c;
  wire v374fbca;
  wire v374f29f;
  wire v375da09;
  wire v3735354;
  wire v3a6fa0d;
  wire v37740f9;
  wire v3a650bb;
  wire v374b1a4;
  wire v3775f56;
  wire v3749c2f;
  wire v3a5fc70;
  wire v376fc80;
  wire v37656c1;
  wire v3729e17;
  wire v375d7df;
  wire v374949d;
  wire v374deab;
  wire v377cf71;
  wire v372b59f;
  wire v3a70a48;
  wire v3740890;
  wire v372e712;
  wire v3a6f56b;
  wire v377e3fe;
  wire v3a6178e;
  wire v3724947;
  wire v377681e;
  wire v373bd8b;
  wire v3747fbc;
  wire v3772bff;
  wire v3807723;
  wire v375c041;
  wire v3726a78;
  wire v377ea73;
  wire v3a5f4b2;
  wire v372df9a;
  wire v37332dd;
  wire v376cf62;
  wire v373ac15;
  wire v3a6ef4e;
  wire v3767cc0;
  wire v3a71398;
  wire v3a5f60f;
  wire v373c164;
  wire v3a57913;
  wire v376fe7d;
  wire b1f79b;
  wire v3a6f657;
  wire v375eef1;
  wire v376f860;
  wire v3743256;
  wire v372825b;
  wire v374d648;
  wire v37567db;
  wire v377b9fd;
  wire v3a6dca6;
  wire v3a5921b;
  wire v3746289;
  wire b00c46;
  wire v3726cd4;
  wire a5f27e;
  wire v374b88a;
  wire v3762f14;
  wire v377d6c5;
  wire v3a6c063;
  wire v3a70d67;
  wire v3a715b0;
  wire v37758d0;
  wire v374f44c;
  wire v3778e46;
  wire b62018;
  wire v23fd8b2;
  wire v3a70a21;
  wire v374cf68;
  wire v3768522;
  wire v373fb32;
  wire v373cb13;
  wire v3a57887;
  wire v3a5a711;
  wire v37537cc;
  wire v3770e43;
  wire v3a5bff1;
  wire v372463a;
  wire v39372da;
  wire v377815d;
  wire v3731f07;
  wire v3377c79;
  wire v373b16f;
  wire v377f3ae;
  wire v37302a2;
  wire v3a6fb00;
  wire v37308bc;
  wire v373a2b4;
  wire v37706ef;
  wire v3a6cd87;
  wire v3736a59;
  wire v373e13a;
  wire v3a6fcb2;
  wire v375be9f;
  wire v372402f;
  wire v35b6c3a;
  wire v3a704ef;
  wire v3807a7d;
  wire v8455c7;
  wire v3a70c77;
  wire v3725c13;
  wire v375e813;
  wire v3a70e09;
  wire c587b2;
  wire v373deb5;
  wire v3a6ffca;
  wire v377989c;
  wire v3a6392b;
  wire v3a6589b;
  wire v3769093;
  wire v3745529;
  wire v37541f4;
  wire v37325a2;
  wire v374d138;
  wire v375f41f;
  wire v3774bed;
  wire v3a7043e;
  wire v372e367;
  wire v3a6a8ee;
  wire v3a716a6;
  wire v373f2e2;
  wire v3a70ff5;
  wire v3a70369;
  wire v3a5dafb;
  wire v375e958;
  wire v3732c56;
  wire v374db8d;
  wire v8455c3;
  wire v376363f;
  wire v3a70ba1;
  wire v375f938;
  wire v373ad95;
  wire v373ab12;
  wire v377230a;
  wire v373f349;
  wire v2acb0d7;
  wire v3a6dae0;
  wire v373c275;
  wire v9af7ec;
  wire v376402f;
  wire v3749cea;
  wire v3379037;
  wire v3a6d4c2;
  wire v372e305;
  wire v372b304;
  wire v374eb89;
  wire v3733df1;
  wire v37721df;
  wire c39398;
  wire v374da61;
  wire v3a71486;
  wire v372e263;
  wire v3763c09;
  wire v3a6fdbc;
  wire v374c679;
  wire v3a70796;
  wire v377ab6b;
  wire v375ccf3;
  wire v3a64058;
  wire v3774bad;
  wire v3a6f270;
  wire v3a6fbf8;
  wire v3779680;
  wire v3752428;
  wire v39eb4ca;
  wire v3a6499e;
  wire v3a569b7;
  wire v3a60b2e;
  wire v37297e8;
  wire v373dd5a;
  wire v3767cc9;
  wire v3a5c983;
  wire v372c85e;
  wire v2acb068;
  wire v3766a64;
  wire v3724d8c;
  wire v3a6fa0a;
  wire v37786c6;
  wire v3762892;
  wire v3a5f21c;
  wire v380760a;
  wire v375a510;
  wire v377981b;
  wire v3769c72;
  wire v3a57e01;
  wire v372c49f;
  wire v3769af4;
  wire v3778ca0;
  wire v374bb64;
  wire v3777b18;
  wire v3a6dea6;
  wire v3a61100;
  wire v37665bf;
  wire v374caab;
  wire v372640f;
  wire v3776e9c;
  wire d5f283;
  wire v37548c4;
  wire v37556fd;
  wire v3a58924;
  wire v377416d;
  wire v37668e9;
  wire v373e209;
  wire v37454a8;
  wire v3a6a07b;
  wire v372edf6;
  wire b0e59c;
  wire v3749f94;
  wire v373a841;
  wire v3a6a129;
  wire v3a64dc2;
  wire v373de4b;
  wire v37433f5;
  wire v3765436;
  wire v3a607af;
  wire v3744fc9;
  wire v3a6ef34;
  wire v377db81;
  wire v35b71da;
  wire v373c22e;
  wire v3a5468d;
  wire v37748b7;
  wire v3a70a5c;
  wire v37635ab;
  wire v3a70f4d;
  wire v3773dc6;
  wire v3773afc;
  wire v3a63f29;
  wire v3a714ab;
  wire v3a6fb21;
  wire v373741d;
  wire v373399e;
  wire v3a6f0f9;
  wire v3740aa7;
  wire v3a70530;
  wire v37422b5;
  wire v377af44;
  wire v3a6f520;
  wire v3747666;
  wire v3a6546b;
  wire v3765e46;
  wire v3729f25;
  wire v3741748;
  wire v37700ee;
  wire v373aaa8;
  wire v372fd0a;
  wire v37720f9;
  wire v377d7dc;
  wire v3748fe0;
  wire v3749004;
  wire v37542d8;
  wire v375c009;
  wire v3a5ab24;
  wire c08050;
  wire v37538af;
  wire v375c94e;
  wire v3a56197;
  wire v3768502;
  wire v3a6ff35;
  wire v376f017;
  wire v377d671;
  wire v376fb92;
  wire v374f645;
  wire v373f262;
  wire v374d54c;
  wire v374e52d;
  wire v375d887;
  wire v3771758;
  wire v3a5fd4a;
  wire v3a67862;
  wire v3a5d5a4;
  wire v37332af;
  wire v3a296dc;
  wire v3a67dd5;
  wire v375649e;
  wire v3a71291;
  wire v3722ac4;
  wire v3a6b78f;
  wire v3749283;
  wire v37645c9;
  wire v373bac2;
  wire v37480b3;
  wire v374e4c0;
  wire v377308e;
  wire v3771394;
  wire v372d8f9;
  wire v3744ef1;
  wire v3a6ad44;
  wire v3730ddd;
  wire v372343e;
  wire v3a71228;
  wire d4d3bb;
  wire v3a6ef2c;
  wire v3a5ab08;
  wire v37747a9;
  wire v372346b;
  wire v3737d90;
  wire v3728ee0;
  wire v372fb2a;
  wire v37c0294;
  wire v3a55a75;
  wire v3a5c41b;
  wire v372f5ca;
  wire v3762e85;
  wire v3a711e6;
  wire v372af06;
  wire v373b837;
  wire v3771e26;
  wire v377f3ba;
  wire v3751b6b;
  wire v377a2d1;
  wire v3747db9;
  wire v37317ba;
  wire v375d304;
  wire v377c7c0;
  wire v376d955;
  wire v373aed4;
  wire v37625f2;
  wire v3768064;
  wire v3a57be6;
  wire ab638b;
  wire v377b774;
  wire v374d184;
  wire v373389a;
  wire v3774524;
  wire v377b4bf;
  wire v375adcd;
  wire v8c5d6a;
  wire v373014d;
  wire v8455bf;
  wire v3a55392;
  wire v3a656ca;
  wire v3777479;
  wire v374b25d;
  wire v374d4ae;
  wire v3a6fd1b;
  wire v3774608;
  wire v375a2ac;
  wire v3a5d1c9;
  wire v3760ab8;
  wire v377caa3;
  wire v372c60a;
  wire v3a5b121;
  wire v372d8e2;
  wire v374b077;
  wire v3a67462;
  wire v3a70db3;
  wire v3761df7;
  wire v37307a7;
  wire v3a5732f;
  wire v375e1de;
  wire v3a5af68;
  wire v3a695f1;
  wire v3a57e1a;
  wire v3a5689e;
  wire v3752000;
  wire v3a710c1;
  wire v377d107;
  wire v35b7168;
  wire v375fa8b;
  wire v377efdc;
  wire v3773982;
  wire v3723542;
  wire v37280b0;
  wire v2acb056;
  wire v3a70e5a;
  wire v3755820;
  wire v3a69dc1;
  wire v374c95a;
  wire v375a94a;
  wire v3776914;
  wire v3a54ebe;
  wire v3a68084;
  wire v3a7029e;
  wire v9e8d30;
  wire v3756ea2;
  wire v3760c3d;
  wire v3a63daa;
  wire v3a707c5;
  wire v377f80c;
  wire v376b7ff;
  wire v375c1d1;
  wire v3a6da8a;
  wire v2092abe;
  wire v3742cd4;
  wire v3762100;
  wire a5c619;
  wire v376bc98;
  wire v3747e71;
  wire v37266b1;
  wire v3766f7d;
  wire v3725198;
  wire v37797a3;
  wire v3a710c6;
  wire v3808f73;
  wire v3762969;
  wire v3732511;
  wire v377419d;
  wire v3736ded;
  wire v3a6b423;
  wire v23fe0be;
  wire v3a57e6d;
  wire v3a61f46;
  wire v3a5857c;
  wire v3774655;
  wire v3a5b289;
  wire v8455bb;
  wire v3728e89;
  wire v3a6f674;
  wire v372f23a;
  wire v3a70e4f;
  wire v377ed5e;
  wire v3743e7b;
  wire v376d85d;
  wire v372f05b;
  wire v375efe0;
  wire v3767561;
  wire v3a71288;
  wire v373cdba;
  wire v373adf1;
  wire v3a6cf15;
  wire v2619b43;
  wire v376b15b;
  wire v3a701a1;
  wire v87be38;
  wire v3729700;
  wire v373f836;
  wire v3744835;
  wire v372adb6;
  wire v3722fc5;
  wire v375dc75;
  wire v374d07a;
  wire v37443ab;
  wire v3727084;
  wire v3760513;
  wire v3770ecc;
  wire v3a70490;
  wire v375a159;
  wire v3a6338d;
  wire v374915c;
  wire v3a713f2;
  wire v3a71284;
  wire v37471cb;
  wire v3724e8e;
  wire v3a707b7;
  wire v372a00b;
  wire v37412f3;
  wire v373c15d;
  wire v3740349;
  wire v375fcfb;
  wire v3a5f0b2;
  wire v3a70f08;
  wire v3a6e13d;
  wire v3a6b9e8;
  wire v3748665;
  wire v3732b75;
  wire v377a083;
  wire v372b60b;
  wire v3751069;
  wire v3750b86;
  wire v374b747;
  wire v373763f;
  wire v376b438;
  wire v3a55e3c;
  wire v373bb3a;
  wire v3763a20;
  wire v373127e;
  wire v3a6fb2b;
  wire v377bbf7;
  wire v37251f1;
  wire v3a6f8f5;
  wire v375d92e;
  wire v3a5bc2c;
  wire v3a6f9c3;
  wire v376730a;
  wire v373f940;
  wire v3776633;
  wire v3a6f012;
  wire v3735bbc;
  wire v374680c;
  wire v3a6aa15;
  wire v3773940;
  wire v3a62c0a;
  wire v3743b12;
  wire v3774641;
  wire v377f883;
  wire cfaa3a;
  wire v374fe49;
  wire v35b773b;
  wire v3764bee;
  wire v373dee7;
  wire v377cd7a;
  wire v374c163;
  wire v3a55bd0;
  wire v3766a8d;
  wire v3725770;
  wire v3a6fc2f;
  wire v374355f;
  wire v3749149;
  wire v3a6c9ab;
  wire v3766b48;
  wire v3a6f53a;
  wire v375977c;
  wire v3a714f6;
  wire v3731487;
  wire v374df14;
  wire v375c334;
  wire v375bb92;
  wire v35b77ec;
  wire v3768b46;
  wire v3a62a96;
  wire v3a68967;
  wire v3759c49;
  wire v377a434;
  wire v3a6f3a2;
  wire v3a5d590;
  wire v37418db;
  wire v3a67d4f;
  wire v3a625b1;
  wire v377bcb3;
  wire v377e442;
  wire cb8cbb;
  wire v3807029;
  wire v3764c4a;
  wire v37465d7;
  wire v9c492b;
  wire v3a6f3ab;
  wire v37716c3;
  wire v3779627;
  wire v373c631;
  wire v37314f2;
  wire v377169f;
  wire v126f91f;
  wire v373d67c;
  wire v3724e64;
  wire v3a704f3;
  wire v3729c6b;
  wire v3732415;
  wire v375fbba;
  wire v372310e;
  wire v375eb97;
  wire v3a6d642;
  wire v28896da;
  wire v3741320;
  wire v373adaa;
  wire v3724e45;
  wire v374f533;
  wire v3a557a1;
  wire v37690fe;
  wire v3a70a2b;
  wire v377854f;
  wire v3806a1c;
  wire v3a7131f;
  wire v3a7084e;
  wire v377bf37;
  wire v3a65da7;
  wire v3760f64;
  wire v37296f5;
  wire v3a5e7fe;
  wire v3756a9e;
  wire bbeeaf;
  wire v3750dd3;
  wire v374eaf4;
  wire v37267f3;
  wire v3a66c66;
  wire v3742275;
  wire v377e406;
  wire v3a5e388;
  wire v3a7007c;
  wire v3a6f031;
  wire v3a6fcea;
  wire v2ff9371;
  wire v3753ee8;
  wire v3808db4;
  wire v3755b07;
  wire v3774937;
  wire v37436e6;
  wire v372dbe7;
  wire v3a57540;
  wire v3762cdf;
  wire v37338d8;
  wire v377e1f6;
  wire v375ed6f;
  wire v3732564;
  wire v3a5c6f9;
  wire v3a6eb2f;
  wire v3742035;
  wire v377fc4b;
  wire v377f584;
  wire v3a56002;
  wire v3a62cb7;
  wire v3778a2f;
  wire v325b591;
  wire v377af09;
  wire v3a6f99c;
  wire v376d0bc;
  wire v3a70364;
  wire v3777009;
  wire v3a5f984;
  wire v380777f;
  wire v3754d88;
  wire v374a41b;
  wire v372d3b2;
  wire v3a5a48f;
  wire v3738e6e;
  wire v3728738;
  wire v3776b22;
  wire v373340f;
  wire v3770ffb;
  wire v3a70c78;
  wire v3750f3b;
  wire v3a6f886;
  wire v3a6c73d;
  wire v372aeef;
  wire v37734cb;
  wire v37539c8;
  wire v377f501;
  wire v3748251;
  wire v3a6fc28;
  wire v372ef56;
  wire v35b70ed;
  wire v3765aa0;
  wire v3a5c1e7;
  wire v377ecec;
  wire v3750b01;
  wire v374d59d;
  wire v3735b64;
  wire v375fe2b;
  wire v3737bd8;
  wire v3a71439;
  wire v3742b92;
  wire v3765248;
  wire v2acb015;
  wire v3a2a422;
  wire v3722b6c;
  wire v3725325;
  wire v3a69631;
  wire v3a70c81;
  wire v3777ac3;
  wire v3769edd;
  wire v3a70f45;
  wire v375671a;
  wire v3727bd4;
  wire v3a5fa29;
  wire v373c0b4;
  wire v3723fa6;
  wire v374e61c;
  wire v3764099;
  wire db32f1;
  wire v3a59cf3;
  wire v3a6e975;
  wire v3a704fe;
  wire v37596f3;
  wire v37244b9;
  wire v3a704e1;
  wire v374bfd6;
  wire v3755774;
  wire v3743094;
  wire v376924d;
  wire v3a5f08f;
  wire v3a668e4;
  wire v3808914;
  wire v3a7078d;
  wire v3a6f114;
  wire v3763c97;
  wire v376fa50;
  wire v3a6f98e;
  wire v372f03c;
  wire v3a70622;
  wire v375a92d;
  wire v3a6f451;
  wire v374193d;
  wire v3a6f9d3;
  wire v3755c3f;
  wire v3a6862e;
  wire v3766607;
  wire v3722af7;
  wire v3a6c555;
  wire v373293c;
  wire v3732e45;
  wire v3a69a42;
  wire v3729b75;
  wire v3a61cb0;
  wire v3a708c9;
  wire v3739c6f;
  wire v3a70c67;
  wire v23fde9c;
  wire v3a5c75c;
  wire v3a5bbaa;
  wire v376f37e;
  wire v3a6667c;
  wire v1e3737f;
  wire v376e0cb;
  wire v372ff96;
  wire v3a6fe76;
  wire v3729a69;
  wire v37263c1;
  wire v87762a;
  wire v373eeec;
  wire v3734810;
  wire v374b2c2;
  wire v37676a5;
  wire v3726bcc;
  wire v377bd17;
  wire v375a76e;
  wire v3a6427b;
  wire v3773ce0;
  wire v372d925;
  wire v3a6d695;
  wire v37257e5;
  wire v3a6fcf1;
  wire v23fdd8d;
  wire v376293f;
  wire v3a656b2;
  wire v37309ae;
  wire v2925cef;
  wire v37445e6;
  wire v3736c86;
  wire v37659e4;
  wire a7b390;
  wire v3a6fb4a;
  wire v37385e9;
  wire v3a296d3;
  wire v376fa86;
  wire v3a6f15d;
  wire v373f394;
  wire v3a63e68;
  wire v3776be5;
  wire v3807072;
  wire v3a70bec;
  wire v374801c;
  wire v3724c8c;
  wire v375fc56;
  wire v3a60030;
  wire v8cf677;
  wire v373ee81;
  wire v3a5cfb0;
  wire v3745dae;
  wire v3766645;
  wire v373f780;
  wire v3743b49;
  wire v372a8d9;
  wire v3747b2b;
  wire v3a70b77;
  wire v3767415;
  wire v376ef2d;
  wire v3a62236;
  wire v3a6f317;
  wire v3a7010c;
  wire v37659c6;
  wire v377632d;
  wire v3a67a02;
  wire v3730bae;
  wire v377984a;
  wire v372d891;
  wire v3757e15;
  wire v3757f07;
  wire v3731159;
  wire v3736e7c;
  wire v3a698d8;
  wire v372d33c;
  wire v3a70a79;
  wire v3a60691;
  wire v3726f6b;
  wire aa9893;
  wire v3a6fc77;
  wire v3a70b5b;
  wire v3a6edf6;
  wire v3a70080;
  wire v373a1d0;
  wire v372588c;
  wire v3a703ba;
  wire v3a7075d;
  wire v3a54519;
  wire v3a6ef60;
  wire v3759519;
  wire v39a53e9;
  wire v3a69057;
  wire v23fe20d;
  wire v3727bc6;
  wire v3728464;
  wire v374cb02;
  wire v375fe7a;
  wire v3746ae3;
  wire v3a5a954;
  wire v3a6cc5f;
  wire v3a70655;
  wire v375930e;
  wire v3724e4b;
  wire v374f6a4;
  wire v3a7013d;
  wire v3732da2;
  wire v3757993;
  wire v374c837;
  wire v9bd777;
  wire v375bc49;
  wire v3749520;
  wire v3a6f6c8;
  wire v374dd11;
  wire v3a70eb8;
  wire v3766f8a;
  wire v3766ef7;
  wire v374e78f;
  wire v372b0ac;
  wire v3749ece;
  wire v374f1a1;
  wire v375f52b;
  wire v372e751;
  wire v3761f22;
  wire v377c34f;
  wire v372d727;
  wire v3729eb0;
  wire v3a633c5;
  wire v3a640c5;
  wire v3757fcc;
  wire v373a2f2;
  wire v373e814;
  wire v3763b0a;
  wire v3776ada;
  wire v1e3737d;
  wire v3a6b266;
  wire v376d680;
  wire v374edba;
  wire v3a6bee8;
  wire v3a70f93;
  wire v3729798;
  wire v1e3778c;
  wire v37341fd;
  wire v3a70c8f;
  wire v3748c75;
  wire v3a5cd20;
  wire v375018e;
  wire v373125c;
  wire v3759abe;
  wire v374e26d;
  wire v3a5cbd8;
  wire v377aa06;
  wire v373141b;
  wire v3a70c3e;
  wire v374a97f;
  wire v3763acf;
  wire v37607e8;
  wire v3737534;
  wire v376b57e;
  wire v372d967;
  wire v3757a57;
  wire v37368e1;
  wire v374b887;
  wire v3a5fc48;
  wire v37430f0;
  wire v376fdbe;
  wire v376f9d3;
  wire v8c9ea7;
  wire v375cebd;
  wire v3a70a22;
  wire v3a5dad5;
  wire v373de86;
  wire v3765463;
  wire v3738a59;
  wire v373664d;
  wire v375609e;
  wire v3808994;
  wire v377a60f;
  wire v373cf66;
  wire v3737f5a;
  wire v376289b;
  wire v3a7125f;
  wire v37387ed;
  wire v3777996;
  wire v373e654;
  wire v374df0b;
  wire v374bf8a;
  wire v3a706b1;
  wire v3a5a824;
  wire v373e642;
  wire v376a2ea;
  wire v3774911;
  wire v3a6f10f;
  wire v37467f3;
  wire v3773016;
  wire v374c062;
  wire v3a71208;
  wire v3758f3c;
  wire v1e37e76;
  wire v3a5b539;
  wire v37737c9;
  wire v3739dae;
  wire v3a6ff87;
  wire v3778648;
  wire v3741216;
  wire v3a6d74f;
  wire v374b47b;
  wire v3752577;
  wire v3733e0a;
  wire v375c41e;
  wire v3739ea3;
  wire v3747ad5;
  wire v375eee3;
  wire v3a5864f;
  wire v374c78e;
  wire v372ba66;
  wire v376e7e8;
  wire v375d00a;
  wire v377fabb;
  wire b68bf2;
  wire v3a71374;
  wire v372b12d;
  wire v3a297f5;
  wire v3757dea;
  wire v987445;
  wire v3756012;
  wire v3a6eb21;
  wire v37316f2;
  wire v37308fc;
  wire v374f754;
  wire v37601d6;
  wire v376bc6a;
  wire v3a5a63c;
  wire v373f91b;
  wire v3a708fa;
  wire v3730e2e;
  wire v3a6f986;
  wire v3773e2a;
  wire v3a615f7;
  wire v374c01f;
  wire v3a70edc;
  wire v372a837;
  wire v374721d;
  wire v3728760;
  wire v3723aea;
  wire v3730ca3;
  wire v373905f;
  wire v3a71682;
  wire v3809a76;
  wire v3a704c9;
  wire v3772c12;
  wire v376c863;
  wire v37748b2;
  wire v37299b3;
  wire v376c235;
  wire v3a5aee5;
  wire v375ec98;
  wire v360d147;
  wire v3a702e8;
  wire v373330f;
  wire v3730e90;
  wire v3730b98;
  wire v3a6c03d;
  wire v373a7ab;
  wire v3a7015e;
  wire v37343d1;
  wire v37501e1;
  wire v3a6fac9;
  wire v376cd02;
  wire v3a5c8c9;
  wire v3a56c1f;
  wire v37265c1;
  wire v37365c6;
  wire v37359cf;
  wire v3772083;
  wire v372ed55;
  wire v372f151;
  wire v3a6e3e0;
  wire v3a71195;
  wire v3730c3c;
  wire v3766222;
  wire v3a6f318;
  wire v3746e94;
  wire v39ebb31;
  wire v372451b;
  wire v3a5d4d0;
  wire v3a6b73c;
  wire v3767a85;
  wire v3a6c09f;
  wire v39ea0c2;
  wire v3a598da;
  wire v3a7140b;
  wire v3743c84;
  wire v3a64612;
  wire v37610ae;
  wire v372eb90;
  wire v3757b39;
  wire v3769559;
  wire v374c0d0;
  wire v3730b8c;
  wire v3809e3c;
  wire v372d827;
  wire v3a6d2e2;
  wire v3743df6;
  wire v374a2b5;
  wire v3a66cee;
  wire v3a7017a;
  wire v3762fc4;
  wire v3a5f308;
  wire v376430b;
  wire v374bb56;
  wire v376442b;
  wire v3a6cdbc;
  wire v377613d;
  wire v3a57ad0;
  wire v3a62550;
  wire v3a603fc;
  wire v3737bb4;
  wire v376dcd0;
  wire v3a69248;
  wire v377e56f;
  wire v3a706b7;
  wire v3a6fac6;
  wire v3752cc5;
  wire v37467a6;
  wire v376f5ef;
  wire v373681a;
  wire v3a5e363;
  wire v3722a7e;
  wire v3734634;
  wire v3761bee;
  wire v3758bfe;
  wire v3a67996;
  wire v3749ab1;
  wire v377ab2c;
  wire v3736a9a;
  wire v3a70315;
  wire v373f2b6;
  wire v3a70967;
  wire v3808870;
  wire v3a70848;
  wire v376a4dd;
  wire v8e4749;
  wire v3769945;
  wire v373222d;
  wire dcb1a9;
  wire v372834d;
  wire v373fa3d;
  wire v1e377bd;
  wire v3a55e7d;
  wire v37345f5;
  wire v375e309;
  wire v37509c7;
  wire v3a6ef74;
  wire a69e17;
  wire v37395f5;
  wire v3a68ef7;
  wire v377574b;
  wire v37531b1;
  wire v3a6f856;
  wire v375e400;
  wire v3a62c12;
  wire v372faf1;
  wire v3734465;
  wire v3779582;
  wire v3760854;
  wire v3a70829;
  wire v3a6f8dc;
  wire v375c771;
  wire v360d080;
  wire v372c706;
  wire v373b8e2;
  wire v2619b04;
  wire v376d1cb;
  wire v3a6f03d;
  wire v372a22d;
  wire v3a71097;
  wire v3a6d569;
  wire v3a6f641;
  wire v3729f41;
  wire v3a5d644;
  wire v3772409;
  wire v2acaeaa;
  wire v3a7169d;
  wire v372690e;
  wire v37289bb;
  wire v3a6fcef;
  wire v37655ac;
  wire v3a5ee12;
  wire v3768d47;
  wire v3a60258;
  wire v37703a5;
  wire v3a7119c;
  wire v377c2d9;
  wire v37474e8;
  wire v1e3732b;
  wire v3757440;
  wire v3a6b4a6;
  wire v3a714f2;
  wire v3739849;
  wire v3a6ebf2;
  wire v3766f14;
  wire v3728f25;
  wire v3777817;
  wire v35ba1cf;
  wire v3777853;
  wire v20930c6;
  wire v3a705bc;
  wire v3767f7f;
  wire v3a6fd0a;
  wire v3809388;
  wire v37685bf;
  wire v3768c2e;
  wire v3a70eb7;
  wire v3745b51;
  wire v3a712ae;
  wire v1e37c22;
  wire v3749e4b;
  wire v372438e;
  wire v3751dd2;
  wire v3751631;
  wire v3a6fd0c;
  wire v23fe37e;
  wire v37370f0;
  wire v3a5fd58;
  wire v372cd37;
  wire v3773340;
  wire v3755539;
  wire v3729382;
  wire v372b33d;
  wire v3778aac;
  wire v3a69714;
  wire v3779070;
  wire v3740161;
  wire v3a55173;
  wire v37645a4;
  wire v3768d3e;
  wire v3771b2c;
  wire v372c503;
  wire v372b790;
  wire v3750269;
  wire v3a299c1;
  wire v376bd2a;
  wire v3777ff3;
  wire v3772e90;
  wire v1e3746e;
  wire v377a2e4;
  wire v373aecf;
  wire v376a4c0;
  wire v2093059;
  wire v3a710bc;
  wire v3741850;
  wire v3a71548;
  wire v375ac48;
  wire v375f8b0;
  wire v3743824;
  wire v372ad53;
  wire v375fbc0;
  wire v37306d8;
  wire v3775165;
  wire v3a575d6;
  wire v3748964;
  wire v37534a4;
  wire v3a6c437;
  wire v3a70a2a;
  wire v3a59833;
  wire v3a7051c;
  wire v373d3dd;
  wire v376ff89;
  wire v37784cc;
  wire v3727347;
  wire v373d7f9;
  wire v3733e62;
  wire v3a5c30f;
  wire v3723477;
  wire v3a710fc;
  wire v3731fc6;
  wire v3a57ed1;
  wire v37331af;
  wire v3a62348;
  wire v375c718;
  wire v3a68e5d;
  wire a708cc;
  wire v3a699a1;
  wire v372bfa1;
  wire v3a664ba;
  wire v373325b;
  wire v373b1cb;
  wire v377e24d;
  wire v376d41b;
  wire v37272df;
  wire v3776715;
  wire v3a5b359;
  wire v372c83f;
  wire v3743546;
  wire v377f21b;
  wire v3734af6;
  wire v372c4c6;
  wire v3a5e7a5;
  wire v3761865;
  wire v3a6305e;
  wire v377b086;
  wire v3a69062;
  wire v3a6124f;
  wire v3a70645;
  wire v3a70e8d;
  wire v377657c;
  wire v373b36c;
  wire v3750c9f;
  wire v3a53329;
  wire v3a5fd34;
  wire v3a705db;
  wire v37581c2;
  wire v3a660b5;
  wire v3743c22;
  wire v3778921;
  wire v3763d79;
  wire v376f409;
  wire v3a66615;
  wire v3776917;
  wire v3a6f1e6;
  wire v373a291;
  wire v3760a2c;
  wire v37733f9;
  wire v3a65aca;
  wire v374f501;
  wire v2acb5c7;
  wire v3a7020b;
  wire v376e3db;
  wire v3754421;
  wire v3a58b8f;
  wire v3767b88;
  wire v375f452;
  wire v373580a;
  wire v373a588;
  wire v3777342;
  wire v3a58907;
  wire v3754a4d;
  wire v37572c1;
  wire v372d51c;
  wire v37411ab;
  wire v3a562b7;
  wire v3754c86;
  wire v3a6480b;
  wire v3a70b2c;
  wire v37414b0;
  wire v37735a0;
  wire v3769cff;
  wire v3a70dc4;
  wire v3a6c355;
  wire v3a6e47f;
  wire v3a68aa8;
  wire v1e3791d;
  wire v373cf4e;
  wire v3743252;
  wire b4fa3c;
  wire v3a6f646;
  wire v3a70e9a;
  wire v37353c0;
  wire v372b4ba;
  wire v374a45c;
  wire v3731258;
  wire v3743745;
  wire v3a5db66;
  wire v3763498;
  wire v39eaa47;
  wire v37359d8;
  wire v376bad8;
  wire v372bf87;
  wire v3755bc2;
  wire v377e14d;
  wire v3a712de;
  wire v3a6006c;
  wire v374815b;
  wire v87cef3;
  wire v377da37;
  wire v376352a;
  wire v3a59351;
  wire v3a70cea;
  wire v3a58a8e;
  wire v3a6b5bc;
  wire v373f954;
  wire abddc4;
  wire v372e562;
  wire v3a6fc96;
  wire v3a7106c;
  wire v377b59e;
  wire v3a70d79;
  wire v376660c;
  wire v373c96e;
  wire v37304b3;
  wire v3725092;
  wire v3a6a831;
  wire v3a709df;
  wire v3732aca;
  wire v375c8e8;
  wire v3739018;
  wire v3a5f20c;
  wire v3733090;
  wire v3a66737;
  wire v3770e2b;
  wire v375a0ff;
  wire v3765b88;
  wire v3749529;
  wire v373b7c8;
  wire v377b68c;
  wire v3a69d81;
  wire v37360b3;
  wire v3734b15;
  wire v3722f16;
  wire v375db62;
  wire v373abdb;
  wire v375bff8;
  wire v3a66d0e;
  wire v3729cfe;
  wire v3724026;
  wire v377682d;
  wire v37794fa;
  wire v3777417;
  wire v377c723;
  wire v3745131;
  wire v375179a;
  wire v374052a;
  wire v39ebab4;
  wire v373262e;
  wire v376954d;
  wire v3753b80;
  wire v3a701fa;
  wire v3a64f2d;
  wire d039bc;
  wire v373a891;
  wire v3a6677e;
  wire v3a70308;
  wire v3727ad4;
  wire v3736e19;
  wire v3778e71;
  wire v376489a;
  wire v37554d5;
  wire v374304d;
  wire v37558e4;
  wire v3a70fa6;
  wire v3a7094f;
  wire v3a6513d;
  wire v3a63831;
  wire v3732701;
  wire v3806db0;
  wire v3a5fee0;
  wire c52384;
  wire v3727f3b;
  wire v37554cd;
  wire v3a5bb4e;
  wire bfae74;
  wire v3a712cc;
  wire v3a685ee;
  wire v3728962;
  wire cd743d;
  wire v3a708d6;
  wire v3a6e844;
  wire v99b721;
  wire v3a5f869;
  wire v3762617;
  wire v3760617;
  wire v3a70b62;
  wire v3a5a4c0;
  wire v374bd23;
  wire v3760bfa;
  wire v3753994;
  wire v37570eb;
  wire v3a6afcd;
  wire v3a5e747;
  wire v3771882;
  wire v372e959;
  wire v37363ae;
  wire v375ba66;
  wire v372e74c;
  wire v372b57a;
  wire v37683bf;
  wire v376592b;
  wire v3a6e721;
  wire v3a5fa45;
  wire v376faf0;
  wire v375c24b;
  wire v3a70f8c;
  wire v3a70298;
  wire v37571c5;
  wire v3a711bd;
  wire v3774161;
  wire v37682d5;
  wire v3773015;
  wire v373a3c3;
  wire v3732849;
  wire v374d218;
  wire v37439b2;
  wire v372fa70;
  wire v377b0f7;
  wire v375cd5d;
  wire v3a7089d;
  wire v372e889;
  wire v3749540;
  wire v3a5ec50;
  wire v3a6fdf7;
  wire v37677d8;
  wire v3a6f7a0;
  wire v3729620;
  wire v3752ac9;
  wire v374877e;
  wire v374586a;
  wire v96dd76;
  wire v3a6eefb;
  wire v3738adf;
  wire v3a5fe2f;
  wire v3725149;
  wire v372ce98;
  wire v3a59609;
  wire v3758c41;
  wire v3731511;
  wire v3a6fc74;
  wire v374e7e6;
  wire ce4abb;
  wire v3757d75;
  wire v375a637;
  wire v3a54c9b;
  wire v3729b4c;
  wire v3771715;
  wire v3a70c91;
  wire v3a6c7e8;
  wire v376e5de;
  wire v375ac26;
  wire v3740546;
  wire v3a711ed;
  wire v3a5ff4b;
  wire v376b3d0;
  wire v3755d20;
  wire v3a67257;
  wire v3a70371;
  wire v376ba62;
  wire v3a6f45a;
  wire v3779e95;
  wire v3778c61;
  wire v3756809;
  wire v3745ce4;
  wire v3754b03;
  wire v3a6fc3f;
  wire v3776fb2;
  wire v3a6f1e7;
  wire v3a6f187;
  wire v2925d06;
  wire v3750f27;
  wire v3a6ec22;
  wire v3a6540f;
  wire v3a60131;
  wire v3a71072;
  wire v375af0b;
  wire v3727581;
  wire v3778619;
  wire v88e7d1;
  wire v3727f9c;
  wire v376a236;
  wire v376d287;
  wire v1e37561;
  wire v3a70877;
  wire v3a62ba4;
  wire v374294f;
  wire v3a56929;
  wire v374803b;
  wire v377bbfc;
  wire v3762aaf;
  wire v376e966;
  wire v39eb033;
  wire v3764a8a;
  wire v3a70642;
  wire v37536b2;
  wire v3736ef2;
  wire v3777d63;
  wire v3770a5b;
  wire v376360a;
  wire v37377d2;
  wire v3a6f07b;
  wire v375b02a;
  wire v3763104;
  wire v3775a4a;
  wire v375c05f;
  wire v3a6f585;
  wire v3725091;
  wire v3a56e79;
  wire v3748e0b;
  wire v3762498;
  wire v3a6fbe4;
  wire v37399b4;
  wire v3a6f147;
  wire v3a5795e;
  wire v3a646f5;
  wire v3745aff;
  wire v2acaf74;
  wire v37720d8;
  wire v375cdb1;
  wire v37316b7;
  wire v3a7145f;
  wire v39a52e6;
  wire v3a70020;
  wire v3760073;
  wire v3723d55;
  wire v3772117;
  wire v3770dcb;
  wire v372ee41;
  wire v3774075;
  wire v372de68;
  wire v3a7143f;
  wire v38099ce;
  wire v37708e7;
  wire v3a6f746;
  wire v3a6e0f4;
  wire v3a70c8c;
  wire v3777f05;
  wire v3746351;
  wire v376f175;
  wire v376b141;
  wire v8c4a86;
  wire v37482be;
  wire v376897b;
  wire v3760279;
  wire v337897a;
  wire v3a6fd11;
  wire v3769041;
  wire v37c0190;
  wire v373a29c;
  wire v374a407;
  wire v3746683;
  wire v37593a1;
  wire v376aaef;
  wire v372d035;
  wire v372c09a;
  wire v3a5eb63;
  wire v375588a;
  wire v3756beb;
  wire v373274f;
  wire v373afd5;
  wire v3a6ff28;
  wire v37538ff;
  wire c7d127;
  wire v37621e9;
  wire v3a5e63b;
  wire v37349ce;
  wire v3a70cf0;
  wire v375e00a;
  wire v3a69f9e;
  wire v3a5a76b;
  wire v3773aa0;
  wire v37431eb;
  wire v3a5b12c;
  wire v373ecae;
  wire v374b0a8;
  wire v3724121;
  wire v376278c;
  wire v3a5988f;
  wire v3766b27;
  wire v3727ec9;
  wire v3a54344;
  wire v372f292;
  wire v3a62986;
  wire v372d1bf;
  wire v3768a57;
  wire v3a68d49;
  wire v3a66387;
  wire v374e1dc;
  wire v3745871;
  wire v3a6a8aa;
  wire v377ce96;
  wire v3770b6e;
  wire v3a5f67d;
  wire v375590f;
  wire v3735afb;
  wire v3a6ff4e;
  wire v3a62bd5;
  wire v3769a71;
  wire v37283c8;
  wire v37638ef;
  wire v375b03c;
  wire v376a87f;
  wire v375e64c;
  wire v3a602a4;
  wire v377a901;
  wire v3730926;
  wire v3755e35;
  wire v3a680b9;
  wire v3a6fa30;
  wire v374fa56;
  wire v374fcf6;
  wire v3a6b688;
  wire v37c038c;
  wire v3a6ff37;
  wire v3a56866;
  wire v3730b62;
  wire v377e52f;
  wire v3a70889;
  wire v374421d;
  wire v374e246;
  wire v3a70349;
  wire v3a6face;
  wire v3759007;
  wire v3a71231;
  wire v374f630;
  wire a6859a;
  wire v375a0ec;
  wire v375c917;
  wire v3771fbb;
  wire v3769c47;
  wire v3a706f6;
  wire v375ac16;
  wire v97ea11;
  wire v3731e16;
  wire v3768b80;
  wire v373683d;
  wire v3723299;
  wire v1e37cab;
  wire v3772362;
  wire v3a6f947;
  wire v374068b;
  wire v3a6f884;
  wire v376c747;
  wire v3757182;
  wire v3731e60;
  wire v3a6065f;
  wire v3764de7;
  wire v373d932;
  wire v3779e66;
  wire v3766d0d;
  wire v3a5cf22;
  wire a89e0c;
  wire v377bf9f;
  wire v360be60;
  wire v3a702cc;
  wire v37590d1;
  wire v3770fef;
  wire v3749dc1;
  wire v376af8d;
  wire v2aca81d;
  wire v372d237;
  wire v3723e00;
  wire v376e822;
  wire v3a6f932;
  wire v3a64361;
  wire v3a6f117;
  wire v375a51f;
  wire v37492d2;
  wire v377bf21;
  wire v377eab5;
  wire v376c31d;
  wire v3a63368;
  wire v3763311;
  wire v3a6fb7b;
  wire v38097c4;
  wire v3a57dbb;
  wire v3a6e031;
  wire v3378fc3;
  wire v3a6eb22;
  wire v3a6fbda;
  wire v375e50c;
  wire v377dfa2;
  wire v3a6fc73;
  wire v3a5e38d;
  wire v3775cca;
  wire v373edb9;
  wire v376fd7a;
  wire v3a63a66;
  wire v376e033;
  wire v33781d5;
  wire v3a5690d;
  wire v3726c5b;
  wire v373c965;
  wire v376c6ed;
  wire v3776b9a;
  wire v3a64045;
  wire v375a99b;
  wire v3a669ae;
  wire v3a6c688;
  wire v3a683a4;
  wire v37558b4;
  wire v377293c;
  wire v3745993;
  wire v3a5fc3c;
  wire v3a715e1;
  wire v3a637ca;
  wire v3a70566;
  wire v373109c;
  wire v3a708c3;
  wire v3a5af82;
  wire v3a652a6;
  wire v3a7159c;
  wire v3a6f647;
  wire v3a66ade;
  wire v3778c64;
  wire v375cc1b;
  wire v3a6f8f6;
  wire v3746e4e;
  wire v3a58dac;
  wire v373cdb0;
  wire a90ef2;
  wire v375647e;
  wire v3a5a2be;
  wire v3749760;
  wire v3a5e55e;
  wire v37c048c;
  wire v3773e17;
  wire v3a6073f;
  wire v377de56;
  wire v373f9eb;
  wire v372b316;
  wire v3756b5c;
  wire v3a70932;
  wire c98bc3;
  wire v37467e9;
  wire v3a6fe0e;
  wire v3a70725;
  wire v2092f41;
  wire v377ec59;
  wire v376b83d;
  wire v377803a;
  wire v37597a4;
  wire v3a57fff;
  wire v3a57c48;
  wire v372bf93;
  wire v3776ca8;
  wire v3747ec5;
  wire v3a6fb8c;
  wire v3a6bc47;
  wire v3a6ffe5;
  wire v3724392;
  wire v37461e1;
  wire v3754229;
  wire v372ac3b;
  wire v3732e59;
  wire v3a71667;
  wire v3a70cf4;
  wire v375b597;
  wire v372b009;
  wire v3773ff0;
  wire v3a6573d;
  wire v376d9c6;
  wire v3764ee3;
  wire v3744898;
  wire v373ef10;
  wire v3a5604a;
  wire v3a6f7b9;
  wire v373dc42;
  wire v3770717;
  wire v376ab51;
  wire v3776e5b;
  wire v3771f9b;
  wire v3a6f2d4;
  wire v2889705;
  wire v3a6be6d;
  wire v3a5fb37;
  wire v3723dae;
  wire v3a6fe58;
  wire v373e2db;
  wire v37627bf;
  wire v3a5a057;
  wire v373f8a7;
  wire v37364d2;
  wire v37329ec;
  wire v3a708e2;
  wire v374e29a;
  wire v375a579;
  wire v3a6546f;
  wire v3a5c50b;
  wire v3a5417e;
  wire v3a7074d;
  wire v3771994;
  wire v37723ce;
  wire v375e21e;
  wire v3a701ec;
  wire v375199a;
  wire v37679d9;
  wire v3a6fe35;
  wire v374d749;
  wire v373cc5c;
  wire v37265d6;
  wire v37311de;
  wire v3757637;
  wire v3a67b28;
  wire v37278c2;
  wire v3757fde;
  wire v3767b98;
  wire v3a70c63;
  wire v3a5fc8d;
  wire v3a6f874;
  wire v374449e;
  wire v37789ca;
  wire v3745aae;
  wire v3a61b59;
  wire v3a7105f;
  wire v376cf96;
  wire v3a63930;
  wire v3758c5e;
  wire v373c00f;
  wire v372bdc2;
  wire v3a67c8e;
  wire v3743b66;
  wire v37626a9;
  wire v3a62f70;
  wire ae4185;
  wire v3771fea;
  wire v37437bb;
  wire v3a5c2f5;
  wire d62ab4;
  wire v372bb5d;
  wire v377734d;
  wire v37701a5;
  wire v3a70d69;
  wire v3733d4f;
  wire v3a6a1e8;
  wire v3a61202;
  wire v3a6f469;
  wire v3a5fc61;
  wire v3a667ba;
  wire v37450aa;
  wire v3763f38;
  wire v3748990;
  wire v3a67899;
  wire v376faf6;
  wire v3a709d3;
  wire v3736e12;
  wire v3762557;
  wire v3747006;
  wire v374723b;
  wire v3776bc7;
  wire v3a6ffce;
  wire v3744ada;
  wire v37701a0;
  wire v376e532;
  wire v3a5f69c;
  wire v37378e5;
  wire v37319cd;
  wire v2092aba;
  wire v3a62f0b;
  wire v3a67729;
  wire v37306cd;
  wire v376305b;
  wire v3a6fe94;
  wire v3742ec4;
  wire v37637d5;
  wire v3a6f3a1;
  wire v380719b;
  wire v3a6f3c4;
  wire v37341b2;
  wire v377222a;
  wire v3a64722;
  wire v372d435;
  wire v3a6ff74;
  wire v375b26a;
  wire v3778352;
  wire v2ff87b0;
  wire v3a5a2e4;
  wire v3764ac0;
  wire v374c0c9;
  wire v3a6f3aa;
  wire v3a6fcfe;
  wire v375f4c8;
  wire v3752d10;
  wire v37237be;
  wire bd3d3d;
  wire v3761c68;
  wire v3a710b7;
  wire v3a702b4;
  wire cd3a92;
  wire v3770a77;
  wire v374ff44;
  wire v374ca41;
  wire v3763004;
  wire v372ea14;
  wire v3750d4c;
  wire v380988c;
  wire v3776492;
  wire v3a665ab;
  wire v3743338;
  wire v3776faf;
  wire v375b2d9;
  wire v373574c;
  wire v3a553db;
  wire v3a6e1ed;
  wire v37656b8;
  wire v37315c5;
  wire v3a70a70;
  wire v3760509;
  wire v3a64c71;
  wire v3743efa;
  wire v3a70c51;
  wire v377f5cb;
  wire v3a6d5e9;
  wire v376aa10;
  wire v3a5f162;
  wire v37496d3;
  wire v3a636d9;
  wire v3a533d3;
  wire v3a2a8f2;
  wire v373fcf4;
  wire v3a713c7;
  wire v3a70e02;
  wire v3a59bb4;
  wire v3742ef6;
  wire v3a70bd0;
  wire v3766572;
  wire v3775c0a;
  wire v377d3e4;
  wire v3743f94;
  wire v373abbe;
  wire v3a6f6fa;
  wire v377abb1;
  wire v373d551;
  wire v374aca8;
  wire v3735134;
  wire v3a70ca7;
  wire v3a70f67;
  wire v3a65503;
  wire v360cfe2;
  wire v3737c13;
  wire v3a6cedc;
  wire v39a4e8f;
  wire v374bec6;
  wire v376c5f5;
  wire v3a712fd;
  wire v37350f9;
  wire v3a70bf6;
  wire v375a938;
  wire v3a70759;
  wire v3754b79;
  wire v375ccc3;
  wire v3749cf7;
  wire v373ecd8;
  wire v372d3ea;
  wire v373f488;
  wire v3775f1f;
  wire v3723614;
  wire v3733fad;
  wire v3806f70;
  wire v1e37d8b;
  wire v8f64f2;
  wire v375a0b3;
  wire v3a5c5b5;
  wire v3750c38;
  wire v373c1d7;
  wire v3740fef;
  wire v3744983;
  wire v3808ed4;
  wire v3776a5c;
  wire v3a6b691;
  wire v373f6c9;
  wire v3749b46;
  wire v3774710;
  wire v3a551d6;
  wire v3a70418;
  wire v376441d;
  wire v3772f4d;
  wire v3a7162e;
  wire v376005f;
  wire v3a5a397;
  wire v3a711e0;
  wire v3777666;
  wire v374b9f9;
  wire v37285a1;
  wire v372b765;
  wire v3a703a4;
  wire v37325ad;
  wire v377cdea;
  wire v3a71660;
  wire v3758187;
  wire v3754d3a;
  wire v3a708e7;
  wire v3730057;
  wire v3a6f505;
  wire v37273d2;
  wire v3728179;
  wire v37622f5;
  wire v33781df;
  wire v28896e3;
  wire v374220d;
  wire v3741357;
  wire v376de5c;
  wire v3a70ee6;
  wire v3a6df5a;
  wire v375baed;
  wire v3728498;
  wire v380954b;
  wire v3a70e69;
  wire v3741384;
  wire v3741c91;
  wire v3759efd;
  wire v377a352;
  wire v3a7088b;
  wire v3a6f237;
  wire v3750113;
  wire v3728ae9;
  wire v3a6eace;
  wire v3a62fc6;
  wire v1e37a06;
  wire v3a5e9e9;
  wire v3a6f78f;
  wire v3761ca6;
  wire v39eb519;
  wire v397fb7c;
  wire v373f537;
  wire v3749a46;
  wire v3756087;
  wire v3a711c6;
  wire v3727a16;
  wire v3730fab;
  wire v3a64eba;
  wire v37364a3;
  wire v376301d;
  wire v377b26a;
  wire v3a68787;
  wire v37784b3;
  wire v3a60b0f;
  wire v376a1c9;
  wire v3a5ff7c;
  wire v372d378;
  wire v3774bc0;
  wire v3a70482;
  wire v3751aab;
  wire v3750d4d;
  wire a9e394;
  wire v377bc8e;
  wire v3a6efc0;
  wire v376964a;
  wire v3769a1c;
  wire v38075cd;
  wire v373580d;
  wire v375495e;
  wire v3a5f891;
  wire v37787dd;
  wire v3a6eb8c;
  wire v3a596c4;
  wire v3a708e3;
  wire v3728ced;
  wire v3a70000;
  wire v373446a;
  wire v3a54b46;
  wire v375babe;
  wire v3a6f5a0;
  wire v37510a5;
  wire v3a5507a;
  wire v37725e7;
  wire v38072fb;
  wire v3a71319;
  wire v375fe5b;
  wire v3a66e4c;
  wire v37235f9;
  wire v3a65368;
  wire v3a5a211;
  wire v372ba45;
  wire v372a823;
  wire v3768c5d;
  wire v3729a2a;
  wire v375a345;
  wire v374e849;
  wire v375492b;
  wire v37658d7;
  wire v3a5a76d;
  wire v37543d8;
  wire v37725f6;
  wire v375185f;
  wire v376073d;
  wire v2092ac0;
  wire v3a5edcb;
  wire v37571f1;
  wire v3a70986;
  wire v37425ad;
  wire v3a70dde;
  wire v1e38288;
  wire v376d935;
  wire v376f661;
  wire v3750b9e;
  wire v3a61482;
  wire v3a6180b;
  wire v37712f8;
  wire v3756f17;
  wire v377960b;
  wire v3a6ee64;
  wire v1e37cd7;
  wire v3725649;
  wire v3762c26;
  wire v376614b;
  wire v3750eb8;
  wire v3a7139f;
  wire v3a6f8a0;
  wire v1e377ba;
  wire aa421e;
  wire v37643e5;
  wire v3806b78;
  wire v3a54350;
  wire v3a582d8;
  wire v372fe8b;
  wire v375626c;
  wire v376d060;
  wire v3766ff3;
  wire v2092a7a;
  wire v3a6ef73;
  wire v374ac72;
  wire v37693a9;
  wire d78807;
  wire v37532ac;
  wire v3a70c5d;
  wire v3723501;
  wire v3735ed2;
  wire v373e28c;
  wire v37400ba;
  wire v37766f3;
  wire v374d92c;
  wire v3731172;
  wire v37c039c;
  wire v376d6f9;
  wire v3a6cfe0;
  wire v3769806;
  wire v377dcbc;
  wire v3738fba;
  wire v372c151;
  wire v373b42b;
  wire v373a101;
  wire v3a56518;
  wire v3729e05;
  wire v372d48d;
  wire v89c52e;
  wire v3743702;
  wire v37467da;
  wire v3a7042a;
  wire v3806e7b;
  wire v3755a84;
  wire v375b65b;
  wire v37491b7;
  wire v3765d2a;
  wire v373cde8;
  wire v375f53a;
  wire v376b4a7;
  wire v3a576d3;
  wire v37507f4;
  wire v3a6d622;
  wire v3777da5;
  wire v373b748;
  wire v3a70210;
  wire v3806798;
  wire v376983e;
  wire v3753eb3;
  wire v375dcac;
  wire v3a70509;
  wire v3a6eb95;
  wire v37715af;
  wire v3764486;
  wire v3a6f386;
  wire v3751d98;
  wire v373a803;
  wire v373b317;
  wire v3725ccb;
  wire v3737ad2;
  wire d0a27e;
  wire v3a6fd95;
  wire v372422d;
  wire v3a57484;
  wire v3762223;
  wire v3742eaf;
  wire v8ad83a;
  wire v3a6f571;
  wire v3a5a5d1;
  wire v3731a5a;
  wire v372c480;
  wire v3743dbc;
  wire v3a70c01;
  wire v37441e0;
  wire v3759605;
  wire v37376c1;
  wire v3735112;
  wire v3a55584;
  wire v373ec98;
  wire v37551b9;
  wire v3a611bd;
  wire v372f202;
  wire v376bf10;
  wire v3750c47;
  wire v3a53c21;
  wire v375314d;
  wire v3a613cc;
  wire v3a71028;
  wire v3728e58;
  wire v37391ac;
  wire v3759d08;
  wire v372c2bf;
  wire v3a705a9;
  wire v3a702e7;
  wire v37607a7;
  wire v374dad0;
  wire v3738ea9;
  wire v37775dd;
  wire v3a6a64a;
  wire v3758291;
  wire v374c3bf;
  wire v3746fdb;
  wire v377296d;
  wire v372aacf;
  wire v37354a9;
  wire v37257e9;
  wire v3744fb6;
  wire v373b91e;
  wire v372f11d;
  wire v374c7e6;
  wire v375dc43;
  wire v3a71448;
  wire v375b24f;
  wire v23fda6c;
  wire v37255e9;
  wire v377609a;
  wire v3a6f7ef;
  wire v3739b5c;
  wire v37731ec;
  wire v374e401;
  wire v3a6fa3c;
  wire v3a70696;
  wire v3a70922;
  wire v3a6fd3f;
  wire v375b5ce;
  wire v37719a9;
  wire v37676cd;
  wire v3a6d7cd;
  wire v373df82;
  wire v37553b9;
  wire v3a6fb1b;
  wire v3728203;
  wire v3754086;
  wire v3a701c4;
  wire v3a62f60;
  wire v37293d5;
  wire v375f74e;
  wire v3a5d2d3;
  wire v3760707;
  wire v3756b39;
  wire v3773d39;
  wire v3743cd6;
  wire v3731aeb;
  wire v3a70e65;
  wire v3754260;
  wire v3a69e8c;
  wire v37778e2;
  wire v3779fb2;
  wire v3779227;
  wire v3765351;
  wire v376bb27;
  wire v3a6ff1a;
  wire v374b15d;
  wire v375444a;
  wire v3a659e5;
  wire v3a6fc43;
  wire v32562a3;
  wire v3748146;
  wire v377015c;
  wire v37547ad;
  wire v3a5641a;
  wire v377c07a;
  wire v374ec91;
  wire v3766924;
  wire v3730217;
  wire v376a9de;
  wire v375b143;
  wire v37662e2;
  wire v37276f2;
  wire v373f410;
  wire v37420bb;
  wire v3a6ef47;
  wire v3751d16;
  wire v37fca8d;
  wire v372cbdb;
  wire v3742241;
  wire v377e60e;
  wire v375cfd7;
  wire v377652b;
  wire v374510e;
  wire v3a70621;
  wire v374fd8d;
  wire v3724a1c;
  wire v373b10f;
  wire v3a70966;
  wire v377814b;
  wire v377773f;
  wire v376a95c;
  wire v2889716;
  wire v377e512;
  wire v374d970;
  wire v3a6152c;
  wire v37610e5;
  wire v3a6fa84;
  wire v3a6c1ac;
  wire v3a6f99d;
  wire v3a6fc30;
  wire v372acab;
  wire v3a65aeb;
  wire v9bbda1;
  wire v3729dfc;
  wire v37511a1;
  wire v376fbe0;
  wire v3a61c49;
  wire v3729ed7;
  wire v3739ba9;
  wire v3751e76;
  wire v37485c0;
  wire v3a70a0e;
  wire v3738f5a;
  wire v3768633;
  wire v3a55844;
  wire v3a70cd3;
  wire v3a6c390;
  wire v372cdc9;
  wire v37282f3;
  wire v373c97a;
  wire v377ef7c;
  wire v3757656;
  wire v3a66ef6;
  wire v374a7ab;
  wire v3778281;
  wire v3763d20;
  wire v3759584;
  wire v3a6f45c;
  wire v377d047;
  wire v377c003;
  wire v3736db8;
  wire v376df24;
  wire v375ced2;
  wire v37460cd;
  wire v3733fd0;
  wire v373c437;
  wire v377a4e5;
  wire v376c17d;
  wire v3378f4e;
  wire v3732736;
  wire v3769a60;
  wire v3a5d015;
  wire v37300d7;
  wire v373924d;
  wire v374ab4b;
  wire v917443;
  wire v3776d32;
  wire v37546a4;
  wire v3a6f2ee;
  wire v37523c6;
  wire v3723ef8;
  wire v3a702c0;
  wire v37454c6;
  wire v3a7144d;
  wire v3770ea8;
  wire v37d8c61;
  wire v3736041;
  wire v375446f;
  wire v377ee33;
  wire v372300f;
  wire v377f180;
  wire v325b59f;
  wire v360d0fd;
  wire v23fdf1b;
  wire v3a707a4;
  wire v3a705fc;
  wire v3a715ca;
  wire v3a602c3;
  wire v374b73b;
  wire v3761fb5;
  wire v375b713;
  wire v373ae91;
  wire v377a478;
  wire v3a70353;
  wire v37272a8;
  wire v376baef;
  wire v376993b;
  wire v3a5de18;
  wire v3a588a0;
  wire v3772a3f;
  wire v3a57118;
  wire v375bd8c;
  wire v3a6bf63;
  wire v372dc51;
  wire v3a67fd9;
  wire v3734cb7;
  wire v3a6ccd6;
  wire v3760fab;
  wire v372afda;
  wire v3a69ad3;
  wire v37480ec;
  wire v3745658;
  wire v373dfec;
  wire v372e05a;
  wire v3a70866;
  wire v375f0af;
  wire db3b98;
  wire v37735cb;
  wire v37734f8;
  wire v33782e5;
  wire v3a702d3;
  wire v375ac50;
  wire v37690af;
  wire v377bfb6;
  wire v3a59df2;
  wire v3a70e9b;
  wire v3728957;
  wire v374700b;
  wire v38090ee;
  wire v37728dc;
  wire v376c335;
  wire v377273d;
  wire v376e605;
  wire v3a5cc9d;
  wire v3a714e9;
  wire v3a68822;
  wire v3a5bc04;
  wire v377b038;
  wire v3a6a54d;
  wire v373144a;
  wire v374a3b7;
  wire v3a704ea;
  wire v373f17f;
  wire v3a5cd88;
  wire v3a70240;
  wire v3739062;
  wire v374a84c;
  wire v3a64417;
  wire v3a6f2cf;
  wire v3725f02;
  wire v3a705ce;
  wire v3a603cf;
  wire v3758418;
  wire v35b724d;
  wire v3774653;
  wire v37615ce;
  wire v3727a2f;
  wire v372d8f7;
  wire v3a6fc83;
  wire v3a6fef1;
  wire v3a715ac;
  wire cbd026;
  wire v37521f6;
  wire v376fdb9;
  wire v3747a53;
  wire v3a6f7fb;
  wire v3a6fc60;
  wire v3734778;
  wire v3774791;
  wire v3732b12;
  wire v3a5b583;
  wire v374a2be;
  wire v3755f9a;
  wire v37297af;
  wire v3a611e6;
  wire v3a6b575;
  wire v377376d;
  wire v3a6fc38;
  wire v3809f5f;
  wire v3735f7a;
  wire v375de2d;
  wire v373dd27;
  wire v3744792;
  wire v376e17a;
  wire v3736b71;
  wire v3a6f164;
  wire v3738844;
  wire v374d695;
  wire v376c1c3;
  wire v3723df0;
  wire v377f37e;
  wire v3a69ef8;
  wire v376c27d;
  wire v3a6fb03;
  wire v372d748;
  wire v375b9a3;
  wire v3772374;
  wire v3a6fe83;
  wire v37371be;
  wire v376fff8;
  wire v23fe152;
  wire v3733b84;
  wire v37334ff;
  wire v3a70d72;
  wire v3760251;
  wire v37683f8;
  wire v3740a9c;
  wire v3a6fc95;
  wire v3734ef4;
  wire v3723023;
  wire v377098c;
  wire v37325e0;
  wire v3a70fd9;
  wire v3727195;
  wire v3736003;
  wire v3a66fb0;
  wire v3725ca4;
  wire v3a6dc57;
  wire v377a337;
  wire v373f1d4;
  wire v3a70f4a;
  wire v375a412;
  wire v3755cc3;
  wire v3735ae4;
  wire v3a63f6d;
  wire v3a70176;
  wire v373178d;
  wire v375a4c4;
  wire v372d772;
  wire v3a71484;
  wire v3732772;
  wire v3a70b3c;
  wire v3a572d0;
  wire v373af6f;
  wire v372efc8;
  wire v3a70b61;
  wire v373bbce;
  wire v3770c0d;
  wire v3809386;
  wire v3722dd6;
  wire v3764a58;
  wire c827f4;
  wire v3a6faf6;
  wire v374e855;
  wire v37414ed;
  wire v3a69eb7;
  wire v3763295;
  wire v1e37b5a;
  wire v3756a59;
  wire v1e37368;
  wire v37284f8;
  wire v3724543;
  wire v3a5c640;
  wire v882147;
  wire v3758a7c;
  wire v3a70e37;
  wire v37261b2;
  wire v8455cb;
  wire v375654b;
  wire v3726838;
  wire v3a6c2a9;
  wire v3a71133;
  wire v3a6e675;
  wire v3773040;
  wire v37559d6;
  wire v375f1db;
  wire v372efb1;
  wire v375f78f;
  wire v375cab5;
  wire v3a70407;
  wire v3724c55;
  wire v3a6be79;
  wire v374478f;
  wire v3a62ad0;
  wire v3a5f648;
  wire v3a70e72;
  wire v375e8c1;
  wire v3a6f470;
  wire v375e21d;
  wire v3749e68;
  wire v3727fa7;
  wire v3a65909;
  wire v374ecd5;
  wire v3a69606;
  wire v37647e3;
  wire v3747243;
  wire v3768551;
  wire v3a61ff9;
  wire v3765f8e;
  wire v37790bd;
  wire v3a6f681;
  wire v3a5520d;
  wire v33789f3;
  wire v3762cf7;
  wire v3a698b7;
  wire v373b6e9;
  wire v376147a;
  wire v3a59cde;
  wire v1e37c6e;
  wire v3777e7d;
  wire v3a609da;
  wire v372e684;
  wire v3a6fe0c;
  wire v3807765;
  wire v3a709fc;
  wire v3744399;
  wire v375830c;
  wire v3a71305;
  wire v3744ad5;
  wire v3a6f86f;
  wire v3723fb3;
  wire v3a6519c;
  wire v3768e48;
  wire v3a68426;
  wire v3a71014;
  wire v3725410;
  wire v373e2f9;
  wire v372311c;
  wire v3a645c2;
  wire v375fa82;
  wire v372ab21;
  wire v3a5a17f;
  wire v3a6b4a2;
  wire v3722f60;
  wire v3771820;
  wire v8455b7;
  wire v377f0fb;
  wire v374e61f;
  wire v3732302;
  wire v374d479;
  wire v3756b48;
  wire v37759b6;
  wire v372433d;
  wire v23fe156;
  wire v3a6393d;
  wire v374eb9c;
  wire v3737554;
  wire v3a70d71;
  wire v37453d8;
  wire v3753418;
  wire v375d9f8;
  wire v3a705f2;
  wire v3a70909;
  wire v376c014;
  wire v1e37acb;
  wire v3773ee6;
  wire v3767b70;
  wire v3a56eb1;
  wire v3a67de3;
  wire v3766dcc;
  wire v3769adb;
  wire v373c404;
  wire v3a6165e;
  wire v380974c;
  wire v3a6eb98;
  wire v37640ff;
  wire v3a6c2d2;
  wire v3768202;
  wire v3a6f533;
  wire v3a7054c;
  wire v3777312;
  wire v3725367;
  wire v3a705d3;
  wire v37678fc;
  wire v3a6faf3;
  wire v3a53e45;
  wire v376dacb;
  wire v3a579da;
  wire v3a6fdd1;
  wire v37306c2;
  wire v3a71394;
  wire v3a707f3;
  wire v373ddfc;
  wire v37430e7;
  wire v37364af;
  wire v3724926;
  wire v374214d;
  wire v3a65acb;
  wire v3a7075c;
  wire v3a5dd98;
  wire v375f42e;
  wire v3748ded;
  wire v3a5844c;
  wire v373ec92;
  wire v360cffa;
  wire v3a6aaea;
  wire v3770187;
  wire v3a61c5a;
  wire v3753d60;
  wire v3a6dcdc;
  wire v37476fd;
  wire v3a6f7a2;
  wire v3742abe;
  wire v3a5bb85;
  wire v3774463;
  wire v3a710cc;
  wire v3761727;
  wire v8e3f65;
  wire v3a617b4;
  wire v3a6c60e;
  wire v375981e;
  wire v3765b3c;
  wire v373f92e;
  wire v3a7010e;
  wire v3a6267f;
  wire v3762475;
  wire v375d3fd;
  wire v3746c1d;
  wire v37269f4;
  wire v3a67905;
  wire v3725901;
  wire v375af43;
  wire v3a6dd29;
  wire v3a6a1af;
  wire v3744593;
  wire v3a6f406;
  wire v376ba56;
  wire v3a5e7f7;
  wire v3a7076a;
  wire v3774438;
  wire v8b1055;
  wire v37285cd;
  wire v3a70e91;
  wire v3767437;
  wire v3760f4e;
  wire v3730553;
  wire v37307dd;
  wire v372ab46;
  wire v3a6f291;
  wire v3764a2c;
  wire v374b3cf;
  wire v37342ef;
  wire v3a5c94c;
  wire v372b6bf;
  wire v376a2d6;
  wire v3a6f360;
  wire v3759c8c;
  wire v372cbdf;
  wire v3777f6f;
  wire v37697d0;
  wire afa913;
  wire v376ccd6;
  wire v373a59e;
  wire v3a705bd;
  wire v3733a1e;
  wire v377f45d;
  wire v3a5b979;
  wire v377444f;
  wire v375d2cf;
  wire v3765615;
  wire v3a6f240;
  wire v3a71631;
  wire v377c5f4;
  wire v3a55ee6;
  wire v3743434;
  wire v373fc36;
  wire v3740a1b;
  wire v3766ce0;
  wire v37291c0;
  wire v3743c40;
  wire v3771971;
  wire v3741b59;
  wire v3737f8d;
  wire v3764539;
  wire v3727dc9;
  wire v377c02f;
  wire v3a6f410;
  wire v3a70d41;
  wire v3723809;
  wire v3a6f298;
  wire v373e419;
  wire v3730e8f;
  wire v374020a;
  wire v377d769;
  wire v376f9ca;
  wire v3a56bb5;
  wire v372667b;
  wire v373ab3d;
  wire v8455d3;
  wire v3778b73;
  wire v8455cf;
  wire v375b0f9;
  wire v376b14c;
  wire v374d972;
  wire v3a6be07;
  wire v3743eed;
  wire v377c06f;
  wire v376c08d;
  wire v3740b58;
  wire v3777186;
  wire v3a5d51a;
  wire v373cb82;
  wire v3a706a8;
  wire v3753921;
  wire v3a70e87;
  wire v3767d4a;
  wire v375d36b;
  wire v375a55d;
  wire v3726111;
  wire v372c7b7;
  wire v3a6d8af;
  wire v377997c;
  wire v37656e5;
  wire v372e4e1;
  wire v377fc89;
  wire v3a6c96a;
  wire v3734d60;
  wire v23fd8a7;
  wire v3725576;
  wire v376f51a;
  wire v3764ecd;
  wire v3a561aa;
  wire v374a7b4;
  wire v372bbab;
  wire v3a70aef;
  wire v3a54478;
  wire v3a5dc2a;
  wire v3a5ec6b;
  wire v3a64102;
  wire v988a3b;
  wire v3765cd5;
  wire v3759fb9;
  wire v3a70c90;
  wire v3a61de8;
  wire v375b787;
  wire v374066d;
  wire v3a70d09;
  wire v3739940;
  wire v3a69f8e;
  wire v37705df;
  wire a27bd0;
  wire v3a6324e;
  wire v3736b12;
  wire v3764811;
  wire v372cf51;
  wire v3a7151f;
  wire bfa92a;
  wire v3772773;
  wire v3741edb;
  wire v3a6fd64;
  wire v380956b;
  wire v3a6a2d7;
  wire v3a713ab;
  wire v3a5f453;
  wire v373e30f;
  wire v3a66e3d;
  wire v3747b81;
  wire v3740bf5;
  wire v3a6f8e1;
  wire v3a70d6b;
  wire v3777070;
  wire v3a68977;
  wire v3778a97;
  wire v3a65aa5;
  wire v3736a50;
  wire v3747fd2;
  wire v3748eff;
  wire v373a228;
  wire v3a6b896;
  wire v374e47e;
  wire v3a6f8f0;
  wire v3a6a352;
  wire v37699c7;
  wire v372cb06;
  wire v374f8da;
  wire v38069c8;
  wire v372416d;
  wire v3a71073;
  wire v374ca02;
  wire v374e34d;
  wire v3a6f62f;
  wire v374cd6b;
  wire v3a66732;
  wire v375159d;
  wire v3a6f2dc;
  wire v375caa0;
  wire v3a6fb28;
  wire v3750a6f;
  wire v37400ab;
  wire c2b7ee;
  wire v2ff87d3;
  wire v3731476;
  wire v372e8ae;
  wire v3a6c6b1;
  wire v3a6f50c;
  wire v375cda1;
  wire v3a5b05d;
  wire v375c003;
  wire v374620b;
  wire v37431a0;
  wire v376cd19;
  wire v3a71546;
  wire v374bce5;
  wire v37347d9;
  wire v89e294;
  wire v976f99;
  wire v3a56b72;
  wire v3730b57;
  wire v3757261;
  wire v3776150;
  wire v3a70a00;
  wire v372ee20;
  wire v3a6fafb;
  wire v37463ef;
  wire v3a6b4ab;
  wire v373449c;
  wire v375542d;
  wire v3a70104;
  wire v376f152;
  wire v37596fd;
  wire v372f22b;
  wire v3a6fd57;
  wire v3753186;
  wire v23fd886;
  wire v37786a4;
  wire v375e47e;
  wire v3a6b4f6;
  wire v3765968;
  wire v3739e70;
  wire v3a708dd;
  wire v3a56688;
  wire v38087c5;
  wire v373ea19;
  wire v3a6fd52;
  wire v3a71093;
  wire v3a54e47;
  wire v3a70956;
  wire v3a6ffa9;
  wire v37739c7;
  wire v3a70278;
  wire v375003c;
  wire v3769d19;
  wire v37497eb;
  wire v3a5979e;
  wire v3a68a30;
  wire v3a6ca82;
  wire v377b49d;
  wire v373ca53;
  wire v377ef09;
  wire v373ec8f;
  wire v375e30f;
  wire v3753fc9;
  wire a72a7c;
  wire v376653d;
  wire v37284a9;
  wire v3a60584;
  wire v3a6f1de;
  wire v3766d11;
  wire v3a606ee;
  wire v372d279;
  wire v3750d09;
  wire v3806c9a;
  wire v3a5c645;
  wire v3743580;
  wire v376078d;
  wire v3a703f6;
  wire v3736dfe;
  wire v3738373;
  wire v376b678;
  wire v3a7089b;
  wire v3a6ff3e;
  wire v377ee74;
  wire v3761472;
  wire v373ad8b;
  wire v377de57;
  wire a15d51;
  wire v3737f8b;
  wire v3767852;
  wire v3a6ec2a;
  wire v372810e;
  wire v3a6abe5;
  wire v3a56d26;
  wire v37727be;
  wire v3743aee;
  wire v372de52;
  wire v3a7168a;
  wire v377c185;
  wire v3a71061;
  wire v3724577;
  wire v3735708;
  wire v3729823;
  wire d22727;
  wire v376e4da;
  wire v37483c5;
  wire v3a5e239;
  wire v3772f85;
  wire v372a1b6;
  wire v3751e07;
  wire v37400fe;
  wire v372ad15;
  wire v3a70367;
  wire v3766260;
  wire v374b024;
  wire v3728d75;
  wire v3809505;
  wire v37712fa;
  wire v3a70778;
  wire v372b77b;
  wire v3a5c00e;
  wire v3a6e6c9;
  wire v37574b0;
  wire v377a9cb;
  wire v37368ce;
  wire v374d3b3;
  wire v3a7044a;
  wire v375da9d;
  wire v3771ddb;
  wire v377011b;
  wire v375fec7;
  wire v374c33a;
  wire v375efa1;
  wire v3773fbb;
  wire v37613d3;
  wire v375dd2b;
  wire v3765758;
  wire v3a70809;
  wire v3a59a05;
  wire v3a704e3;
  wire v376b1b7;
  wire v3a637a5;
  wire v374e9b8;
  wire v375989b;
  wire v3772696;
  wire v373bf09;
  wire v3a6727a;
  wire v3a6fa8b;
  wire v37556c1;
  wire v3a6b7e9;
  wire v3a7127e;
  wire v37721e3;
  wire v3741e68;
  wire v372594c;
  wire v372ff68;
  wire v3a6f94e;
  wire v3a68848;
  wire v3736968;
  wire v37560b4;
  wire v374e0a4;
  wire v3a63966;
  wire v377ed2d;
  wire v374afa3;
  wire v375b8a2;
  wire v3a71271;
  wire v375c608;
  wire v3746ab6;
  wire v3755744;
  wire v375895e;
  wire v3a70674;
  wire v3773262;
  wire v373e2e5;
  wire v373ae6a;
  wire v373ae4a;
  wire v37729fa;
  wire v375a319;
  wire v373b08f;
  wire v377e431;
  wire v3a6337a;
  wire v3a70588;
  wire v375f46d;
  wire v377af8e;
  wire v374d409;
  wire v3a66920;
  wire v37405a3;
  wire v372f98a;
  wire v37708bb;
  wire v37599b8;
  wire b7dcc5;
  wire v375888e;
  wire v3a6f5b3;
  wire v3a6e124;
  wire v3a5a2c6;
  wire v375da36;
  wire v3a63d83;
  wire v3a5bf21;
  wire v3a62b09;
  wire v3a6eef7;
  wire v39eb413;
  wire v37654e7;
  wire v3a6bb65;
  wire v3a702d0;
  wire v3a58f20;
  wire v3749fd7;
  wire v3a5c2d7;
  wire v23fde7c;
  wire v3a5d04e;
  wire v374ed4f;
  wire v3770751;
  wire v3752c61;
  wire b41a29;
  wire v3755c8b;
  wire v372cfdf;
  wire v3a5f07a;
  wire v3756018;
  wire v375ec0b;
  wire v373dfcc;
  wire v372834c;
  wire v3757601;
  wire v3a5acd5;
  wire v3778da6;
  wire v377e0b8;
  wire v3a70b7d;
  wire v3a6fb29;
  wire v1e379d2;
  wire v3a70cfe;
  wire v3768857;
  wire v377ee3c;
  wire v372bdca;
  wire v375d1d9;
  wire v899d31;
  wire v3a5b3d8;
  wire v3a7129b;
  wire v3a7163e;
  wire v372aed1;
  wire v377a35c;
  wire v37316bb;
  wire v372ba0f;
  wire v37449b3;
  wire v3742655;
  wire v37790df;
  wire v3a6f408;
  wire v3736cdb;
  wire d8a786;
  wire v375f504;
  wire v3779316;
  wire v3728d2a;
  wire v372bcb0;
  wire v376fa94;
  wire v3a7071b;
  wire v3a6ef2a;
  wire v3a6d367;
  wire v376d76c;
  wire v3763c0a;
  wire v3a58eed;
  wire v3742c87;
  wire v3777bf9;
  wire v37343bc;
  wire v376382c;
  wire v3764d0b;
  wire v23fd8c6;
  wire v3756996;
  wire v37474df;
  wire v3a5f642;
  wire v3728fe7;
  wire v3a7169e;
  wire v375c170;
  wire v3a6bdd7;
  wire v372a201;
  wire v3a66460;
  wire v3a67927;
  wire v373602d;
  wire v3a69d9b;
  wire v3a66559;
  wire v38079ff;
  wire v3740e49;
  wire v3a6ab8d;
  wire v3769de7;
  wire v3a62d54;
  wire v377d4dc;
  wire v3a66a6c;
  wire v3762db3;
  wire v376a4d3;
  wire v3a6f07e;
  wire v3a65212;
  wire v3255a31;
  wire v3a701d3;
  wire v3a70a95;
  wire v3733542;
  wire v3a5f5e8;
  wire v37258b7;
  wire v3743c7e;
  wire v38097d8;
  wire v3a6fbe1;
  wire v3a5d63f;
  wire v3751238;
  wire v375a930;
  wire v3743c89;
  wire v373f94e;
  wire v3a67458;
  wire v377f865;
  wire v3740672;
  wire v32559c3;
  wire v377d78b;
  wire v3a70b60;
  wire v3752e8e;
  wire v3734046;
  wire v3774a8f;
  wire v3730452;
  wire v3a7154e;
  wire v3753b7d;
  wire v3739f1f;
  wire v3767578;
  wire v374d4ca;
  wire v373ee41;
  wire v3a61220;
  wire v3a6fee1;
  wire v37543a0;
  wire v3771bed;
  wire v3a6145f;
  wire v3a548f2;
  wire v373d9d3;
  wire v3a5cd5c;
  wire v3a6e548;
  wire v3a6eebb;
  wire v377282c;
  wire v3a6eba9;
  wire v3808eed;
  wire v3779d33;
  wire v3a67e67;
  wire v3a65369;
  wire v373e5a7;
  wire v377f61e;
  wire v374e519;
  wire v3a5e859;
  wire v376156f;
  wire v377e16a;
  wire v37689be;
  wire v3a6e130;
  wire v3a71658;
  wire v3a5ba58;
  wire v3a6ffc0;
  wire v3725ad3;
  wire v3777586;
  wire v3747429;
  wire v3a5ce35;
  wire v377b3be;
  wire v3a702f1;
  wire v37386c0;
  wire v3a626da;
  wire v3755508;
  wire v3741d7c;
  wire v3a64868;
  wire v372e2eb;
  wire v3774d2a;
  wire v376e0f5;
  wire v374cfd8;
  wire v3a6e82d;
  wire v372b32f;
  wire v3729189;
  wire v372bbc7;
  wire v3a64ba3;
  wire v3763ad3;
  wire v3a7136f;
  wire v380713a;
  wire v3752fe9;
  wire v3732128;
  wire v3a6f77a;
  wire v37403ea;
  wire v3a70b39;
  wire v374a233;
  wire v3a62a68;
  wire v37494ee;
  wire v3a6efce;
  wire v3a6fda7;
  wire v3a70c54;
  wire v397d85e;
  wire v3a54497;
  wire v38088e1;
  wire v3748656;
  wire v3734ec1;
  wire v373ee51;
  wire v372642c;
  wire v3762a9f;
  wire v375297d;
  wire v3a55347;
  wire v375c6c7;
  wire v374dafa;
  wire v3a6f145;
  wire v376067f;
  wire v37683c2;
  wire v3a6fc05;
  wire v3774c55;
  wire v373ff9a;
  wire v3a64293;
  wire v377ae0c;
  wire v3a63f49;
  wire v3726980;
  wire v3a63d5f;
  wire v3767e38;
  wire v3765f99;
  wire v3773697;
  wire v3a70d43;
  wire v375e94c;
  wire v3a6f62b;
  wire v377115d;
  wire v3a7130e;
  wire v374326f;
  wire v3759501;
  wire v375634b;
  wire v376081b;
  wire v37bfd10;
  wire v37535e7;
  wire v37640fd;
  wire v377b0a0;
  wire v3a7160f;
  wire v3808e85;
  wire v3a705f4;
  wire v3737c86;
  wire v3a63df6;
  wire v372d366;
  wire v3a6f767;
  wire v3727662;
  wire v375ed63;
  wire v3728230;
  wire v376981e;
  wire v3745e51;
  wire v3735f9b;
  wire v376803b;
  wire v3731478;
  wire v374f126;
  wire v3a6c549;
  wire v2acaf2d;
  wire v376e17e;
  wire v92acd8;
  wire v3a60cbd;
  wire v3a60e7e;
  wire v3724be1;
  wire v3756de3;
  wire v8e4f94;
  wire v3748016;
  wire v372f231;
  wire v3a6a78c;
  wire v3a56bf0;
  wire v3760bfd;
  wire v3a544de;
  wire v373f883;
  wire v35b9d5e;
  wire v377e639;
  wire v2aca264;
  wire v373c2a2;
  wire v375fe03;
  wire v3758ee1;
  wire v376755f;
  wire v3750797;
  wire v3a67d83;
  wire v374c3ff;
  wire v3a69390;
  wire v3767e55;
  wire v3a5f12b;
  wire v3a6f537;
  wire v3a71373;
  wire v3a700c1;
  wire v372eaf3;
  wire v3750ce8;
  wire v3a6aaaa;
  wire v37571c0;
  wire v374cbc4;
  wire v376c5af;
  wire v3a53f85;
  wire v3762f98;
  wire v3a702a8;
  wire v33790e4;
  wire v3748f17;
  wire v3a588ec;
  wire v37755d5;
  wire v377472b;
  wire v3738c2e;
  wire v3760aa7;
  wire v373f401;
  wire da4c01;
  wire v3726865;
  wire v3a6f29c;
  wire v3760d46;
  wire v376c4e8;
  wire v3759bd0;
  wire v3732775;
  wire v3761433;
  wire v3736ee0;
  wire v3809487;
  wire v37267a5;
  wire v1e37b74;
  wire v37c014f;
  wire v375aceb;
  wire v377b626;
  wire v3779337;
  wire v373f125;
  wire v3a6b572;
  wire v3735153;
  wire v37435a9;
  wire v373324d;
  wire v37280b7;
  wire v376ed30;
  wire v3a6f579;
  wire v3a5a853;
  wire v97f405;
  wire v3a6c91f;
  wire v3a5e2b9;
  wire v3768aa4;
  wire v3745d8c;
  wire v3a5aaed;
  wire v376b908;
  wire v3a60c05;
  wire v37509a3;
  wire v3a70e62;
  wire v3a6f5fe;
  wire v373422b;
  wire v3a69bfd;
  wire v3731737;
  wire v375d42d;
  wire v376e9fd;
  wire v375a463;
  wire v3a6fd5a;
  wire dafc4e;
  wire v3a70894;
  wire v3a6f11e;
  wire v375da6a;
  wire v372f739;
  wire v3a71483;
  wire v864fe4;
  wire v376e358;
  wire v3745fd1;
  wire v377845d;
  wire v3759602;
  wire v372da7e;
  wire v374f6c0;
  wire v3a61661;
  wire v3a63fd5;
  wire v3a6f4e0;
  wire v3745f63;
  wire v37511f6;
  wire v38076b3;
  wire v3a71241;
  wire v3a71156;
  wire v3a71442;
  wire v3723de9;
  wire v373f418;
  wire v37378a3;
  wire v3a5c9d7;
  wire v374d042;
  wire v375b247;
  wire v3a6f7e4;
  wire v3a5aff3;
  wire v3a67182;
  wire v3a6e40f;
  wire v375fbae;
  wire v377c35c;
  wire v3a6ebd0;
  wire v3a5cb92;
  wire v373908c;
  wire v375f67d;
  wire v37508c4;
  wire v3a6eb91;
  wire v3a6ecd1;
  wire v37462ee;
  wire v3771be6;
  wire v3a69c64;
  wire v3725d5a;
  wire v3a6f411;
  wire v374247d;
  wire v3a6fb07;
  wire v3a6fd02;
  wire v3a64355;
  wire v37232aa;
  wire v3771cac;
  wire v3a5b660;
  wire v375982a;
  wire v37592c9;
  wire v3774b2b;
  wire v3729263;
  wire v373f461;
  wire v3a5e999;
  wire v3377b0f;
  wire v3a5a210;
  wire v3a6dfec;
  wire v37c36cb;
  wire v3a70efe;
  wire v360d177;
  wire v3773c10;
  wire v3a57fa1;
  wire v3a5fe00;
  wire v3762f27;
  wire v37435b7;
  wire v3730f34;
  wire v375e516;
  wire v3733940;
  wire v373395b;
  wire v3756afd;
  wire v37434c6;
  wire v3a58fe2;
  wire v37332bf;
  wire v3740451;
  wire v3a6eee3;
  wire v3a5b333;
  wire v1e378ce;
  wire v3a5aef2;
  wire v3a614df;
  wire v376d4cb;
  wire v376fe0c;
  wire v374d6dd;
  wire v3739896;
  wire v375306b;
  wire v37379fc;
  wire v3a714bd;
  wire v3a62524;
  wire v373cdb7;
  wire ae7027;
  wire v372beb8;
  wire d0a687;
  wire v3a5cfdb;
  wire v3a65546;
  wire v3777749;
  wire v3754543;
  wire v3764381;
  wire v373899b;
  wire v3740ee1;
  wire v3a29842;
  wire v3748fba;
  wire v375b878;
  wire v3a6b6ef;
  wire v3a711e5;
  wire v3765c1f;
  wire v3a64f54;
  wire v3763952;
  wire v376ee65;
  wire v37300a5;
  wire v375f2ec;
  wire v3a6c580;
  wire v3a56aeb;
  wire v37301f5;
  wire v3774e64;
  wire v3a71130;
  wire v376ef3f;
  wire v3728b05;
  wire v3772dc6;
  wire v3a6fe5d;
  wire v8d428b;
  wire v372f87f;
  wire v37674a5;
  wire v3731e31;
  wire v3723701;
  wire v3756ef1;
  wire v3751d9c;
  wire v373c627;
  wire v3a6f972;
  wire v37772bf;
  wire v3a66ff2;
  wire v1e3825d;
  wire v3a5759a;
  wire v3738766;
  wire v377b5c4;
  wire v23fe10f;
  wire v2acafdf;
  wire b6ae10;
  wire v377db88;
  wire v3728813;
  wire v37623f5;
  wire v37519bf;
  wire v3a5dd70;
  wire v37286e7;
  wire v372d525;
  wire v3760237;
  wire v3738457;
  wire v3a6a48e;
  wire v374ab22;
  wire v3a6178c;
  wire v3736f61;
  wire v374a2f3;
  wire v3771c85;
  wire v357742d;
  wire v3730055;
  wire v3a6f831;
  wire v3a55b39;
  wire v3a70267;
  wire v3258dd9;
  wire v377a470;
  wire d09db6;
  wire ab11fe;
  wire v3765cf3;
  wire v9d4353;
  wire v3771607;
  wire v3737028;
  wire v3a6f378;
  wire v380956d;
  wire v3765ef0;
  wire v3a709f8;
  wire v372cab6;
  wire v37251e7;
  wire v376ef7a;
  wire v375937f;
  wire v3a53cfe;
  wire v3724475;
  wire v3a6cab1;
  wire v37521af;
  wire v3a60618;
  wire v37523f4;
  wire v3a6f9a8;
  wire v374720c;
  wire v3772d27;
  wire v3a64f9b;
  wire v3a61237;
  wire v3a6ebe7;
  wire v375d182;
  wire v3a67e2e;
  wire v37443d6;
  wire v3a63f05;
  wire v3751b0e;
  wire v376da28;
  wire v37625b7;
  wire v3a6f748;
  wire v3733da3;
  wire v377149d;
  wire v3741ae7;
  wire v3a6f9c4;
  wire v373d27f;
  wire v3a5b0dd;
  wire v372dffe;
  wire v3a6406d;
  wire v377286e;
  wire v37676b8;
  wire v3762700;
  wire v3a6f22b;
  wire v3724112;
  wire v3a65f3e;
  wire v3773871;
  wire v3747346;
  wire v3a594a5;
  wire v3767d1b;
  wire v3767a93;
  wire v372988e;
  wire v3a6581b;
  wire v39ebb7b;
  wire v37533e5;
  wire v3a65b3e;
  wire v376de99;
  wire v3731a1f;
  wire v376fb60;
  wire v3736fb6;
  wire v3779797;
  wire v372b10b;
  wire v377a13b;
  wire v3a57108;
  wire v3746d57;
  wire v375f83b;
  wire v3a61f9b;
  wire v3757adc;
  wire v3a59b8a;
  wire v3726905;
  wire v377aa7a;
  wire v3a70912;
  wire v3743879;
  wire v3a662c7;
  wire v377c671;
  wire v37722e5;
  wire v3756206;
  wire v3a63bdb;
  wire v3723676;
  wire v372d3e8;
  wire v3722b42;
  wire v37459dd;
  wire v3a704b1;
  wire v9aa8f3;
  wire v37619dc;
  wire v3806912;
  wire v3a6f22f;
  wire v3a704ee;
  wire v3a6ff4f;
  wire v372a3af;
  wire v3746641;
  wire v3746d49;
  wire bf5753;
  wire v373ae02;
  wire v37bfd3a;
  wire v373cc82;
  wire v375a1a7;
  wire v377ef58;
  wire v373e27e;
  wire v3770f97;
  wire v3759eb6;
  wire v3a6bcf9;
  wire v3a5a220;
  wire v23fd98d;
  wire v37271f9;
  wire v3a71456;
  wire v3a67d2e;
  wire v3a5d673;
  wire v3745020;
  wire v3749207;
  wire v373132b;
  wire c0b4d9;
  wire v3763eac;
  wire v372fa02;
  wire v3768573;
  wire v3731099;
  wire v37701fd;
  wire v3766285;
  wire v3a705b9;
  wire v3734062;
  wire v3a68f5f;
  wire v3728399;
  wire v3760bdd;
  wire v375168a;
  wire v3a6c6aa;
  wire v3a5b9ea;
  wire v37736ad;
  wire v3773856;
  wire v3a6fc7b;
  wire v3750134;
  wire v372d9e0;
  wire v37574d3;
  wire v3a7029f;
  wire v375ecff;
  wire v374f178;
  wire v37698a1;
  wire v3a6f388;
  wire v375eba9;
  wire v2ff9189;
  wire v31c3043;
  wire v3a5d41e;
  wire v3a54242;
  wire v376ba96;
  wire v37283c0;
  wire v375243f;
  wire v3a6d6ff;
  wire v3733083;
  wire b77306;
  wire v37756ef;
  wire v376f45b;
  wire v3765960;
  wire v3806bd9;
  wire v3a705e1;
  wire v3a706d1;
  wire v3a6fa6e;
  wire v377934a;
  wire v37362fc;
  wire v3a70dd6;
  wire v3a62a8c;
  wire v373ccc7;
  wire v3772185;
  wire v360d036;
  wire v376eb3f;
  wire v3a6f968;
  wire v373e933;
  wire v3a6eb2d;
  wire v374f677;
  wire v3a6ebcd;
  wire v3a715e2;
  wire v3a70f3e;
  wire v376dcdc;
  wire v3a70832;
  wire v37617de;
  wire v372526a;
  wire v2925ce0;
  wire v3737415;
  wire v3a70a96;
  wire v3762072;
  wire v3a6ec0a;
  wire v3743b98;
  wire v37c023b;
  wire v8a9c95;
  wire v3a7014c;
  wire v376b33c;
  wire v3a56f66;
  wire v3741f39;
  wire v3a5948d;
  wire v3765a98;
  wire v372f747;
  wire v373449a;
  wire v3743ada;
  wire v377a5df;
  wire v373f10d;
  wire v3722a9c;
  wire v3737c3f;
  wire v3755ffc;
  wire v3a6377a;
  wire v376a3cb;
  wire v3a67524;
  wire v3733c82;
  wire v3777d79;
  wire v3a6a7b4;
  wire v376ef36;
  wire v3a70d42;
  wire v3a59d47;
  wire v3a6f4f1;
  wire v3a584f1;
  wire v3762a49;
  wire v3a60c38;
  wire v3a6ca4e;
  wire v377b734;
  wire v3a6a435;
  wire v372745b;
  wire b95be3;
  wire v376a220;
  wire v3a591b4;
  wire v3a70952;
  wire v3746dc9;
  wire v3a6f93a;
  wire v3779df7;
  wire dac24d;
  wire v3745939;
  wire v3a6a52b;
  wire v3a70929;
  wire v373227a;
  wire v375582f;
  wire v3a6f5d2;
  wire v3a71460;
  wire v3a59ffa;
  wire v3a6d18a;
  wire v372a0bd;
  wire v3741dce;
  wire v3a6a1f4;
  wire v37671ad;
  wire v325b5e0;
  wire v2619b54;
  wire v375e03c;
  wire v3a6c860;
  wire v374e418;
  wire v3a706b5;
  wire v3a703e0;
  wire v373d62b;
  wire v373619d;
  wire v86d306;
  wire v37777ba;
  wire v3a2a14e;
  wire v3762245;
  wire b318d6;
  wire v376b031;
  wire v37478bc;
  wire v374bf0f;
  wire v376d57d;
  wire v37581d2;
  wire v3a65b64;
  wire af345a;
  wire v3a6e543;
  wire v372b2aa;
  wire v372f853;
  wire v3a70b4a;
  wire v374a91e;
  wire v3767adc;
  wire v37535c4;
  wire v3747ed4;
  wire v374d153;
  wire v3775e2e;
  wire v38087ba;
  wire v3746dbf;
  wire v3763846;
  wire v3777b5b;
  wire v3776fc5;
  wire v2acb06f;
  wire v3753093;
  wire v3734419;
  wire v23fdf76;
  wire v3756506;
  wire v374d52a;
  wire v3a71243;
  wire v3765305;
  wire v3a6ff29;
  wire v37286e9;
  wire v373c04a;
  wire v377faae;
  wire v374074a;
  wire v37502f1;
  wire v373aca2;
  wire v3739815;
  wire v3769bdb;
  wire v372fb58;
  wire v376bb7a;
  wire v37357ce;
  wire v3766b26;
  wire v3a6d627;
  wire v3a6c7ab;
  wire v376ccdf;
  wire v376761d;
  wire v3a70f4e;
  wire v3731fd2;
  wire v3778628;
  wire v3a6f36f;
  wire v3a5fd6a;
  wire v3722e5e;
  wire v3755312;
  wire v377dfec;
  wire v3743ef0;
  wire v3a2ad1b;
  wire v3a6f2d7;
  wire v372797f;
  wire v3a62d7d;
  wire v3a6f402;
  wire v3a564a8;
  wire v373cb2d;
  wire v3a5fe72;
  wire v37321b8;
  wire v3766238;
  wire v3a622d0;
  wire v37658b1;
  wire v1e37ab9;
  wire v376b734;
  wire v3775aea;
  wire v373687f;
  wire v3a68e39;
  wire v3a62041;
  wire v374f3e3;
  wire v373fd72;
  wire v3735ecd;
  wire v372cdb8;
  wire v3765ab2;
  wire v375c7a9;
  wire v3a6f365;
  wire v3a67cfe;
  wire v373f82c;
  wire v3a6f64e;
  wire v3750613;
  wire v3a61445;
  wire v3727bca;
  wire v3737a29;
  wire v3735906;
  wire v3a57cd0;
  wire v3a651b5;
  wire v3a56b19;
  wire v3768bbc;
  wire v376d2f4;
  wire v3764ad1;
  wire v377e70d;
  wire v377623c;
  wire v377d6f9;
  wire v3a6143f;
  wire v3753e00;
  wire v3739386;
  wire v3a70ad4;
  wire v3a6f17e;
  wire v3759b11;
  wire v3a701a6;
  wire v375c379;
  wire v376d817;
  wire v377fc87;
  wire v3737e8c;
  wire v37288db;
  wire v3a65b53;
  wire v3747c3d;
  wire v3a6f0bc;
  wire v375d4aa;
  wire v3a60332;
  wire v3a55cf2;
  wire v3723b86;
  wire v3749cdf;
  wire v372cb28;
  wire v37274ef;
  wire v372298c;
  wire v3a7096e;
  wire v372ce88;
  wire v375deaa;
  wire v375b01a;
  wire v1e37dd9;
  wire v377c7b2;
  wire v377327b;
  wire v39a53b3;
  wire v372c565;
  wire v377bdbe;
  wire c22b44;
  wire v3758c35;
  wire v3a70e49;
  wire v3767642;
  wire v3807ddf;
  wire v372ac5c;
  wire v3773ba2;
  wire v3755e29;
  wire v376bb64;
  wire v3755aef;
  wire v376655b;
  wire v372fb60;
  wire v3809112;
  wire v3a71308;
  wire v3763424;
  wire v3a5e1ab;
  wire v3a60181;
  wire v3723aa8;
  wire v3a68f04;
  wire v373b548;
  wire v3a60f18;
  wire v3772b7e;
  wire v3763e44;
  wire v37360d1;
  wire v3a6fad5;
  wire v3a70e45;
  wire v377a0da;
  wire v3a60a9b;
  wire v3776923;
  wire v372e99c;
  wire v3a5bbc1;
  wire be181b;
  wire v374ac2e;
  wire v37500ae;
  wire v3728fa6;
  wire v3a54677;
  wire v2ff87a0;
  wire v3774063;
  wire v3a5d2f0;
  wire v39eb4e4;
  wire v376d3e2;
  wire v373c8bb;
  wire v37429d9;
  wire v374eddc;
  wire v374b7f6;
  wire v375685c;
  wire v37536fd;
  wire v3779c8e;
  wire v375b400;
  wire v37650e4;
  wire v3a611b0;
  wire v375eaac;
  wire v37555cd;
  wire v37344c6;
  wire v374189b;
  wire v3759623;
  wire v3a60a40;
  wire v3777e0a;
  wire v376c687;
  wire v3760748;
  wire v3a71455;
  wire v374d926;
  wire v3a70ee9;
  wire v374bd6a;
  wire v3732202;
  wire v372bffa;
  wire v3756f42;
  wire v375409b;
  wire v37520c4;
  wire v3726f89;
  wire v373fbb6;
  wire v3a701d1;
  wire v3a70397;
  wire v3a5c350;
  wire v376aad2;
  wire v373d27a;
  wire v3759de1;
  wire v3756ecd;
  wire v373a02b;
  wire v374d9fe;
  wire v374bfa2;
  wire v3a63938;
  wire v3a643a0;
  wire v3a6f2a2;
  wire v377e142;
  wire v3a57e40;
  wire v374b5d9;
  wire v373bb0f;
  wire v3a6a1e9;
  wire v3740374;
  wire v3728a12;
  wire v3a71283;
  wire v37328da;
  wire v37545ea;
  wire v3a5be6d;
  wire v374f75e;
  wire v3a6a6eb;
  wire v3a5ed4b;
  wire v3775654;
  wire v3733aa5;
  wire v374ac24;
  wire v3726a7e;
  wire v3a6fe5f;
  wire v3a5e985;
  wire v372967b;
  wire v3a6e614;
  wire v3734632;
  wire v3a705d0;
  wire v3a53f1c;
  wire v3768c98;
  wire v375b777;
  wire v3726a09;
  wire v375889d;
  wire v3749b2e;
  wire v3a6c40d;
  wire v1e382dc;
  wire v3a7112d;
  wire v3a674a8;
  wire v376ee08;
  wire v3a6fbee;
  wire v374b393;
  wire v3a53e30;
  wire v3760c1b;
  wire v3735675;
  wire v377da10;
  wire v37320f4;
  wire v37535d9;
  wire v372f7b4;
  wire v23fe295;
  wire v37514c2;
  wire v37563cf;
  wire v3a708f7;
  wire v377dd0d;
  wire v3775723;
  wire v3757f96;
  wire v39a52b7;
  wire v3728650;
  wire v3a56eeb;
  wire v3a64a83;
  wire v23fde7b;
  wire v37546c9;
  wire v3768a7b;
  wire v377aaba;
  wire v376ad77;
  wire v3722d5a;
  wire v3731eca;
  wire v374df25;
  wire v3a6ff56;
  wire v3a6eab8;
  wire v38090e9;
  wire v3a701c7;
  wire v3724394;
  wire v3a6fdd2;
  wire v37529d9;
  wire v37326a0;
  wire v3a6e118;
  wire v377e2e3;
  wire v374d121;
  wire v375161a;
  wire v3744577;
  wire v3748900;
  wire v376cd91;
  wire v373c978;
  wire v3a6fb27;
  wire v374165a;
  wire v3a6b2c9;
  wire v3748b43;
  wire v3a6f9e7;
  wire v376673b;
  wire v3724908;
  wire v375e099;
  wire c45930;
  wire v374ddef;
  wire v3743dff;
  wire v3a714b4;
  wire v37551b0;
  wire v3a71161;
  wire v372b902;
  wire v3a584be;
  wire v3a59979;
  wire v3729b52;
  wire v39ebb63;
  wire v3750c57;
  wire v3a5f853;
  wire v905dc4;
  wire v373a560;
  wire v3a6ac26;
  wire v373c151;
  wire v3749a89;
  wire v3a70cc0;
  wire v3767d4e;
  wire v377ddae;
  wire v3a56864;
  wire v3744417;
  wire v3a714aa;
  wire v373959b;
  wire v3a6fbd0;
  wire v37238b1;
  wire v3a70c34;
  wire v374a6a5;
  wire v372a98e;
  wire v3a6ef18;
  wire v3a601a0;
  wire v376a08d;
  wire v3a6a895;
  wire v375d5ac;
  wire v3760ba3;
  wire v3a66c20;
  wire v3a702ce;
  wire v3750f20;
  wire v37795d9;
  wire v93c94e;
  wire v3a6efcd;
  wire v37374a1;
  wire v376c652;
  wire v376c4c9;
  wire v372ef7c;
  wire v337793f;
  wire v3773fdc;
  wire v3a608b9;
  wire v376b6c8;
  wire v3a70e0f;
  wire v3a714fd;
  wire v373e21a;
  wire v1e379fe;
  wire v374ab4f;
  wire v374e77f;
  wire v374fe0f;
  wire v3734a92;
  wire v3a5be15;
  wire bbba6b;
  wire v37549cd;
  wire v3a6fe41;
  wire v39ebb2e;
  wire v3a6a036;
  wire v372e27b;
  wire v377ecac;
  wire v37266df;
  wire v3a6f54b;
  wire v374d010;
  wire v376e7a5;
  wire v375a12e;
  wire v3a70ff7;
  wire v37278f5;
  wire v3751a94;
  wire v3762db6;
  wire v3a6681e;
  wire v375139a;
  wire v3a641c0;
  wire v37742ca;
  wire v3733711;
  wire v373373d;
  wire v377050c;
  wire v3769310;
  wire v3727cec;
  wire v37715b9;
  wire v3a6fa97;
  wire v372a450;
  wire v3729ddd;
  wire v3a6b1ab;
  wire v3a6255b;
  wire v3731300;
  wire v3760b3d;
  wire v3a6f817;
  wire v3753ccf;
  wire v3a5acc7;
  wire v3a713b7;
  wire v375a2ff;
  wire v3a63d05;
  wire v37419fa;
  wire ce7a16;
  wire v3741286;
  wire v372b0cd;
  wire b09623;
  wire v372ef9b;
  wire v95d97e;
  wire v3732034;
  wire v1e37869;
  wire v3a6fd47;
  wire v375a18e;
  wire v37367da;
  wire v3a6f8f9;
  wire v3a6e468;
  wire v374df64;
  wire a34d2b;
  wire v37592d0;
  wire v3a683e2;
  wire v3766a28;
  wire v374a97c;
  wire v3738745;
  wire v3a5d80f;
  wire c8a454;
  wire v3752f78;
  wire v3774074;
  wire v373a391;
  wire v374c937;
  wire v3758233;
  wire v3760549;
  wire v2aca978;
  wire v372c6cb;
  wire v3a62251;
  wire v1e37481;
  wire v3a6fad0;
  wire v3a5b850;
  wire v3732d4b;
  wire v3a70626;
  wire v3a6ec7a;
  wire v3749caa;
  wire v374074d;
  wire v373ddca;
  wire v3378c57;
  wire v37541a7;
  wire v3a5ba28;
  wire v3a5cf5e;
  wire v3756810;
  wire bad3a6;
  wire v374961f;
  wire v3a5d923;
  wire v3736a37;
  wire v376ebdd;
  wire v3768931;
  wire v3727eca;
  wire v2092ab0;
  wire v3737ea9;
  wire v3a65bad;
  wire v372e4cf;
  wire v3a70513;
  wire v376eeea;
  wire v3728a6a;
  wire v2619ae8;
  wire v2acaff4;
  wire v3772d9a;
  wire v3739c30;
  wire v374d85e;
  wire v3760bf8;
  wire v372c9ac;
  wire v37606e5;
  wire v376938e;
  wire v3767b75;
  wire v3a5c33d;
  wire v372c46e;
  wire v3764ddc;
  wire v376a2df;
  wire v8f7302;
  wire v3a6eff8;
  wire v3a6f85a;
  wire v3724249;
  wire v3754bc9;
  wire v374b362;
  wire v3a6aef7;
  wire v3756045;
  wire v3a62ad8;
  wire v3a6dd4d;
  wire v376b8f1;
  wire v3a6008f;
  wire v3a6f7b0;
  wire v3765c35;
  wire v373d9e4;
  wire v375567c;
  wire v3a542c0;
  wire v372d842;
  wire v89a228;
  wire v3748301;
  wire v377d850;
  wire v37798da;
  wire v3779403;
  wire v3a703ab;
  wire v375c724;
  wire v3a6ca15;
  wire v376f858;
  wire v3a676ce;
  wire v3a6fb68;
  wire v376bbbe;
  wire v37342e7;
  wire v374a0b1;
  wire v3769ba9;
  wire v374bab6;
  wire v37782de;
  wire v37518e7;
  wire v374472d;
  wire v3a711fd;
  wire v373df91;
  wire v3768e31;
  wire v3742fbf;
  wire v9d97fe;
  wire v373afb4;
  wire v3a6efe8;
  wire v372ac49;
  wire v374c5b2;
  wire v372f173;
  wire v374d01c;
  wire v3769a16;
  wire v3a61853;
  wire v3736785;
  wire v3726ef1;
  wire v3730181;
  wire v37672ac;
  wire v376b087;
  wire v3723af9;
  wire v377041c;
  wire v37266d1;
  wire v377a27f;
  wire v37347cd;
  wire v375dd80;
  wire v37499a9;
  wire v3779e38;
  wire v3766f13;
  wire v3a5e80e;
  wire v373edbe;
  wire v373b381;
  wire v3a7112c;
  wire v372d8ff;
  wire v3748f81;
  wire v377adf7;
  wire v3a5c064;
  wire v3738641;
  wire v3a56d2e;
  wire v9259bc;
  wire v3764c4c;
  wire v3a67d66;
  wire v377bdb8;
  wire v3770415;
  wire v374430e;
  wire v3a6f426;
  wire v3a67aa1;
  wire v3779e70;
  wire v3a6bd87;
  wire v3a6b714;
  wire v373fbb4;
  wire ca01e4;
  wire v3758a96;
  wire v372dfc3;
  wire v374d741;
  wire v3a56118;
  wire v3776f42;
  wire v3778998;
  wire v376bfe6;
  wire v3762729;
  wire v377824e;
  wire v380714c;
  wire v3a6f97b;
  wire v375f852;
  wire v3a6f35b;
  wire v3a65607;
  wire v3a7080c;
  wire v373461a;
  wire v37482f5;
  wire v372509d;
  wire v3a56dff;
  wire v3770621;
  wire v376bb04;
  wire v375f020;
  wire v376e1c4;
  wire v3a709a6;
  wire v375b902;
  wire v3a6f598;
  wire v3730122;
  wire v3727eb8;
  wire v3739336;
  wire v37560ff;
  wire v3756820;
  wire v37684b7;
  wire v3749ea2;
  wire v3748ca5;
  wire v375338a;
  wire v374af0d;
  wire v3752e65;
  wire v37646c7;
  wire v3a6ac60;
  wire v3a702d9;
  wire v3767f52;
  wire v3a62973;
  wire v3a704a8;
  wire v372d8fa;
  wire v376cc20;
  wire v376e1ed;
  wire v3a6eb2b;
  wire v3a56049;
  wire v3806ce9;
  wire v372ccbe;
  wire v3a712e7;
  wire v3735c51;
  wire v3774a13;
  wire v3a61392;
  wire v372ccbb;
  wire v375ca08;
  wire v2acb5a7;
  wire v3a5e591;
  wire v3809f65;
  wire v3755c7c;
  wire v3a6f434;
  wire v37284d5;
  wire v3748179;
  wire v3a7104e;
  wire v3a6d614;
  wire v37511c6;
  wire v3a6f740;
  wire v3765109;
  wire v3a6f749;
  wire v373f06c;
  wire v3a6be05;
  wire v374c8b8;
  wire v360d0fb;
  wire v373db5d;
  wire v375a52a;
  wire v3774737;
  wire v3a7079a;
  wire v37582e7;
  wire v3808f2f;
  wire v375398e;
  wire v37770ab;
  wire v3759421;
  wire v377244a;
  wire v380a188;
  wire v3a6f57c;
  wire v3a5beb5;
  wire v3744131;
  wire v3a70e46;
  wire v377f13c;
  wire v372545e;
  wire v325c94d;
  wire v376f5e1;
  wire v3774dbe;
  wire v376ba33;
  wire v377ef47;
  wire v372d851;
  wire v375cbdf;
  wire v3a70ba8;
  wire v372a53e;
  wire v375069a;
  wire v3730d6c;
  wire v3745734;
  wire v372bc4c;
  wire v3a7033f;
  wire v3a6ff5e;
  wire v3a6f568;
  wire v3a6a9cf;
  wire v3776aa8;
  wire v3a60711;
  wire v3755806;
  wire v360cdfe;
  wire v3a6e94b;
  wire v375c7b6;
  wire v3a58cc0;
  wire v3a6ee22;
  wire v372706d;
  wire v3776fa4;
  wire v3a6f052;
  wire v372ac83;
  wire v3a69bf4;
  wire v3750775;
  wire v3729991;
  wire v376a96b;
  wire v372b1b5;
  wire v3744380;
  wire v373a772;
  wire v9f9402;
  wire v3745539;
  wire v374fe44;
  wire v3a71297;
  wire v3a71417;
  wire v37522d3;
  wire v3a5bcfd;
  wire c88c38;
  wire v3a70ad2;
  wire v3a712a8;
  wire v372cfec;
  wire v376e9b7;
  wire v372c095;
  wire v377506b;
  wire v3746745;
  wire v3763efc;
  wire v3a612a3;
  wire v376fd05;
  wire v3764af7;
  wire v3745053;
  wire v374e459;
  wire v3a6963f;
  wire v3777642;
  wire v3771dda;
  wire v375a086;
  wire v3753dbd;
  wire v372658a;
  wire v3754981;
  wire v373257d;
  wire v3a680bd;
  wire v375706b;
  wire v37452e7;
  wire v3a5936a;
  wire v3a706eb;
  wire v372a79d;
  wire v3a5a035;
  wire v35ba1a5;
  wire v3a71611;
  wire v374bdea;
  wire v377c620;
  wire v3752348;
  wire v3a6fe22;
  wire v3774e33;
  wire v3a5f439;
  wire v374e7b5;
  wire v3a616f0;
  wire v3a5f485;
  wire v374cab5;
  wire v3a2a13a;
  wire v3730cde;
  wire v373769f;
  wire v375501e;
  wire v3737e2e;
  wire v377a10f;
  wire v3a67ffd;
  wire v372ff72;
  wire v3a5be57;
  wire v3736cb3;
  wire v3759fd0;
  wire v2092bdc;
  wire v376bad7;
  wire v3a68e46;
  wire v37324da;
  wire v3724b26;
  wire v376d191;
  wire v3809e71;
  wire v3726994;
  wire v3771da0;
  wire v37699ec;
  wire v374e3c1;
  wire v3730a22;
  wire v376644e;
  wire v376d432;
  wire v3734473;
  wire v3a709db;
  wire v375ad9f;
  wire v3770a68;
  wire v3750b5b;
  wire v3a711df;
  wire v1e37cf9;
  wire v3a702f2;
  wire v375cbe2;
  wire v2092ac3;
  wire v372e40f;
  wire v37710fb;
  wire v3a704cb;
  wire v377ce1c;
  wire v37702a1;
  wire v3a588e5;
  wire v3a7092f;
  wire v37656cd;
  wire v3a606e6;
  wire v376df9f;
  wire v32558c4;
  wire v35b70fa;
  wire v3a70311;
  wire v3a29760;
  wire v3a5f030;
  wire v3736dc2;
  wire v3a7125c;
  wire v377163d;
  wire v3747a5f;
  wire v3a6fbf1;
  wire v3764b6e;
  wire v3753fb7;
  wire v3750e0b;
  wire v3a6184c;
  wire v3a6fb56;
  wire v3743f4d;
  wire v3724a65;
  wire v3a616fb;
  wire v374e05d;
  wire v3757858;
  wire v3764fe1;
  wire v376ae69;
  wire v3a65096;
  wire v372e479;
  wire v3a69063;
  wire v3728916;
  wire v37424a9;
  wire v3767919;
  wire v1e37c44;
  wire v377324f;
  wire v37555cb;
  wire v37471a7;
  wire v374ddc7;
  wire v3a715fa;
  wire v375d06d;
  wire v3773524;
  wire v375e64d;
  wire v3a6f356;
  wire v3771ea7;
  wire v372a4c1;
  wire v376652f;
  wire v3a70647;
  wire v375cfaa;
  wire v3a70afe;
  wire v3744151;
  wire v3a6ff6e;
  wire v377e905;
  wire v3772f3c;
  wire v3a5cb20;
  wire v3a56a2c;
  wire v3a70f51;
  wire v3a6f944;
  wire v374be0c;
  wire v376b063;
  wire v376f4b9;
  wire v3760ac5;
  wire v377a75f;
  wire v372d24d;
  wire v3a70bc8;
  wire v373cb54;
  wire v376e72d;
  wire v3724b1c;
  wire v37293ee;
  wire v372b231;
  wire v37754e6;
  wire v373f012;
  wire v3a6fb24;
  wire v3a61604;
  wire v372c614;
  wire v3a58057;
  wire v3756a04;
  wire v3743f3b;
  wire v37302b7;
  wire v3778baf;
  wire v3a7032a;
  wire v3a6fc67;
  wire v374fe51;
  wire v3737695;
  wire v37252c2;
  wire v360d136;
  wire v3741869;
  wire v372309d;
  wire v37258b4;
  wire v37611fb;
  wire v372fd4a;
  wire v3728f0a;
  wire v377504f;
  wire v37303aa;
  wire v3a6f668;
  wire v375833e;
  wire v3a70142;
  wire v374a3db;
  wire v375604f;
  wire v3757f09;
  wire v3729b33;
  wire v377b1db;
  wire v3779cb7;
  wire v3a5788f;
  wire v376ba53;
  wire v376187f;
  wire v374233c;
  wire v3a6fd91;
  wire v3a6f13e;
  wire v376e3a0;
  wire v3760ba8;
  wire v3726077;
  wire v3737a76;
  wire v3a709e1;
  wire v376773f;
  wire v3739a53;
  wire v375feba;
  wire v3a6f09f;
  wire v374d847;
  wire v3809390;
  wire v3755f2d;
  wire v3a6a0c4;
  wire v3724e61;
  wire v377f730;
  wire v3766c97;
  wire v3731e91;
  wire v373f2d8;
  wire v3a71561;
  wire v3a5538a;
  wire v372a0f7;
  wire v3a6823d;
  wire v377362f;
  wire v3a563ba;
  wire v3757ec8;
  wire v3a6f782;
  wire v3753f37;
  wire v37375bc;
  wire v3a70b9e;
  wire v3a615c8;
  wire v3a5f4b8;
  wire v3a6eaef;
  wire v3a7124c;
  wire v373dfff;
  wire v37240a4;
  wire v3751c68;
  wire v372fe10;
  wire v3a6ef42;
  wire v375ab17;
  wire v3a6f3a3;
  wire v374ec22;
  wire v3a70f14;
  wire v372e30c;
  wire v3a70212;
  wire v377e51b;
  wire v375ac09;
  wire v3776767;
  wire v3757cd1;
  wire v376d8fd;
  wire v374089d;
  wire v3a70099;
  wire v3a56f9d;
  wire v3749bc0;
  wire v376f8ea;
  wire v3734e0b;
  wire v1e37915;
  wire v3a69529;
  wire v3a5c779;
  wire v372a20f;
  wire v374fa21;
  wire v1e38305;
  wire v37463bc;
  wire v3732949;
  wire v3a6b405;
  wire v376a3ca;
  wire v3738d43;
  wire v3a66088;
  wire v372ec32;
  wire v1e37e82;
  wire v373583d;
  wire v375cde6;
  wire v3752f21;
  wire v375034b;
  wire v3737423;
  wire v3a70507;
  wire v3770fa1;
  wire v3a6f726;
  wire v3724325;
  wire v3738270;
  wire v3a71674;
  wire v3745239;
  wire v374de25;
  wire v3779003;
  wire v3a6f2fd;
  wire v3739e0e;
  wire v3a53dfc;
  wire v92aebd;
  wire v376c712;
  wire v375cd3f;
  wire v377a36e;
  wire v3a5b5c4;
  wire v37229c2;
  wire v377038e;
  wire v372f74f;
  wire v3a6fb7a;
  wire v3a679ae;
  wire v3767121;
  wire v3764219;
  wire v37235ee;
  wire v3a6a489;
  wire v3a706f1;
  wire v37605e6;
  wire v3779f67;
  wire v3a6324b;
  wire v377f46d;
  wire v3753097;
  wire v3740490;
  wire v372e91a;
  wire v3a67118;
  wire v37367f1;
  wire v3737d38;
  wire v3a6d040;
  wire v3a6fc48;
  wire v3a58a39;
  wire v3775179;
  wire v37767e6;
  wire v3a6bdaa;
  wire v3a61ce7;
  wire v374fb8d;
  wire v3764f27;
  wire v3a6a880;
  wire v373481c;
  wire v3a6fcc8;
  wire v3a56e7a;
  wire v3752eda;
  wire v3725578;
  wire v374f6f9;
  wire v376204f;
  wire v3746496;
  wire v3a6f387;
  wire v2092a9a;
  wire v377dfbf;
  wire v376d979;
  wire v3a6f122;
  wire v3a70134;
  wire v374704d;
  wire v376e2ac;
  wire v3a6ff67;
  wire v375a38b;
  wire v377a7e9;
  wire v372c546;
  wire v3a658c0;
  wire v37577d7;
  wire v375e973;
  wire v3a6f1e4;
  wire v3a703b1;
  wire v372cdef;
  wire v3a64879;
  wire v3a70f30;
  wire v373823e;
  wire v3a6f30a;
  wire v373a0e2;
  wire v3729f32;
  wire v374df1b;
  wire v3762f51;
  wire v372f326;
  wire v3725a21;
  wire v372404f;
  wire v3736b43;
  wire v3735236;
  wire v372bcf2;
  wire v3a6eab2;
  wire v372beb6;
  wire v3a71361;
  wire v37593cb;
  wire v3a57ce9;
  wire v377a51b;
  wire v374f691;
  wire v3a299cd;
  wire v3a661d0;
  wire v372cace;
  wire v3a6d89d;
  wire v3a6f680;
  wire v38079c2;
  wire v374b9ee;
  wire v37307d4;
  wire v3a70902;
  wire v3776f8c;
  wire v3a5bfe6;
  wire v37549e2;
  wire v3741627;
  wire v373a0db;
  wire v3a6efc8;
  wire v372eab1;
  wire v373e74b;
  wire v3a7039a;
  wire v37291e7;
  wire v3737b54;
  wire v3765b77;
  wire v3a661f8;
  wire v3a71353;
  wire v3779cc0;
  wire v3723c3f;
  wire v3a6f896;
  wire v37554b1;
  wire v37643e6;
  wire v3a6eee8;
  wire v3a6f1c1;
  wire v3a64d7c;
  wire v3a60195;
  wire v373c9c1;
  wire v3764805;
  wire v3a70695;
  wire v3a5f5dd;
  wire v373a41e;
  wire v3766a69;
  wire v372c353;
  wire v3a675b2;
  wire v3762ec5;
  wire v37525e0;
  wire v37299d5;
  wire v373ce66;
  wire v37573d2;
  wire v377a65c;
  wire v3a70239;
  wire v3a625ee;
  wire v3769ae2;
  wire v37419a9;
  wire v3730627;
  wire v37311fa;
  wire v3a6f63a;
  wire v3747280;
  wire v37664f6;
  wire v374f96e;
  wire v3742121;
  wire v2092b2c;
  wire v3a5e7bf;
  wire v37654bc;
  wire v37755b2;
  wire v37505a2;
  wire v992750;
  wire v37385fc;
  wire v375a135;
  wire v373453a;
  wire v37574f8;
  wire v3772698;
  wire v3a6de90;
  wire v3a538b4;
  wire v376999f;
  wire v373e91a;
  wire v3a61dca;
  wire v3772dd2;
  wire v3a571de;
  wire v8d3fe3;
  wire v3740923;
  wire v3738e45;
  wire v373e877;
  wire v37570f8;
  wire v37652a5;
  wire v3724af9;
  wire v3a5d8bc;
  wire v3748b15;
  wire v373d49c;
  wire v3724204;
  wire v3757a88;
  wire v3725e0d;
  wire v3a65e6a;
  wire v3a5575e;
  wire v3a6fc5c;
  wire v3a5c75a;
  wire v373d5e7;
  wire v3a70623;
  wire v37784a9;
  wire v374f106;
  wire v3750178;
  wire v3736fc4;
  wire v3726f10;
  wire v3a6fd3e;
  wire v377437d;
  wire v3726826;
  wire v37582c2;
  wire v3a5455e;
  wire v3a71050;
  wire v3807550;
  wire v3a6d80d;
  wire v3a6fc81;
  wire v3752e80;
  wire v3a6fde8;
  wire v3a5980d;
  wire v374b57c;
  wire v3a6ebbc;
  wire v3a6a261;
  wire v3734982;
  wire v37533ae;
  wire v3a5efb2;
  wire v3a6bf6d;
  wire v3a6fff0;
  wire v3746b6e;
  wire v3a70635;
  wire v3732c72;
  wire v3a6e93d;
  wire v3745c84;
  wire v3725932;
  wire v374d751;
  wire v3a6fdc7;
  wire v37c006d;
  wire v372689b;
  wire v373ff4a;
  wire v3725ba8;
  wire v3a69796;
  wire v375c621;
  wire v375b97a;
  wire v3735974;
  wire v373285d;
  wire v377730a;
  wire v376c198;
  wire v3a6c179;
  wire v3770f76;
  wire v9fc6a0;
  wire v375d78f;
  wire v375682e;
  wire v3778176;
  wire v3a55d66;
  wire v3747892;
  wire v37519a8;
  wire v3757b0f;
  wire v374aab3;
  wire v3723dc3;
  wire v376fa43;
  wire v373af15;
  wire v3767a08;
  wire v3762802;
  wire v37649ab;
  wire v3776751;
  wire v372e6a1;
  wire v3768ba1;
  wire v375a023;
  wire v3743393;
  wire v373aeb3;
  wire v3a6f90a;
  wire v374a86a;
  wire v3755417;
  wire v3a6fdea;
  wire v376ce06;
  wire v3724f4f;
  wire v37676dc;
  wire v377152e;
  wire v37232bd;
  wire bdc54c;
  wire v2092f59;
  wire v374bcac;
  wire v3a6c55a;
  wire v3a6f0d1;
  wire v376e3d3;
  wire v3733b0c;
  wire v3744cb5;
  wire v3756cb8;
  wire v3a676aa;
  wire v3a6498e;
  wire v3577318;
  wire v3a71333;
  wire v3a5b03b;
  wire v3767830;
  wire v3a61c41;
  wire v3724418;
  wire v374f0e7;
  wire v375df77;
  wire v37386da;
  wire v3a5b27f;
  wire v3a5ddea;
  wire v372c1cf;
  wire v3a64969;
  wire v3739ac1;
  wire v37256d2;
  wire v39ea7a8;
  wire v3735eb8;
  wire v3a67261;
  wire v3a6784d;
  wire v373a303;
  wire v3a6ef24;
  wire v3a6614b;
  wire v372c91d;
  wire v376856b;
  wire v372c638;
  wire v374dc6d;
  wire v37425a0;
  wire v37343dc;
  wire v3747a97;
  wire v3768f0c;
  wire v37281fb;
  wire v37532ee;
  wire v3a65d93;
  wire v3758466;
  wire v3a70ca5;
  wire v3748360;
  wire v3a674b3;
  wire v377a2f3;
  wire v372fa9d;
  wire v3777527;
  wire v3773098;
  wire v373064e;
  wire v3762ea7;
  wire v37572d0;
  wire v374a0ac;
  wire v3a6fc5d;
  wire v3809fbb;
  wire v3778ecc;
  wire v380a170;
  wire v3a6f00d;
  wire v3763a29;
  wire b1f7c8;
  wire v3a63d55;
  wire v3757da6;
  wire v37504f9;
  wire v3761136;
  wire v3a706a0;
  wire v372d19a;
  wire v374b6ba;
  wire v377926d;
  wire v3778aa6;
  wire v3a70fa3;
  wire v3a70c52;
  wire v3a5d46c;
  wire v3a5f744;
  wire v3774e41;
  wire v3a6a998;
  wire v377816f;
  wire v3a5a6cc;
  wire v373fd58;
  wire v37571fc;
  wire v377053a;
  wire v373ba93;
  wire v375e29c;
  wire v3a7003d;
  wire v3a7008a;
  wire v3745c20;
  wire v374fa2a;
  wire v377455b;
  wire v374f12c;
  wire v37250af;
  wire d1331f;
  wire v3a6757a;
  wire v376b0e6;
  wire v3a6efaa;
  wire v3731688;
  wire v37249f1;
  wire v373fbca;
  wire v3a6f3bb;
  wire v3757966;
  wire v3724579;
  wire v377b690;
  wire v372bdef;
  wire v3771720;
  wire v377320f;
  wire v375adaa;
  wire v3a6f3af;
  wire v3a6f2af;
  wire v37400aa;
  wire v3761071;
  wire v3759e9d;
  wire v3a6ec0d;
  wire v3758ef5;
  wire v373b31d;
  wire v375ed5a;
  wire v3770651;
  wire v2ff8e00;
  wire v372d10e;
  wire v37480f1;
  wire v37617dd;
  wire v377843d;
  wire v372f478;
  wire v37547c9;
  wire v374a5a9;
  wire v3764ba8;
  wire v376bbe8;
  wire v372c6fb;
  wire v3a5affd;
  wire v3754940;
  wire v377e698;
  wire v3775688;
  wire v3a57672;
  wire v3742cd5;
  wire v374c288;
  wire v3727e56;
  wire v377894f;
  wire v377119f;
  wire v3a6f8c1;
  wire v372f576;
  wire v3a70b0d;
  wire v3735580;
  wire v3766d04;
  wire v3725678;
  wire v35b7769;
  wire v3a6ecf6;
  wire v37761fe;
  wire v3a56da3;
  wire v3a5c4e8;
  wire v37242cb;
  wire v373198c;
  wire v3a6e884;
  wire v3741ea8;
  wire v374e078;
  wire v8a1014;
  wire v3767885;
  wire v374c1c3;
  wire v3a693bf;
  wire v3a711f1;
  wire v375c5a1;
  wire v376a6d7;
  wire v37488ed;
  wire v3769f95;
  wire v3a5ef37;
  wire v37452d5;
  wire v3738910;
  wire v374ff5a;
  wire v3760453;
  wire v374b522;
  wire v3a6f4a4;
  wire v376b035;
  wire v3761781;
  wire v3756416;
  wire v373c924;
  wire v3766b11;
  wire v372a711;
  wire v8c890d;
  wire v3747c0b;
  wire v376ee7c;
  wire v3769cd7;
  wire v373f42d;
  wire v375d17c;
  wire v3752d9f;
  wire v3730c49;
  wire v3737f16;
  wire v373eb05;
  wire v373be4d;
  wire v376dd91;
  wire v3a5f8b6;
  wire v376d9ad;
  wire v376b5ac;
  wire v3809e5c;
  wire v3a66aa4;
  wire v37351bc;
  wire v372c3df;
  wire v377d19f;
  wire v37381af;
  wire v372b386;
  wire v35b774b;
  wire v372e93d;
  wire v377c2ac;
  wire v375ff95;
  wire v3a6f213;
  wire v3773b18;
  wire v3a70620;
  wire v37727f9;
  wire v3a70618;
  wire v374174c;
  wire v373b80b;
  wire v3a6fe0d;
  wire v3a540f3;
  wire v3754ec1;
  wire v3756de7;
  wire v3a6e127;
  wire v37255a2;
  wire v3a6f909;
  wire v37656ec;
  wire v373c755;
  wire v3a6f574;
  wire v3774109;
  wire v3a6fe1a;
  wire v3728202;
  wire v3a707b1;
  wire v3772cc3;
  wire v3a57f64;
  wire v3a62c37;
  wire v3774ad3;
  wire v3a662f7;
  wire v37282cf;
  wire v3728608;
  wire v37728d0;
  wire v3a5e817;
  wire v373b599;
  wire v3a6fccc;
  wire v3a66b8a;
  wire cc809f;
  wire v9230c3;
  wire v37c0382;
  wire v3a6f5a5;
  wire v3a6a6c6;
  wire v373e924;
  wire v89df94;
  wire v374a9cd;
  wire v373ed37;
  wire v3a711b7;
  wire v373997b;
  wire v37270d9;
  wire v37686af;
  wire v3752a45;
  wire v37738fc;
  wire v3a6773a;
  wire v3760512;
  wire v37578d4;
  wire v3775750;
  wire v3a710c3;
  wire v3740d05;
  wire v3750e23;
  wire v373badc;
  wire d3af9c;
  wire v3763191;
  wire v3a58d68;
  wire v38093c2;
  wire v3744d99;
  wire v3a70100;
  wire v37242b9;
  wire v373e712;
  wire d58c24;
  wire v373f691;
  wire v372e550;
  wire v3a66ba8;
  wire v3a71424;
  wire v3a6143b;
  wire v375bc4b;
  wire v3a6254e;
  wire v39a4ca8;
  wire v3a55cd6;
  wire v3a70ec7;
  wire v377abd6;
  wire v3a6fdc9;
  wire v3a6bc9a;
  wire v3a69f0e;
  wire v3742d95;
  wire d68a4d;
  wire v376b2e9;
  wire v37274c2;
  wire v3a610a4;
  wire v3a62ccf;
  wire v376da3f;
  wire v3a70a3a;
  wire v377cb41;
  wire v2acb0ef;
  wire v37374e5;
  wire v3a6ef38;
  wire v3738b4c;
  wire v3778484;
  wire v3a62a14;
  wire v3a6eb8f;
  wire v372f046;
  wire v373fa8c;
  wire v372a4e5;
  wire v3766852;
  wire v376dad0;
  wire v3745e0d;
  wire v3a69239;
  wire v374fd1f;
  wire v3730617;
  wire v3808cf5;
  wire v3737ab4;
  wire v376abd1;
  wire v3a701ac;
  wire v372bf1d;
  wire v3a65a52;
  wire v3766048;
  wire v3741c3d;
  wire v377435f;
  wire v35b776e;
  wire v37605a5;
  wire v3a6b161;
  wire v375b61a;
  wire v3776196;
  wire v3a5c5e5;
  wire v374b4ef;
  wire v3a5a307;
  wire v372bb82;
  wire v376848c;
  wire v3732d8f;
  wire v3a623cb;
  wire v376fbfe;
  wire v3a64320;
  wire v380a189;
  wire v3a7027a;
  wire v3778901;
  wire v3736320;
  wire v37362fd;
  wire v37642fa;
  wire v372b1ed;
  wire v3745069;
  wire v3766cd5;
  wire v3a5749f;
  wire v3a68697;
  wire v3770bc0;
  wire v3a6c610;
  wire da7312;
  wire v373e5e7;
  wire v3a713e8;
  wire v37384cb;
  wire v3a6f626;
  wire v377e896;
  wire v373fe1f;
  wire v37313e4;
  wire v377e9c9;
  wire v3739b18;
  wire v3a6f22a;
  wire v3a5dec3;
  wire v3a67f12;
  wire cae8ef;
  wire v3a6f769;
  wire v3a6f01d;
  wire v3739514;
  wire v3a71608;
  wire v377c2ff;
  wire v375e04e;
  wire v3a6f692;
  wire v3763f30;
  wire v3768ed2;
  wire v3760a6e;
  wire v373dee0;
  wire v373cf73;
  wire v3731ab1;
  wire v374e55f;
  wire v373f9bf;
  wire v375e8d9;
  wire v3a6f20c;
  wire v3776fb8;
  wire v37284f3;
  wire v3a71082;
  wire v3a67c34;
  wire v3747212;
  wire v372a0ed;
  wire v373d5af;
  wire v37429cc;
  wire v3736b55;
  wire v3767baa;
  wire v3a60e78;
  wire v3757231;
  wire v37434b2;
  wire v37642e6;
  wire v3a561f0;
  wire v375b0cd;
  wire v3762153;
  wire v37670dd;
  wire v3739368;
  wire v376702c;
  wire v374ae4e;
  wire v3746138;
  wire v3a558be;
  wire v3770071;
  wire v3a71530;
  wire v377a8c3;
  wire v3779470;
  wire v377aae4;
  wire v372f1e9;
  wire v3756dd6;
  wire v372a0a1;
  wire v3a674e2;
  wire v37578f3;
  wire v3763cfa;
  wire v374f95d;
  wire v3734b80;
  wire v3a6f89d;
  wire v3728d84;
  wire v3761cd3;
  wire v3766485;
  wire v3771137;
  wire v3a6efdd;
  wire v3740655;
  wire v372ffd2;
  wire v3741d2d;
  wire v374d260;
  wire v377de41;
  wire v375f077;
  wire v3a61310;
  wire v3727a6c;
  wire v3a711f0;
  wire v3773a9d;
  wire v3729513;
  wire v374e6ec;
  wire v3769c2e;
  wire v375a234;
  wire v3a64c10;
  wire v3734256;
  wire v3751f28;
  wire v3a69ada;
  wire v3732515;
  wire v3a6827b;
  wire v3a5bf5f;
  wire v3749001;
  wire v3735f25;
  wire v3a69ed9;
  wire v374a192;
  wire v3a70fdf;
  wire v3736f2a;
  wire v3a557b1;
  wire v3744590;
  wire v374f617;
  wire v3722b74;
  wire v39a536d;
  wire v3a5f9f2;
  wire v375f74a;
  wire v3a7069e;
  wire v3a6e9b1;
  wire v375dbc6;
  wire v3757082;
  wire v3775a84;
  wire v3752511;
  wire v3a5d90a;
  wire v37419fd;
  wire v1e3780f;
  wire v372a786;
  wire v3a5d6a6;
  wire v3a700ac;
  wire v372610a;
  wire v3766b95;
  wire v3a70097;
  wire v3738dc0;
  wire v3a7132e;
  wire v375faac;
  wire v375d15c;
  wire v3a6f08d;
  wire v373cada;
  wire v3755ad0;
  wire v372e096;
  wire v3774f3b;
  wire v3a7048e;
  wire v37503ec;
  wire v3a63f27;
  wire v3759b6f;
  wire v377bd97;
  wire v373acce;
  wire dbdbc5;
  wire v375c7f8;
  wire c17897;
  wire v3779dae;
  wire v375a288;
  wire v377c186;
  wire bbbe50;
  wire v374b383;
  wire v3a6e8fa;
  wire v3724ee0;
  wire v3a5bded;
  wire v377dfe2;
  wire v372eecf;
  wire v37576d1;
  wire v3a71138;
  wire v3a56f9f;
  wire v3a5fe9e;
  wire v37317f2;
  wire v3741c4b;
  wire v3730895;
  wire v3a6f5e6;
  wire v3a6fb49;
  wire v3778a4f;
  wire v372a9a5;
  wire v37390d5;
  wire v3771a62;
  wire v376ea59;
  wire v3a6fb40;
  wire v373040b;
  wire v3a5fc33;
  wire v37728b9;
  wire v3a6f792;
  wire v3768343;
  wire v3a70264;
  wire v3a66835;
  wire v37534da;
  wire v3a62322;
  wire v37c1a73;
  wire v3731fab;
  wire v3755502;
  wire v374eb3b;
  wire v3a71415;
  wire v37676d0;
  wire v37286d3;
  wire v39eb5ab;
  wire v37462e3;
  wire v375d877;
  wire v372f73c;
  wire v374a4ea;
  wire v3a5e221;
  wire v376df43;
  wire v3723e5f;
  wire v372f6a1;
  wire v3a671f4;
  wire v3a6885a;
  wire v3a568f7;
  wire v3a63af6;
  wire c60044;
  wire v3a69515;
  wire v373aea0;
  wire v1e37bab;
  wire v3806818;
  wire v3a5df97;
  wire v3a712f0;
  wire v373c6a2;
  wire v373d506;
  wire v373342f;
  wire v373b5b8;
  wire v37667f9;
  wire v373df3d;
  wire v3a58554;
  wire v3722f10;
  wire v3a715a7;
  wire v3a67d2f;
  wire v375d7fc;
  wire v3768f7f;
  wire v3a69430;
  wire v3a6feb3;
  wire v38097f6;
  wire v376648e;
  wire v37433ff;
  wire v3755785;
  wire v23fe098;
  wire v373e09b;
  wire v3a5c2df;
  wire v373c768;
  wire v375f9ec;
  wire v3a6f05e;
  wire v37580d5;
  wire v375c910;
  wire v3a7025d;
  wire v3a57bb0;
  wire v376730e;
  wire v3a5e7c0;
  wire v3a5fa25;
  wire v3723747;
  wire v3765b28;
  wire v375e8a2;
  wire v3a66671;
  wire v377a039;
  wire v3a5757f;
  wire v37463e5;
  wire v3807ac6;
  wire v37375f3;
  wire v3a5cf78;
  wire v3a6f3fb;
  wire v377df9c;
  wire v3a5bcf5;
  wire v37586d3;
  wire v3a5d6aa;
  wire v373c8d0;
  wire v3738e72;
  wire v377586c;
  wire v374a0c5;
  wire v3a61753;
  wire c0990a;
  wire v3a672cb;
  wire v3761866;
  wire v3a61acf;
  wire v375685b;
  wire v3775d1d;
  wire v37781ac;
  wire v37647aa;
  wire v37673dd;
  wire v3a6fd27;
  wire v373df71;
  wire v3a69671;
  wire v3764d17;
  wire v3a5996e;
  wire v3762cff;
  wire v3a6ff43;
  wire v3753cc4;
  wire v3a6d525;
  wire v375591f;
  wire v372f4f1;
  wire v3771d2d;
  wire v3727638;
  wire v3731bcf;
  wire v3a6c0e4;
  wire v3a67d59;
  wire v37643eb;
  wire v372b388;
  wire v3a6fb86;
  wire v374916a;
  wire v3a65752;
  wire v3a70616;
  wire v2619aa5;
  wire v3a70fa8;
  wire v3a63812;
  wire v3a6f19d;
  wire v3722b5c;
  wire v375d577;
  wire v3a70cf6;
  wire v3a6f629;
  wire v374b873;
  wire v3744a56;
  wire v3737c04;
  wire v3a702ef;
  wire v376beb3;
  wire v373531a;
  wire v3765798;
  wire v37345e9;
  wire v373fff3;
  wire v3a6eac1;
  wire v3747552;
  wire v3a62a51;
  wire v3a55785;
  wire v3a70bf2;
  wire v3775f0b;
  wire v374c9e9;
  wire v3724a6d;
  wire v3a7036b;
  wire v3768c19;
  wire v37419d7;
  wire v3727de3;
  wire v372826c;
  wire v3a67880;
  wire v3769617;
  wire v3773613;
  wire v3a627a8;
  wire v37418b3;
  wire v3744982;
  wire v37681fa;
  wire v3a576c0;
  wire v3774200;
  wire v3a7103c;
  wire v3a5e9a3;
  wire v3a7092a;
  wire v3a65f15;
  wire v39eb57c;
  wire v3a6f48b;
  wire v37777ad;
  wire v37277a5;
  wire v1e3778d;
  wire v374893c;
  wire v374cfd9;
  wire v3a70010;
  wire v37721e6;
  wire v372cc25;
  wire v3a711ec;
  wire v373d2e3;
  wire v3a5ee85;
  wire v37264a2;
  wire v3a70089;
  wire v35b9d52;
  wire v3738eb6;
  wire v376887c;
  wire v3a6fdb4;
  wire v1e37a34;
  wire v3a5ef0c;
  wire v3733ea2;
  wire v3763f8b;
  wire v377d408;
  wire v372ade8;
  wire v3755c31;
  wire v3763fdf;
  wire v37749b7;
  wire v37c011c;
  wire v3761224;
  wire v3a65f1f;
  wire v373d357;
  wire v3a6fd79;
  wire v3769df4;
  wire v37568c8;
  wire v3a6557d;
  wire v3a5c5ca;
  wire v3754a27;
  wire v3760f62;
  wire v3730aaf;
  wire v377a88e;
  wire v373b98a;
  wire v372b7a5;
  wire v3a6cb5b;
  wire v374f8a1;
  wire v375fa66;
  wire v3735436;
  wire v37697e2;
  wire v373edc8;
  wire v3a55039;
  wire v37740e0;
  wire v37708f1;
  wire v377d2e7;
  wire v377d770;
  wire b62916;
  wire v3a6ff46;
  wire v376d9f8;
  wire v3a5c687;
  wire v377e090;
  wire v3a6e3d1;
  wire v3756925;
  wire v3a6f3ec;
  wire v3765a69;
  wire v3a6797d;
  wire v3a6faab;
  wire v3a6bd5a;
  wire v3a5e776;
  wire v3a68c63;
  wire v377bb93;
  wire v3a6f039;
  wire v3a6b0a1;
  wire v37258d0;
  wire v3a6c127;
  wire v3a70d60;
  wire v37443e0;
  wire v372ed93;
  wire v3739ed3;
  wire v374d12f;
  wire v37548be;
  wire v375a71d;
  wire v375b752;
  wire v3768adf;
  wire v3759e3c;
  wire v3a690c2;
  wire v377957a;
  wire b1feb1;
  wire v2acaff1;
  wire v3762f6e;
  wire cb0c12;
  wire v3742132;
  wire v3a6b89e;
  wire v3a7053b;
  wire v37462ed;
  wire v35b7805;
  wire v3741608;
  wire v3744751;
  wire v3730fb9;
  wire v3a5d6f9;
  wire v373ec72;
  wire c29340;
  wire v3777deb;
  wire v39ebae8;
  wire v3a6f66a;
  wire v377e033;
  wire v3a6f050;
  wire v3a57012;
  wire v375ec4e;
  wire v372f93c;
  wire cceefd;
  wire v377209b;
  wire v3a55861;
  wire v3a6267a;
  wire v374ae67;
  wire v3755898;
  wire v3a62ef1;
  wire v3753445;
  wire v376062b;
  wire v3a710d1;
  wire v3760912;
  wire v3a6f5df;
  wire v3a57584;
  wire v37773c4;
  wire v3a6f32f;
  wire v3763055;
  wire v373f47b;
  wire v1e38291;
  wire v372fca8;
  wire v3a7101b;
  wire v3730e75;
  wire v3a59431;
  wire v3731977;
  wire v3723c25;
  wire v3763793;
  wire v3a5952d;
  wire v3728fd0;
  wire v3a70f33;
  wire v375ef7b;
  wire v37585e6;
  wire v3a707c4;
  wire v3a6f84c;
  wire v374d8c9;
  wire v375e8d2;
  wire v3a299ba;
  wire v3a70a44;
  wire v37415ea;
  wire v38073d4;
  wire v372b982;
  wire v377a7d7;
  wire v372b24d;
  wire v37764d7;
  wire v3a5968c;
  wire v3a6d749;
  wire v3a5614c;
  wire v373f1a5;
  wire v3726d7a;
  wire v3a67e64;
  wire v3734f9f;
  wire v3746fce;
  wire v3726791;
  wire v373fa24;
  wire v3a707d5;
  wire v3a713c9;
  wire v3a71381;
  wire v3759a21;
  wire v3a66a6e;
  wire v3a63172;
  wire v376ce37;
  wire v3a71689;
  wire v3a577f2;
  wire v3a687ea;
  wire v3758539;
  wire v377f34a;
  wire a33229;
  wire v376cebe;
  wire v3a706ce;
  wire v3a6431f;
  wire v3772827;
  wire v3a613f4;
  wire v3a70a6d;
  wire v3a6b97b;
  wire v373a696;
  wire v374f9f5;
  wire v3a70d66;
  wire v3a6e4cd;
  wire v3a6ef30;
  wire v3a6c1d3;
  wire v3769ca2;
  wire v37661dc;
  wire v375e183;
  wire v3a705b2;
  wire v3772007;
  wire v372b798;
  wire v375e167;
  wire v376ad8c;
  wire v374039d;
  wire v3742034;
  wire v3759dda;
  wire v374bf36;
  wire v375eefe;
  wire v373e0b1;
  wire v3732eaa;
  wire v3a70af6;
  wire v3737928;
  wire v1e37a35;
  wire v373de18;
  wire v3a5b23c;
  wire v3a684ee;
  wire v3a61b13;
  wire v3a29856;
  wire v3733412;
  wire v3a587f6;
  wire v3a7007e;
  wire v3a714ef;
  wire v3756471;
  wire v377ebc9;
  wire v372b313;
  wire v37275f8;
  wire v3a6ff62;
  wire v3759664;
  wire v3a70680;
  wire v3a6f3d6;
  wire v374b4d6;
  wire v2093127;
  wire v372a406;
  wire v3724e98;
  wire v3779412;
  wire v3a71659;
  wire v3726c8e;
  wire v2093069;
  wire v3757047;
  wire v35b6167;
  wire v3a6a8c5;
  wire v375feb1;
  wire v9a07a5;
  wire v376513c;
  wire v377ea20;
  wire v3a69203;
  wire v3775ee8;
  wire v3a626ea;
  wire v3a6fa36;
  wire v3761587;
  wire v3a6bb45;
  wire v37526a5;
  wire v3739904;
  wire v37627ec;
  wire v373357d;
  wire v3a7145e;
  wire v377ba29;
  wire v375b84e;
  wire v3a7168c;
  wire v3749f49;
  wire v3a6fea3;
  wire v3a6f581;
  wire v374a23a;
  wire v372a5fc;
  wire v375dbf3;
  wire v3766b94;
  wire v3732b3c;
  wire d3482c;
  wire v3a6f4cc;
  wire v3a5e755;
  wire v376cb9d;
  wire v3766126;
  wire v3739e0d;
  wire v3752a05;
  wire v37711cd;
  wire v376079a;
  wire v372a64f;
  wire v3a71031;
  wire v3a69957;
  wire v3a629fb;
  wire v3a64c32;
  wire v3a5ecb9;
  wire v373fc52;
  wire adaeff;
  wire v3a6d198;
  wire v958697;
  wire v3742441;
  wire v3a68391;
  wire v37346c5;
  wire v8455df;
  wire v31c329f;
  wire v3a6521e;
  wire v39378d6;
  wire v3a58b3f;
  wire v375c50a;
  wire v3776eff;
  wire v3730a6a;
  wire v376858c;
  wire v377b221;
  wire v3a70945;
  wire v3937409;
  wire v3793188;
  wire v3730712;
  wire v3725872;
  wire v3751a4f;
  wire v372cd7e;
  wire v379318f;
  wire v3766e62;
  wire v37772c0;
  wire v373e8e3;
  wire v3a6fe4a;
  wire v3a29814;
  wire v37788d5;
  wire v3a55aa3;
  wire v374d781;
  wire v3752e29;
  wire v375c7cd;
  wire v374a39f;
  wire v3806a7a;
  wire v3773165;
  wire v377065f;
  wire v9684f8;
  wire v375571d;
  wire v3751369;
  wire v377a975;
  wire v373172e;
  wire v3773c62;
  wire v3727eda;
  wire v3760a58;
  wire v372ee4b;
  wire v3a7093d;
  wire v3729555;
  wire v372dbe1;
  wire v3a6fbc2;
  wire v374bd13;
  wire v3739d49;
  wire v377e0c6;
  wire v3a6acd3;
  wire v38076b7;
  wire v37726d9;
  wire v3a6f1ef;
  wire v3a680cd;
  wire v3741920;
  wire v3a5cae1;
  wire v375c525;
  wire v372a25a;
  wire v375e9c0;
  wire v374e692;
  wire bc8871;
  wire v37260fc;
  wire v37261b3;
  wire v372a958;
  wire v3a558c2;
  wire v3a705d7;
  wire v8f695f;
  wire v3770fb7;
  wire c7ba89;
  wire v3a63f55;
  wire v3746f89;
  wire v372cf41;
  wire v375efe8;
  wire v375ace5;
  wire v376d766;
  wire v372aff0;
  wire v3a70ca8;
  wire v3763c04;
  wire v373abe2;
  wire v375e2ab;
  wire v372adb5;
  wire v372bc50;
  wire v3a70a25;
  wire v37395d4;
  wire v377d999;
  wire v3a57796;
  wire v372fe64;
  wire v3778354;
  wire v3a6d098;
  wire v3a707ee;
  wire v3a702f0;
  wire v375722a;
  wire v3a6adb8;
  wire v373bb89;
  wire v3733b4b;
  wire v3a6a332;
  wire v3a64288;
  wire v3a70f15;
  wire v374ab76;
  wire v374de47;
  wire v3a70cd0;
  wire v3757fdd;
  wire v8686c3;
  wire v3a6f619;
  wire v3a618f6;
  wire v37550ac;
  wire v3759ff9;
  wire v374aa67;
  wire v92a8d7;
  wire v374b40e;
  wire v3a5ff26;
  wire v3a5f60c;
  wire v3a5897a;
  wire v3737411;
  wire v3a6caab;
  wire v3a7141d;
  wire v3723a1d;
  wire v3735f03;
  wire d9fd79;
  wire v3a7039b;
  wire v3731859;
  wire v3726d94;
  wire v373759d;
  wire v8fdd0d;
  wire v373642c;
  wire v3a5a807;
  wire v375ff74;
  wire v376b651;
  wire v3a6efe3;
  wire v374c02e;
  wire v3a572ea;
  wire v3754d67;
  wire v3762199;
  wire v3731376;
  wire v3a54d04;
  wire v373087c;
  wire v3a70760;
  wire v376da21;
  wire v3a70ff2;
  wire v3a6eb4f;
  wire v2ff8e8b;
  wire v3723ac4;
  wire v3a5bb57;
  wire v3a5e874;
  wire v3a6f41f;
  wire v37334c2;
  wire v377a0be;
  wire v3a708ed;
  wire v3732ef8;
  wire v3743c45;
  wire v3727f67;
  wire v374fe7f;
  wire v3a70e06;
  wire v374f593;
  wire v37684ed;
  wire v3a7116b;
  wire v3a6d92f;
  wire v372ac19;
  wire v376f718;
  wire v3a53e5c;
  wire v3a63e51;
  wire v3a65dbb;
  wire v3a55456;
  wire v3a6f70a;
  wire v372e868;
  wire v3a7132d;
  wire v372d905;
  wire v3739faf;
  wire v375ef36;
  wire v377955b;
  wire v3a6f36d;
  wire v372fb3c;
  wire v3723ddc;
  wire v3734b5a;
  wire v3765d05;
  wire v3a6fca0;
  wire v376ac47;
  wire v3722e59;
  wire v372ed79;
  wire v377bde3;
  wire v3771df4;
  wire v3774662;
  wire v3a66b6e;
  wire v37367e3;
  wire v374a650;
  wire v3737700;
  wire v3a6e9fc;
  wire v372aafa;
  wire v3a71342;
  wire v3a6c6c3;
  wire v373c071;
  wire v3a71392;
  wire v3a5397f;
  wire v373da7d;
  wire v375874f;
  wire v3740f25;
  wire v3a6fc84;
  wire v3a66a8e;
  wire v3a7031a;
  wire v377ac0f;
  wire v3734041;
  wire v3a703c9;
  wire v37795eb;
  wire v3a5a8f6;
  wire v3a712b9;
  wire v3a6f7b6;
  wire v372fff7;
  wire v3a6becc;
  wire v3756fd9;
  wire v37395e6;
  wire v37473af;
  wire v373b589;
  wire v3776441;
  wire v3a6fd67;
  wire v372fe58;
  wire v3767f33;
  wire v3a713f0;
  wire v376bcaa;
  wire v375925f;
  wire aab2b0;
  wire v3753a65;
  wire v3757556;
  wire v3a61480;
  wire v376dad4;
  wire v3749139;
  wire v3a5fed1;
  wire v3a6c3ae;
  wire v3777216;
  wire v373c82f;
  wire v3746d89;
  wire v3a54b5d;
  wire v3737a21;
  wire v376c224;
  wire v376fd84;
  wire v37512f6;
  wire v375b278;
  wire v3743ab6;
  wire v376faa6;
  wire v3778395;
  wire v376581d;
  wire v3765978;
  wire v3733dea;
  wire v3738726;
  wire v3a715a4;
  wire v3a63fbc;
  wire v374df88;
  wire v373aa76;
  wire v3a55b91;
  wire v3a65ee0;
  wire v372b034;
  wire v3a6f52a;
  wire v23fe21d;
  wire v37299ef;
  wire v3a6c9c7;
  wire v37742c5;
  wire v373714f;
  wire v3a71286;
  wire v3a6eb5b;
  wire v375534d;
  wire v373755a;
  wire v3a70990;
  wire v3731d06;
  wire v375527f;
  wire v3731f3c;
  wire v3753576;
  wire a2a6f3;
  wire v373346a;
  wire v3a57891;
  wire v375bb11;
  wire v374e7c5;
  wire v3a58732;
  wire v37609d7;
  wire v3734b35;
  wire v3a554a6;
  wire v3741b28;
  wire v376fbcd;
  wire v3a6b6d2;
  wire v372d1a4;
  wire v3744752;
  wire v3a70182;
  wire v3a6432d;
  wire v374d140;
  wire v3774f45;
  wire v376b0fb;
  wire v376563d;
  wire v374bbbf;
  wire v3a70bbc;
  wire v380853c;
  wire v372c4bd;
  wire v3751196;
  wire v3741cda;
  wire v37476f7;
  wire v1e3741b;
  wire v3255a07;
  wire v37569ec;
  wire v376a1a3;
  wire v374c88a;
  wire v3a6f942;
  wire v3a61e33;
  wire v376c611;
  wire v3a6fc57;
  wire v377b8c5;
  wire v3744af7;
  wire v372b29d;
  wire v372c762;
  wire v372e53f;
  wire v374a664;
  wire v3a71688;
  wire v3767a5b;
  wire v37506d8;
  wire v3a594f1;
  wire v372580e;
  wire v3a70b98;
  wire v374c69c;
  wire v3753c8c;
  wire v3a67c6d;
  wire v3a714f8;
  wire v3771214;
  wire v377de72;
  wire v3a70596;
  wire v376e115;
  wire v376226e;
  wire v3733993;
  wire v8db8b7;
  wire v375095a;
  wire v376c1d6;
  wire v3732510;
  wire v373db50;
  wire v3774ae5;
  wire v3a6e09b;
  wire v3a5cc14;
  wire v3777825;
  wire v374f1e9;
  wire v3a6d3b6;
  wire v372b2ab;
  wire v372b780;
  wire v1e37846;
  wire v3a65716;
  wire v377e618;
  wire v376847d;
  wire v3a700f8;
  wire v3738be9;
  wire v372af46;
  wire v375f3bd;
  wire v376218c;
  wire v3a7031d;
  wire v377a6ce;
  wire v372fbf4;
  wire v3727fd0;
  wire v3a70710;
  wire v3736ab1;
  wire v375eb78;
  wire v374270d;
  wire v376bf04;
  wire v373b744;
  wire v3a56396;
  wire v373f8fb;
  wire v3a63197;
  wire v374bee4;
  wire v3809427;
  wire v3a70bfa;
  wire v374b60b;
  wire v3a70d90;
  wire v373b2ce;
  wire v377437f;
  wire v372546e;
  wire v3a5d93f;
  wire v3751cc4;
  wire v92e6f3;
  wire v3a70d3e;
  wire v3773f83;
  wire v37767cd;
  wire v3a5ee62;
  wire v3757024;
  wire v37434f6;
  wire v3747167;
  wire v373ba4a;
  wire v376c017;
  wire v3778a89;
  wire v3a5ff76;
  wire v3809282;
  wire v3744fa5;
  wire v3a710e9;
  wire v37565ae;
  wire v372f192;
  wire v3731a29;
  wire v3774d15;
  wire v3755b54;
  wire v373ec0f;
  wire v3a5e1bc;
  wire v3a70190;
  wire v37741ca;
  wire v37419bc;
  wire v3778492;
  wire v3725931;
  wire v374f4a3;
  wire v3773e34;
  wire v3750c0d;
  wire v3a598a9;
  wire v8615d7;
  wire v3a7108a;
  wire v376fac8;
  wire v37520db;
  wire v374e5ac;
  wire v372923a;
  wire v373621d;
  wire v8cdbc1;
  wire v3733a19;
  wire v3a6f331;
  wire v23fd804;
  wire v2ff91fe;
  wire v372a9c7;
  wire v3722ae9;
  wire v3a6fcc9;
  wire v3773bbc;
  wire v377aa2e;
  wire v3a7106e;
  wire v3a66014;
  wire v3763011;
  wire v3741acc;
  wire v37636e4;
  wire v3752af0;
  wire v3751931;
  wire v377d393;
  wire v3a6fee8;
  wire v3a70351;
  wire v3758b3f;
  wire v3a5a0b3;
  wire v374c4e1;
  wire v3771ee8;
  wire v373dcb0;
  wire v90a00a;
  wire v377e52e;
  wire v3a714e6;
  wire v373d8c0;
  wire ae6485;
  wire v1e37921;
  wire v375f4fd;
  wire v3774a7e;
  wire v3a7062e;
  wire v3a704c0;
  wire v3a699f5;
  wire v375ed9f;
  wire v375bcf2;
  wire v372f2b7;
  wire v3723a00;
  wire v3768c97;
  wire v35b710e;
  wire v373409f;
  wire v3a70e35;
  wire v377a036;
  wire v377a343;
  wire v3777d95;
  wire v3a7138d;
  wire v372c86a;
  wire v372984c;
  wire v3739e25;
  wire v376e844;
  wire v3725580;
  wire v3a6ef00;
  wire v3a6f902;
  wire v3a57b88;
  wire v375e261;
  wire v376096f;
  wire v375d861;
  wire v3725252;
  wire v3a71379;
  wire v3a6b129;
  wire v373a3e4;
  wire v3a5af86;
  wire v3774416;
  wire v360bb9f;
  wire c51df8;
  wire v3736d51;
  wire v3a6f562;
  wire v373c331;
  wire v3a6f8bb;
  wire v373f028;
  wire v3809879;
  wire v3723cc2;
  wire v3a6f110;
  wire v3a6442f;
  wire v373f051;
  wire v37407f5;
  wire v373b46b;
  wire v377c4b7;
  wire v377317d;
  wire v3a6ef7f;
  wire v372dcac;
  wire v377e934;
  wire v3a6830a;
  wire c8ab71;
  wire v376d268;
  wire v374a6ce;
  wire v3730be3;
  wire v374e86a;
  wire v37306ec;
  wire v3762116;
  wire v3a70ecc;
  wire v375cc8b;
  wire v3a6fa33;
  wire v3807587;
  wire v3756943;
  wire v3751f67;
  wire v3a6f5d1;
  wire v3749686;
  wire v3734827;
  wire v37487f5;
  wire v3744dd2;
  wire v3a70568;
  wire v3773a45;
  wire v3a7088d;
  wire v374fc82;
  wire v3764586;
  wire v374d674;
  wire v3a70a41;
  wire v3737d95;
  wire v3a6c8cc;
  wire v3731b72;
  wire v3a5872b;
  wire v37765fb;
  wire v3a68607;
  wire v3738251;
  wire v3741dea;
  wire v3a6826d;
  wire v3766105;
  wire v3743c44;
  wire v375e9a7;
  wire v3a65e1e;
  wire v377a657;
  wire v376151e;
  wire v376cedc;
  wire v375380a;
  wire v3a70c13;
  wire v875999;
  wire v377e5fd;
  wire v376efda;
  wire v3a5b4c1;
  wire v3a6f328;
  wire v3726806;
  wire v37619b8;
  wire v3758f6d;
  wire v3a6f4dc;
  wire v3731389;
  wire c8d28b;
  wire v3a6c004;
  wire v375f6c7;
  wire v3748d55;
  wire v3a70be4;
  wire v3a7074c;
  wire v3a6d3bc;
  wire v375b929;
  wire v3a705e0;
  wire v37655c5;
  wire v3a6fe75;
  wire v3a5a805;
  wire v3a6f4ee;
  wire v37518c9;
  wire v3a706a1;
  wire v3747554;
  wire v374366a;
  wire v3a5dab7;
  wire v3750f1e;
  wire v3a694a5;
  wire v3722f8e;
  wire v3a6764b;
  wire v375c2e2;
  wire v3a6f69c;
  wire v3775630;
  wire v3744b16;
  wire v3747d51;
  wire v3a6f459;
  wire v373a0ea;
  wire v3a625ac;
  wire v3a61be2;
  wire v3a715d7;
  wire v3a675bb;
  wire v374bec2;
  wire v37322a9;
  wire v372771e;
  wire v3a6f1ad;
  wire v3776dcd;
  wire v3747a3f;
  wire v3a67f0c;
  wire v3769245;
  wire v37c00f6;
  wire v3a6c908;
  wire v373d62f;
  wire v3742e25;
  wire v373951e;
  wire v3a60e6d;
  wire v3774882;
  wire v375a563;
  wire cdcddf;
  wire v3a6fab5;
  wire v3a62072;
  wire v373b4ce;
  wire v3a615a2;
  wire v3a70112;
  wire v3731b60;
  wire v3a6cc65;
  wire v377529a;
  wire v3a5fd0a;
  wire v3a576bd;
  wire v373d235;
  wire v3756343;
  wire v3728b47;
  wire v3a6f729;
  wire v377b61e;
  wire v3773804;
  wire d9e2a4;
  wire v3a583cd;
  wire v37507be;
  wire v3776996;
  wire v3a6f918;
  wire v3a64fe0;
  wire v377e08c;
  wire v3745291;
  wire v3744fbb;
  wire v3771656;
  wire v3a6f880;
  wire v3a53a8a;
  wire v3748829;
  wire v3728f66;
  wire v3740da1;
  wire v3a70d59;
  wire v376596c;
  wire v37493c7;
  wire v3a7009f;
  wire v37532a8;
  wire v2acb0c1;
  wire v3726df4;
  wire v3a5ec2d;
  wire v372886c;
  wire v3a57d40;
  wire v3a5a4a0;
  wire v3737053;
  wire v375ecd5;
  wire v3a712d0;
  wire v3733557;
  wire v376d9f3;
  wire v337904a;
  wire v3a5d0d3;
  wire v372d764;
  wire v376c9a5;
  wire v3a6b372;
  wire v3733bed;
  wire v376afb1;
  wire v372e754;
  wire v37379a2;
  wire v3a70713;
  wire v2ff8c78;
  wire v376285a;
  wire v37635de;
  wire v3765927;
  wire v3a62027;
  wire v39eb56d;
  wire v374ba3c;
  wire v3a712a6;
  wire v94ce87;
  wire v3a6958b;
  wire v373dcad;
  wire v3a709e2;
  wire v3769c70;
  wire v3a7143c;
  wire v3739bb2;
  wire v3a6c40f;
  wire v3a700ec;
  wire v37733e3;
  wire v3a60c82;
  wire v3726aa5;
  wire v3a63bb0;
  wire v3765d84;
  wire v3740df7;
  wire v3a5e60c;
  wire v37661b2;
  wire v3a5cc1a;
  wire v376f4b2;
  wire v37439ad;
  wire v3769ad7;
  wire v374b68a;
  wire v377e869;
  wire v3727141;
  wire v3742b88;
  wire v37360c0;
  wire v3a57bd7;
  wire v3a70ea1;
  wire v3a6380f;
  wire v3745458;
  wire v3749a4c;
  wire v3777efb;
  wire v3a6b1b9;
  wire v3758b78;
  wire v3a6f2ba;
  wire v969d5b;
  wire v3a66ad2;
  wire v3736ecc;
  wire v377e6f5;
  wire v373b59f;
  wire v375795d;
  wire v3725b9b;
  wire v3a585d1;
  wire v3a6854c;
  wire v3a712af;
  wire v3733767;
  wire v375859a;
  wire v3732ecb;
  wire v3a5fc05;
  wire v37480ad;
  wire v3a58ca1;
  wire v375f708;
  wire v374b36f;
  wire v3732926;
  wire v377d126;
  wire v3751807;
  wire v37390c5;
  wire v3a71248;
  wire v375585e;
  wire v3a7129d;
  wire v375d102;
  wire v37758d3;
  wire v373db07;
  wire v37353c6;
  wire v3a6f456;
  wire v3a709ea;
  wire v3a5acd9;
  wire v375c939;
  wire v37388ce;
  wire v376093b;
  wire v3a6dcf0;
  wire v377a876;
  wire v372b75b;
  wire v375a08b;
  wire v3757684;
  wire v37670ac;
  wire v3763224;
  wire v2ff9362;
  wire v375c3b0;
  wire v3759158;
  wire v377a2f2;
  wire v377acae;
  wire v37588c4;
  wire v374820d;
  wire v3724a6e;
  wire v23fdeaf;
  wire v3755914;
  wire v375f368;
  wire v3771931;
  wire v3a60301;
  wire v3774df5;
  wire v375e8aa;
  wire v3773c70;
  wire v3a61bac;
  wire v3a63624;
  wire v373822e;
  wire v3a56847;
  wire v374daa9;
  wire v3730829;
  wire v372b8a5;
  wire v37258d6;
  wire v3a6eeb9;
  wire v372a352;
  wire v380714f;
  wire v374ad96;
  wire v3752446;
  wire v3a71505;
  wire v377b48b;
  wire v376d1b3;
  wire v3750e94;
  wire v374be59;
  wire v373fb71;
  wire v37411c6;
  wire v3732bb6;
  wire v37380e2;
  wire v377f61c;
  wire v3739ab2;
  wire v37686c7;
  wire v3a5c998;
  wire v375b5eb;
  wire v3a7043d;
  wire v374fcac;
  wire v3a6fb38;
  wire v3a709d6;
  wire v375041a;
  wire v372b715;
  wire v3a64f1f;
  wire v3806cd2;
  wire v3a6f8af;
  wire v3768a3c;
  wire v91ebb9;
  wire v3a6094a;
  wire v37609a8;
  wire v376b1ad;
  wire v3a67312;
  wire v3740922;
  wire v3748f40;
  wire v3729d65;
  wire v3754450;
  wire v8bc7a8;
  wire v3745717;
  wire v3a707ef;
  wire v3a674c4;
  wire v37788d6;
  wire v3a5b0ea;
  wire v3a5ccab;
  wire v3758e73;
  wire v3a70063;
  wire v3a6f684;
  wire v3746676;
  wire v374c22d;
  wire v377f71d;
  wire d7cff8;
  wire v375d1d0;
  wire v3a5b00a;
  wire v3739bd5;
  wire v373c665;
  wire v376c22c;
  wire v3a6b29f;
  wire v376f542;
  wire v37329e1;
  wire v3760e75;
  wire v3766b05;
  wire v3747e73;
  wire v3725d48;
  wire v3a6924e;
  wire v3a600a8;
  wire v375986d;
  wire v3a6d4cd;
  wire v3728382;
  wire v9f56fd;
  wire v375a025;
  wire v37676e0;
  wire v372766c;
  wire v3a6fa13;
  wire v37236b3;
  wire v372c5a0;
  wire v3765c70;
  wire b3a152;
  wire v374837b;
  wire v374f8a5;
  wire v3a7110f;
  wire v37693ce;
  wire v3a6f96e;
  wire v360d029;
  wire v3762121;
  wire v2092b90;
  wire v3a6f766;
  wire v372775f;
  wire v375a0ed;
  wire v380877d;
  wire v3a61ad3;
  wire v375e52f;
  wire v376f4a6;
  wire v374d03f;
  wire v375b265;
  wire v3729bd7;
  wire v37c101a;
  wire v3806f67;
  wire v37308bf;
  wire v377dcf5;
  wire v3a6b798;
  wire v376230d;
  wire v3a70efb;
  wire v372c702;
  wire v3769cc2;
  wire v3a6422d;
  wire v3a7128e;
  wire v3766014;
  wire v3a6e404;
  wire v372dc35;
  wire v3a6f040;
  wire v3a5e82d;
  wire v3a58d2e;
  wire v377260b;
  wire v372c6b3;
  wire v8f2b25;
  wire v37499c4;
  wire v3734c75;
  wire v3776fae;
  wire v37293c2;
  wire v8455f9;
  wire v3a28da6;
  wire v372c046;
  wire v376a25e;
  wire v37666b4;
  wire v397d860;
  wire v3a6ebf9;
  wire v3728d9c;
  wire v3a70ae5;
  wire v3769f5f;
  wire v3a69727;
  wire v37504fd;
  wire v3a66667;
  wire v3a57aad;
  wire v3a709a4;
  wire v3a71685;
  wire v373e827;
  wire v374be5d;
  wire v372f38e;
  wire v376dea1;
  wire v372e365;
  wire v3a7093a;
  wire v3a5c0d4;
  wire v3a712b1;
  wire v376e3fb;
  wire v374486d;
  wire v375929c;
  wire v3774f56;
  wire v376c4ef;
  wire v3a6c322;
  wire v3a710e0;
  wire v376d45e;
  wire v1e38241;
  wire v3772c7a;
  wire v3a6cd35;
  wire v37781b8;
  wire v3a62b5f;
  wire v377ae32;
  wire v374ec35;
  wire v37796bf;
  wire v3772112;
  wire v3a6843c;
  wire v373c0a8;
  wire v372d411;
  wire v3774175;
  wire v372d83d;
  wire v373d35f;
  wire v373b76d;
  wire v3a6df32;
  wire v3a70375;
  wire v3a67e13;
  wire v3a70863;
  wire v3738a5e;
  wire v3a6fbd8;
  wire v373261f;
  wire v3777ee9;
  wire v377297e;
  wire v3a57c0b;
  wire v3775a29;
  wire v3a5491d;
  wire v3726c8c;
  wire v3738263;
  wire v3748256;
  wire v375d3da;
  wire v376a70f;
  wire v3a65a2e;
  wire v3a6b49a;
  wire v37751b2;
  wire v374a134;
  wire v9450a2;
  wire v3a70987;
  wire v374249f;
  wire v3746d2a;
  wire v373026f;
  wire v376a3aa;
  wire v37751cb;
  wire v3726a38;
  wire v377b3cf;
  wire v374f547;
  wire v3a6f56a;
  wire v3a6b6a3;
  wire v3a5c733;
  wire v375408d;
  wire v3a71524;
  wire v3a70209;
  wire v37771e3;
  wire v3735012;
  wire v3a712ed;
  wire v377a01a;
  wire v38094fb;
  wire v37770ed;
  wire v3776b09;
  wire v3756d53;
  wire v3808d0f;
  wire v3771804;
  wire v3a6e7a4;
  wire v360c3d7;
  wire v372ae9d;
  wire v377fb81;
  wire v376a755;
  wire v377eac3;
  wire v374b65e;
  wire ae317f;
  wire v37327c5;
  wire v377672d;
  wire v37366da;
  wire v3778362;
  wire v3730ba6;
  wire v375fbf2;
  wire v377d76b;
  wire v3a6b916;
  wire v3a71330;
  wire v3a70318;
  wire v372ef17;
  wire v3a5a8a4;
  wire v374d162;
  wire v3a640a0;
  wire v374e0f6;
  wire v3773ee7;
  wire v3768c3e;
  wire v3a6f23a;
  wire v374e4ec;
  wire v3a70556;
  wire v376d4f3;
  wire v3a7022a;
  wire v37556c0;
  wire v37449d1;
  wire v3a6ec10;
  wire v37601df;
  wire v3255a16;
  wire v3739d88;
  wire v374e056;
  wire v3725d73;
  wire v3757c7f;
  wire v375959a;
  wire v3a570f5;
  wire v3722d81;
  wire v37438b9;
  wire v3a70476;
  wire v3a60dfb;
  wire v377b9ab;
  wire v3724db7;
  wire v376a056;
  wire v376142c;
  wire v372383a;
  wire v3a6fb71;
  wire v373f6ee;
  wire v3758cf5;
  wire v3743040;
  wire v375022e;
  wire acc1e3;
  wire v37509a9;
  wire v372e36d;
  wire v373505c;
  wire v3a70d63;
  wire v3731349;
  wire v3740cd2;
  wire v3733998;
  wire v3a58d22;
  wire v3a57325;
  wire v3764978;
  wire v3754d82;
  wire v3a68cc4;
  wire v3a70b1e;
  wire v3a539bf;
  wire v3807183;
  wire v377359f;
  wire v374e542;
  wire v3a6f84a;
  wire v3a58353;
  wire v373325f;
  wire v3a6a2f3;
  wire v377e181;
  wire v3a667e7;
  wire v3a6ebac;
  wire v3a65402;
  wire v3a6f765;
  wire v376af1a;
  wire v377f640;
  wire v3745e0e;
  wire v3a70386;
  wire v3a6c5e5;
  wire v3768048;
  wire v3762f2d;
  wire v3a61a37;
  wire v377be72;
  wire v3a61714;
  wire v373d97a;
  wire v375e961;
  wire v3a6f8a7;
  wire v3a6d874;
  wire v376f271;
  wire v3a70f70;
  wire v375bed5;
  wire v3742fc4;
  wire v3a70025;
  wire v375d9b1;
  wire v376ecc8;
  wire v37389d5;
  wire v3730d1e;
  wire v3a5fe39;
  wire v3a70cda;
  wire v3a6bbc6;
  wire v375dd02;
  wire v3a6e7ce;
  wire v373a755;
  wire v3a6eb6e;
  wire v372def3;
  wire v3a6f91e;
  wire v375331e;
  wire v372a071;
  wire v3a56b7c;
  wire v372bb0f;
  wire v373b7dd;
  wire v375facf;
  wire v37280f3;
  wire v3772200;
  wire v37509fc;
  wire v3a60bae;
  wire v3725470;
  wire v377cd9c;
  wire v3a6cad7;
  wire v3a6fe57;
  wire v37522e8;
  wire v3a6c7f2;
  wire v372f58a;
  wire v3a62079;
  wire v3a700e9;
  wire v375c4ab;
  wire v373651a;
  wire v3a70137;
  wire v374bb9f;
  wire ca095d;
  wire v377c9f3;
  wire v377c4bf;
  wire v375f8b1;
  wire v377e6fc;
  wire v373e944;
  wire v3a6375b;
  wire v3a71124;
  wire v3a6fbad;
  wire v3a70cd6;
  wire v33782fe;
  wire v374e5ab;
  wire v372dd2a;
  wire v374fda1;
  wire v35b987f;
  wire v372b813;
  wire v3737517;
  wire v35b91ba;
  wire v374b86c;
  wire v37366b7;
  wire v377c0fa;
  wire v3751c1c;
  wire v373ff17;
  wire v3765121;
  wire v3749f78;
  wire v3a6efe1;
  wire v377c9bd;
  wire v377700a;
  wire v3a65a0f;
  wire v3a67f49;
  wire v3a61992;
  wire v372757f;
  wire v3a7101d;
  wire v3747f46;
  wire v3735d6f;
  wire v3a6fcb7;
  wire v373518a;
  wire v3a6f44a;
  wire v37341ff;
  wire v3750faa;
  wire v375cf11;
  wire v35b86d1;
  wire v3a6953d;
  wire v3777d7c;
  wire v373264f;
  wire v375c28e;
  wire v376209f;
  wire v37689b5;
  wire v37626cc;
  wire v37c36c4;
  wire v3749f2e;
  wire v375e944;
  wire v37273f6;
  wire v372ec9f;
  wire v377cbf0;
  wire v3751929;
  wire v3a5d6b7;
  wire v373f364;
  wire v3a6879a;
  wire v3a695ec;
  wire dc57c8;
  wire v1e37489;
  wire v3738906;
  wire v375d640;
  wire v3a6ef7d;
  wire v377cb05;
  wire v3a6d926;
  wire v3a715f8;
  wire v3756c19;
  wire v3a6bc32;
  wire v375580b;
  wire v3760ba7;
  wire v373bca5;
  wire v3750a17;
  wire v35b7096;
  wire v373c050;
  wire v3a64624;
  wire v3a713e2;
  wire v373dc11;
  wire v3a715bb;
  wire v3756031;
  wire v3a5de32;
  wire v3731123;
  wire v376a8c8;
  wire v3731549;
  wire v377d256;
  wire v37733c0;
  wire v3a58da1;
  wire v372cda0;
  wire v3a6fb7c;
  wire v3a710f6;
  wire v372be59;
  wire v375a766;
  wire v377af34;
  wire v3741f5e;
  wire v3a6f6d3;
  wire v3745181;
  wire v377ef6e;
  wire v3a53f53;
  wire v373828a;
  wire v372cfad;
  wire v39eb536;
  wire v373f224;
  wire v3755f4a;
  wire v373c8ff;
  wire v37586c0;
  wire v3743f5a;
  wire v372f570;
  wire v374679f;
  wire v37600c0;
  wire v3a6f700;
  wire v3a6f838;
  wire v3a6f7d2;
  wire v37271fd;
  wire v377bdec;
  wire v3733b46;
  wire v37490ae;
  wire v39eb44e;
  wire v3727c1d;
  wire v3a573cc;
  wire v3a6e2d0;
  wire v3a55ecf;
  wire v3a5acca;
  wire v3732939;
  wire v3a59e74;
  wire v3772e46;
  wire v377e71d;
  wire v3a53c50;
  wire v3a6000d;
  wire v3a5e96b;
  wire v3740f5d;
  wire v3a6fe5e;
  wire v377b0a3;
  wire v3a65ae2;
  wire v3750254;
  wire v377ea3c;
  wire v3778ab7;
  wire v376daf2;
  wire v3a713f1;
  wire v1e37daf;
  wire v3751862;
  wire v373b295;
  wire v3a5a04c;
  wire v376ed2b;
  wire v3a706af;
  wire v377ddc1;
  wire v3a67a41;
  wire v3742b6a;
  wire v3760927;
  wire v3a701bc;
  wire v3a5b58e;
  wire v3a69bdc;
  wire v23fde66;
  wire v3a6f773;
  wire v376b94a;
  wire v2acaeee;
  wire v3a6ffdd;
  wire v374f3a9;
  wire v3758e9e;
  wire v3731c79;
  wire v37361e7;
  wire v372ed88;
  wire v3a6e57f;
  wire v3a70453;
  wire v3761333;
  wire v377a653;
  wire cb85ef;
  wire v3a643d6;
  wire v372fe28;
  wire v3a7041c;
  wire v373b717;
  wire v3a5f5f5;
  wire v3722ad4;
  wire v3a61246;
  wire v373a945;
  wire v3a29da0;
  wire v3729cfa;
  wire v373d199;
  wire v3757ca4;
  wire v37b64f8;
  wire v373cd8a;
  wire v37720ce;
  wire v3a6f07f;
  wire v3723add;
  wire v3a6355c;
  wire v37709ec;
  wire v375fcab;
  wire v3724c25;
  wire v377bca1;
  wire v3a652de;
  wire v3750674;
  wire v376a7b5;
  wire v3a7062c;
  wire v377ac4c;
  wire v373c01a;
  wire v37785a8;
  wire v374b894;
  wire b3f461;
  wire v37584c6;
  wire v3a67fea;
  wire v3724784;
  wire v3722d9d;
  wire v3a60cdb;
  wire v3809400;
  wire v3a7045b;
  wire v3a6600c;
  wire v3a6fbdd;
  wire v3a70ac7;
  wire v372aa55;
  wire v3734dd8;
  wire v3a694bb;
  wire v376af2d;
  wire v3a7146f;
  wire v3733343;
  wire v3762d06;
  wire v37651b2;
  wire v3a53f42;
  wire v375b4d8;
  wire v3a5a68d;
  wire v3743da3;
  wire v3a586f1;
  wire v3779f6b;
  wire v377873a;
  wire v3731c72;
  wire v3a55755;
  wire be2682;
  wire v376c490;
  wire d648e4;
  wire v3777c59;
  wire v376c6ba;
  wire v3a5b8b0;
  wire v3a70ca3;
  wire v3748a87;
  wire v3751968;
  wire v375e3d1;
  wire v375946b;
  wire v372d9ad;
  wire v3a6eb1d;
  wire v374f304;
  wire v372992f;
  wire v3a715e3;
  wire v37663b5;
  wire v3a6f09a;
  wire v3768c2a;
  wire v3755bbd;
  wire v3a71563;
  wire v3723e77;
  wire v377970b;
  wire v3a6ef5c;
  wire v3a57106;
  wire v37775ff;
  wire v3735ff7;
  wire v3a5ae8d;
  wire v3a708c1;
  wire v37424b8;
  wire v372ea2d;
  wire v3727f68;
  wire v3a69dbd;
  wire v37737b9;
  wire v373f0d2;
  wire v37299de;
  wire v3807754;
  wire v3a61ff4;
  wire v372cfc2;
  wire v3a6a40b;
  wire v3a6333a;
  wire v37330d3;
  wire v3807020;
  wire v3a2976f;
  wire v1e37407;
  wire v3771e6d;
  wire v3a70503;
  wire v3741566;
  wire v3a66273;
  wire v3a6a0aa;
  wire v3a70a04;
  wire v3a70462;
  wire v3a60620;
  wire v3741609;
  wire v3a5e8a0;
  wire v3a707f5;
  wire v3758f02;
  wire v3768dbc;
  wire v374df4b;
  wire v3761e19;
  wire v3a6912a;
  wire v3726699;
  wire v3a65526;
  wire v372f216;
  wire v373339b;
  wire v3a5c59f;
  wire v3729f6c;
  wire v375c1d9;
  wire v37565ce;
  wire v377b706;
  wire v3a66210;
  wire v376277f;
  wire v3a6e0ab;
  wire v3765395;
  wire v3752091;
  wire v3a71592;
  wire v377b0fb;
  wire v3a6897b;
  wire v3a6f8c6;
  wire v3a612a9;
  wire v372c35a;
  wire v3768454;
  wire v3735461;
  wire v3747c10;
  wire v3a5dfe8;
  wire v3723485;
  wire v37662ac;
  wire v373f684;
  wire v360d144;
  wire v373daac;
  wire v376fdd6;
  wire v373351d;
  wire v3a6d32c;
  wire v3a6d0ec;
  wire v37718cc;
  wire v375899a;
  wire v3a70377;
  wire v3a5d186;
  wire v373c72a;
  wire v3774131;
  wire v3a6ecee;
  wire v3a5d8f6;
  wire v37556ce;
  wire v37503e7;
  wire v3a70658;
  wire v377311c;
  wire v3732f65;
  wire v3a70200;
  wire v3767018;
  wire v372b6db;
  wire v373bf74;
  wire v3a67a73;
  wire v372870d;
  wire v374fcd2;
  wire v3a579a3;
  wire v37413fc;
  wire v376348c;
  wire v3a70d9c;
  wire v3a6f0c9;
  wire v3a66dc0;
  wire v3757740;
  wire v3a60a2b;
  wire v377f4d5;
  wire v377ed8e;
  wire v3731eb5;
  wire v373f647;
  wire v372809d;
  wire v3a5d8a9;
  wire v3775064;
  wire v377ceb5;
  wire v374474d;
  wire v374caae;
  wire v37496b5;
  wire v37723a2;
  wire v3a70caf;
  wire v3779544;
  wire v3a602d7;
  wire v3759970;
  wire v373b4e6;
  wire v377fb43;
  wire v37525b0;
  wire v3a59c12;
  wire v3745928;
  wire v3765f61;
  wire v3763a1e;
  wire v3a54853;
  wire v3a70abc;
  wire v3749ddf;
  wire v375fba5;
  wire v3a55454;
  wire v373425d;
  wire v376cc45;
  wire v380663a;
  wire v3727e59;
  wire v377b6fc;
  wire v376ace2;
  wire v37556ae;
  wire v376740f;
  wire v3757e4a;
  wire v376c3f8;
  wire v3a70d5c;
  wire v3a6f04f;
  wire v3a5f89e;
  wire v3a700cd;
  wire v3744bfc;
  wire v3776ca9;
  wire v3a6cc78;
  wire v3a62cb5;
  wire v3a67beb;
  wire v3a6205a;
  wire v3767631;
  wire v377a968;
  wire v3a65c81;
  wire v3744539;
  wire v372dc20;
  wire cfe6df;
  wire v377aa17;
  wire v3a6206d;
  wire v3a714c7;
  wire v3a6ebe2;
  wire v3a59b6d;
  wire v3a712d5;
  wire v3750371;
  wire v1e37cec;
  wire v3754e5e;
  wire v9edb6a;
  wire v3a59424;
  wire v372ee0e;
  wire v37532c8;
  wire v37345a5;
  wire v3739915;
  wire v3733c7f;
  wire v3768e37;
  wire v3746e30;
  wire v376d657;
  wire v37298b2;
  wire v3a70214;
  wire v3a6c4e4;
  wire v3743d23;
  wire v375139d;
  wire v3728fcd;
  wire v3a56cdc;
  wire v3a6eb29;
  wire v3a7039e;
  wire v3a70ac8;
  wire v3728e1d;
  wire v37581a6;
  wire v376ff46;
  wire v3767ea6;
  wire v3a6650e;
  wire v372adaa;
  wire v373e484;
  wire v3a666bb;
  wire v376ab53;
  wire v3768c01;
  wire v3765f0a;
  wire v3775790;
  wire v3725d14;
  wire v3761470;
  wire v3769280;
  wire v3770af6;
  wire v3a68b25;
  wire v372f071;
  wire v3767dc8;
  wire v376d68d;
  wire v3768500;
  wire v37622aa;
  wire v37739ba;
  wire v3739b80;
  wire v3733de8;
  wire v373e72e;
  wire a5c257;
  wire v3a5b7c2;
  wire v375eb29;
  wire v3a700ea;
  wire v376d66c;
  wire v375070a;
  wire v3765627;
  wire v377d1a3;
  wire v3761fda;
  wire v3a60e38;
  wire v3a713ef;
  wire v3774757;
  wire v377a376;
  wire v3764881;
  wire v3a659b2;
  wire v3a7055a;
  wire v3a603f3;
  wire v3742476;
  wire v3741c39;
  wire v3a66819;
  wire v374c2e1;
  wire v374139a;
  wire v37590fb;
  wire v3a70ac4;
  wire v3a5c3c4;
  wire v3a67fc6;
  wire v3807315;
  wire v3774f38;
  wire v3740bcb;
  wire v879494;
  wire v37743c6;
  wire v374ce2a;
  wire v23fde41;
  wire v3a5cebe;
  wire v3775bca;
  wire v3752fbc;
  wire v3a711ea;
  wire v3724aaf;
  wire v3a70425;
  wire v37750f7;
  wire v3a6ff47;
  wire v37533c8;
  wire v3a6c82f;
  wire v374188e;
  wire v3766ff7;
  wire v37355ea;
  wire v375c2b1;
  wire v3a6fce5;
  wire v3768a41;
  wire v375449f;
  wire v3a575dc;
  wire v3a70978;
  wire v374d5c0;
  wire v376c62d;
  wire v374a2cc;
  wire v92e5bb;
  wire v374742c;
  wire v3729b2e;
  wire v3a70af5;
  wire v37594c5;
  wire v3a6cc72;
  wire v372c3a4;
  wire v3a70443;
  wire v376041f;
  wire v3a6fa19;
  wire v3779eea;
  wire v3a6607f;
  wire v3738365;
  wire v372fa7b;
  wire v3a61081;
  wire v3767897;
  wire v3a6f2c2;
  wire v3769d07;
  wire v3a644cd;
  wire v3a6f2c0;
  wire v3a60f71;
  wire v325c93e;
  wire v37706b3;
  wire v375f169;
  wire v372475d;
  wire v3766f1c;
  wire v375c06a;
  wire v377d8b7;
  wire v3a6f4eb;
  wire v377211f;
  wire v3750d19;
  wire v3761d7d;
  wire v3809f0e;
  wire v376c789;
  wire v3a6e0cc;
  wire v376219d;
  wire v3a700ce;
  wire v37678bd;
  wire v3a70a7e;
  wire v373112c;
  wire v373b6ba;
  wire v372f9b4;
  wire v3a709b5;
  wire v37375ed;
  wire v3749fdc;
  wire v3a56531;
  wire v3a59cae;
  wire v373ed5c;
  wire v3a708ce;
  wire v3a661c2;
  wire v3809e90;
  wire v2acaee4;
  wire v375cd7b;
  wire v3767483;
  wire v37290fa;
  wire v37498bd;
  wire v3a70cb2;
  wire v37424df;
  wire v372fecd;
  wire v3a5f2c0;
  wire v3a679b5;
  wire v3a706b8;
  wire v376e3a3;
  wire v3769b1d;
  wire v375b046;
  wire v3a658f7;
  wire v3753d03;
  wire v3a6ff36;
  wire v375f0d4;
  wire v374aa4f;
  wire v372c83a;
  wire v2acb094;
  wire v374478a;
  wire v3747a36;
  wire v3a6f3ac;
  wire v377380a;
  wire v3740fe2;
  wire v3749bba;
  wire v373feaa;
  wire v3a62dfa;
  wire ab808e;
  wire v37398e5;
  wire v3771739;
  wire v373e6eb;
  wire v372bc46;
  wire v3a70c1d;
  wire v373a4ea;
  wire v37343e7;
  wire v37403cc;
  wire v3736eee;
  wire v37283f8;
  wire v3746ce0;
  wire v375c600;
  wire v3a6f9cd;
  wire v3763183;
  wire v3765e5b;
  wire v3a70f1e;
  wire v375b99c;
  wire v3a5f447;
  wire v3770a82;
  wire v376cfae;
  wire v3a67f5b;
  wire v3a5d11d;
  wire v376d780;
  wire v23fe316;
  wire v37659c5;
  wire v3a6fa58;
  wire v3a6ef56;
  wire v3766a37;
  wire v3a6f7fe;
  wire v376069d;
  wire v3a6d8f4;
  wire v3739983;
  wire v3a60ac5;
  wire v3a63f77;
  wire v3723447;
  wire v376f468;
  wire v3774af1;
  wire v37363fd;
  wire v3a6feca;
  wire v3a6ebaf;
  wire v3a7033d;
  wire v3a57d41;
  wire v3a6fc18;
  wire v3a5c40b;
  wire v37621b5;
  wire v3a65241;
  wire v3a55fc6;
  wire v372c5e4;
  wire v375e624;
  wire v3757169;
  wire v3a5b517;
  wire v23fdaf1;
  wire v3a6f9bb;
  wire v375d366;
  wire v9342d1;
  wire v3a7099f;
  wire v3a7124f;
  wire v376b962;
  wire v376ad46;
  wire v3a689b8;
  wire v37629db;
  wire v3a70d4a;
  wire v37bfff7;
  wire v3a6fb9f;
  wire v376afff;
  wire v376b662;
  wire v376a7ac;
  wire v3a6f336;
  wire v3767419;
  wire v376a863;
  wire v374b3b5;
  wire v3744887;
  wire v373cbc5;
  wire v3a7091e;
  wire v3a6fae3;
  wire v3728906;
  wire v3757569;
  wire v38072f0;
  wire v3a70149;
  wire v3a5c4e1;
  wire v3750cfa;
  wire v3724665;
  wire v3378f5b;
  wire v3a6f929;
  wire v3a700d9;
  wire v372cb9d;
  wire v3770827;
  wire v3732558;
  wire v3a70606;
  wire v3772c8e;
  wire v35ba1c6;
  wire v3a713cd;
  wire v373a072;
  wire v374bc97;
  wire v3a70700;
  wire v3a70e5c;
  wire v373fecb;
  wire v3a6f9ab;
  wire v377a887;
  wire v373e55b;
  wire v3736ea9;
  wire v3723749;
  wire v38093a8;
  wire v373700d;
  wire v3a70570;
  wire v372b172;
  wire v3756cf2;
  wire v3752913;
  wire v3a58e15;
  wire v3744c88;
  wire v376b87b;
  wire v3a6eb28;
  wire v3771d70;
  wire v3a7042d;
  wire v3a5fc9c;
  wire v3a70b12;
  wire v3772464;
  wire v375fcfa;
  wire v377b848;
  wire v3a6f8ec;
  wire v373862e;
  wire v3a5948f;
  wire v377dca9;
  wire v3a6f601;
  wire v3a6deaa;
  wire v3a6fc42;
  wire v3a6f106;
  wire v3749580;
  wire v3a7018b;
  wire v3a6fa1c;
  wire v3a5a2cd;
  wire v3a2abf4;
  wire v3a70878;
  wire v3a575e5;
  wire v3765268;
  wire v372954d;
  wire v3a6f70f;
  wire v372ed89;
  wire v373f4cf;
  wire v3808884;
  wire a0715f;
  wire v3738e62;
  wire v3a6ed55;
  wire v372704f;
  wire v377074b;
  wire v377f66c;
  wire v3a70a9e;
  wire v373a265;
  wire v374373a;
  wire v3778023;
  wire v3a59283;
  wire v373738e;
  wire v3a6582d;
  wire v376dd80;
  wire v3a6443f;
  wire v37293f2;
  wire v3a6ff8d;
  wire v3a70380;
  wire v3a702d8;
  wire v37469ba;
  wire v3a6f945;
  wire v374cc43;
  wire v3755e1f;
  wire v3728dd0;
  wire bca64b;
  wire v3a6199f;
  wire v3755967;
  wire v37312f4;
  wire v3a6f427;
  wire v3735930;
  wire v373f88a;
  wire v3a6c6ac;
  wire v3a62ce4;
  wire bb3b0a;
  wire v3733a0e;
  wire v3738279;
  wire v372a27f;
  wire v3743012;
  wire v3a6869f;
  wire v3a6b4db;
  wire v372e8f2;
  wire v37241a0;
  wire v3a571e5;
  wire v3761f74;
  wire v3776ce3;
  wire v376766e;
  wire v3a6a990;
  wire v3a5ac8b;
  wire v3a62cac;
  wire v3a7059e;
  wire v3759b09;
  wire v376fbff;
  wire v3769e01;
  wire v3a2951d;
  wire v37368bb;
  wire v3744bed;
  wire v372d24a;
  wire v3735da7;
  wire v3775c24;
  wire v3a64032;
  wire v38069e7;
  wire v374d3b0;
  wire v37723ed;
  wire v3a6aaed;
  wire v3745b71;
  wire v3a5c7ca;
  wire v3749658;
  wire v3726ddb;
  wire v3a6fcdf;
  wire v3a62f72;
  wire v3769db7;
  wire v3767c16;
  wire v3730a90;
  wire v3a7166e;
  wire v3729370;
  wire v374dba6;
  wire v3a6fb42;
  wire v3a6fe15;
  wire v372da95;
  wire v375d1e1;
  wire v373a2cc;
  wire v3a6fd3d;
  wire v375b483;
  wire v3a7130f;
  wire c6fb51;
  wire v3a6eb26;
  wire v3a6ff75;
  wire v376babf;
  wire v3727342;
  wire v37793d4;
  wire v372c0de;
  wire v374e1fd;
  wire v3a61b45;
  wire v377cc6d;
  wire v3727889;
  wire v3a53ae0;
  wire v3a7121a;
  wire bb0568;
  wire v374fc3b;
  wire v375e62f;
  wire v373a4b2;
  wire v3745b5b;
  wire v3a6f073;
  wire v376e79d;
  wire v372a77a;
  wire v373f996;
  wire v374bc63;
  wire v372580c;
  wire v376a6ae;
  wire v3a653d5;
  wire v37470e6;
  wire v3a617a2;
  wire v37392e2;
  wire v3755786;
  wire v375994d;
  wire v3a5cca9;
  wire v374e109;
  wire v372571e;
  wire v3741438;
  wire v1e38262;
  wire v375792c;
  wire v3a704be;
  wire v3723d73;
  wire v377104a;
  wire v3a5caf4;
  wire v3a5e922;
  wire v3723abc;
  wire v374352b;
  wire v375d134;
  wire v3a6d81d;
  wire v375e527;
  wire v376eea3;
  wire v37660f2;
  wire v3a7083c;
  wire v3755bbf;
  wire v3a71557;
  wire v373b747;
  wire v3a715fc;
  wire v3756263;
  wire v3a70235;
  wire v377bae8;
  wire v373d3ec;
  wire v3a5bbbb;
  wire v3724b5a;
  wire v3a693dc;
  wire v9a88fd;
  wire v3740f65;
  wire v3747b02;
  wire v376ecde;
  wire v375dd87;
  wire v3807386;
  wire v3772214;
  wire v375f798;
  wire v3a675df;
  wire v3a70c8e;
  wire v37555fd;
  wire v3a65174;
  wire v3a65652;
  wire v372c6ce;
  wire v376de00;
  wire v3729bd1;
  wire v3a6046d;
  wire v374e788;
  wire v377b017;
  wire v3764f01;
  wire v372a02b;
  wire v23fde69;
  wire v3744aaa;
  wire v373f53e;
  wire v3a6ba88;
  wire v3738a87;
  wire v3765c08;
  wire v3a70c87;
  wire v3a6e8b1;
  wire v376373e;
  wire v3755640;
  wire v3a5e3f1;
  wire v372d4d4;
  wire v3743a49;
  wire v3764f5c;
  wire v377ad63;
  wire v3734374;
  wire v372505f;
  wire v3772231;
  wire v3728fd2;
  wire v373cc9a;
  wire v376ba63;
  wire v3a5c46a;
  wire v373b732;
  wire v3a70103;
  wire v3a71245;
  wire v3a61dd0;
  wire v37655ff;
  wire v3a6f89b;
  wire v373e76c;
  wire v374f2fb;
  wire v374d14a;
  wire v37274a1;
  wire v3a71461;
  wire v376634b;
  wire v3763387;
  wire v375f848;
  wire v374e745;
  wire v3740825;
  wire v376497a;
  wire v37465c7;
  wire v373c7af;
  wire v375b676;
  wire v3778f32;
  wire v374c000;
  wire v3a714b0;
  wire v3a58e79;
  wire v375583c;
  wire v3a5b46d;
  wire v3a56d04;
  wire v3a6f826;
  wire v37460de;
  wire v37617b9;
  wire v3759758;
  wire v3753e8e;
  wire v3a691fb;
  wire v373bfd8;
  wire v3778fae;
  wire cc9e54;
  wire v3255a0f;
  wire v3a61d9f;
  wire v3a70041;
  wire v37664c5;
  wire v3a56130;
  wire v3a5f717;
  wire v374307e;
  wire v3a71116;
  wire v375f071;
  wire v372773c;
  wire v90b307;
  wire v3a6f253;
  wire v373556f;
  wire v3a6f1db;
  wire v373471a;
  wire v3a5d7f7;
  wire v372b840;
  wire v3a70d5f;
  wire v373ec1f;
  wire v374bd38;
  wire v376abd3;
  wire v375c07c;
  wire v3a6f3df;
  wire v3a70581;
  wire v3a54cd9;
  wire v97c94a;
  wire v373f11a;
  wire v37510b9;
  wire v3755045;
  wire v373a452;
  wire v374a9a0;
  wire v3736e7d;
  wire v3a57fb8;
  wire v3a669bc;
  wire v3759f77;
  wire v375cd8b;
  wire v91f9a4;
  wire v3a69f4e;
  wire v3746cc3;
  wire v3745473;
  wire v373d203;
  wire b69f28;
  wire v376726e;
  wire v3a5beb8;
  wire v3a550c2;
  wire a85c8e;
  wire v3a70e2f;
  wire v3a673fa;
  wire v3a6eb0d;
  wire v373ab06;
  wire v37781d4;
  wire v373b2ba;
  wire v374aa0f;
  wire v372facf;
  wire v372d538;
  wire v37368c8;
  wire v3a705cc;
  wire v2acaed7;
  wire v3762806;
  wire v3a5ce55;
  wire v3724872;
  wire v3764331;
  wire v3a70743;
  wire v3a5cc79;
  wire v3752d24;
  wire v3747e1f;
  wire v3772c95;
  wire v3a55c8f;
  wire v3a5b571;
  wire v377faa6;
  wire v37324e7;
  wire v3a5db83;
  wire v372cf2e;
  wire v3a6cd89;
  wire v3a70306;
  wire v3809e41;
  wire v3a702dd;
  wire v3770359;
  wire v3773bd7;
  wire v3754a8e;
  wire v3a6fbec;
  wire v375db64;
  wire v375647b;
  wire v377be84;
  wire v3a659eb;
  wire v373520f;
  wire v374efb3;
  wire v3745072;
  wire v3739e31;
  wire v3a70081;
  wire v37665e2;
  wire v23fe324;
  wire v37317ec;
  wire v3747a5b;
  wire v3747c4c;
  wire v3730749;
  wire v3a7096f;
  wire v3a67c50;
  wire v372a22f;
  wire v3a6ff6f;
  wire v37253dc;
  wire v375aa9b;
  wire v3736958;
  wire v3736b1d;
  wire v3769a34;
  wire v373dd36;
  wire v3a701f2;
  wire v376c0d8;
  wire v37494ed;
  wire d9e97c;
  wire v374fdeb;
  wire v376e562;
  wire v37463d4;
  wire v3a5a484;
  wire v3754392;
  wire v3a59c1d;
  wire v3779e29;
  wire v3a2a0e9;
  wire v374d1d7;
  wire v37432e2;
  wire v3764677;
  wire v3a6ae04;
  wire v3a67e25;
  wire b46885;
  wire v373a6bf;
  wire v375dc5f;
  wire v372750b;
  wire v376af8c;
  wire v37485df;
  wire v3a611cf;
  wire v376ea50;
  wire v3745e71;
  wire v376bc5b;
  wire v3777140;
  wire v3751f34;
  wire v377df2e;
  wire v374bc02;
  wire v377b7ad;
  wire v37414d1;
  wire v3726204;
  wire v3a705f0;
  wire v3a6fd5c;
  wire baccec;
  wire v3a6c970;
  wire v3a6ef95;
  wire v3767b6e;
  wire v3a6848c;
  wire v3752281;
  wire v3760eb8;
  wire v375648e;
  wire v375efa4;
  wire v375fcbf;
  wire a8c5c5;
  wire v373afc3;
  wire v374e380;
  wire v3738169;
  wire v377de50;
  wire v374fc20;
  wire v37263c3;
  wire v375820a;
  wire v376d1b4;
  wire v376462a;
  wire v377597f;
  wire v3a6ead8;
  wire v3a56580;
  wire v3765d74;
  wire v2925cbb;
  wire v3a6581d;
  wire v3a6fdde;
  wire v3736806;
  wire v37690bf;
  wire v3a7137c;
  wire v3a6ea66;
  wire v3732e09;
  wire v3a6f3b8;
  wire v3a603c1;
  wire c79715;
  wire v37316ec;
  wire v373bbb4;
  wire v3a7088a;
  wire d0c237;
  wire v3a5d929;
  wire v3a53c63;
  wire v3a6b306;
  wire v3a68232;
  wire v374bace;
  wire v3a7012a;
  wire v3a70b3f;
  wire v3761953;
  wire v3762a37;
  wire v3a70d07;
  wire v375c3f6;
  wire v3a698ed;
  wire v374cb24;
  wire v37280a0;
  wire v3a70a57;
  wire v376d3cb;
  wire v2acae60;
  wire v3741ba8;
  wire v3a70706;
  wire v374f0af;
  wire v373ab7e;
  wire v373653b;
  wire v3736adf;
  wire v374e207;
  wire v377f24b;
  wire v374216a;
  wire v3a56ebd;
  wire v3a6db95;
  wire v3a715e5;
  wire v37604d6;
  wire v2092abf;
  wire v373ae27;
  wire v377e710;
  wire v3a6f3ef;
  wire v3a5ab05;
  wire v376d48b;
  wire v37730ec;
  wire v3a6f047;
  wire v3750519;
  wire v861ce0;
  wire v37599a4;
  wire v3769101;
  wire b6a7cc;
  wire v377cc7b;
  wire v3a6f61a;
  wire v3746fcb;
  wire v375c2d0;
  wire v374c556;
  wire v372c959;
  wire v87f2ea;
  wire v374fde8;
  wire v376654b;
  wire v375bab8;
  wire v373bcdd;
  wire v3a59c21;
  wire v3767471;
  wire v374407c;
  wire v373a3e7;
  wire v373dc5a;
  wire v37356a7;
  wire v3778211;
  wire v3725dbb;
  wire v3a704e9;
  wire v3a7037a;
  wire v3754488;
  wire v3a70b9f;
  wire v3a6fac3;
  wire v3a70daf;
  wire v3a61e79;
  wire v3a6c0b7;
  wire v3735fe8;
  wire v3762fdb;
  wire v3a65b39;
  wire v3a6e916;
  wire v3730f21;
  wire v3777e59;
  wire v3a70a58;
  wire v37433e6;
  wire v3a711a8;
  wire v375aa0d;
  wire v3a60b56;
  wire v373335b;
  wire v37507a8;
  wire v38078ea;
  wire v3a700d3;
  wire v3809b53;
  wire v2092bfc;
  wire v376dee4;
  wire v373a85c;
  wire v3725612;
  wire v3a6f40a;
  wire v375016d;
  wire v3a6f2c6;
  wire v3a70194;
  wire v3754ddd;
  wire v372df76;
  wire v3a57e27;
  wire v3a7058d;
  wire v3733384;
  wire v372b971;
  wire v3735302;
  wire v37793cd;
  wire v377b735;
  wire v377664f;
  wire v3a541f5;
  wire v373c916;
  wire v3a6f43b;
  wire v3724b20;
  wire v3768a11;
  wire v3a70b26;
  wire v3737897;
  wire v374763e;
  wire v376e4c5;
  wire v372715f;
  wire v3a6c0f1;
  wire v376fbd0;
  wire v3a6fb30;
  wire v3765385;
  wire v3a5d527;
  wire v3735936;
  wire v3723f71;
  wire v3759c80;
  wire v3a6de3a;
  wire v372700e;
  wire v3a532f2;
  wire v3a70a85;
  wire v3a715a2;
  wire v380700f;
  wire v373d119;
  wire v3a53962;
  wire v3a70c4c;
  wire v3730288;
  wire v375dda4;
  wire v3762847;
  wire v3725804;
  wire v1e37d14;
  wire v3a6faed;
  wire v3738336;
  wire v3752845;
  wire v377a886;
  wire v3768172;
  wire v3778b83;
  wire v3772e3f;
  wire v375facd;
  wire v3755dfa;
  wire v3a6d3c9;
  wire v375c6cc;
  wire v3a59656;
  wire v374743a;
  wire v3748851;
  wire v8455f3;
  wire v3a70f2a;
  wire v3a5d9bc;
  wire v360ba91;
  wire v3a7166b;
  wire v3a6f0f4;
  wire v3a6903e;
  wire v377c9b3;
  wire v37348e5;
  wire v374cad6;
  wire v3747462;
  wire v3775544;
  wire v3744aca;
  wire v377e7f8;
  wire v3753f36;
  wire v3903ee2;
  wire v375025f;
  wire v372fe3d;
  wire v3a66e7f;
  wire v3a5ef0d;
  wire v3a5f375;
  wire v8455b1;
  wire v3a63de8;
  wire v3a6ff68;
  wire d95e20;
  wire v3a6fc50;
  wire v375f689;
  wire v3a5e0dd;
  wire v380a20c;
  wire v8455e3;
  wire v375956a;
  wire v376f693;
  wire v3732170;
  wire v3a63e82;
  wire v376e914;
  wire v3724398;
  wire v37503bd;
  wire v37231e5;
  wire v373f497;
  wire v3756234;
  wire v3a637dc;
  wire v3a637dd;
  wire v3a653e4;
  wire v3759dfb;
  wire v3a705cb;
  wire v373327e;
  wire v3730601;
  wire v37300ba;
  wire v375d23b;
  wire v3a64e13;
  wire v3a68b0a;
  wire v2ff87c6;
  wire v3a6fdec;
  wire v3776cda;
  wire v37594ae;
  wire v37346be;
  wire v3738686;
  wire v3a6ef50;
  wire v209310e;
  wire v937864;
  wire v375fb00;
  wire v3a6b873;
  wire v3a554d8;
  wire v3a71232;
  wire v374b962;
  wire v3750d06;
  wire v374514c;
  wire v3a6f5cd;
  wire v8a94c2;
  wire v3809892;
  wire v3a5cf3c;
  wire v3a7137d;
  wire v20930c9;
  wire v3a6f563;
  wire v37797f4;
  wire v3773daf;
  wire v3754bb9;
  wire v3a5a2d0;
  wire v3808db7;
  wire v375023c;
  wire v3a709d9;
  wire v373d381;
  wire v3a62a2d;
  wire v3a594e8;
  wire v374831d;
  wire v3a5ba8f;
  wire v373b5c1;
  wire v3740777;
  wire v3771901;
  wire v3750e4f;
  wire v37651e0;
  wire v3a5f97f;
  wire v373ee66;
  wire v3a6eb88;
  wire v37363f8;
  wire v373ff97;
  wire v376243f;
  wire v37322d8;
  wire v372c23f;
  wire v372a9c2;
  wire v3737c21;
  wire v3a61988;
  wire v3a6feed;
  wire v3732a41;
  wire v37687ce;
  wire v374f0c1;
  wire v3a57330;
  wire v372692d;
  wire v3a6cf18;
  wire v376f45e;
  wire v37356ce;
  wire v3a5fa18;
  wire v374e753;
  wire v374fe73;
  wire v376a39c;
  wire v3a709ee;
  wire v37323a2;
  wire v3a71273;
  wire v37270b5;
  wire v3765583;
  wire v376b561;
  wire v3728a45;
  wire v372f0ee;
  wire v3746d75;
  wire v3807b40;
  wire v3a54f04;
  wire v3a6fadd;
  wire v3a7145b;
  wire v376a1d7;
  wire v3a6fca5;
  wire v372fc77;
  wire v3779f13;
  wire v37425a1;
  wire v37290a1;
  wire v3727986;
  wire v377c7ae;
  wire v3a6fa11;
  wire v3a553aa;
  wire v37313fa;
  wire v37435e9;
  wire v373ac65;
  wire v3a618ea;
  wire v3a58fe9;
  wire v3a711f7;
  wire v3750746;
  wire v3763961;
  wire v373df14;
  wire v37328a1;
  wire v3a66140;
  wire v3a70208;
  wire d27546;
  wire v3a70a92;
  wire v37373af;
  wire v3a696a7;
  wire v3a62efa;
  wire bde868;
  wire v3a6f891;
  wire v3a676f1;
  wire v372b7a8;
  wire v37695c7;
  wire v373da1b;
  wire v3a7023d;
  wire v3745536;
  wire v3749dad;
  wire v3a7048a;
  wire v3a568ac;
  wire v374f4a0;
  wire v37717f4;
  wire v37509af;
  wire b8006a;
  wire v37497b1;
  wire v3a6e236;
  wire v376640b;
  wire v3a70286;
  wire v3753317;
  wire v3a60bbf;
  wire v372c197;
  wire v3a66037;
  wire v377e784;
  wire v3757dd1;
  wire v3a6b27e;
  wire v3a61336;
  wire v3722b17;
  wire v372f71f;
  wire v374d1ad;
  wire v3a70617;
  wire v3773847;
  wire v3a6f508;
  wire v3a712f6;
  wire v3a7124d;
  wire v37385ee;
  wire v37421bd;
  wire v3a6f290;
  wire v3726cf7;
  wire v377f342;
  wire v3734f09;
  wire v3739f84;
  wire v3750c59;
  wire v3a66a01;
  wire v2092f0f;
  wire v3a6f3a8;
  wire v3765fcf;
  wire v37739c6;
  wire v3758c65;
  wire v37630d9;
  wire v3a5baaf;
  wire v3764114;
  wire v3a5fbad;
  wire v3a6f244;
  wire v375d507;
  wire v3729238;
  wire v377e8be;
  wire v3a6f7de;
  wire v3a6b083;
  wire v3a5ea7b;
  wire v3755296;
  wire v375b04f;
  wire v3743e83;
  wire v375518f;
  wire v3761769;
  wire v3723296;
  wire v3a6faeb;
  wire v3a53d1e;
  wire v3759c2e;
  wire v375b203;
  wire v377911e;
  wire v3a6effa;
  wire v3a64e40;
  wire v377d2a0;
  wire v3a70cab;
  wire v376c2d6;
  wire v3a6a516;
  wire v1e37dcd;
  wire v3728040;
  wire v3a7164f;
  wire v372cd8b;
  wire v3a635b1;
  wire v3744039;
  wire v372a93f;
  wire b02944;
  wire dc33c0;
  wire v3728389;
  wire v376d774;
  wire v3a715d1;
  wire d7e38d;
  wire v37621e0;
  wire v3766bdf;
  wire v374554d;
  wire v3a6f54f;
  wire v37487b0;
  wire v376c72f;
  wire v377cc25;
  wire v375603c;
  wire v3777573;
  wire v374109e;
  wire v375c769;
  wire v37560f7;
  wire v3a53da1;
  wire v373554b;
  wire v3a6a289;
  wire v3733887;
  wire v3a70c0b;
  wire v372dab0;
  wire v375dd29;
  wire v3a6da3b;
  wire v3a64977;
  wire v37419b4;
  wire v3732f00;
  wire v3727f86;
  wire v37426ed;
  wire v373f56b;
  wire v3729a9f;
  wire v3a7003e;
  wire v3a671a2;
  wire v372e4b3;
  wire v37259e6;
  wire v377f67b;
  wire v3750cae;
  wire v3a70f20;
  wire v3a70401;
  wire v372aafb;
  wire v374c9ee;
  wire v3765b30;
  wire v3a5a798;
  wire v374cb90;
  wire v3738419;
  wire v360d07a;
  wire v3750b61;
  wire v3778277;
  wire v3a715d6;
  wire v9b63b0;
  wire v3736d97;
  wire v3a6a33a;
  wire v3a68ad7;
  wire v2ff8bb1;
  wire v372e268;
  wire v3a6992f;
  wire v373f7ef;
  wire v3a6ac2c;
  wire v3737bfe;
  wire v3725088;
  wire v35b70d2;
  wire v3739916;
  wire v372fe43;
  wire v3a6de5e;
  wire v3a7038d;
  wire v3a5e0c9;
  wire v374c144;
  wire v3774c98;
  wire v3a58761;
  wire v377f2bb;
  wire v3a6f64a;
  wire v37680de;
  wire v2092eb6;
  wire v3a66c49;
  wire v3739e4c;
  wire v377f6ff;
  wire v374e248;
  wire v3a669ac;
  wire v376e1b7;
  wire v377cbc9;
  wire v23fe061;
  wire v374a556;
  wire v3a692f6;
  wire v3a6eb36;
  wire v3763bc4;
  wire v3a6f191;
  wire v3766bbb;
  wire v374e2a0;
  wire v3a710c4;
  wire v3769cac;
  wire v3a70472;
  wire v39a4ef6;
  wire v3a7079b;
  wire v3755d23;
  wire v373923a;
  wire v3725b1f;
  wire v3765322;
  wire v3729e65;
  wire v3761ad8;
  wire v3a706d3;
  wire v3a69f17;
  wire v374e531;
  wire v3a66d7e;
  wire v3a609bb;
  wire v3a706e3;
  wire v3a6b8a0;
  wire v3a6767a;
  wire v3a56c66;
  wire v3741baf;
  wire v37450a5;
  wire v3759a34;
  wire v2ff8e1f;
  wire v3a702e9;
  wire v377246b;
  wire v374cc40;
  wire v3807b2e;
  wire v3756740;
  wire v3a551d7;
  wire v3a6f2be;
  wire v377795a;
  wire v37444c9;
  wire v3768d7e;
  wire v3a634fa;
  wire v3743407;
  wire v3a5ebde;
  wire v3770ccf;
  wire v3779be2;
  wire v376110e;
  wire v372cfeb;
  wire v37385de;
  wire v3775626;
  wire v3a5ed4a;
  wire v3a65b2b;
  wire v3758c64;
  wire v376db07;
  wire v2678c40;
  wire v3a5bc35;
  wire v3759fca;
  wire v377855f;
  wire v3a565ef;
  wire v3750403;
  wire v3a6e8bc;
  wire v376bf97;
  wire v1e37e4f;
  wire v3a602cd;
  wire v37605ab;
  wire v3764210;
  wire v3735a94;
  wire v375637c;
  wire v376c784;
  wire v372f357;
  wire v3742cce;
  wire v3729caa;
  wire v3a56abc;
  wire v373ec4c;
  wire v3806828;
  wire v3a64c73;
  wire v376233b;
  wire v3778a91;
  wire v3773430;
  wire v372dd14;
  wire v3a6eaea;
  wire v3a712a1;
  wire v3751981;
  wire v3732cf6;
  wire v3a66a86;
  wire v3767dac;
  wire v3773091;
  wire v3754586;
  wire v3750deb;
  wire v376e76f;
  wire v3747467;
  wire v3a57496;
  wire v375c883;
  wire v3a582c5;
  wire v3a665b3;
  wire v3a71307;
  wire v372f6f9;
  wire v3a67b3c;
  wire v3755670;
  wire v374c1a0;
  wire v377af5d;
  wire v3a70342;
  wire v373a3a7;
  wire v3a70bdf;
  wire v3a71312;
  wire v373a982;
  wire v3a70ff9;
  wire v3749c91;
  wire v3778fa0;
  wire v37580b3;
  wire v376a91d;
  wire v372dfc1;
  wire v3730118;
  wire v3a70e2a;
  wire v3a6fe21;
  wire v3729996;
  wire v376ebc6;
  wire v3a6b17e;
  wire v373ae2e;
  wire v3733350;
  wire v3a7044c;
  wire v3a70df1;
  wire v374d552;
  wire v375538a;
  wire v374ad82;
  wire v3728dc7;
  wire v3762455;
  wire v3767d55;
  wire v3774061;
  wire v374fb93;
  wire v3764e95;
  wire v37765d0;
  wire v376888c;
  wire v3a6f6cf;
  wire v3739938;
  wire v3761e62;
  wire v374385c;
  wire v375d1d4;
  wire v3a68e10;
  wire v374f834;
  wire v377d496;
  wire v3a64854;
  wire v374fac9;
  wire v37712e5;
  wire v3a6accb;
  wire v3730862;
  wire v375d7bc;
  wire v37464f0;
  wire v37762b6;
  wire v37500c2;
  wire v37326a1;
  wire v375787b;
  wire v3809d87;
  wire v3a71601;
  wire v1e37a26;
  wire v3740db1;
  wire v37539ef;
  wire v373ca5f;
  wire v375a858;
  wire v3a6f6df;
  wire v3a703ca;
  wire v3a5a374;
  wire v372a9bd;
  wire v3759590;
  wire v3a683d2;
  wire v3777386;
  wire v3a6f52e;
  wire v377c44f;
  wire v375de43;
  wire v376f29d;
  wire v39eb517;
  wire v3733fd8;
  wire v377903f;
  wire v376b99f;
  wire v3747d37;
  wire v3745704;
  wire v3757c7d;
  wire v376d81c;
  wire v372ab80;
  wire v374a9eb;
  wire v3a714da;
  wire v374fcde;
  wire v373a267;
  wire v375b282;
  wire v3a6a2ab;
  wire v37519e5;
  wire v372e865;
  wire v37287fa;
  wire v377740c;
  wire v3a713d7;
  wire v3a6dea7;
  wire v37500e2;
  wire v373812a;
  wire v372b2cb;
  wire v3753a8a;
  wire v374b394;
  wire v375a268;
  wire v377de6f;
  wire v376a85d;
  wire v3747b30;
  wire v3764276;
  wire v3727a4d;
  wire v3a700fa;
  wire v37730df;
  wire v3a65335;
  wire v374fb58;
  wire v37648af;
  wire v3750ea5;
  wire v3746806;
  wire v376d882;
  wire v3a708a7;
  wire v3a70592;
  wire v3726139;
  wire v3a70806;
  wire v3751c4c;
  wire v3775107;
  wire v372aacd;
  wire v3726434;
  wire v373f022;
  wire v3736048;
  wire v3739a23;
  wire v37420de;
  wire v377d497;
  wire v375d1a1;
  wire v3a6eecb;
  wire v3a70cfa;
  wire v37691b8;
  wire v3743c90;
  wire v3732be9;
  wire v377a9fc;
  wire v372f320;
  wire v3756764;
  wire v3a6f48a;
  wire v377a4bd;
  wire v3771be4;
  wire v3a710a3;
  wire v37781fe;
  wire v3a6f774;
  wire v3742a8b;
  wire v372e47b;
  wire v37650c4;
  wire v3a56b80;
  wire v3a6f8be;
  wire v3733cfb;
  wire v3a675b9;
  wire v373ee19;
  wire v3764530;
  wire v3770b33;
  wire v3740f89;
  wire v3a70d88;
  wire v3771a36;
  wire v377d320;
  wire v37583f2;
  wire v3808658;
  wire v3a65161;
  wire v23fdbdc;
  wire v375da17;
  wire v3764df7;
  wire v3a70f48;
  wire v375d337;
  wire v3767e66;
  wire v373ebac;
  wire v3a683f9;
  wire v372664e;
  wire v3730de9;
  wire v374f033;
  wire v374053e;
  wire v376e9e2;
  wire v3a713dc;
  wire v37565a0;
  wire v3766e29;
  wire v372d8e8;
  wire a3d29c;
  wire v375a5f9;
  wire v3a6f487;
  wire v3a5907f;
  wire v3a690ff;
  wire v377a018;
  wire v3a6f656;
  wire v3a684af;
  wire v37758ce;
  wire v375fd38;
  wire v374e314;
  wire v3750e32;
  wire v3743113;
  wire v3735cfb;
  wire v3751a0d;
  wire v3770a83;
  wire v376ff42;
  wire v3a55c48;
  wire v3728992;
  wire v374a9e7;
  wire v375bd9c;
  wire v3744e11;
  wire v37325f4;
  wire v3a5755b;
  wire v3a53ffa;
  wire v377564a;
  wire v377754d;
  wire v3771360;
  wire v2925c5b;
  wire v3a710d0;
  wire v372f770;
  wire v373a1f2;
  wire v374262d;
  wire v3733234;
  wire v3750b03;
  wire v3a6d175;
  wire v37330b1;
  wire v375ad1d;
  wire v3729c37;
  wire v3747035;
  wire v372fd45;
  wire v37391e8;
  wire v37310c2;
  wire v3a6fc2d;
  wire v3a6462c;
  wire v3378996;
  wire v3a60fa7;
  wire v3a6fe31;
  wire v376acd9;
  wire v3a6ef91;
  wire v375c5cf;
  wire v37292f4;
  wire v3763299;
  wire v373ce74;
  wire v3744a0c;
  wire v3a70ded;
  wire v3730f77;
  wire v3a623f2;
  wire v3a6d806;
  wire v3766eef;
  wire v3a682a1;
  wire v3765699;
  wire v374394c;
  wire v3731079;
  wire v374dcbd;
  wire v3a63135;
  wire v375bdf0;
  wire v3725bea;
  wire v3a5e6b2;
  wire v3774cde;
  wire v376b5a4;
  wire v3763ce3;
  wire v3a6f48c;
  wire v375401a;
  wire v376a21c;
  wire v3808d42;
  wire v3a701cd;
  wire v1e379f7;
  wire v3a6f0ed;
  wire v3775b82;
  wire v3739ea5;
  wire v374c9c2;
  wire v3a71497;
  wire v376ee82;
  wire v3763716;
  wire v3a70d2b;
  wire v35ba2cb;
  wire v3a6f55a;
  wire v37781b7;
  wire v3a6f173;
  wire v3725269;
  wire v3a715eb;
  wire v376978e;
  wire v377463d;
  wire v377b5aa;
  wire v372ef62;
  wire v37726b0;
  wire v373e8de;
  wire v3a55352;
  wire v3a70111;
  wire v373139d;
  wire v3a63994;
  wire v39ed7e4;
  wire v376e5ef;
  wire v3742ed3;
  wire v3a71352;
  wire v39ed7ea;
  wire v3985138;
  wire v2ff8d08;
  wire v37530d1;
  wire v372debd;
  wire v3a70772;
  wire v373fc77;
  wire v3985143;
  wire v3a70f3f;
  wire v3a61a1d;
  wire v39af33c;
  wire v3a70641;
  wire v374b51f;
  wire v372c524;
  wire v3a6373e;
  wire v375b258;
  wire v3a56346;
  wire v3a690ec;
  wire v3806db7;
  wire v3a677ce;
  wire v3a71509;
  wire v3a6e431;
  wire v372b7fb;
  wire v3732eca;
  wire v377ba55;
  wire v3a6e91e;
  wire v37637d4;
  wire v23fdead;
  wire v3a70ce4;
  wire v3729ca6;
  wire v3a6869d;
  wire v372fba5;
  wire v3746211;
  wire v3747192;
  wire v8455d5;
  wire v3722f37;
  wire v3742b0e;
  wire v3a5ca7b;
  wire v3724940;
  wire v3747a7b;
  wire v3a70b15;
  wire v3a67b93;
  wire v3739a05;
  wire v377e310;
  wire v3a70f23;
  wire v37435f1;
  wire v3a6ec30;
  wire v3778bb4;
  wire v3a71604;
  wire v3735da3;
  wire v37612d0;
  wire v372ae4f;
  wire v3750fa9;
  wire v373fdce;
  wire v374c6aa;
  wire v3a6a81f;
  wire v373cdb4;
  wire v3727345;
  wire v3a5d532;
  wire v376a14f;
  wire v3a61d83;
  wire v3777197;
  wire v3a6fa7a;
  wire v3a54c77;
  wire v3a70248;
  wire v3a6fc27;
  wire v372b6bc;
  wire d5bac5;
  wire v3a6294e;
  wire v3756e87;
  wire v374f87c;
  wire v3754f6b;
  wire v3a5a573;
  wire v3727f14;
  wire v3a67d3d;
  wire v37302fa;
  wire v3752f15;
  wire v3736107;
  wire v3763175;
  wire v3763f95;
  wire v3a70c39;
  wire v373380d;
  wire v3a5ce0f;
  wire v37470fc;
  wire v3a704cc;
  wire v3a6744e;
  wire v3255a34;
  wire v373b8c6;
  wire v37695c1;
  wire v3756ebf;
  wire v373d452;
  wire v376c9ee;
  wire v3a6dc08;
  wire v373f694;
  wire v3a70820;
  wire v3755783;
  wire v3744a67;
  wire v3a625a1;
  wire v37741bd;
  wire v3a6eec5;
  wire v3753f35;
  wire v375de66;
  wire v372b6a1;
  wire v3a64a7b;
  wire v37374bc;
  wire v3a70abe;
  wire v3760681;
  wire v3762b52;
  wire v3735f9a;
  wire v376d896;
  wire v3731974;
  wire v3735ad7;
  wire v3a6ed49;
  wire v3738c33;
  wire v3a6e221;
  wire v3722f65;
  wire v376dc26;
  wire v3735ed0;
  wire v2619b26;
  wire v3733383;
  wire v3733c46;
  wire v3778993;
  wire v3724621;
  wire v8f6518;
  wire v3a7058a;
  wire v372dcfb;
  wire v376b11a;
  wire v373dd77;
  wire v373dd66;
  wire v3a6f9d1;
  wire v375b05e;
  wire v3a6910c;
  wire v3731e7b;
  wire v3730fcd;
  wire v374e28d;
  wire v3a6ff23;
  wire v3a6230b;
  wire v37596de;
  wire v3a660f2;
  wire v35772c9;
  wire v372ca2a;
  wire v3a67f31;
  wire v37287d8;
  wire v3a6d1a5;
  wire v3766c8c;
  wire v37366d0;
  wire v3a646f8;
  wire v3a715d2;
  wire v380992b;
  wire v3a57b3c;
  wire v375b5b4;
  wire v372700a;
  wire v3a6f4f3;
  wire v3a7033a;
  wire v374d8ac;
  wire v3a5d259;
  wire v375cd50;
  wire v3724798;
  wire v3a70bc0;
  wire v3a62009;
  wire v3753dab;
  wire v3a6672b;
  wire v3753329;
  wire v3743966;
  wire v375e682;
  wire v3777adb;
  wire bbab81;
  wire v37751d9;
  wire v376d21d;
  wire v376086c;
  wire v3a6fa39;
  wire v37386cb;
  wire v377348f;
  wire v37485bd;
  wire v377b8ee;
  wire v373ef01;
  wire v35b7771;
  wire v374cd2c;
  wire v373f4a9;
  wire v3a53fb5;
  wire v37551eb;
  wire v3a70892;
  wire v3a6eefa;
  wire v3a63a21;
  wire v37644ff;
  wire v377d904;
  wire v3a66da0;
  wire v3753825;
  wire v3809cc0;
  wire v3a6f8b5;
  wire v374af1f;
  wire v37658de;
  wire v376fc23;
  wire v96c77f;
  wire v3a71150;
  wire v376bc75;
  wire v3a635eb;
  wire v3a70a6f;
  wire v3a6a41e;
  wire v3746c51;
  wire v377f01a;
  wire v37373ea;
  wire v3778834;
  wire v3777311;
  wire v3a70db0;
  wire v37269bf;
  wire v3a708f9;
  wire v3734291;
  wire v372f7d4;
  wire v3a5a5ec;
  wire v3a56642;
  wire v373165b;
  wire v3744806;
  wire v3a5d33e;
  wire v37605db;
  wire v37356f0;
  wire adf78a;
  wire v3722dfb;
  wire v37356ec;
  wire v37500db;
  wire v3730ffe;
  wire v3741a83;
  wire v3a6f1f5;
  wire v3a6194e;
  wire v3a54059;
  wire v3742c64;
  wire v3a67ab5;
  wire v3a5d417;
  wire v3a68057;
  wire v37c028d;
  wire v3a70f55;
  wire v3a70dcd;
  wire v3a654fb;
  wire v3759031;
  wire v372b726;
  wire v3a5ab9d;
  wire v377a393;
  wire v3a687be;
  wire v3742b9d;
  wire v3744da3;
  wire cda4f0;
  wire v373b983;
  wire v37592d6;
  wire v3754eb1;
  wire v3742122;
  wire v3a6dc60;
  wire v3777d6c;
  wire v3a63d0f;
  wire v3a663d6;
  wire v3a63ea7;
  wire v373f058;
  wire v3a711c0;
  wire v3a54264;
  wire v374e74c;
  wire v375d616;
  wire v376cfd9;
  wire v3a6fc1c;
  wire v3753838;
  wire v3a6eb4e;
  wire v3726fff;
  wire v3773729;
  wire v373abd0;
  wire v374608b;
  wire v3a6e152;
  wire v23fdbfc;
  wire v3746d92;
  wire v924b19;
  wire v3a70893;
  wire v3728c5b;
  wire v375928d;
  wire v373cd16;
  wire v8907fb;
  wire v373b5d8;
  wire v3a70666;
  wire v3726ea3;
  wire v3a71263;
  wire v3761181;
  wire v3a70edb;
  wire v377961f;
  wire v3a6669b;
  wire v3a6f4f8;
  wire v375c0cb;
  wire v3a59b5c;
  wire v3a6cb50;
  wire v3a5b037;
  wire v375355a;
  wire v37510fb;
  wire v3a67447;
  wire v37591bc;
  wire v3774399;
  wire v37685fe;
  wire v3767a2f;
  wire v3a63dbb;
  wire v3734af2;
  wire v3a5f495;
  wire v94faa4;
  wire v372b5f5;
  wire v374571a;
  wire v376029a;
  wire v3a70e03;
  wire v376e056;
  wire v3a70980;
  wire v373318b;
  wire v3a65711;
  wire v372dfba;
  wire v3a5740f;
  wire v3746a45;
  wire v3a6fa57;
  wire v374048c;
  wire v3a71159;
  wire v380987d;
  wire v3a581fb;
  wire v37296a5;
  wire v372d561;
  wire v3a6d8a9;
  wire v376af81;
  wire v377d23c;
  wire v3a667d2;
  wire v3a6ec0e;
  wire v1e37932;
  wire v35772a2;
  wire v3778425;
  wire v3748d3e;
  wire v372c502;
  wire v3a67967;
  wire v372b9e9;
  wire v37666bd;
  wire v3a70cc3;
  wire v3a714b1;
  wire v3774878;
  wire v3726339;
  wire v3743dfc;
  wire v372c8d1;
  wire v374da4a;
  wire v377928c;
  wire v37328b0;
  wire v37466d4;
  wire v37318da;
  wire v3763e88;
  wire v374102a;
  wire v3a71314;
  wire v377a985;
  wire v375fdb5;
  wire v3778a5a;
  wire v37551ac;
  wire v372e749;
  wire b4389d;
  wire v3a5e4e3;
  wire v373ee80;
  wire v3a5c473;
  wire v3729004;
  wire v37738ae;
  wire v3a704e5;
  wire v37793a6;
  wire v3779cd7;
  wire v37290af;
  wire v3775100;
  wire v3a65d33;
  wire v372a1b5;
  wire v3a6daed;
  wire v3a6a73a;
  wire v3748efb;
  wire v3767704;
  wire v3a70d29;
  wire v3768873;
  wire v3a56cfd;
  wire v3771d56;
  wire v3730b84;
  wire v3772c5a;
  wire v37281ca;
  wire v3754eb4;
  wire v3a6bde4;
  wire v3a6ebe8;
  wire v372eec6;
  wire v3a5902d;
  wire ade6f1;
  wire v37419f2;
  wire v377c72c;
  wire v3a53e46;
  wire v37611f5;
  wire v3a5e998;
  wire v3778627;
  wire v3a682e5;
  wire v37362e9;
  wire v37640e2;
  wire v955d7b;
  wire v377e851;
  wire v3a63cf3;
  wire v3746b91;
  wire v3765763;
  wire v3a61cb5;
  wire v3a5c93e;
  wire v376b28c;
  wire v3738f8a;
  wire v3a71560;
  wire v3728d1d;
  wire v37593c6;
  wire v3753e74;
  wire v3734930;
  wire v37407ef;
  wire v375377b;
  wire v3a6fb53;
  wire v3a58ef3;
  wire v3a7066b;
  wire v3728164;
  wire v3754a39;
  wire v3736012;
  wire v3a68dcb;
  wire v372c0cc;
  wire v3a5a5c4;
  wire v3735c06;
  wire v3768da7;
  wire v372cf1f;
  wire v3748a16;
  wire v37246d9;
  wire v3a71235;
  wire v376640a;
  wire v3a71535;
  wire v3a70f2e;
  wire v373eadd;
  wire v3a701b7;
  wire v3724488;
  wire v3773076;
  wire v3a704c4;
  wire v3a709eb;
  wire v3a6e69d;
  wire v3807472;
  wire v37631bf;
  wire a64c20;
  wire v376e661;
  wire v38072dc;
  wire v373c2e3;
  wire v37707b6;
  wire v375841a;
  wire v3a7050a;
  wire v3a70777;
  wire v374544f;
  wire v374e5ad;
  wire v3768082;
  wire v37506fe;
  wire v377d27f;
  wire v380913f;
  wire v376c79a;
  wire v3774f39;
  wire v376054c;
  wire v3757066;
  wire v3777ad7;
  wire v372b72d;
  wire v3a6cb96;
  wire v3a299ea;
  wire v37488cb;
  wire v3a66d2e;
  wire v373a782;
  wire v3a6b213;
  wire v3a70280;
  wire v374a075;
  wire v3750d8e;
  wire v3742e54;
  wire v3734f60;
  wire v375ed19;
  wire v3730d77;
  wire v3a70d7d;
  wire v3a7161f;
  wire v375eac3;
  wire v377c22b;
  wire v375a475;
  wire v3a670e4;
  wire v39a53eb;
  wire v375439c;
  wire v377c487;
  wire v3767dd2;
  wire v3a6eed1;
  wire d66718;
  wire v3a5ce54;
  wire v37503c2;
  wire v374ad23;
  wire v374704e;
  wire v3a689d1;
  wire v375c6cd;
  wire v3a71294;
  wire v372ef80;
  wire v3a6fb8d;
  wire v845765;
  wire v3765b5a;
  wire v3a70a33;
  wire v372e332;
  wire v8f9a63;
  wire v376e9e1;
  wire v3a5e5ec;
  wire v3a5fcc2;
  wire v37332b8;
  wire v38072bc;
  wire v3730d18;
  wire v374e99f;
  wire v3a5baf5;
  wire v3a6fe8d;
  wire v3a555ae;
  wire v3a62f14;
  wire v375dbda;
  wire v374aabf;
  wire v374a8e2;
  wire v3a70bf0;
  wire v377e5a6;
  wire v375eb37;
  wire v375067d;
  wire v3a6fa70;
  wire v3723089;
  wire v39748fd;
  wire v3a5a24d;
  wire v3a6f433;
  wire v3a5f3f0;
  wire v3770fff;
  wire v3a701b9;
  wire v3770ee4;
  wire v37770ae;
  wire v3a71140;
  wire v3772098;
  wire v374d313;
  wire v3a7110d;
  wire v37297ac;
  wire v3747804;
  wire v35b70ee;
  wire v3a548a0;
  wire a18d54;
  wire v3a6ded8;
  wire d23562;
  wire v3a6c4b3;
  wire v3a6a045;
  wire v3a64aa2;
  wire v377f6af;
  wire v374cb5e;
  wire v92bc1e;
  wire v3748443;
  wire v3a70c83;
  wire v375e459;
  wire v3759570;
  wire v3a6fcd4;
  wire v37531af;
  wire v374a3b2;
  wire v376142a;
  wire v3a57444;
  wire v3a63f66;
  wire v3769f7f;
  wire v3726b90;
  wire v375f888;
  wire v377db89;
  wire v3726634;
  wire v3a6fb1d;
  wire v3a6f069;
  wire v3a7133d;
  wire v3a6ae2d;
  wire v377938d;
  wire v377182c;
  wire v360d1cb;
  wire v3a69ac0;
  wire v375cd0c;
  wire v23fd970;
  wire v377e976;
  wire v3724994;
  wire v37328bf;
  wire v3a6f84d;
  wire v373178e;
  wire v372981e;
  wire v3746e79;
  wire v3725c02;
  wire v375b9c3;
  wire v3724200;
  wire v376cc23;
  wire v3a711a9;
  wire v377c29f;
  wire v3778ac6;
  wire v3a704a9;
  wire v3a569a9;
  wire v3770f96;
  wire v3a5c511;
  wire v376f980;
  wire v3a647b8;
  wire v373dcb6;
  wire v3770548;
  wire v3a6ffbe;
  wire v375803a;
  wire v3a7045c;
  wire v37693cf;
  wire v3769f88;
  wire v373343b;
  wire v3730cda;
  wire v37538e4;
  wire v3a712d6;
  wire v376011a;
  wire v3767650;
  wire v37784b9;
  wire v3761c1a;
  wire v375abc2;
  wire d3a479;
  wire v3a6f6cb;
  wire v373a1dc;
  wire v3776d72;
  wire v374410c;
  wire v3a6f632;
  wire v3a6fc35;
  wire v3756683;
  wire v3741435;
  wire v37693fe;
  wire v3739646;
  wire v3737dee;
  wire v3a70b2f;
  wire v3a60b1b;
  wire v3a5ad4f;
  wire v373b077;
  wire v3a6d951;
  wire v372fa0f;
  wire v3771fb3;
  wire v3a71567;
  wire v375ca6c;
  wire v3764dc2;
  wire v376ace9;
  wire v37490cb;
  wire v3730e71;
  wire v3a6f113;
  wire v373df21;
  wire v372456f;
  wire v372373f;
  wire v375c956;
  wire v374a63c;
  wire v3a6b18a;
  wire v373b197;
  wire v3a54a76;
  wire v3a6ff4c;
  wire v37565c7;
  wire v375f653;
  wire v375d80d;
  wire v3723ac5;
  wire v373d7fe;
  wire v3766df9;
  wire v374fac6;
  wire v3a6cdd4;
  wire v37314cb;
  wire v377a751;
  wire v3761af1;
  wire v375e551;
  wire v377de92;
  wire v375a116;
  wire v3a693af;
  wire v3a7028d;
  wire v3a70b55;
  wire v373b0be;
  wire v37577e7;
  wire v376db8f;
  wire v373510a;
  wire v3a5818a;
  wire v3762e13;
  wire v3754fd2;
  wire v376004c;
  wire v3a5e1a5;
  wire v37384fa;
  wire v374ab5b;
  wire v3a6f7f0;
  wire v374c718;
  wire v37709bb;
  wire v3741f69;
  wire v37756e8;
  wire v3a5e2b2;
  wire v377af98;
  wire v3a70799;
  wire v3730bf5;
  wire v373c441;
  wire v3757e28;
  wire v3a6ebaa;
  wire v3a6a3ac;
  wire aba148;
  wire v3a6935c;
  wire v3a6f54c;
  wire v372d30b;
  wire v375b9dc;
  wire v3a6f634;
  wire v37264cb;
  wire v3a704b6;
  wire v38079d5;
  wire v3774901;
  wire v3a70365;
  wire v3a5d6e3;
  wire v373be21;
  wire v3806f24;
  wire v91cdff;
  wire v3a699d3;
  wire v3a632f4;
  wire v3725994;
  wire v37669b4;
  wire v372b931;
  wire v3767abc;
  wire v373ead4;
  wire v3a5dbb7;
  wire v3766035;
  wire v3760bb4;
  wire v375323b;
  wire v373dafc;
  wire v3743698;
  wire v3a5da57;
  wire v37592f8;
  wire v377c842;
  wire v37244e7;
  wire v3743f47;
  wire v3743b79;
  wire v373cc51;
  wire v3735a71;
  wire v37654f4;
  wire v375e262;
  wire v377e419;
  wire v374a0ae;
  wire v37486e9;
  wire v3a70dfa;
  wire v37279dc;
  wire v39eb30a;
  wire v3779910;
  wire v3738e79;
  wire v3734bc3;
  wire v3745dc7;
  wire v3762949;
  wire v3768364;
  wire v3a6f723;
  wire v3a6f591;
  wire v375da95;
  wire v37386c5;
  wire v3723012;
  wire v3a5d830;
  wire v377a801;
  wire v3728f64;
  wire v375318f;
  wire v3a6dfc6;
  wire v3a6f8d1;
  wire v373a496;
  wire v3a6f4f5;
  wire v3a6fce0;
  wire v3a6f76a;
  wire v3775b3a;
  wire v373d091;
  wire v3a6fc65;
  wire v38097fc;
  wire v3746ac7;
  wire bf6063;
  wire v3a5be6a;
  wire v3a70f6b;
  wire v376f167;
  wire v372c00b;
  wire v3741022;
  wire v37c2b31;
  wire v374a99e;
  wire v3a63408;
  wire v3a2a144;
  wire v37782ff;
  wire v372d96e;
  wire v37254d2;
  wire v3779fbd;
  wire v3767fa5;
  wire v3a714e8;
  wire v3762f1a;
  wire v3a53e50;
  wire v374bb9c;
  wire v372d9ae;
  wire v372c8d0;
  wire v376f07c;
  wire v3740fc3;
  wire v3a6edfb;
  wire v8a0a3d;
  wire v3378fca;
  wire v3a668ec;
  wire v37655d3;
  wire v373d440;
  wire v373e10c;
  wire v375d1a6;
  wire v38065aa;
  wire v3a64087;
  wire v37513b7;
  wire v3a59d07;
  wire v3a6c0c5;
  wire v3a712c2;
  wire v2acaf41;
  wire v3a714b2;
  wire v374a3c5;
  wire v372672f;
  wire v376311f;
  wire v3760d74;
  wire v372cd91;
  wire v3768e79;
  wire v376ba4d;
  wire v3759cce;
  wire v3a6b3df;
  wire v3a6ff5c;
  wire v3772f26;
  wire v373f63e;
  wire v3724a2c;
  wire v37696a2;
  wire v374e124;
  wire v376b1a1;
  wire v37315af;
  wire v3809f61;
  wire v3762790;
  wire v377bdb2;
  wire v373dd82;
  wire v3a70f83;
  wire v39e9c6f;
  wire v372a7c9;
  wire v376cf85;
  wire v3a6d0ef;
  wire v372c577;
  wire v372396a;
  wire v372ae4c;
  wire v372de43;
  wire v3737ac6;
  wire v37721b2;
  wire v374b8ad;
  wire v377b68e;
  wire v373bb50;
  wire v3a6595f;
  wire v360d1b0;
  wire v37447e1;
  wire v3a703c0;
  wire v3a6d2df;
  wire v375d067;
  wire v377b5f6;
  wire v372fc9d;
  wire v3a66e5d;
  wire v37699c9;
  wire v376d240;
  wire v3a54393;
  wire v3a69e18;
  wire v37296f0;
  wire v374f485;
  wire v3a70d57;
  wire v3a70b8a;
  wire v3a70204;
  wire v3a6ff9e;
  wire v3a70fae;
  wire v373a8c0;
  wire v3a6b462;
  wire v3a6f73c;
  wire v3a70550;
  wire v37293e9;
  wire v3764eff;
  wire v2acb006;
  wire v3a64df4;
  wire v3728729;
  wire v3808e5b;
  wire v37358d5;
  wire v3a63198;
  wire v375e444;
  wire v3a6fe3d;
  wire v3774103;
  wire v3a6fc66;
  wire v3732d0f;
  wire v3a6fe59;
  wire v3776c87;
  wire v3a56a79;
  wire v3a5e784;
  wire v377997f;
  wire v3a6bff5;
  wire v3a62424;
  wire v3727626;
  wire v377b2b6;
  wire v375ced9;
  wire v3741f22;
  wire v37500ac;
  wire v375d12e;
  wire v3a548b2;
  wire v3748932;
  wire v3739417;
  wire v3a6f627;
  wire v377e9c4;
  wire v37629e2;
  wire v377cbcb;
  wire v373eb4d;
  wire v375e01c;
  wire v3743eae;
  wire v3779e45;
  wire v37396eb;
  wire v3a6999c;
  wire v37645ec;
  wire v3759470;
  wire v3730fd2;
  wire v3761bb6;
  wire v3764c57;
  wire v3779002;
  wire v3a645df;
  wire v375a02d;
  wire v3751faf;
  wire v3769d5c;
  wire v3a5d08a;
  wire v3a6e463;
  wire v3751e09;
  wire v37384ee;
  wire v3a6ef6d;
  wire v3a6f24c;
  wire v3a6487f;
  wire v3a6dd5a;
  wire v3a6d958;
  wire v37747f8;
  wire v37762cd;
  wire v3746efb;
  wire v3745452;
  wire v374760a;
  wire v37418ac;
  wire v3a6f687;
  wire v375913f;
  wire v3777a6c;
  wire v38064a2;
  wire v3a69146;
  wire v3723549;
  wire v374b0bc;
  wire v3a6af71;
  wire v3722e90;
  wire v3754e70;
  wire v3a647e3;
  wire v3743285;
  wire v373acc2;
  wire v375f423;
  wire v37248c1;
  wire v3a68407;
  wire v37317c4;
  wire v3a6e29c;
  wire v3a68b34;
  wire v3762886;
  wire v3739884;
  wire v3736913;
  wire v37538f5;
  wire v3742ce8;
  wire v376b5f8;
  wire v373243e;
  wire v2ff9268;
  wire v3730de2;
  wire v372d397;
  wire v375f3e2;
  wire v37711c8;
  wire v3a6ac7e;
  wire v3732d55;
  wire v372b4d7;
  wire v372b512;
  wire v3777a8c;
  wire v372a536;
  wire v3a64ad2;
  wire d1f2e2;
  wire v375d715;
  wire v3a70327;
  wire v37782af;
  wire v3779081;
  wire v374d402;
  wire v377cd6c;
  wire v3761d06;
  wire v3a6aa9f;
  wire v372b4a0;
  wire v3759a27;
  wire v3a68cec;
  wire v372ef39;
  wire v3725152;
  wire v3735c95;
  wire v3725fe1;
  wire v373ab4a;
  wire v372f09a;
  wire v3a6f1a4;
  wire v37331e7;
  wire v37600af;
  wire v3775442;
  wire v3777705;
  wire v360d1ca;
  wire v3a539ee;
  wire v376e139;
  wire v37526e0;
  wire v3a5c559;
  wire v373fc30;
  wire v377ae65;
  wire v3a6fff7;
  wire v3a6f485;
  wire v377a965;
  wire v3756b78;
  wire v3a702bb;
  wire v3739ca8;
  wire v3759842;
  wire v3744d52;
  wire v3a29803;
  wire v3a6f1c6;
  wire v3a56417;
  wire v376f148;
  wire v37675f4;
  wire v374b43d;
  wire v374b18c;
  wire v375c44b;
  wire v3a710aa;
  wire v373be9e;
  wire v3a701e7;
  wire v9644fd;
  wire v374d99a;
  wire v3730cc8;
  wire v3a6fa5e;
  wire v3a5a52a;
  wire v3a5f20d;
  wire v3a711ac;
  wire v3732b1e;
  wire v37643b5;
  wire v3728a77;
  wire v3730b6c;
  wire v376ea64;
  wire v377757b;
  wire v3a70408;
  wire v3a5cb5f;
  wire v3a5de50;
  wire v375c55a;
  wire v3a69765;
  wire v37c1a6f;
  wire v37536df;
  wire v3753edb;
  wire v37461ac;
  wire v376e364;
  wire v3757746;
  wire v3768eb1;
  wire v3737bc8;
  wire v373146d;
  wire v37308a8;
  wire v3a6f18f;
  wire v37699a0;
  wire v38070c1;
  wire v3a6faac;
  wire v3a6fb64;
  wire v3a5ef59;
  wire v37508a4;
  wire v3806b35;
  wire v3741401;
  wire v3a6f4ec;
  wire v373f42f;
  wire v372baaf;
  wire v3808c39;
  wire v376bc4b;
  wire v3a7036a;
  wire v375c463;
  wire v37474da;
  wire v3745b32;
  wire v3a5eac0;
  wire v373f23c;
  wire v3769f0f;
  wire v377ea59;
  wire v3732f03;
  wire v372818d;
  wire v373e0d3;
  wire v3a6fec9;
  wire v37672aa;
  wire v3a5cdc1;
  wire v3725058;
  wire v37230ec;
  wire v376bf83;
  wire b52e7d;
  wire v3a6fc33;
  wire v3a5b819;
  wire v3a6fdcb;
  wire v3726ee7;
  wire v1e37a8d;
  wire v3a7096d;
  wire v377316f;
  wire v3a6de60;
  wire v3a57422;
  wire v373b7be;
  wire v3725e33;
  wire v3741abd;
  wire v3731202;
  wire v3a5dffe;
  wire v3751b9a;
  wire v3764fad;
  wire v3a71279;
  wire v376fbe5;
  wire v3a6ffeb;
  wire v3a6f47d;
  wire v374e304;
  wire v3a6a557;
  wire v377bd77;
  wire v37656f7;
  wire v3a6f2fc;
  wire v3a71110;
  wire v37472b9;
  wire v3725d18;
  wire v37609e3;
  wire v3a5bda4;
  wire v3a6b68e;
  wire v3a7150f;
  wire d7f8bb;
  wire v373bf79;
  wire v3a5e46d;
  wire v3a6f696;
  wire v37603b3;
  wire v377e1d0;
  wire v3756149;
  wire v376306b;
  wire v3a6f02f;
  wire v376a936;
  wire v3a5e91b;
  wire v377aacd;
  wire v3a55d2f;
  wire v3a6ef6e;
  wire v3769f2f;
  wire v3748347;
  wire v3a6fa64;
  wire v3760101;
  wire v3778937;
  wire v37273d7;
  wire v3748bf9;
  wire v3775fae;
  wire v377389f;
  wire v3726f38;
  wire v3a5fe3c;
  wire v3a707e9;
  wire v373173e;
  wire v377dee0;
  wire v3a70649;
  wire v3a704f1;
  wire v3a6ba6a;
  wire v3a59275;
  wire v3a70bc7;
  wire v3757c37;
  wire v374b07a;
  wire v3a6fafa;
  wire v3a5a41c;
  wire v375461f;
  wire v3745a47;
  wire v3764d9e;
  wire v37706bf;
  wire v3a584bf;
  wire v37331b5;
  wire v3761932;
  wire v3758eae;
  wire v380749d;
  wire v373e09c;
  wire v3745e1f;
  wire v372372d;
  wire v1e3735b;
  wire v3730169;
  wire v374f979;
  wire v374e4bd;
  wire v3767b77;
  wire v373cd5d;
  wire v373a9ac;
  wire v3a71470;
  wire v376bc6b;
  wire v372993f;
  wire v3a6ffc3;
  wire v3776022;
  wire v37247f2;
  wire v3745ac6;
  wire v3a60f22;
  wire v3737571;
  wire v376c02d;
  wire v3a53f43;
  wire v3752943;
  wire c32250;
  wire v37501fd;
  wire v376b3bc;
  wire v376fb6b;
  wire v3731e0f;
  wire v3727293;
  wire v372d59e;
  wire v94e000;
  wire v375f8dd;
  wire v3a55b1d;
  wire v3a70ecb;
  wire v37759ff;
  wire v3a7005d;
  wire v3a7135e;
  wire a13040;
  wire v3a704e0;
  wire v3a6efd9;
  wire v3776756;
  wire v37247b3;
  wire v39eb5b0;
  wire v37241db;
  wire v374e210;
  wire v37625a0;
  wire v37480c6;
  wire v377af0b;
  wire v374ec37;
  wire v373c1ed;
  wire v3a551f9;
  wire v377eb00;
  wire v375e99f;
  wire v3a6f238;
  wire v377d310;
  wire v3739f07;
  wire v373c49e;
  wire v373929f;
  wire v3744794;
  wire v3a6968b;
  wire v373e113;
  wire v3a54ba5;
  wire v3a70c96;
  wire v3723f1a;
  wire v374b724;
  wire v3756559;
  wire v3777cae;
  wire v373bfd9;
  wire v37435a8;
  wire v37710c7;
  wire v3a63b57;
  wire v3772c7d;
  wire v37606b8;
  wire v3a7038e;
  wire v374f6a0;
  wire v3743ded;
  wire v3733f1c;
  wire v3a5f292;
  wire v37502d4;
  wire v3a7047f;
  wire v3a6f91a;
  wire v377defb;
  wire v3772ae7;
  wire v3728e25;
  wire v3759fe8;
  wire v376b5bc;
  wire v3a70055;
  wire v375cd00;
  wire v3761cdb;
  wire v3775eee;
  wire v3746f11;
  wire v3a545a7;
  wire v3a62ee2;
  wire v376eaed;
  wire v3a645ac;
  wire v374153d;
  wire v37738ca;
  wire v375ee43;
  wire v374db0f;
  wire v3729808;
  wire v3728d5a;
  wire v376c484;
  wire v3a64112;
  wire v37332c8;
  wire v3a6f481;
  wire v3a67bff;
  wire v3a7057f;
  wire v375a771;
  wire v3a70e85;
  wire v3764b3f;
  wire v37487a4;
  wire v3a6504e;
  wire v37686f3;
  wire v3a5c85c;
  wire v23fdad1;
  wire v35b779c;
  wire v3a70df6;
  wire v374464b;
  wire v375dfc6;
  wire v3a6ebd4;
  wire v3a5605f;
  wire v3a715df;
  wire v3a5f066;
  wire v3a5ec68;
  wire v3a701de;
  wire v3751253;
  wire v374d94e;
  wire v3755af9;
  wire v380971d;
  wire v373186a;
  wire v372a966;
  wire v3a69ead;
  wire v376d091;
  wire v37409c7;
  wire v9ae45c;
  wire v3a6fd4e;
  wire v3a619b8;
  wire v3769948;
  wire v3a57733;
  wire v3a6fab6;
  wire v3a557ea;
  wire v3a7131c;
  wire v3a6d809;
  wire v3a5d3af;
  wire v3742f28;
  wire v374113d;
  wire v3725dc4;
  wire v3a5cb45;
  wire v377459d;
  wire c3d672;
  wire v3737511;
  wire v375cb83;
  wire v3a67ee6;
  wire v375144b;
  wire v3a6ac2e;
  wire v3764898;
  wire v3769e94;
  wire a3cddb;
  wire v3a5ffbf;
  wire v372a51d;
  wire v3770d6d;
  wire v375d40b;
  wire v3a6f37c;
  wire v3742c52;
  wire v375d1fa;
  wire v3808ee4;
  wire v37612dd;
  wire v3732bc0;
  wire v377eba4;
  wire v3a6fd9d;
  wire v376cdf3;
  wire v376629a;
  wire v390071e;
  wire v3722dcd;
  wire v3a69c05;
  wire v3a68bb1;
  wire v37774e4;
  wire v3724c77;
  wire v37362d7;
  wire v3748e9d;
  wire v3a5bd58;
  wire v37c02a0;
  wire v375dd60;
  wire v373c5f5;
  wire v3768486;
  wire v374a7f0;
  wire v377722d;
  wire v37503c9;
  wire v3740dc6;
  wire v377312f;
  wire v3a70971;
  wire v374c190;
  wire v3a5a2a7;
  wire v3a7048d;
  wire v3745e72;
  wire v3754fac;
  wire v377535a;
  wire v3735d71;
  wire v376d658;
  wire v375ab6d;
  wire v3748792;
  wire v3772cf2;
  wire v3a6ebfd;
  wire v3737ada;
  wire v37470d6;
  wire v3a6bbed;
  wire v377b2ce;
  wire v37680af;
  wire v2acafff;
  wire v372538b;
  wire v1e37d2a;
  wire v3a6859a;
  wire v3a70f37;
  wire v3a6ebd3;
  wire v375924f;
  wire v377070e;
  wire v3770f75;
  wire v3a5c369;
  wire v3743a66;
  wire v3728196;
  wire v3779734;
  wire v3a67f60;
  wire v37444b4;
  wire v373ebf9;
  wire v373f95b;
  wire v3a6fce1;
  wire v3809127;
  wire v37386fb;
  wire v3a6fb66;
  wire v3a6fe9f;
  wire v3a6f3d9;
  wire v3745a0a;
  wire v372f9c3;
  wire v3a5adfd;
  wire v3a7081b;
  wire v3731ed2;
  wire v3757388;
  wire v3749408;
  wire a7f6c5;
  wire v37650e3;
  wire c7f1d0;
  wire v376eca3;
  wire v3a70219;
  wire v3740409;
  wire v3a6831c;
  wire dac346;
  wire v37719c6;
  wire v3772828;
  wire v2092aaa;
  wire v3775684;
  wire v3a6fa45;
  wire v3a625eb;
  wire v2acaecc;
  wire v3a70ef4;
  wire v3749831;
  wire v3733f28;
  wire d90332;
  wire v374672f;
  wire v3a6fa88;
  wire v3577392;
  wire v373f08d;
  wire v373d957;
  wire v3734c5c;
  wire v37247b5;
  wire v3762642;
  wire v3a6ea2b;
  wire v372e1bb;
  wire v3a6fcb5;
  wire v375e33e;
  wire v375fbef;
  wire v3a7046e;
  wire v377efe1;
  wire v37577ab;
  wire v3a613e6;
  wire v3729720;
  wire v3772229;
  wire v373f834;
  wire v3755d19;
  wire v37640dc;
  wire v37411c1;
  wire v373b571;
  wire v373bce1;
  wire v3752a43;
  wire v3a6f321;
  wire v3a70ed4;
  wire v3a695c2;
  wire bc3d4a;
  wire v1e38260;
  wire v377f2ec;
  wire v375d1d1;
  wire v374ad5f;
  wire v373bb90;
  wire v37790c6;
  wire v3a70448;
  wire v3722e04;
  wire v23fde61;
  wire v373e32c;
  wire v3763b37;
  wire v3a69a4c;
  wire v3736358;
  wire v376530c;
  wire v3a56c6d;
  wire v3770163;
  wire v3a5cd53;
  wire v376e9c5;
  wire v3751f46;
  wire v3a59b9e;
  wire v377e2e2;
  wire v3a66027;
  wire v3a6f975;
  wire v3779d16;
  wire v37578a2;
  wire v3a66279;
  wire v3769758;
  wire v3a5e020;
  wire v3a5ba97;
  wire v37280de;
  wire v3740e7d;
  wire v3a622f5;
  wire v3752523;
  wire v3747a41;
  wire v3735b31;
  wire v3a6851f;
  wire v3a5e5f3;
  wire v376ab5d;
  wire v3a58b4c;
  wire v3a6dc33;
  wire v3a6f898;
  wire v3a6fe71;
  wire v377f7e1;
  wire v3a6cd0f;
  wire v372339a;
  wire v373ffa0;
  wire v3a6f447;
  wire v376beaa;
  wire v3734f04;
  wire v3775219;
  wire v375f90e;
  wire v373db8f;
  wire v3a6770f;
  wire v37526cd;
  wire v3767463;
  wire v3a59d59;
  wire v3a595b8;
  wire v3763030;
  wire a97cd0;
  wire v3a59dd6;
  wire v37398ac;
  wire v374f654;
  wire v375a918;
  wire v3a6e857;
  wire v376944c;
  wire v3a5b581;
  wire v3a7083b;
  wire v3a665dd;
  wire v3760f1e;
  wire v375ff5c;
  wire v3a70ffb;
  wire v3a6f6b8;
  wire v3a62082;
  wire v377e288;
  wire v375eff3;
  wire v2092eaf;
  wire v3a70232;
  wire v374429f;
  wire v37480fe;
  wire v376f8bf;
  wire v3a600f3;
  wire v372ddf8;
  wire v325b5fd;
  wire v375556d;
  wire v3a7024b;
  wire v376a348;
  wire v3a6d48c;
  wire v3774a12;
  wire v3a66ada;
  wire v373ac67;
  wire v3749b62;
  wire v3a6f4de;
  wire v376ca93;
  wire v373a542;
  wire v377bd79;
  wire v3750714;
  wire v3a59545;
  wire v3756716;
  wire v3a57829;
  wire v3746e47;
  wire v3754f0f;
  wire v37336f0;
  wire v376773b;
  wire v375c482;
  wire v3a70a08;
  wire v3a5a34e;
  wire v373de53;
  wire v3733599;
  wire v372edd9;
  wire v3a706cb;
  wire v376a94e;
  wire v3a68c23;
  wire v37609d6;
  wire v3738fe2;
  wire v374b30b;
  wire v3742dce;
  wire v374880c;
  wire v377bea3;
  wire v37384a3;
  wire v3749a06;
  wire v3a6f2e5;
  wire v3742582;
  wire v372945c;
  wire v3a5749e;
  wire v376140e;
  wire v373db68;
  wire v3a5c653;
  wire v372e5a8;
  wire v3a6fabf;
  wire v373e6bc;
  wire v3756577;
  wire v373edd6;
  wire v3771ce8;
  wire v3a62c28;
  wire v372b390;
  wire v375fe02;
  wire aeff0f;
  wire v377e36c;
  wire v3a70c37;
  wire v3a6ef61;
  wire v376fdfb;
  wire v1e37938;
  wire v3756bd1;
  wire v376114f;
  wire v3758cc6;
  wire v376b934;
  wire v373b16e;
  wire v3a63004;
  wire v373859a;
  wire v377eb2d;
  wire v376ae07;
  wire v37431d8;
  wire v3a627a1;
  wire v98d1dc;
  wire v375c8c4;
  wire v375f354;
  wire v3767059;
  wire v3741e61;
  wire v377df77;
  wire v3a7056e;
  wire v3730d6e;
  wire v3a65dce;
  wire v37383b1;
  wire v37649e9;
  wire v3735049;
  wire v1e382f1;
  wire v3a66d74;
  wire v3735c5f;
  wire v377f298;
  wire v375ad90;
  wire v3761da2;
  wire v3a70898;
  wire v376b829;
  wire v37451c0;
  wire v3753b93;
  wire v3a6f511;
  wire v3a62841;
  wire v3738832;
  wire v35b70c9;
  wire v373d268;
  wire v3a66e63;
  wire v23fdbce;
  wire v3729beb;
  wire v3a6ff0c;
  wire v3a67f8e;
  wire v3a5a01b;
  wire v37677a3;
  wire v3a563d3;
  wire v3a700c7;
  wire v37527f2;
  wire v373676d;
  wire v3722bfc;
  wire v3a6f612;
  wire v3a5ff09;
  wire v37315da;
  wire v3737d2f;
  wire v374677f;
  wire v3808dcb;
  wire v372f5e5;
  wire v3a702c2;
  wire v372a20b;
  wire v3a6f87e;
  wire v2ff8f77;
  wire v3752987;
  wire v376b4a2;
  wire v3a71504;
  wire v3a71096;
  wire v37635d6;
  wire v3a6ef27;
  wire v37271e7;
  wire v37731d8;
  wire v3a6a4b0;
  wire v373e04e;
  wire v3735758;
  wire v372dd94;
  wire v37434bc;
  wire v37795e0;
  wire v3a71292;
  wire v376c898;
  wire c536d5;
  wire v3a5d2c5;
  wire v377ecf0;
  wire v3809ee4;
  wire v3a57e58;
  wire v372630c;
  wire v376e0cd;
  wire v372549f;
  wire beab35;
  wire v373e57b;
  wire v3a55e75;
  wire v3745e29;
  wire v3750883;
  wire v3763fec;
  wire v3a712d8;
  wire v3a7157b;
  wire v3751d7d;
  wire v3a6ab7f;
  wire v375be54;
  wire v3773b30;
  wire v3a652a2;
  wire v3729ed5;
  wire v3730df7;
  wire v3776084;
  wire v375101b;
  wire v376495c;
  wire v3a64bc8;
  wire v3774a7d;
  wire v372e083;
  wire v376d5a7;
  wire v3a71609;
  wire v375897d;
  wire v1e3780e;
  wire v3a5912f;
  wire v3a661f3;
  wire v375e0cc;
  wire dc571e;
  wire v372b627;
  wire b412f3;
  wire v380929f;
  wire v375c691;
  wire v376f0c2;
  wire v37261a6;
  wire v3747042;
  wire v374f31d;
  wire v3a715c5;
  wire v3a640d1;
  wire v372ad6d;
  wire v373c545;
  wire v37335ff;
  wire v3756f8c;
  wire v3769ec3;
  wire v374abbf;
  wire v37720ee;
  wire v38097ee;
  wire v37645bc;
  wire v372e95b;
  wire v3779f51;
  wire v372ec65;
  wire v3a66bc6;
  wire v3a68821;
  wire v3724600;
  wire v3767c92;
  wire v374b00b;
  wire v372b219;
  wire v3a6fd21;
  wire v3a7113f;
  wire v3a6f371;
  wire v3a6242b;
  wire v376f92c;
  wire v372dc77;
  wire v3a6fc76;
  wire v3a6731d;
  wire v37625d5;
  wire v9a641e;
  wire v3a6756b;
  wire v3770517;
  wire v3775303;
  wire v3739d51;
  wire v3a60c77;
  wire v374c6df;
  wire v3a6c23b;
  wire v3a5bf75;
  wire v37651cc;
  wire v3a7024a;
  wire v3a6f81f;
  wire v3722dba;
  wire v3a5a452;
  wire v375bf9a;
  wire v376c945;
  wire v37433d5;
  wire v3a6feab;
  wire v3772590;
  wire v3a63805;
  wire v3a710b4;
  wire v23fda7e;
  wire v1e3780d;
  wire v374a46d;
  wire v37381c2;
  wire v3a69973;
  wire v376945e;
  wire v3a69ce6;
  wire v380880f;
  wire v3a5d90d;
  wire v373b003;
  wire v37563eb;
  wire v3752407;
  wire v3a7042b;
  wire v3749435;
  wire v3a6ff25;
  wire v377378e;
  wire v3743da0;
  wire v3a70da3;
  wire v375941a;
  wire v3771555;
  wire v3a71581;
  wire v3770fb6;
  wire v3a6f5ea;
  wire v3a2975f;
  wire v373ea29;
  wire v377f06c;
  wire v3775d6e;
  wire v375e2de;
  wire v373cca3;
  wire v3a58218;
  wire v37406d2;
  wire v3730fc4;
  wire v37350c3;
  wire v3a6f6d1;
  wire v380881d;
  wire v3742efb;
  wire v37299dc;
  wire v3779c26;
  wire v3a63ef6;
  wire v3753ee5;
  wire v3a6f249;
  wire v3a706be;
  wire v374e58f;
  wire v377ab40;
  wire v3770578;
  wire v3a6f778;
  wire v3769cd3;
  wire v375a10d;
  wire v377030a;
  wire v3727acb;
  wire v3a573a7;
  wire v3a707a1;
  wire v373be40;
  wire v376648d;
  wire v372d0ad;
  wire v3770769;
  wire v3758e7b;
  wire v3a6fcb0;
  wire v3771e6f;
  wire v3a6e08c;
  wire v3a7097f;
  wire b79c3c;
  wire v3a7054d;
  wire v377d607;
  wire v3777c6f;
  wire v37670b6;
  wire v3a5f8d0;
  wire v3749907;
  wire v373c828;
  wire v3a5cb57;
  wire v377c38c;
  wire v372f9cf;
  wire v3a70fe6;
  wire v375fa7a;
  wire v3756203;
  wire v3a6c725;
  wire v3760740;
  wire v3a59905;
  wire v3728270;
  wire v375e5bb;
  wire v372b9d7;
  wire v37474e1;
  wire v375ca45;
  wire v374da21;
  wire v375ac23;
  wire v3768d11;
  wire v3a6b94f;
  wire v3a6a075;
  wire v3763c9c;
  wire v3730e01;
  wire v3a6e123;
  wire v3745075;
  wire v3733471;
  wire v37684c3;
  wire v374e4fd;
  wire v372f0c7;
  wire v376055d;
  wire v3737298;
  wire v37343bd;
  wire v3a693ca;
  wire v3776a3e;
  wire v3a5cff8;
  wire v3a5a8e6;
  wire v3a70f52;
  wire v3a6f094;
  wire v3a705ba;
  wire v376a9f5;
  wire v3760066;
  wire v374d41e;
  wire b0b0c6;
  wire v3770be6;
  wire v3758b25;
  wire v3742259;
  wire v373d78b;
  wire v3732dac;
  wire v3a6fcb9;
  wire v3a6f5fb;
  wire v372ec78;
  wire v3a6f359;
  wire v3a66606;
  wire v372ee06;
  wire v372dd09;
  wire v3776b2a;
  wire v377904f;
  wire v37638fe;
  wire v3775557;
  wire v3747994;
  wire v373a415;
  wire v3759ad6;
  wire v3731210;
  wire v3a56df7;
  wire v94e9e0;
  wire v374edd8;
  wire v3a70609;
  wire v3807601;
  wire v3a563c1;
  wire v3a69ba1;
  wire v372c298;
  wire v3a6f993;
  wire v9de657;
  wire v3748cce;
  wire v375f98a;
  wire v3736184;
  wire v3752cac;
  wire v37796c6;
  wire v372bcd0;
  wire v3a6c605;
  wire v3747de2;
  wire v3807ae8;
  wire v3a614fe;
  wire v3764daf;
  wire v3771a24;
  wire v375b22c;
  wire v3a70042;
  wire v3750296;
  wire v3a606a0;
  wire v3a612fa;
  wire v374183f;
  wire v3a683c1;
  wire v3a70528;
  wire v3a5544e;
  wire v3a6eee2;
  wire v3a62da7;
  wire v37284b7;
  wire cee4af;
  wire v372989d;
  wire v38073b0;
  wire v3732c51;
  wire v372c9b0;
  wire d03df7;
  wire v3754025;
  wire v372f49f;
  wire v375c652;
  wire v37604e1;
  wire v3735a77;
  wire v374e463;
  wire v3728bd6;
  wire v3a70e5f;
  wire v3767651;
  wire v376b86f;
  wire v375d889;
  wire v3a700b9;
  wire v3a6924d;
  wire v3a6dd8f;
  wire v377e031;
  wire v374b7b2;
  wire v373a8be;
  wire v3779015;
  wire v372af35;
  wire v372f039;
  wire v3a6eb9d;
  wire v37761d1;
  wire v3773b4b;
  wire v8ac439;
  wire v375c648;
  wire v3a58307;
  wire v376ef3d;
  wire v3a701cb;
  wire v37635a4;
  wire v3723d31;
  wire v3a7064e;
  wire v374fe2d;
  wire v3a657d3;
  wire v3a6f121;
  wire v3751539;
  wire v3769a2a;
  wire v3a63866;
  wire v3733e4f;
  wire v373c2e1;
  wire v377d3bf;
  wire v3a6fec5;
  wire v375aa44;
  wire bf2cd1;
  wire v375e566;
  wire v3737de9;
  wire v3751154;
  wire v37571d0;
  wire v3726a8d;
  wire v373a3b9;
  wire v3a63039;
  wire v3744daa;
  wire v3739c76;
  wire v3a58d7a;
  wire v374a343;
  wire v3731fae;
  wire v2acafaa;
  wire v3a701ad;
  wire v3807008;
  wire v3a6f90f;
  wire v3a556ab;
  wire v37782a8;
  wire v3735fb2;
  wire v3a565bc;
  wire v37256b3;
  wire v35b6dae;
  wire v3a5ec1a;
  wire v373cde5;
  wire v376d876;
  wire v3a6d34c;
  wire v3a6f3dc;
  wire v3a6f737;
  wire v3761d7e;
  wire v3756960;
  wire v3a6fc1a;
  wire v375f862;
  wire v3748446;
  wire v37262ad;
  wire v3763f8e;
  wire v3a70236;
  wire v3758c07;
  wire v3a6b5ea;
  wire v37c01ec;
  wire v3a6f072;
  wire v37677e2;
  wire v377346e;
  wire v3a68a8b;
  wire v3a6f7a3;
  wire v374e55d;
  wire v37376dd;
  wire v38076cf;
  wire v372faf3;
  wire v377cb0b;
  wire v3a63cce;
  wire v373024e;
  wire v3a60815;
  wire v376dc03;
  wire v3762fd0;
  wire v374ef97;
  wire v3740233;
  wire v376f920;
  wire v3765d5e;
  wire v3732c6a;
  wire v373443d;
  wire v375d43d;
  wire v374c91a;
  wire v37793c8;
  wire v373d41a;
  wire v3a70948;
  wire v3752a7a;
  wire v3747824;
  wire v3a6f8bd;
  wire v376a11d;
  wire v3a5b6b0;
  wire v3a5e035;
  wire v3744cf1;
  wire v374215e;
  wire v3a7060c;
  wire bdb538;
  wire v373d5f4;
  wire v3a6de06;
  wire v372c92c;
  wire v3a6cf91;
  wire v3a69036;
  wire v3806f1f;
  wire v374c6de;
  wire v3a5b0f5;
  wire v376a662;
  wire v3a6f3b5;
  wire v3a7151b;
  wire v2acaf4f;
  wire v1e37d35;
  wire v3a6f8a8;
  wire v377c5f8;
  wire v3764ec5;
  wire v23fdadd;
  wire v3a6abcb;
  wire v375a269;
  wire v3756f41;
  wire v3a5b3e6;
  wire v3a61d67;
  wire v373e2aa;
  wire v3a6233b;
  wire v3a5907a;
  wire v375bde1;
  wire v37543c2;
  wire v37275a7;
  wire v3761611;
  wire v37417f6;
  wire v376fa80;
  wire v2acaeb7;
  wire v3a663c7;
  wire v3a59b5f;
  wire v3a6eab0;
  wire v2aca789;
  wire v3a71261;
  wire v9e2dd1;
  wire v3741c76;
  wire v3748451;
  wire v372a246;
  wire v3a6ab55;
  wire v3725c60;
  wire v377ef0b;
  wire v3722be8;
  wire v3a6f9a0;
  wire v3a6fed2;
  wire v376ed1f;
  wire v3749e96;
  wire v37710d4;
  wire v3724581;
  wire v3a5d448;
  wire v3a71378;
  wire v3a6fe0a;
  wire v3a5d836;
  wire v376beed;
  wire v3a68728;
  wire v373cddc;
  wire v377e283;
  wire v37721cb;
  wire v3778ab3;
  wire v3a53c87;
  wire v3a71251;
  wire v373a263;
  wire v37694a0;
  wire v3a68915;
  wire v3a6cdcd;
  wire v373dafe;
  wire v3a68825;
  wire v375cd8c;
  wire v37615c5;
  wire v3724d99;
  wire v3723211;
  wire v3774b12;
  wire v3a64b9b;
  wire v3a574bf;
  wire v372e466;
  wire v3a703a7;
  wire v3759265;
  wire v37350a4;
  wire v3776b93;
  wire v3761cd5;
  wire v3a68d70;
  wire v377ed6c;
  wire v3a5a226;
  wire v3a70682;
  wire v375818a;
  wire v3771b8a;
  wire v37346fe;
  wire v3a5bc5f;
  wire d383e7;
  wire v3726eb4;
  wire v3a6fb17;
  wire v372b9a2;
  wire v377225c;
  wire v3a6fdbf;
  wire v37314f0;
  wire v3a69674;
  wire v3764334;
  wire v3a624d7;
  wire v3747d3d;
  wire v373da33;
  wire v372316a;
  wire v3a6570f;
  wire v3723f0c;
  wire v3778d9d;
  wire v37637db;
  wire v39a5382;
  wire v3769061;
  wire v37747fc;
  wire v3765a43;
  wire v375b269;
  wire v376b1bf;
  wire v3a70512;
  wire v3777962;
  wire v37331ef;
  wire v3a65e52;
  wire v20930c2;
  wire v375fdf5;
  wire v37318d7;
  wire v377a577;
  wire v3a68c7d;
  wire v3a708b6;
  wire v8e4471;
  wire v3577388;
  wire v3760af0;
  wire v3a618b7;
  wire v375978a;
  wire v374a95d;
  wire v3a715ab;
  wire v375f30d;
  wire v37400bc;
  wire v3776f7f;
  wire v37473a3;
  wire v3a6fa3f;
  wire v3a71293;
  wire v374f820;
  wire v3a59a2b;
  wire v3758a23;
  wire v3a5da31;
  wire v3778595;
  wire v3a5520a;
  wire v3a55b16;
  wire v37739af;
  wire v376c94b;
  wire v373705f;
  wire v3a59e1b;
  wire v373e679;
  wire v374e402;
  wire v37252ee;
  wire v3a708a0;
  wire v3761915;
  wire v3a57b46;
  wire v376ffb4;
  wire v375ebc3;
  wire v3a6f48e;
  wire v3a70052;
  wire v373bdd9;
  wire v3778355;
  wire v3735cb3;
  wire v3a673d6;
  wire v3725bf4;
  wire v37282ac;
  wire v37724f9;
  wire v373f79d;
  wire v376eb1f;
  wire v3a6c0fb;
  wire v3751b42;
  wire v3a6f75c;
  wire v209312a;
  wire v3a5a72a;
  wire v37331df;
  wire v3a60c86;
  wire v376c2da;
  wire v3744640;
  wire v374b923;
  wire v3754c8d;
  wire v3a6f68f;
  wire v377a461;
  wire v3749caf;
  wire v374518b;
  wire v3a5ec7a;
  wire v372cac6;
  wire v3a6f195;
  wire v373a791;
  wire v3a6f8b9;
  wire v3756202;
  wire v3a5971e;
  wire v377ce47;
  wire d2ccfa;
  wire v3743c35;
  wire v3738f1b;
  wire v3a7135a;
  wire v374e032;
  wire v3751022;
  wire v3a5aac9;
  wire v3a705df;
  wire v3a57c78;
  wire v23fe20c;
  wire v3a660c0;
  wire v3a6602e;
  wire v372995e;
  wire v9ed0ba;
  wire v3a6b090;
  wire v377ca40;
  wire v3a7016b;
  wire v3a708fb;
  wire v3a569c8;
  wire v3a711d5;
  wire v372e96f;
  wire v3a6f6b9;
  wire v3807afa;
  wire v37258c9;
  wire v3806fa6;
  wire v3776a27;
  wire v3a7145a;
  wire v3a65436;
  wire v3a5a1ba;
  wire v37381eb;
  wire v377ca8e;
  wire v374fe39;
  wire v3734916;
  wire v37644ce;
  wire v376dc91;
  wire v372a954;
  wire v377aa81;
  wire v3728526;
  wire v3753e49;
  wire v375aaf3;
  wire v374eda5;
  wire v2925ca9;
  wire v37470c7;
  wire v3724f5d;
  wire v375a32c;
  wire v3a70363;
  wire v3a7091c;
  wire v376d328;
  wire v3a61895;
  wire v3762934;
  wire v3a70057;
  wire v3a5e4f4;
  wire v3a6fbca;
  wire v372ea9b;
  wire v3379430;
  wire v3a6fc0f;
  wire v375b9b2;
  wire v375f3f4;
  wire v3766ff1;
  wire v3744c95;
  wire v3730bb7;
  wire v3a70a68;
  wire v372ae0b;
  wire v3a654c4;
  wire v3722a0a;
  wire v375a2b5;
  wire v376faad;
  wire v3a6f42c;
  wire v377ce30;
  wire v3751073;
  wire v3a61739;
  wire v3770bd5;
  wire v372ddde;
  wire v377193a;
  wire v3a6f043;
  wire v3a5db41;
  wire v377e57f;
  wire v37788fc;
  wire v3a70f7f;
  wire v377af47;
  wire v3a5ad12;
  wire v3771042;
  wire v3a6f849;
  wire a12203;
  wire v373ee70;
  wire v3a6fd82;
  wire v375d707;
  wire v3a71429;
  wire v373d34e;
  wire v37299e2;
  wire v3a6802b;
  wire v3733be1;
  wire v3767d4b;
  wire v3764568;
  wire v3a57912;
  wire v374bc9c;
  wire v3a70950;
  wire v3767e79;
  wire v372b3ca;
  wire v3a5551b;
  wire v3800ee4;
  wire v37608ba;
  wire v98068b;
  wire v3779da3;
  wire v372c334;
  wire v3a70737;
  wire v3a70f01;
  wire v376efdb;
  wire v3734913;
  wire v374890e;
  wire v375b534;
  wire v3a70b74;
  wire v3a6ec1f;
  wire v3a6f9b3;
  wire v3a61e10;
  wire v3722da3;
  wire v37456d2;
  wire v3738cab;
  wire v376fd9a;
  wire v374b95f;
  wire v37368df;
  wire v3727165;
  wire v3a647f3;
  wire v377dae6;
  wire v3752c99;
  wire v376455c;
  wire v374cd51;
  wire v3760d54;
  wire v373bf6a;
  wire v373ca8d;
  wire v3a71387;
  wire v3749e33;
  wire v3770be3;
  wire v37658f5;
  wire v3a6b20a;
  wire v377e9cd;
  wire v3a5a52d;
  wire v376c573;
  wire v3776352;
  wire v372871c;
  wire v3a6fb23;
  wire v3a61e9f;
  wire v37360c8;
  wire v3a62d1c;
  wire v3740b8b;
  wire v376c1f7;
  wire v3723555;
  wire v2678c95;
  wire v3a63690;
  wire v3767258;
  wire v3a6eec9;
  wire v374813d;
  wire v3755bb0;
  wire v374d810;
  wire v377d8eb;
  wire v38063dd;
  wire v372807c;
  wire v372b5a8;
  wire v376865d;
  wire v3745366;
  wire v3a60a75;
  wire v3752869;
  wire v3a5c3ba;
  wire v3733174;
  wire v952f44;
  wire v374db48;
  wire v375e574;
  wire v3736894;
  wire v375a9c1;
  wire v3775adf;
  wire v373f247;
  wire v376d488;
  wire v37506d6;
  wire v37785b8;
  wire v3a671de;
  wire v3732f8d;
  wire v37427f8;
  wire v37479ef;
  wire v3769283;
  wire v23fe03a;
  wire v377bbd1;
  wire v3750f4b;
  wire v3767e15;
  wire v3808dca;
  wire v3a66476;
  wire v39a4db0;
  wire v372475e;
  wire v375a65f;
  wire v3738ad8;
  wire v3738c0a;
  wire v1e37c38;
  wire v3a6fd4a;
  wire v3734fa5;
  wire v3a6fcb8;
  wire v372d70c;
  wire v3a6f192;
  wire v3a647df;
  wire v3a6eb62;
  wire v373f5d3;
  wire v3a68c1c;
  wire v3732246;
  wire v372dddc;
  wire v37773fa;
  wire v37463a6;
  wire v3758a10;
  wire v372f91d;
  wire v37331ff;
  wire v377d742;
  wire v377c261;
  wire v3a608fe;
  wire v3a68c72;
  wire v372449f;
  wire v3a5fbd6;
  wire v3763bb8;
  wire v372ea02;
  wire v372a49a;
  wire v372b418;
  wire v3a5fd18;
  wire v3741872;
  wire v3745d0a;
  wire v3a6addc;
  wire v377fab4;
  wire v375c358;
  wire v3732871;
  wire v3a70421;
  wire v3738ab6;
  wire v39eb3d2;
  wire v3726ba5;
  wire v3a71580;
  wire v374fa8c;
  wire v3a63c3b;
  wire v3a6fc9c;
  wire v3a60147;
  wire v3a60594;
  wire v372f04d;
  wire v3a5d438;
  wire v3762079;
  wire v3a5fe51;
  wire v3a6ff2e;
  wire v373498b;
  wire v3a6f9e3;
  wire v37623dd;
  wire v377135e;
  wire v375aa2d;
  wire v37611c3;
  wire v3a6ef75;
  wire v3730e54;
  wire v3a5ca44;
  wire v374448e;
  wire v3768358;
  wire v375301b;
  wire v3731599;
  wire v3727849;
  wire v3724c35;
  wire v37353b5;
  wire v375d9a7;
  wire v372a902;
  wire v3a6b8d8;
  wire v3a58d63;
  wire v3a709e5;
  wire v372a674;
  wire db1dc4;
  wire v3a6113b;
  wire v3a5a36d;
  wire v3806e88;
  wire v3a61120;
  wire v372e03f;
  wire v3a70d86;
  wire v377c258;
  wire v3a57d2f;
  wire v377dae8;
  wire v373a3fa;
  wire v374ac8c;
  wire v373935b;
  wire v376e513;
  wire v3a714fc;
  wire v3a6616c;
  wire v3a71410;
  wire v376245d;
  wire v372adc8;
  wire v37520a9;
  wire v3a7022e;
  wire v3a71632;
  wire v3a7033b;
  wire a2e8c8;
  wire v3a71092;
  wire v3a6ad00;
  wire v374f968;
  wire v374f397;
  wire v37301dd;
  wire v3a58ea7;
  wire v3a5b1a3;
  wire v37639b1;
  wire v3a6f0bd;
  wire v3a682f0;
  wire v3764049;
  wire v375a6a7;
  wire v3a715c3;
  wire v3a705e4;
  wire v37567ef;
  wire v373dd7f;
  wire v372aa71;
  wire v375abdb;
  wire v377c690;
  wire v3a5ad83;
  wire v3a54b2b;
  wire v3a6f414;
  wire v3a714a3;
  wire v3a6fa17;
  wire v372b8da;
  wire v3756c2e;
  wire v373ae84;
  wire v376d078;
  wire v3a6e581;
  wire v3754eca;
  wire v3743fea;
  wire v3a5567a;
  wire v377fb09;
  wire v376e580;
  wire v373cae8;
  wire v37247b2;
  wire v37266a0;
  wire v3a6f73f;
  wire v375fbc6;
  wire v3759a7f;
  wire v3779988;
  wire v3a70347;
  wire v375c062;
  wire v376704f;
  wire v3a6f2b7;
  wire v3a6f8b7;
  wire v3756b7b;
  wire v3a63dde;
  wire v3a6f8ce;
  wire v3775da1;
  wire v373cedb;
  wire v37769d5;
  wire v3a6d003;
  wire v372a599;
  wire v3a70e80;
  wire v372bb35;
  wire v374f832;
  wire v3741816;
  wire v3a62959;
  wire v3a6fc6b;
  wire v37471c2;
  wire v3752552;
  wire v374f003;
  wire v37333a4;
  wire v375a878;
  wire v3733239;
  wire v374802b;
  wire v3a674c9;
  wire v3a6f590;
  wire v3a643ef;
  wire v3732d3e;
  wire v375415d;
  wire v373d26a;
  wire a36719;
  wire v3773a25;
  wire v3772140;
  wire v3734aa5;
  wire v37586ed;
  wire v3a712d2;
  wire v375e051;
  wire v3776a2e;
  wire v3a65155;
  wire v3a6fb6f;
  wire v3a664ed;
  wire v38071c7;
  wire v3a6f6f0;
  wire v3738f36;
  wire v37229db;
  wire v38063ce;
  wire v3a5ddef;
  wire v37688bf;
  wire v3731839;
  wire v374d163;
  wire d973ae;
  wire v376e0b5;
  wire v3a60b69;
  wire v377a2b2;
  wire v375055f;
  wire v3a6effd;
  wire v3738aa6;
  wire v3724bdd;
  wire v892398;
  wire v3a63fd2;
  wire v3a6f292;
  wire v3760592;
  wire a94d63;
  wire v3729180;
  wire v37758e6;
  wire v3761947;
  wire v373a327;
  wire v3749ca6;
  wire v3a5e3d1;
  wire v3a6167d;
  wire v3a5f6c2;
  wire v37438ba;
  wire v3a5bfbd;
  wire v377d23d;
  wire v37303f0;
  wire v37273f4;
  wire v3740627;
  wire v373b7b5;
  wire v3773c5d;
  wire v3a71167;
  wire v37649a5;
  wire v3763502;
  wire v3760ca3;
  wire v3741bd4;
  wire v3739a33;
  wire v3a6fbcc;
  wire v3776135;
  wire v3a53b76;
  wire v3a675dc;
  wire v37736b4;
  wire v37586e4;
  wire v3a6f93b;
  wire v3747389;
  wire v3a711d1;
  wire v3a715cd;
  wire v373b0b2;
  wire v3763d10;
  wire v375cdee;
  wire v3a70297;
  wire v3a62b8d;
  wire v3a7051a;
  wire v377d4a0;
  wire v374f20c;
  wire v374383b;
  wire v3a65596;
  wire v3a70293;
  wire v3a70c61;
  wire v3a62ed6;
  wire v3a6ebdb;
  wire v3a6eb94;
  wire v3749e5a;
  wire v37711e2;
  wire v3778345;
  wire v3769a36;
  wire v372b4c0;
  wire v374776e;
  wire v373e6d2;
  wire v3733ec6;
  wire v3a622c0;
  wire v374cda5;
  wire v35b70a0;
  wire v37241cc;
  wire v372618d;
  wire v3758adb;
  wire v3743d21;
  wire v374edff;
  wire v376e65d;
  wire v374f658;
  wire v372f2fe;
  wire v3741e5c;
  wire v374a23b;
  wire v3769bec;
  wire v3a70ed6;
  wire v37642f9;
  wire v377c147;
  wire v3750e83;
  wire v3731666;
  wire v3a6fcc0;
  wire v3a7032d;
  wire v3a70a3c;
  wire v3a7000e;
  wire v3733be0;
  wire v373a374;
  wire v377636a;
  wire v3749586;
  wire v3a707ae;
  wire v3757598;
  wire v3724887;
  wire v37591ae;
  wire v3748858;
  wire v372424e;
  wire v372dcff;
  wire v3a53b8b;
  wire v3763a4a;
  wire v3726521;
  wire v3743b2c;
  wire v373940c;
  wire v3808eb8;
  wire v37584fe;
  wire v3a58a16;
  wire v3a60882;
  wire v3a63d63;
  wire v37747b4;
  wire v375f0ba;
  wire v3777e69;
  wire v3a70d94;
  wire v374f5e0;
  wire v3a705e2;
  wire v373240c;
  wire v3723988;
  wire v3a71149;
  wire v3a6ed27;
  wire v3a6261c;
  wire v3770338;
  wire v373de83;
  wire v375808f;
  wire v37717d0;
  wire v373e475;
  wire v3a5d96d;
  wire v374819d;
  wire v3a6906e;
  wire v376af64;
  wire v3a674fd;
  wire v3a67bbd;
  wire v37743e0;
  wire v374558a;
  wire v3732688;
  wire v3774cc2;
  wire v3a59d80;
  wire v37637ef;
  wire v373104a;
  wire v375d3bc;
  wire v374fa4f;
  wire v3a631b4;
  wire v3a5e95a;
  wire v3a6c066;
  wire v3a6ecd9;
  wire v376c569;
  wire v3a6f4c5;
  wire v377e867;
  wire v372ba4d;
  wire v3a71630;
  wire v3755b5e;
  wire v3a6f2ef;
  wire v3a6de33;
  wire v37764a5;
  wire v3735826;
  wire v375d635;
  wire v373f661;
  wire v3a58fef;
  wire v3760e7b;
  wire v375a7fc;
  wire v3776c09;
  wire v3a708af;
  wire v373e369;
  wire v375e948;
  wire v374a19d;
  wire v373fad7;
  wire v3a66d94;
  wire v37549eb;
  wire v377c2ce;
  wire v3773a84;
  wire v373fe10;
  wire v3754cf4;
  wire v3751af0;
  wire v377d7db;
  wire v3778967;
  wire v374ba65;
  wire v3a710d2;
  wire v3a6f6ba;
  wire v3a6cef4;
  wire cf1ae7;
  wire v3724f9c;
  wire v372bcbc;
  wire v39a4dd4;
  wire v3a5ee99;
  wire v374125a;
  wire v373fb30;
  wire v3a66f0d;
  wire v37704dc;
  wire v3737e2d;
  wire v377e8e4;
  wire v37676c3;
  wire v3a6009a;
  wire v377444e;
  wire v3a69547;
  wire v377c0d5;
  wire v3a6fd66;
  wire v3a63bb7;
  wire v3a6ab5e;
  wire v377a6fe;
  wire v372f0bb;
  wire v3a70b8f;
  wire v3807b27;
  wire v375c423;
  wire v3754fc8;
  wire v375af57;
  wire v3731320;
  wire v3776592;
  wire v3727d95;
  wire v372ff2c;
  wire v37511c0;
  wire v3a6f9ca;
  wire v3a6505b;
  wire v37703c6;
  wire v3758c62;
  wire v3a6eeca;
  wire v3a69b5c;
  wire v3a6f70c;
  wire v3757f01;
  wire v3a71377;
  wire v372e213;
  wire v3768c08;
  wire v3772a4f;
  wire v375d849;
  wire v3a5b855;
  wire v3a5cd4c;
  wire v2889706;
  wire v3a628cf;
  wire v3a610f8;
  wire v3740352;
  wire v374fe63;
  wire v3a6eb7d;
  wire v3725626;
  wire v3a712c5;
  wire v3a7113a;
  wire v377cf67;
  wire v376f48d;
  wire v3a5cc17;
  wire v3809583;
  wire v377db21;
  wire v37480a7;
  wire cb9412;
  wire v3a63260;
  wire v37263bc;
  wire v37556cb;
  wire v3732f66;
  wire ac438c;
  wire v3806b87;
  wire v37391b4;
  wire v3a62539;
  wire v3734c7e;
  wire v3a57156;
  wire v3a6a713;
  wire v3765265;
  wire v3758180;
  wire v3726bb8;
  wire v37355db;
  wire v3a5b6ca;
  wire v2092bae;
  wire v3a68240;
  wire v3733dd3;
  wire v3775aef;
  wire v375b8b9;
  wire v377ceea;
  wire v374c75e;
  wire v3a70f1c;
  wire v3a5fde5;
  wire v3768dd8;
  wire v3a70c28;
  wire v3a6f7f2;
  wire v3a61bef;
  wire v373fb40;
  wire v372cc3d;
  wire v374a36a;
  wire v3a6eff3;
  wire v37295ce;
  wire v374b035;
  wire v376b2a3;
  wire v37603d4;
  wire v3808d47;
  wire v3a5f4e0;
  wire v3a7087d;
  wire v372e426;
  wire v3730dc4;
  wire v3763fdc;
  wire v3a6f75d;
  wire v3724733;
  wire v374602f;
  wire v374c007;
  wire v372b31a;
  wire v373d245;
  wire v3a54ac1;
  wire v3771cf0;
  wire v376157e;
  wire v3a656d0;
  wire v37776b6;
  wire v3773fd1;
  wire v37711cc;
  wire v37700b9;
  wire v372d490;
  wire v3a6f46a;
  wire v377dc87;
  wire v3a67a06;
  wire v3a70cdb;
  wire v37502d9;
  wire v377222b;
  wire v3777d41;
  wire v3a709c1;
  wire v3a71400;
  wire v3a5d717;
  wire v3776be1;
  wire v37297b2;
  wire v3a68ad8;
  wire v2ff8f0a;
  wire v376022e;
  wire v3751338;
  wire v3a5e070;
  wire v3760799;
  wire v372bd23;
  wire v375265e;
  wire v3731c6f;
  wire v3a6fbd9;
  wire v3a6f3f9;
  wire v3a6cb19;
  wire v3739d45;
  wire v375ecf5;
  wire v376dba6;
  wire v3741f3c;
  wire v3a6c717;
  wire v3a6fcda;
  wire v3a71018;
  wire v3739892;
  wire v3a714e4;
  wire v3a5aa3a;
  wire v3775fb0;
  wire v3a6f38c;
  wire v3a53fa4;
  wire v3750aea;
  wire v3a5f991;
  wire v3743e29;
  wire v3742033;
  wire v372a4c4;
  wire v3a6f72a;
  wire v374e19c;
  wire v375d4f9;
  wire v375f98c;
  wire v37404b3;
  wire v375791b;
  wire v3a6ebb3;
  wire v374974e;
  wire v3744b3d;
  wire a6f8c7;
  wire v37bfcae;
  wire v3756bc2;
  wire v374551a;
  wire v373e1a6;
  wire v3a58b28;
  wire v374638c;
  wire v3756883;
  wire v38092e6;
  wire v375ceff;
  wire v3738114;
  wire v376fe96;
  wire v3a55d7c;
  wire v3765474;
  wire v37539bc;
  wire v3a5de8f;
  wire v3a6da5a;
  wire v375361a;
  wire v375783c;
  wire v37401ce;
  wire v20930ad;
  wire v3772c21;
  wire v3764c8a;
  wire v3a6f309;
  wire v37406e8;
  wire v3a7062d;
  wire v372476f;
  wire v3731beb;
  wire v37771ed;
  wire v3a6fd2d;
  wire v39ea0c5;
  wire v377d1cd;
  wire v3a70ac9;
  wire v37592a3;
  wire v37513fa;
  wire v3a7139c;
  wire aca44a;
  wire v3a6eaf3;
  wire v3768985;
  wire v3727369;
  wire v372aadd;
  wire v3737ca3;
  wire v3a5afe8;
  wire v3a6db06;
  wire v3a6f940;
  wire v37281d0;
  wire v3a69c6f;
  wire v3a714c6;
  wire v3a711c9;
  wire v3a638e9;
  wire v375ff98;
  wire v3a713ae;
  wire v3a5be72;
  wire v3757f9b;
  wire v372526e;
  wire v373b666;
  wire v3a6817a;
  wire v3763aec;
  wire v3a706e4;
  wire v375d77d;
  wire v3a64483;
  wire v3751100;
  wire v376604f;
  wire v375f147;
  wire v3a59461;
  wire v3a71503;
  wire v3a65053;
  wire v3a6297f;
  wire v3746404;
  wire v375635b;
  wire v374ac3f;
  wire v3a6ce42;
  wire v372eec5;
  wire v3730ad2;
  wire v8b51d2;
  wire v374000d;
  wire v372a6c8;
  wire v3749381;
  wire v373c5a6;
  wire v372bdcf;
  wire v3a6f1ea;
  wire v3a6eec8;
  wire v3761bd6;
  wire v377a681;
  wire v372641e;
  wire v3a712e4;
  wire v3a6eb19;
  wire v3a63c12;
  wire v37796e9;
  wire v376b7e1;
  wire v375133a;
  wire v3769090;
  wire v3808db6;
  wire v373d0d3;
  wire v3a5514a;
  wire v375df5a;
  wire v37239a5;
  wire v3a6bce9;
  wire v3740742;
  wire v377dc82;
  wire v372ea5d;
  wire v3744b87;
  wire v37335e0;
  wire v3a54952;
  wire v23fd9af;
  wire v37510d7;
  wire v3a5a8ce;
  wire v372ff6d;
  wire v3a59c91;
  wire v37520d9;
  wire v3735331;
  wire v3a62ad5;
  wire v3742953;
  wire v37691e2;
  wire v375a5e3;
  wire v3a574d6;
  wire v3a6ff69;
  wire v373ecb2;
  wire v3754018;
  wire v375624e;
  wire a8fef2;
  wire v3a53904;
  wire v37730ff;
  wire v37371df;
  wire v37531fd;
  wire v3a6fe4e;
  wire v3754685;
  wire v373c526;
  wire v3a67f13;
  wire v3a70c04;
  wire c4699e;
  wire v3777670;
  wire v3a702b0;
  wire v3a58773;
  wire v3a6c39b;
  wire v3749eb2;
  wire v3758e05;
  wire v374a4a0;
  wire v375d22f;
  wire v3a6dae2;
  wire v3777a7e;
  wire v373a188;
  wire v376ddfb;
  wire v375b8b2;
  wire v3a6dc32;
  wire v373421c;
  wire v373f42a;
  wire v3a62037;
  wire v374047a;
  wire v3a70788;
  wire v39ed7e6;
  wire v3731803;
  wire v377f32e;
  wire v37365ce;
  wire v3a70beb;
  wire v3772a9b;
  wire v3a709f3;
  wire v37331a1;
  wire v3726f57;
  wire v373e9a5;
  wire v3a716a3;
  wire v372c713;
  wire v377d714;
  wire v3a62c7d;
  wire v3a6e159;
  wire v373ffa9;
  wire v3755ec0;
  wire v374cb9e;
  wire v375ca93;
  wire v3a6f29a;
  wire v3768622;
  wire v37492bc;
  wire v3777f86;
  wire v3a2978d;
  wire v3a53f2b;
  wire v3a71411;
  wire v377efac;
  wire v376021f;
  wire v3a6ee06;
  wire d35b26;
  wire v37512a0;
  wire v3728f87;
  wire v3a70629;
  wire v3a5f9d2;
  wire v3a5d134;
  wire v3a70f9c;
  wire v3a70101;
  wire v3a6f8fb;
  wire v37558eb;
  wire v374f559;
  wire v3759d3c;
  wire v3a62508;
  wire v374bcb4;
  wire v3a299d7;
  wire v3729127;
  wire v377fb84;
  wire v3758950;
  wire v37721cd;
  wire v37528b9;
  wire v376f911;
  wire v8f30ee;
  wire v3a592f7;
  wire v376f6d1;
  wire b254e2;
  wire v375c541;
  wire v3771bb9;
  wire v3773aa9;
  wire v3a6f5da;
  wire v3a70409;
  wire v3a5b4be;
  wire v3a715b2;
  wire v3a290f9;
  wire v37453dd;
  wire v373cee7;
  wire v3751d30;
  wire v3750df3;
  wire v3740e5a;
  wire afa7f5;
  wire v372eeda;
  wire v373af21;
  wire v3a62fc4;
  wire v37526af;
  wire v3766573;
  wire v3a6eec4;
  wire v372bb72;
  wire v3a70f1d;
  wire v374122a;
  wire v3a60013;
  wire v3a6fbd3;
  wire v375e6a0;
  wire v3746cc1;
  wire v372893a;
  wire v375c4e0;
  wire v3743792;
  wire v375a688;
  wire v3a65b79;
  wire v994115;
  wire v3741d52;
  wire v3741d24;
  wire v376d522;
  wire v37287fb;
  wire v375595c;
  wire v373b610;
  wire v37588a3;
  wire v3a5d4ac;
  wire v3a70540;
  wire v3a70dfc;
  wire v3757044;
  wire v3738a70;
  wire v374ef66;
  wire v360bcf2;
  wire v3a6d156;
  wire v3a6feaa;
  wire v209324e;
  wire v3a6f1ee;
  wire v3723048;
  wire v37785be;
  wire v3a6fe74;
  wire v3758f19;
  wire v376cfc1;
  wire v3a6f0d9;
  wire v3a59c87;
  wire v377c32f;
  wire v3765dda;
  wire v3a7146b;
  wire v3255b23;
  wire v3777bde;
  wire v3a586d0;
  wire v3772c92;
  wire v374cc74;
  wire v3756ec2;
  wire v3a5f5b3;
  wire v374096a;
  wire v374ebc5;
  wire v37681f3;
  wire v374892a;
  wire v3a69123;
  wire v3750e89;
  wire v376c0a0;
  wire d2728f;
  wire v3a57122;
  wire v3a6fcae;
  wire v376acbb;
  wire v3806821;
  wire bb611d;
  wire v373a25b;
  wire v3768726;
  wire v3739c05;
  wire v3a6fc2e;
  wire v3a5a980;
  wire v3a71402;
  wire v374d7ce;
  wire v377add5;
  wire v3a59517;
  wire v376b903;
  wire v372a886;
  wire v3808874;
  wire v1e37442;
  wire v3744a21;
  wire v3746846;
  wire v3a7104d;
  wire v3744dca;
  wire v3377c6a;
  wire v3a6e8d2;
  wire v3a633ac;
  wire v3809eab;
  wire v373e750;
  wire v376c590;
  wire v3258760;
  wire v377583c;
  wire v372b2b4;
  wire v3741714;
  wire v37750e0;
  wire v375cce7;
  wire v3767c3e;
  wire v3a610f7;
  wire v3a65383;
  wire v3a5f4a8;
  wire v374094a;
  wire v376147f;
  wire v3755002;
  wire v3a6fd24;
  wire v374067c;
  wire v3a7152b;
  wire v3a5600a;
  wire v3739934;
  wire v3743327;
  wire v37386f2;
  wire v375eb9c;
  wire v3748ca3;
  wire v375100c;
  wire v3762552;
  wire v3728abd;
  wire c17a4a;
  wire v372794f;
  wire v372791c;
  wire v3761480;
  wire v375444e;
  wire v372f694;
  wire v373b3fb;
  wire v37375ee;
  wire v3a5fdfc;
  wire v3a70116;
  wire v3771fec;
  wire v3739bfa;
  wire v373006f;
  wire v3a709b9;
  wire v377c500;
  wire v374da93;
  wire v3a7070c;
  wire v3a70d30;
  wire v3727dab;
  wire v2acafeb;
  wire v23fd858;
  wire v3a6eb0e;
  wire v3742e40;
  wire v3757ee7;
  wire v3751159;
  wire v3a6a03c;
  wire v3a7101a;
  wire v23fde7f;
  wire v3a6e5f0;
  wire v3a5d494;
  wire v3a6f6a4;
  wire v3a7004f;
  wire v2acaedd;
  wire c41ef0;
  wire v373dceb;
  wire v37757e0;
  wire v375e373;
  wire v3773b23;
  wire v3258d68;
  wire v3766ea9;
  wire v3730cce;
  wire v3a57309;
  wire v37626d5;
  wire v3741aca;
  wire v3a5690e;
  wire v95a0a1;
  wire v37576b1;
  wire v3a656dd;
  wire v377ce1a;
  wire v3767e7e;
  wire v374b025;
  wire v374e92a;
  wire v3a669c6;
  wire v3759586;
  wire v377d04f;
  wire v3a6857b;
  wire v375ecd4;
  wire v3724e14;
  wire v3a6fde6;
  wire v375d388;
  wire v376b856;
  wire v3a70016;
  wire v3734a93;
  wire v325b59d;
  wire v376c25b;
  wire v3747b55;
  wire v376c85c;
  wire v3735e69;
  wire v374ffc1;
  wire v3a5f946;
  wire c5ed52;
  wire v3a6818c;
  wire v373d687;
  wire v375e737;
  wire v3a6dd80;
  wire v3a6f40f;
  wire v3a64ff4;
  wire v3a708d7;
  wire v376ee62;
  wire v37399ef;
  wire v3a549f0;
  wire v376604d;
  wire d70cde;
  wire v3728b1d;
  wire v3a5ed64;
  wire v3759f8b;
  wire v373fa07;
  wire v374ebb0;
  wire v3745b07;
  wire v375b012;
  wire v3770116;
  wire v3a5a03f;
  wire v3a63659;
  wire v374aae0;
  wire v3756e01;
  wire v3744724;
  wire v3a69a04;
  wire v373d136;
  wire v372ef16;
  wire v3757d70;
  wire v373f4ce;
  wire v3a61603;
  wire v376b81b;
  wire v3a6f96f;
  wire v3a658be;
  wire v3a7094d;
  wire v3772ad5;
  wire v3a5ddee;
  wire v3a66750;
  wire v377ccba;
  wire v3727b0e;
  wire v376d07b;
  wire v37437c1;
  wire v377d99d;
  wire v3a71350;
  wire v373ce6d;
  wire v3750078;
  wire v375db7f;
  wire v3a6d1ce;
  wire v375d25d;
  wire v3759daf;
  wire v3a5ef76;
  wire v3a6d3f2;
  wire v374131b;
  wire v3740d32;
  wire v37470c6;
  wire v3a562ea;
  wire v3a620e2;
  wire v376ddc6;
  wire v377ce00;
  wire v375d5f3;
  wire v37685bb;
  wire v3773e5f;
  wire v3739395;
  wire v377d652;
  wire v3a713cc;
  wire v3a71554;
  wire v373f52e;
  wire v376ce4d;
  wire v3a5f0cf;
  wire v3a57f42;
  wire v3a70bf7;
  wire v3a5dd7f;
  wire v3761ed2;
  wire v376f449;
  wire v3771102;
  wire v3774055;
  wire v3a70b97;
  wire v3a70a24;
  wire v373f503;
  wire v3a57506;
  wire v3a58a90;
  wire v3a70d45;
  wire v3a6f837;
  wire v3732c95;
  wire v3a66514;
  wire v37233f1;
  wire v37375e2;
  wire v37440e4;
  wire v374cff2;
  wire v3765f9e;
  wire v37718fb;
  wire v3a709ed;
  wire v3a58967;
  wire v3723c99;
  wire v3779b9c;
  wire v3a70dca;
  wire v373efee;
  wire v3759b20;
  wire v3730568;
  wire v3a5445c;
  wire v372c03b;
  wire v3a5f9d5;
  wire v3a29d87;
  wire v3a6fbac;
  wire v3724ff0;
  wire v3753b1b;
  wire v372b8a0;
  wire v3a5bcfa;
  wire v3766b23;
  wire v3a704ca;
  wire v3761a32;
  wire v3774e8d;
  wire v380777c;
  wire v372de8f;
  wire v375f60e;
  wire v3767ed6;
  wire v2aca770;
  wire v374f78c;
  wire v376a8d5;
  wire v3a69d06;
  wire v3a65f0f;
  wire v3748e81;
  wire v3766025;
  wire v37339c8;
  wire v3752dd0;
  wire v376e431;
  wire v3a7081e;
  wire v3a6146a;
  wire v376dd3d;
  wire v3a5bab6;
  wire v373472c;
  wire v374ec8b;
  wire v37573f4;
  wire v3a66a3b;
  wire v373d262;
  wire v2acb095;
  wire v376223b;
  wire v374f871;
  wire v23fe06e;
  wire v3a6a1b9;
  wire v376ac9b;
  wire v377c57a;
  wire v372ea48;
  wire v3727ee4;
  wire b038e6;
  wire v37341d3;
  wire v377e4b4;
  wire b56d1b;
  wire v3762815;
  wire v37401f0;
  wire v3762414;
  wire v373720a;
  wire v374ea45;
  wire v3728b2f;
  wire v3759c5d;
  wire v3a655c3;
  wire v3737d55;
  wire v3a6fe46;
  wire v3a6ff9f;
  wire v3763056;
  wire v3750a9c;
  wire v3742dac;
  wire v377d2bc;
  wire v3a7037c;
  wire v3746f84;
  wire v3757264;
  wire v3756fba;
  wire v3a5b213;
  wire v3757575;
  wire v3a6b102;
  wire v3a6f5a1;
  wire v3765321;
  wire v3757ffa;
  wire v374dfe1;
  wire v374ae00;
  wire v3770367;
  wire v3729fa4;
  wire v376589f;
  wire v3779477;
  wire v3a65b87;
  wire v372dd98;
  wire v374dfad;
  wire v3746818;
  wire v38072fe;
  wire v376e441;
  wire v3a6895d;
  wire v3779860;
  wire v373cbc2;
  wire v373114f;
  wire v2ff8ce3;
  wire v3a70b35;
  wire v3755d10;
  wire v3a570cd;
  wire v3a70dd9;
  wire v37494ce;
  wire v3a55bd3;
  wire v3745706;
  wire v3a711ab;
  wire v3724df8;
  wire v37448a7;
  wire v376ec0d;
  wire v3768636;
  wire v3773708;
  wire v3a6fa77;
  wire v376cb10;
  wire v3a5dba4;
  wire v374fb30;
  wire v374e800;
  wire v3757ab6;
  wire v372ef36;
  wire v372e885;
  wire v3809561;
  wire v3a707e3;
  wire v3a6ffb2;
  wire v3a5f47b;
  wire v3a70d4e;
  wire v3a5d834;
  wire v9014db;
  wire v376a92f;
  wire v3a5f55e;
  wire v372e02d;
  wire v991591;
  wire v3a5dcd4;
  wire v377af48;
  wire v3a6a635;
  wire v3737edc;
  wire v377bb3a;
  wire v3a6320d;
  wire v372d203;
  wire v3a70222;
  wire v3a6c016;
  wire v3775932;
  wire v2092eac;
  wire v37720e5;
  wire v3a6fac5;
  wire v376de4e;
  wire v374b0c1;
  wire v3a6f314;
  wire v39eb569;
  wire v3742a78;
  wire v3724a4b;
  wire v37545a0;
  wire v374d645;
  wire v3741ac2;
  wire v374c2b4;
  wire v3a6f539;
  wire v3a61f4c;
  wire v374ad7d;
  wire v372c0d6;
  wire v3a6c0ba;
  wire v372b4b4;
  wire v3751925;
  wire v3a6f455;
  wire v3a70135;
  wire v372dc39;
  wire v3730595;
  wire v376ae94;
  wire v375eea5;
  wire v376d19f;
  wire v8ebe6e;
  wire v3a5509a;
  wire v376dad7;
  wire v3a5c7a6;
  wire v944e42;
  wire v374aa46;
  wire v376a2de;
  wire v373a6d9;
  wire v3a7152a;
  wire v3750bc4;
  wire v3736f6d;
  wire v3a5a2e5;
  wire v3a54120;
  wire v373a7b4;
  wire v37430c6;
  wire v3a68276;
  wire v3a68838;
  wire v3751d6f;
  wire v3a63bd4;
  wire v3756546;
  wire v37732a0;
  wire v3a299d4;
  wire v3a2a2ee;
  wire v37c0297;
  wire v3a708d1;
  wire v377de7b;
  wire v3a5ee6b;
  wire v3727540;
  wire v3a66724;
  wire v372af30;
  wire v373b5f5;
  wire v377a121;
  wire v3751004;
  wire v376b67d;
  wire v3743d30;
  wire v3754a54;
  wire v375d8a6;
  wire v3a64082;
  wire v375240c;
  wire v3a64d8f;
  wire v374dc3c;
  wire v373496c;
  wire v3a593cc;
  wire v37787d1;
  wire v3a70c12;
  wire v373e88f;
  wire v374ba88;
  wire v3a6fa5d;
  wire v3255b27;
  wire v3a6fe4d;
  wire v373796a;
  wire v3a7157d;
  wire v375e120;
  wire v3a61519;
  wire v3a6ae12;
  wire v3a6fba2;
  wire v374726f;
  wire v375c2e6;
  wire v3a6f9bf;
  wire v37706e9;
  wire v3766a74;
  wire v3a5a8bf;
  wire v3a70279;
  wire v3a6a910;
  wire v3738855;
  wire v3a6219d;
  wire v372554a;
  wire v3730c69;
  wire v3746caf;
  wire v3776c95;
  wire v372d35f;
  wire v3737c0a;
  wire v377a4f1;
  wire v3759dd9;
  wire v3778fb2;
  wire v377bb86;
  wire v3771e18;
  wire v3a70d05;
  wire v3a5a6f4;
  wire v3a6f0f6;
  wire v8a21c4;
  wire v375153e;
  wire v3a678d2;
  wire v337900b;
  wire v37451ad;
  wire v3a58b1f;
  wire v3a707d1;
  wire v37302ea;
  wire v2925c67;
  wire v23fdbca;
  wire v3745d21;
  wire v374f12d;
  wire v372dbf1;
  wire a11f42;
  wire v376aa6d;
  wire v377b218;
  wire v377c0fe;
  wire v373e49f;
  wire v3737721;
  wire v376b2ab;
  wire v372e250;
  wire v3a7045d;
  wire v372ca24;
  wire v374a277;
  wire v3a6e39a;
  wire v377ad9b;
  wire v375d152;
  wire v374ed5a;
  wire v376ce6f;
  wire v3a6f809;
  wire v373d32e;
  wire v97b684;
  wire v374ae3d;
  wire v375aca9;
  wire v37457b1;
  wire v373a1d7;
  wire v3763a33;
  wire v3a70265;
  wire v3a6fb9e;
  wire v3767690;
  wire v3a6efac;
  wire v37728b1;
  wire v375e1a1;
  wire v3753f62;
  wire v3a64d60;
  wire v375bfd5;
  wire v3752e13;
  wire v373f172;
  wire v3a5bd69;
  wire v376c3fd;
  wire v3777460;
  wire v3a6ec76;
  wire v3a712f2;
  wire v3770c96;
  wire v374e345;
  wire v3760954;
  wire v374e758;
  wire v37237a8;
  wire v3a652b6;
  wire v3a5d45c;
  wire v3a71602;
  wire v3a709b2;
  wire v3731d2d;
  wire v3a6ffd2;
  wire v374aed5;
  wire v375a187;
  wire v374fc17;
  wire v372874e;
  wire v373be73;
  wire v3a5770f;
  wire v3a7158e;
  wire v373852b;
  wire v373eba7;
  wire v3a61280;
  wire v373ba25;
  wire v37477b7;
  wire v376bbc5;
  wire v3a700eb;
  wire v3762e8d;
  wire v3a572ee;
  wire v374a565;
  wire v3765ed6;
  wire v372f96d;
  wire v3a6af4d;
  wire v3a70e71;
  wire v2092f90;
  wire v3a6528b;
  wire v376725a;
  wire v3748645;
  wire v3746feb;
  wire v375070c;
  wire v372d939;
  wire v375a750;
  wire v3a58dc1;
  wire v3a6eae6;
  wire v3a71395;
  wire v3752aa5;
  wire v37270b9;
  wire v3a634fd;
  wire v3737e21;
  wire v3731945;
  wire v373e524;
  wire v3776685;
  wire v3a6f5c8;
  wire v373f8d4;
  wire v3a6df9a;
  wire v380922b;
  wire v3a5b079;
  wire v3377c6c;
  wire v374fef7;
  wire v3a64ca0;
  wire v374b70d;
  wire v3731df6;
  wire v374d173;
  wire v37495f2;
  wire v3a702e5;
  wire v3751cd1;
  wire v379318b;
  wire v3743613;
  wire v3a6a312;
  wire v3a6f86b;
  wire v3751de0;
  wire v3770957;
  wire v37558c7;
  wire v3a5d8b5;
  wire v375456e;
  wire v37538ca;
  wire v377d7a0;
  wire v3a68ee5;
  wire v8a7af6;
  wire v374771c;
  wire v377e586;
  wire v3a6e327;
  wire v3728604;
  wire v3a65c2a;
  wire v35b7b3b;
  wire v3a70e42;
  wire v377281c;
  wire v372a3cb;
  wire v377ea01;
  wire v377c470;
  wire v3744713;
  wire v374f319;
  wire v3769f01;
  wire v3a63bde;
  wire v3760d53;
  wire v3a71046;
  wire v3a6dbaa;
  wire v373f950;
  wire v3747f81;
  wire v1e378ea;
  wire v3a296d8;
  wire v3a705f5;
  wire v3a6fdee;
  wire c4dd17;
  wire v3773089;
  wire v3a6f90e;
  wire v374949f;
  wire v3a70515;
  wire v375c90c;
  wire v375aacf;
  wire v37330ca;
  wire v3a709f1;
  wire v3a6f369;
  wire v377933b;
  wire v374cb62;
  wire v375870e;
  wire v374e82c;
  wire v3723185;
  wire v38087e5;
  wire v37728cd;
  wire v3752d31;
  wire v373d4d1;
  wire v3746cbf;
  wire v3a6f506;
  wire v3a556f8;
  wire v375d661;
  wire v3a60e5d;
  wire v376ed36;
  wire v3752edb;
  wire v3a70ebb;
  wire v372d49e;
  wire v3771dd8;
  wire v3a5c317;
  wire v3a6bbe5;
  wire v3a6f47f;
  wire v376e6e2;
  wire v3a5724f;
  wire v3a6f7a6;
  wire v3a6f710;
  wire v37403fe;
  wire v3a666e8;
  wire v375c505;
  wire v377adf0;
  wire v3747bfe;
  wire v3739c66;
  wire v3733a17;
  wire v3726983;
  wire v3a67a48;
  wire v3a5bd76;
  wire v9a3ffa;
  wire v375eef0;
  wire v372be56;
  wire v3a6eb3e;
  wire v37c0296;
  wire v3770e0e;
  wire v3a6fef5;
  wire v372f99a;
  wire v3738a2b;
  wire v373aa91;
  wire v373c5b5;
  wire v375a6d8;
  wire v3743d03;
  wire v37388d6;
  wire bb49f9;
  wire v372cb2c;
  wire v3744410;
  wire v3750b9b;
  wire v375abf4;
  wire v3a6ff24;
  wire v375921f;
  wire v37419b2;
  wire v374980f;
  wire v373c583;
  wire v372bd5e;
  wire v3776cb6;
  wire v3774e5a;
  wire v3a70bee;
  wire v37671d3;
  wire v3807969;
  wire v3735ad0;
  wire v3a6ddb3;
  wire v377f35c;
  wire v3a6146c;
  wire v3a6f049;
  wire v372706f;
  wire v37649c2;
  wire v375bfa6;
  wire v3a6eb44;
  wire v3756eaf;
  wire v3a7000a;
  wire v1e38283;
  wire v373d0a3;
  wire v3771536;
  wire v3a7084c;
  wire v3763327;
  wire v374e288;
  wire v37597c4;
  wire v3776d6e;
  wire v3725a73;
  wire v3a61462;
  wire v374f0bf;
  wire v377e2b3;
  wire v374c23f;
  wire v374bff0;
  wire v373aee6;
  wire v3749942;
  wire v33789d2;
  wire v3a6376d;
  wire v3a5b4a0;
  wire v35b7070;
  wire cc8eeb;
  wire v376b6fb;
  wire v3763188;
  wire v2acb5c8;
  wire v35b7808;
  wire v376b870;
  wire v3a70d4d;
  wire v376c51e;
  wire v374244e;
  wire v377d7a4;
  wire v3723eef;
  wire v37362ff;
  wire v3a70427;
  wire v377afb7;
  wire v3775476;
  wire v372b3cf;
  wire v3a707c2;
  wire v3a54c2e;
  wire v3a59e1c;
  wire v3a6fc75;
  wire v3a7142a;
  wire v3a7069a;
  wire v3a67983;
  wire v377eb9d;
  wire v3a68834;
  wire v375d4e5;
  wire v377c71d;
  wire v372e031;
  wire v3768828;
  wire v376e2fb;
  wire v3a572bd;
  wire v375da52;
  wire v3778674;
  wire v376f319;
  wire v3a6ba54;
  wire v37351f6;
  wire v3a6a95a;
  wire v3257354;
  wire v3a545c8;
  wire v3a5bc27;
  wire v3a714e0;
  wire v3a5aaf9;
  wire v3a6f810;
  wire v37551b8;
  wire v375b1a0;
  wire v3758435;
  wire v3a6dcbf;
  wire v3a5b9c3;
  wire v3731d66;
  wire v3725e12;
  wire v375515c;
  wire v3771182;
  wire v3751983;
  wire v3a661fe;
  wire aa5556;
  wire v3a713df;
  wire v377a615;
  wire v3772bb3;
  wire v35b70c3;
  wire v3740f7d;
  wire v374535e;
  wire v3a5be93;
  wire v375d832;
  wire v3727c3c;
  wire v3742adb;
  wire v373bcea;
  wire v374d057;
  wire v360d2ce;
  wire v23fd799;
  wire v376486a;
  wire v373c1a2;
  wire v3a6602d;
  wire v3746f58;
  wire v3a700b2;
  wire v3744b55;
  wire v3752115;
  wire v37567f5;
  wire v373013d;
  wire v3a6fcd2;
  wire v3729708;
  wire v3742bc3;
  wire v377eb8b;
  wire v376db27;
  wire v3a56f0b;
  wire v3a61d5b;
  wire v3808d85;
  wire v3a5f0d0;
  wire v3762de5;
  wire v37289bc;
  wire v372b870;
  wire v375f123;
  wire v376297b;
  wire v99b6f5;
  wire v373bbc1;
  wire v377929d;
  wire v3a70aae;
  wire v3774c25;
  wire v3a6177b;
  wire v3a6fd81;
  wire v37425c6;
  wire v3a711db;
  wire v376ac56;
  wire v372e3e7;
  wire v3728343;
  wire v372f520;
  wire v376b504;
  wire v375c99d;
  wire v3740e8d;
  wire v3a65104;
  wire v3a6eae9;
  wire v3a6ffd9;
  wire v38070ea;
  wire v375f742;
  wire v3a68317;
  wire v3776337;
  wire v3724974;
  wire v377acde;
  wire v3a6ef64;
  wire v3a6f816;
  wire v373e6d8;
  wire v3a6c467;
  wire v37581c0;
  wire v3a57836;
  wire v377cb2b;
  wire v37615d8;
  wire v1e382c4;
  wire v373e046;
  wire v3a645d7;
  wire v3768a88;
  wire v3739509;
  wire v3730b23;
  wire v3779d86;
  wire v3a6f4e8;
  wire v37299dd;
  wire c3f48e;
  wire v374e34f;
  wire v3a64e05;
  wire v3754c5e;
  wire v3a6cc9a;
  wire v3a6268c;
  wire v3a70ee5;
  wire v3a6fd7b;
  wire v3727b41;
  wire v3a58134;
  wire v37453f0;
  wire v373594b;
  wire v375bb26;
  wire v3779c38;
  wire v3738f35;
  wire v3a6ff39;
  wire v3a65c2c;
  wire v377086c;
  wire v372c433;
  wire v3a5fb9e;
  wire v372c9eb;
  wire v3a5ae9f;
  wire v3764261;
  wire v3a6a8d2;
  wire v3a70e86;
  wire v376bf69;
  wire v372f391;
  wire v37571a9;
  wire v3748a4f;
  wire v3736739;
  wire v3a63c47;
  wire v37425c0;
  wire v3a5beb6;
  wire v37693af;
  wire v380971a;
  wire v3743cb5;
  wire v3a70065;
  wire v373712d;
  wire v3762d5f;
  wire v375d8ea;
  wire v375b912;
  wire v37319d5;
  wire v374077c;
  wire v3764e58;
  wire v37585a0;
  wire v3a70316;
  wire v3a5bd48;
  wire v3a651b8;
  wire v375ac98;
  wire v3a6bc78;
  wire v373313b;
  wire v373bf45;
  wire v3a63ee6;
  wire v375a16d;
  wire v372ccc4;
  wire v374465a;
  wire v3a7148e;
  wire v374b697;
  wire v375c7d3;
  wire v3a5a258;
  wire v3a65aba;
  wire v376be50;
  wire v3a6f3b9;
  wire v2092a68;
  wire v37507d6;
  wire v373449d;
  wire v3769ad5;
  wire v3776da7;
  wire v3744abe;
  wire v3a57486;
  wire v373d5ac;
  wire v37429c5;
  wire v3a7010a;
  wire v376d0d8;
  wire v3769199;
  wire v3a6f7fa;
  wire v3a6847c;
  wire v3726efb;
  wire v3a5f40e;
  wire v3a6c8c0;
  wire v3761362;
  wire v376a166;
  wire v38074ac;
  wire v3a70574;
  wire v3728a3d;
  wire v3a65afa;
  wire v37627bd;
  wire v376d374;
  wire v3762759;
  wire v3a704d5;
  wire v3a63545;
  wire v3a5f371;
  wire v3762ffa;
  wire v372587b;
  wire v37787ac;
  wire v374424e;
  wire v3a6fbd4;
  wire v3766202;
  wire v3a5e665;
  wire v3a70468;
  wire v376e4a6;
  wire v3a634db;
  wire v3809240;
  wire v3a70f8f;
  wire v375af5d;
  wire v3744a60;
  wire v372ff9e;
  wire v3a57660;
  wire v374061b;
  wire v372912f;
  wire b2ea29;
  wire v3a5a854;
  wire v37564a2;
  wire v377dc65;
  wire v377c79a;
  wire v375cdd7;
  wire b2271d;
  wire v376a6bc;
  wire v373632a;
  wire v3a70348;
  wire v3a6336e;
  wire v372d92b;
  wire v375355c;
  wire v3747d82;
  wire v3a7163c;
  wire v3a59ee0;
  wire v3a621cb;
  wire v3a606b7;
  wire v374af92;
  wire v3a6fa86;
  wire v3741240;
  wire v3764a94;
  wire v3a6fc90;
  wire v373055c;
  wire v3a66822;
  wire v373d4a6;
  wire v3a5d2a6;
  wire v3a6e6a7;
  wire v373a9a9;
  wire v3a703a3;
  wire v3a65388;
  wire v3a6f37d;
  wire v23fdc4f;
  wire v3a6f937;
  wire v3a6eb4b;
  wire v37581f6;
  wire v3740194;
  wire v3a6a6b4;
  wire v374571d;
  wire v3739ec9;
  wire v377d077;
  wire v374a65c;
  wire c6053a;
  wire v3729f64;
  wire v3758924;
  wire v373b95e;
  wire v3a6fdab;
  wire v37756df;
  wire v375b92a;
  wire v3a55f42;
  wire v3a6d625;
  wire v376a8ee;
  wire v3a667a7;
  wire v3a5665e;
  wire v3754727;
  wire v3770c1a;
  wire v3a6512d;
  wire v3747a68;
  wire v3735f51;
  wire v9ecbe0;
  wire v3775931;
  wire v3770a3b;
  wire v3762873;
  wire v37686c2;
  wire v3750625;
  wire v3758636;
  wire v37773a0;
  wire v3a6f379;
  wire v3746061;
  wire v3a568e8;
  wire v3a5923e;
  wire v3a5e541;
  wire v3737421;
  wire v3733e56;
  wire v37738be;
  wire v37650d7;
  wire v375a8d5;
  wire v374dfe3;
  wire v37331e1;
  wire v37716b0;
  wire v3a70b71;
  wire v37410bd;
  wire v3a6cd8b;
  wire v2acae99;
  wire v3a70296;
  wire v374248e;
  wire v375bca7;
  wire v3726e7b;
  wire v376a907;
  wire v3a697d2;
  wire v37451b8;
  wire v376ee43;
  wire ac043d;
  wire v3741e09;
  wire v3742d2a;
  wire v373e2b7;
  wire v3a6ec28;
  wire v373b18b;
  wire v374b549;
  wire v3a6f7d0;
  wire v3a6f2f5;
  wire v3a71506;
  wire v3758f89;
  wire v375ff11;
  wire v3a71285;
  wire v3a5c2d6;
  wire v376746b;
  wire v3740380;
  wire v3a7087f;
  wire v3755d8e;
  wire v374e08e;
  wire v374b5a8;
  wire a26fed;
  wire v374ae7a;
  wire v3a6fa41;
  wire v37384a6;
  wire v375e75d;
  wire v3a63033;
  wire v3768888;
  wire v3746e8b;
  wire v3a6dfa3;
  wire v3a71105;
  wire v375b12b;
  wire v3a70a1f;
  wire v374287d;
  wire v373d68a;
  wire v3a68399;
  wire v1e37bde;
  wire v3766d07;
  wire v3736d58;
  wire v3761b24;
  wire v3a6bce0;
  wire v373d964;
  wire v37327c3;
  wire v376fcd6;
  wire v372981a;
  wire v3a7015b;
  wire v3a6f847;
  wire v37289b0;
  wire v3a6f951;
  wire v37561e0;
  wire v3a715e8;
  wire v3a5842b;
  wire v377b679;
  wire v37626ae;
  wire v3761ac9;
  wire v3763eb0;
  wire v3a5eb0f;
  wire v3737ca0;
  wire v376b5f2;
  wire v375b429;
  wire v2acaef3;
  wire v37624a2;
  wire v37574c0;
  wire v37355c9;
  wire v37592d5;
  wire v3773df0;
  wire v374668d;
  wire v37749f0;
  wire v3730e98;
  wire v3760be5;
  wire v3738ed2;
  wire v3725bb3;
  wire v3741500;
  wire v377e85e;
  wire v372ed51;
  wire v377d142;
  wire v3a71399;
  wire cc2999;
  wire v375ba6d;
  wire v3a62d82;
  wire v374c0a4;
  wire v3770700;
  wire v3739d2a;
  wire v376e8e3;
  wire v3744b11;
  wire v9864ec;
  wire v3a6ff98;
  wire v37340b4;
  wire v3757fa5;
  wire v3a6f888;
  wire v3a6ee50;
  wire v375be57;
  wire v373cc68;
  wire v3741f4b;
  wire v376a40d;
  wire v376265d;
  wire v373fcbf;
  wire v376600a;
  wire v3808f75;
  wire v38067bb;
  wire v2092f1b;
  wire v372ee8a;
  wire v374ea7e;
  wire v374057a;
  wire v3a705f6;
  wire v372feb2;
  wire v375ac20;
  wire v3a5b8b9;
  wire v3746063;
  wire v377f526;
  wire v3776c9c;
  wire v3a70eeb;
  wire v375eeaf;
  wire v3a67d6f;
  wire v374b3bf;
  wire v3a64f7e;
  wire v3a64fb4;
  wire v3778aa0;
  wire v3a7160a;
  wire v3a5d8e8;
  wire v3a6a197;
  wire v3a56e53;
  wire v3a5f51c;
  wire v377918a;
  wire v3775610;
  wire v3a67fe2;
  wire v990999;
  wire v37614fa;
  wire v3a6f818;
  wire v3a701ce;
  wire v3a613f2;
  wire v3a70e3c;
  wire v3a5b6a3;
  wire v39ebad8;
  wire v374717a;
  wire v376b7a8;
  wire v3761825;
  wire v3a6e7e1;
  wire v376b47d;
  wire v3a7153a;
  wire aefb3e;
  wire v3755381;
  wire v3a6de8c;
  wire v377ef4a;
  wire v3a710bd;
  wire v3a70a23;
  wire v3a71019;
  wire v3a55526;
  wire v3a647e2;
  wire v37550d4;
  wire v3a6ebb0;
  wire v3a6f9f6;
  wire v374d04b;
  wire v3729864;
  wire v88d9b8;
  wire v375c48c;
  wire v37765cf;
  wire v39a4f09;
  wire v372ae6a;
  wire v3778572;
  wire v360d048;
  wire v3a61b9c;
  wire v372f6ab;
  wire v3a6d69b;
  wire v3a57d9f;
  wire v37390c9;
  wire v374774a;
  wire v3a540f8;
  wire v3a65911;
  wire v3a707d0;
  wire v3a62481;
  wire v372eb5c;
  wire v3737fca;
  wire v3722fe6;
  wire v3731e50;
  wire v3a712e9;
  wire v38064e3;
  wire v37464f3;
  wire v37673f7;
  wire v3747956;
  wire v3769be7;
  wire v376db9c;
  wire v3a702be;
  wire v3a712bb;
  wire v3a5d20a;
  wire v380701a;
  wire v37617a9;
  wire v373dc73;
  wire v37317f1;
  wire v3806ff6;
  wire v373086c;
  wire v3771ea6;
  wire v3a6211e;
  wire v37313e5;
  wire v374d339;
  wire v373568b;
  wire v372e59e;
  wire v3a59f74;
  wire v3a6a609;
  wire v37682fc;
  wire v376c5b2;
  wire v3a6ffbc;
  wire v375b233;
  wire v377cf7f;
  wire v3754bb1;
  wire v375559b;
  wire v373276f;
  wire v37705c0;
  wire v37591ac;
  wire v376fad7;
  wire v37527dc;
  wire v37694f9;
  wire v37573f5;
  wire v3a61a75;
  wire v3a66161;
  wire v3a59f7d;
  wire v3a6faae;
  wire v3a66170;
  wire v373a9c4;
  wire v3a71249;
  wire v3759b46;
  wire v3a6c15c;
  wire v3757dd4;
  wire v375bdd6;
  wire v372f3b1;
  wire v3a7010d;
  wire v3a5f5db;
  wire v3a7071a;
  wire v3733d60;
  wire v3a7006e;
  wire v3a68789;
  wire v37280b2;
  wire v377d745;
  wire v377cebd;
  wire v3a70a78;
  wire v3a6088f;
  wire v39a53a1;
  wire v375b3b7;
  wire v3a5f5ec;
  wire v3743e3c;
  wire v3a70f80;
  wire v3a6eb83;
  wire v3759f4c;
  wire v372904d;
  wire v3732359;
  wire v377e453;
  wire v3a6ff85;
  wire v3a70d77;
  wire v3a70f78;
  wire v3737280;
  wire v2ff8f8e;
  wire v377a99d;
  wire v3a600b8;
  wire v3a6a0b0;
  wire v377144d;
  wire v3775d59;
  wire v37c02a9;
  wire v3728fda;
  wire v3779ff0;
  wire v377374f;
  wire v376e040;
  wire v3769374;
  wire v3771fb7;
  wire v3a6f347;
  wire v3763f6f;
  wire v3731b02;
  wire v3a70a7d;
  wire v37772d5;
  wire v377422b;
  wire a0cf3e;
  wire v3a7004b;
  wire v376583c;
  wire v37691e6;
  wire v3a6faff;
  wire v3a6bf05;
  wire v375351d;
  wire v3761db0;
  wire v3a6eeb0;
  wire v375cbcb;
  wire v3759aec;
  wire v3751887;
  wire v3a709ae;
  wire v37402ee;
  wire v3763d2c;
  wire v377831d;
  wire v37390ce;
  wire v372adfd;
  wire v3a6793d;
  wire v374a289;
  wire v3a64e18;
  wire v3726e1f;
  wire v375f159;
  wire v372700b;
  wire v373abc5;
  wire v3a70675;
  wire v37532cd;
  wire v3a55c44;
  wire v3a6501d;
  wire v375fb71;
  wire v3378fb8;
  wire v373650c;
  wire v3a5a73d;
  wire v373a331;
  wire v372ab8d;
  wire v3a713c3;
  wire v372bf9f;
  wire v3a59ba9;
  wire v374bbcc;
  wire v3a6ebed;
  wire v3758f58;
  wire v374bfc8;
  wire v375e91f;
  wire v372dd0c;
  wire v377eb45;
  wire v3758c72;
  wire v3a6a693;
  wire v3a5d76d;
  wire v3a5df94;
  wire v3a6051a;
  wire v3a6ef5f;
  wire v3a6f3d5;
  wire v3745f8d;
  wire v3755e97;
  wire v377988b;
  wire v3761d4c;
  wire v37717a4;
  wire v37551ec;
  wire v376c5f3;
  wire v37697ed;
  wire v878208;
  wire v3a6eb7e;
  wire v3738b70;
  wire v3a70ed3;
  wire v377c977;
  wire v3777989;
  wire v374eb9e;
  wire v23fd7e1;
  wire v3749091;
  wire v3a701bf;
  wire v3a5db7d;
  wire v3756526;
  wire v3a6a25c;
  wire v380985a;
  wire v375d85b;
  wire d5c12b;
  wire v3a703a9;
  wire v3a70a7b;
  wire v376b3a9;
  wire v3a712be;
  wire v3a70ce3;
  wire v3751860;
  wire v3a65206;
  wire v3a617fa;
  wire v373ff99;
  wire v376dbdf;
  wire v3a6a2f8;
  wire v375818b;
  wire v3761fd7;
  wire v3a5afd7;
  wire v3777c4e;
  wire v376bcad;
  wire v3a5b585;
  wire v374ee47;
  wire v3a70fa5;
  wire v3a6f71d;
  wire v3a713e1;
  wire v372fc81;
  wire v3731741;
  wire v3a69d8f;
  wire v3766786;
  wire v3a70021;
  wire v3a701d2;
  wire v374b9bb;
  wire v3a58b5a;
  wire v3724270;
  wire v3a6facb;
  wire v377bd63;
  wire d18baa;
  wire v3766d10;
  wire v3a70f5e;
  wire v1e37bb4;
  wire v3a70ff4;
  wire v3a6f670;
  wire v37569b8;
  wire v3a5db7b;
  wire v376f2f8;
  wire v3745ece;
  wire v374ad16;
  wire v37436bc;
  wire v3745b9c;
  wire v3a6feb4;
  wire v374cbc3;
  wire v3a706c2;
  wire v3a696ed;
  wire v3a706dc;
  wire v3a6074d;
  wire b9f474;
  wire v3725230;
  wire v3a6fcab;
  wire v376fd32;
  wire v3727385;
  wire v373e055;
  wire v3a59c73;
  wire v3a6f926;
  wire v3a66d47;
  wire v372feea;
  wire v373fd7b;
  wire v372fdfd;
  wire v373e86e;
  wire v3a5f239;
  wire v3a6d590;
  wire v3765c6d;
  wire v374ab8d;
  wire v3a71066;
  wire v3a667b8;
  wire v3760eb3;
  wire v3740c8e;
  wire v3a5bb6a;
  wire v372a520;
  wire v373823d;
  wire v3725819;
  wire v375f61e;
  wire v3765aee;
  wire v376ac74;
  wire v376d306;
  wire v3741b5e;
  wire v3775533;
  wire v377cc69;
  wire v3752df5;
  wire v37615d0;
  wire v37439ef;
  wire v375db57;
  wire v373e553;
  wire v372d782;
  wire v3758f17;
  wire v3a71650;
  wire v373cc48;
  wire v3a6f7a5;
  wire v374513e;
  wire v376e370;
  wire v3724882;
  wire v376376a;
  wire aadac1;
  wire v37392ad;
  wire v372754b;
  wire v3759144;
  wire v3a6f964;
  wire v3a62f0f;
  wire v35b71ca;
  wire v3752fe6;
  wire v373a8b4;
  wire v39eb4a5;
  wire v3a6fbc4;
  wire v374fbcf;
  wire v37234c3;
  wire v3724e7d;
  wire v375b4cb;
  wire v3a59c72;
  wire v377dbdc;
  wire v3a647c6;
  wire v3806d42;
  wire v377097a;
  wire v376b015;
  wire v3a62184;
  wire v37484e0;
  wire v3a714d5;
  wire v37475d9;
  wire v377fb9d;
  wire v3a5e544;
  wire v3731c7b;
  wire v373133d;
  wire v37549e1;
  wire v375b7bd;
  wire v3a5c3d3;
  wire v374a8bb;
  wire v3764f48;
  wire v37533f6;
  wire v376f051;
  wire v3767fd7;
  wire v375620b;
  wire v3a70b50;
  wire v3a6f66d;
  wire v3725f4a;
  wire v37728a5;
  wire v373d99d;
  wire v3729f14;
  wire v376342f;
  wire v3a6ff32;
  wire v3761c61;
  wire v3a679e2;
  wire v3a70d2c;
  wire v3775537;
  wire v377aefe;
  wire v3a5d9e7;
  wire v3a6f3b1;
  wire v37395e8;
  wire v3a58b9f;
  wire v3725882;
  wire v374190f;
  wire v37315a3;
  wire v37629b0;
  wire v377aecd;
  wire v37797d5;
  wire v3a65b0a;
  wire v37491af;
  wire v3377b02;
  wire v3775a25;
  wire v372b46a;
  wire v3a6f64c;
  wire v3a6842c;
  wire bf6c15;
  wire v3a60f9b;
  wire v37560b0;
  wire v37c025b;
  wire v3a558e5;
  wire v8af425;
  wire v3a6fe7e;
  wire v3a5aef8;
  wire v372ddea;
  wire v376c841;
  wire v37667c6;
  wire v3728419;
  wire v3768fba;
  wire v374948b;
  wire v3a5cb9d;
  wire v373359b;
  wire v3769a00;
  wire v376e7e4;
  wire v3764d40;
  wire v372a1a9;
  wire v3779239;
  wire v3a6f6d5;
  wire v3727d45;
  wire v373540f;
  wire v380952f;
  wire v3730d16;
  wire v373bc8f;
  wire v3742358;
  wire v3753f85;
  wire v376013c;
  wire v372879d;
  wire v375750d;
  wire v1e37b48;
  wire v3a7157f;
  wire v9af5fc;
  wire v3a55c2f;
  wire v3771162;
  wire v372363e;
  wire v3736948;
  wire v3a6ff93;
  wire v3a6fee7;
  wire v3a6ecdf;
  wire v37606b1;
  wire v3a5642f;
  wire v377f46e;
  wire v37512d2;
  wire v39a4d8a;
  wire v3a70154;
  wire v23fe1ca;
  wire v377a7f8;
  wire v3724aa0;
  wire v373d0a2;
  wire v3a7046f;
  wire v3a6f850;
  wire v372a7e7;
  wire v3768b2d;
  wire v3766e3a;
  wire v372f85e;
  wire v372efbe;
  wire v373ac39;
  wire v37639c3;
  wire v37737aa;
  wire v3a6ebc9;
  wire v3a56b92;
  wire v3746a78;
  wire v375863a;
  wire v3a6e438;
  wire v374bf71;
  wire v3a5b7b5;
  wire v37bfc8c;
  wire v9f823e;
  wire v373eff1;
  wire v377f64b;
  wire v39ebacc;
  wire v374776b;
  wire v374e538;
  wire cc70ad;
  wire v3a70d6f;
  wire v373e67e;
  wire v3807107;
  wire v1e3755f;
  wire v3732cb4;
  wire v37770c9;
  wire v373366b;
  wire v3a70d3f;
  wire v3a6396b;
  wire v3756d57;
  wire v375b9b0;
  wire v37294c5;
  wire v377c348;
  wire v3a63383;
  wire v3a59e5e;
  wire v375ee73;
  wire v3a6f781;
  wire v3729186;
  wire v372ab23;
  wire v37646e1;
  wire v373c8c5;
  wire v3a58fa7;
  wire v374a9db;
  wire v372a652;
  wire v3739594;
  wire c0b985;
  wire v3a70147;
  wire v376c854;
  wire v3779491;
  wire v373578d;
  wire v377329f;
  wire v3a70497;
  wire v376b18f;
  wire v373197e;
  wire v3a6f0ee;
  wire v37251cc;
  wire v37705de;
  wire v3a6fd37;
  wire v37314fa;
  wire v37445a8;
  wire v3737223;
  wire v374b0a9;
  wire v375b64b;
  wire v3a6fe96;
  wire v37709d2;
  wire v373b6ca;
  wire v3a6f431;
  wire v3739aa6;
  wire v37627c3;
  wire v3776cbb;
  wire v37752be;
  wire v376a619;
  wire v98bccb;
  wire v377dc15;
  wire v3752ef1;
  wire v377913f;
  wire ccdd71;
  wire v3a57cb4;
  wire v3a6b77d;
  wire v3774b56;
  wire v1e3795b;
  wire v3a5b978;
  wire v3723fec;
  wire v3a6c21d;
  wire v3a62cff;
  wire v375dc01;
  wire v3a6e592;
  wire v3a59b87;
  wire v3a702a5;
  wire v3a6325a;
  wire v3a70a8a;
  wire v3a6e622;
  wire v37489ea;
  wire v375cbe3;
  wire v372c029;
  wire v3744cd7;
  wire v3a6fc04;
  wire v3a5e537;
  wire b9675e;
  wire v3a6fd87;
  wire v380921b;
  wire v376f237;
  wire v373a4ef;
  wire v3735077;
  wire v3732a75;
  wire v23fde6d;
  wire v376fb37;
  wire v376d81a;
  wire v3a71186;
  wire v37784a0;
  wire v3779a06;
  wire v3a71637;
  wire v375993d;
  wire v372642b;
  wire v1e38282;
  wire v375026b;
  wire v37631d9;
  wire v3a700e0;
  wire v3a59158;
  wire v375b82d;
  wire v3765e03;
  wire v3a6f97d;
  wire be9654;
  wire v377a3da;
  wire v374c5c5;
  wire v3a7161a;
  wire v373bf3c;
  wire v374d859;
  wire v3809a6a;
  wire v3745803;
  wire v3a70373;
  wire v3a70850;
  wire v3a6911d;
  wire v3a6cf46;
  wire v3749993;
  wire v3a6fa3a;
  wire v360d0a9;
  wire v3a6c573;
  wire v3737e57;
  wire v3726bdb;
  wire v373b71f;
  wire v3735891;
  wire v3a6f352;
  wire v375ed43;
  wire v3a63f43;
  wire v1e37ae9;
  wire v37444ae;
  wire v3776e23;
  wire v374ed07;
  wire v3a70268;
  wire v375af3c;
  wire v3a711dd;
  wire v377dae3;
  wire v3a71678;
  wire v372a414;
  wire v3a7109d;
  wire v3723f24;
  wire v3a53c9d;
  wire v3a6f801;
  wire v376e717;
  wire v372a92a;
  wire v3767efa;
  wire v3735bef;
  wire v3a6f794;
  wire v3a70c97;
  wire v374253f;
  wire v37c0077;
  wire v3a708f0;
  wire v3750c52;
  wire v37674f6;
  wire v3756aaa;
  wire v3a5a381;
  wire v3748eaa;
  wire v373f057;
  wire v375ca80;
  wire v374bb02;
  wire v3737101;
  wire v3776db6;
  wire v373a972;
  wire v374d4e6;
  wire v372ad1d;
  wire v377340e;
  wire v3a70988;
  wire v37707d5;
  wire v3a70bf4;
  wire v3a707f9;
  wire v373cfd0;
  wire v375b234;
  wire v374fb2f;
  wire v3745451;
  wire v3776c44;
  wire v1e37a04;
  wire v3a6faef;
  wire v3a7142f;
  wire v3a6dded;
  wire v37363da;
  wire v3736c7e;
  wire v37519e2;
  wire v377ce91;
  wire v3a5fd2f;
  wire v3a619a2;
  wire v3776c82;
  wire v3754a41;
  wire v372abb9;
  wire v37695f7;
  wire v377d59e;
  wire v377e630;
  wire v3744142;
  wire v3a70bf5;
  wire v3a59ff7;
  wire v1e3828a;
  wire v3a70303;
  wire v3a655a3;
  wire v3748870;
  wire v37282c1;
  wire v37390f9;
  wire v377b556;
  wire v372fc6c;
  wire v3777870;
  wire v37378ca;
  wire v3744c29;
  wire v3a70e01;
  wire v3776d7d;
  wire v3a70096;
  wire v377bb0e;
  wire v3a6ef98;
  wire v1e37ebb;
  wire v3a55c0c;
  wire c75852;
  wire v374a681;
  wire v3745c8f;
  wire v3a71265;
  wire v377ce7d;
  wire v3772935;
  wire v3a66292;
  wire v375523d;
  wire v377839c;
  wire v1e37579;
  wire v3a5efc4;
  wire v3724987;
  wire v3a70deb;
  wire v3a6f19b;
  wire v3a5b6ac;
  wire v374da8a;
  wire v37252b7;
  wire v3a706c8;
  wire v372a56e;
  wire v3751891;
  wire v3776a59;
  wire v3a6a678;
  wire v3a57e56;
  wire v376a411;
  wire v3a710bf;
  wire v372324a;
  wire v3744c9d;
  wire v3a70074;
  wire v3764703;
  wire v37249cc;
  wire v377d891;
  wire v3a658a9;
  wire v3769c95;
  wire v374f1ae;
  wire v3757e2f;
  wire v3a5c026;
  wire v3a6ffa1;
  wire v3765013;
  wire v375ef1e;
  wire v929796;
  wire v3a6ffd5;
  wire v376f903;
  wire v3a7000f;
  wire v3a7018e;
  wire v3a6f3ee;
  wire v3a539ae;
  wire v3a57378;
  wire v37767d8;
  wire v373c628;
  wire v3a5de35;
  wire v3a5fff6;
  wire v377e0d2;
  wire v3741197;
  wire v3a562a7;
  wire v3735afe;
  wire v3a69ad9;
  wire v3a6e37f;
  wire v372f8af;
  wire v3747b4e;
  wire v375fc83;
  wire v3a70a65;
  wire v375d8af;
  wire v3765d27;
  wire v360c3cc;
  wire v3a6312c;
  wire v3724976;
  wire v375fb86;
  wire v3a62f59;
  wire v3a56e15;
  wire v376610a;
  wire v3a6fdb1;
  wire v376e113;
  wire v376f549;
  wire v37661e4;
  wire v3723686;
  wire v374ce46;
  wire v37738d4;
  wire v1e3787a;
  wire v3a6d9ac;
  wire v373ce4e;
  wire v3769ba0;
  wire v374c9cf;
  wire v3a703c3;
  wire v3a66d14;
  wire v37621d5;
  wire v374d95f;
  wire v373e5f3;
  wire v373083d;
  wire v3a56644;
  wire v3a62a25;
  wire v374bf07;
  wire v3741280;
  wire v3773f88;
  wire v374c870;
  wire v376dce5;
  wire v37695e0;
  wire v3a5a4ce;
  wire v3a55ec0;
  wire v374b21a;
  wire v376ac08;
  wire v373691d;
  wire v3739ddf;
  wire v3a6dafc;
  wire v377d4a6;
  wire v3731bc8;
  wire v3a713a7;
  wire v37784d0;
  wire v3a6fa50;
  wire v37466cb;
  wire v3a6fb6d;
  wire v3752d2c;
  wire v3725947;
  wire v377b94f;
  wire v374c164;
  wire v3778ac2;
  wire v3a59299;
  wire v23fd84e;
  wire v3a6f33e;
  wire v3a655d2;
  wire v3777628;
  wire v3757d76;
  wire v37271ad;
  wire v3728bff;
  wire v374a528;
  wire v23fdbe6;
  wire v3724dfb;
  wire a5679d;
  wire v375e657;
  wire v374834b;
  wire v37296cd;
  wire v374ce04;
  wire v3a6667e;
  wire v3a69591;
  wire v375fcd6;
  wire v377acc6;
  wire v8be8ac;
  wire v3773341;
  wire v37493ce;
  wire v3a6f682;
  wire v373414c;
  wire v37779ea;
  wire v1e37e66;
  wire v37261df;
  wire v3a6f42e;
  wire v3a710f0;
  wire v377b9a2;
  wire v372a1ab;
  wire v375fed2;
  wire v3758615;
  wire v90fd44;
  wire v3a5ae7d;
  wire v3755252;
  wire v3730e43;
  wire v376f321;
  wire v3a5df70;
  wire v3773796;
  wire v37390ca;
  wire v376045b;
  wire v3a62826;
  wire v37598ab;
  wire v3a567b7;
  wire v374a950;
  wire v3a6c97d;
  wire v3758c58;
  wire v3777bfc;
  wire v37693e7;
  wire v375b0d5;
  wire v372d65f;
  wire v3a67403;
  wire v3731bb5;
  wire v37377cf;
  wire v3766e31;
  wire v3a70f10;
  wire v3a6f7ae;
  wire v3a70051;
  wire v3a29a44;
  wire v3767fa4;
  wire v3731e5c;
  wire v372ec1c;
  wire v376ce77;
  wire v372f02f;
  wire v37541ff;
  wire v375cec2;
  wire v377ad57;
  wire a7adce;
  wire v3a63028;
  wire v3738006;
  wire v3a7163a;
  wire v372ca6e;
  wire v372919a;
  wire v373c21c;
  wire v37287f6;
  wire v3731dfd;
  wire v3750088;
  wire v3a636ce;
  wire v3a6eb6a;
  wire v3726379;
  wire v374610d;
  wire v372d732;
  wire v3a7085e;
  wire v3a5fae2;
  wire v3738bdf;
  wire v372bf72;
  wire v372ab45;
  wire v3758a11;
  wire v37348c9;
  wire v3a6f7b7;
  wire v2acaf9d;
  wire v372f649;
  wire v8fa780;
  wire v37234d5;
  wire v374d7fc;
  wire v3a5c1a1;
  wire v3a70766;
  wire v3a7049d;
  wire v3a5da8f;
  wire v3722ebc;
  wire v372c4cd;
  wire v375dc63;
  wire v373a494;
  wire v37730b9;
  wire v37677b4;
  wire v3806ec9;
  wire v376f8ba;
  wire v376e150;
  wire v3378535;
  wire v3767872;
  wire v3761912;
  wire v375745a;
  wire v3a55fc1;
  wire v3770ee9;
  wire v377cf20;
  wire v3742d6c;
  wire v3a62cf3;
  wire v3a70962;
  wire v360d099;
  wire v3735907;
  wire v3a7077a;
  wire v3a6c001;
  wire v3749fd0;
  wire v376046c;
  wire v373e743;
  wire v3a5998b;
  wire v375d455;
  wire v3a6f9f7;
  wire v3761065;
  wire v3a60b37;
  wire v3764983;
  wire v374bf93;
  wire v3a71591;
  wire v3730587;
  wire v3727d77;
  wire v3a6f578;
  wire v3722e49;
  wire v373754d;
  wire v3a660a5;
  wire v377a308;
  wire v38073ff;
  wire v373da6d;
  wire v37313a7;
  wire v375ec1d;
  wire v3806f21;
  wire v3a6f225;
  wire v376d6d9;
  wire v20930fa;
  wire v374f48b;
  wire v3739d69;
  wire v3a70c1b;
  wire v3a62582;
  wire ade0d8;
  wire v3a5a6e6;
  wire v3a61eea;
  wire v3731e3a;
  wire v3a7157e;
  wire v374158d;
  wire v372421d;
  wire v375f77f;
  wire v373fde1;
  wire v3728cb3;
  wire v3763a84;
  wire v376cd14;
  wire v377b2d0;
  wire v3a6f4ba;
  wire v3a6f4f0;
  wire v3761954;
  wire v3a7072d;
  wire v373c56f;
  wire v377da08;
  wire v3a65521;
  wire v3a69409;
  wire v3a7117c;
  wire v3745754;
  wire v3a6f087;
  wire v3750700;
  wire v3776445;
  wire v3a6909f;
  wire v372f2ce;
  wire ae5f9e;
  wire v376f576;
  wire v372e759;
  wire v3a70259;
  wire v3764109;
  wire v37673d6;
  wire v3a56d06;
  wire v3a70e0c;
  wire v3759387;
  wire v377d7a8;
  wire v375e7aa;
  wire v3737193;
  wire v3733734;
  wire v3a59178;
  wire v3a6aa59;
  wire v37c073f;
  wire v372cd3f;
  wire v3a661b5;
  wire v3771913;
  wire v1e37519;
  wire v3a5473a;
  wire v3a6fea9;
  wire v3a6b14a;
  wire v3766c60;
  wire v3a70113;
  wire v3770173;
  wire v377e8ca;
  wire v37796c5;
  wire v3747971;
  wire v3a6b73b;
  wire v3a6f94c;
  wire v3a6f948;
  wire v374d7dc;
  wire v3808c5f;
  wire v37497a5;
  wire v3a60a56;
  wire v377108d;
  wire aa783c;
  wire v3a601cd;
  wire v3a5c65d;
  wire v3738d86;
  wire v3768ec3;
  wire v375a2a7;
  wire v3751c00;
  wire v3763b09;
  wire v3a70b87;
  wire v372b607;
  wire v3736b0e;
  wire v3737ca2;
  wire v8e06bc;
  wire v3753bb4;
  wire v373a4a8;
  wire v37639a1;
  wire v3774a1b;
  wire v3a6dfdb;
  wire v37582a2;
  wire v3a57759;
  wire v37667ed;
  wire v374ab34;
  wire v374e590;
  wire v3a6471e;
  wire v375d0d2;
  wire v3a6256a;
  wire v3776081;
  wire v377df7d;
  wire v372cc69;
  wire v3776f25;
  wire v3a70816;
  wire v37607c6;
  wire v3a70dad;
  wire v2093005;
  wire v3a71476;
  wire v373eedf;
  wire v3a6ebb1;
  wire v375b974;
  wire v3741aa1;
  wire v3735c92;
  wire v3753eb2;
  wire v3a6f5c0;
  wire v3a70cc5;
  wire v3a5eeb4;
  wire v3a6e699;
  wire v3743de1;
  wire v3a65dcf;
  wire v372ba93;
  wire v1e3733c;
  wire v37611df;
  wire v3a70c57;
  wire v3a70607;
  wire v3776fe2;
  wire v377bb62;
  wire v37542af;
  wire v372cc0a;
  wire v373891b;
  wire v380911e;
  wire v373098e;
  wire v3a569dd;
  wire v3a709cb;
  wire v3724a15;
  wire v3726d00;
  wire v373d8e5;
  wire v3750859;
  wire v3729f6a;
  wire v376a715;
  wire v3807604;
  wire v3a712e2;
  wire v376d15d;
  wire v3774e8c;
  wire v377dabc;
  wire v3726d2a;
  wire v3a6fb51;
  wire v37759e3;
  wire v3736026;
  wire v3a6c631;
  wire v3a6eb11;
  wire v373a999;
  wire v3a71380;
  wire v3a703cc;
  wire v3736fdd;
  wire v3a6ef1f;
  wire v373867c;
  wire v3a71454;
  wire v3a626e4;
  wire v9bf1d8;
  wire v3a62092;
  wire v373ee3e;
  wire v3a6f7e1;
  wire v3a6ebea;
  wire v37332ca;
  wire v3732df3;
  wire v3752333;
  wire v37497ce;
  wire v37519cb;
  wire v376a4ba;
  wire v37415c3;
  wire v3773530;
  wire v373efc2;
  wire v376c4fe;
  wire v3a709c4;
  wire v3773a6b;
  wire v3740b8d;
  wire v377b030;
  wire v3a707cf;
  wire v373cc95;
  wire v3745b15;
  wire v3a56318;
  wire v375a9d0;
  wire v3a6f99e;
  wire v37369e4;
  wire v3757e4b;
  wire v375581b;
  wire v3a6c8b4;
  wire v37653d1;
  wire v3a56230;
  wire v3748db2;
  wire v3758d3f;
  wire v373d214;
  wire v3a7059b;
  wire v3a5fdab;
  wire v3731678;
  wire v37256c4;
  wire v3774cd5;
  wire v3a644ab;
  wire v3778d07;
  wire v38076ec;
  wire v3732938;
  wire v3a70f9a;
  wire v3a6f475;
  wire v3a6f235;
  wire v3770eeb;
  wire v374b225;
  wire v37583ea;
  wire v3a57139;
  wire v377c125;
  wire v3a6e790;
  wire v37426bf;
  wire v3a71204;
  wire v372ff37;
  wire v3a5c7be;
  wire v3a67971;
  wire v3a70463;
  wire v3739acd;
  wire v3743f5b;
  wire v373fe39;
  wire v3745236;
  wire v3a70d22;
  wire v3a703f1;
  wire v37276a5;
  wire v376e4bd;
  wire v3740b01;
  wire v374eedb;
  wire v3739d23;
  wire v3726be0;
  wire v3745df8;
  wire v3758f94;
  wire v376575c;
  wire v3a6f99b;
  wire v37605c1;
  wire v3772b2b;
  wire v376132e;
  wire v3753fea;
  wire v871244;
  wire v3737a5a;
  wire v3a6f7bc;
  wire v377050f;
  wire v3a6fcc1;
  wire v372df69;
  wire v3a70a60;
  wire v3773100;
  wire v3806fbf;
  wire v373d139;
  wire v3a70976;
  wire v37315d5;
  wire v3a6c6d6;
  wire v375c1df;
  wire v377e19d;
  wire v3769e49;
  wire v375562a;
  wire v376681a;
  wire v377c6dc;
  wire v37585d8;
  wire v3a62b13;
  wire v3738b0b;
  wire v3a70650;
  wire v37658d9;
  wire v37717ed;
  wire v37503ce;
  wire v372dd77;
  wire v3a53b85;
  wire v3745ced;
  wire v3a71309;
  wire v376ab0f;
  wire v3752cc4;
  wire v3a5d176;
  wire v37351a7;
  wire v3740bba;
  wire v3a708cd;
  wire v377b4fa;
  wire v3769524;
  wire v3a70400;
  wire v374f307;
  wire v375238e;
  wire v373e376;
  wire db20f4;
  wire v376189a;
  wire v3a68f62;
  wire d44200;
  wire v3739f75;
  wire v377521b;
  wire v3760b46;
  wire v374e1f6;
  wire v2092abd;
  wire v3775ca5;
  wire v376beee;
  wire v23fdab8;
  wire v3a7151d;
  wire v376af20;
  wire v3736d0d;
  wire v38088b6;
  wire v3a7051d;
  wire v374f094;
  wire v3759ec7;
  wire v3741069;
  wire v376501e;
  wire v3a7088f;
  wire v3a716a0;
  wire v372dcaa;
  wire v3a6f772;
  wire v3746acf;
  wire v3a6ffc6;
  wire v3a6f081;
  wire v372b3b0;
  wire v3a64eac;
  wire v3a7090b;
  wire v3773f70;
  wire v374fe65;
  wire v3a7156d;
  wire v3777226;
  wire v3a63eaf;
  wire v373ee17;
  wire v2092ec6;
  wire v376c7f9;
  wire v37725d6;
  wire v377b456;
  wire v3723b00;
  wire v3a54b31;
  wire v374b1bc;
  wire v3727eb2;
  wire v376495e;
  wire d26e1e;
  wire v3a67092;
  wire v3807dc9;
  wire v372bd2b;
  wire v373285a;
  wire v3722de8;
  wire v37534c6;
  wire v3a5e2a9;
  wire v3732b15;
  wire v3774058;
  wire v3734c0f;
  wire v3a668a4;
  wire v3a7153c;
  wire v37636e3;
  wire v3768e0c;
  wire v35ba2da;
  wire v3756f06;
  wire v375c671;
  wire b05db7;
  wire v376c2e6;
  wire v3a70bc6;
  wire v3730a3d;
  wire v3a6fa9a;
  wire v372ff70;
  wire v376c1de;
  wire v3a583b0;
  wire v3744d2b;
  wire v3809d49;
  wire v3754dd0;
  wire v3a7167d;
  wire v3a6ca0b;
  wire v373adb9;
  wire v376ef47;
  wire v3758d2a;
  wire v3a564d9;
  wire v373c38b;
  wire v374f749;
  wire v90a475;
  wire v377115c;
  wire v37618e0;
  wire v3807f45;
  wire v3764979;
  wire v3809ebc;
  wire v376eaf1;
  wire v3a60dd5;
  wire v3728373;
  wire v375bd16;
  wire v3727976;
  wire v3a6a536;
  wire v3766803;
  wire v3a6ff04;
  wire v3a621d5;
  wire v374c47e;
  wire v37245f8;
  wire v372e6ee;
  wire v3a6fdd6;
  wire v377609f;
  wire v3a700c6;
  wire v3744cf7;
  wire v3a70319;
  wire v374e28f;
  wire bddd83;
  wire v3723ee4;
  wire v374abb5;
  wire v3a6277d;
  wire v3767e6a;
  wire v3a710b5;
  wire v3a70b17;
  wire v37408e1;
  wire v374d6b2;
  wire v3a6e8d9;
  wire v2093132;
  wire v3762fc3;
  wire v3a5cfac;
  wire v3a70479;
  wire v3a6fafd;
  wire v3760933;
  wire v3a71164;
  wire v375fb03;
  wire v373e0d8;
  wire v3736969;
  wire v373dcdd;
  wire v37229e6;
  wire v3809d8e;
  wire v3725b69;
  wire v37447b9;
  wire v3722968;
  wire v37798bd;
  wire v3750eaa;
  wire v37369b2;
  wire v3a6fafe;
  wire v3764efe;
  wire v2ff9314;
  wire v3a6f1ab;
  wire v3726991;
  wire v3a7046c;
  wire v37598a3;
  wire v3759379;
  wire v3a70c30;
  wire v37423d1;
  wire v3745eab;
  wire v3a6eeef;
  wire v372b7a3;
  wire v3a70252;
  wire v3a6fa22;
  wire v37435fd;
  wire v3738826;
  wire v3a6680b;
  wire v3a57ccf;
  wire v3a6f51e;
  wire v3722d85;
  wire v375043b;
  wire v3a6ff9c;
  wire v3752986;
  wire v3a6f548;
  wire v372b679;
  wire v377f579;
  wire v3a5949f;
  wire v3a64e01;
  wire v372bef4;
  wire v3740614;
  wire v3a566c0;
  wire v375c4ef;
  wire v3a59bf7;
  wire v37273b1;
  wire v3a68b8a;
  wire v375d98c;
  wire v376196f;
  wire v375e06b;
  wire v376d52a;
  wire v375a56b;
  wire v3762c8e;
  wire v3749649;
  wire v3748ff3;
  wire v3771204;
  wire v375a4a0;
  wire v374d1ed;
  wire v3742698;
  wire v3a6f9a1;
  wire v3762cd8;
  wire v3a63fe2;
  wire v372d07b;
  wire v373eea8;
  wire v374b160;
  wire v37797c2;
  wire v3764ef1;
  wire v377a236;
  wire v3a709c3;
  wire v377adbd;
  wire v37664aa;
  wire v3770a1c;
  wire v374ed80;
  wire v376f80c;
  wire v377c71e;
  wire v373f6b1;
  wire v3727e33;
  wire v3a71405;
  wire v3743dc4;
  wire v3739731;
  wire v3745186;
  wire v373bd3d;
  wire v3728876;
  wire v37512b3;
  wire v3767ef0;
  wire v3731780;
  wire v37738e9;
  wire v377a916;
  wire v3a61410;
  wire v376832f;
  wire v3751210;
  wire v372baa1;
  wire v3a6a478;
  wire v3740328;
  wire v3a711f8;
  wire v377094d;
  wire v3a70f8b;
  wire v377f829;
  wire v375f15c;
  wire v3a6f556;
  wire v3735cb2;
  wire v3735ee1;
  wire v3754956;
  wire v37602b1;
  wire v3754740;
  wire v3a70d97;
  wire v3a6c793;
  wire v373483e;
  wire v376f9ac;
  wire v3a67af1;
  wire v3a6eb45;
  wire v3a6eb81;
  wire v3a70e52;
  wire v23fd7d9;
  wire v374ad1e;
  wire v3773d82;
  wire v3723ace;
  wire v374314f;
  wire v375e177;
  wire v37763bd;
  wire v3740c92;
  wire v3a7130b;
  wire v3730d64;
  wire v3a6cae3;
  wire v375780e;
  wire v3774e48;
  wire v3a5f281;
  wire v3734502;
  wire v3754d47;
  wire v3746069;
  wire v3735fb3;
  wire v3749165;
  wire v3a714c9;
  wire v3743e56;
  wire v37677ee;
  wire b6390c;
  wire v3722e7a;
  wire v3a700e2;
  wire v375b828;
  wire v375ea85;
  wire v377edd6;
  wire v377abe1;
  wire v3a7143d;
  wire v374c34d;
  wire v3a6f40d;
  wire v37476b8;
  wire v2e5fb38;
  wire v3724696;
  wire v373f687;
  wire v374a058;
  wire v373c263;
  wire v377c4d7;
  wire v3777239;
  wire v3753f77;
  wire v3a65df3;
  wire c0d797;
  wire v3a6f5e9;
  wire v3731f6b;
  wire b736f4;
  wire v375be11;
  wire v3a605d3;
  wire v373ea00;
  wire ae60a0;
  wire v37326be;
  wire v3734aae;
  wire v3772d6e;
  wire v8cb684;
  wire v3748f09;
  wire v37469c4;
  wire v373ff5c;
  wire v3752183;
  wire v377a9b8;
  wire v3765b9b;
  wire v3a577de;
  wire v375e9c8;
  wire v373c239;
  wire v38098b0;
  wire v374999b;
  wire v1e3771d;
  wire v3a6556a;
  wire v3a7154f;
  wire adf1da;
  wire v2ff8c74;
  wire v3a708c8;
  wire v375460c;
  wire v3a7149d;
  wire v3a681e8;
  wire v3772f0f;
  wire v37767fa;
  wire d2afa4;
  wire v374bcb5;
  wire v3a70e99;
  wire v3737b19;
  wire v3a666a9;
  wire v37723c6;
  wire v3739e21;
  wire v372c17e;
  wire v3741dee;
  wire dc5fea;
  wire v373e8df;
  wire v372dcc0;
  wire v3740af7;
  wire v3a6856a;
  wire v3771160;
  wire v374b7e8;
  wire v3a5a219;
  wire v37736b3;
  wire v373c76c;
  wire v374170e;
  wire v373ba84;
  wire v373046c;
  wire v3a63f57;
  wire v3724e60;
  wire v3a66f83;
  wire v3a6f425;
  wire v3770f3a;
  wire v3a6ff3f;
  wire v3a6fe3e;
  wire v3752862;
  wire v3758133;
  wire v3768421;
  wire v373f392;
  wire v374dd24;
  wire v373a0bf;
  wire v374e35e;
  wire v374eb6a;
  wire v3a60576;
  wire v374ab1e;
  wire v3a6f0e7;
  wire v372936a;
  wire v3a5727d;
  wire v3773048;
  wire v3a6cf5d;
  wire v3761b3d;
  wire v3a6f4d0;
  wire v3773bb0;
  wire v3756c5d;
  wire v376db34;
  wire v3a70a37;
  wire v3a712c6;
  wire v377bac2;
  wire v3a6eb63;
  wire v373d4e8;
  wire v373a2fc;
  wire v3730f98;
  wire v3750037;
  wire v3a5e81d;
  wire v3723493;
  wire v374616d;
  wire b66167;
  wire v375be63;
  wire v3739fff;
  wire v373ef69;
  wire v376d509;
  wire v3a6de03;
  wire v37747c0;
  wire v3a7008b;
  wire v3a61b63;
  wire v3a713d8;
  wire v37798c3;
  wire v3729ae4;
  wire v3a67904;
  wire v3751215;
  wire v3723e64;
  wire v376f9d9;
  wire v376102a;
  wire v3765cfd;
  wire v377ae9c;
  wire v375c4a1;
  wire v3a703ad;
  wire v3a7008c;
  wire v3736a23;
  wire v3a6995c;
  wire v3746e85;
  wire v375c76b;
  wire v3a5a81d;
  wire v3a6f4c9;
  wire v3769d79;
  wire v374069b;
  wire v3806c04;
  wire v3a67dab;
  wire v3a5637b;
  wire v377beba;
  wire v377a1ef;
  wire v37360df;
  wire v37644b7;
  wire v3a6f28b;
  wire v3779069;
  wire v3a63556;
  wire v3736260;
  wire v375058a;
  wire v37411ca;
  wire v377e852;
  wire v3774d9c;
  wire v3a5902f;
  wire v3a673d3;
  wire v3a6c68c;
  wire v376b4e5;
  wire v374838d;
  wire v3a6fa44;
  wire v3a540a1;
  wire v3a712a2;
  wire v37474d6;
  wire v3a70217;
  wire v3734ab5;
  wire v374f543;
  wire v375d4d4;
  wire v3775e81;
  wire v377d7bd;
  wire v3a5d40d;
  wire v3a5b903;
  wire v372be16;
  wire v9773b9;
  wire v372ad4e;
  wire v3a706a4;
  wire v37445ff;
  wire v375777d;
  wire v377c700;
  wire v3a577fe;
  wire v37769cc;
  wire v3a6f833;
  wire v3a6b41e;
  wire v3a7149e;
  wire v89a0d1;
  wire v3a62415;
  wire v374c840;
  wire v374953c;
  wire v377d06b;
  wire v376a0f6;
  wire v3742efa;
  wire v23fd817;
  wire v37645eb;
  wire v3770aa1;
  wire v377055c;
  wire v377584f;
  wire v3749106;
  wire v37419ca;
  wire v377f113;
  wire v3a5a637;
  wire v3a6b31c;
  wire v3725dd5;
  wire v3a713bf;
  wire v3773f26;
  wire v37588cf;
  wire v372a738;
  wire v3738f37;
  wire v375e510;
  wire v3756da3;
  wire v3809dcb;
  wire v3757dad;
  wire v37647e7;
  wire v375082a;
  wire v3a6f9f8;
  wire v373568c;
  wire v3a5ff5a;
  wire v3a5c80e;
  wire v3779183;
  wire v3a6f736;
  wire v3a70501;
  wire v374801f;
  wire v3809e72;
  wire v3a5db94;
  wire v3a59f8c;
  wire v376a5c1;
  wire v37520b7;
  wire v3a70159;
  wire v37617d4;
  wire v3741e80;
  wire v372a831;
  wire v377497c;
  wire v37740fd;
  wire d1e3dd;
  wire v3a6802f;
  wire v372c221;
  wire v3a7098f;
  wire v3a573af;
  wire v3a60358;
  wire v3a6f6c7;
  wire v373e34e;
  wire v3747514;
  wire v373419f;
  wire v374d643;
  wire v376a58a;
  wire v3765a4a;
  wire v3a7083e;
  wire v376b0d6;
  wire v37313b6;
  wire v3741dab;
  wire v3746ffa;
  wire v375f2ba;
  wire v377dbd7;
  wire v375705a;
  wire v3728bc3;
  wire v374e3ab;
  wire v3a6f901;
  wire v3a6aea3;
  wire beb41d;
  wire v374de3d;
  wire v3a70a2d;
  wire v3a6f703;
  wire v39a4e7e;
  wire v3a66c22;
  wire v3729844;
  wire v372be4a;
  wire v3a710e1;
  wire v374c671;
  wire v3a56bd5;
  wire v3a62a53;
  wire v375ba37;
  wire v37640e9;
  wire v374c5c6;
  wire v3743018;
  wire v373052f;
  wire v3985142;
  wire v3a6fec8;
  wire v37477d3;
  wire v3755423;
  wire v3a7157c;
  wire v3764caf;
  wire v3a65ca8;
  wire v373c983;
  wire v3a64225;
  wire v3a61535;
  wire v375f94a;
  wire v3a6e52e;
  wire v3a70853;
  wire v3808899;
  wire v377e156;
  wire v373d55f;
  wire v37582e1;
  wire v3759ce2;
  wire v377db66;
  wire v3741fe8;
  wire v3a6a73d;
  wire v3734d58;
  wire v3747b78;
  wire v37658af;
  wire v3a7010f;
  wire v3a6fc54;
  wire v3727486;
  wire v3747d68;
  wire v3a6f495;
  wire v377ea64;
  wire v3a71057;
  wire v3a58b04;
  wire v3761178;
  wire v376b40c;
  wire v3807729;
  wire v374e8a2;
  wire v3a553bc;
  wire v3a59cce;
  wire v3a6bba5;
  wire v3738b0f;
  wire v3a66998;
  wire v3806624;
  wire v3a69892;
  wire v37524b2;
  wire v3731eb8;
  wire v3738510;
  wire v3a6fb95;
  wire v8bc0e2;
  wire v3a603b6;
  wire v376cbbe;
  wire v372f441;
  wire v3760c32;
  wire ca32a1;
  wire be145a;
  wire v3a6f39b;
  wire v3a61e59;
  wire v372f475;
  wire v3a705fb;
  wire v372f236;
  wire v3a627a4;
  wire v373744b;
  wire v3a6ff59;
  wire v3722bcf;
  wire v3a6ef86;
  wire v3766ddb;
  wire v373015f;
  wire v374549a;
  wire v3a64ebb;
  wire v37729ac;
  wire v37596c8;
  wire v3739311;
  wire v374b429;
  wire v3a6fedc;
  wire v3a711f9;
  wire v3a6605d;
  wire v375aafe;
  wire v377498e;
  wire v3a6439a;
  wire v375e6b2;
  wire v377b461;
  wire v37482c8;
  wire v3729d1b;
  wire v376a898;
  wire v3a6f547;
  wire v372d8c9;
  wire cb89d9;
  wire v373ca0e;
  wire v2ff8be4;
  wire v372d3e5;
  wire v37331c0;
  wire v3a701a5;
  wire v3a6f054;
  wire v3764d26;
  wire v374640f;
  wire v3a6dcf5;
  wire v375b8cf;
  wire v374e968;
  wire v3a70a3e;
  wire v3769b7e;
  wire v3a6b90e;
  wire v3a70a2c;
  wire v37776eb;
  wire v377ed25;
  wire v3a64b87;
  wire v3a6cf44;
  wire v3a7018d;
  wire v372b0b0;
  wire v3766c86;
  wire v3742afe;
  wire v372d59d;
  wire v3a71030;
  wire v373f5b1;
  wire v376801c;
  wire v3753bfb;
  wire v3a63d7a;
  wire v373ea71;
  wire v3766da7;
  wire v3a6f462;
  wire v3a5d3fc;
  wire v3a71388;
  wire v37291f4;
  wire v3a706f4;
  wire v377e319;
  wire v376e093;
  wire v375ea72;
  wire v3a70cd9;
  wire v377021d;
  wire v3744df8;
  wire v374b35e;
  wire v3a70937;
  wire beb1cf;
  wire v377cdee;
  wire v374d183;
  wire v37643af;
  wire v3a71250;
  wire v372c14d;
  wire v375d078;
  wire v3a6fa15;
  wire v3a70a55;
  wire v3764af3;
  wire v37246a5;
  wire v3767848;
  wire v3a6e846;
  wire v37629cf;
  wire v374409a;
  wire v39a5420;
  wire v3a706a6;
  wire v3a59d5f;
  wire v377de0d;
  wire v376071e;
  wire v3a5b774;
  wire v3754b83;
  wire v3a6f764;
  wire v3742dc6;
  wire v372d434;
  wire v3755305;
  wire v3a702b6;
  wire v3768fe7;
  wire v37766fb;
  wire v373ec34;
  wire v3733c53;
  wire v377c0bd;
  wire v37745eb;
  wire v3a6effc;
  wire v375e486;
  wire v3a60e4c;
  wire ab4f60;
  wire bdc0a1;
  wire v3735486;
  wire v37524cf;
  wire v3779852;
  wire v39a5359;
  wire v3a606b9;
  wire v3a53d98;
  wire v3766307;
  wire v3a70db1;
  wire v376eef5;
  wire v3a62cda;
  wire v3807d51;
  wire v374a795;
  wire v3731edf;
  wire v3738cd4;
  wire v3a67c41;
  wire v3a6c022;
  wire v3a68e0d;
  wire v3a70fde;
  wire v3756d56;
  wire v37645f6;
  wire v3a5b3dc;
  wire v3a7001c;
  wire v374b867;
  wire v3752b6d;
  wire v374fdc8;
  wire v377a0e7;
  wire v377c77a;
  wire v3775dbc;
  wire a75a41;
  wire v374eab4;
  wire v37301d8;
  wire v3a5b1ca;
  wire v3a5bc5d;
  wire v3a6d2ae;
  wire v3777790;
  wire v3742f52;
  wire v3774391;
  wire v3a70a97;
  wire v377a883;
  wire v3a61123;
  wire v3729a7a;
  wire v376d66b;
  wire v375f2f3;
  wire v3a58c15;
  wire v3747c23;
  wire v3a5c576;
  wire v35b77ab;
  wire v3723f33;
  wire v3a5664b;
  wire v3747367;
  wire v376a015;
  wire v376b4ad;
  wire v3a6c6ad;
  wire v3729801;
  wire v39eb590;
  wire v3729793;
  wire v377e4d8;
  wire v372b59d;
  wire v3a71016;
  wire v3a6df14;
  wire v377ec28;
  wire v3728c23;
  wire v3771a11;
  wire v3a6c98c;
  wire v3724e30;
  wire v3758ff0;
  wire v3a70105;
  wire v3a6ff61;
  wire v3749628;
  wire v3734d9a;
  wire v3809380;
  wire v37377df;
  wire v3766d4b;
  wire v39a4ca6;
  wire v37652ae;
  wire v3765324;
  wire v3a701f0;
  wire v374ee76;
  wire v3751a0b;
  wire v3a6ffb6;
  wire v37724ca;
  wire v372c3d4;
  wire v3a661f1;
  wire v3770a8c;
  wire v3a696ee;
  wire v377a275;
  wire v3a5ef5c;
  wire v3749ec1;
  wire v3a5a806;
  wire v37628f6;
  wire v374431a;
  wire v377dc0c;
  wire v3a682b1;
  wire v37782c9;
  wire v3a705ad;
  wire v375c675;
  wire v37396f7;
  wire v3753cf6;
  wire v374ef62;
  wire v37450cb;
  wire v3a64349;
  wire v3a71645;
  wire v372b551;
  wire v376d88f;
  wire v3766a7d;
  wire v3733392;
  wire db0673;
  wire v9ed516;
  wire v3730e2a;
  wire v3a639a2;
  wire c51aa0;
  wire v3a70bd6;
  wire v374677a;
  wire v373732f;
  wire v3735417;
  wire v3753189;
  wire v3752a0d;
  wire v3a6af83;
  wire v3744efc;
  wire v3a6ac17;
  wire v3a55d64;
  wire v375918d;
  wire v3763c0d;
  wire v377cc52;
  wire v3776864;
  wire v3a70fcd;
  wire v37370a1;
  wire v375d288;
  wire v3a645ca;
  wire v374693f;
  wire v37705f3;
  wire v37660dd;
  wire v3a65e3c;
  wire v373f8f8;
  wire v3743de6;
  wire v372f1d4;
  wire v3744280;
  wire v377a42f;
  wire v3a63a7a;
  wire dc47a7;
  wire v37416c6;
  wire v3a6f55b;
  wire v376df4c;
  wire v3a5e2c8;
  wire v3a5ae76;
  wire v3a6a199;
  wire v376abdf;
  wire v373bfd3;
  wire v374b03c;
  wire v3a5762d;
  wire v3807bfa;
  wire v3726efd;
  wire v3768ac9;
  wire v372de49;
  wire v3729440;
  wire v37751ae;
  wire v372bccc;
  wire v3a6f7d4;
  wire v23fdbc1;
  wire v373f3dd;
  wire v375f5c1;
  wire v3777631;
  wire v3a29835;
  wire v3a6f0ca;
  wire v373501a;
  wire v3a69d78;
  wire v3a6efb7;
  wire v372953c;
  wire v3a5bd12;
  wire v3a6f827;
  wire v3775cc9;
  wire v374f16d;
  wire v373a6ba;
  wire v3762a26;
  wire v3a578ef;
  wire v3a6fe3f;
  wire v376fd85;
  wire v37378d4;
  wire v3a65af6;
  wire v3a6eaf6;
  wire v37247cf;
  wire v3a67bce;
  wire v3a5f714;
  wire v375e346;
  wire v3775dfb;
  wire v3749ed5;
  wire v374888e;
  wire v377abbe;
  wire v3749762;
  wire v3a67f5c;
  wire v3766658;
  wire v3778eed;
  wire v3a70107;
  wire v3737711;
  wire v3a7165a;
  wire v3758b45;
  wire v3a556df;
  wire v3a56827;
  wire v3a62fc9;
  wire v376e9ed;
  wire v3a6f226;
  wire v3a6f4f7;
  wire v3a71664;
  wire v3a702f9;
  wire v374182b;
  wire v3a70bbd;
  wire v3a6367f;
  wire v3a5fa09;
  wire v37318cb;
  wire v3a585d3;
  wire v372f2ae;
  wire v373ec38;
  wire v3734331;
  wire v374d490;
  wire v376e31a;
  wire v3763cef;
  wire v28896cd;
  wire v3769323;
  wire v375d6b4;
  wire v940c77;
  wire v377aa5d;
  wire aa8b86;
  wire v3a5c73c;
  wire v37403ef;
  wire v3742623;
  wire v3a6f3f2;
  wire v372351f;
  wire v3a70e68;
  wire v3a6257d;
  wire v373d40c;
  wire v3732f4d;
  wire v377e568;
  wire v377673f;
  wire v3779d6b;
  wire v375aea8;
  wire v372f765;
  wire v372c921;
  wire v3a6ffc5;
  wire v3738a45;
  wire v37418ab;
  wire v375a513;
  wire v3761d84;
  wire v375e439;
  wire v3768727;
  wire v3a6f7e2;
  wire v37624e5;
  wire v376dffd;
  wire v3779195;
  wire v374bd7d;
  wire v3a71610;
  wire v86d727;
  wire v3a710d3;
  wire v3752b90;
  wire v3a6ff0b;
  wire v3806f68;
  wire v373b209;
  wire v37518fb;
  wire v3a70504;
  wire v3a62070;
  wire v3a6f7dd;
  wire v3757735;
  wire v37754f6;
  wire v3a70f3b;
  wire v3a6fda8;
  wire v3a6f957;
  wire v3a58dfc;
  wire v3806579;
  wire v375269c;
  wire v3735f0b;
  wire v3a70cb6;
  wire v375a312;
  wire v3a568e4;
  wire v3a70fe8;
  wire v3769d48;
  wire v3746200;
  wire v3a5c6d0;
  wire v3773f2b;
  wire v37524b4;
  wire v377c065;
  wire v3a6c4a4;
  wire v37654e0;
  wire v3a6274c;
  wire v376a556;
  wire v3725a6e;
  wire v374a262;
  wire v376ce90;
  wire v3762333;
  wire v374bdfe;
  wire v373d735;
  wire v375e721;
  wire v3769424;
  wire v38073b5;
  wire v375783b;
  wire v3a71101;
  wire v3a70941;
  wire v374b2f5;
  wire v3a6fc70;
  wire v3727ee9;
  wire v3806542;
  wire v3764f6a;
  wire v3807414;
  wire v373d142;
  wire v37419da;
  wire v9864a7;
  wire v3733886;
  wire v3750a45;
  wire v3a6fed7;
  wire v37585bd;
  wire v37472ea;
  wire v37446b1;
  wire v3a6af23;
  wire v3a6eef5;
  wire v3732c0a;
  wire v3a555d7;
  wire v37334a3;
  wire v377c58e;
  wire v3a64f63;
  wire v37276d6;
  wire v377a477;
  wire v3a706c1;
  wire v373a26b;
  wire v3808d74;
  wire v373a4f7;
  wire v3774add;
  wire b7df2b;
  wire v374e1c3;
  wire v3a70124;
  wire v9cbad6;
  wire v3a6f1f2;
  wire ce4c9b;
  wire v3762cca;
  wire v377402f;
  wire v37678eb;
  wire v374bcfb;
  wire v3a66c2f;
  wire v3733726;
  wire v376e35e;
  wire v3760452;
  wire v377445c;
  wire v374195f;
  wire v37706fd;
  wire v3771fd8;
  wire v3a6fcad;
  wire v37439c2;
  wire v3759d52;
  wire v3a63f06;
  wire v3a701d9;
  wire v3a70ec9;
  wire v374db32;
  wire v376cbb7;
  wire v3a70cfc;
  wire v373058e;
  wire v3a6fd12;
  wire v3a63ae9;
  wire v3724060;
  wire v3749242;
  wire v3a680e1;
  wire v3746008;
  wire v372ee5a;
  wire v376ce59;
  wire v3a555e5;
  wire v360c5d9;
  wire v3748e5a;
  wire v3808cbf;
  wire v3a6fb8a;
  wire v3758559;
  wire v37408e4;
  wire v375a500;
  wire v3a702c5;
  wire v377312b;
  wire v3744e62;
  wire v374c05b;
  wire v3722e52;
  wire v376a0d2;
  wire v376bded;
  wire v2ff8ee1;
  wire v3a5ace8;
  wire v377c8fd;
  wire v37621c1;
  wire v377ba78;
  wire v3a683d9;
  wire v376bd96;
  wire v3767640;
  wire v3757888;
  wire v375bc70;
  wire v3a6fc07;
  wire v3a70994;
  wire v375f2b3;
  wire v372fef2;
  wire v37291c7;
  wire v3a65760;
  wire v37355d6;
  wire v377007d;
  wire v374731f;
  wire v3a701c6;
  wire v3a639e7;
  wire v37678f8;
  wire v380958f;
  wire v373a756;
  wire v375f8f2;
  wire v3758526;
  wire v37447df;
  wire v3775942;
  wire v3771252;
  wire v3a6eb37;
  wire v3a628ef;
  wire v3a629a9;
  wire v3a59c0b;
  wire v374b07b;
  wire v374fc6c;
  wire v3a6f6de;
  wire v373ccb9;
  wire v374d2dd;
  wire v377702c;
  wire v3755928;
  wire v3a7002c;
  wire v3a65934;
  wire v376ed91;
  wire v373bff4;
  wire v374e9ac;
  wire v3735ea8;
  wire v376158d;
  wire v377a8ea;
  wire v2acafb4;
  wire v3746b22;
  wire v377a0cb;
  wire v3736613;
  wire v3a6d930;
  wire v3a70b90;
  wire c80162;
  wire v37663a2;
  wire v373c428;
  wire d39337;
  wire v377c546;
  wire v375602e;
  wire v3a701ab;
  wire v377ed24;
  wire v375d263;
  wire v376eb68;
  wire v3a703f2;
  wire v3760765;
  wire v37485cb;
  wire bb4062;
  wire v3767f9a;
  wire v3a70d26;
  wire v3753e23;
  wire v3728a6d;
  wire v375ab92;
  wire v372e02c;
  wire v374fd0b;
  wire v37441b5;
  wire v372e27f;
  wire v3736f3b;
  wire v3a702e1;
  wire v3764dc0;
  wire v37587fa;
  wire v375c60f;
  wire v375e9ef;
  wire v372a965;
  wire v37775d9;
  wire v374dfea;
  wire v3770f6e;
  wire v3a70088;
  wire v3a7005f;
  wire v3a60b88;
  wire v3a701e0;
  wire v3a57de9;
  wire v3744aa9;
  wire v375ed37;
  wire v373ce36;
  wire v375e6fc;
  wire v37476d9;
  wire v377bc9f;
  wire v3759aea;
  wire v3a6900c;
  wire v3a6fcaa;
  wire v37531ff;
  wire v374037a;
  wire v3a70b08;
  wire v3a5a1ff;
  wire v3735bdc;
  wire ad3125;
  wire v373350e;
  wire v3743ff2;
  wire v3a6f008;
  wire v376d33b;
  wire v3a7079d;
  wire v377a855;
  wire v375f84b;
  wire v3736f36;
  wire v3a70656;
  wire v3a6eb9e;
  wire v93144b;
  wire v372edf8;
  wire v3745db5;
  wire v3a7028a;
  wire v3774492;
  wire v3a71002;
  wire v3767a21;
  wire v373d8c3;
  wire v3753900;
  wire v376bc9b;
  wire v373db25;
  wire v3a57ef6;
  wire v3767c44;
  wire v373b17c;
  wire v3745484;
  wire v3a5f315;
  wire v3772513;
  wire v374eaeb;
  wire v3a5c562;
  wire v374e019;
  wire v374546c;
  wire v3772612;
  wire v3a711c8;
  wire v3a66e30;
  wire v3a6f79f;
  wire v3764dda;
  wire v3779958;
  wire v3769980;
  wire v373fe8f;
  wire v3a6f95b;
  wire v3a616aa;
  wire v374cb86;
  wire v3a551bd;
  wire v3773950;
  wire v3a6fa62;
  wire v375984e;
  wire v3760f87;
  wire v377b07a;
  wire v3a6f829;
  wire v3a61f83;
  wire v374254d;
  wire v376b012;
  wire v373f27d;
  wire b58331;
  wire v3a70c36;
  wire v37741bc;
  wire v375d4fa;
  wire v3764a1c;
  wire d3c22f;
  wire v3731d89;
  wire v372a1d6;
  wire v3756a6f;
  wire v3743ea8;
  wire v209323b;
  wire v3741d99;
  wire v374874a;
  wire v3a6becb;
  wire v3a6f4c3;
  wire v3a70e21;
  wire v37291d1;
  wire v375964f;
  wire v3a60130;
  wire v373cf60;
  wire v3747787;
  wire v373af66;
  wire v37557a0;
  wire v37770f5;
  wire v3a68004;
  wire v3a708f2;
  wire v37250fa;
  wire v3a6fc7a;
  wire v377f548;
  wire v3778f83;
  wire v3a5a80c;
  wire v3777ca9;
  wire v3a70a1a;
  wire v376c13c;
  wire v372d86a;
  wire v3772af6;
  wire v3808553;
  wire v373c668;
  wire v374e3c2;
  wire v377e9aa;
  wire v3a7035a;
  wire v374572e;
  wire v373893a;
  wire v374e0a9;
  wire v3751d41;
  wire v37438fc;
  wire v3a7156e;
  wire v3754fcc;
  wire v376e7cf;
  wire v8e42b4;
  wire v3a62812;
  wire v3a6a413;
  wire v3a70e6a;
  wire v3740bb7;
  wire v374ac57;
  wire v3a6cfa1;
  wire v373a832;
  wire v39ebb20;
  wire v37463de;
  wire v3770d93;
  wire v3756aea;
  wire v3738d51;
  wire v373d4c6;
  wire v3a6fde9;
  wire v3a705a5;
  wire v37397f0;
  wire v375ea89;
  wire v377d69c;
  wire v3746a7e;
  wire v372c676;
  wire v3a6f7f9;
  wire v376c1cc;
  wire v373c387;
  wire v3257329;
  wire v37297e4;
  wire v375bf93;
  wire v3756ef4;
  wire v3746bce;
  wire v3a70ea5;
  wire v3a7062f;
  wire v3a29810;
  wire v3a70c1f;
  wire a26159;
  wire v3745dac;
  wire v3a5e686;
  wire v3766c7b;
  wire v377226d;
  wire v3751719;
  wire v3a65e9a;
  wire v3a71614;
  wire v3731381;
  wire v37634cf;
  wire v3755883;
  wire v3a6f0f5;
  wire v374b5b6;
  wire v3a5d09b;
  wire v372a744;
  wire v377d545;
  wire v3a6c38a;
  wire v377bdd1;
  wire v3a5e975;
  wire v373c183;
  wire v3762a68;
  wire v377af89;
  wire v3a70bba;
  wire v3753e6f;
  wire v2acb0e4;
  wire v3772aaf;
  wire v374ab03;
  wire v3a672a8;
  wire v3a7006d;
  wire v3a5877f;
  wire v3a6f526;
  wire v37358f3;
  wire v3773c40;
  wire v3a6ef70;
  wire v3a6fe8c;
  wire a1b632;
  wire v38099a4;
  wire v964c47;
  wire v1e3824a;
  wire v3774829;
  wire v3a60d11;
  wire v3a6fd75;
  wire v374ea29;
  wire v3732c0d;
  wire v372ef3e;
  wire v375afbf;
  wire v3774550;
  wire v376e06b;
  wire v3725f48;
  wire v3a70e36;
  wire v3a70a43;
  wire v3a67e79;
  wire v3764809;
  wire v37711c3;
  wire v3772962;
  wire v37243e6;
  wire v3a6f22e;
  wire v3775de3;
  wire v3764462;
  wire v3a2abd2;
  wire v3751359;
  wire v372386d;
  wire v37280c8;
  wire v3755026;
  wire v374cf20;
  wire v3a70f26;
  wire v374270e;
  wire v3a69ca2;
  wire v376d98d;
  wire v3723be4;
  wire v3a6f1a6;
  wire v1e37bdd;
  wire v372b6c4;
  wire v372989c;
  wire v3a56593;
  wire v3a69bbd;
  wire v3758850;
  wire v3727e66;
  wire v375945f;
  wire v377f486;
  wire v373ce49;
  wire v3744637;
  wire v373d032;
  wire v37647ce;
  wire v3a7112a;
  wire v3751913;
  wire v37429c2;
  wire v3a6f65e;
  wire v3a6b100;
  wire v3747926;
  wire v37697ca;
  wire v3a60c4f;
  wire v3a5fa82;
  wire v3a299f8;
  wire v3a7047b;
  wire v3a639a1;
  wire v37717ea;
  wire v37656be;
  wire v3a6fdca;
  wire v372d5ba;
  wire v3759e04;
  wire v3776cad;
  wire v374e985;
  wire v3a60888;
  wire v2acaeeb;
  wire v3725bdd;
  wire v3a70ad1;
  wire v35b7d97;
  wire v3762817;
  wire v372b689;
  wire v3a6fa56;
  wire v3a6f6dd;
  wire v3a6ec1b;
  wire v3a7092b;
  wire v374a526;
  wire b15d44;
  wire v3903ee6;
  wire v3806640;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hbusreq2_p;
  input hbusreq2;
  reg hlock2_p;
  input hlock2;
  reg hbusreq3_p;
  input hbusreq3;
  reg hlock3_p;
  input hlock3;
  reg hbusreq4_p;
  input hbusreq4;
  reg hlock4_p;
  input hlock4;
  reg hbusreq5_p;
  input hbusreq5;
  reg hlock5_p;
  input hlock5;
  reg hbusreq6_p;
  input hbusreq6;
  reg hlock6_p;
  input hlock6;
  reg hbusreq7_p;
  input hbusreq7;
  reg hlock7_p;
  input hlock7;
  reg hbusreq8_p;
  input hbusreq8;
  reg hlock8_p;
  input hlock8;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmaster1_p;
  output hmaster1;
  reg hmaster2_p;
  output hmaster2;
  reg hmaster3_p;
  output hmaster3;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg hgrant2_p;
  output hgrant2;
  reg hgrant3_p;
  output hgrant3;
  reg hgrant4_p;
  output hgrant4;
  reg hgrant5_p;
  output hgrant5;
  reg hgrant6_p;
  output hgrant6;
  reg hgrant7_p;
  output hgrant7;
  reg hgrant8_p;
  output hgrant8;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg stateG10_2_p;
  output stateG10_2;
  reg stateG10_3_p;
  output stateG10_3;
  reg stateG10_4_p;
  output stateG10_4;
  reg stateG10_5_p;
  output stateG10_5;
  reg stateG10_6_p;
  output stateG10_6;
  reg stateG10_7_p;
  output stateG10_7;
  reg stateG10_8_p;
  output stateG10_8;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;
  reg jx2_p;
  output jx2;
  reg jx3_p;
  output jx3;

assign v3a701f0 = hmaster3_p & v3a61123 | !hmaster3_p & v3765324;
assign v3727580 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3747a0e;
assign v372a450 = hmaster2_p & v375e53a | !hmaster2_p & v3760513;
assign a8afe1 = hgrant2_p & v8455ab | !hgrant2_p & v375a235;
assign v3756eaf = hbusreq6_p & v3a6eb44 | !hbusreq6_p & v8455b0;
assign v376f4a6 = hmaster0_p & v8455ab | !hmaster0_p & v375e52f;
assign v3a541ec = hmaster0_p & v375646d | !hmaster0_p & v3a5524f;
assign v3770c66 = hlock6 & v3759d78 | !hlock6 & v3a6f4bc;
assign v3a544c4 = hlock8 & v3a5c40e | !hlock8 & v3757a2b;
assign v373d753 = hbusreq4 & v376b1be | !hbusreq4 & v3778f6c;
assign v38073e8 = hmaster0_p & v3a7162a | !hmaster0_p & v3a6fb81;
assign v377a7d7 = hburst0 & v3a6ac26 | !hburst0 & v372b982;
assign v375d1a6 = hgrant6_p & v377938d | !hgrant6_p & v373e10c;
assign v3724c95 = hbusreq0_p & v37621ee | !hbusreq0_p & v3a706c7;
assign v3751e5e = hbusreq6 & v376f501 | !hbusreq6 & v372462b;
assign v3a703c9 = hbusreq7 & v3734041 | !hbusreq7 & !v8455ab;
assign v3a70062 = hgrant6_p & v377e13b | !hgrant6_p & !v3a62a71;
assign v3750375 = hlock5 & v37558d3 | !hlock5 & v3a6f47a;
assign v3728870 = hmaster1_p & v3728903 | !hmaster1_p & v374bd4a;
assign dc33c0 = hgrant5_p & v3a635b1 | !hgrant5_p & b02944;
assign v37512dc = hlock4 & v372ead6 | !hlock4 & v37667b3;
assign v3753189 = hbusreq0_p & v35b774b | !hbusreq0_p & v9ed516;
assign v3a6fc6d = hmaster1_p & v3a6e31f | !hmaster1_p & v3a67315;
assign v3a6f776 = busreq_p & v3a715fd | !busreq_p & !v3a5ead2;
assign v373d4d1 = hmaster0_p & v3723185 | !hmaster0_p & v3769f01;
assign v37533ac = hgrant0_p & v8455ab | !hgrant0_p & v3760d83;
assign v377c690 = hbusreq5 & v372aa71 | !hbusreq5 & v375abdb;
assign be0bbd = hlock4_p & v3a624da | !hlock4_p & v35772a6;
assign v3a5b4de = hlock6 & v3a6fa76 | !hlock6 & v3809de2;
assign v376ba2b = hmaster2_p & v3a635ea | !hmaster2_p & v3740d3b;
assign v376a7bf = jx0_p & v37667e4 | !jx0_p & v375e91e;
assign v8e3f65 = hbusreq8_p & v360cffa | !hbusreq8_p & v3761727;
assign v3764463 = locked_p & v3771ae3 | !locked_p & !v8455ab;
assign v372d9e8 = hmaster0_p & v3a6fe18 | !hmaster0_p & v3752ade;
assign v375bdd6 = hbusreq8 & v3a5d20a | !hbusreq8 & v3757dd4;
assign v3a7066b = hmaster0_p & v3a58ef3 | !hmaster0_p & v3a70641;
assign v3747453 = hlock5_p & v906a66 | !hlock5_p & v3751285;
assign v376b0d6 = hbusreq3_p & v3a7083e | !hbusreq3_p & v8455ab;
assign v376fcc3 = hbusreq2_p & v3a70e33 | !hbusreq2_p & !v8455ab;
assign v3a6123a = hgrant0_p & v376c03e | !hgrant0_p & a38ed7;
assign v3a6cb4e = hlock0 & v373f3b5 | !hlock0 & v3a714e1;
assign v1e3731f = stateG10_1_p & v3a5deb7 | !stateG10_1_p & !v3a71109;
assign v3a6eb8f = hbusreq8 & v3a62a14 | !hbusreq8 & v372e550;
assign v9773b9 = hbusreq4 & v3773bb0 | !hbusreq4 & v8455ab;
assign v3744e13 = hmaster2_p & v35772a6 | !hmaster2_p & v3a62a08;
assign v3754eb1 = hlock2_p & v373b983 | !hlock2_p & v37592d6;
assign v372ad53 = hbusreq3_p & v3a710bc | !hbusreq3_p & v3743824;
assign v3a5f453 = hbusreq5 & v3a6fd64 | !hbusreq5 & !v3a713ab;
assign v373d66c = hmaster0_p & v3a70ddd | !hmaster0_p & v375d2b3;
assign v37266e1 = hbusreq0_p & v372b351 | !hbusreq0_p & bef73a;
assign v374f304 = hbusreq4_p & v372d9ad | !hbusreq4_p & v3a6eb1d;
assign v375be9f = hlock5_p & v8455ab | !hlock5_p & v3a6fcb2;
assign ce4c9b = hgrant6_p & v8455ab | !hgrant6_p & v3a6f1f2;
assign v3727b03 = hbusreq4_p & v37617ef | !hbusreq4_p & v35772a6;
assign v377efe7 = hmaster0_p & v375058e | !hmaster0_p & v3775928;
assign v3752304 = hbusreq6_p & v373142a | !hbusreq6_p & !v3a6fdae;
assign v3724d99 = hbusreq0 & v3a6cdd4 | !hbusreq0 & v373b0be;
assign v376a936 = hbusreq3 & v373b197 | !hbusreq3 & v8455ab;
assign v376cc20 = hbusreq3_p & v372d8fa | !hbusreq3_p & v8455ab;
assign v372354b = hbusreq5 & v374d255 | !hbusreq5 & v3a6eaf8;
assign v376730e = hbusreq6 & v3a6fdc9 | !hbusreq6 & !v8455b5;
assign v375f2c7 = hlock7 & v3742a8e | !hlock7 & v3a70d36;
assign v3764ac0 = hbusreq6 & v3a5a2e4 | !hbusreq6 & v3a56e79;
assign v3a67524 = hbusreq5_p & v376f45b | !hbusreq5_p & v3a5bb85;
assign v376e954 = hbusreq7_p & v3a6f7b8 | !hbusreq7_p & v3777474;
assign v3726ba5 = hbusreq5_p & v3738ab6 | !hbusreq5_p & v39eb3d2;
assign v37365c6 = hbusreq5_p & v3756012 | !hbusreq5_p & v37265c1;
assign v37392d7 = hbusreq8_p & v3a6a5a8 | !hbusreq8_p & v3743477;
assign v37487a6 = hbusreq7 & v3753231 | !hbusreq7 & v3a6c81d;
assign v373173b = hbusreq5_p & v3a5c3a0 | !hbusreq5_p & v3731a49;
assign a875ea = hbusreq2 & v372dccf | !hbusreq2 & v3a69487;
assign v3a70988 = hgrant2_p & v8455ab | !hgrant2_p & v377340e;
assign v3a6c33a = hbusreq2_p & v37455c2 | !hbusreq2_p & v377c5c2;
assign v2ff8bb1 = hgrant5_p & v3a6f54f | !hgrant5_p & v3a68ad7;
assign v37356cc = hbusreq4_p & v39a5265 | !hbusreq4_p & v8455e1;
assign v376d3d1 = hgrant6_p & v3a6c7fe | !hgrant6_p & v3762d3e;
assign v377e14d = hbusreq2 & v372bf87 | !hbusreq2 & v3755bc2;
assign d305e8 = hbusreq6_p & v3747302 | !hbusreq6_p & v3775d04;
assign v374af1f = hbusreq8 & v3a6f8b5 | !hbusreq8 & v8455ab;
assign v3a5b960 = hlock7 & v37325b9 | !hlock7 & v3a70b20;
assign v3739ca5 = hbusreq6_p & v375b16e | !hbusreq6_p & !v3768be2;
assign v3a68c72 = hbusreq4_p & v3a608fe | !hbusreq4_p & !v8455c2;
assign v373df21 = hready & v3a6f113 | !hready & !v8455ab;
assign v373f4dd = hbusreq5_p & v3a7122f | !hbusreq5_p & v3a71372;
assign v3a6efef = hbusreq0 & v372567b | !hbusreq0 & v3a62b11;
assign v3a59c91 = hmaster0_p & v372ff6d | !hmaster0_p & v377904f;
assign v38072fb = hbusreq6_p & v337897a | !hbusreq6_p & v3731e60;
assign v377b3a2 = hmaster1_p & v3772b8a | !hmaster1_p & v37249ff;
assign v373e2f2 = hbusreq8_p & v3a70578 | !hbusreq8_p & v3a7050f;
assign v37583f2 = hgrant1_p & v375a268 | !hgrant1_p & v377d320;
assign v3a5c7a8 = hlock4_p & v3770559 | !hlock4_p & v35772a6;
assign v92c996 = hmaster0_p & v37261be | !hmaster0_p & !v37590f4;
assign v373ef4b = hburst0 & v8455ab | !hburst0 & !v3740690;
assign v374ddc7 = hmaster0_p & v374502e | !hmaster0_p & v37471a7;
assign v373b17c = hgrant0_p & v8455ab | !hgrant0_p & v3767c44;
assign v37447e9 = hgrant4_p & v8455c2 | !hgrant4_p & v376051c;
assign v3a63873 = hlock0 & v3763209 | !hlock0 & v373e4db;
assign v3738b0f = hbusreq8 & v3a58b04 | !hbusreq8 & v3a6bba5;
assign v375c75c = hbusreq0 & v3748560 | !hbusreq0 & v3a6b18b;
assign bdb538 = hlock5_p & v3754a39 | !hlock5_p & !v8455d9;
assign v3a693dc = hmaster1_p & v373b747 | !hmaster1_p & v3724b5a;
assign v373946b = hbusreq5 & v3a6fa53 | !hbusreq5 & v3a62a6d;
assign v3a6256a = hmaster0_p & v375d0d2 | !hmaster0_p & v3a7163a;
assign v3a53c63 = hmaster2_p & v37390c5 | !hmaster2_p & v375efa4;
assign v3a6cf18 = hgrant1_p & v3a6ffae | !hgrant1_p & v3a57330;
assign v3767b70 = hbusreq0 & v3773ee6 | !hbusreq0 & v8455ab;
assign v37416b5 = hlock1 & v373dd8a | !hlock1 & v3a6a195;
assign v372fc7e = hgrant5_p & v374f0f1 | !hgrant5_p & v3a5ebc8;
assign v936e47 = hbusreq6_p & v3730646 | !hbusreq6_p & v3a541ee;
assign v9aa8f3 = hbusreq3_p & v3a704b1 | !hbusreq3_p & v37459dd;
assign v3732f00 = hlock1_p & v3a653e4 | !hlock1_p & !v8455ab;
assign stateG3_0 = !v2ff87db;
assign v3773b66 = hbusreq8 & v376e507 | !hbusreq8 & v372fdd0;
assign v372b373 = hgrant3_p & v3a7082a | !hgrant3_p & v3806388;
assign v372b89e = hlock2 & v374355d | !hlock2 & v372d078;
assign v3774e4f = hmaster2_p & v3a6f501 | !hmaster2_p & v3761175;
assign v375d364 = hlock5 & v3725c6c | !hlock5 & v3738f30;
assign v3774000 = hgrant6_p & v3729214 | !hgrant6_p & v3a711a4;
assign v373b381 = hbusreq6_p & v3a6efe8 | !hbusreq6_p & v373edbe;
assign v3759172 = hmaster2_p & v3736afd | !hmaster2_p & v3a710c8;
assign v3775cc9 = hbusreq7 & v8455ab | !hbusreq7 & v376e66e;
assign v372efb4 = hbusreq0 & v37346dc | !hbusreq0 & v3752556;
assign v3a6efc6 = hbusreq3_p & v3a5891c | !hbusreq3_p & !v3809adf;
assign v376d285 = hbusreq6_p & v3759032 | !hbusreq6_p & v3733e9e;
assign v374611e = hbusreq6_p & v3a70a05 | !hbusreq6_p & v374ea27;
assign v3732aab = hready_p & v3a70dc1 | !hready_p & !v374b64d;
assign v3a66447 = hbusreq0_p & v20d166d | !hbusreq0_p & v3751db0;
assign v3749a06 = hmaster0_p & v372ddf8 | !hmaster0_p & v37384a3;
assign v3a6dae5 = hbusreq6_p & v374faa9 | !hbusreq6_p & v3767266;
assign v3767dac = jx1_p & v380a20c | !jx1_p & v3a66a86;
assign v3746496 = hmaster2_p & v8455cb | !hmaster2_p & v3737d38;
assign v37729ac = hbusreq3 & v3750037 | !hbusreq3 & v8455ab;
assign v3778b60 = hbusreq4_p & v377818c | !hbusreq4_p & v8455ab;
assign d8a75b = hlock1 & v3a6d5b3 | !hlock1 & v3a5ef54;
assign v3a5d763 = hmaster2_p & v372455c | !hmaster2_p & v3a70e2e;
assign v3769cc4 = hbusreq5 & v3a7017d | !hbusreq5 & v2925d03;
assign v376f45b = hbusreq5 & v3a6d6ff | !hbusreq5 & v37756ef;
assign v37654ea = hbusreq7_p & v3a6d4f8 | !hbusreq7_p & v3a6f8ef;
assign v3746818 = hbusreq5 & v3729fa4 | !hbusreq5 & v374dfad;
assign v9e8a9c = hmaster2_p & v35772b3 | !hmaster2_p & v3a642cf;
assign v3a63a2a = hbusreq2 & v3a5610f | !hbusreq2 & v38072fd;
assign v3a6f259 = hmaster1_p & v374156a | !hmaster1_p & v37675f1;
assign v374306c = locked_p & v3a6f210 | !locked_p & v3a6ffae;
assign v373301d = hbusreq2_p & v3a713e3 | !hbusreq2_p & v3a53dbf;
assign v3774dbe = hbusreq2_p & v3748ca5 | !hbusreq2_p & v376f5e1;
assign v37724f9 = hgrant6_p & v8455ab | !hgrant6_p & v37282ac;
assign v3748ab9 = hmaster1_p & v377dbd3 | !hmaster1_p & v9ca2d6;
assign v3760748 = hbusreq4_p & v373fd72 | !hbusreq4_p & v376c687;
assign v3769adb = hmaster0_p & v3767b70 | !hmaster0_p & v3766dcc;
assign v37244b9 = hbusreq7_p & v37596f3 | !hbusreq7_p & v8455c7;
assign v3740466 = hlock5 & v3a6ae0f | !hlock5 & v3770425;
assign v3771252 = hmaster1_p & v3775942 | !hmaster1_p & !v376abdf;
assign v3763478 = hbusreq5 & v3730688 | !hbusreq5 & v3a62f50;
assign v373a7a5 = hgrant4_p & v377b946 | !hgrant4_p & v373eaee;
assign v380946e = hbusreq8_p & v2acb0b1 | !hbusreq8_p & v3761f2b;
assign v376a95c = hbusreq2_p & v377773f | !hbusreq2_p & v8455ab;
assign v3748d67 = hbusreq3_p & v3747302 | !hbusreq3_p & v3743b9e;
assign v3a62fa7 = hbusreq6 & v3a710e4 | !hbusreq6 & v3a6f71a;
assign v375df4f = hbusreq8_p & v3a6f2f8 | !hbusreq8_p & v374e620;
assign v376b2e9 = hbusreq0_p & v3a6143b | !hbusreq0_p & !v39a4ca8;
assign v373e491 = jx0_p & v37684c0 | !jx0_p & v3a6f6f8;
assign v3729a9f = hbusreq1_p & v3727f86 | !hbusreq1_p & !v373f56b;
assign v3807ac6 = hbusreq2_p & v372a786 | !hbusreq2_p & v372eecf;
assign v3734af2 = hbusreq2_p & adf78a | !hbusreq2_p & v3753dab;
assign v373e37c = hbusreq3_p & v376ef42 | !hbusreq3_p & v3a70c07;
assign v37302fb = hmaster1_p & v3757100 | !hmaster1_p & v374f526;
assign v373a8c0 = hmaster0_p & v360d1b0 | !hmaster0_p & v3a70fae;
assign v3744a21 = hgrant4_p & v3a6fcae | !hgrant4_p & v1e37442;
assign v3738906 = hmaster2_p & v1e37489 | !hmaster2_p & v3728d9c;
assign v375b269 = hgrant3_p & v37669b4 | !hgrant3_p & v3765a43;
assign v377094d = hmaster2_p & v3a6fdd6 | !hmaster2_p & v37369b2;
assign v3779fbd = hgrant0_p & v3724940 | !hgrant0_p & v8455ab;
assign v3a70b85 = hlock8 & v3737808 | !hlock8 & v3758357;
assign v376245d = hlock6_p & v376d240 | !hlock6_p & v372d96e;
assign v3a6fd24 = hlock5_p & v3755002 | !hlock5_p & !v8455ab;
assign v377723a = hbusreq4 & v3769a1e | !hbusreq4 & v373abde;
assign v3a6f57c = hbusreq4_p & v3a709a6 | !hbusreq4_p & v380a188;
assign v3767ef0 = hmaster0_p & v37245f8 | !hmaster0_p & v37512b3;
assign v3740951 = hmaster2_p & v8455ab | !hmaster2_p & !v376aa98;
assign v3a703ab = hmaster1_p & v3779403 | !hmaster1_p & v3a62ad8;
assign v375daac = hmaster2_p & v3771a80 | !hmaster2_p & v3a691eb;
assign v3746406 = hmaster0_p & v37295e7 | !hmaster0_p & v3728cdc;
assign v37518e7 = hmaster0_p & v374bab6 | !hmaster0_p & v37782de;
assign v37240e6 = hbusreq6_p & v37535bd | !hbusreq6_p & v3728cd0;
assign v375ff98 = hgrant2_p & v3a6db06 | !hgrant2_p & v3a638e9;
assign v3731ed2 = hbusreq3 & v37508a4 | !hbusreq3 & v8455ab;
assign v3a70e42 = hmaster1_p & v35b7b3b | !hmaster1_p & v8a7af6;
assign v372ccbe = hbusreq4_p & v3806ce9 | !hbusreq4_p & v8455bf;
assign v3a5e618 = hbusreq5 & v376dc6f | !hbusreq5 & v3a5e030;
assign v3a56c2e = hlock6 & v375c9ea | !hlock6 & v374cf79;
assign v3747fd2 = hbusreq5_p & v3736a50 | !hbusreq5_p & v3a5d644;
assign v3a5cdef = hbusreq5_p & v3a5df66 | !hbusreq5_p & v375ede6;
assign v37440c3 = hmastlock_p & v3a5ff81 | !hmastlock_p & v8455ab;
assign v3737411 = hbusreq7 & v374b40e | !hbusreq7 & v3a5897a;
assign v377c29b = hmaster3_p & v377541e | !hmaster3_p & v3a5857e;
assign v372fc17 = hmastlock_p & v8455ff | !hmastlock_p & !v8455ab;
assign v3761334 = hmaster0_p & v372ff09 | !hmaster0_p & v37584e6;
assign v3762fc2 = hbusreq3_p & v2092ffc | !hbusreq3_p & bdda12;
assign v372d9e0 = hbusreq6_p & v3a704ee | !hbusreq6_p & v3750134;
assign v377de50 = hmaster2_p & v373afc3 | !hmaster2_p & v3738169;
assign v3a6ebf8 = hlock6 & v3743dae | !hlock6 & v3a70734;
assign v3a6a990 = hlock5_p & v372fe58 | !hlock5_p & v376581d;
assign v3764f8a = hbusreq0_p & v37682a8 | !hbusreq0_p & v35772a6;
assign v3a5e1bc = hbusreq6_p & v372d630 | !hbusreq6_p & v373ec0f;
assign v3a6f1ef = hlock8_p & v37726d9 | !hlock8_p & !v8455ab;
assign v376905f = hlock3 & v3743366 | !hlock3 & v3a6f77c;
assign v3772d2f = hbusreq8 & v3776395 | !hbusreq8 & v3a67b58;
assign busreq = v23fdb05;
assign v372efcd = hmaster2_p & v3769921 | !hmaster2_p & v377d1dc;
assign v3a6e93d = hmaster2_p & v3a6fff0 | !hmaster2_p & v3732c72;
assign v3779ac0 = hbusreq5_p & v8d2bbf | !hbusreq5_p & !v375931f;
assign v373578d = hmaster1_p & v3a6f781 | !hmaster1_p & v3779491;
assign v3a700a5 = locked_p & v3a61254 | !locked_p & v3807bf8;
assign v3735ec7 = hmaster2_p & v3a5e24e | !hmaster2_p & !v37745a0;
assign v373a07f = hbusreq0_p & v8455e7 | !hbusreq0_p & v3751c87;
assign v3a70d66 = hbusreq0 & v3a6b97b | !hbusreq0 & !v374f9f5;
assign v3a70afe = hmaster2_p & v2aca977 | !hmaster2_p & v372a4c1;
assign v372df43 = hbusreq6_p & v38072fd | !hbusreq6_p & v3a6a236;
assign v3a55456 = hbusreq0 & v373fe5e | !hbusreq0 & v8455e7;
assign v3809487 = hbusreq4_p & v377b0a0 | !hbusreq4_p & v3a702a8;
assign v374a668 = hmaster2_p & v2acafcc | !hmaster2_p & v3a6fa8e;
assign v3a6469c = hlock0_p & v37583be | !hlock0_p & v8455ab;
assign v3a62949 = hlock5_p & v37249c7 | !hlock5_p & !v3a71541;
assign v3759edb = hlock4 & v374e353 | !hlock4 & v3a6f0e9;
assign v37229b8 = hgrant6_p & v377b6ce | !hgrant6_p & v35b7189;
assign v374f78c = hbusreq3_p & v2aca770 | !hbusreq3_p & v8455b0;
assign v3a6fd90 = hbusreq7_p & v372fe57 | !hbusreq7_p & v376db6d;
assign v37705df = hbusreq5 & v374b887 | !hbusreq5 & v3a5fc48;
assign v37599b1 = hlock1 & v374197c | !hlock1 & v3a70a12;
assign v375a76e = hmaster1_p & v377c7c0 | !hmaster1_p & v377bd17;
assign v3a69feb = hmaster3_p & v3a6fd86 | !hmaster3_p & v3a62e7b;
assign v3725367 = hbusreq8 & v3a6c2d2 | !hbusreq8 & v3777312;
assign v375dc75 = hbusreq5_p & v373cdba | !hbusreq5_p & v3722fc5;
assign v374a650 = hmaster0_p & v372d905 | !hmaster0_p & v37367e3;
assign v372ee6a = hmaster2_p & v3a60077 | !hmaster2_p & v3a5b68a;
assign v8615d7 = hbusreq2 & v374362e | !hbusreq2 & !v3a568f7;
assign v373e419 = hmaster3_p & v375f42e | !hmaster3_p & v3a6f298;
assign v2092aba = hlock6_p & v373aed4 | !hlock6_p & v8455bf;
assign cfaa3a = hmaster0_p & v3763a20 | !hmaster0_p & v377bbf7;
assign v3a70dca = hlock5_p & v3a58967 | !hlock5_p & v3779b9c;
assign a25d5b = hgrant6_p & v3a6ab8c | !hgrant6_p & v374fda4;
assign v3a5c73c = hbusreq5 & v940c77 | !hbusreq5 & aa8b86;
assign v37404d0 = hmaster0_p & v3a70da4 | !hmaster0_p & v377ce5e;
assign v377ce3f = hmaster2_p & v3a635ea | !hmaster2_p & v375da10;
assign v3725931 = hbusreq4 & v3a56e63 | !hbusreq4 & !v8455ab;
assign v3a70ba1 = hmaster0_p & v374db8d | !hmaster0_p & v376363f;
assign v374c936 = hbusreq1_p & v3a70c73 | !hbusreq1_p & !v373e16a;
assign v376e772 = hbusreq0 & v3a636fe | !hbusreq0 & v3746f46;
assign v376e041 = hbusreq3_p & v3747302 | !hbusreq3_p & v37496fa;
assign v375e2d3 = hgrant3_p & v3a5c945 | !hgrant3_p & v376d28f;
assign v3725cbf = hgrant0_p & v8455ab | !hgrant0_p & v3a5e3d3;
assign v374e6ec = hgrant3_p & v372ffd2 | !hgrant3_p & v3729513;
assign v1e37af7 = hbusreq7 & v373f909 | !hbusreq7 & v3765e47;
assign v372c219 = hgrant6_p & v377f09a | !hgrant6_p & v376fe88;
assign v372d608 = hbusreq2 & v37288b6 | !hbusreq2 & v372e83f;
assign v38097a9 = hbusreq0 & v3730d6a | !hbusreq0 & v3723400;
assign v3749c4b = hbusreq4_p & v3a6814a | !hbusreq4_p & !v3a672c9;
assign v375f74a = hlock0_p & v373997b | !hlock0_p & v3a6143b;
assign v3774c77 = hlock6 & v377476b | !hlock6 & v375859f;
assign v37664aa = hbusreq7_p & v3764ef1 | !hbusreq7_p & !v377adbd;
assign v373ea10 = hbusreq4_p & v380678d | !hbusreq4_p & v3809ec3;
assign v3a71456 = hgrant1_p & v3a57445 | !hgrant1_p & v37271f9;
assign v3a5e3bb = hbusreq3_p & v2092ffc | !hbusreq3_p & v3726006;
assign v376fed4 = hlock7_p & v374f0f1 | !hlock7_p & !v377478a;
assign v373601e = hbusreq6 & v3734db5 | !hbusreq6 & v3765e79;
assign v372eb1a = hbusreq4 & v3727580 | !hbusreq4 & v3a5fc82;
assign v3739190 = hbusreq4_p & v3a66e96 | !hbusreq4_p & v375af58;
assign v37368bb = hbusreq7 & v3a7059e | !hbusreq7 & v3a2951d;
assign v3a707c5 = hbusreq5_p & v37307a7 | !hbusreq5_p & v9e8d30;
assign v374c8a8 = hmaster2_p & v375f619 | !hmaster2_p & v3746540;
assign v3a6fc17 = hbusreq3_p & v375bdd4 | !hbusreq3_p & v8455e1;
assign v3730688 = hmaster0_p & v37338bb | !hmaster0_p & v3a7090f;
assign v377598a = hmaster2_p & v3a6d684 | !hmaster2_p & v37432c6;
assign v3a67257 = hbusreq4_p & v372e562 | !hbusreq4_p & v3757a57;
assign v9f56fd = hbusreq8_p & v3728382 | !hbusreq8_p & v8455ab;
assign v1e37e04 = hmaster3_p & v8455ab | !hmaster3_p & v38074c0;
assign v37398eb = hlock2 & v3a618b3 | !hlock2 & v376a34d;
assign v3a70403 = hbusreq2_p & v3a6962d | !hbusreq2_p & v3754871;
assign v375d3da = jx0_p & v3738a5e | !jx0_p & v3748256;
assign v3808fc2 = hgrant2_p & v8455ab | !hgrant2_p & v3753b90;
assign v372a1b4 = hbusreq6_p & v8455ab | !hbusreq6_p & v8455b9;
assign v3a6c803 = hmaster2_p & v3730755 | !hmaster2_p & v375a4fa;
assign v3740c94 = hbusreq7 & v3a6cc2a | !hbusreq7 & v37612a3;
assign v2acaed3 = hlock4 & v373fde6 | !hlock4 & v373a6c8;
assign v373d12a = hbusreq0 & v372af57 | !hbusreq0 & v3723dac;
assign v375e356 = hlock0 & v3759361 | !hlock0 & v373ace1;
assign v376c3c2 = jx1_p & v374b237 | !jx1_p & !v3753198;
assign v3a6a197 = hmaster2_p & v3a5b8b9 | !hmaster2_p & v3763fdc;
assign v3a70322 = hlock4 & v373f6d5 | !hlock4 & v3a5dc82;
assign v3777adb = hlock4_p & v375e682 | !hlock4_p & !v8455ab;
assign v3a6fba8 = hlock4 & v3a709ba | !hlock4 & v374291b;
assign v3742a4d = hbusreq7 & v3a53977 | !hbusreq7 & v3a6fba3;
assign v376b654 = hmaster0_p & v375a3dd | !hmaster0_p & v373cde7;
assign v3744982 = hlock1_p & v37418b3 | !hlock1_p & !v8455ab;
assign v37336b4 = hlock8 & v3a711be | !hlock8 & v377b481;
assign v377670f = stateA1_p & v8455ab | !stateA1_p & v3726dfa;
assign v3727387 = hbusreq5_p & v3a706d9 | !hbusreq5_p & v37390f0;
assign v3746cc3 = hgrant5_p & v3a69f4e | !hgrant5_p & !v8455ab;
assign v3a6f84d = hgrant1_p & v375cd0c | !hgrant1_p & v37328bf;
assign v372ec4e = hbusreq4_p & v38097db | !hbusreq4_p & v3a64374;
assign v37484ac = hlock5 & v372bcd3 | !hlock5 & v37713e8;
assign v882147 = hmaster2_p & v374e855 | !hmaster2_p & v3a5c640;
assign v3a6c628 = hmaster2_p & v3a70a7f | !hmaster2_p & v3779cf9;
assign v3a7142f = hgrant4_p & v3a70d99 | !hgrant4_p & v3a6faef;
assign v3723400 = hgrant6_p & v1e37cd6 | !hgrant6_p & v3809d6a;
assign v372ea9b = hgrant4_p & v3a70363 | !hgrant4_p & v3a6fbca;
assign v3745291 = hlock3_p & v3a64fe0 | !hlock3_p & v377e08c;
assign v373a59e = hmaster1_p & v376ccd6 | !hmaster1_p & v3a5e7f7;
assign v3a69727 = hgrant4_p & v8455ab | !hgrant4_p & !v3769f5f;
assign v3a6fc1d = hlock4 & v37458d2 | !hlock4 & v3a6dbf0;
assign v3a62fc9 = hmaster1_p & v3758b45 | !hmaster1_p & v3a56827;
assign v3766830 = jx0_p & v3a68af5 | !jx0_p & v8455ab;
assign v377f2a9 = hgrant4_p & v3a53eeb | !hgrant4_p & v3a5986c;
assign v377168f = jx0_p & v374c154 | !jx0_p & v376614e;
assign v372afe7 = hmaster0_p & v3a70fd6 | !hmaster0_p & v3a59ea2;
assign v3a693bf = hlock1_p & v374c1c3 | !hlock1_p & !v8455ab;
assign v376944c = hbusreq6 & v377928c | !hbusreq6 & v8455ab;
assign v3a65c47 = hbusreq8_p & v3a5be8a | !hbusreq8_p & c39ea5;
assign v37423d1 = hbusreq4_p & v3a70d99 | !hbusreq4_p & v2ff9314;
assign v3a61739 = hbusreq0 & v375a2b5 | !hbusreq0 & v3751073;
assign v372f5e7 = hgrant1_p & v372af91 | !hgrant1_p & v8455e7;
assign v3a5d185 = hmaster1_p & v3778fb5 | !hmaster1_p & v373fb22;
assign v3a6edfa = hburst0 & v3a64235 | !hburst0 & v8455ab;
assign v3a66b2b = hlock0_p & v3a635ea | !hlock0_p & !v374bae0;
assign v3a56d0a = hgrant2_p & v3a5e3c0 | !hgrant2_p & v376daf6;
assign v3a70547 = hgrant0_p & v3753e6a | !hgrant0_p & v3738de9;
assign v374fc82 = hgrant4_p & v1e37b99 | !hgrant4_p & v3a7088d;
assign v3a6fdb1 = hbusreq7 & v376610a | !hbusreq7 & v8455ab;
assign v3a6fa41 = hbusreq5 & v376ee43 | !hbusreq5 & v374ae7a;
assign v3a67b86 = hbusreq6 & v3a69488 | !hbusreq6 & v23fd967;
assign v3a7153a = hbusreq1_p & v376b47d | !hbusreq1_p & v8455ab;
assign v37439b2 = hgrant2_p & v8455ab | !hgrant2_p & v374d218;
assign v3a700ab = hready_p & v3763f05 | !hready_p & v39a4ce0;
assign v37328b0 = hmaster2_p & v35772a2 | !hmaster2_p & v377928c;
assign v3755c7c = hbusreq2_p & v372ccbb | !hbusreq2_p & v3809f65;
assign v3a5ed4a = hmaster2_p & v372cfeb | !hmaster2_p & v3775626;
assign v3776715 = hgrant4_p & v8455ab | !hgrant4_p & v37272df;
assign v37326be = hbusreq8_p & v3777239 | !hbusreq8_p & ae60a0;
assign v372b24d = hburst1 & v3a6ac26 | !hburst1 & v377a7d7;
assign v3735974 = hmaster2_p & v8455b7 | !hmaster2_p & v8455ab;
assign v37654e0 = hmaster0_p & v3a5c6d0 | !hmaster0_p & v377c065;
assign v3750f27 = hbusreq5 & v3756809 | !hbusreq5 & v2925d06;
assign v3724028 = hbusreq5 & v375f963 | !hbusreq5 & v3a6fb73;
assign v35b70c3 = hmaster1_p & v3a661fe | !hmaster1_p & v3772bb3;
assign v37782de = hmaster2_p & v3774bad | !hmaster2_p & v3a5c33d;
assign v373931a = hmaster2_p & v377746e | !hmaster2_p & v376dc44;
assign v3a68838 = hbusreq2_p & v3a68276 | !hbusreq2_p & v8455ab;
assign v373aee6 = hbusreq5_p & v374bff0 | !hbusreq5_p & v3725a73;
assign v375aa2d = hlock6_p & v3a64087 | !hlock6_p & v3762949;
assign v3378996 = hmaster1_p & v372f770 | !hmaster1_p & v3a6462c;
assign v3754c8d = hgrant6_p & v8455ab | !hgrant6_p & v374b923;
assign v3a5affd = hgrant3_p & v8455ab | !hgrant3_p & v372c6fb;
assign v37315c5 = hgrant4_p & v37319cd | !hgrant4_p & v37656b8;
assign v374193d = hmaster0_p & v3a6f451 | !hmaster0_p & v3a5fd4a;
assign v377b0fb = hmaster3_p & v376b94a | !hmaster3_p & v3a71592;
assign v3a6e4ec = hmaster2_p & v3a635ea | !hmaster2_p & v3748d67;
assign v3a709f0 = hgrant5_p & v376130f | !hgrant5_p & v3772afb;
assign v3a65c2a = hmaster2_p & v3728604 | !hmaster2_p & v375070c;
assign v9259bc = hbusreq8_p & v3766f13 | !hbusreq8_p & v3a56d2e;
assign v3747585 = hgrant4_p & v375c7b9 | !hgrant4_p & v3735554;
assign v3a6f781 = hgrant4_p & v8455ab | !hgrant4_p & v375ee73;
assign v375bebd = hbusreq0_p & v375fbd7 | !hbusreq0_p & v3a706c7;
assign v3762d80 = hbusreq3 & a9f66a | !hbusreq3 & v375039e;
assign v375841a = hmaster0_p & v37707b6 | !hmaster0_p & v8455ab;
assign v37316ec = hbusreq5 & v3a603c1 | !hbusreq5 & c79715;
assign v376801c = hmaster2_p & v3a6fdd6 | !hmaster2_p & v3759379;
assign v3a7145e = hgrant5_p & v8455ab | !hgrant5_p & v373357d;
assign v3a70cb3 = hbusreq7 & v3776e33 | !hbusreq7 & v3a5fc34;
assign v3753d03 = hmaster0_p & v3a658f7 | !hmaster0_p & v375449f;
assign v3757311 = hlock8 & v3a5c040 | !hlock8 & v3a5b960;
assign v3a70c59 = hmaster0_p & v3a66110 | !hmaster0_p & !v3a57f59;
assign v377903f = hgrant2_p & v3750d06 | !hgrant2_p & v3733fd8;
assign v3743de6 = hbusreq0 & v373f8f8 | !hbusreq0 & v8455ab;
assign v372a92a = hmaster2_p & v3a71678 | !hmaster2_p & v376e717;
assign v1e37776 = hmaster1_p & v3a5a510 | !hmaster1_p & v37473c5;
assign v375c976 = hgrant6_p & v8455ab | !hgrant6_p & v374fb40;
assign v3a6c82f = hlock6_p & v37388ce | !hlock6_p & v375aaca;
assign v377359f = hlock6_p & v3728e09 | !hlock6_p & !v8455ab;
assign v3a5bb64 = hlock0_p & v3747302 | !hlock0_p & v3a709ef;
assign v374282f = hbusreq2_p & v373c830 | !hbusreq2_p & !v8455ab;
assign v3a6feed = hmastlock_p & v3a61988 | !hmastlock_p & v8455ab;
assign v3722bb0 = hmaster1_p & v3a635ea | !hmaster1_p & v37512c1;
assign v1e38275 = stateA1_p & v8455ab | !stateA1_p & !v373c3bd;
assign v3a54519 = hbusreq7_p & v3a67a02 | !hbusreq7_p & v3a7075d;
assign v3777c7f = hmaster1_p & v3778cba | !hmaster1_p & v376a3f5;
assign v3a704b0 = hlock6 & v3770e30 | !hlock6 & v3a70fd2;
assign c81b97 = hmaster0_p & b88b06 | !hmaster0_p & v3a57741;
assign v375f4fd = hgrant3_p & v3a70351 | !hgrant3_p & v1e37921;
assign v3778f81 = hmaster3_p & v374d0ad | !hmaster3_p & v3763590;
assign v3a55aba = hbusreq3_p & v3a5a6db | !hbusreq3_p & v8455e7;
assign v3739fc8 = hgrant7_p & v3a6f046 | !hgrant7_p & v374494b;
assign v373ed5c = hmaster0_p & v3a59cae | !hmaster0_p & !v3a6ff47;
assign v37250af = jx2_p & v37699ec | !jx2_p & v374f12c;
assign v37595c8 = hgrant0_p & v8455ab | !hgrant0_p & v3a59883;
assign v374421d = hbusreq6_p & v37708e7 | !hbusreq6_p & v3a70889;
assign v37649a0 = hgrant6_p & v2acaf72 | !hgrant6_p & !v373b012;
assign v3a714c8 = hbusreq5 & v372b794 | !hbusreq5 & v3760bda;
assign v3776352 = hmaster1_p & v374b95f | !hmaster1_p & v376c573;
assign v3756f42 = hbusreq0 & v372bffa | !hbusreq0 & v372d967;
assign v37675e9 = hmaster0_p & v37560f1 | !hmaster0_p & v3a6a9d7;
assign v3743a8a = hlock5 & v3a6ebc7 | !hlock5 & v3258dc5;
assign v3743a4d = hlock4_p & v376c176 | !hlock4_p & !v8455ab;
assign v376db87 = hmaster2_p & v8455ab | !hmaster2_p & v372abb1;
assign v372b794 = hmaster0_p & v3a635ea | !hmaster0_p & v3a70761;
assign v3a6ffcc = hgrant6_p & v8455ab | !hgrant6_p & v3770735;
assign v3a6fe81 = hgrant5_p & v8455c6 | !hgrant5_p & v3a57fa3;
assign v3752523 = hbusreq0 & v3a66279 | !hbusreq0 & v3a622f5;
assign v3a71119 = hmaster1_p & v372b1dc | !hmaster1_p & v3a71230;
assign v3a5bbc2 = hmaster2_p & v8455ab | !hmaster2_p & v37314fc;
assign v3771a80 = hgrant4_p & v8455ab | !hgrant4_p & v3745012;
assign v944e42 = hmaster1_p & v377bb3a | !hmaster1_p & v3a5c7a6;
assign v376945e = hbusreq8 & v1e3780d | !hbusreq8 & v3a69973;
assign v3a5c2df = hbusreq6_p & v3a5d6a6 | !hbusreq6_p & v37576d1;
assign v3772f09 = hgrant7_p & v3a70c80 | !hgrant7_p & v3a6a9cd;
assign v3a70490 = hbusreq8 & v374d07a | !hbusreq8 & v3770ecc;
assign v373f909 = hmaster1_p & v8455b0 | !hmaster1_p & v3a607fa;
assign v3743d5d = hbusreq5 & v377f1ff | !hbusreq5 & v3a57ee9;
assign v39eb4d4 = hgrant2_p & v374d542 | !hgrant2_p & v3a7119e;
assign v3a60dfb = hmaster0_p & v375959a | !hmaster0_p & v3a70476;
assign v374ad17 = hmaster0_p & v37440c0 | !hmaster0_p & v374d4d3;
assign v373d99d = hbusreq2 & v376f2f8 | !hbusreq2 & v8455ab;
assign v374ce04 = hmaster1_p & v35b774b | !hmaster1_p & v37296cd;
assign v376eb3f = hlock6_p & v3725410 | !hlock6_p & v8455b7;
assign v3a708f6 = hbusreq4 & v3a6f496 | !hbusreq4 & v3a69487;
assign v3a70010 = hbusreq1 & v8455e1 | !hbusreq1 & v8455ab;
assign v3a7010e = hbusreq0 & v373f92e | !hbusreq0 & v8455ab;
assign v375a9d7 = hmaster1_p & v374a296 | !hmaster1_p & v374cab1;
assign v372ddfa = hgrant6_p & v1e37cd6 | !hgrant6_p & v376b5c6;
assign v375efe0 = hlock8_p & v3774655 | !hlock8_p & v372f05b;
assign v3735c06 = hmaster2_p & v374f87c | !hmaster2_p & v8455ab;
assign v3a6ef98 = hbusreq4_p & v374513e | !hbusreq4_p & !v37392ad;
assign v3770425 = hmaster0_p & v3a70fbf | !hmaster0_p & v3a6b4e8;
assign v377d10c = hgrant6_p & v3a5dc35 | !hgrant6_p & v376572c;
assign v3735e39 = locked_p & v3a5bd24 | !locked_p & v39a537f;
assign v3769280 = hmaster2_p & v3a6c4e4 | !hmaster2_p & v3761470;
assign dbc26f = hlock0 & v3748797 | !hlock0 & v3779008;
assign v28896cd = hbusreq5_p & v374d490 | !hbusreq5_p & !v3763cef;
assign v3a5e3f1 = hmaster0_p & v3a6d098 | !hmaster0_p & v8455e7;
assign v3a71294 = hbusreq7_p & v375c6cd | !hbusreq7_p & v3a689d1;
assign v3a675bb = hbusreq5_p & v3a625ac | !hbusreq5_p & v3a715d7;
assign v3761f78 = hbusreq5 & v37386f5 | !hbusreq5 & !v8455b9;
assign v3a66e41 = hlock4 & v3a5d06d | !hlock4 & v3764ca0;
assign v373a3c8 = hmaster2_p & v3a6b860 | !hmaster2_p & v3a66ea9;
assign v3745ce8 = hbusreq0 & v3a712d3 | !hbusreq0 & v373b286;
assign v3a715a9 = hlock4 & a53cf9 | !hlock4 & v375e12d;
assign v3722bc2 = hgrant2_p & v3a58762 | !hgrant2_p & v3727482;
assign v3a63198 = hmaster2_p & v372b6bc | !hmaster2_p & v37287d8;
assign v374efeb = hgrant8_p & v8455b5 | !hgrant8_p & v3a5f8b2;
assign v375c60f = hmaster0_p & v3a7002c | !hmaster0_p & v37587fa;
assign v375e2de = hbusreq8 & v3a71581 | !hbusreq8 & v3775d6e;
assign v375b9a3 = hmaster1_p & v376c27d | !hmaster1_p & v372d748;
assign v37fca8d = hbusreq4 & v3751d16 | !hbusreq4 & v3a63a66;
assign v3a6ef01 = hgrant4_p & v8455ab | !hgrant4_p & v3730e74;
assign v3770ad8 = hmaster0_p & v375a86a | !hmaster0_p & v37328f1;
assign v376aa5e = hlock6_p & v3770559 | !hlock6_p & v35772a6;
assign v3a709af = hbusreq6_p & v374d2b3 | !hbusreq6_p & v3a55349;
assign v3733b90 = hgrant5_p & v3723d79 | !hgrant5_p & v209306f;
assign v377b774 = hbusreq3_p & ab638b | !hbusreq3_p & v8455ab;
assign v377282c = hmaster0_p & v3743c7e | !hmaster0_p & v3a6eebb;
assign v37414be = hbusreq8_p & aeaf7c | !hbusreq8_p & v3a61b9d;
assign v3a70f63 = hmaster1_p & v3752dc7 | !hmaster1_p & v37705ec;
assign v3745b85 = start_p & v3746bdb | !start_p & v3a5a496;
assign v3741850 = hbusreq3 & v3a6d4c2 | !hbusreq3 & v8455ab;
assign v376b743 = hlock5 & v3741bd8 | !hlock5 & v33789ef;
assign v3a6cb69 = hbusreq3_p & v37b6451 | !hbusreq3_p & !v8455ab;
assign v3738750 = hbusreq5 & v3739ec6 | !hbusreq5 & v3a6f158;
assign v37586bb = hmaster0_p & v376a254 | !hmaster0_p & v37508b9;
assign v38095b1 = hbusreq5 & v3a71574 | !hbusreq5 & v3764761;
assign v3a61c5a = hlock0_p & v8455b7 | !hlock0_p & v3770187;
assign v3a6ffa9 = busreq_p & v373d9e5 | !busreq_p & !v37481c3;
assign v3763f95 = hlock4_p & v3763175 | !hlock4_p & !v8455ab;
assign v2619ada = hbusreq2_p & v38072fd | !hbusreq2_p & v373dec1;
assign v3a55755 = hbusreq6 & v3731c72 | !hbusreq6 & v8455ab;
assign v372f7b4 = hmaster1_p & v3a53e30 | !hmaster1_p & v37535d9;
assign v3a6dfec = hbusreq7 & v373f461 | !hbusreq7 & v3a5a210;
assign v37b6451 = hbusreq3 & v3a703df | !hbusreq3 & !v8455ab;
assign v37472b9 = hmaster0_p & v37356f0 | !hmaster0_p & v374a075;
assign d0c237 = hmaster2_p & v374ccb7 | !hmaster2_p & v377df2e;
assign v3756416 = hbusreq2 & v3766d04 | !hbusreq2 & v3a5affd;
assign v3735539 = hmaster0_p & v377940a | !hmaster0_p & v377e241;
assign hgrant1 = !v35b6167;
assign v3770e2b = hlock0_p & v8455ab | !hlock0_p & v3a66737;
assign v292555a = hbusreq2_p & v3a7162d | !hbusreq2_p & v3778528;
assign v37287fa = hbusreq7_p & v374fcde | !hbusreq7_p & !v372e865;
assign v3756960 = jx0_p & v8455ab | !jx0_p & v3761d7e;
assign v375a0ff = hgrant0_p & v3733090 | !hgrant0_p & v3770e2b;
assign v3751073 = hgrant6_p & v3725fe1 | !hgrant6_p & v377ce30;
assign v3762c44 = hgrant2_p & v8455ab | !hgrant2_p & !v3808cee;
assign v37676d0 = hbusreq4 & v3a55cd6 | !hbusreq4 & !v8455b5;
assign v3a70665 = hmaster2_p & v3a635ea | !hmaster2_p & v377c931;
assign v372954d = hlock5_p & v37655c5 | !hlock5_p & v8455e7;
assign v372f5ca = hmaster1_p & v3a5ab08 | !hmaster1_p & v3a5c41b;
assign v3a652c7 = hmaster2_p & v8455ab | !hmaster2_p & !v3a62396;
assign v374fe0f = hbusreq0 & v373e21a | !hbusreq0 & !v374e77f;
assign v377097e = jx0_p & v3730b3a | !jx0_p & v373fcc7;
assign v3a6fa2c = hlock2 & v3726d97 | !hlock2 & v372da76;
assign v377463d = jx0_p & v3a60fa7 | !jx0_p & !v376978e;
assign v3a6c8dc = hbusreq2 & v3a64703 | !hbusreq2 & v3a5ab6e;
assign v375d85b = hmaster3_p & v376b7a8 | !hmaster3_p & v380985a;
assign v37480a7 = hbusreq3 & v373cca3 | !hbusreq3 & v8455ab;
assign v372455c = hbusreq2_p & v377018e | !hbusreq2_p & v8455ab;
assign v3a6817a = hgrant6_p & v372aadd | !hgrant6_p & v373b666;
assign v3749cf4 = hmaster0_p & v375b0d4 | !hmaster0_p & !v2ff9391;
assign v3a70414 = hlock6 & v37305b9 | !hlock6 & v375aeca;
assign v3a6f5bf = hlock5 & v375b563 | !hlock5 & v374fab7;
assign v2889716 = hgrant2_p & v8455ab | !hgrant2_p & v376a95c;
assign v3808e56 = hbusreq7_p & a0a219 | !hbusreq7_p & v3775709;
assign v3a646ae = hbusreq4 & v372456c | !hbusreq4 & v3752cf6;
assign v376430d = hmaster0_p & v3a635ea | !hmaster0_p & v37650b8;
assign v373ca4f = hlock0_p & b0c091 | !hlock0_p & !v8455ab;
assign v3a71293 = hgrant4_p & v37615c5 | !hgrant4_p & v3a6fa3f;
assign v3739940 = hbusreq5_p & v375b787 | !hbusreq5_p & !v3a70d09;
assign v3a70147 = hgrant4_p & v8455ab | !hgrant4_p & c0b985;
assign v3740e4c = hmaster2_p & v3774276 | !hmaster2_p & be166e;
assign v372ee7e = hlock0_p & v3a70c07 | !hlock0_p & v37307de;
assign v3767e03 = hmaster1_p & v3a70cb0 | !hmaster1_p & !v3768ae9;
assign v3a67880 = hgrant7_p & v3a558be | !hgrant7_p & v372826c;
assign v375f069 = hmaster3_p & v8455ab | !hmaster3_p & v3a70ffe;
assign v373698b = hbusreq6 & v3a6f03f | !hbusreq6 & v3a70a7f;
assign v37553f5 = hbusreq5 & v3a6087b | !hbusreq5 & v3757ad8;
assign v374478a = hbusreq7_p & v37290fa | !hbusreq7_p & !v2acb094;
assign v372bc6c = hmaster0_p & v37447f7 | !hmaster0_p & v375c65a;
assign v3a6837d = hbusreq6_p & v374faa9 | !hbusreq6_p & v37789da;
assign v3a71644 = hgrant0_p & v8455ab | !hgrant0_p & !v3744b38;
assign v37519bf = hbusreq5_p & v3765c1f | !hbusreq5_p & v37623f5;
assign v373aa77 = hlock0_p & v375098f | !hlock0_p & v3762244;
assign v38097fc = hlock1_p & v3a6fc65 | !hlock1_p & !v8455ab;
assign v375e1a2 = hbusreq2_p & v377bc89 | !hbusreq2_p & v3a6feb9;
assign v373f88a = hlock5_p & v3735930 | !hlock5_p & v8455e7;
assign v376780f = hlock6 & v3731c1c | !hlock6 & v374bc3e;
assign v376aa76 = hbusreq0 & v3a715a9 | !hbusreq0 & v37629bf;
assign v3a70fa2 = hbusreq3 & v374cab9 | !hbusreq3 & !v8455ab;
assign v3378fb8 = hbusreq3_p & v3759f4c | !hbusreq3_p & v8455b0;
assign v20930c6 = hgrant4_p & v3774bad | !hgrant4_p & v37368e1;
assign v374d617 = hmaster1_p & v3a635ea | !hmaster1_p & v3a70582;
assign v372cace = hmaster1_p & v3a57ce9 | !hmaster1_p & v373823e;
assign v3741fc9 = hbusreq0 & v372a79f | !hbusreq0 & v3735fdc;
assign v3778b19 = hgrant4_p & v3a70969 | !hgrant4_p & v3728127;
assign v3779a9c = hbusreq5 & v37565a6 | !hbusreq5 & v375ee2e;
assign v3779be2 = hmaster2_p & v3a637dd | !hmaster2_p & v3770ccf;
assign v377a8ea = hmaster2_p & v3a7002c | !hmaster2_p & v376158d;
assign v3a6f947 = hbusreq2 & v377cd7a | !hbusreq2 & v375c1d1;
assign v37567ef = hbusreq5 & v37301dd | !hbusreq5 & v3a705e4;
assign v372de52 = stateG10_1_p & v8455ab | !stateG10_1_p & v3743aee;
assign v374a8db = hmaster2_p & v3a635ea | !hmaster2_p & v3756304;
assign v372acd0 = hmaster2_p & v3753a06 | !hmaster2_p & v8455ab;
assign v3778fae = hbusreq8_p & v373bfd8 | !hbusreq8_p & v373c7af;
assign v37366eb = hmaster1_p & v372b9c5 | !hmaster1_p & v373e674;
assign v3724600 = hmaster1_p & v37645bc | !hmaster1_p & v3a68821;
assign v3a70734 = hgrant2_p & v377a291 | !hgrant2_p & v8455ab;
assign v3750b9b = hlock7_p & v3743d03 | !hlock7_p & v3744410;
assign v3a548f2 = hgrant2_p & v3a709df | !hgrant2_p & v3a6145f;
assign v3a64a14 = hbusreq5 & v38072a2 | !hbusreq5 & v3a54466;
assign v3a70cd2 = hbusreq0_p & v3806507 | !hbusreq0_p & v3a63621;
assign v374061b = hbusreq6_p & v3a57660 | !hbusreq6_p & v8455ab;
assign v3a5a374 = stateG10_1_p & v8455ab | !stateG10_1_p & !v3a703ca;
assign v3731c72 = hlock6_p & v375ed9f | !hlock6_p & v375e9a7;
assign v37258b7 = hgrant4_p & v375c170 | !hgrant4_p & v3a5f5e8;
assign v3a5d4d0 = hgrant4_p & v8455c1 | !hgrant4_p & v372451b;
assign v1e37759 = hbusreq8 & v3a6ffd7 | !hbusreq8 & v37565d3;
assign v376fe6e = hgrant4_p & v3753429 | !hgrant4_p & v3a6fdcc;
assign v3759d98 = jx1_p & v377e04a | !jx1_p & v3730d52;
assign v3776fb8 = hmaster2_p & v3a6f213 | !hmaster2_p & v35b774b;
assign v3a5ba58 = hbusreq5 & v37689be | !hbusreq5 & v3a71658;
assign v3a71630 = hbusreq3 & v3a58218 | !hbusreq3 & v8455ab;
assign v2092ee9 = hmaster1_p & v3a587be | !hmaster1_p & v376314e;
assign v3738f04 = hbusreq1_p & v3a6f316 | !hbusreq1_p & v8455ab;
assign v377eb8b = hbusreq5 & v3729708 | !hbusreq5 & v3742bc3;
assign v3735f9a = hbusreq5 & v3762b52 | !hbusreq5 & v8455ab;
assign v3a5f41b = hbusreq4_p & v8455ab | !hbusreq4_p & v375dab2;
assign v374c718 = hgrant3_p & v3a5e1a5 | !hgrant3_p & v3a6f7f0;
assign v37261be = hmaster2_p & v3756f10 | !hmaster2_p & !v373d2bd;
assign v39eb44e = hmaster1_p & v3a715bb | !hmaster1_p & v37490ae;
assign v1e37b5a = hmaster2_p & v374e855 | !hmaster2_p & v3763295;
assign v372fbf8 = hbusreq2 & v3729421 | !hbusreq2 & v8455bd;
assign v3731079 = hmaster2_p & v3a6d806 | !hmaster2_p & v374394c;
assign v374ba05 = hbusreq0 & v3a7136a | !hbusreq0 & v374e6e3;
assign v3767b6e = hbusreq4_p & v3a700ec | !hbusreq4_p & v3757684;
assign v3778fb5 = hlock5 & v3a56789 | !hlock5 & v3a70f62;
assign v3a6f31f = hmaster2_p & v8455ca | !hmaster2_p & v8455ba;
assign v3725947 = hbusreq6 & v3725230 | !hbusreq6 & v8455ab;
assign v3754c2d = hgrant0_p & v3a71647 | !hgrant0_p & v3762bf1;
assign v3756740 = hlock5_p & v377246b | !hlock5_p & !v3807b2e;
assign v373a7d4 = hmastlock_p & v3a6446a | !hmastlock_p & v8455ab;
assign v374a35d = hmaster1_p & v3a68cb5 | !hmaster1_p & !v375eb79;
assign v372d2cd = hgrant5_p & v3a6eca6 | !hgrant5_p & v3743057;
assign v373f7b7 = hbusreq6 & v377b84e | !hbusreq6 & v38072fd;
assign v377a4f1 = hbusreq3 & v3a6fe46 | !hbusreq3 & v8455ab;
assign v3a6cf91 = hmaster1_p & v3a7060c | !hmaster1_p & v372c92c;
assign v373aaca = stateG3_1_p & v845601 | !stateG3_1_p & !v8455ab;
assign v37629bf = hlock0 & v3765e79 | !hlock0 & v3a715a9;
assign v3750866 = hlock3 & v377b292 | !hlock3 & v3a70321;
assign v37603a3 = hbusreq2_p & v3a5d555 | !hbusreq2_p & !v377408e;
assign v3a711da = hbusreq6_p & v3a55349 | !hbusreq6_p & v372bbb3;
assign v3752446 = hbusreq6_p & v374ad96 | !hbusreq6_p & !v8455ab;
assign v3749762 = hmaster3_p & v3a6eaf6 | !hmaster3_p & v377abbe;
assign v3a70626 = hbusreq3_p & v3a6ac26 | !hbusreq3_p & v3732d4b;
assign v376f51a = hgrant5_p & v3725576 | !hgrant5_p & v377fc89;
assign v37588a3 = hbusreq4_p & v375624e | !hbusreq4_p & v373b610;
assign v3a5b571 = hbusreq5 & v3752d24 | !hbusreq5 & v3a55c8f;
assign v3761930 = hmaster3_p & v3a5a52f | !hmaster3_p & v3a70931;
assign v3a6b560 = hbusreq3_p & v376d34b | !hbusreq3_p & v3748797;
assign v3751bf3 = hbusreq8 & v37479c3 | !hbusreq8 & v372b396;
assign v3a682cb = hlock3_p & v3a5b5d3 | !hlock3_p & v3a658bf;
assign v375937f = hbusreq6 & v37251e7 | !hbusreq6 & v376ef7a;
assign v3730693 = hbusreq3_p & v375d7b6 | !hbusreq3_p & v377d34b;
assign v3a6b2c9 = hbusreq4_p & v374165a | !hbusreq4_p & v8455ab;
assign v2ff8e61 = hbusreq8_p & v3726638 | !hbusreq8_p & !v3a698e1;
assign v37395d4 = hmaster1_p & v3a70ca8 | !hmaster1_p & v3a70a25;
assign v376d76c = hmaster0_p & v3a70b7d | !hmaster0_p & v3a6d367;
assign v372c470 = hgrant5_p & v8455ab | !hgrant5_p & d4044f;
assign v3729f6c = hbusreq4_p & v372d9ad | !hbusreq4_p & v3a5c59f;
assign v373c755 = locked_p & v37656ec | !locked_p & v8455ab;
assign v8e42b4 = hbusreq5_p & v3a7156e | !hbusreq5_p & v376e7cf;
assign v377c174 = hmaster0_p & v3768fc7 | !hmaster0_p & v8455ab;
assign v374eb3b = hmaster1_p & v3771a62 | !hmaster1_p & v3755502;
assign v39eaa47 = hbusreq1_p & b4fa3c | !hbusreq1_p & v3763498;
assign v3755f9d = hmaster0_p & v37516ba | !hmaster0_p & v8455ab;
assign v3a649da = jx0_p & v373b6dd | !jx0_p & v3727a6b;
assign v376725a = hbusreq2 & v3a6528b | !hbusreq2 & v8455ab;
assign v377d74c = hgrant4_p & v3754df4 | !hgrant4_p & v3a296e8;
assign v3727a2b = hbusreq8_p & v376bb81 | !hbusreq8_p & v372deb9;
assign v3752aa5 = hbusreq6_p & v3a6eae6 | !hbusreq6_p & v3a71395;
assign v375d2b3 = hmaster2_p & v3747ac9 | !hmaster2_p & v3a5a0d2;
assign v3777a8c = hgrant6_p & v375f3e2 | !hgrant6_p & v372b512;
assign v374056e = hgrant3_p & v3a5872a | !hgrant3_p & v2acaf23;
assign v3a70f27 = hlock5 & v376a47e | !hlock5 & v3a70d21;
assign v3a70941 = hmaster2_p & v3769d48 | !hmaster2_p & v375e721;
assign v373e07e = hmaster1_p & v3a635ea | !hmaster1_p & v3a61c80;
assign v376a0e6 = hbusreq7_p & v377de4d | !hbusreq7_p & !v37738b2;
assign v37522ea = hlock4 & v3a7019a | !hlock4 & v375cf55;
assign v3a706ba = hbusreq8_p & v3737456 | !hbusreq8_p & v3a691ca;
assign v3739ea3 = hbusreq0 & v3778648 | !hbusreq0 & v375c41e;
assign v377eea3 = hmaster2_p & v3774a95 | !hmaster2_p & v3a5bfc8;
assign v372919e = hbusreq7_p & v3736dfd | !hbusreq7_p & v3725688;
assign v3769cad = hburst1 & v39ebac7 | !hburst1 & v3a709c6;
assign v3722f60 = hmaster1_p & v3a68426 | !hmaster1_p & v3a6b4a2;
assign v3a6fb43 = hbusreq5 & v3773078 | !hbusreq5 & v3a705d4;
assign v377f113 = hmaster0_p & v37419ca | !hmaster0_p & v37445ff;
assign v3a70f2a = hgrant7_p & v8455ab | !hgrant7_p & !v8455f3;
assign v376b706 = hgrant7_p & v3a6e708 | !hgrant7_p & v373ac95;
assign v3741ab9 = hmaster0_p & v3a6fe5c | !hmaster0_p & v3a580fb;
assign v3734473 = hbusreq7_p & v8455ab | !hbusreq7_p & v376d432;
assign v3770def = hbusreq5 & v3763076 | !hbusreq5 & v3a6ff12;
assign v3772a4f = hmaster1_p & v3a66d94 | !hmaster1_p & v3768c08;
assign v37c0382 = hbusreq1_p & v9230c3 | !hbusreq1_p & !v8455ab;
assign v9da9d2 = hbusreq2_p & v3736ebd | !hbusreq2_p & v3a6cb69;
assign v3a6f389 = hmaster1_p & v3a6b924 | !hmaster1_p & v3743e4f;
assign v3a6de90 = hbusreq2_p & v3769ae2 | !hbusreq2_p & v3772698;
assign v37590a2 = hbusreq0 & v37510e0 | !hbusreq0 & v373a9ee;
assign v377851b = hmaster2_p & v3a60787 | !hmaster2_p & v3a6a213;
assign v3741365 = hmaster2_p & v3a6e7b3 | !hmaster2_p & v2925c39;
assign v3a5fb9e = hbusreq5 & v3a6ff39 | !hbusreq5 & v372c433;
assign v3770548 = hgrant1_p & v3755791 | !hgrant1_p & v8455ab;
assign v376c2e6 = hmaster0_p & v37636e3 | !hmaster0_p & b05db7;
assign v3a296e8 = hbusreq0 & v3767385 | !hbusreq0 & v37664a1;
assign v373c111 = hbusreq4_p & v3a63559 | !hbusreq4_p & v3a6157d;
assign v3a6fb37 = hmaster2_p & v3a5f6d5 | !hmaster2_p & v3a64ded;
assign v3772020 = hgrant3_p & v373e37c | !hgrant3_p & v37707eb;
assign v3a706d3 = hmaster2_p & v3a63e82 | !hmaster2_p & v3761ad8;
assign v37605bb = hbusreq3 & v3a6edab | !hbusreq3 & v376bade;
assign v3a614dd = jx0_p & v372c79f | !jx0_p & v374e455;
assign v3767561 = hlock2_p & v3379037 | !hlock2_p & !v8455ab;
assign v377c4bd = hgrant0_p & c7f8d6 | !hgrant0_p & !v3767527;
assign v3a7056c = hbusreq4 & v3727713 | !hbusreq4 & v3a57959;
assign v3756a04 = hmaster2_p & v376e72d | !hmaster2_p & v3a58057;
assign v375c6d6 = hready_p & v23fda46 | !hready_p & v37587a6;
assign v373b4ad = hgrant3_p & v377eaf2 | !hgrant3_p & v8455ab;
assign v373dd3c = hlock5_p & v373a2f4 | !hlock5_p & v3a5b25f;
assign v37686f3 = hbusreq0 & v375a771 | !hbusreq0 & v3a6504e;
assign v376a056 = hbusreq6_p & v3724db7 | !hbusreq6_p & v8455ab;
assign v3a71388 = hmaster2_p & v374e28f | !hmaster2_p & !v3759379;
assign v3a58cf7 = hbusreq6 & v3806c41 | !hbusreq6 & v3a5b6de;
assign v3755aef = hgrant3_p & v3758c35 | !hgrant3_p & v376bb64;
assign v3756a59 = hmaster0_p & v374e855 | !hmaster0_p & v1e37b5a;
assign v3a2981d = hbusreq7_p & v377dfbd | !hbusreq7_p & v3a612df;
assign v3751090 = hbusreq4 & v1e37b3f | !hbusreq4 & v372b5a3;
assign v92141c = hgrant2_p & v8455ba | !hgrant2_p & v373e0ad;
assign v373ed95 = hbusreq2_p & v3745149 | !hbusreq2_p & v3a712e3;
assign v377ecf0 = hmaster2_p & v3a70641 | !hmaster2_p & v3a660f2;
assign v375cddb = hmaster2_p & v3747302 | !hmaster2_p & v374acbe;
assign v3a70727 = hmaster1_p & v3a61a7f | !hmaster1_p & v374fa11;
assign v3727b0e = hgrant4_p & v377ccba | !hgrant4_p & v3a7094d;
assign v3749d58 = hgrant2_p & v3775b81 | !hgrant2_p & v8455ab;
assign v3a60576 = hbusreq6_p & v374eb6a | !hbusreq6_p & !v3a7151d;
assign v3726434 = hmaster2_p & v3751c4c | !hmaster2_p & v372aacd;
assign v3a6c0ba = hmaster0_p & v3a61f4c | !hmaster0_p & v374ad7d;
assign v3a6fdd8 = hbusreq6 & v3768ecc | !hbusreq6 & v8455e7;
assign v3776c09 = hlock0_p & v3760e7b | !hlock0_p & v375a7fc;
assign v3a70762 = hgrant8_p & v8455ab | !hgrant8_p & v3749a98;
assign v3728957 = hbusreq0 & v3a70353 | !hbusreq0 & v3a70e9b;
assign v3a6fd50 = hgrant2_p & v3747c3e | !hgrant2_p & v8455ab;
assign v376d810 = hbusreq8_p & v373d4f7 | !hbusreq8_p & v377c831;
assign v373de53 = hgrant6_p & v377bd79 | !hgrant6_p & v3a5a34e;
assign v3768c5d = hbusreq4_p & v3a64722 | !hbusreq4_p & v372a823;
assign v3762121 = hbusreq8 & v360d029 | !hbusreq8 & !v8455ab;
assign v375cec6 = hgrant1_p & v3a619c0 | !hgrant1_p & v376ba47;
assign v3751c4b = hbusreq2 & v373c01b | !hbusreq2 & v3a5b6de;
assign v376285a = hburst1 & v3771ce2 | !hburst1 & v2ff8c78;
assign v3985143 = decide_p & v373fc77 | !decide_p & v3a70772;
assign v3a5e541 = hbusreq5 & v3746061 | !hbusreq5 & v3a5923e;
assign v3772513 = hgrant6_p & v375d288 | !hgrant6_p & v3a5f315;
assign v37508a4 = hgrant0_p & v3a6faac | !hgrant0_p & v3a5ef59;
assign v3a70a37 = hmaster0_p & v3768421 | !hmaster0_p & v376db34;
assign v1e379c4 = hmaster0_p & v374e6c7 | !hmaster0_p & v3727e58;
assign v373501a = hbusreq8 & v3a6f0ca | !hbusreq8 & v8455ab;
assign v8f559e = hlock6 & v373fe7b | !hlock6 & v376d081;
assign v3a6fd57 = hbusreq1_p & v376f152 | !hbusreq1_p & v372f22b;
assign v3a58ba8 = hlock6 & v3a70bff | !hlock6 & v372cb77;
assign v37409f4 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v3a5dd17;
assign v3a69a9f = hmaster0_p & v3a6a8c0 | !hmaster0_p & a1bc5b;
assign v377cd68 = hmaster1_p & v3a5c3d6 | !hmaster1_p & v35b91b9;
assign v3a572e2 = hbusreq7 & v3a567ea | !hbusreq7 & v375538e;
assign v3a68bf8 = hlock3 & v3a6fc64 | !hlock3 & v3759b7c;
assign v377e2ae = hbusreq4 & v3754422 | !hbusreq4 & v38072fd;
assign v360d1cd = hmaster2_p & v3a57f59 | !hmaster2_p & !v3735e39;
assign v3a6bf41 = hgrant6_p & v8455ab | !hgrant6_p & v391331d;
assign v3768b81 = hgrant0_p & v373ca4f | !hgrant0_p & !v8455ab;
assign v3772e44 = hbusreq7 & v37690e7 | !hbusreq7 & v3a70242;
assign v375fd29 = hgrant4_p & v8455ab | !hgrant4_p & v1e37762;
assign v375d8e0 = hlock6 & v374ba04 | !hlock6 & v377d41d;
assign v3a70122 = jx0_p & v3779d24 | !jx0_p & v360caba;
assign v3739f07 = hbusreq6_p & v3a6f238 | !hbusreq6_p & v377d310;
assign v37408b7 = hlock7 & v373280e | !hlock7 & v3a58673;
assign v3727369 = hbusreq6 & v3733471 | !hbusreq6 & v8455ab;
assign v3732c6a = hbusreq5 & v8455b0 | !hbusreq5 & v373eadd;
assign v3a6f2fc = hbusreq5 & v37356f0 | !hbusreq5 & v8455ab;
assign v374383b = hbusreq3_p & v374f20c | !hbusreq3_p & v3a60132;
assign v3a5a711 = jx2_p & v373c164 | !jx2_p & v3a57887;
assign v3a65dc4 = hgrant2_p & v8455ba | !hgrant2_p & v374b918;
assign v377a5a9 = hlock6 & v375a41b | !hlock6 & v3a60008;
assign v377e85a = hbusreq4 & v3a53d12 | !hbusreq4 & v377b946;
assign v3a708a8 = hlock2 & v372ee70 | !hlock2 & v3a61f82;
assign a792d5 = hmaster1_p & v3a67269 | !hmaster1_p & v3a66a3a;
assign v3741d99 = hbusreq6 & v374e9ac | !hbusreq6 & v37542af;
assign v2678c95 = hgrant6_p & v3a69146 | !hgrant6_p & v3723555;
assign v3a7136e = hbusreq0 & v37790ef | !hbusreq0 & v8455ab;
assign v3a71687 = hbusreq5 & v3724c63 | !hbusreq5 & v3753f1d;
assign v3771804 = hbusreq8 & v377a01a | !hbusreq8 & !v3808d0f;
assign v3a56d30 = hmaster0_p & v3a58cfc | !hmaster0_p & v373cd8f;
assign c2e325 = hlock5_p & v376c4ba | !hlock5_p & v375b2af;
assign v377b423 = hbusreq4_p & v37367a0 | !hbusreq4_p & v3761ca9;
assign v8fdd0d = hmaster1_p & v8455e7 | !hmaster1_p & v373759d;
assign v3a702e8 = hbusreq4 & v360d147 | !hbusreq4 & v8455ab;
assign v3735f51 = hmaster0_p & v373632a | !hmaster0_p & v3754727;
assign d03e23 = hmaster3_p & v377e9c1 | !hmaster3_p & !v3a681f5;
assign v3767e7e = hbusreq0 & v3a6e5f0 | !hbusreq0 & v377ce1a;
assign v37343f6 = hlock8 & v3737265 | !hlock8 & v374ffb8;
assign v3a6a66f = hgrant6_p & v8455ab | !hgrant6_p & v3a6e8a4;
assign v3773091 = hgrant1_p & v374306c | !hgrant1_p & v3a57330;
assign v374f7cb = hmaster0_p & v3a7106b | !hmaster0_p & v3742bc1;
assign v37705be = hmaster3_p & v8455ab | !hmaster3_p & v3a6a720;
assign v3745b20 = hlock6 & v3a6f338 | !hlock6 & v35b779f;
assign v3752cc5 = hgrant4_p & v3a53eeb | !hgrant4_p & v3a6fac6;
assign v376d81c = hmaster2_p & v3a637dd | !hmaster2_p & !v377c44f;
assign v37332af = hmaster2_p & v3774bad | !hmaster2_p & v3a5d5a4;
assign v373b241 = hlock8 & v376ae9f | !hlock8 & v3739c89;
assign v374fa0d = hgrant2_p & v8455ab | !hgrant2_p & v3a63dcc;
assign v3a6f07d = hgrant4_p & v3a6ef0e | !hgrant4_p & v3577421;
assign v3728230 = hgrant4_p & v372b77b | !hgrant4_p & v375ed63;
assign v3739594 = hbusreq4 & v37770c9 | !hbusreq4 & v8455ab;
assign v3741d00 = stateG10_1_p & d8a75b | !stateG10_1_p & v3732817;
assign v3a6a63c = hmaster2_p & v8455ab | !hmaster2_p & !v3a62abc;
assign v377a8e0 = hlock4 & v374e3a9 | !hlock4 & v3a6f8d5;
assign v374f871 = hlock2_p & v376223b | !hlock2_p & v8455b0;
assign v3757f54 = hmaster2_p & v373cf9c | !hmaster2_p & v37786a6;
assign v3378fca = hbusreq3 & v3806db7 | !hbusreq3 & v372fba5;
assign v3770719 = hbusreq0 & v3778a76 | !hbusreq0 & v377d042;
assign v373c1a0 = hmaster2_p & v3a5e696 | !hmaster2_p & !v8455ab;
assign v3a57c0d = hbusreq5 & v372c85f | !hbusreq5 & v3a6d0af;
assign v3729fa4 = hlock5_p & v374dfe1 | !hlock5_p & v3770367;
assign v3743dbc = hbusreq3_p & v372b765 | !hbusreq3_p & !v3a5cd20;
assign v3764e37 = hmaster2_p & v8455ab | !hmaster2_p & v3a6f9f9;
assign v3a5d8b5 = hmaster2_p & v373f058 | !hmaster2_p & v3776685;
assign v374c9cf = hbusreq6 & v372fc81 | !hbusreq6 & !v8455ab;
assign v3a6ffda = hgrant6_p & v8455ca | !hgrant6_p & v3a6e0f2;
assign v3766658 = hmaster2_p & v374314f | !hmaster2_p & v8455ab;
assign v3a64b83 = hbusreq4 & v3760a55 | !hbusreq4 & v3a65d01;
assign v3748f09 = hbusreq4_p & v8cb684 | !hbusreq4_p & v8455b0;
assign v3a58038 = hlock4 & v3737681 | !hlock4 & v377221f;
assign v373e72e = hmaster0_p & v3a6c4e4 | !hmaster0_p & v3733de8;
assign v37563fe = hgrant3_p & v2acb088 | !hgrant3_p & !v3a6acab;
assign v376865d = hgrant2_p & v3732d55 | !hgrant2_p & v372b5a8;
assign v3752fe6 = hbusreq2_p & v35b71ca | !hbusreq2_p & v8455ab;
assign v3a70316 = hlock1_p & v37585a0 | !hlock1_p & v8455b0;
assign v37769ee = hbusreq1_p & v3a635ea | !hbusreq1_p & !v3728b9d;
assign v3741320 = hmaster2_p & v372310e | !hmaster2_p & v28896da;
assign v3a6f6e8 = hbusreq7 & v3762ac3 | !hbusreq7 & v376a06d;
assign v375b26a = hbusreq4 & v3a6ff74 | !hbusreq4 & v3763104;
assign v374fac9 = hmaster0_p & v3a64854 | !hmaster0_p & v376ebc6;
assign v3807072 = hbusreq7 & v3776be5 | !hbusreq7 & v3736ded;
assign v3730d1e = hmaster2_p & v375d9b1 | !hmaster2_p & !v37389d5;
assign v3a6deea = hlock5 & v3a5d405 | !hlock5 & v377653f;
assign v375d3bb = hmaster1_p & v3748ac8 | !hmaster1_p & v3a58803;
assign v372b69c = jx3_p & v374f2d1 | !jx3_p & v3a62dec;
assign v3a5c210 = hgrant2_p & v3768b99 | !hgrant2_p & !v3a6f4f4;
assign v3736cb8 = hbusreq4 & v3753bb2 | !hbusreq4 & v3a67cff;
assign v3a5d94f = jx0_p & v376bce3 | !jx0_p & v37242f1;
assign v377395b = hbusreq2 & a29a96 | !hbusreq2 & v8455ab;
assign v3a56a86 = hbusreq5 & v3768495 | !hbusreq5 & v3a55cda;
assign v3a5ec91 = hgrant6_p & v3729214 | !hgrant6_p & v374b2f7;
assign v372a56e = hbusreq7_p & v3a70deb | !hbusreq7_p & v3a706c8;
assign v375f0f8 = hmaster0_p & v377766c | !hmaster0_p & v375754a;
assign v3a5b909 = hlock1 & v380693e | !hlock1 & v373f19e;
assign v3737ceb = hlock5 & v3a63f9a | !hlock5 & v3a5cb0e;
assign v375adcd = hmaster1_p & v377b774 | !hmaster1_p & v377b4bf;
assign v3736b4a = hbusreq5 & v376b38c | !hbusreq5 & v375517b;
assign v374cd10 = hbusreq6 & v3727615 | !hbusreq6 & v375de7f;
assign v3760ce0 = jx2_p & v3a6b368 | !jx2_p & v3767010;
assign v376dcbe = hmaster2_p & v376c7d1 | !hmaster2_p & v376358f;
assign v3a6f0d1 = hbusreq3_p & v3725ba8 | !hbusreq3_p & v3a6c55a;
assign v3771ddb = hgrant4_p & v372b77b | !hgrant4_p & v375da9d;
assign v3a6fa76 = hbusreq6 & v3809de2 | !hbusreq6 & v38072fd;
assign v373c071 = hmaster3_p & v376ac47 | !hmaster3_p & v3a6c6c3;
assign v3740655 = hbusreq3 & v3a6fe0d | !hbusreq3 & !v8455b5;
assign v376d328 = hgrant2_p & v376b5f8 | !hgrant2_p & v3a7091c;
assign v3a5b3d8 = hbusreq6_p & v8455ab | !hbusreq6_p & v376e4da;
assign v3a70f15 = hbusreq8 & v8455e7 | !hbusreq8 & v3a64288;
assign v3a61dca = hmaster2_p & v376999f | !hmaster2_p & v372433d;
assign v3761a96 = hbusreq4 & v38097ca | !hbusreq4 & v3a70c74;
assign v3746ffa = hgrant6_p & v3a70b17 | !hgrant6_p & v3741dab;
assign v374b68a = hmaster2_p & v376f4b2 | !hmaster2_p & v3769ad7;
assign v372d842 = hmaster2_p & v8455c3 | !hmaster2_p & a34d2b;
assign v372879a = hlock6 & v3a5ef6e | !hlock6 & v37745b8;
assign v375e035 = hmaster1_p & v3a63777 | !hmaster1_p & v37476c2;
assign b21e3c = hbusreq4 & v3723635 | !hbusreq4 & v373bd6c;
assign v3a6f7d2 = hmaster1_p & v3745181 | !hmaster1_p & v3a6f838;
assign v3a6f959 = hmaster2_p & v3a635ea | !hmaster2_p & v375bb51;
assign v1e38288 = hgrant6_p & v37658d7 | !hgrant6_p & v3a70dde;
assign v3725470 = hbusreq8 & v375facf | !hbusreq8 & v3a60bae;
assign v3735db2 = hlock5 & v3775526 | !hlock5 & v3806def;
assign v3763d2c = hmaster1_p & v3779ff0 | !hmaster1_p & v37402ee;
assign v3762873 = hbusreq5 & v3747a68 | !hbusreq5 & v3770a3b;
assign v3a6268c = hlock4_p & v3723eef | !hlock4_p & v8455b0;
assign v9d7045 = hmaster2_p & v39ea76e | !hmaster2_p & v3733e9e;
assign v3765a98 = hlock0_p & v3a706d1 | !hlock0_p & v8455b7;
assign v3723780 = hgrant5_p & v3a70e38 | !hgrant5_p & v375a79d;
assign v2acb006 = hmaster0_p & v3743966 | !hmaster0_p & v3a6230b;
assign v375b5ca = hmaster2_p & v3760353 | !hmaster2_p & v8455ab;
assign v37350f9 = hgrant4_p & v3a5f162 | !hgrant4_p & v3a712fd;
assign v3a62539 = hbusreq6_p & v375e948 | !hbusreq6_p & v37391b4;
assign bd3d3d = hbusreq2 & v8455bf | !hbusreq2 & !v374b25d;
assign v3761c1a = hmaster2_p & v3770f96 | !hmaster2_p & v37784b9;
assign v3766df8 = hmaster2_p & v3a5fabd | !hmaster2_p & v35772a6;
assign v37431ac = hmaster1_p & v3a61a7f | !hmaster1_p & v3a5c3ef;
assign v3736382 = hbusreq7_p & v3749975 | !hbusreq7_p & !v373b938;
assign v3a714aa = hgrant4_p & v3744417 | !hgrant4_p & v3a70cc0;
assign v3a5ccfd = hgrant3_p & v8455b5 | !hgrant3_p & v374a7cd;
assign v3a61668 = hbusreq3 & v3736e1d | !hbusreq3 & v3748797;
assign v3730e2e = hbusreq2_p & v3a708fa | !hbusreq2_p & v373f91b;
assign v3a70d05 = hbusreq3_p & v3771e18 | !hbusreq3_p & v8455ab;
assign v373ff9a = hmaster1_p & v3748656 | !hmaster1_p & v3774c55;
assign v3766709 = hgrant3_p & v3a57f59 | !hgrant3_p & v374dfd9;
assign v3746877 = hbusreq7 & v3a5bc72 | !hbusreq7 & v372721d;
assign v3771171 = hbusreq5 & v3770bcd | !hbusreq5 & v3a6eb3d;
assign v3765b5c = hmaster1_p & v37386c6 | !hmaster1_p & v2ff8f33;
assign v97c94a = hbusreq7_p & v3a54cd9 | !hbusreq7_p & v373c7af;
assign v3760bd6 = hlock0_p & v3a5db8a | !hlock0_p & v8455ab;
assign v375bb26 = hmaster0_p & v3a6cc9a | !hmaster0_p & v373594b;
assign v3a6a6b4 = hbusreq6 & v3740194 | !hbusreq6 & v8455ab;
assign v3a6cac4 = jx0_p & v8455bd | !jx0_p & v8455ab;
assign v373c8a4 = jx0_p & v3a636c0 | !jx0_p & v3a61964;
assign v3a71545 = hmaster3_p & v3a68183 | !hmaster3_p & v3735350;
assign v3771720 = hgrant0_p & v8455ab | !hgrant0_p & !v372bdef;
assign v3a6f32a = stateG10_1_p & v1e38224 | !stateG10_1_p & v3770b89;
assign v3a6dc08 = hready & v376c9ee | !hready & !v8455ab;
assign v3a70b0e = hlock6 & v3a63e87 | !hlock6 & v3a5dbc7;
assign v373d8f2 = hlock4 & v3730451 | !hlock4 & v3740a38;
assign v374d41e = hlock8_p & v3a70f52 | !hlock8_p & v3760066;
assign v374d01c = hmaster0_p & v3a6efe8 | !hmaster0_p & v372f173;
assign v3743dce = hmaster1_p & v3a635ea | !hmaster1_p & v3769639;
assign v372992f = hlock6_p & v373f028 | !hlock6_p & v3a5b4c1;
assign v3742723 = hlock4 & v374e353 | !hlock4 & v373340d;
assign v3776592 = hbusreq6 & v3a6fcb9 | !hbusreq6 & v8455ab;
assign v3a703ca = hgrant1_p & v3a653e4 | !hgrant1_p & v3a637dd;
assign v3776eef = hmaster1_p & v3734967 | !hmaster1_p & v373c642;
assign v3750f3b = hbusreq8_p & v3762cdf | !hbusreq8_p & v3a70c78;
assign v3a70ce5 = hmaster0_p & v3a5e7dc | !hmaster0_p & !v374da92;
assign v374fa11 = hlock5 & v3a70586 | !hlock5 & v377a0d8;
assign v37256c4 = hgrant0_p & v3731678 | !hgrant0_p & v373eedf;
assign v377e11d = hlock0 & v3779cf9 | !hlock0 & v373059e;
assign v3a70538 = hmaster2_p & v2092faa | !hmaster2_p & v372493b;
assign v3a6046c = stateA1_p & v37295fe | !stateA1_p & v3a71085;
assign v3a673d6 = hlock6_p & v3724200 | !hlock6_p & v37531af;
assign v374457a = hmaster0_p & v375bce7 | !hmaster0_p & v3a70716;
assign v37607e8 = hbusreq2_p & v3757fcc | !hbusreq2_p & v3763acf;
assign v3748460 = hmaster0_p & v3745cc6 | !hmaster0_p & v3a7060a;
assign v3a6f86b = hmaster0_p & v3a6a312 | !hmaster0_p & v379318b;
assign v23fd9f9 = hmaster2_p & v3a635ea | !hmaster2_p & v3a5af28;
assign v372d943 = hbusreq0_p & v3759032 | !hbusreq0_p & v3733e9e;
assign v3a6f47a = hmaster0_p & v377c5de | !hmaster0_p & v37328f1;
assign v376e3fb = hgrant4_p & v8455ab | !hgrant4_p & !v3a712b1;
assign v3a70a43 = hgrant2_p & v3a645ca | !hgrant2_p & v3a70e36;
assign v3745a0a = hbusreq2 & v3a5b037 | !hbusreq2 & v8455ab;
assign v3a5cd51 = hbusreq6_p & v3a5c945 | !hbusreq6_p & !v3a66110;
assign v3725882 = hmaster0_p & v377aefe | !hmaster0_p & v3a58b9f;
assign v3a582d6 = hlock2 & v3752fb7 | !hlock2 & v3a603bb;
assign v373b303 = hbusreq3 & v3a6fe90 | !hbusreq3 & !v8455ab;
assign v373f42d = hmaster2_p & v3757966 | !hmaster2_p & v3769cd7;
assign v374d14a = jx0_p & v3a5c46a | !jx0_p & v374f2fb;
assign c2b7ee = hbusreq5 & v37400ab | !hbusreq5 & v3809388;
assign v3a6f99e = hbusreq2_p & v375e657 | !hbusreq2_p & !v3a69591;
assign v377c9f3 = hbusreq7 & ca095d | !hbusreq7 & !v8455ca;
assign v3a7091e = hmaster1_p & v376b662 | !hmaster1_p & v373cbc5;
assign v377aede = hgrant2_p & v31c3694 | !hgrant2_p & v3a583dc;
assign v3a7025f = hlock2 & v3745039 | !hlock2 & v23fd923;
assign v372647d = hgrant4_p & v3a6ffea | !hgrant4_p & v374ad44;
assign v3732b63 = hmaster2_p & v3747c3e | !hmaster2_p & v8455ab;
assign c51aa0 = hbusreq6_p & v35b774b | !hbusreq6_p & v9ed516;
assign v37407ef = hbusreq7_p & v3734930 | !hbusreq7_p & v3753e74;
assign v37443a2 = hmaster0_p & v377adf5 | !hmaster0_p & v3a5e1e8;
assign v3a64dbb = hgrant5_p & d62aa6 | !hgrant5_p & v3a6f100;
assign v3758924 = hmaster1_p & v3729f64 | !hmaster1_p & v3a65388;
assign v3a70d4d = hmaster0_p & v8455b0 | !hmaster0_p & v376b870;
assign v3809ee4 = hbusreq4_p & v3a70641 | !hbusreq4_p & v3733383;
assign v376e979 = hbusreq5 & v3a6ed2b | !hbusreq5 & v3a705d4;
assign v3756ecd = hgrant4_p & v373fbb6 | !hgrant4_p & v3759de1;
assign v3a554f0 = hbusreq5 & v373b380 | !hbusreq5 & v377e018;
assign v3755207 = hbusreq5 & v3a6329a | !hbusreq5 & v375d417;
assign v3757dc4 = hlock5 & v3722b91 | !hlock5 & v3760644;
assign v3a6ac2e = hbusreq4 & v373b5d8 | !hbusreq4 & v8455ab;
assign v3a58ddb = hgrant4_p & v8455ab | !hgrant4_p & v3729bf3;
assign v374ae4e = jx0_p & v376702c | !jx0_p & v8455ab;
assign v3728f3a = hlock4 & v3763186 | !hlock4 & v3768870;
assign v374b8e2 = hgrant2_p & v376b307 | !hgrant2_p & v3a6b1e4;
assign v3a6811a = hmaster0_p & v373cd03 | !hmaster0_p & v3a5ac38;
assign v3a71560 = hmaster2_p & v3763f95 | !hmaster2_p & v3753dab;
assign v37686c2 = hlock4_p & v374d057 | !hlock4_p & v3a6fd81;
assign v372f2ff = hgrant5_p & v374407e | !hgrant5_p & d193f7;
assign v3a65053 = hbusreq4_p & v375f147 | !hbusreq4_p & v3a71503;
assign v3a6f750 = hmaster1_p & v3a635ea | !hmaster1_p & ca50c0;
assign v3725dc4 = hbusreq6 & v3a6dc08 | !hbusreq6 & adf78a;
assign v3740a94 = hgrant5_p & a80fe2 | !hgrant5_p & v372437d;
assign v3a6e975 = hbusreq5_p & v3a59cf3 | !hbusreq5_p & v8455ab;
assign v3732246 = hgrant6_p & v3743eae | !hgrant6_p & v3a68c1c;
assign v374d7a7 = hmaster1_p & v99797a | !hmaster1_p & v374ef4a;
assign v37758e6 = hbusreq7 & v3a6f292 | !hbusreq7 & v3729180;
assign v377d831 = jx0_p & v374f252 | !jx0_p & v3a6f931;
assign v375585a = hmaster0_p & v376da5f | !hmaster0_p & v3a7090f;
assign v373c5dc = hmaster2_p & v374729b | !hmaster2_p & !v372ee7e;
assign v37390c5 = hburst1 & v37295fe | !hburst1 & v3751807;
assign v3a70a54 = hmaster1_p & v8455ab | !hmaster1_p & !v3a6ebc5;
assign v373cb89 = hlock5 & v3774d6e | !hlock5 & v3770ad8;
assign v3742adb = hlock6_p & v373b3fb | !hlock6_p & v373006f;
assign v373c0a8 = hmaster3_p & v3a70ae5 | !hmaster3_p & v3a6843c;
assign v376a65b = hbusreq8 & v377cb85 | !hbusreq8 & v374c2aa;
assign v372ea5d = hbusreq5 & v372f0c7 | !hbusreq5 & v377dc82;
assign v377de57 = hbusreq5 & v373ad8b | !hbusreq5 & v8455ab;
assign v374190f = hmaster2_p & v3a70d99 | !hmaster2_p & v3775537;
assign v3741925 = hbusreq4_p & v377ba37 | !hbusreq4_p & !v8455ab;
assign v3a62589 = hlock6 & v376bb05 | !hlock6 & v376b4a8;
assign v374cbc3 = hbusreq5 & v3a6feb4 | !hbusreq5 & v8455ab;
assign v373dfec = hgrant4_p & v372dc51 | !hgrant4_p & v3745658;
assign v38098bf = hmaster0_p & v3a5af94 | !hmaster0_p & !v3730876;
assign v37798bb = hmaster1_p & v8455ab | !hmaster1_p & v377a91a;
assign v3a5e687 = hbusreq8_p & v373ca17 | !hbusreq8_p & v3a6299c;
assign v360d105 = hbusreq7 & v3772b81 | !hbusreq7 & v3a635ea;
assign v3749149 = hbusreq2_p & v8455bf | !hbusreq2_p & v377cd7a;
assign v3a63a7a = hbusreq0 & v377a42f | !hbusreq0 & v8455ab;
assign v3a6e231 = hbusreq7 & v3765203 | !hbusreq7 & v3723d79;
assign v376a08d = hbusreq2 & v3a6ab5f | !hbusreq2 & !v3a6ac2a;
assign v3737ce3 = hmaster0_p & v374b116 | !hmaster0_p & v375f014;
assign v377623c = hbusreq4 & v372ab46 | !hbusreq4 & v8455b3;
assign v37652f1 = hlock4 & v377af10 | !hlock4 & v3a67691;
assign v3772c5a = hmaster2_p & v3753dab | !hmaster2_p & v373ee80;
assign v3a6d1aa = hmaster2_p & v376f569 | !hmaster2_p & v3a7136e;
assign v3a71442 = hlock7_p & v3a68426 | !hlock7_p & v8455b7;
assign v3a6ebc9 = hbusreq5 & v37737aa | !hbusreq5 & v8455ab;
assign v3726806 = hlock0_p & v377395f | !hlock0_p & !v8455ab;
assign v380956e = hbusreq6_p & v3a6f61f | !hbusreq6_p & v377b860;
assign v376195f = hbusreq2 & v37251b9 | !hbusreq2 & v375da10;
assign v3a71350 = hlock3_p & v377d99d | !hlock3_p & !v8455ab;
assign v3a6fa18 = hmaster3_p & v38067ba | !hmaster3_p & v8455ab;
assign v3a60815 = hgrant5_p & v3a63cce | !hgrant5_p & v373024e;
assign v3a58d7a = hbusreq6 & v3739c76 | !hbusreq6 & v8455ab;
assign v372b5bc = hmaster0_p & v3732bff | !hmaster0_p & v3a71498;
assign v3766b27 = hgrant6_p & v3a69f9e | !hgrant6_p & v3a5988f;
assign v374fae5 = hbusreq2_p & v37765e1 | !hbusreq2_p & v373ed9a;
assign v37497d6 = hbusreq5_p & v37681a3 | !hbusreq5_p & v3a5f4c6;
assign v376ebbf = hbusreq6_p & v3a63eff | !hbusreq6_p & v373b288;
assign v373f247 = hbusreq5 & v3775adf | !hbusreq5 & bdb538;
assign v372c638 = hmaster2_p & v3724af9 | !hmaster2_p & v376856b;
assign v3a58541 = hbusreq7_p & v37c0282 | !hbusreq7_p & v3a66c14;
assign v372dd94 = hbusreq8 & v8455b0 | !hbusreq8 & v3735758;
assign v3754086 = hmaster1_p & v3a6fa3c | !hmaster1_p & v3728203;
assign v3770fdb = hbusreq5_p & v3777647 | !hbusreq5_p & v3a674fa;
assign v375d966 = hbusreq7 & v3a6f6f1 | !hbusreq7 & !v377a571;
assign v3778619 = hmaster0_p & v3727581 | !hmaster0_p & !v37c0294;
assign v3761912 = jx0_p & v8455ab | !jx0_p & v3767872;
assign v3a69ce6 = hlock8_p & v3772590 | !hlock8_p & v376945e;
assign v3757ab6 = hbusreq7 & v376cb10 | !hbusreq7 & v374e800;
assign v292500d = decide_p & v3a563aa | !decide_p & v3771fe5;
assign v376e16e = hgrant4_p & v8455ab | !hgrant4_p & v3a6bab9;
assign v3a6fe3f = hmaster2_p & v3775dbc | !hmaster2_p & v3728c23;
assign v375f798 = hbusreq7_p & v9a88fd | !hbusreq7_p & v3772214;
assign v37419e7 = hmaster2_p & v3a5ace5 | !hmaster2_p & v3a6febd;
assign v3752af0 = hbusreq2 & v3728e09 | !hbusreq2 & !v8455ab;
assign v376b8e9 = hgrant0_p & v8455ab | !hgrant0_p & v3a70fc0;
assign v39eb1df = hmaster2_p & v374502e | !hmaster2_p & !v3a7127f;
assign a1b632 = hmaster2_p & v375c675 | !hmaster2_p & v3a63a7a;
assign v37749fd = hgrant0_p & v8455ab | !hgrant0_p & v3a6dcb2;
assign v3770e95 = hbusreq0 & v23fe27f | !hbusreq0 & v373cdea;
assign v3a56866 = hbusreq3_p & v3760073 | !hbusreq3_p & v3a5cd20;
assign v3756524 = hgrant6_p & v8455ab | !hgrant6_p & !v3a7148c;
assign v373a902 = hmaster0_p & v8455ab | !hmaster0_p & v3765a79;
assign v377696a = hbusreq3 & v39a537f | !hbusreq3 & !v8455ab;
assign v3a70b9f = hbusreq5 & v374fde8 | !hbusreq5 & !v3754488;
assign v375911a = hbusreq3_p & v376d1e2 | !hbusreq3_p & v37348ee;
assign v3763b37 = hmaster0_p & v373e32c | !hmaster0_p & v3775100;
assign v374892a = hgrant4_p & v3777f86 | !hgrant4_p & v37681f3;
assign v3a5a057 = hgrant6_p & v3a6f2d4 | !hgrant6_p & v37627bf;
assign v3a57733 = hmaster1_p & v3a701de | !hmaster1_p & v3769948;
assign v3738e79 = hbusreq3 & v377ba55 | !hbusreq3 & v3724940;
assign v372300f = hgrant2_p & v8455ab | !hgrant2_p & v377ee33;
assign v37780e2 = hmaster0_p & v3731a49 | !hmaster0_p & v3a550cd;
assign v3776e85 = hgrant2_p & v8455ba | !hgrant2_p & v3a713e3;
assign v373d955 = hbusreq5 & v3a5e496 | !hbusreq5 & v3a5e4e5;
assign v374c9db = hbusreq2_p & v3a70aa2 | !hbusreq2_p & v2acae68;
assign v3732c95 = hmaster2_p & v3a70d45 | !hmaster2_p & v3a6f837;
assign v3a7042b = hready & v3752407 | !hready & v8455e7;
assign v3742b24 = hlock6 & v3a654af | !hlock6 & v376b7db;
assign v3a6f19b = hmaster1_p & v375620b | !hmaster1_p & v37695f7;
assign v3766dfb = hlock8 & v3a6ac9e | !hlock8 & v3a6faf0;
assign v3777bd6 = hbusreq6_p & v3a5dfad | !hbusreq6_p & v35772a6;
assign v376dcca = hbusreq4 & v3743c51 | !hbusreq4 & v375b349;
assign v3a61bfd = hgrant4_p & v3762924 | !hgrant4_p & !v3752e1b;
assign v372779c = hbusreq8_p & v3808c89 | !hbusreq8_p & v37475be;
assign v3a59424 = hbusreq6 & v3a70200 | !hbusreq6 & !v9edb6a;
assign v3a66fb0 = hbusreq8 & v3727195 | !hbusreq8 & v3736003;
assign v3a710c6 = hbusreq2_p & v37797a3 | !hbusreq2_p & v8455ab;
assign v3768768 = hgrant4_p & v37528fd | !hgrant4_p & v8455ab;
assign v37bfd10 = hlock6_p & v8455ab | !hlock6_p & v3a57ad0;
assign v3732775 = hmaster0_p & v3738c2e | !hmaster0_p & v3759bd0;
assign v374c5f6 = hbusreq8 & b9d061 | !hbusreq8 & v3a7016e;
assign v376e914 = locked_p & v3a63e82 | !locked_p & !v35772a6;
assign v3a5bc2c = hbusreq4_p & v8455bf | !hbusreq4_p & v3763a20;
assign v3734f60 = hbusreq7 & v3742e54 | !hbusreq7 & v8455ab;
assign v3a593bb = hgrant2_p & v3a5eadd | !hgrant2_p & v3a7133f;
assign v3755f80 = hgrant5_p & v3a70578 | !hgrant5_p & v375eb1b;
assign v374d674 = hbusreq6 & v372eaaf | !hbusreq6 & v377395f;
assign v37775c4 = hbusreq1_p & v1e37d3f | !hbusreq1_p & v3a70c07;
assign v3a6fd71 = hgrant1_p & v373a66d | !hgrant1_p & v3740171;
assign v3a6faab = jx0_p & v3a5c687 | !jx0_p & v3a6797d;
assign v3761065 = hmaster0_p & v3a6f9f7 | !hmaster0_p & v3744cd7;
assign v373f2e2 = hbusreq4 & v3a716a6 | !hbusreq4 & v8455ab;
assign v374e1c3 = hgrant4_p & v376b4ad | !hgrant4_p & b7df2b;
assign v372310e = hbusreq4_p & v3736ded | !hbusreq4_p & v377169f;
assign v372d3ea = hbusreq4_p & v3754b79 | !hbusreq4_p & v373ecd8;
assign v3732564 = hbusreq2_p & v3a7084e | !hbusreq2_p & !v8455ab;
assign v37647aa = hbusreq2 & v3763191 | !hbusreq2 & v35b774b;
assign v3747367 = hbusreq7_p & v3a5664b | !hbusreq7_p & v8455ab;
assign v375897d = hmaster0_p & v372e083 | !hmaster0_p & v3a71609;
assign v3a6e6c2 = hmaster2_p & v3a635ea | !hmaster2_p & v3a6f3c6;
assign v3778676 = hlock8 & v3a6f55c | !hlock8 & v3a6a0e4;
assign v37532c8 = hmaster2_p & v372ee0e | !hmaster2_p & !v8455ab;
assign v3734aef = hgrant6_p & v8455ab | !hgrant6_p & v3757b32;
assign ac4b49 = hbusreq8 & v37517f7 | !hbusreq8 & v375af91;
assign v3a649fd = hgrant6_p & v8455ab | !hgrant6_p & v3a62f13;
assign v3744f86 = hbusreq4 & v3730755 | !hbusreq4 & !v8455ab;
assign v3728382 = hlock8_p & v3a6d4cd | !hlock8_p & v8455ab;
assign v39ebb2e = hbusreq5 & v3a6fe41 | !hbusreq5 & v8455ab;
assign v3a708a4 = hbusreq0 & v374b274 | !hbusreq0 & v3762037;
assign v375c944 = hlock0 & v3a70b92 | !hlock0 & v2aca778;
assign v38097c0 = hmaster0_p & v372f885 | !hmaster0_p & v372e58c;
assign v3a57fb8 = hmaster2_p & v3736e7d | !hmaster2_p & v3a5a807;
assign v373e93e = hmaster0_p & v375a4eb | !hmaster0_p & v3a5e371;
assign v3a6f64a = hmaster2_p & v374f0c1 | !hmaster2_p & v35772a6;
assign v1e37e76 = hgrant0_p & v376a2ea | !hgrant0_p & v3758f3c;
assign v37c37ed = hbusreq7_p & v3a5dfa3 | !hbusreq7_p & v373cba8;
assign v37736b3 = hbusreq5 & v374b7e8 | !hbusreq5 & v3a5a219;
assign v37327ee = hbusreq4 & v37772db | !hbusreq4 & v37651c2;
assign a16ae7 = hlock6 & v38072fd | !hlock6 & v373f7b7;
assign v3a6b213 = jx0_p & a64c20 | !jx0_p & v373a782;
assign v3746efa = hbusreq5_p & v3766c68 | !hbusreq5_p & v3a60767;
assign v3a5a2a7 = hbusreq4 & v377961f | !hbusreq4 & v8455ab;
assign v3765960 = hbusreq5_p & v376f45b | !hbusreq5_p & v8455b7;
assign v3a6f1de = hbusreq1_p & v37284a9 | !hbusreq1_p & !v3a60584;
assign v375f2f3 = hmaster2_p & v8455e7 | !hmaster2_p & v3723b00;
assign v372c17e = hbusreq4 & v3723ace | !hbusreq4 & v8455ab;
assign v380877d = jx1_p & v375a0ed | !jx1_p & v37676e0;
assign v3741e9f = hgrant5_p & v3779a9a | !hgrant5_p & v3a6eb53;
assign v3729844 = hbusreq8_p & v3765a4a | !hbusreq8_p & v3a66c22;
assign v3a70c01 = hgrant3_p & v8455bd | !hgrant3_p & !v3743dbc;
assign v3742cfe = hbusreq2 & v3a712b6 | !hbusreq2 & v37730bf;
assign v3742655 = hbusreq2_p & v8455ab | !hbusreq2_p & v3a71061;
assign v3a64e3e = hbusreq5 & v3a6d2d7 | !hbusreq5 & v1e37405;
assign v372ae6a = hlock4_p & v3a7153a | !hlock4_p & v3a63805;
assign v3776f93 = hmaster1_p & v373173b | !hmaster1_p & v3a7121f;
assign v23fd869 = hbusreq7_p & v37386af | !hbusreq7_p & !v372bdb1;
assign v3a69bf4 = hbusreq3_p & v372ac83 | !hbusreq3_p & !v8455ab;
assign v373fa3d = hbusreq5_p & v3749ab1 | !hbusreq5_p & v372834d;
assign v3a5efc4 = hbusreq5_p & v375523d | !hbusreq5_p & v1e37579;
assign v3773a96 = hbusreq7 & v37655bf | !hbusreq7 & v374d6f6;
assign v23fe361 = hgrant4_p & v8455ab | !hgrant4_p & v3a6c2df;
assign v3a64624 = hlock5_p & v3a5a807 | !hlock5_p & !v373c050;
assign v373617a = hbusreq8_p & v3725948 | !hbusreq8_p & v3a62e3c;
assign v373a374 = hgrant0_p & v3733be0 | !hgrant0_p & v8455ab;
assign v37587a4 = hbusreq5_p & v38067ea | !hbusreq5_p & v3769740;
assign v3a6f4ca = hbusreq5 & v376cda5 | !hbusreq5 & !v8455ab;
assign v3759f23 = hlock4 & v3743604 | !hlock4 & v376992a;
assign v37419fd = hgrant6_p & v3736f2a | !hgrant6_p & v3a5d90a;
assign v372a9a6 = hbusreq4 & v3a6f79b | !hbusreq4 & v3a6bf41;
assign v375f8b0 = hgrant3_p & v3a71548 | !hgrant3_p & v375ac48;
assign v3743b12 = hmaster0_p & v3a62c0a | !hmaster0_p & v37412f3;
assign v3a6d8f4 = jx0_p & v23fde41 | !jx0_p & v376069d;
assign v372be74 = hlock5 & v3a713b5 | !hlock5 & v373fa48;
assign v3a70b91 = hlock4 & v3a6f8f7 | !hlock4 & v3729e32;
assign v375f5f0 = hlock5 & v3a63f9a | !hlock5 & v37551b2;
assign v372bf9f = hbusreq6 & v8455b0 | !hbusreq6 & v372d0ad;
assign v3757261 = hbusreq5_p & v3a56b72 | !hbusreq5_p & v3730b57;
assign v3723447 = hmaster3_p & v8455ab | !hmaster3_p & v3a63f77;
assign v3a6312c = jx0_p & v372a56e | !jx0_p & v360c3cc;
assign v3777642 = hbusreq2_p & v3a6963f | !hbusreq2_p & v8455b3;
assign v373d025 = hlock3_p & v37625a8 | !hlock3_p & v3a5ace5;
assign v3741a07 = hmaster0_p & v376374b | !hmaster0_p & v3a70f68;
assign v3764d17 = hbusreq3_p & v373df71 | !hbusreq3_p & v3a69671;
assign v3a5e7bf = hmaster1_p & v3769ae2 | !hmaster1_p & v2092b2c;
assign v1e37915 = hbusreq3 & v3a6ab5f | !hbusreq3 & !v3748900;
assign v3a56118 = hbusreq8 & v3a67aa1 | !hbusreq8 & v374d741;
assign v37477aa = hbusreq0 & v375bd37 | !hbusreq0 & v1e37cd6;
assign v3a645c2 = hmaster1_p & v3a68426 | !hmaster1_p & v372311c;
assign v3a5f546 = hbusreq7 & v3741736 | !hbusreq7 & v376ae9f;
assign v3750ac3 = hmaster1_p & v3734967 | !hmaster1_p & v3725ceb;
assign v372cde4 = hmaster2_p & v3728685 | !hmaster2_p & v37763d1;
assign v3a5baaf = hbusreq2_p & v37630d9 | !hbusreq2_p & !v3a658bf;
assign v3731e0e = hbusreq5 & v376ea5c | !hbusreq5 & v3753f1d;
assign v375517b = hmaster0_p & v3a5a039 | !hmaster0_p & v375f2f2;
assign v376ba2e = hgrant6_p & v3809e93 | !hgrant6_p & v377da26;
assign v3a6fc42 = hbusreq8 & v3a6deaa | !hbusreq8 & v38076b7;
assign v375e7bb = jx0_p & v3750e8a | !jx0_p & v3755596;
assign v377109a = hmaster0_p & v377e089 | !hmaster0_p & v3761fd6;
assign v3771ad8 = hmaster1_p & v3a6b60d | !hmaster1_p & v376b8c2;
assign v3807a92 = hbusreq0_p & v35772a5 | !hbusreq0_p & !v3a635ea;
assign v3a6dd8f = hbusreq8 & v3a6924d | !hbusreq8 & v8455ab;
assign v3a57d40 = hbusreq1_p & v2aca977 | !hbusreq1_p & v372886c;
assign v3a701a1 = hbusreq4_p & v3a5b289 | !hbusreq4_p & v376b15b;
assign v3a68d70 = hbusreq0 & v3741f69 | !hbusreq0 & v373c441;
assign v377b556 = hmaster2_p & v1e3828a | !hmaster2_p & v37390f9;
assign v3a6d749 = hlock1_p & v37764d7 | !hlock1_p & v3a5968c;
assign v3775626 = hbusreq2_p & v37385de | !hbusreq2_p & v3a637dd;
assign v3a5afd7 = hbusreq5_p & v3761fd7 | !hbusreq5_p & v8455ab;
assign v3a6f044 = hgrant6_p & v376d8d1 | !hgrant6_p & v8455ab;
assign v374bf69 = hmaster3_p & v3765d94 | !hmaster3_p & v3769a63;
assign v377d6e5 = hgrant3_p & v8455ab | !hgrant3_p & v3773c57;
assign v374407e = hmaster1_p & v377a18b | !hmaster1_p & v3728435;
assign v3762e66 = hlock0 & v3775999 | !hlock0 & v3730c0a;
assign v3a6fb4f = hlock7 & v3734279 | !hlock7 & v3748a0a;
assign v374f5e3 = hlock6 & v3768c4c | !hlock6 & v3a6beb6;
assign v3751931 = hbusreq2_p & v37636e4 | !hbusreq2_p & v3752af0;
assign v374094a = jx2_p & v376b934 | !jx2_p & v3a5f4a8;
assign v37682fc = hmaster2_p & v3769be7 | !hmaster2_p & v3a6a609;
assign v37598e6 = hgrant1_p & v8455b0 | !hgrant1_p & !v3723430;
assign v3a6fb23 = hbusreq7 & v3800ee4 | !hbusreq7 & v372871c;
assign v373c064 = hlock3 & v372f8c1 | !hlock3 & v375be64;
assign v377e156 = hbusreq5 & v3a6e52e | !hbusreq5 & v3808899;
assign v3a6ec1e = hbusreq2_p & v3748797 | !hbusreq2_p & v3764312;
assign v380911c = hbusreq4_p & v376daec | !hbusreq4_p & v3729c7e;
assign v380701a = hlock6_p & v3730e98 | !hlock6_p & v373cc68;
assign v3a712e9 = hbusreq5 & v3a540f8 | !hbusreq5 & v3737fca;
assign v373c978 = hgrant3_p & v376cd91 | !hgrant3_p & v2aca977;
assign v377bb66 = hgrant2_p & v374e6a5 | !hgrant2_p & v372731e;
assign cecaa5 = hgrant6_p & v3748d67 | !hgrant6_p & v3a6ed79;
assign v3a70a7e = hmaster2_p & v3a5b7c2 | !hmaster2_p & !v374a2cc;
assign v37c01ec = hbusreq5 & v3a6b5ea | !hbusreq5 & v8455ab;
assign v373f2b6 = hgrant4_p & v8455ab | !hgrant4_p & v3a70315;
assign v3a6fd47 = hbusreq3_p & v1e37869 | !hbusreq3_p & v8455ab;
assign v3728fee = hbusreq7_p & v373f8c4 | !hbusreq7_p & v1e37eb7;
assign v37717ea = hmaster2_p & v9bf1d8 | !hmaster2_p & v37711c3;
assign v37276a8 = hmaster2_p & v3a614b1 | !hmaster2_p & !v3a5dbd1;
assign v3753b6a = hbusreq0 & v3757695 | !hbusreq0 & v3768304;
assign v376cad6 = hlock2 & v373e7d9 | !hlock2 & v3809516;
assign v37499a0 = hbusreq5 & v32574c7 | !hbusreq5 & v3a6ff12;
assign v3a656b2 = hbusreq5_p & v372d925 | !hbusreq5_p & v376293f;
assign v377bf37 = hmaster2_p & v8455bb | !hmaster2_p & v3a7084e;
assign v372bbb3 = hgrant2_p & v3a5eadd | !hgrant2_p & v3a6e5f4;
assign v3a5dd7f = hlock0_p & v373b3fb | !hlock0_p & v8455b0;
assign v3a5dc5c = hlock8 & v3732a04 | !hlock8 & v373b17e;
assign v3a60638 = hbusreq2_p & v3747d3c | !hbusreq2_p & c0d46a;
assign v3a70cc3 = hbusreq2_p & v37666bd | !hbusreq2_p & v8455ab;
assign v3739731 = hbusreq8_p & v373f6b1 | !hbusreq8_p & v3743dc4;
assign v3748fba = hgrant2_p & v3a62524 | !hgrant2_p & v3a29842;
assign v374f9c5 = hgrant6_p & v3729214 | !hgrant6_p & v3758fe4;
assign v3724e67 = hbusreq3 & v3a6fbfc | !hbusreq3 & v372842d;
assign v3a29835 = hbusreq8_p & v3777631 | !hbusreq8_p & v376e66e;
assign v3a62424 = hbusreq5_p & v3a56a79 | !hbusreq5_p & v3a6bff5;
assign v3806828 = jx3_p & v3a5f375 | !jx3_p & !v373ec4c;
assign v3a6f07e = hgrant6_p & v37414b0 | !hgrant6_p & v3a66a6c;
assign v3722f85 = hbusreq2_p & a7afd8 | !hbusreq2_p & v8455ab;
assign v37577ab = hbusreq5 & v37296a5 | !hbusreq5 & v8455ab;
assign v377a343 = hbusreq6 & v37270d9 | !hbusreq6 & v8455e7;
assign v3772ae7 = hbusreq2 & v37538e4 | !hbusreq2 & v8455ab;
assign v377c2ce = hbusreq0 & v37549eb | !hbusreq0 & v8455ab;
assign v2092a89 = hlock7 & v3a70d78 | !hlock7 & v3a6f55d;
assign v375c9b9 = hlock5 & v3a5ae05 | !hlock5 & v377772d;
assign v39eb5ab = hbusreq6 & v3a6773a | !hbusreq6 & v35b774b;
assign v373632a = hmaster2_p & v376a6bc | !hmaster2_p & v3766202;
assign v3728867 = hbusreq5 & v3a66ca0 | !hbusreq5 & aac06c;
assign v376b47d = hlock1_p & v3761825 | !hlock1_p & v3a6e7e1;
assign v372b88d = hbusreq4 & v374362e | !hbusreq4 & v8455ab;
assign v377fada = hgrant4_p & b2eec3 | !hgrant4_p & v2092be1;
assign v3a653e4 = locked_p & v3a637dd | !locked_p & !v8455ab;
assign v3a68cc4 = hlock6_p & v3a56e63 | !hlock6_p & !v8455ab;
assign v3765ad4 = jx2_p & v3759203 | !jx2_p & v3a70583;
assign v3809ab5 = hlock7 & v3a5fbcb | !hlock7 & v374c28e;
assign v3a5b25b = hmaster0_p & v373a27c | !hmaster0_p & v3747afb;
assign v3a708c9 = hbusreq5 & v3a69a42 | !hbusreq5 & v3a61cb0;
assign v3a6c449 = hlock2 & v375a00a | !hlock2 & v376b6c9;
assign v3729dea = hbusreq5 & v3a60feb | !hbusreq5 & v3a6ff12;
assign be9654 = hbusreq4_p & v3a6f97d | !hbusreq4_p & v8455ab;
assign v3a6e581 = hmaster0_p & v376d078 | !hmaster0_p & v372a674;
assign v3a5e4e3 = hbusreq8 & b4389d | !hbusreq8 & v8455ab;
assign v3a5a48f = hmaster1_p & v3778a2f | !hmaster1_p & v372d3b2;
assign v8727d2 = hmaster3_p & v373fede | !hmaster3_p & !v3759d9c;
assign v3768343 = hlock5_p & v3a5fc33 | !hlock5_p & !v3a6f792;
assign v3754272 = hlock2_p & v3a6f343 | !hlock2_p & !v8455ab;
assign v3a61310 = hbusreq1 & v375f077 | !hbusreq1 & v8455ab;
assign v3a6fc03 = hbusreq4 & v3751734 | !hbusreq4 & !v8455ab;
assign v373bc30 = hlock0 & v373bd6c | !hlock0 & b5f474;
assign v3731aeb = hbusreq2 & v375fbc0 | !hbusreq2 & v8455ab;
assign v3a5fa81 = hbusreq0 & v3a67de4 | !hbusreq0 & v3a70722;
assign v3a6eb91 = hbusreq7 & v37508c4 | !hbusreq7 & v8455b3;
assign v373f687 = hbusreq5_p & v2e5fb38 | !hbusreq5_p & v3724696;
assign v377c4b8 = hgrant6_p & v8455ab | !hgrant6_p & !v377f118;
assign v376b269 = hlock0_p & v3a7126a | !hlock0_p & v3a635ea;
assign v3748f87 = hlock2_p & b4f302 | !hlock2_p & !v8455ab;
assign v3740923 = hbusreq7_p & v992750 | !hbusreq7_p & v8d3fe3;
assign v3a54ac1 = hmaster1_p & v37603d4 | !hmaster1_p & v373d245;
assign v3a6708d = hbusreq5 & v3740762 | !hbusreq5 & v3a5395c;
assign v3743ded = hbusreq6_p & v3a7038e | !hbusreq6_p & v374f6a0;
assign v3737202 = hmaster2_p & v3a635ea | !hmaster2_p & v3a62caa;
assign v3741abd = hgrant5_p & v3a6de60 | !hgrant5_p & v3725e33;
assign v373daa8 = hbusreq4_p & v377834b | !hbusreq4_p & v3a6f8de;
assign v3739915 = hmaster1_p & v37345a5 | !hmaster1_p & v8455ab;
assign v375309f = hlock0_p & v3a6b6f3 | !hlock0_p & v8455ab;
assign v376dd48 = hmaster0_p & v372fa3a | !hmaster0_p & v377d1dc;
assign v3a6b4ab = hlock4_p & v377989c | !hlock4_p & v3a6ffca;
assign v376a85d = hmaster0_p & v375a268 | !hmaster0_p & v377de6f;
assign v3735272 = hgrant4_p & v8455ab | !hgrant4_p & v3749a32;
assign v37791a7 = hbusreq2 & v3761909 | !hbusreq2 & v3a6fee9;
assign v3749207 = hlock0_p & v3751b0e | !hlock0_p & v3745020;
assign v374a681 = hbusreq3_p & c75852 | !hbusreq3_p & v8455ab;
assign v3732be9 = hmaster3_p & v3a65335 | !hmaster3_p & !v3743c90;
assign v375ef49 = hlock4 & v3a61a71 | !hlock4 & v3a5f7d7;
assign v3767c16 = hbusreq5_p & v3745b71 | !hbusreq5_p & !v8455ab;
assign v3a6f68f = hlock6_p & v3a712d6 | !hlock6_p & v8455ab;
assign v375f326 = hgrant2_p & v8455e7 | !hgrant2_p & !v3a6f0b2;
assign v375a51f = hbusreq5_p & v3756beb | !hbusreq5_p & v3a6f117;
assign v3a6ffa0 = hgrant3_p & v376015e | !hgrant3_p & v8455ab;
assign v3759de1 = hbusreq4_p & v3747c3d | !hbusreq4_p & v373d27a;
assign v3a5f55e = hmaster1_p & v9014db | !hmaster1_p & v376a92f;
assign v37424b8 = hmaster1_p & v37651b2 | !hmaster1_p & v3a708c1;
assign v376fbe3 = hmaster0_p & v3a6f63c | !hmaster0_p & v8455ab;
assign v3757b32 = hgrant2_p & v8455ab | !hgrant2_p & v373291c;
assign v37343dc = hbusreq4 & v374dc6d | !hbusreq4 & v37425a0;
assign v376a252 = hmaster1_p & v37333de | !hmaster1_p & v3a5b4ca;
assign v37699c7 = hbusreq5 & v3a6a352 | !hbusreq5 & v3778a97;
assign v373627b = hmaster3_p & v375452a | !hmaster3_p & v37449e7;
assign v3a5b8b0 = hlock4_p & v374f547 | !hlock4_p & v37770ed;
assign v372f6ab = hlock0_p & v37624a2 | !hlock0_p & v8455b0;
assign v37730ab = hbusreq7_p & v3726ec0 | !hbusreq7_p & v373824d;
assign v37291f4 = hmaster0_p & v3a71388 | !hmaster0_p & !v372b7a3;
assign v377ba29 = hmaster1_p & v377ea20 | !hmaster1_p & v3739904;
assign v374d42c = hbusreq3_p & v375068c | !hbusreq3_p & !v8455ab;
assign v360d18d = hbusreq2 & v3a6ffa0 | !hbusreq2 & v3a5b614;
assign v374158f = jx1_p & v376fb6e | !jx1_p & v374e06d;
assign v3a5ef9d = hmaster0_p & v3a58f56 | !hmaster0_p & v376cd84;
assign v37577d7 = hbusreq6 & v3a658c0 | !hbusreq6 & v8455ab;
assign v3a6e733 = hgrant7_p & v3a6ffde | !hgrant7_p & v375e3a1;
assign b1feb1 = hmaster0_p & v377957a | !hmaster0_p & v8455ab;
assign v376c31d = hmaster1_p & v377bf21 | !hmaster1_p & v377eab5;
assign v3a69961 = hgrant5_p & v3a60cf8 | !hgrant5_p & v3a68116;
assign v377bdd6 = hlock0_p & v377094b | !hlock0_p & v35b91b6;
assign v3723c99 = hmaster2_p & v373006f | !hmaster2_p & v3a71350;
assign v3a61237 = hbusreq1 & v3a70d71 | !hbusreq1 & v8455ab;
assign v2092aaa = hbusreq0 & c7f1d0 | !hbusreq0 & v3772828;
assign v3776d6e = hmaster2_p & v8455b0 | !hmaster2_p & v37685bb;
assign v375c170 = hbusreq4_p & v3728fe7 | !hbusreq4_p & v3a7169e;
assign c4d63a = hmaster0_p & v3747797 | !hmaster0_p & !v3777f6e;
assign v3754b6c = hbusreq0_p & v37502b7 | !hbusreq0_p & v3735e39;
assign v3a6af23 = hbusreq7_p & v37446b1 | !hbusreq7_p & v8455ab;
assign v3a54ba5 = hgrant6_p & v3739f07 | !hgrant6_p & v373e113;
assign v3722f16 = hgrant2_p & v3a709df | !hgrant2_p & v3734b15;
assign v3a6f8c7 = hbusreq5_p & v3777647 | !hbusreq5_p & v377b0b0;
assign v377a51b = hmaster2_p & v8455cb | !hmaster2_p & v3a706f1;
assign v3a6fc29 = hbusreq3 & v3a58429 | !hbusreq3 & v3736679;
assign v3a5b46d = hmaster2_p & v376430b | !hmaster2_p & !v8455e7;
assign v3732e39 = stateG10_1_p & v39ebac7 | !stateG10_1_p & v3a5ddd4;
assign v3a712ac = hbusreq6_p & v3747302 | !hbusreq6_p & v3a70905;
assign v375571e = hlock7 & a0a219 | !hlock7 & v3a6f4ea;
assign v3a6f83a = hgrant4_p & v8455ab | !hgrant4_p & v3a620d3;
assign v375f94a = hgrant4_p & v37245f8 | !hgrant4_p & v3a61535;
assign v3a54f04 = hbusreq0_p & v37356ce | !hbusreq0_p & v3807b40;
assign v3a70462 = hmaster2_p & v3a67a41 | !hmaster2_p & v3a70a04;
assign v376f9ac = hbusreq5_p & v373483e | !hbusreq5_p & v3a58c07;
assign v3764d26 = hmaster2_p & v377b461 | !hmaster2_p & v3a6f054;
assign v3758d1e = hbusreq5_p & v3a63f9a | !hbusreq5_p & v3737ceb;
assign v372be8e = hbusreq2_p & v377b24b | !hbusreq2_p & v375987b;
assign v3a5b581 = hbusreq6 & v3a704e5 | !hbusreq6 & v8455ab;
assign v37269f4 = hlock0_p & v373a841 | !hlock0_p & v8455e7;
assign v3a62236 = hmaster1_p & v376ef2d | !hmaster1_p & v377b774;
assign a56488 = hmaster3_p & v377a12e | !hmaster3_p & v374335b;
assign v37255e9 = hbusreq7_p & v3756087 | !hbusreq7_p & v23fda6c;
assign v37614c1 = hmaster2_p & v377bf77 | !hmaster2_p & v3a7129f;
assign v360bcf2 = hbusreq3_p & v3a5ee99 | !hbusreq3_p & v37355db;
assign v3777bcf = hbusreq5 & v3a7107e | !hbusreq5 & v374e4fa;
assign v3a546a2 = hmaster0_p & v3734dd6 | !hmaster0_p & v375f145;
assign v3a7041e = hbusreq2_p & v3736319 | !hbusreq2_p & v3a63597;
assign v373e219 = hmaster0_p & v372ab19 | !hmaster0_p & v373185b;
assign v37383c0 = hgrant2_p & v8455ab | !hgrant2_p & v376fc98;
assign v373164a = hbusreq4_p & v3a71077 | !hbusreq4_p & !v3764b0a;
assign v374f979 = hmaster0_p & v3a5fe3c | !hmaster0_p & v3730169;
assign v3763961 = locked_p & v3750746 | !locked_p & v3a637dc;
assign v3a70e01 = hgrant2_p & v3a5e544 | !hgrant2_p & v3744c29;
assign v3733dd3 = hgrant2_p & v37511c0 | !hgrant2_p & v3a68240;
assign v372995e = hmaster0_p & v372e083 | !hmaster0_p & v3a57e58;
assign v3a715c1 = hgrant4_p & v8455c2 | !hgrant4_p & v3740174;
assign v373059e = hlock4 & v373cdca | !hlock4 & v3a70e75;
assign v3a716a3 = hlock6_p & v3a6f5ea | !hlock6_p & v37406d2;
assign v3728d28 = hmaster1_p & v3736610 | !hmaster1_p & v3749a17;
assign v28896c8 = hgrant0_p & v376ea4a | !hgrant0_p & !v3a59720;
assign v37482be = hlock3_p & v8455ab | !hlock3_p & v37598c6;
assign v3a6ebb3 = hgrant4_p & v3a5aa3a | !hgrant4_p & v375791b;
assign v3744ef1 = hmaster2_p & v377308e | !hmaster2_p & v372d8f9;
assign v3723b33 = hmaster1_p & v3a635ea | !hmaster1_p & v3a70106;
assign v3a6ac7e = hlock2_p & v37711c8 | !hlock2_p & !v8455ab;
assign v372984c = hgrant6_p & v3a7138d | !hgrant6_p & v373ec0f;
assign v3724734 = hmaster2_p & v39ea76e | !hmaster2_p & v3759032;
assign v3a6425d = hbusreq4_p & v3725c63 | !hbusreq4_p & !v38074c2;
assign v3776b22 = hbusreq5_p & v8455bb | !hbusreq5_p & v3728738;
assign v372d8e8 = hgrant4_p & v3764276 | !hgrant4_p & v3766e29;
assign v37673a3 = hgrant7_p & v373ee8b | !hgrant7_p & v372b5ed;
assign v3a572e9 = hlock0 & v37496fa | !hlock0 & v377910a;
assign v37597f4 = hbusreq5_p & v3771cf7 | !hbusreq5_p & v373e873;
assign v3754ddd = hmaster2_p & v3a6ab5f | !hmaster2_p & !v8455ab;
assign v3a6f4c7 = hbusreq0 & v3a6f9c7 | !hbusreq0 & v373ca1a;
assign v3a660af = hgrant4_p & v3806b0a | !hgrant4_p & v8455ab;
assign v375208a = hgrant2_p & v3768b99 | !hgrant2_p & !v3740f70;
assign v3a6f309 = hbusreq0 & v374e19c | !hbusreq0 & v3764c8a;
assign v37431c0 = hgrant5_p & v3a714b7 | !hgrant5_p & v37358ae;
assign v3a6f081 = hbusreq4_p & v3a6ffc6 | !hbusreq4_p & !v8455ab;
assign v374cff2 = hmaster1_p & v37470c6 | !hmaster1_p & v37440e4;
assign v373a999 = hmaster1_p & v3a712e2 | !hmaster1_p & v3a6eb11;
assign v3a6f3be = hlock8 & v377fb55 | !hlock8 & v3724d8b;
assign v373b08f = hmaster1_p & v377ed2d | !hmaster1_p & v375a319;
assign v37391a1 = hbusreq6 & v3a58530 | !hbusreq6 & v3748797;
assign v376897b = hbusreq3_p & v37482be | !hbusreq3_p & v8455ab;
assign v3a6c15d = hbusreq7_p & v3a70cf5 | !hbusreq7_p & !v3a70bf9;
assign v3768500 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v376d68d;
assign v2619aa7 = hmaster0_p & v376894a | !hmaster0_p & v3a6f9a4;
assign v3808cf1 = hlock0 & v374a637 | !hlock0 & v3730043;
assign v3807472 = hbusreq7 & v8455b0 | !hbusreq7 & v3a6e69d;
assign v3a70820 = hmaster0_p & v3763f95 | !hmaster0_p & v373f694;
assign v372ab21 = hbusreq1_p & v375fa82 | !hbusreq1_p & v8455ab;
assign v376d680 = hmaster2_p & v372d727 | !hmaster2_p & v374b8fa;
assign v3768727 = hmaster1_p & v374314f | !hmaster1_p & v3734502;
assign v3a70097 = hmaster2_p & v3a5bf5f | !hmaster2_p & v3766b95;
assign v3a6599b = hgrant2_p & v375e7cc | !hgrant2_p & v375cab0;
assign v376d9ad = locked_p & v8455ab | !locked_p & v3a619c0;
assign v3772d8b = hgrant5_p & v8455c6 | !hgrant5_p & v372ba1c;
assign v3756f8c = hmaster0_p & v3a5a01b | !hmaster0_p & v373c545;
assign v375444a = hgrant4_p & v3a5d2d3 | !hgrant4_p & v374b15d;
assign v3771303 = hmaster1_p & v8455ab | !hmaster1_p & v375eeb9;
assign v3771933 = hmaster1_p & v374a36b | !hmaster1_p & v372c23b;
assign v375f014 = hmaster2_p & v375c8e6 | !hmaster2_p & v376e25b;
assign v3729139 = jx1_p & v374f7f8 | !jx1_p & v3a5de1e;
assign v374da7f = hgrant6_p & v377f09a | !hgrant6_p & v377915c;
assign v3a56200 = hlock5 & v37389ba | !hlock5 & v3a60924;
assign v372e332 = hmaster0_p & v3a63ea7 | !hmaster0_p & v3a70a33;
assign v3745db5 = hmaster0_p & v3743ff2 | !hmaster0_p & v372edf8;
assign v3759284 = hmaster1_p & v3a635ea | !hmaster1_p & v3806636;
assign b62018 = hmaster2_p & v8455ab | !hmaster2_p & !b1ca9b;
assign v3753353 = stateG10_1_p & v8455ab | !stateG10_1_p & v37551f2;
assign v3a6fd4e = hmaster0_p & v9ae45c | !hmaster0_p & v376e056;
assign v37796f6 = hlock2 & v3a6c8dc | !hlock2 & v375efc9;
assign v3777362 = hmaster0_p & v376058c | !hmaster0_p & v372dcf7;
assign v377acde = hbusreq8 & v377929d | !hbusreq8 & v3724974;
assign v374bc10 = hbusreq6_p & v372bf35 | !hbusreq6_p & !v38094e9;
assign v3a5642f = hmaster0_p & v37606b1 | !hmaster0_p & !v3a714d5;
assign v372d782 = hmaster1_p & v373e553 | !hmaster1_p & v37615d0;
assign v372f6f9 = hmaster1_p & v3a582c5 | !hmaster1_p & v3a71307;
assign v3734c5c = hmaster2_p & v3a70ecb | !hmaster2_p & v3770f75;
assign v3a6f0c9 = hbusreq4_p & v3a579a3 | !hbusreq4_p & v3a70d9c;
assign v3764de1 = hlock7_p & v3778e2d | !hlock7_p & !v3a6fb3e;
assign v3758c46 = hgrant0_p & v372493b | !hgrant0_p & !v374fa94;
assign v3a5a1e8 = hmaster0_p & v3a6f92f | !hmaster0_p & v99aa13;
assign v3a7148e = hlock0_p & v35b7808 | !hlock0_p & v8455b0;
assign v37784cc = hlock4_p & v376ff89 | !hlock4_p & v3a62550;
assign v3756ff6 = hlock7 & v372c5bc | !hlock7 & v3a6ff9a;
assign v374e3c1 = hbusreq8 & v3771ce2 | !hbusreq8 & v8455ab;
assign v375fa16 = hmaster2_p & v372391f | !hmaster2_p & !v376ea4a;
assign v37466a5 = hbusreq7_p & v37654a9 | !hbusreq7_p & v3777d70;
assign v3729e0b = hbusreq4 & v3a6f8de | !hbusreq4 & v3a62a6d;
assign v23fd84e = hmaster0_p & v3a59299 | !hmaster0_p & v374c164;
assign v372468b = hlock4_p & v35772b3 | !hlock4_p & v35772a6;
assign v3a65a52 = hmaster1_p & v3757966 | !hmaster1_p & v377843d;
assign v3a710fc = hlock6_p & v8455ab | !hlock6_p & !v373ad95;
assign v3a582ea = hbusreq5_p & v375a4d0 | !hbusreq5_p & v3a6f0d5;
assign v376d374 = hbusreq6_p & v37627bd | !hbusreq6_p & v8455ab;
assign v373a26e = busreq_p & v376f978 | !busreq_p & !v377c47d;
assign v3761fb5 = hbusreq6_p & v3756b39 | !hbusreq6_p & v374b73b;
assign v375e958 = hmaster1_p & v3a6a8ee | !hmaster1_p & v3a5dafb;
assign v375cfaa = hmaster1_p & v374502e | !hmaster1_p & v3a70647;
assign v372e83f = hbusreq3_p & v3a635ea | !hbusreq3_p & v375cf36;
assign v376ed36 = hbusreq8 & v3752d31 | !hbusreq8 & v3a60e5d;
assign v2092ac0 = hbusreq2_p & v3761c68 | !hbusreq2_p & v376073d;
assign v375d98c = hmaster1_p & v376501e | !hmaster1_p & v3a68b8a;
assign v374e26d = hgrant2_p & v8455b9 | !hgrant2_p & v3759abe;
assign v3773950 = hmaster2_p & v372c3d4 | !hmaster2_p & v8455ab;
assign v3762557 = hmaster2_p & v374b077 | !hmaster2_p & v3a6f8f5;
assign v3778962 = hgrant2_p & v8455ab | !hgrant2_p & v3753ca0;
assign v374170e = hgrant5_p & v376d52a | !hgrant5_p & v373c76c;
assign v376d658 = hbusreq2 & v377961f | !hbusreq2 & v8455ab;
assign v374d010 = hmaster1_p & v376c4c9 | !hmaster1_p & v3a6f54b;
assign v3a5bf28 = hgrant4_p & v8455c2 | !hgrant4_p & v3a5618d;
assign v3a6eee6 = hgrant3_p & v3733d6e | !hgrant3_p & v37485f0;
assign v3748d55 = hmaster0_p & v376151e | !hmaster0_p & v375f6c7;
assign v376f5ef = hlock2_p & v37467a6 | !hlock2_p & !v8455ab;
assign v3a6b4d7 = hgrant3_p & v8455be | !hgrant3_p & v3750025;
assign v374048c = hmaster2_p & v373cd16 | !hmaster2_p & v8455ab;
assign v3730ddd = hbusreq4_p & v3a6ad44 | !hbusreq4_p & !v8455ab;
assign v373e625 = hgrant4_p & v8455c2 | !hgrant4_p & v3a5fa81;
assign v37624e5 = hbusreq7 & v3a6f7e2 | !hbusreq7 & v376e9ed;
assign v3777197 = hbusreq4 & v3a61d83 | !hbusreq4 & v8455ab;
assign v375ec51 = hmaster1_p & v374fedc | !hmaster1_p & !v37350b2;
assign v3722a6f = hmaster0_p & v37390d6 | !hmaster0_p & v3a712d4;
assign v3725c60 = hmaster1_p & v3748451 | !hmaster1_p & v3a6ab55;
assign v3808658 = stateG10_1_p & v377d320 | !stateG10_1_p & v37583f2;
assign v32574c7 = hmaster0_p & v375a202 | !hmaster0_p & v3a6991b;
assign v376b0fd = hlock1_p & v20d166d | !hlock1_p & v8455ab;
assign v374d54c = hbusreq4_p & v3a6f0f9 | !hbusreq4_p & !v8455ab;
assign v3755ab8 = hlock8_p & v3779fbc | !hlock8_p & v3778ae9;
assign v37438ba = hmaster0_p & v3a5f6c2 | !hmaster0_p & v3736184;
assign v3a706b7 = hbusreq6_p & v377e56f | !hbusreq6_p & !v8455ab;
assign v2acae60 = hmaster2_p & v376b4e1 | !hmaster2_p & !v377df2e;
assign v3764e55 = hmaster1_p & v3807aa1 | !hmaster1_p & v3a6d329;
assign v3a70f1c = hgrant4_p & v3731320 | !hgrant4_p & v374c75e;
assign v3a612a4 = hlock4 & v375431d | !hlock4 & v377d6ba;
assign v374f52f = hmaster0_p & v375da9f | !hmaster0_p & v3774a9c;
assign v372e443 = hgrant4_p & v8455c2 | !hgrant4_p & v3a71213;
assign v376ab51 = hbusreq4 & v376b15b | !hbusreq4 & v3727084;
assign v3a54919 = hbusreq6_p & v3a635ea | !hbusreq6_p & v375d8e0;
assign v37481f3 = hgrant0_p & v3756261 | !hgrant0_p & v8455ab;
assign v376ae07 = hmaster2_p & v8455ab | !hmaster2_p & v377eb2d;
assign v377d491 = hbusreq5 & v3a6f6ea | !hbusreq5 & v372b5bc;
assign v375ced2 = hgrant4_p & v377ec59 | !hgrant4_p & v376df24;
assign v373e674 = hbusreq5_p & v37485e2 | !hbusreq5_p & v3757188;
assign v3a5ef3e = hbusreq4_p & v37259c7 | !hbusreq4_p & v35772a6;
assign v372b313 = hmaster3_p & v37415ea | !hmaster3_p & v377ebc9;
assign v3a669ae = hbusreq2 & v372e751 | !hbusreq2 & v8455ab;
assign v37598dc = hbusreq2_p & v3379035 | !hbusreq2_p & v35772a6;
assign v372da76 = hlock3 & v376be4c | !hlock3 & v3a6ca99;
assign v3a6186a = hbusreq6_p & v373f785 | !hbusreq6_p & v3a700fe;
assign v3765763 = hbusreq7_p & v3746b91 | !hbusreq7_p & v3a63cf3;
assign v3a6402e = hmaster2_p & v3a65b4a | !hmaster2_p & !v8455ab;
assign v3a5992f = hmaster2_p & v3a66534 | !hmaster2_p & v3757956;
assign v3a6fbb4 = hbusreq2_p & v37300b7 | !hbusreq2_p & v3a5f9ad;
assign v374e968 = hbusreq5 & v374640f | !hbusreq5 & v375b8cf;
assign v3732b12 = hbusreq2_p & v377ef7c | !hbusreq2_p & v3763acf;
assign v3739bfa = stateA1_p & v8455ab | !stateA1_p & !v3722f37;
assign v372dfc1 = hgrant6_p & v376e914 | !hgrant6_p & !v376fafe;
assign v3727889 = hmaster2_p & v3a6f942 | !hmaster2_p & v372b780;
assign v3a6fb03 = hbusreq5 & v37454c6 | !hbusreq5 & v3760513;
assign v3772c12 = hgrant6_p & v3a5a63c | !hgrant6_p & v3a704c9;
assign v376da5f = hmaster2_p & v3760881 | !hmaster2_p & v377d58d;
assign v374253f = hbusreq3_p & v3a70c97 | !hbusreq3_p & v8455ab;
assign v3a707f3 = hmaster0_p & v3a6fdd1 | !hmaster0_p & v3a71394;
assign v3a6fd9d = hgrant6_p & v372a51d | !hgrant6_p & v377eba4;
assign v3745fd1 = hmaster1_p & v864fe4 | !hmaster1_p & v376e358;
assign v3745abb = hbusreq5 & v3a67577 | !hbusreq5 & v8455ab;
assign v3724d8c = hmaster1_p & v3752428 | !hmaster1_p & v3766a64;
assign v37503f5 = hbusreq7 & v3775903 | !hbusreq7 & v3740a94;
assign v376f0cd = hbusreq8 & v3a6be38 | !hbusreq8 & v376ae9f;
assign v373f13e = hmaster3_p & v3a70430 | !hmaster3_p & !v376b1ee;
assign v37295a5 = hbusreq8 & v37710f3 | !hbusreq8 & !v37565d3;
assign v37645aa = jx1_p & v3738a94 | !jx1_p & v37662d7;
assign v3778ac6 = hgrant2_p & v377182c | !hgrant2_p & v377c29f;
assign v375a4eb = hmaster2_p & v3a635ea | !hmaster2_p & v3a710c8;
assign v3a6f766 = hbusreq7_p & v373db07 | !hbusreq7_p & !v2092b90;
assign v3a6e13d = hbusreq4_p & v377b774 | !hbusreq4_p & v3724e8e;
assign v3753097 = hmaster2_p & v8455ab | !hmaster2_p & v377f46d;
assign v374e3fa = hmaster1_p & v3a55081 | !hmaster1_p & v3733641;
assign v35b91b9 = hbusreq5_p & v3777647 | !hbusreq5_p & v3766309;
assign v37729db = hlock4 & v377d3b9 | !hlock4 & v3a55efa;
assign v3723f71 = hbusreq5 & v372715f | !hbusreq5 & !v3735936;
assign ae7027 = hbusreq3_p & v373cdb7 | !hbusreq3_p & v8455b7;
assign v3a6498e = hmaster0_p & v37676dc | !hmaster0_p & v3a676aa;
assign v3778ca0 = hbusreq5 & v3769af4 | !hbusreq5 & v8455ab;
assign v3756f17 = hbusreq4_p & v375b2d9 | !hbusreq4_p & v37712f8;
assign v3a63805 = hlock1_p & v8455b0 | !hlock1_p & !v8455ab;
assign v37656e5 = hmaster2_p & v8455ab | !hmaster2_p & v3776ada;
assign v8f64f2 = hlock6_p & v3732b75 | !hlock6_p & v3a6f9c3;
assign v3772c19 = hbusreq1_p & v373a8d6 | !hbusreq1_p & v377538f;
assign v3766996 = hbusreq3 & v375c806 | !hbusreq3 & v8455ab;
assign v3a6db7f = hlock5 & v3a62bcf | !hlock5 & v375a4ba;
assign v373c553 = jx2_p & v3776974 | !jx2_p & v3a5b945;
assign v3730818 = hbusreq3_p & v3753638 | !hbusreq3_p & v8455ab;
assign v3a5c57a = hbusreq5_p & v3733d3f | !hbusreq5_p & v3a70786;
assign v3738a5e = hgrant5_p & v8455ab | !hgrant5_p & v3a70863;
assign v373df91 = hbusreq7_p & v377d850 | !hbusreq7_p & v3a711fd;
assign v3779cf9 = hbusreq3_p & v375da10 | !hbusreq3_p & v376bb26;
assign v3a6ff2d = hgrant2_p & v8455ab | !hgrant2_p & v3741325;
assign v3a6d500 = hlock4 & v374748f | !hlock4 & v3a6f04c;
assign v373262e = hbusreq4_p & v39ebab4 | !hbusreq4_p & v373e814;
assign v375fe2b = hbusreq7 & v3735b64 | !hbusreq7 & v3774bad;
assign v3a6a199 = hmaster0_p & v3a5ae76 | !hmaster0_p & v376df4c;
assign v3a70525 = hbusreq4 & v3768349 | !hbusreq4 & v3a67cff;
assign v3a67221 = hbusreq6 & v372d2ad | !hbusreq6 & v8455ab;
assign v3a6fc83 = hbusreq4_p & v3a65aeb | !hbusreq4_p & v372d8f7;
assign v3a70504 = hbusreq6_p & v37518fb | !hbusreq6_p & v8455b0;
assign v3a7054c = hmaster0_p & v8455b3 | !hmaster0_p & v3a6f533;
assign v3777479 = hmaster1_p & v373014d | !hmaster1_p & v3a656ca;
assign v3a6fb0e = hbusreq5_p & v3a6e7ed | !hbusreq5_p & v3a707b2;
assign v374514c = hmaster2_p & v3a71232 | !hmaster2_p & v3750d06;
assign v373e21a = hlock0_p & v3a6ab5f | !hlock0_p & !v8455ab;
assign v3a6f1ae = hgrant2_p & v8455ba | !hgrant2_p & v3a6e138;
assign v376dc44 = hgrant4_p & v1e378b4 | !hgrant4_p & v374d63f;
assign v375431d = hbusreq4 & v377d6ba | !hbusreq4 & v38078ed;
assign v3a6f454 = hbusreq6_p & v3774c1b | !hbusreq6_p & !v38099c1;
assign v373d55f = hmaster2_p & v375f94a | !hmaster2_p & v3a7142f;
assign v374b364 = hmaster3_p & v3a635ea | !hmaster3_p & v377386a;
assign v3a6f748 = hgrant0_p & v8455ab | !hgrant0_p & v37625b7;
assign v372fe43 = jx1_p & v380a20c | !jx1_p & v3739916;
assign v377a571 = hmaster0_p & v8455b2 | !hmaster0_p & v8455ab;
assign v3755883 = hbusreq5 & v3731381 | !hbusreq5 & v37634cf;
assign v37376c1 = hbusreq6_p & v377cdea | !hbusreq6_p & v3759605;
assign v37720d8 = hlock3_p & v3745aff | !hlock3_p & v2acaf74;
assign v23fd8b2 = hmaster0_p & b62018 | !hmaster0_p & v8455ab;
assign v374a4cc = hgrant5_p & v3746f9d | !hgrant5_p & v3a647e0;
assign v376fad7 = hbusreq0 & v372f6ab | !hbusreq0 & v37591ac;
assign v375b7dc = hbusreq3 & v3a70a45 | !hbusreq3 & v376c343;
assign v3a5bb57 = hmaster1_p & v3723ac4 | !hmaster1_p & v3a5a807;
assign v3a595fd = hlock7 & v3a715b8 | !hlock7 & v37736c4;
assign v377e310 = hbusreq5_p & v3739a05 | !hbusreq5_p & v8455ab;
assign v3734810 = hbusreq7 & v3777479 | !hbusreq7 & v8455bf;
assign v3a67370 = hbusreq1_p & v37533d5 | !hbusreq1_p & v8455ab;
assign v375c8b0 = hgrant0_p & v3808e0d | !hgrant0_p & v8455ab;
assign v3a6f61c = hbusreq5 & v372ca99 | !hbusreq5 & v3a6f5eb;
assign v374b5d9 = hbusreq3_p & v376bb64 | !hbusreq3_p & v3a57e40;
assign v3a6fda8 = hgrant5_p & v3a578ef | !hgrant5_p & v3a70f3b;
assign v3769384 = hmaster1_p & v3778e3f | !hmaster1_p & v375b389;
assign v3766307 = hmaster2_p & v3747d68 | !hmaster2_p & v3744df8;
assign v3a6fbd7 = hlock0 & v37283bb | !hlock0 & v3756430;
assign v3750b86 = hmaster0_p & v3751069 | !hmaster0_p & v377a083;
assign v3a5eb0f = hmaster3_p & v3a6f710 | !hmaster3_p & v3763eb0;
assign v37235f1 = hbusreq8_p & v376a65b | !hbusreq8_p & da0ed3;
assign v3a606ee = hgrant3_p & v377dd3b | !hgrant3_p & v3766d11;
assign v3a6fe0c = hlock8_p & v372e684 | !hlock8_p & v8455cb;
assign v373ee70 = hgrant0_p & v3753edb | !hgrant0_p & a12203;
assign v3a62a68 = hmaster2_p & v8455ab | !hmaster2_p & v374a233;
assign v3a6ef4a = hgrant4_p & v3734067 | !hgrant4_p & v3a6fc46;
assign v3a628d4 = hmaster2_p & v3a7159a | !hmaster2_p & v3760700;
assign v3742d95 = hmaster2_p & v3a6143b | !hmaster2_p & v8455ab;
assign v3728127 = hbusreq0 & v373b88a | !hbusreq0 & v377c31d;
assign v37696b6 = hbusreq6_p & v3a635ea | !hbusreq6_p & v375cf36;
assign v3764825 = hbusreq0 & v3759edb | !hbusreq0 & v37454cc;
assign v3726980 = hbusreq7_p & v3a63f49 | !hbusreq7_p & v3a6b896;
assign v29256bb = hlock3 & v377b8b9 | !hlock3 & v3776ce0;
assign v3729933 = hlock5 & v3742a4b | !hlock5 & v373e93e;
assign v3a66cad = hbusreq5_p & v3766c68 | !hbusreq5_p & v2ff87d2;
assign v3741500 = hbusreq1 & v3755002 | !hbusreq1 & v8455ab;
assign v373fcae = hbusreq6_p & v373f704 | !hbusreq6_p & v3a6bbee;
assign v3757bf1 = hmaster1_p & v3779595 | !hmaster1_p & v3a6836a;
assign v3740df7 = hbusreq1_p & v3765d84 | !hbusreq1_p & !v3a5bbed;
assign v377aeba = hlock6 & v3740232 | !hlock6 & v373d91f;
assign v37440ff = hbusreq3_p & v374d3d7 | !hbusreq3_p & v3a5903a;
assign v9dc858 = stateG10_1_p & v372c11d | !stateG10_1_p & v373918a;
assign v2acb015 = hbusreq7 & v3765248 | !hbusreq7 & v3a6a8ee;
assign v3751440 = hmaster1_p & v8455ab | !hmaster1_p & v375e431;
assign v3765e5b = hbusreq5 & v375c600 | !hbusreq5 & v3763183;
assign v3a6008f = hbusreq4 & v376b8f1 | !hbusreq4 & v8455ab;
assign v376f9b5 = hbusreq6 & v3a6f30f | !hbusreq6 & v372462b;
assign v3a6a413 = hgrant5_p & b58331 | !hgrant5_p & v3a62812;
assign v3a6ef6f = hmaster0_p & v37444d4 | !hmaster0_p & v3a70caa;
assign v3a5b39d = hgrant6_p & v1e37cd6 | !hgrant6_p & v375a990;
assign v37586c0 = hbusreq6 & v373c8ff | !hbusreq6 & v8455ab;
assign v2ff9362 = hbusreq1 & v37482f8 | !hbusreq1 & !v3a709ea;
assign v3767537 = hbusreq7_p & v3a71618 | !hbusreq7_p & !v8455ab;
assign v377d428 = hmaster1_p & v3a635ea | !hmaster1_p & v3a6eb69;
assign v3a70376 = hlock3 & v3769404 | !hlock3 & v3776b61;
assign v3773729 = hmaster2_p & v3a63ea7 | !hmaster2_p & v3a6dc08;
assign v3763a86 = hgrant4_p & v3a70b92 | !hgrant4_p & v376c76d;
assign v3a67c8e = hbusreq5 & v373ee81 | !hbusreq5 & v3760513;
assign v3730e90 = hbusreq4_p & v373330f | !hbusreq4_p & v3763b0a;
assign v3754956 = jx0_p & v3a711f8 | !jx0_p & v3735ee1;
assign v37407f5 = hgrant2_p & v3a6b129 | !hgrant2_p & v373f051;
assign v3a65ea7 = hgrant5_p & v8455ab | !hgrant5_p & !v3773103;
assign v3751196 = hgrant3_p & v3a6432d | !hgrant3_p & v372c4bd;
assign v373a560 = jx0_p & v3a6eab8 | !jx0_p & v905dc4;
assign v37384ee = hgrant2_p & v3779e45 | !hgrant2_p & v3751e09;
assign v3773847 = hbusreq8_p & v3a676f1 | !hbusreq8_p & v3a70617;
assign v377e89a = hgrant7_p & v3773071 | !hgrant7_p & v375d57e;
assign v3774e41 = hbusreq4_p & v3747a97 | !hbusreq4_p & v37430e7;
assign v3a6eb47 = hbusreq6_p & v3762502 | !hbusreq6_p & v3a5bb64;
assign v377636a = hgrant3_p & v3a7000e | !hgrant3_p & v373a374;
assign v376575a = hmaster0_p & v8455ab | !hmaster0_p & v3a6fe6c;
assign v37474f3 = hgrant2_p & v3a5fdd3 | !hgrant2_p & !v3a569e1;
assign v374ddcd = hbusreq4_p & v3a66e96 | !hbusreq4_p & v3764998;
assign v3728c46 = hlock3_p & v3a6f882 | !hlock3_p & !v8455ab;
assign v377f4d5 = hlock5_p & v3a67a73 | !hlock5_p & v3a60a2b;
assign v3a703a0 = hgrant5_p & v3734579 | !hgrant5_p & v3740cb5;
assign v3a6ff25 = hbusreq0 & v3749435 | !hbusreq0 & v8455ab;
assign v377444e = hgrant5_p & v3a59d80 | !hgrant5_p & v3a6009a;
assign v377836a = hready & v3a593ee | !hready & v37496fa;
assign v3a70d43 = hmaster0_p & v3a706a8 | !hmaster0_p & v374e855;
assign v3a6ae19 = hbusreq8 & v373f6e7 | !hbusreq8 & v3a69b91;
assign v3743a49 = hbusreq5 & v372c6c4 | !hbusreq5 & v372d4d4;
assign v37536df = hbusreq0_p & v8455b0 | !hbusreq0_p & v3a6dc08;
assign v377696e = hlock8 & v377ace4 | !hlock8 & v3767153;
assign v2092b01 = hgrant2_p & v8df61b | !hgrant2_p & v3a5f9ad;
assign v38072dc = hmaster0_p & v376e661 | !hmaster0_p & v3a6230b;
assign v3759a7f = hgrant4_p & v375fbc6 | !hgrant4_p & v3a5ec7a;
assign v3a578e2 = hgrant4_p & v372b96c | !hgrant4_p & v3a6fc21;
assign v3a616cb = hmaster1_p & v372abd2 | !hmaster1_p & v372f7ca;
assign v372ff9e = hlock6_p & v3a57f42 | !hlock6_p & v373006f;
assign v3777e59 = hmaster1_p & v8455ab | !hmaster1_p & !v3730f21;
assign v3731857 = hbusreq4_p & v377766c | !hbusreq4_p & v374a8a5;
assign v3770174 = hmaster2_p & v3a5d678 | !hmaster2_p & v3a54eae;
assign v3a6f0f5 = hmaster0_p & v3754fcc | !hmaster0_p & v3a71614;
assign v3773341 = hbusreq8_p & v374ce04 | !hbusreq8_p & v8be8ac;
assign v3a582bc = hmaster1_p & v3a58cfc | !hmaster1_p & v374f52a;
assign v3a708ec = hbusreq1_p & v3725ef7 | !hbusreq1_p & v37728a4;
assign v3a7168c = jx0_p & v3a7145e | !jx0_p & v375b84e;
assign v373ec92 = hmaster1_p & v3a68426 | !hmaster1_p & v3a5844c;
assign v37255de = hbusreq6_p & v372cb42 | !hbusreq6_p & v37668e2;
assign v37645da = hgrant5_p & v8455c6 | !hgrant5_p & v373becf;
assign v374d802 = hgrant7_p & v3a70b4c | !hgrant7_p & v372cd50;
assign v3758ce2 = hmaster2_p & v374aec2 | !hmaster2_p & v37431ec;
assign b6b4ea = hgrant1_p & v3a6f333 | !hgrant1_p & v375aa47;
assign v376ee65 = hbusreq5_p & v376d4cb | !hbusreq5_p & v372433d;
assign v375c541 = hbusreq0_p & v3a56417 | !hbusreq0_p & v8455ab;
assign v39ebb64 = hbusreq4_p & v372abf1 | !hbusreq4_p & v376e0df;
assign v3744713 = hbusreq6_p & v377ea01 | !hbusreq6_p & v377c470;
assign v3a6efb2 = hlock0 & v3a6b53f | !hlock0 & v376f5b3;
assign v3730e01 = hmaster0_p & v3768d11 | !hmaster0_p & v3763c9c;
assign v37519e2 = hgrant5_p & v3a70d99 | !hgrant5_p & v3736c7e;
assign v3a67c41 = hgrant7_p & v3754740 | !hgrant7_p & v3738cd4;
assign v3a5d8bb = hmaster2_p & v373ff04 | !hmaster2_p & v372ba1c;
assign v376d896 = hbusreq5_p & v3735f9a | !hbusreq5_p & v8455ab;
assign v376629b = jx3_p & v3767a42 | !jx3_p & v3808904;
assign v3a64349 = hbusreq0 & v37450cb | !hbusreq0 & !v8455ab;
assign v37386c0 = hbusreq5_p & v3a62b09 | !hbusreq5_p & v3a702f1;
assign v3a6c64d = hbusreq5 & v3809968 | !hbusreq5 & v376508b;
assign v3a713b8 = hmaster2_p & v8455ab | !hmaster2_p & v3a6f910;
assign v373b3a8 = hbusreq4_p & v3a6a213 | !hbusreq4_p & !v373e8ad;
assign v372b77b = hbusreq4_p & v3a70778 | !hbusreq4_p & v8455cb;
assign v98bccb = hbusreq5_p & v376a619 | !hbusreq5_p & v8455ab;
assign v3a71402 = hbusreq3_p & v3773aa9 | !hbusreq3_p & v3a5a980;
assign v3a5b567 = hmaster0_p & v3a70fcf | !hmaster0_p & v3a7045e;
assign v374bfd2 = hgrant4_p & v3770032 | !hgrant4_p & v3a5cccf;
assign cb85ef = hgrant5_p & v8455ab | !hgrant5_p & v377a653;
assign v375e03c = hgrant6_p & v3a6f5d2 | !hgrant6_p & v2619b54;
assign v37466b7 = hmaster2_p & v3a6dc83 | !hmaster2_p & v3759c1f;
assign b05db7 = hmaster2_p & v35ba2da | !hmaster2_p & v375c671;
assign v372fca8 = hbusreq1 & v3a6fe6a | !hbusreq1 & !v8455ab;
assign v3735e84 = hgrant4_p & v8455c2 | !hgrant4_p & v3a565a8;
assign v3765e03 = hgrant4_p & v8455ab | !hgrant4_p & v375b82d;
assign v3728e1d = hbusreq6_p & v3a70ac8 | !hbusreq6_p & !v8455ab;
assign v3769199 = hlock7_p & v3a7010a | !hlock7_p & v376d0d8;
assign v3a6b72a = hgrant5_p & v37654e1 | !hgrant5_p & v377a57a;
assign v37510b1 = hbusreq2_p & v39a537f | !hbusreq2_p & !v9181c9;
assign v35b70a0 = hgrant1_p & v3733ec6 | !hgrant1_p & v374cda5;
assign v37c073f = hmaster0_p & v377d7a8 | !hmaster0_p & v3a6aa59;
assign v3a6fe1a = hbusreq1_p & v3774109 | !hbusreq1_p & !v8455ab;
assign v3a6efeb = hgrant4_p & v374db21 | !hgrant4_p & v3758e1c;
assign v3a651fc = hlock6 & v3774aa2 | !hlock6 & v375cf7d;
assign v3a6bf22 = hgrant4_p & v3a632aa | !hgrant4_p & v3a6fe33;
assign v3a706a4 = hgrant4_p & v8455ab | !hgrant4_p & v372ad4e;
assign v372361c = hready & v372e34d | !hready & v8455ab;
assign v3a63abb = hlock0_p & v37482f8 | !hlock0_p & v3a6eef6;
assign v3a56e15 = hgrant8_p & v3a6f64c | !hgrant8_p & v3a62f59;
assign v37668e2 = hgrant2_p & v3a5eadd | !hgrant2_p & v3729829;
assign v3a64293 = hgrant5_p & v3a6e82d | !hgrant5_p & v373ff9a;
assign v3730d6e = hmaster0_p & v8455e7 | !hmaster0_p & v3a7056e;
assign v37c014f = hmaster0_p & v1e37b74 | !hmaster0_p & v3759bd0;
assign v37571ad = hbusreq6_p & v3a6f43e | !hbusreq6_p & v372935c;
assign v3774209 = hbusreq6 & v3a6cf19 | !hbusreq6 & v3a70c74;
assign v3a700c1 = hmaster1_p & v3a69390 | !hmaster1_p & v3a71373;
assign v3a6fd20 = hgrant5_p & v3740bf7 | !hgrant5_p & v376a252;
assign v3725649 = hbusreq2_p & v375baed | !hbusreq2_p & v3779e66;
assign v3a618f6 = hbusreq8 & v8455e7 | !hbusreq8 & v8455ab;
assign v3733a1e = hmaster2_p & v3767437 | !hmaster2_p & v3760f4e;
assign v3a70658 = jx3_p & v3a6f8c6 | !jx3_p & v37503e7;
assign v376e074 = hmaster0_p & v3a5e24e | !hmaster0_p & v373afd0;
assign v3779ff0 = hmaster0_p & v377e453 | !hmaster0_p & v3728fda;
assign v3748443 = hmaster3_p & v38072bc | !hmaster3_p & v92bc1e;
assign v374e0a9 = hmaster2_p & v377f548 | !hmaster2_p & v373893a;
assign v3740052 = hmaster1_p & v8455ab | !hmaster1_p & v3a63f9a;
assign v3a6fc66 = hbusreq0 & v3a70c39 | !hbusreq0 & v3a704cc;
assign v3743ab6 = hbusreq8 & v375b278 | !hbusreq8 & v8455ab;
assign v3722ee2 = hlock3_p & v2ff9190 | !hlock3_p & v8455ab;
assign v376021f = hlock2_p & v377efac | !hlock2_p & v37406d2;
assign v37695c1 = hbusreq8 & v37470fc | !hbusreq8 & v373b8c6;
assign v3779316 = hbusreq4 & d8a786 | !hbusreq4 & v375f504;
assign v3a5455e = hmaster0_p & v377437d | !hmaster0_p & v37582c2;
assign v3a7165b = hbusreq4 & v3768ecc | !hbusreq4 & v8455e7;
assign v3a6ea3b = hbusreq4_p & v37337d2 | !hbusreq4_p & v3731230;
assign v376fbfd = hlock5 & v38095b1 | !hlock5 & v3a71574;
assign v3723f45 = hbusreq8 & v3a69761 | !hbusreq8 & v3a71478;
assign v374016f = hbusreq5_p & v37297c0 | !hbusreq5_p & v3766d53;
assign v3728a6d = hmaster1_p & v37485cb | !hmaster1_p & v3753e23;
assign v3a6e592 = hbusreq0_p & v376dbdf | !hbusreq0_p & !v372fc81;
assign v3767c46 = hbusreq4 & v3a6f567 | !hbusreq4 & v374a637;
assign v3a5d431 = hmaster0_p & v3757568 | !hmaster0_p & v3a5e8a1;
assign v3a6fe8c = hbusreq7_p & v3762a68 | !hbusreq7_p & v3a6ef70;
assign v376e89b = hbusreq2_p & v373e689 | !hbusreq2_p & v8455ab;
assign v3a7115e = hmaster2_p & v3a6f998 | !hmaster2_p & v37431ec;
assign v3a66051 = hlock3 & v3a6fed3 | !hlock3 & v376c8ea;
assign v3a708dd = hgrant6_p & v3777996 | !hgrant6_p & v3739e70;
assign v3750859 = hgrant3_p & v3a69487 | !hgrant3_p & v373d8e5;
assign v3779c33 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v292555a;
assign v3a71096 = hbusreq8 & v2ff8f77 | !hbusreq8 & v3a71504;
assign v37766cf = hmaster0_p & v3777149 | !hmaster0_p & !v373e15b;
assign v373b42d = hbusreq7 & v37702e0 | !hbusreq7 & v3768734;
assign v3a67833 = hlock0 & v372348c | !hlock0 & v377c079;
assign v373bd24 = hlock0_p & v373a27c | !hlock0_p & v37566b2;
assign v3726d2a = hgrant2_p & v372ec1c | !hgrant2_p & v377dabc;
assign v3759cce = hlock2_p & v376ba4d | !hlock2_p & v8455b0;
assign v3738d0b = hlock2 & v376195f | !hlock2 & v37251b9;
assign v3a6f940 = hbusreq3 & v3760740 | !hbusreq3 & v8455ab;
assign v372c83f = hbusreq6 & v3a5b359 | !hbusreq6 & v8455ab;
assign v37667f8 = hbusreq5_p & v375e512 | !hbusreq5_p & v3a713ad;
assign v375a94d = hready_p & v3773343 | !hready_p & !v3a58546;
assign v3740f7d = hlock6_p & v375444e | !hlock6_p & v373006f;
assign v3a5c473 = hmaster2_p & v373f058 | !hmaster2_p & v373ee80;
assign v375c3b6 = hlock5 & v3736fb4 | !hlock5 & v376e74b;
assign v3a6d4cd = hbusreq8 & v375d1d0 | !hbusreq8 & v375986d;
assign v376fcd6 = hbusreq5_p & v3762873 | !hbusreq5_p & v37327c3;
assign v3a71077 = hbusreq0 & v3a68f16 | !hbusreq0 & v8455ab;
assign v3a70719 = hbusreq8 & v374cffd | !hbusreq8 & v3737808;
assign v3a6f833 = hmaster2_p & v3a6f781 | !hmaster2_p & v37769cc;
assign v3750ef8 = hgrant6_p & v3a6fd6a | !hgrant6_p & v3a62589;
assign v3776196 = hgrant4_p & v8455ab | !hgrant4_p & v35b7769;
assign v3a66039 = hmaster3_p & v376a74a | !hmaster3_p & !v376b1ee;
assign v373f75b = hmaster2_p & v377d9aa | !hmaster2_p & !v3777a00;
assign v3a6356b = hgrant2_p & v375c7b9 | !hgrant2_p & !v3a6e9c0;
assign v3a601cd = hmaster1_p & aa783c | !hmaster1_p & v374d7dc;
assign v3774c98 = hmaster2_p & v374f0c1 | !hmaster2_p & !v3a63e82;
assign v375d8ea = hbusreq2_p & v3762d5f | !hbusreq2_p & v8455b0;
assign v377568c = hbusreq3_p & v8455ab | !hbusreq3_p & v3a714c3;
assign b04260 = hbusreq4 & v373c7a5 | !hbusreq4 & v3775999;
assign v3a64103 = hmaster3_p & v375fea8 | !hmaster3_p & v3a70122;
assign v3731517 = hbusreq7 & v375f2e8 | !hbusreq7 & v3a6f1c8;
assign v372c197 = hgrant6_p & v3a637dc | !hgrant6_p & v3a60bbf;
assign v3a58a39 = hlock6_p & v8455ab | !hlock6_p & !v3a6ac26;
assign v373fef5 = hgrant2_p & v377eaf2 | !hgrant2_p & v8455ab;
assign v3764994 = hlock2 & v373a802 | !hlock2 & v377c929;
assign v376b8f8 = hbusreq0 & v3a5e3be | !hbusreq0 & v3a57d9e;
assign v3a59217 = hgrant4_p & v325c9cb | !hgrant4_p & !v3a715f2;
assign v3757ffa = hmaster2_p & v8455ab | !hmaster2_p & v3765321;
assign v3a70ad3 = hmaster2_p & v37696fe | !hmaster2_p & v3751491;
assign v377de29 = hmaster0_p & v374306c | !hmaster0_p & v3a6db2d;
assign v3a6f9d3 = hbusreq5 & v375a92d | !hbusreq5 & v374193d;
assign v372525e = hmaster2_p & v37566b2 | !hmaster2_p & !v39a5381;
assign v3a6a367 = hlock7 & v3735ba1 | !hlock7 & v3a71556;
assign v374083d = hmaster0_p & v3a5e24e | !hmaster0_p & v3a704b4;
assign v3a70392 = hmaster3_p & v3a70d48 | !hmaster3_p & v3750e8a;
assign v3a645df = hbusreq4 & v3779002 | !hbusreq4 & v8455ab;
assign v3a70e3f = hmaster2_p & v8455ab | !hmaster2_p & v3a62015;
assign v3746b7f = hmaster2_p & v3a5b5d3 | !hmaster2_p & v3a6eb39;
assign v373f6e7 = hlock7 & v374a189 | !hlock7 & v3a710ea;
assign b1ca9b = hbusreq3_p & v3a5ba6d | !hbusreq3_p & !v8455ab;
assign v3a651c8 = hlock8 & v3a70e54 | !hlock8 & v3a5d6f3;
assign v37712aa = hmaster2_p & v3a70374 | !hmaster2_p & v3722bca;
assign v375b344 = jx0_p & v3a701f3 | !jx0_p & v37392d7;
assign v37425a7 = hlock2 & v37791a7 | !hlock2 & v3761909;
assign v3a66c34 = hmaster1_p & v374d383 | !hmaster1_p & !v8455ab;
assign v372a886 = hgrant6_p & v3806821 | !hgrant6_p & v376b903;
assign v3a6fe57 = jx0_p & v8455ab | !jx0_p & v3a6cad7;
assign v3749336 = hmaster2_p & v373ee52 | !hmaster2_p & v3750adf;
assign v3757c37 = hbusreq2_p & v3a59275 | !hbusreq2_p & v3a70bc7;
assign v373cdca = hbusreq4 & v3a70e75 | !hbusreq4 & v3779cf9;
assign v377c58e = hmaster2_p & v37334a3 | !hmaster2_p & v3a71016;
assign v3773871 = hgrant0_p & v8455ab | !hgrant0_p & v3a65f3e;
assign v375a30e = hmaster1_p & v37653a2 | !hmaster1_p & v377d080;
assign v3a5d30d = hbusreq7_p & v373d64d | !hbusreq7_p & !v3577344;
assign v3752e71 = hlock2 & v37430c2 | !hlock2 & v37300c9;
assign v372a9c2 = hmaster3_p & v374831d | !hmaster3_p & !v372c23f;
assign v377936c = hbusreq5_p & v3738d19 | !hbusreq5_p & !v37443a2;
assign v37693cf = hgrant3_p & v360d1cb | !hgrant3_p & v3a7045c;
assign v3738f1b = hgrant5_p & v3761915 | !hgrant5_p & v3743c35;
assign v37592ca = hbusreq0 & v3a711de | !hbusreq0 & v373a68a;
assign v374e078 = jx0_p & v377119f | !jx0_p & v3741ea8;
assign v3a56d26 = hbusreq4_p & v372810e | !hbusreq4_p & v3a6abe5;
assign v37778a2 = hgrant4_p & v8455ab | !hgrant4_p & v3726344;
assign v33782fe = hmaster1_p & v3a70209 | !hmaster1_p & v3a70cd6;
assign v374a407 = hgrant6_p & v376f175 | !hgrant6_p & v373a29c;
assign v37659c6 = hmaster1_p & v3a7010c | !hmaster1_p & !v8455bf;
assign v377cf67 = hbusreq4_p & v373104a | !hbusreq4_p & v3a7113a;
assign v3809400 = hbusreq4_p & v3722d9d | !hbusreq4_p & v3a60cdb;
assign v3a6f061 = hbusreq4_p & v3757009 | !hbusreq4_p & v375a677;
assign v3726088 = hmaster1_p & v372cdde | !hmaster1_p & c4d24d;
assign v373c99b = hbusreq2_p & v3a66d7b | !hbusreq2_p & v3a56094;
assign v375cb72 = hbusreq2_p & v3a64b41 | !hbusreq2_p & v372e88a;
assign v375d15c = hbusreq5 & v3a71608 | !hbusreq5 & v3a71530;
assign v3a68f4d = hlock2 & v3a5a2e2 | !hlock2 & v3a6d810;
assign v376d23f = hlock8 & d950cb | !hlock8 & v37629fc;
assign v3808f73 = hmaster2_p & v3725198 | !hmaster2_p & v3a710c6;
assign v37242fa = hbusreq7 & v3a70d7e | !hbusreq7 & v3a635ea;
assign v372673d = hgrant4_p & v3a635ea | !hgrant4_p & v377704c;
assign v3759947 = hgrant0_p & v3a6fdef | !hgrant0_p & v3748cbd;
assign v3745e5e = hmaster1_p & v8455ab | !hmaster1_p & v373300a;
assign v3777a00 = hbusreq4 & v376b21a | !hbusreq4 & v8455ab;
assign v377c0bd = hmaster0_p & v3733c53 | !hmaster0_p & v37766fb;
assign v89b450 = hmaster0_p & v377d766 | !hmaster0_p & v372840a;
assign v3732706 = hgrant2_p & v8455ab | !hgrant2_p & v3a637e0;
assign v2ff8e8b = hmaster2_p & v8455ab | !hmaster2_p & v3a5a807;
assign v3a701ad = hmaster1_p & v2acafaa | !hmaster1_p & v8455ab;
assign v375452a = jx0_p & v375c551 | !jx0_p & v3750e4b;
assign v38071c1 = hgrant1_p & v3a5c945 | !hgrant1_p & !v376ba47;
assign v376f48d = hbusreq6 & v3a6f778 | !hbusreq6 & v8455ab;
assign v3743f94 = hlock3_p & v377d3e4 | !hlock3_p & v37509c7;
assign v3a5d548 = hmaster2_p & v3733da4 | !hmaster2_p & v37786a6;
assign v377fabc = hbusreq1_p & v3378a0a | !hbusreq1_p & v3742f38;
assign v39a4dac = hbusreq4_p & v373f7ff | !hbusreq4_p & !v8455ab;
assign v38072a2 = hmaster0_p & v3772347 | !hmaster0_p & v3a5ae95;
assign dbdbc5 = hbusreq2_p & v377bd97 | !hbusreq2_p & !v373acce;
assign v375bca7 = hmaster1_p & v37410bd | !hmaster1_p & v3a6f937;
assign v3a59b5f = hgrant6_p & v3771fb3 | !hgrant6_p & v3a663c7;
assign d284a6 = hbusreq3_p & v38072fd | !hbusreq3_p & v3a64474;
assign v3772ab6 = hmaster0_p & v8455ab | !hmaster0_p & v3a68b6c;
assign d9767c = hlock0_p & v3a5e3d3 | !hlock0_p & v373541f;
assign v38079d5 = hbusreq5 & v3a704b6 | !hbusreq5 & v8455ab;
assign v35b7189 = hgrant2_p & v377b6ce | !hgrant2_p & v373ff58;
assign v3730ae3 = hbusreq6_p & v3745f76 | !hbusreq6_p & v3a701e4;
assign v3741c4b = hmaster0_p & v3a5bf5f | !hmaster0_p & v37317f2;
assign v372f391 = hlock3_p & v376bf69 | !hlock3_p & v8455b0;
assign v37235ee = hlock6_p & v8455ab | !hlock6_p & v3a56864;
assign v373dbfe = hmaster2_p & v3a5b469 | !hmaster2_p & v3a6ff2c;
assign v3a63c3b = hlock5_p & v3a71580 | !hlock5_p & v374fa8c;
assign v3754d67 = hmaster1_p & v3a5a807 | !hmaster1_p & v3a572ea;
assign v377ad8f = hgrant0_p & v372802c | !hgrant0_p & v3742101;
assign v376f332 = hlock0_p & v373ad3c | !hlock0_p & v377a63c;
assign v377eab7 = hlock5 & v3724b8c | !hlock5 & v3a711cb;
assign v375dfc6 = hbusreq8_p & v376eaed | !hbusreq8_p & v374464b;
assign a6f1de = hbusreq2_p & v377bc89 | !hbusreq2_p & v3735c5d;
assign v374da1a = hmaster2_p & v8455c2 | !hmaster2_p & v3a5d94a;
assign v3a5a47b = hbusreq5 & v3a5b9d6 | !hbusreq5 & v373790d;
assign v3754892 = hmaster0_p & v37233a2 | !hmaster0_p & v3a71420;
assign v377376d = hmaster2_p & v3a715ac | !hmaster2_p & v3a6b575;
assign v3a70065 = hbusreq2_p & v3743cb5 | !hbusreq2_p & v8455b0;
assign v377349f = hgrant6_p & v8455ab | !hgrant6_p & v374d2b3;
assign v3a674c9 = hbusreq7 & v3a6f6d1 | !hbusreq7 & v8455ab;
assign v374b18c = hgrant6_p & v3a702bb | !hgrant6_p & v374b43d;
assign v37351f5 = hgrant4_p & v8455ab | !hgrant4_p & v3758c06;
assign v3736421 = hbusreq5 & v372f309 | !hbusreq5 & v3a5fc34;
assign v374e28d = hbusreq4 & v3730fcd | !hbusreq4 & v8455ab;
assign v3746f9d = hmaster1_p & v3a635ea | !hmaster1_p & v3a5584b;
assign v3754e33 = hbusreq8_p & v3730289 | !hbusreq8_p & v3a5d30d;
assign v377d004 = hmaster0_p & v3a6f9cb | !hmaster0_p & v3a6fbd1;
assign v3a5dfa3 = hgrant5_p & v8455ab | !hgrant5_p & v3a703e2;
assign v37317b4 = hgrant7_p & v8455ce | !hgrant7_p & v374c058;
assign v3730646 = hgrant2_p & v3a5f50e | !hgrant2_p & v375b506;
assign v37296cd = hmaster0_p & v35b774b | !hmaster0_p & v374834b;
assign v377097a = hbusreq3_p & v3806d42 | !hbusreq3_p & v8455ab;
assign v377167e = hbusreq2_p & v373ac52 | !hbusreq2_p & !v8455ab;
assign v3753f37 = hlock2_p & v3a6f782 | !hlock2_p & !v8455ab;
assign v377a75f = hbusreq7_p & v376b063 | !hbusreq7_p & v376d432;
assign v373d09a = hlock7_p & v3a714b7 | !hlock7_p & !v3748984;
assign v3769fa2 = hbusreq7_p & v377b920 | !hbusreq7_p & v3a66373;
assign v372b8a0 = hbusreq5_p & v3753b1b | !hbusreq5_p & v8455ab;
assign v3730a90 = hmaster1_p & v3767c16 | !hmaster1_p & !v373a265;
assign v3741c03 = hbusreq1_p & v375f6f6 | !hbusreq1_p & !v3a6f133;
assign v372998e = hmaster0_p & v376dafa | !hmaster0_p & !v373a3c8;
assign v375790e = hmaster1_p & v37735b8 | !hmaster1_p & v3a70bbe;
assign v375a8ad = hlock4 & v3735ad2 | !hlock4 & v3a5dc35;
assign v377f584 = hbusreq4_p & v3760f64 | !hbusreq4_p & v377fc4b;
assign v3a71486 = hmaster2_p & v9af7ec | !hmaster2_p & v374da61;
assign v37749c3 = hgrant6_p & v8455ab | !hgrant6_p & v3a6f151;
assign v3763c1f = hbusreq8 & v3a7031e | !hbusreq8 & v374a4c2;
assign v374c2e1 = hbusreq8_p & v37739ba | !hbusreq8_p & v3a66819;
assign v374d88f = hbusreq4 & d305e8 | !hbusreq4 & v376498f;
assign v3a543c5 = hmaster0_p & v3771507 | !hmaster0_p & v377d280;
assign v374212c = hbusreq2 & v37674c1 | !hbusreq2 & !v8455ab;
assign v3731de2 = hbusreq4 & v372ee9a | !hbusreq4 & v3a6be44;
assign v3a6f0e9 = hbusreq6_p & v3a56c2e | !hbusreq6_p & v3778528;
assign v3a714f0 = hlock0_p & v8a7f7e | !hlock0_p & v373040e;
assign v3759b11 = hbusreq2 & v375d9f8 | !hbusreq2 & !v3766238;
assign v377aecd = hmaster1_p & v3a679e2 | !hmaster1_p & v37629b0;
assign v3a6d922 = stateG10_1_p & v8455e7 | !stateG10_1_p & v3774c11;
assign v3a6d2d7 = hmaster0_p & v3a6fbcb | !hmaster0_p & v3a6fb52;
assign v377d280 = hmaster2_p & v3771507 | !hmaster2_p & v8455ab;
assign v3729b6a = hgrant6_p & v8455ab | !hgrant6_p & v3753b3f;
assign v3a5dc2a = hmaster1_p & v372d727 | !hmaster1_p & v3a54478;
assign v377bbf7 = hmaster2_p & v373127e | !hmaster2_p & v3a6fb2b;
assign v3a6ffab = hbusreq6 & v374944b | !hbusreq6 & v374f35a;
assign v3756430 = hlock4 & v3a540a4 | !hlock4 & v3a712ac;
assign v3750797 = hgrant5_p & v375634b | !hgrant5_p & v376755f;
assign v373dc53 = hmaster1_p & v8455ab | !hmaster1_p & v3747d42;
assign v1e38239 = hgrant2_p & v8455ba | !hgrant2_p & v3767feb;
assign v3a69bbd = hgrant6_p & v377a42f | !hgrant6_p & v3a56593;
assign v3a67519 = hgrant6_p & v3a70283 | !hgrant6_p & !v377c3ea;
assign v3a642cf = hbusreq1_p & v3a5b9ba | !hbusreq1_p & v35772a6;
assign v377514f = hgrant0_p & v8455b5 | !hgrant0_p & v3a6d93d;
assign v3a70902 = hmaster2_p & v3a71133 | !hmaster2_p & v37307d4;
assign v3a5e7c4 = hmaster2_p & v37432cd | !hmaster2_p & v3a71026;
assign v3a5b719 = hmaster0_p & v37400d2 | !hmaster0_p & !v374da92;
assign v3a70d76 = hmaster3_p & v3a706ef | !hmaster3_p & v2acaf12;
assign v372869e = hgrant3_p & v8455be | !hgrant3_p & v374ed51;
assign v376866e = hlock0_p & v37502b7 | !hlock0_p & v3732c52;
assign v3a5d46c = hbusreq4_p & v376856b | !hbusreq4_p & v3a70c52;
assign v374e2a1 = hready & v3a7098c | !hready & v3748797;
assign v3764998 = hbusreq0 & v37322ca | !hbusreq0 & v1e37cd6;
assign v3a708bd = hbusreq6_p & v377094b | !hbusreq6_p & v3a71422;
assign v372c3c7 = hmaster0_p & v380909e | !hmaster0_p & v3769923;
assign v3a70c1a = hgrant6_p & v8455ab | !hgrant6_p & v3776bb6;
assign v3745cf8 = hmaster1_p & v3a6f6bc | !hmaster1_p & v3765d2b;
assign v3a59461 = hbusreq4 & v8455b0 | !hbusreq4 & v3755791;
assign v3a71410 = hgrant4_p & v3a6616c | !hgrant4_p & v3a5ec7a;
assign v37794fa = hgrant0_p & v377682d | !hgrant0_p & !v3770e2b;
assign v3772af6 = hbusreq0_p & v3760f87 | !hbusreq0_p & !v3a5ef5c;
assign v373da6d = hmaster1_p & v37737aa | !hmaster1_p & v377f64b;
assign v3775269 = hbusreq4_p & v3a6efef | !hbusreq4_p & v8455ab;
assign v325c976 = hgrant3_p & v375a293 | !hgrant3_p & v8455ab;
assign v3a6d625 = hbusreq0 & v3a634db | !hbusreq0 & v3a55f42;
assign c6598e = hgrant2_p & v8455e7 | !hgrant2_p & !v3768d79;
assign v372e4ac = hbusreq5 & v372e4a7 | !hbusreq5 & v374a369;
assign v3a68ad8 = hgrant3_p & v3a709c1 | !hgrant3_p & v8455ab;
assign v377a6e2 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3a6d665;
assign v372c345 = hbusreq8 & v376d36a | !hbusreq8 & v3733b90;
assign v377a2f2 = hmaster2_p & v37482f8 | !hmaster2_p & v3759158;
assign v374e784 = hmaster0_p & v3748489 | !hmaster0_p & v377291b;
assign v3750746 = busreq_p & v3a637dc | !busreq_p & v372fc17;
assign v3779a9a = hmaster1_p & v3a587be | !hmaster1_p & v3745b39;
assign v3a65161 = hbusreq1_p & v37583f2 | !hbusreq1_p & v3808658;
assign v373b14a = hlock0 & v3a6fba8 | !hlock0 & v3a70b91;
assign v3748f48 = hgrant3_p & v3a5872a | !hgrant3_p & v3a6fd17;
assign v3a6fcf5 = hlock7 & v3748e6a | !hlock7 & v372f1a8;
assign v3a7079d = hmaster1_p & v3743ff2 | !hmaster1_p & v376d33b;
assign v374776b = hbusreq5_p & v39ebacc | !hbusreq5_p & v8455ab;
assign v3a682f7 = hmaster1_p & a747d7 | !hmaster1_p & v3a5aa33;
assign v37390d5 = hbusreq5 & v3a69f0e | !hbusreq5 & !v8455b5;
assign v37278c8 = hbusreq3_p & v3a68523 | !hbusreq3_p & v3770f51;
assign v3a58588 = hmastlock_p & v3a6affa | !hmastlock_p & v8455ab;
assign v3a6f210 = busreq_p & v35772a5 | !busreq_p & v3577306;
assign v3765d27 = hgrant5_p & v3747b4e | !hgrant5_p & v375d8af;
assign v3a6f692 = hmaster2_p & v3a6fe0d | !hmaster2_p & !v39a4ca8;
assign v3a667a7 = hbusreq0 & v3809240 | !hbusreq0 & v376a8ee;
assign v3a6d1ce = hbusreq6 & v3750078 | !hbusreq6 & v375db7f;
assign v373b78b = hgrant6_p & v3807bf7 | !hgrant6_p & v8455ab;
assign v1e37daf = hmaster1_p & v3778ab7 | !hmaster1_p & v3a713f1;
assign v373ccc7 = hgrant6_p & v37379fc | !hgrant6_p & v3a62a8c;
assign v375c7cb = hbusreq7_p & v3a6471a | !hbusreq7_p & v3744940;
assign v3745dba = stateG10_1_p & v3741e12 | !stateG10_1_p & v375104f;
assign v373be40 = hmaster1_p & v377030a | !hmaster1_p & v3a707a1;
assign v3a57311 = jx0_p & v374c885 | !jx0_p & v3a6fc08;
assign v375bd8a = hbusreq1 & v377836a | !hbusreq1 & v37496fa;
assign v3a6f8f0 = hmaster0_p & v374e47e | !hmaster0_p & dcb1a9;
assign v377e2b3 = hmaster0_p & v374f0bf | !hmaster0_p & v374e288;
assign v3a6ec88 = hmaster1_p & v3770733 | !hmaster1_p & v373ed57;
assign v374d184 = hlock3_p & v8455ab | !hlock3_p & !v3753f1a;
assign v37708bb = hbusreq8_p & v3a637a5 | !hbusreq8_p & v372f98a;
assign v377c103 = hlock3 & v377f149 | !hlock3 & v374b424;
assign v3740fe2 = hmaster2_p & v377d1a3 | !hmaster2_p & !v3a60f71;
assign v3a5aa8e = hmaster3_p & v3a6844c | !hmaster3_p & v376b1ee;
assign v3775a25 = jx0_p & v3a6f66d | !jx0_p & v3377b02;
assign v3a66e96 = hbusreq0 & v373af1f | !hbusreq0 & v8455ab;
assign v1e37bb4 = hmaster2_p & v377234d | !hmaster2_p & !v3a70f5e;
assign v3a712b7 = hlock8 & v3753278 | !hlock8 & v3a61c73;
assign v3776d7d = hgrant6_p & v3a5e544 | !hgrant6_p & v3a70e01;
assign v3a6ec04 = hbusreq4 & v377c3a1 | !hbusreq4 & !v8455ab;
assign v3a6fb7b = hbusreq8 & v3763311 | !hbusreq8 & v3a63368;
assign v3773ee7 = hbusreq5_p & v8455ca | !hbusreq5_p & v374e0f6;
assign v3378f4e = hlock5_p & v2ff9371 | !hlock5_p & v3774937;
assign v3748234 = hmaster2_p & v372e0b0 | !hmaster2_p & v3737c0d;
assign v3779bde = hlock5 & v3a6add2 | !hlock5 & v3a712c0;
assign bdbe8b = hmaster3_p & v3a68183 | !hmaster3_p & v37766d3;
assign v37284a9 = hgrant1_p & v3a57445 | !hgrant1_p & !v376653d;
assign v374e78f = locked_p & v373d9e5 | !locked_p & !v8455ab;
assign v37482c3 = hmaster2_p & v377b429 | !hmaster2_p & !v8455ab;
assign v373c275 = hlock8_p & v3732c56 | !hlock8_p & v3a6dae0;
assign v376129a = hgrant0_p & v3a708fd | !hgrant0_p & v37777bf;
assign v3a6f3f9 = hlock6_p & v375bf9a | !hlock6_p & v8455b0;
assign v8f7302 = hmaster0_p & v376a2df | !hmaster0_p & v372c46e;
assign v374535e = hbusreq6 & v3740f7d | !hbusreq6 & v8455ab;
assign v3a70ac8 = hbusreq6 & v3a7039e | !hbusreq6 & !v8455ab;
assign v3757066 = hbusreq7_p & v377d27f | !hbusreq7_p & v376054c;
assign v3a6eb5a = hgrant3_p & v35b7299 | !hgrant3_p & !v3a5f0a7;
assign v376827d = hlock8 & v37682bc | !hlock8 & v3769bb0;
assign v3a5b978 = hgrant4_p & v3a696ed | !hgrant4_p & v1e3795b;
assign v3a5468d = hlock4_p & v37665bf | !hlock4_p & v8455e7;
assign v3728826 = hbusreq1_p & v376f56d | !hbusreq1_p & !v8455ab;
assign v3808f44 = hbusreq0 & v3741b6c | !hbusreq0 & v37477ca;
assign v37297ce = hmaster2_p & v3a64421 | !hmaster2_p & v3740d3b;
assign v3758180 = hbusreq5_p & v3a66d94 | !hbusreq5_p & v3765265;
assign v377a104 = hmaster0_p & v3a6a4e6 | !hmaster0_p & !v8455ab;
assign v3776e33 = hmaster1_p & v372f309 | !hmaster1_p & v3a5af26;
assign v373478e = hgrant5_p & v8455ab | !hgrant5_p & v377b732;
assign v325c9cb = hbusreq4_p & v372391f | !hbusreq4_p & !v375c5a8;
assign v3a70204 = hbusreq0 & v3a54393 | !hbusreq0 & v3a70b8a;
assign v3729127 = hbusreq6_p & v374bcb4 | !hbusreq6_p & v3a299d7;
assign v376158e = hlock5 & v3a6f8a9 | !hlock5 & v3a67f58;
assign v3a65069 = hmaster2_p & v3a712dd | !hmaster2_p & v373b02e;
assign cc70ad = hgrant5_p & v8455ab | !hgrant5_p & v374e538;
assign v3732b75 = hbusreq3_p & v3748665 | !hbusreq3_p & v8455ab;
assign v3723247 = hgrant0_p & v3735f14 | !hgrant0_p & v3a6f7c0;
assign v377a63c = hbusreq0_p & v373ad3c | !hbusreq0_p & v376bb26;
assign v3a70752 = hbusreq2 & v3747527 | !hbusreq2 & v377ba5a;
assign v375dd87 = hbusreq5_p & v376ecde | !hbusreq5_p & v8455ab;
assign v3730651 = hbusreq5 & ae0bd0 | !hbusreq5 & v375b0ad;
assign v374de48 = hbusreq6 & v3a713f4 | !hbusreq6 & v380730d;
assign v375b563 = hbusreq5 & v374fab7 | !hbusreq5 & v377de7f;
assign v9d7b97 = hgrant0_p & v3722e5c | !hgrant0_p & v37682a8;
assign v376b4a2 = hmaster0_p & v8455ab | !hmaster0_p & v3752987;
assign v3775442 = hbusreq1 & v3806db7 | !hbusreq1 & v374f87c;
assign v3a704eb = hlock7_p & v3a6535f | !hlock7_p & !v3a662a2;
assign v373ff5c = hmaster2_p & v37469c4 | !hmaster2_p & v3a6f781;
assign v37c0282 = hgrant5_p & v3731c27 | !hgrant5_p & v3a6f706;
assign v3a675ad = hmaster2_p & v3a6b924 | !hmaster2_p & v3735d9c;
assign v373c7a5 = hgrant6_p & v375cfa5 | !hgrant6_p & v37792cf;
assign v37536fd = hmaster0_p & v375685c | !hmaster0_p & v3737f8d;
assign v37571d0 = hbusreq8_p & bf2cd1 | !hbusreq8_p & v3751154;
assign v3a69b5f = hlock0_p & v3a635ea | !hlock0_p & v373339c;
assign v3760e78 = hlock7_p & v3a6450a | !hlock7_p & !v8455ab;
assign v3a70016 = hmaster0_p & v3a6e5f0 | !hmaster0_p & v376b856;
assign v374350d = hmaster1_p & v3a6f4f9 | !hmaster1_p & !v3a6f446;
assign v3a551bd = jx0_p & v3759aea | !jx0_p & v374cb86;
assign v375a79d = hmaster1_p & v372d249 | !hmaster1_p & v3a70601;
assign v3a6f77a = hgrant3_p & v3732128 | !hgrant3_p & v37598c6;
assign v3731a1f = hbusreq0 & v3767437 | !hbusreq0 & v373e814;
assign v377632d = hbusreq7 & v374680c | !hbusreq7 & !v37659c6;
assign v3a711e2 = hgrant6_p & v8455ab | !hgrant6_p & v3740f92;
assign v3a70311 = hlock7_p & v37656cd | !hlock7_p & !v35b70fa;
assign v377150c = hlock4 & v3757091 | !hlock4 & v372b906;
assign v3a70513 = hmaster2_p & v37326a0 | !hmaster2_p & v372e4cf;
assign v373e8b5 = hbusreq1_p & v3a6fc6c | !hbusreq1_p & v373c059;
assign v3a66b8a = hmaster1_p & v3a6fe0d | !hmaster1_p & v3a6fccc;
assign v3a5c5ae = hgrant1_p & v3a5891c | !hgrant1_p & !v3809adf;
assign v3726013 = hmaster0_p & v3a70e3f | !hmaster0_p & v3a70be7;
assign v376aaef = hmaster2_p & v3a70c8c | !hmaster2_p & v37593a1;
assign v3255a34 = hmaster0_p & v8455ab | !hmaster0_p & v3a6744e;
assign v376a411 = hbusreq5_p & v3776a59 | !hbusreq5_p & !v3a57e56;
assign v3a6f6e0 = hmaster1_p & v3a635ea | !hmaster1_p & v3a6d6fb;
assign v376c198 = hmaster2_p & v374f96e | !hmaster2_p & v8455ab;
assign v374047a = hgrant3_p & v373f42a | !hgrant3_p & v3a62037;
assign v2acb0a5 = hmaster2_p & v3747302 | !hmaster2_p & v23fd83f;
assign v376614b = hbusreq6_p & v3728498 | !hbusreq6_p & v3762c26;
assign v37571da = hgrant2_p & v3a5eadd | !hgrant2_p & v3760629;
assign v37257cf = hmaster1_p & v3a5e696 | !hmaster1_p & v3756813;
assign v375a990 = hbusreq6_p & v3766218 | !hbusreq6_p & v39eb4a7;
assign v3a6ff97 = hmaster2_p & v3a5fe5e | !hmaster2_p & v3a6ef06;
assign v37774e4 = hbusreq6 & v3a6dc08 | !hbusreq6 & v3730ffe;
assign v377e933 = hgrant6_p & v8455b5 | !hgrant6_p & v37286a2;
assign v377a901 = hbusreq6 & v3752000 | !hbusreq6 & v3a6da8a;
assign v3772d0e = hmaster1_p & v37576f6 | !hmaster1_p & v372c467;
assign v377296d = hbusreq5_p & v3727a16 | !hbusreq5_p & v3746fdb;
assign v377a2b2 = hmaster1_p & v3a60b69 | !hmaster1_p & v8455ab;
assign v373096c = hgrant4_p & v372e708 | !hgrant4_p & v8455ab;
assign v3758700 = hgrant6_p & v3733d6e | !hgrant6_p & v37728d3;
assign v37316fd = hgrant2_p & v8455ba | !hgrant2_p & v3765626;
assign v3a71285 = hmaster1_p & v375ff11 | !hmaster1_p & v3737421;
assign v3807587 = hmaster1_p & v372b29d | !hmaster1_p & v3a6fa33;
assign v3a6918e = hbusreq1_p & v3779709 | !hbusreq1_p & !v3732e39;
assign v3a71026 = hgrant4_p & v373d11f | !hgrant4_p & v3a58db9;
assign v3740625 = hbusreq0_p & v8455b6 | !hbusreq0_p & v377e928;
assign v3a69146 = hbusreq6_p & v38064a2 | !hbusreq6_p & !v8455ab;
assign v3729e05 = hbusreq2_p & v3a6f6fa | !hbusreq2_p & v372c151;
assign v3a6ff18 = hlock6 & v3a5ef6e | !hlock6 & v372fd12;
assign v3a71576 = hmaster1_p & v37757cb | !hmaster1_p & v3778657;
assign v3777f6e = hmaster2_p & v374c3f2 | !hmaster2_p & v3737d44;
assign v3742132 = hbusreq7 & v2acaff1 | !hbusreq7 & cb0c12;
assign v3729b63 = hlock3_p & v38073fd | !hlock3_p & !v8455ab;
assign v3a70a83 = stateG2_p & v3a5a496 | !stateG2_p & v3745b85;
assign v3745241 = hbusreq0 & v3a71188 | !hbusreq0 & v37501f3;
assign v3745b36 = hgrant1_p & v38072fd | !hgrant1_p & v8455ab;
assign v3738365 = hmaster0_p & v92e5bb | !hmaster0_p & v3a6607f;
assign v3a67cf0 = hmaster2_p & v3a702ee | !hmaster2_p & !v8455ab;
assign v3a55f42 = hbusreq4 & v3a70468 | !hbusreq4 & v375b92a;
assign v3768678 = hbusreq7 & v3a663dd | !hbusreq7 & v3a66f40;
assign v3a6fd10 = hbusreq5_p & v377d1dc | !hbusreq5_p & v37763d1;
assign v3a6279c = hlock5 & v3777888 | !hlock5 & v3774385;
assign v376ebc6 = hmaster2_p & v3730118 | !hmaster2_p & v3729996;
assign v373c853 = hgrant3_p & v3a55aba | !hgrant3_p & !v8455ab;
assign v377a5cc = hbusreq7_p & v374d669 | !hbusreq7_p & v3a70652;
assign v37bfc35 = hgrant4_p & v374ddcd | !hgrant4_p & v377eda6;
assign v376b0cc = hmaster1_p & v375dff6 | !hmaster1_p & v376b2f4;
assign v3a62968 = hgrant4_p & v3a6ff99 | !hgrant4_p & v3a6dcb9;
assign v372cfbf = hgrant6_p & v8455ab | !hgrant6_p & v3a621be;
assign v3a6f722 = hgrant6_p & v3760a55 | !hgrant6_p & v3a605f1;
assign v3a55673 = hgrant2_p & v376df02 | !hgrant2_p & v3758d37;
assign v3a6e622 = hgrant3_p & v3725230 | !hgrant3_p & v3a70a8a;
assign v37603af = stateG3_1_p & v8455ab | !stateG3_1_p & v845601;
assign v373a4e4 = hbusreq2_p & v377852a | !hbusreq2_p & v8455ab;
assign v3727a82 = hlock7_p & v37648fb | !hlock7_p & !v8455ab;
assign v3a6b5ea = hlock5_p & v375d889 | !hlock5_p & v3758c07;
assign v3a6faf6 = hbusreq6 & c827f4 | !hbusreq6 & v8455ab;
assign v3a60cd0 = hmaster2_p & v3a55033 | !hmaster2_p & !v3735b3e;
assign v3a6dcb2 = hlock0_p & v372b351 | !hlock0_p & v376605a;
assign v3a705d3 = hlock8_p & v3a6165e | !hlock8_p & v3725367;
assign v376da22 = hgrant4_p & v3a6f43e | !hgrant4_p & v37235bd;
assign v374473f = hgrant1_p & v37422d8 | !hgrant1_p & v8455e7;
assign v3a70265 = hmaster1_p & v3763a33 | !hmaster1_p & v373d32e;
assign v3761866 = hbusreq4 & v37274c2 | !hbusreq4 & !v8455b5;
assign v3a6b07b = hmaster2_p & v1e38224 | !hmaster2_p & !v3a695fc;
assign v3a5ade4 = hmaster2_p & v3768c3c | !hmaster2_p & v3a5fdd3;
assign v3776c6b = hbusreq8_p & v3a635ea | !hbusreq8_p & v3728e91;
assign v3a5e1a5 = hbusreq3_p & v924b19 | !hbusreq3_p & !v8455ab;
assign v3a707e0 = hmaster0_p & v3a5c3a0 | !hmaster0_p & v373e5d9;
assign v372a49a = hmaster2_p & v3a71293 | !hmaster2_p & v3a5fbd6;
assign v37354a9 = hmaster0_p & v372aacf | !hmaster0_p & v3a6f3a2;
assign a52d64 = hbusreq5_p & v373c1ff | !hbusreq5_p & v375517b;
assign v372fe05 = busreq_p & v377d219 | !busreq_p & !v376a967;
assign v3a70617 = hbusreq7_p & v3a7023d | !hbusreq7_p & v374d1ad;
assign v3a60b69 = hmaster0_p & v376e0b5 | !hmaster0_p & v8455ab;
assign v37650dd = hbusreq3_p & b66740 | !hbusreq3_p & !v2092faa;
assign v373014d = hlock3_p & v3a6ffca | !hlock3_p & !v8455ab;
assign v374db8d = hlock4_p & v3a6ffca | !hlock4_p & !v8455ab;
assign v376c573 = hmaster0_p & v3760d54 | !hmaster0_p & v3a5a52d;
assign v375367c = hlock5 & v377de7f | !hlock5 & v375b563;
assign v37247e2 = hgrant1_p & v3769f4a | !hgrant1_p & v8455ab;
assign v3a555b3 = hmaster2_p & v376618c | !hmaster2_p & v3731142;
assign v360c6f5 = hgrant1_p & v37422d8 | !hgrant1_p & v37457fb;
assign v3a6eff7 = hbusreq6_p & v3a635c3 | !hbusreq6_p & v3737acd;
assign v3a703c0 = hlock4_p & v372fba5 | !hlock4_p & v8455b0;
assign v3736217 = hlock4 & v3a552f7 | !hlock4 & cb1cc0;
assign v3a5bd99 = hgrant4_p & v8455ab | !hgrant4_p & v3757818;
assign v3a5ef54 = hready & v37386a9 | !hready & v3a635ea;
assign v377311c = hgrant8_p & v372f58a | !hgrant8_p & v3a70658;
assign v3a6b688 = hgrant2_p & v3a680b9 | !hgrant2_p & v374fcf6;
assign v3742a27 = hlock0 & v3a65d01 | !hlock0 & v37621eb;
assign v3733dea = hmaster2_p & v377395f | !hmaster2_p & v8455e7;
assign v3729c28 = hbusreq7_p & v3727651 | !hbusreq7_p & v3a70df8;
assign v374e758 = hmaster2_p & v3760954 | !hmaster2_p & v373e49f;
assign v37295e7 = hmaster2_p & v3a705c5 | !hmaster2_p & v3a70d99;
assign v37782af = hbusreq2_p & v3a70799 | !hbusreq2_p & v3a7028d;
assign v3a5fb15 = hbusreq6_p & v372defe | !hbusreq6_p & v8455e7;
assign v3756981 = hmaster0_p & v3a5e2a3 | !hmaster0_p & v3742938;
assign v37468e5 = hgrant4_p & v3a70f7a | !hgrant4_p & v8455ab;
assign hmastlock = v2619368;
assign v3a70ed3 = hbusreq5 & v878208 | !hbusreq5 & v3738b70;
assign v3a7058d = hmaster2_p & v372a4c1 | !hmaster2_p & v8455ab;
assign v372998a = hgrant6_p & v375564e | !hgrant6_p & v3a5c858;
assign v3a62027 = hmaster1_p & v376285a | !hmaster1_p & v3765927;
assign v3a64e13 = hlock8_p & v373327e | !hlock8_p & v375d23b;
assign v37545a5 = hgrant6_p & v3748194 | !hgrant6_p & !v3a6eeba;
assign v3a70472 = hmaster1_p & v3750746 | !hmaster1_p & v3769cac;
assign v3756780 = hbusreq7 & v3a2a105 | !hbusreq7 & !v3765e47;
assign v3a6f703 = hgrant5_p & v3743dc4 | !hgrant5_p & v3a70a2d;
assign v3759b6f = hbusreq6_p & v37503ec | !hbusreq6_p & !v3a63f27;
assign v37721cb = hgrant4_p & v8455ab | !hgrant4_p & v376beed;
assign v375f238 = hbusreq8_p & v3a71254 | !hbusreq8_p & v375fcac;
assign v3a70f4e = hmaster0_p & v376761d | !hmaster0_p & v37286e9;
assign v3a6fd2f = hmaster0_p & v3a62a6d | !hmaster0_p & v3775782;
assign v3731ca8 = hbusreq5_p & v3a6b924 | !hbusreq5_p & v375b7b0;
assign v3a6aea3 = hmaster0_p & v3779183 | !hmaster0_p & v3a6f901;
assign v3a6fee7 = hmaster0_p & v3a6ff93 | !hmaster0_p & v3a714d5;
assign v375da3a = hlock0_p & v3729724 | !hlock0_p & v3732aa6;
assign v375733e = hbusreq6 & v372e9f3 | !hbusreq6 & v373c2ec;
assign v37667b3 = hgrant6_p & v373a333 | !hgrant6_p & v3742521;
assign v3a7081c = hlock0_p & v3a635ea | !hlock0_p & v376c777;
assign v3a551d7 = hbusreq5_p & v3756740 | !hbusreq5_p & !v3807b2e;
assign v35ba1c6 = hmaster2_p & v8455ab | !hmaster2_p & v373c755;
assign v3738700 = hbusreq0_p & v374c693 | !hbusreq0_p & v372998c;
assign v376c0a0 = hbusreq5_p & v3741d24 | !hbusreq5_p & v3750e89;
assign v37244e7 = hgrant0_p & v8455ab | !hgrant0_p & v375323b;
assign d08a74 = hbusreq3_p & v375825a | !hbusreq3_p & v37504b9;
assign v373dceb = stateA1_p & v3a6ffe0 | !stateA1_p & v3a5cf0b;
assign v35b7299 = hbusreq3_p & v8455e7 | !hbusreq3_p & !v8455ab;
assign v372b819 = stateG10_1_p & v2aca977 | !stateG10_1_p & v376f665;
assign v37645ec = hbusreq3_p & v3a6999c | !hbusreq3_p & !v8455ab;
assign v377a10f = hmaster0_p & v3730cde | !hmaster0_p & v3737e2e;
assign v373a822 = hgrant4_p & v8455ab | !hgrant4_p & v3a656b6;
assign v37594c5 = hbusreq4_p & v3729b2e | !hbusreq4_p & !v3a70af5;
assign v3a70348 = hmaster0_p & v373632a | !hmaster0_p & b2ea29;
assign v37730b3 = hmaster1_p & v8455ab | !hmaster1_p & v3775072;
assign v377db81 = hbusreq4_p & v3a6ef34 | !hbusreq4_p & v8455ab;
assign v3a6fb1d = hbusreq5_p & v3726634 | !hbusreq5_p & v8455ab;
assign v374f36b = hmaster1_p & v3751e0a | !hmaster1_p & v373f6f0;
assign v3a64862 = hmaster0_p & v3a6604e | !hmaster0_p & !v3776b20;
assign v374a509 = hbusreq5 & v3a70467 | !hbusreq5 & v377077a;
assign v3a66349 = hmaster3_p & v376b1d4 | !hmaster3_p & v8455ab;
assign v3744d99 = hmaster2_p & v37738fc | !hmaster2_p & v8455ab;
assign v3a707ea = hbusreq6_p & v3732d82 | !hbusreq6_p & v3a69946;
assign v3730402 = hlock5 & v3a698ab | !hlock5 & v28896f0;
assign v3770338 = hgrant5_p & v37736b4 | !hgrant5_p & v3a6261c;
assign v37418b3 = hbusreq1 & v39a5265 | !hbusreq1 & !v2acb5a2;
assign v373c3ba = hbusreq0 & v374ad24 | !hbusreq0 & !v37298b9;
assign v375d453 = hbusreq0_p & v3a562a9 | !hbusreq0_p & v37674c1;
assign v374b23d = hmaster0_p & v28896dc | !hmaster0_p & v37662e7;
assign v374a134 = hlock6_p & v376d9ad | !hlock6_p & v8455e7;
assign v376e661 = hmaster2_p & v372b6bc | !hmaster2_p & v3a7058a;
assign v3738279 = hlock5_p & v376eed1 | !hlock5_p & !v8455ab;
assign v3a6b6a3 = hmaster0_p & v3a5a807 | !hmaster0_p & v3a6f56a;
assign v3769d4c = hmaster0_p & v3a6fab8 | !hmaster0_p & v37662e7;
assign v3a67de4 = hgrant6_p & v8455ca | !hgrant6_p & v3758fc7;
assign v37342cd = hmaster1_p & v375646d | !hmaster1_p & v373833b;
assign v3a5ba1a = hgrant6_p & v8455ab | !hgrant6_p & v3a66fb3;
assign v373ec24 = hlock4_p & v39a4dbb | !hlock4_p & v3736847;
assign v3a6eeb5 = hlock0_p & v3779060 | !hlock0_p & !v3a6dfb2;
assign v3775533 = hmaster0_p & v3765aee | !hmaster0_p & v3741b5e;
assign v3a57122 = hbusreq0 & d2728f | !hbusreq0 & v8455ab;
assign v3732cf6 = jx0_p & v3740777 | !jx0_p & v373ee66;
assign v3a71118 = hbusreq5 & v37384a9 | !hbusreq5 & !v3a5b955;
assign v37359cb = hlock5 & v37548e9 | !hlock5 & v3a5c4c6;
assign v375803a = hbusreq1_p & v373dcb6 | !hbusreq1_p & v3a6ffbe;
assign v373c7aa = hlock7 & v3a5dff7 | !hlock7 & v3a64200;
assign v376c3f8 = jx0_p & v376cc45 | !jx0_p & v3757e4a;
assign v37512d2 = hbusreq7_p & v3a6ecdf | !hbusreq7_p & !v377f46e;
assign v3a71473 = hlock0 & v3748797 | !hlock0 & v3a70960;
assign v3a63c8e = hmaster1_p & v377b3df | !hmaster1_p & v3774359;
assign a90ef2 = hgrant6_p & v3a6f8f6 | !hgrant6_p & v373cdb0;
assign v3760951 = hmaster2_p & v3733467 | !hmaster2_p & v375898f;
assign v3768d7e = hmaster1_p & v37444c9 | !hmaster1_p & !v3a551d7;
assign v3a6ec08 = hgrant7_p & v374ac8a | !hgrant7_p & v3778c9a;
assign v3a6d926 = hmaster1_p & v375929c | !hmaster1_p & v3728d9c;
assign v3734e69 = hlock4 & v3a701c3 | !hlock4 & v3a6fe44;
assign v3731a3b = hbusreq6 & v373d4fc | !hbusreq6 & v391331d;
assign v37522e8 = hmaster3_p & v37601df | !hmaster3_p & v3a6fe57;
assign v374d965 = hbusreq4 & v3725494 | !hbusreq4 & v37763c2;
assign v373184e = hbusreq3 & v374f76a | !hbusreq3 & v3a708c2;
assign v3734a79 = hbusreq3 & v3768ecc | !hbusreq3 & v8455e7;
assign v373f9db = hgrant6_p & v3a55efa | !hgrant6_p & v3730fc0;
assign c0d797 = hmaster1_p & v37763bd | !hmaster1_p & v3a65df3;
assign v376072e = hmaster0_p & v372883e | !hmaster0_p & v3764ed7;
assign v3a63bbc = hlock0_p & v39a5381 | !hlock0_p & v8455ab;
assign v3a542c0 = hbusreq7 & v3a6dd4d | !hbusreq7 & v375567c;
assign v37606bb = jx3_p & v3a5690f | !jx3_p & v375f883;
assign v3a7156b = hgrant5_p & aeaf7c | !hgrant5_p & v3807abe;
assign bad3a6 = hbusreq1 & v3a6ab5f | !hbusreq1 & !v2aca977;
assign v3727eda = hbusreq4 & v3773c62 | !hbusreq4 & v8455ab;
assign v372c3d7 = hmaster0_p & v373ac08 | !hmaster0_p & v377cccb;
assign v3a5e2b2 = hbusreq4 & v37756e8 | !hbusreq4 & v8455ab;
assign v3760c3d = hbusreq5_p & v3a5732f | !hbusreq5_p & v3756ea2;
assign v373fbb6 = hbusreq4_p & v377e70d | !hbusreq4_p & v3726f89;
assign v3a6c004 = hgrant4_p & v1e37b99 | !hgrant4_p & c8d28b;
assign v3a6ac81 = hbusreq3 & v39a5265 | !hbusreq3 & !v2acb5a2;
assign v3a71161 = hmaster1_p & v3724394 | !hmaster1_p & v37551b0;
assign v372abb1 = hgrant4_p & v8455ab | !hgrant4_p & v3a714bf;
assign v3a704e9 = hmaster2_p & v3a6ac26 | !hmaster2_p & v8455ab;
assign v3806f68 = hbusreq6 & v8455ab | !hbusreq6 & v8455b0;
assign v375b7b0 = hgrant4_p & v376d2b7 | !hgrant4_p & v3761d0c;
assign v37401ce = hbusreq2 & v8455b0 | !hbusreq2 & v3755791;
assign v3a70646 = hgrant5_p & v3a61b9d | !hgrant5_p & v3a7121e;
assign v3723a1d = hlock8_p & v3a7141d | !hlock8_p & !v8455ab;
assign v37781b8 = hbusreq4_p & v3a6cd35 | !hbusreq4_p & v3a712b1;
assign v3a62e92 = hbusreq5 & v376e1fd | !hbusreq5 & v37493b4;
assign v3768690 = hmaster1_p & a568f8 | !hmaster1_p & v3a6f4ce;
assign v3a70ca6 = jx2_p & v3a56114 | !jx2_p & v3807b9c;
assign v3a70950 = hmaster2_p & v37318d7 | !hmaster2_p & v3770bd5;
assign v3747971 = hmaster2_p & v3766c60 | !hmaster2_p & v37796c5;
assign v3a56a2c = hmaster2_p & v2aca977 | !hmaster2_p & v8455ab;
assign v377c71e = hmaster0_p & v3807f45 | !hmaster0_p & v376f80c;
assign v3a68426 = hbusreq1_p & v3768e48 | !hbusreq1_p & v8455ab;
assign v3774d13 = hbusreq8_p & v3735fc8 | !hbusreq8_p & !v3744202;
assign v3a70306 = jx1_p & v3a6cd89 | !jx1_p & v373c7af;
assign v374e855 = hbusreq6_p & v3a6faf6 | !hbusreq6_p & v8455ab;
assign v37537cc = hready_p & v3a5ada2 | !hready_p & v3a5a711;
assign v373e933 = hbusreq6 & v376eb3f | !hbusreq6 & v3a6f968;
assign v8f4f53 = hbusreq7_p & v3777b84 | !hbusreq7_p & v373c342;
assign v2acb5bc = jx0_p & v3a68757 | !jx0_p & v3a592bb;
assign v377f27f = hgrant0_p & v377eaf2 | !hgrant0_p & v8455ab;
assign v3a596df = hbusreq5_p & v3747aa5 | !hbusreq5_p & !v38097ae;
assign v372a599 = hmaster0_p & v3775303 | !hmaster0_p & v3a6d003;
assign v3a67899 = hmaster2_p & v374b25d | !hmaster2_p & !v8455bf;
assign v37524b2 = hmaster0_p & v3a69892 | !hmaster0_p & v375fb03;
assign v3a6e6a7 = hmaster2_p & v3a702c2 | !hmaster2_p & v3a621cb;
assign v89df94 = hbusreq8 & v3a66b8a | !hbusreq8 & !v373e924;
assign v3747b15 = hgrant4_p & v376498f | !hgrant4_p & v3a6fba6;
assign v3a70cb0 = hmaster0_p & v37755ff | !hmaster0_p & !v373cde7;
assign v3a66b6e = hbusreq8_p & v3774662 | !hbusreq8_p & !v8455ab;
assign v3a65532 = hgrant0_p & v3778ed4 | !hgrant0_p & !v8455ab;
assign v3a5b448 = hbusreq7 & v377b4b0 | !hbusreq7 & v3774452;
assign v377989c = locked_p & v8455ab | !locked_p & v3a6ffca;
assign v3743477 = hbusreq7_p & v3a6a5a8 | !hbusreq7_p & v376ea80;
assign v3775e03 = hmaster2_p & v8455ab | !hmaster2_p & v3a70ff8;
assign v3a70af6 = hmaster2_p & v3a5952d | !hmaster2_p & !v3a713c9;
assign v845603 = stateG3_1_p & v8455ab | !stateG3_1_p & !v8455ab;
assign v3a6ffec = hbusreq5_p & v3a60bfb | !hbusreq5_p & v3a692da;
assign v3a715e5 = hbusreq5 & v377f24b | !hbusreq5 & !v3a6db95;
assign v3a6f4dc = hgrant2_p & v3758472 | !hgrant2_p & v3758f6d;
assign v3a6f3a9 = hbusreq5 & v3745790 | !hbusreq5 & v3746e10;
assign v3741e68 = hbusreq6_p & v3a6e6c9 | !hbusreq6_p & v3737534;
assign v39eb536 = hbusreq6 & v372cfad | !hbusreq6 & v8455ab;
assign v23fd799 = hmaster0_p & v3a661fe | !hmaster0_p & v360d2ce;
assign d62ab4 = hbusreq8 & v3a5c2f5 | !hbusreq8 & v37437bb;
assign v3a6d140 = hmaster0_p & v3a6f443 | !hmaster0_p & v3747816;
assign v3769510 = hgrant0_p & v3724f54 | !hgrant0_p & v3a635ea;
assign v377cf71 = hbusreq5_p & v376fc80 | !hbusreq5_p & !v374deab;
assign v8455c5 = hbusreq5_p & v8455ab | !hbusreq5_p & !v8455ab;
assign v3774f35 = hgrant4_p & v3a6a295 | !hgrant4_p & v3a70dfe;
assign v3a68cec = hmaster2_p & v3a6e29c | !hmaster2_p & v3759a27;
assign v3a70f68 = hgrant4_p & v8455ab | !hgrant4_p & v3777ce4;
assign v3761ba8 = hlock0 & v373d4ff | !hlock0 & v375afc7;
assign v3761aa3 = hgrant8_p & v37580b6 | !hgrant8_p & v374ee77;
assign v3779081 = hgrant2_p & v3732d55 | !hgrant2_p & v37782af;
assign v374f92e = hmaster2_p & v375c5a8 | !hmaster2_p & v375641f;
assign v3774757 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v3a713ef;
assign v892398 = hmaster2_p & v3a70da3 | !hmaster2_p & v372ec78;
assign v372be4a = hbusreq2 & v8455ab | !hbusreq2 & v8455b0;
assign v3a65503 = hbusreq4 & v3a70ca7 | !hbusreq4 & v3a70f67;
assign v3745509 = busreq_p & v3724744 | !busreq_p & !v3727e15;
assign v3745ced = hmaster0_p & v3a53b85 | !hmaster0_p & v3a6f7bc;
assign v37349d3 = hgrant2_p & v3a6c80b | !hgrant2_p & v3a6900b;
assign v374e5ad = hmaster0_p & v374544f | !hmaster0_p & v8455ab;
assign v3770eb9 = hgrant6_p & v8455ab | !hgrant6_p & v374b1ea;
assign v37734cb = hlock7_p & v37302a2 | !hlock7_p & v8455c7;
assign v3a6274c = hbusreq5 & v3a6c4a4 | !hbusreq5 & v37654e0;
assign v3750cfd = hmaster1_p & v373f14d | !hmaster1_p & v3a5f587;
assign v37358d5 = hbusreq5_p & v3728729 | !hbusreq5_p & v3808e5b;
assign v3a61753 = hbusreq4_p & v372610a | !hbusreq4_p & v3a56f9f;
assign v3734d60 = hlock5_p & v8455ab | !hlock5_p & v372e4e1;
assign v376fddc = hlock7 & v3752215 | !hlock7 & v3743dce;
assign v3745c75 = hbusreq4 & v3743c51 | !hbusreq4 & v3a635ea;
assign v3a6ec52 = hbusreq6 & v3a71078 | !hbusreq6 & v376711c;
assign v2acadfb = hbusreq3 & v8455e1 | !hbusreq3 & v8455ab;
assign v3743a66 = hlock4_p & v3777311 | !hlock4_p & adf78a;
assign v3776f7d = hmaster1_p & v376b374 | !hmaster1_p & v3735d84;
assign v3a5a226 = hmaster2_p & v3723211 | !hmaster2_p & v377ed6c;
assign v377db66 = hbusreq5 & v37582e1 | !hbusreq5 & v3759ce2;
assign v3751f72 = hlock2 & v377c6e8 | !hlock2 & v3722b64;
assign v3a5ae7d = hbusreq0_p & v90fd44 | !hbusreq0_p & !v8455ab;
assign v374f4d4 = hmaster0_p & v3776340 | !hmaster0_p & v3752684;
assign v375d22f = hbusreq6 & v3a6f993 | !hbusreq6 & v8455ab;
assign v376e5ef = hgrant7_p & v8455c5 | !hgrant7_p & v39ed7e4;
assign v375fa66 = hmaster3_p & v8455ab | !hmaster3_p & v374f8a1;
assign v375b0cd = hmaster2_p & v37c0382 | !hmaster2_p & v8455b5;
assign v3725e0d = hmaster2_p & v37570f8 | !hmaster2_p & v3757a88;
assign v374a806 = hbusreq5 & v3a6f2d8 | !hbusreq5 & v3730b15;
assign v37730df = hmaster1_p & v3764276 | !hmaster1_p & v3a700fa;
assign v3758f17 = hbusreq7_p & v37439ef | !hbusreq7_p & v372d782;
assign v3a556f8 = hbusreq5 & v373d4d1 | !hbusreq5 & v3a6f506;
assign v3732c86 = hmaster2_p & v37386c6 | !hmaster2_p & v3a61517;
assign v37548e7 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3a7125d;
assign v37542af = hgrant2_p & v35b774b | !hgrant2_p & v377bb62;
assign v3760088 = hlock4 & v3a6ead6 | !hlock4 & v3a70d04;
assign v3a5c7a3 = hmaster2_p & v3730e7d | !hmaster2_p & v377834b;
assign v3726156 = hbusreq8 & v373d223 | !hbusreq8 & v3731cc6;
assign v376497a = hbusreq5 & v372c6c4 | !hbusreq5 & v3740825;
assign v375a766 = hbusreq6 & v372be59 | !hbusreq6 & v8455ab;
assign v3a714b2 = hlock6_p & v372fba5 | !hlock6_p & v8455b0;
assign v372d249 = hmaster0_p & v374b759 | !hmaster0_p & v3766d24;
assign v3a6f40d = hmaster2_p & v375ea85 | !hmaster2_p & v8455ab;
assign v3728392 = hmaster0_p & v375e53a | !hmaster0_p & v376a6f1;
assign v3808d74 = hmaster1_p & v377e4d8 | !hmaster1_p & v373a26b;
assign v3763a33 = hmaster0_p & v373a1d7 | !hmaster0_p & v3776c95;
assign v372b386 = hmaster1_p & v3a66aa4 | !hmaster1_p & v37381af;
assign v3a6932d = hbusreq2_p & v38088f5 | !hbusreq2_p & !v1e38224;
assign v3765ab2 = hlock4_p & v373f92e | !hlock4_p & v37307dd;
assign v372a3de = hmaster2_p & v35772b3 | !hmaster2_p & v3778b8c;
assign v3766bdf = hmaster0_p & v37621e0 | !hmaster0_p & !v374514c;
assign v9c9282 = hbusreq7_p & v375e70f | !hbusreq7_p & !v8455ab;
assign v37265b3 = stateG10_1_p & v8455ab | !stateG10_1_p & v3a635ea;
assign v3a6d09c = hbusreq4_p & v3726d1f | !hbusreq4_p & v3a6f4ed;
assign v3a6f7a5 = hbusreq3 & v376dbdf | !hbusreq3 & v8455ab;
assign v3a5e388 = hmaster1_p & v37296f5 | !hmaster1_p & v377e406;
assign v3724b94 = hbusreq8_p & v3a715e6 | !hbusreq8_p & b4f354;
assign v377d6f9 = hbusreq0 & v377623c | !hbusreq0 & v8455ab;
assign v3a70898 = hbusreq8 & v3761da2 | !hbusreq8 & v3750fa9;
assign v373e743 = hmaster1_p & v3a6feb4 | !hmaster1_p & v376046c;
assign v3a64aa2 = hmaster1_p & v3a6a045 | !hmaster1_p & v3a6a73a;
assign v37587a6 = jx2_p & v3a5e3e2 | !jx2_p & v37606bb;
assign v3a6f47d = jx0_p & v3764eff | !jx0_p & v3a6ffeb;
assign v3735c92 = hgrant6_p & v35b774b | !hgrant6_p & v3741aa1;
assign v373f4ce = hbusreq6_p & v3757d70 | !hbusreq6_p & v8455b0;
assign v3774e32 = hlock0 & v37496fa | !hlock0 & v373d8ec;
assign v3766ff7 = hbusreq6_p & v374188e | !hbusreq6_p & v8455ab;
assign v3a70786 = hmaster0_p & v23fdf1a | !hmaster0_p & v3731b41;
assign v3a69946 = hlock0_p & v3a635ea | !hlock0_p & !v377744b;
assign v372d378 = hmaster1_p & v3a68787 | !hmaster1_p & v39eb519;
assign v3a5e74c = hmaster1_p & v3a709d1 | !hmaster1_p & !v376ca02;
assign v3766d53 = hmaster0_p & v3a57f59 | !hmaster0_p & v360d1cd;
assign v375161a = stateA1_p & v37440c3 | !stateA1_p & a81487;
assign v3a7035f = hgrant6_p & v3a69ae7 | !hgrant6_p & v373d1bb;
assign v3779486 = hbusreq8_p & v377d91c | !hbusreq8_p & v374f0f1;
assign v3a70680 = jx2_p & v3a5e776 | !jx2_p & v3759664;
assign v3a68b6c = hmaster2_p & v8455ab | !hmaster2_p & v3775b81;
assign v3a701b9 = hbusreq7_p & v375eb37 | !hbusreq7_p & v3770fff;
assign v3a64722 = hbusreq0 & v3a6f3c4 | !hbusreq0 & v377222a;
assign v3a6bbe3 = hbusreq5 & v3a709fb | !hbusreq5 & v3731720;
assign v360c5d9 = hmaster2_p & v3a6f4ba | !hmaster2_p & v374e1c3;
assign v374bc97 = hbusreq5 & v373a072 | !hbusreq5 & !v8455ab;
assign v3a703cb = hbusreq5 & v3a700a3 | !hbusreq5 & bb70de;
assign v3766b95 = hgrant4_p & v3a69ed9 | !hgrant4_p & v372610a;
assign v37350b2 = hbusreq5_p & v3807474 | !hbusreq5_p & !v3a5c188;
assign v3a6cd8b = hmaster2_p & v8455b0 | !hmaster2_p & v376d374;
assign v3746825 = hmaster1_p & v37753dc | !hmaster1_p & v374bac7;
assign v376f07c = hlock5_p & v8455ab | !hlock5_p & v372c8d0;
assign v38088f5 = hlock2_p & v1e38275 | !hlock2_p & v39a537f;
assign v373531a = hbusreq7_p & v3722b5c | !hbusreq7_p & v376beb3;
assign v373b03b = hmaster2_p & v377cfd9 | !hmaster2_p & v3a6febd;
assign v3762eeb = hmaster0_p & v3766c5c | !hmaster0_p & v372acd0;
assign v37644ff = hmaster0_p & v3a63a21 | !hmaster0_p & v3a6230b;
assign v3a6f1c1 = hbusreq5_p & v3a57ce9 | !hbusreq5_p & v3a6eee8;
assign v3734bd2 = hmaster2_p & v37745c3 | !hmaster2_p & v2ff937f;
assign v3a6fa64 = hbusreq3 & v3761af1 | !hbusreq3 & v8455ab;
assign v377ca49 = hbusreq0 & v3a6ff8f | !hbusreq0 & v377a3ec;
assign v375da82 = hbusreq2_p & v3747302 | !hbusreq2_p & v37496fa;
assign v375b18e = hgrant6_p & v3a7099b | !hgrant6_p & v8455ab;
assign v3771b63 = hmaster2_p & v374502e | !hmaster2_p & v37482f8;
assign v8e6c5f = hbusreq4 & v3a70480 | !hbusreq4 & v3a5fc82;
assign v37782c9 = hbusreq0 & v3a682b1 | !hbusreq0 & v8455b0;
assign v374d12f = hbusreq8 & v3739ed3 | !hbusreq8 & v37258d0;
assign v3a7157f = hbusreq8_p & v1e37b48 | !hbusreq8_p & v3a62a6d;
assign v3a71195 = hgrant4_p & v8455c1 | !hgrant4_p & v3a6e3e0;
assign v3a70186 = hbusreq6 & v3a6f9a2 | !hbusreq6 & v3755a05;
assign v35b91ba = hbusreq7 & v3737517 | !hbusreq7 & !v3773ee7;
assign v372cda0 = hbusreq6 & v3a58da1 | !hbusreq6 & v8455ab;
assign v3a71548 = hbusreq3_p & v3a710bc | !hbusreq3_p & v3741850;
assign v3a6fa70 = hmaster1_p & v375067d | !hmaster1_p & v372dfba;
assign v3809259 = hgrant2_p & v3a5c700 | !hgrant2_p & v376942f;
assign v38098b0 = hgrant5_p & v375d98c | !hgrant5_p & v373c239;
assign v37441fb = hmaster2_p & v3a5af94 | !hmaster2_p & v376d856;
assign v3a63329 = hbusreq2_p & v3a565eb | !hbusreq2_p & v8455ab;
assign v3a70962 = hbusreq8 & v3a62cf3 | !hbusreq8 & v8455ab;
assign v372dc77 = hbusreq7_p & v374b00b | !hbusreq7_p & v376f92c;
assign v37796c3 = hmaster0_p & v3a6f7c5 | !hmaster0_p & !v376ff85;
assign v3a6f22f = hgrant3_p & v9aa8f3 | !hgrant3_p & v3806912;
assign v3774bdf = hmaster2_p & v374ba05 | !hmaster2_p & v375c98d;
assign v3a61532 = hbusreq5_p & v37566c9 | !hbusreq5_p & !v3770a6d;
assign v37749f0 = hlock1_p & v3773df0 | !hlock1_p & v374668d;
assign v3a655cb = hlock0_p & v8455b6 | !hlock0_p & v3740625;
assign d8fb57 = hbusreq5 & v3740d4e | !hbusreq5 & v3758eb3;
assign v3745158 = hbusreq2 & v37566b2 | !hbusreq2 & v8455ab;
assign v376c5b2 = hmaster0_p & v37682fc | !hmaster0_p & v374d339;
assign v374815b = hbusreq6 & v3a712de | !hbusreq6 & v3a6006c;
assign v3773ca9 = hburst1 & v376c211 | !hburst1 & v374de7f;
assign v373ab60 = hmaster1_p & v374decf | !hmaster1_p & v37750e4;
assign v3759628 = hbusreq7_p & v377209d | !hbusreq7_p & !v3764378;
assign v3a5e0dd = jx0_p & v3773536 | !jx0_p & !v375f689;
assign v3725ec4 = hgrant6_p & v8455ab | !hgrant6_p & v3a6f243;
assign v3757b9b = hbusreq6_p & v9015e2 | !hbusreq6_p & v8455ab;
assign v372c85f = hmaster0_p & v3a635ea | !hmaster0_p & v3a5e620;
assign v376b0f2 = hgrant4_p & v37402cd | !hgrant4_p & v8455ab;
assign v3762642 = hmaster0_p & v3734c5c | !hmaster0_p & v3577392;
assign v9b81ab = hmaster0_p & v3a5e24e | !hmaster0_p & v1e37784;
assign v3a6fc90 = hbusreq6 & v3764a94 | !hbusreq6 & v8455ab;
assign v3727638 = hbusreq0_p & v3a6fe1a | !hbusreq0_p & v37c0382;
assign v375dd4c = hbusreq8 & v3a664e6 | !hbusreq8 & v3756a20;
assign v38072f0 = hmaster0_p & v8455e7 | !hmaster0_p & v3757569;
assign v373705f = hlock7_p & v3577388 | !hlock7_p & v376c94b;
assign v3755901 = hbusreq8 & v3779cda | !hbusreq8 & v3737808;
assign v372a3dc = hmaster3_p & v3a59f5a | !hmaster3_p & v3724a10;
assign v373d5e7 = hmaster0_p & v37570f8 | !hmaster0_p & v3a5c75a;
assign v3a6efe3 = hbusreq6_p & v376b651 | !hbusreq6_p & !v8455ab;
assign v377e618 = hbusreq4_p & v1e37846 | !hbusreq4_p & v3a65716;
assign v376c1e4 = hlock4 & v3a70d0f | !hlock4 & v375f6ef;
assign v3777b00 = hgrant4_p & v3758aec | !hgrant4_p & v3a57db8;
assign v3768c97 = hmaster2_p & v372b780 | !hmaster2_p & v3723a00;
assign v3a6f4e0 = hbusreq7_p & v3750797 | !hbusreq7_p & v3a63fd5;
assign v3a62092 = hmaster2_p & v3a712e2 | !hmaster2_p & v9bf1d8;
assign v376f9eb = hbusreq4 & v3768ecc | !hbusreq4 & v8455ab;
assign v375c67c = hmaster1_p & v39ea76e | !hmaster1_p & v377c490;
assign v3a68255 = hlock6 & v3a711fa | !hlock6 & v377b4b9;
assign v3a6bbee = hgrant2_p & v3a71121 | !hgrant2_p & v23fe10d;
assign v3761cdb = hbusreq0 & v377defb | !hbusreq0 & v375cd00;
assign v3723db5 = hlock7 & v3a69391 | !hlock7 & v375ceb9;
assign v3735f03 = hbusreq7_p & v3723a1d | !hbusreq7_p & v37550ac;
assign v3769ecf = hbusreq0 & v3738e63 | !hbusreq0 & v37765a3;
assign v377e889 = hgrant4_p & v372b8eb | !hgrant4_p & v373690a;
assign v3a6f28a = hbusreq5 & v3a6934e | !hbusreq5 & v3a7126e;
assign v373bd76 = hbusreq0 & v374733b | !hbusreq0 & v3a6eba0;
assign v37243dc = hgrant6_p & v3a6ef4c | !hgrant6_p & !v37607d2;
assign v3a6866f = hgrant4_p & v376a6f1 | !hgrant4_p & v3a6ebc3;
assign v377ef4a = hbusreq3_p & v3a6de8c | !hbusreq3_p & v3755381;
assign v375d366 = hmaster3_p & v8455ab | !hmaster3_p & v3a67beb;
assign v3745539 = hbusreq6_p & v9f9402 | !hbusreq6_p & v8455bb;
assign v2acb5a7 = hbusreq3 & v374d85e | !hbusreq3 & !v8455ab;
assign v374f0a4 = hbusreq3_p & v3a6efd1 | !hbusreq3_p & v3776c9a;
assign v372a520 = hmaster2_p & v3760eb3 | !hmaster2_p & v3a5bb6a;
assign v3731b60 = hbusreq4 & v3a70112 | !hbusreq4 & !v8455ab;
assign v3a6bc9a = hmaster2_p & v377abd6 | !hmaster2_p & v3a6fdc9;
assign v3736f36 = hmaster0_p & v3743ff2 | !hmaster0_p & v375f84b;
assign v374b3af = hgrant4_p & v8455ab | !hgrant4_p & v37717ac;
assign v3a6e152 = hbusreq8 & v374608b | !hbusreq8 & v3753838;
assign v3769de7 = hgrant3_p & v3a68aa8 | !hgrant3_p & v38079ff;
assign v3724703 = hmaster2_p & v8455ab | !hmaster2_p & bb97e8;
assign v2acb5c7 = hmaster2_p & v3740161 | !hmaster2_p & v374f501;
assign v3a5ea57 = hmaster1_p & v3a6f662 | !hmaster1_p & v373b130;
assign v1e38283 = hmaster0_p & v37649c2 | !hmaster0_p & v3a7000a;
assign v3775abc = hgrant0_p & v3770559 | !hgrant0_p & c1a4f5;
assign v2e5fb38 = hbusreq5 & v3734502 | !hbusreq5 & v37476b8;
assign v3a6f441 = hmaster2_p & v8455ab | !hmaster2_p & !v3750d37;
assign v3775f0b = hmaster2_p & v3757966 | !hmaster2_p & v3a70bf2;
assign v3a62fc6 = hmaster2_p & v377caa3 | !hmaster2_p & v3a6f8f5;
assign v373b4aa = hmaster2_p & v3a5ace5 | !hmaster2_p & v373e8ad;
assign v3a679e7 = hbusreq4 & v37775f9 | !hbusreq4 & v3a635ea;
assign v373bcb6 = hgrant4_p & v8455ab | !hgrant4_p & v3746259;
assign v37507d0 = hbusreq3_p & v3753f1a | !hbusreq3_p & !v8455ab;
assign v3762729 = hlock8_p & v3a56118 | !hlock8_p & v376bfe6;
assign v375cab5 = hmaster0_p & v372efb1 | !hmaster0_p & v375f78f;
assign v377938d = hbusreq6_p & v3a6ae2d | !hbusreq6_p & v3a708a2;
assign v3a6fbf6 = hlock7 & v3734279 | !hlock7 & v37484b6;
assign v37359d8 = hgrant0_p & v1e3791d | !hgrant0_p & v39eaa47;
assign v37655ac = hbusreq2_p & v377ab2c | !hbusreq2_p & v3a6fcef;
assign v3a6d21e = hgrant4_p & v3777d29 | !hgrant4_p & !v3a5c0ac;
assign v3a70556 = hmaster0_p & v374e0f6 | !hmaster0_p & v374e4ec;
assign v3767a5b = hgrant3_p & v35b7299 | !hgrant3_p & v3a71688;
assign v3765305 = hbusreq4_p & v3736f61 | !hbusreq4_p & v376de99;
assign v377f21b = hbusreq6_p & v372c83f | !hbusreq6_p & v3743546;
assign v3738e63 = hlock4 & v3a7165c | !hlock4 & v376beb4;
assign v372defe = hlock6_p & v3778ed4 | !hlock6_p & v8455e7;
assign v3751081 = hbusreq0 & v374d2e5 | !hbusreq0 & v374b6ac;
assign v3a6f9bd = hmaster2_p & v8455ab | !hmaster2_p & v375d84e;
assign v376954d = hgrant4_p & v8455ab | !hgrant4_p & v373262e;
assign v3a70816 = hbusreq7_p & v3776081 | !hbusreq7_p & !v3776f25;
assign v3734634 = hgrant4_p & v3a53eeb | !hgrant4_p & v3722a7e;
assign v376d935 = hbusreq4 & v37425ad | !hbusreq4 & v1e38288;
assign v3a538ba = hbusreq5_p & v375c01e | !hbusreq5_p & v374457a;
assign v3a620fd = hlock8_p & v376c477 | !hlock8_p & v3a6ebc6;
assign v37531ca = hbusreq7_p & v3734279 | !hbusreq7_p & v376d23f;
assign v3a705f2 = hbusreq0 & v375d9f8 | !hbusreq0 & v8455ab;
assign v3a709ec = hlock0 & v376e041 | !hlock0 & v3a70a03;
assign v372adfd = hmaster2_p & v37390ce | !hmaster2_p & v3732359;
assign v3737c2f = hbusreq0_p & v3a70f6a | !hbusreq0_p & v8455ab;
assign v3729381 = hmaster0_p & v3761719 | !hmaster0_p & v3751c73;
assign v374677a = hmaster2_p & c51aa0 | !hmaster2_p & v3a70bd6;
assign v3735ac0 = hbusreq5 & v3755691 | !hbusreq5 & v37366d5;
assign v3773071 = jx1_p & v377a68a | !jx1_p & v8455ab;
assign v3a6ff3f = hgrant3_p & v3a66f83 | !hgrant3_p & v3770f3a;
assign v377c6dc = hgrant4_p & v375562a | !hgrant4_p & v376681a;
assign v3a71647 = hlock0_p & v376ef42 | !hlock0_p & v37307de;
assign v374ecf9 = hgrant5_p & v3765203 | !hgrant5_p & v376ecae;
assign v373b779 = hgrant4_p & v8455ab | !hgrant4_p & v377463a;
assign v3a620f1 = hgrant4_p & v8455ab | !hgrant4_p & v372ab8f;
assign v374802b = hbusreq7 & v3733239 | !hbusreq7 & v8455ab;
assign v3a70b50 = hmaster1_p & v375620b | !hmaster1_p & v376f051;
assign v37271ad = hmaster1_p & v3757d76 | !hmaster1_p & v3a6f33e;
assign v375c55a = hbusreq2_p & v37318da | !hbusreq2_p & v3a5de50;
assign v377340e = hbusreq2_p & v372ad1d | !hbusreq2_p & v8455ab;
assign v3a6d040 = hmaster2_p & v372b231 | !hmaster2_p & v3737d38;
assign v3a6f837 = hbusreq0 & v3748ca3 | !hbusreq0 & v373006f;
assign v3728646 = hmaster2_p & v35772a6 | !hmaster2_p & v3a642cf;
assign v380662a = hburst1 & v8455ab | !hburst1 & v3779b03;
assign v3a6f882 = hbusreq3 & b0c091 | !hbusreq3 & !v3768ac7;
assign v3a6d768 = hmaster2_p & v3a56cdb | !hmaster2_p & !v3a627cc;
assign v376f032 = hmaster3_p & v374510a | !hmaster3_p & v8455ab;
assign v3a5a34e = hgrant2_p & v8455ab | !hgrant2_p & v3a70a08;
assign v374f252 = hbusreq7_p & v377a525 | !hbusreq7_p & v374ca2e;
assign v372e92b = hbusreq3_p & v3759b9a | !hbusreq3_p & v3a6eb01;
assign v373b197 = hgrant0_p & v37490cb | !hgrant0_p & v3a6b18a;
assign v3a6f0d3 = hgrant6_p & v3760e2e | !hgrant6_p & v3758824;
assign v8ef654 = hbusreq2_p & v377eaf2 | !hbusreq2_p & v372e38f;
assign v372d397 = hbusreq6 & v3731e7b | !hbusreq6 & v8455ab;
assign v375ace5 = hmaster2_p & v8455e7 | !hmaster2_p & d99853;
assign v3777817 = hmaster2_p & v374b887 | !hmaster2_p & v3728f25;
assign v3a611be = hgrant6_p & v8455ab | !hgrant6_p & v374b4da;
assign v3a67d4f = hmaster1_p & v3a714f6 | !hmaster1_p & v37418db;
assign v360c3cc = hbusreq7_p & v372f8af | !hbusreq7_p & v3765d27;
assign v2092ba8 = hbusreq6_p & v3742aff | !hbusreq6_p & !v1e38224;
assign v376fd85 = hmaster0_p & v3775dbc | !hmaster0_p & v3a6fe3f;
assign v37719f2 = hlock2 & v3258db3 | !hlock2 & v3750866;
assign v37770ab = hmaster1_p & v375398e | !hmaster1_p & v374c8b8;
assign v3a70c3a = hgrant6_p & v3a70fa7 | !hgrant6_p & v3742657;
assign v3751a0d = hmaster1_p & v372d8e8 | !hmaster1_p & v3735cfb;
assign v37795eb = hbusreq8 & v3a703c9 | !hbusreq8 & v8455ab;
assign v3751891 = hmaster2_p & v3752fe6 | !hmaster2_p & v3775537;
assign v3755e61 = hmaster0_p & v3a64421 | !hmaster0_p & v374581a;
assign v3a6f49f = hmaster2_p & v3726c61 | !hmaster2_p & v3a6fa93;
assign v3754f6b = hlock4_p & v374f87c | !hlock4_p & v377ba55;
assign v37692c1 = hbusreq0 & v37239ed | !hbusreq0 & v3736e06;
assign v376773a = hbusreq0_p & v39a4e5f | !hbusreq0_p & v3a68d2e;
assign v3a57f04 = hlock7 & v3732b30 | !hlock7 & v3753b70;
assign v3a588a0 = hbusreq0 & v3a70353 | !hbusreq0 & v3a5de18;
assign v374410c = hgrant5_p & v3a6f069 | !hgrant5_p & v3776d72;
assign v372a732 = hbusreq0_p & v376f56d | !hbusreq0_p & !v8455ab;
assign v3a583ee = hgrant2_p & v37672a5 | !hgrant2_p & v3758972;
assign v37530cf = hmaster3_p & v8455ab | !hmaster3_p & v3a673d9;
assign v37341ff = hlock7_p & v3a61992 | !hlock7_p & v3a6f44a;
assign v375ae3d = hlock8 & v3257687 | !hlock8 & v373f3e4;
assign v373e225 = hbusreq7_p & v1e37a9d | !hbusreq7_p & v372b6b9;
assign v3a6f910 = hgrant4_p & v8455ab | !hgrant4_p & v372408b;
assign v3a701b1 = hbusreq5 & v2ff918d | !hbusreq5 & v377de7f;
assign v3a71391 = hbusreq3 & v376b4e1 | !hbusreq3 & !v8455ab;
assign v3808d47 = hmaster2_p & v3a6c23b | !hmaster2_p & v8455ab;
assign v1e37558 = hlock0 & v3a5aacb | !hlock0 & v3739e7a;
assign v3a706f1 = hbusreq6_p & v3a6a489 | !hbusreq6_p & v8455bf;
assign v3a68bdb = hbusreq5 & v376c5de | !hbusreq5 & v92c996;
assign v3a569dd = hmaster1_p & v3753eb2 | !hmaster1_p & v373098e;
assign v3778e71 = hgrant6_p & v37304b3 | !hgrant6_p & v375db62;
assign v3765351 = hbusreq2_p & v3779227 | !hbusreq2_p & v377ab2c;
assign v3761ca9 = hbusreq0 & v375d0ed | !hbusreq0 & !v1e37cd6;
assign v3a6f6b9 = hbusreq4 & v3a6672b | !hbusreq4 & v8455ab;
assign v3756fd9 = hbusreq8_p & v3a6becc | !hbusreq8_p & v8455ab;
assign v3758ff0 = hmaster2_p & v3771a11 | !hmaster2_p & v3724e30;
assign v3a7161a = hmaster0_p & v3a700e0 | !hmaster0_p & v374c5c5;
assign v3740d36 = hbusreq1_p & b33e26 | !hbusreq1_p & v3a6fcd1;
assign v3a6843e = jx0_p & v3a6f860 | !jx0_p & v3740dc8;
assign v377dfbf = hmaster2_p & v3a58057 | !hmaster2_p & v3737d38;
assign v3a61344 = hbusreq4 & v3a714be | !hbusreq4 & v3a70d32;
assign v375805a = hbusreq4_p & v372c8bc | !hbusreq4_p & !v8455ab;
assign v3779a06 = hmaster2_p & v3a70f5e | !hmaster2_p & !v375f61e;
assign v3768d3e = hbusreq6 & v373399e | !hbusreq6 & v8455ab;
assign v3724e64 = hmaster0_p & v3779627 | !hmaster0_p & v373d67c;
assign v3a5d2d3 = hbusreq4_p & v37293d5 | !hbusreq4_p & v375f74e;
assign v37721eb = hbusreq2_p & v38072fd | !hbusreq2_p & v3a615bb;
assign v3723e15 = hmaster2_p & v3762929 | !hmaster2_p & v37745c3;
assign v3744637 = hbusreq4_p & v373ce49 | !hbusreq4_p & !v3a64349;
assign v3a71563 = hbusreq6_p & v3755bbd | !hbusreq6_p & v8455ab;
assign v37343e7 = hmaster0_p & v373a4ea | !hmaster0_p & v3a6ff47;
assign v375d616 = hlock2_p & v3a5d5d3 | !hlock2_p & !v8455ab;
assign v3a70d2a = hbusreq5 & v3770a5a | !hbusreq5 & v372a465;
assign v377a57a = hmaster1_p & v3a6fcfa | !hmaster1_p & v3a68dab;
assign v3a6d6fb = hmaster0_p & v3a635ea | !hmaster0_p & v375c19b;
assign v3770f75 = hgrant4_p & v3745e72 | !hgrant4_p & v377070e;
assign v3724718 = hmaster1_p & v3a56027 | !hmaster1_p & v3a6fd9f;
assign v3a7117c = hmaster2_p & v8455ab | !hmaster2_p & v37314fa;
assign v3a7098c = locked_p & v3a6a539 | !locked_p & v8455ab;
assign v3a66645 = hmaster0_p & v374502e | !hmaster0_p & v37407cb;
assign v376baad = jx0_p & v375a251 | !jx0_p & v3725c95;
assign v3a6f0a2 = hlock6 & v3a71582 | !hlock6 & v3a62d59;
assign v3725612 = hmaster0_p & v373a85c | !hmaster0_p & v8455ab;
assign v37c0297 = hbusreq2 & v3a57309 | !hbusreq2 & v8455ab;
assign v375fa82 = hlock1_p & v8455ab | !hlock1_p & !v3753f1a;
assign v3a6f5f9 = hgrant5_p & v372a264 | !hgrant5_p & v375bb06;
assign v3772775 = hmaster2_p & v2678bee | !hmaster2_p & v3a6d93d;
assign v373a984 = hgrant3_p & v3759512 | !hgrant3_p & !v374efee;
assign v3a6eb3d = hmaster0_p & v374bfcf | !hmaster0_p & v3770bcd;
assign v3753eb3 = hbusreq4_p & v3746683 | !hbusreq4_p & v360be60;
assign v372e263 = hmaster0_p & v9af7ec | !hmaster0_p & v3a71486;
assign v3377b02 = hbusreq7_p & v377aecd | !hbusreq7_p & v37491af;
assign v3a59e1b = hbusreq7_p & v373705f | !hbusreq7_p & v8455ab;
assign v373908c = hmaster2_p & v380974c | !hmaster2_p & v3767437;
assign v375a878 = hmaster0_p & v3a6ff25 | !hmaster0_p & v37333a4;
assign v3744bed = hlock5_p & v3a54b5d | !hlock5_p & !v8455ab;
assign v373178e = hgrant1_p & v3755791 | !hgrant1_p & v37328bf;
assign v3a6a48e = hbusreq0 & v380974c | !hbusreq0 & v373e814;
assign v37556c0 = hbusreq8 & v374d162 | !hbusreq8 & !v3a7022a;
assign v3a296d8 = hmaster2_p & v1e378ea | !hmaster2_p & v3751cd1;
assign v3a6fe9a = hmaster2_p & v3a57046 | !hmaster2_p & v3769740;
assign v3738f30 = hmaster0_p & v37392ae | !hmaster0_p & v23fe28c;
assign v3a5bd83 = hgrant4_p & v8455ab | !hgrant4_p & v3734d8a;
assign v373b51b = hbusreq4 & v3a704b0 | !hbusreq4 & v3a7162d;
assign v3765443 = hmaster3_p & v8455ab | !hmaster3_p & v3a708bc;
assign v3a564d9 = hmaster0_p & v3758d2a | !hmaster0_p & b05db7;
assign v3728b9d = stateG10_1_p & v35772a5 | !stateG10_1_p & !v375be5b;
assign v3a70d9c = hbusreq6_p & v376348c | !hbusreq6_p & !v8455ab;
assign v37759a7 = hmaster0_p & v3a635ea | !hmaster0_p & v3774d86;
assign v37305e3 = hgrant5_p & v3754107 | !hgrant5_p & v3750cfd;
assign v3a56cfd = hmaster0_p & v3768873 | !hmaster0_p & v3774878;
assign v37489a0 = hmaster2_p & v3a5af94 | !hmaster2_p & v39a537f;
assign v375ee43 = hbusreq5 & v372e332 | !hbusreq5 & v8455ab;
assign v3a557ea = hbusreq4 & v8907fb | !hbusreq4 & v8455ab;
assign v37435fd = hmaster0_p & v3a6fa22 | !hmaster0_p & v372b7a3;
assign v3732871 = hmaster0_p & v38097ee | !hmaster0_p & v3a715c5;
assign v3772112 = hgrant5_p & v8455ab | !hgrant5_p & v37796bf;
assign v3a6f736 = hmaster2_p & v3779183 | !hmaster2_p & v3a71678;
assign v3a647df = hbusreq4_p & v3a6f192 | !hbusreq4_p & !v8455c2;
assign v3a7154f = hbusreq0 & v8455b0 | !hbusreq0 & v3a6556a;
assign v372b3f6 = hmaster2_p & v37428ac | !hmaster2_p & v3a62aef;
assign v375583c = hbusreq8 & v3a58e79 | !hbusreq8 & v373c7af;
assign v2ff9189 = hmaster1_p & v3a68f5f | !hmaster1_p & v375eba9;
assign v37419bc = hgrant4_p & v3a5ee62 | !hgrant4_p & v37741ca;
assign v39ea76e = hbusreq2_p & v3a5c945 | !hbusreq2_p & v3a57f59;
assign v37649d3 = hbusreq6 & v3a646fb | !hbusreq6 & v372348c;
assign v376dafa = hmaster2_p & v37536ae | !hmaster2_p & !v3a7136e;
assign v3771a0d = hgrant4_p & v3a53eeb | !hgrant4_p & v374da7f;
assign v3a561f0 = hmaster1_p & v37642e6 | !hmaster1_p & !v377cb41;
assign v3a6f541 = hgrant4_p & v376a6f1 | !hgrant4_p & v3a7076d;
assign v3770ccf = hbusreq3_p & v3a5ebde | !hbusreq3_p & v3a637dd;
assign v3754dd0 = hbusreq4_p & v3809d49 | !hbusreq4_p & v8455ab;
assign v3a708d3 = hbusreq4_p & v373ac50 | !hbusreq4_p & v3734bf8;
assign v374e542 = hbusreq6 & v377359f | !hbusreq6 & v8455ab;
assign v3255b23 = hbusreq4_p & v3755ec0 | !hbusreq4_p & v3a7146b;
assign v3778a97 = hlock5_p & v8455ab | !hlock5_p & v372834d;
assign v375750d = hmaster0_p & v3a62a6d | !hmaster0_p & v372879d;
assign v373141b = hbusreq4_p & v8455ab | !hbusreq4_p & v377aa06;
assign v3774175 = hlock6_p & v8f695f | !hlock6_p & !v8455ab;
assign v3762934 = hbusreq2_p & v37538e4 | !hbusreq2_p & v37331ef;
assign v372862a = hmaster2_p & v373cbf9 | !hmaster2_p & v8455ab;
assign v3a6fcab = hmaster2_p & v3a6074d | !hmaster2_p & v3725230;
assign v3754b58 = hbusreq4_p & v3a5c7a8 | !hbusreq4_p & v35772a6;
assign v377410f = hmaster0_p & v377b24b | !hmaster0_p & v3775c03;
assign v374da8a = hmaster0_p & v3a5b6ac | !hmaster0_p & v377b556;
assign v3a63812 = hbusreq5_p & v3a70616 | !hbusreq5_p & v3a70fa8;
assign v375200e = hlock4 & v3744ae4 | !hlock4 & v3a5408c;
assign v3740d9a = hbusreq5 & v3740975 | !hbusreq5 & v3a2a107;
assign v37311d8 = hbusreq4_p & v3a71467 | !hbusreq4_p & !v376cdf6;
assign v3739b17 = hbusreq3 & v3a6772f | !hbusreq3 & v3728fb5;
assign v3727df1 = hbusreq0 & v3a63a46 | !hbusreq0 & v375ab99;
assign v37708f1 = hlock3_p & v3a55039 | !hlock3_p & v37740e0;
assign v3a6fce6 = hlock6_p & v8455e7 | !hlock6_p & !v8455ab;
assign v377375f = hbusreq7 & v3a700be | !hbusreq7 & v3773f27;
assign v3753bb2 = hbusreq6_p & v3747302 | !hbusreq6_p & v3726e81;
assign v3751b42 = hgrant6_p & v8455ab | !hgrant6_p & v3a6c0fb;
assign v3a5b310 = hmaster0_p & v3745bdf | !hmaster0_p & v3a6fb52;
assign v374457b = hmaster1_p & v8455ab | !hmaster1_p & v3a6f12b;
assign v3a6ef7f = hmaster2_p & v3725580 | !hmaster2_p & v377317d;
assign v374f272 = hbusreq7 & v3755bb4 | !hbusreq7 & v376002d;
assign v3a56027 = hbusreq5_p & v37566c9 | !hbusreq5_p & !v374fd32;
assign v3773ccd = hmaster1_p & v376c0c8 | !hmaster1_p & v3773ab1;
assign v3a6f7d5 = hbusreq7 & v375d997 | !hbusreq7 & v3a71146;
assign v373ff91 = hbusreq4_p & v3a5c945 | !hbusreq4_p & !v3a619c0;
assign v373623d = hbusreq5 & v3766101 | !hbusreq5 & v3769023;
assign v37297c0 = hmaster0_p & v3a5c945 | !hmaster0_p & v3a6cfc5;
assign v374e00b = hlock8 & v3a5cf57 | !hlock8 & v373a0f8;
assign v380853c = hbusreq1_p & v376b0fb | !hbusreq1_p & v3a70bbc;
assign v3771fd8 = hbusreq4_p & v37706fd | !hbusreq4_p & v373d735;
assign v3a64f9b = hbusreq3_p & v3772d27 | !hbusreq3_p & v374720c;
assign v376140e = hbusreq5 & v372945c | !hbusreq5 & v3a5749e;
assign v3a711f9 = hgrant4_p & v3a5cfac | !hgrant4_p & v3a6fedc;
assign v3a6f337 = hgrant8_p & v3a6aea2 | !hgrant8_p & v3a6ec08;
assign v374d810 = hbusreq4_p & v3755bb0 | !hbusreq4_p & !v8455c2;
assign v3a7109b = hbusreq8_p & v37240c0 | !hbusreq8_p & v3a70da8;
assign v3735050 = hmaster0_p & v3a70fd5 | !hmaster0_p & v3a61ab0;
assign v3730dea = stateA1_p & v3a67241 | !stateA1_p & v3a6a939;
assign v373a263 = hmaster0_p & v37710d4 | !hmaster0_p & v3a71251;
assign v3753186 = hgrant0_p & v376a2ea | !hgrant0_p & v3a6fd57;
assign v376e0df = hgrant6_p & v8455ab | !hgrant6_p & v376bb7b;
assign v372912f = hbusreq0 & v3744a60 | !hbusreq0 & v374061b;
assign v373a692 = hmaster0_p & v377adf5 | !hmaster0_p & !v376f6e4;
assign v375d113 = hbusreq7 & v3730ae6 | !hbusreq7 & v372eb5b;
assign v3739517 = hmaster2_p & v3a71416 | !hmaster2_p & v3775bd3;
assign v3a539bb = hlock6 & v37540e7 | !hlock6 & v3773b7b;
assign v3763cef = hmaster0_p & v376e31a | !hmaster0_p & !d26e1e;
assign v375d304 = hlock3_p & v37317ba | !hlock3_p & v8455e7;
assign v3756bde = hmaster0_p & v377766c | !hmaster0_p & v3a70bcd;
assign v3a65596 = hlock0_p & v3775303 | !hlock0_p & v8455b0;
assign v3a6eb26 = hmaster2_p & v372580e | !hmaster2_p & v3734827;
assign v3a6fbee = hlock5_p & v8455ab | !hlock5_p & v3771ce2;
assign b62916 = hgrant2_p & v377d770 | !hgrant2_p & v373edc8;
assign v373173e = hbusreq4 & adf78a | !hbusreq4 & v8455ab;
assign v3a708f7 = hbusreq5 & v37563cf | !hbusreq5 & v8455ab;
assign v377f424 = hmaster2_p & v3759119 | !hmaster2_p & !v8455ab;
assign v373055c = hbusreq6_p & v3a6fc90 | !hbusreq6_p & v8455ab;
assign v374a5a9 = hlock1_p & v37547c9 | !hlock1_p & !v8455ab;
assign v3745704 = hmaster2_p & v376f29d | !hmaster2_p & !v3747d37;
assign v377535e = hmaster0_p & v3a6c9c2 | !hmaster0_p & v377306c;
assign v3a64b87 = hmaster1_p & v377ed25 | !hmaster1_p & v3a6b90e;
assign v373dbb0 = hbusreq2_p & v3a6a233 | !hbusreq2_p & v23fda6a;
assign v372f292 = hbusreq3_p & v3a54344 | !hbusreq3_p & v3a640c5;
assign v374b6e8 = hmaster2_p & v8455ab | !hmaster2_p & v3730695;
assign v377050f = hmaster0_p & v3739d23 | !hmaster0_p & v3a6f7bc;
assign v3a70137 = hmaster2_p & v3a70209 | !hmaster2_p & v3a58d22;
assign v3a6ed2b = hmaster0_p & v372838e | !hmaster0_p & v3748b9d;
assign v37653bf = hlock5 & v376a9aa | !hlock5 & v3a6fc89;
assign v3a70910 = hbusreq3 & v3733cca | !hbusreq3 & v3a70452;
assign v3a6bfea = locked_p & v375ed52 | !locked_p & v8455ab;
assign v3763e88 = hbusreq2 & v3a715d2 | !hbusreq2 & v8455ab;
assign v3747c93 = hbusreq3 & v374cc2a | !hbusreq3 & v3a7162d;
assign v380881d = hbusreq0 & v37406d2 | !hbusreq0 & v8455ab;
assign v3a58d2e = jx0_p & v372c702 | !jx0_p & v3a5e82d;
assign v3a60a56 = hmaster1_p & v3757d76 | !hmaster1_p & v3a70259;
assign v3779cda = hlock7 & v23fe209 | !hlock7 & v375fae9;
assign v3a6a8ee = hbusreq4_p & v372e367 | !hbusreq4_p & v8455ab;
assign v3a6f66a = hmaster0_p & v39ebae8 | !hmaster0_p & v8455ab;
assign v376a63f = hmaster2_p & v3772e0c | !hmaster2_p & v374fe54;
assign v3258762 = hgrant4_p & v377ea72 | !hgrant4_p & v3755451;
assign v375602e = hgrant2_p & v3a6ffb6 | !hgrant2_p & v377c546;
assign v3729d0b = hbusreq5_p & v3a6692b | !hbusreq5_p & !v377439e;
assign v372c4cd = hmaster1_p & v3a5a807 | !hmaster1_p & v3722ebc;
assign v37767d8 = hbusreq2_p & v3a57378 | !hbusreq2_p & v8455ab;
assign v374518e = hmaster0_p & v3a635ea | !hmaster0_p & v3a5e647;
assign v3734e0b = hmaster1_p & v3a6eaef | !hmaster1_p & !v376f8ea;
assign v3a62fa3 = hlock3 & v37408a3 | !hlock3 & v3a71452;
assign v3a6da59 = hmaster1_p & v3723021 | !hmaster1_p & v9e78af;
assign v3a5b47c = hlock6 & v3a5f75a | !hlock6 & v376b082;
assign v3722a42 = jx0_p & v3a6f834 | !jx0_p & v8455ab;
assign v3774f56 = hbusreq5 & v372e365 | !hbusreq5 & v375929c;
assign v375a92b = hbusreq4 & v373eecc | !hbusreq4 & v3a635ea;
assign v372437c = hbusreq6_p & v3737c2f | !hbusreq6_p & v3a6ca53;
assign v3a70a46 = hlock8 & v374990a | !hlock8 & v3745ee1;
assign v35b779c = hmaster0_p & v37710c7 | !hmaster0_p & v23fdad1;
assign v376db34 = hmaster2_p & v3a5727d | !hmaster2_p & v3756c5d;
assign v3747587 = hlock7 & v3772ac1 | !hlock7 & v23fe345;
assign v3739f49 = hmaster1_p & v3a67471 | !hmaster1_p & v8455e7;
assign v23fdaed = hgrant6_p & v8455ca | !hgrant6_p & v3a5b91d;
assign v377c67b = hmaster0_p & v377849a | !hmaster0_p & !d6aeaf;
assign v39a53a1 = hbusreq7 & v3a5f5db | !hbusreq7 & v3a6088f;
assign v374b894 = hbusreq6_p & v37785a8 | !hbusreq6_p & v8455ab;
assign v3774c3f = hbusreq3 & v3a71422 | !hbusreq3 & v8455ab;
assign v3a6ef1e = hlock3 & v37518fa | !hlock3 & v3776ce0;
assign v3a70382 = hmaster0_p & v37483f9 | !hmaster0_p & !v375af99;
assign v3729b9f = hlock0 & v373f3b5 | !hlock0 & v372cfd5;
assign v3a713c9 = hbusreq3_p & v373fa24 | !hbusreq3_p & !v3a707d5;
assign v377c160 = hlock2 & v375b0e8 | !hlock2 & v3a6c7c6;
assign v3725494 = hgrant6_p & v3762385 | !hgrant6_p & v3737628;
assign v3a71071 = hlock6_p & v20d166d | !hlock6_p & v8455ab;
assign v3777989 = hmaster1_p & v3a5d76d | !hmaster1_p & v377c977;
assign v3a6f040 = hlock8_p & v372dc35 | !hlock8_p & v8455ab;
assign v3a6f068 = hmaster1_p & v3a61323 | !hmaster1_p & v372c28d;
assign v3a5a637 = hmaster1_p & v377f113 | !hmaster1_p & v377055c;
assign v3a6fe7c = hbusreq8_p & v3a65b10 | !hbusreq8_p & v3738a2a;
assign v3770abd = hgrant4_p & v1e37996 | !hgrant4_p & v3a6a1b4;
assign v377479e = hbusreq6 & v377e089 | !hbusreq6 & !v8455bd;
assign v373d5f4 = hlock5_p & v3748a16 | !hlock5_p & !v8455d9;
assign v377af0b = hbusreq5 & v3a54264 | !hbusreq5 & v8455ab;
assign v3758a0c = hgrant2_p & v8455ab | !hgrant2_p & v375c01d;
assign v3a71455 = hgrant4_p & v375eaac | !hgrant4_p & v3760748;
assign v3a6dc83 = hbusreq4_p & v3a64792 | !hbusreq4_p & v8455ab;
assign v3a5b5d3 = locked_p & v35772b3 | !locked_p & v35772a6;
assign v1e37d71 = hmaster0_p & v3a5e24e | !hmaster0_p & v3744314;
assign v377e241 = hmaster2_p & v376b397 | !hmaster2_p & v37316c9;
assign v374c009 = hbusreq8_p & v3a67755 | !hbusreq8_p & v37666d7;
assign v373510a = hbusreq0 & v377a751 | !hbusreq0 & v376db8f;
assign v3a7163e = hbusreq0 & v899d31 | !hbusreq0 & v3a7129b;
assign v3a6f238 = hbusreq6 & v3759031 | !hbusreq6 & v8455ab;
assign v3a691fb = hbusreq8 & v3753e8e | !hbusreq8 & v373c7af;
assign v377506b = hbusreq4 & c88c38 | !hbusreq4 & v372c095;
assign v375b8b2 = hbusreq3 & v3743da0 | !hbusreq3 & v3a6f5ea;
assign v380714c = hbusreq6_p & v3a67d66 | !hbusreq6_p & v377824e;
assign v3a57b46 = hmaster0_p & v8455b0 | !hmaster0_p & v3a63866;
assign v3762f51 = hbusreq6_p & v374df1b | !hbusreq6_p & v8455ab;
assign v3807414 = hbusreq7 & v3a71101 | !hbusreq7 & v3764f6a;
assign v3760644 = hmaster0_p & v3754164 | !hmaster0_p & v372efee;
assign v372fd97 = hgrant3_p & v3779060 | !hgrant3_p & v3a69adb;
assign v3759fb4 = hgrant6_p & v3770c9d | !hgrant6_p & v37349d3;
assign v3a5de32 = hbusreq5 & v374bb9f | !hbusreq5 & !v8455ca;
assign v376bb7b = hbusreq6_p & v37308b0 | !hbusreq6_p & v3764bca;
assign v3723bac = hbusreq4 & v376ebbf | !hbusreq4 & v373628e;
assign v376b3bc = hgrant2_p & v3a53f43 | !hgrant2_p & v37501fd;
assign v3a7145b = hgrant0_p & v3753e6a | !hgrant0_p & v3a6fadd;
assign v372a636 = hmaster1_p & v3a70874 | !hmaster1_p & v37735aa;
assign v373a7a1 = hmaster0_p & v3a7006c | !hmaster0_p & v3744d60;
assign v372d336 = hgrant6_p & v3756057 | !hgrant6_p & v3a70b0e;
assign v3a66d74 = hlock7_p & v377df77 | !hlock7_p & v1e382f1;
assign v377cd7e = hlock0 & v375cf36 | !hlock0 & v3736217;
assign v8455ba = hbusreq2 & v8455ab | !hbusreq2 & !v8455ab;
assign v3a6678b = hbusreq5 & v3740c5f | !hbusreq5 & v3a635ea;
assign v373327e = hmaster1_p & v3a637dc | !hmaster1_p & v3a705cb;
assign v37655bf = hmaster1_p & v37364bd | !hmaster1_p & v37249ff;
assign v3a5bb98 = hbusreq2_p & v3a6900b | !hbusreq2_p & v374c4bc;
assign v3a56d06 = hbusreq6_p & v37673d6 | !hbusreq6_p & v8455ab;
assign v3763086 = hgrant5_p & v8455ab | !hgrant5_p & v37744a3;
assign v372954c = hmaster2_p & v38072fd | !hmaster2_p & v8455ab;
assign v3752831 = hlock3 & v37605bb | !hlock3 & v3a6edab;
assign v3a62f72 = hbusreq7 & v3a5c7ca | !hbusreq7 & v3a6fcdf;
assign v373d43a = hmaster2_p & v3761175 | !hmaster2_p & v3755a05;
assign v3a5b28d = hmaster2_p & v8455ab | !hmaster2_p & v374f528;
assign v375b9cc = hmaster0_p & v376aa57 | !hmaster0_p & v374a0eb;
assign v3a6fceb = hmaster3_p & v2678bee | !hmaster3_p & v3737b1a;
assign v376b3d4 = hmaster1_p & v375f906 | !hmaster1_p & v3a62a6d;
assign v3a65160 = hgrant5_p & v37541d4 | !hgrant5_p & v3a6ff07;
assign v3a6e31f = hbusreq6_p & v3a5c945 | !hbusreq6_p & v3a57f59;
assign v37658af = hbusreq2 & v374ad1e | !hbusreq2 & v8455ab;
assign v375adaa = hgrant2_p & v8455ab | !hgrant2_p & v377320f;
assign v37795a3 = hbusreq7_p & v373a373 | !hbusreq7_p & v376d972;
assign v373d3e5 = hmaster0_p & v3a5e2a3 | !hmaster0_p & v3a62f75;
assign v3a6ef4e = hmaster0_p & v373ac15 | !hmaster0_p & v8455ab;
assign v3725b75 = hbusreq4 & v37564e4 | !hbusreq4 & !v8455bd;
assign v37432cd = hgrant4_p & v3769f61 | !hgrant4_p & v376aedb;
assign v3758a02 = hbusreq4 & v3737d44 | !hbusreq4 & !v8455ab;
assign v372a417 = hmaster2_p & v3a635ea | !hmaster2_p & v376bade;
assign v3807550 = hmaster1_p & v3726826 | !hmaster1_p & v3a71050;
assign v373e521 = hlock3 & v377ec08 | !hlock3 & v3a71452;
assign v3a636ce = hmaster0_p & v37287f6 | !hmaster0_p & v3750088;
assign v3a71618 = hlock7_p & v374b08d | !hlock7_p & !v8455ab;
assign v3735afe = hmaster0_p & v3a562a7 | !hmaster0_p & v377e0d2;
assign v3a65f1f = stateA1_p & v37440c3 | !stateA1_p & v3757c6f;
assign v377acc6 = hmaster0_p & v35b774b | !hmaster0_p & v375fcd6;
assign v3a6f192 = hbusreq4 & v3778993 | !hbusreq4 & v8455ab;
assign v3779f0a = hgrant5_p & v37472f4 | !hgrant5_p & v3a71090;
assign v374bfd6 = hbusreq8_p & v37244b9 | !hbusreq8_p & v3a704e1;
assign v3a6f7b6 = hlock8_p & v3a5a8f6 | !hlock8_p & v3a712b9;
assign v3a5d6c6 = hbusreq4 & d2e9f6 | !hbusreq4 & v3a6c5ee;
assign v373bdd1 = hmaster2_p & v3a658bf | !hmaster2_p & v35772a6;
assign v3a71574 = hmaster0_p & v3749336 | !hmaster0_p & v372f07d;
assign v3a68ed1 = hbusreq6 & v372b89e | !hbusreq6 & v376e90a;
assign v37641b8 = hmaster0_p & v37520ee | !hmaster0_p & v3a67b7f;
assign v3724418 = hbusreq3 & v37652a5 | !hbusreq3 & v3a61c41;
assign v372bdb1 = hbusreq7 & v376d559 | !hbusreq7 & v3a581f1;
assign v3737909 = hbusreq0 & v373291e | !hbusreq0 & v373bd6c;
assign v3a6ffd5 = hgrant6_p & v3775537 | !hgrant6_p & v929796;
assign v3776fa4 = hbusreq1_p & v2aca977 | !hbusreq1_p & v372706d;
assign v3770e43 = hgrant2_p & v8455ab | !hgrant2_p & !v8455ef;
assign v3773524 = hmaster0_p & v2aca977 | !hmaster0_p & v375d06d;
assign v37467f7 = hbusreq2_p & v3733d6e | !hbusreq2_p & v372ee7e;
assign v3a6f922 = hlock4_p & v3750d37 | !hlock4_p & !v8455ab;
assign v37462ca = hgrant0_p & v8455ab | !hgrant0_p & !v3741c03;
assign v3a5b286 = hgrant2_p & v37234e0 | !hgrant2_p & !v375cb72;
assign v3a70da2 = hmaster2_p & v8455ab | !hmaster2_p & !v37358ab;
assign v3763043 = hmaster0_p & v376aa57 | !hmaster0_p & v3a5a6fb;
assign v3a5ba95 = jx3_p & v3a66940 | !jx3_p & v373070b;
assign v3806a78 = hmaster2_p & v3753ee0 | !hmaster2_p & v8455ab;
assign v8be8ac = hmaster1_p & v35b774b | !hmaster1_p & v377acc6;
assign v3a617a2 = hlock5_p & v37470e6 | !hlock5_p & !v8455ab;
assign v37758ce = hgrant3_p & v374fb58 | !hgrant3_p & v3a684af;
assign v377e355 = hlock5 & v3a538b3 | !hlock5 & v3a62d5d;
assign v3a63628 = hmaster0_p & v3726458 | !hmaster0_p & v37481bf;
assign v373f8c4 = hgrant5_p & v3a607bd | !hgrant5_p & !v374eb2d;
assign v3770f7a = hready & v3734a99 | !hready & v3a635ea;
assign v377e87e = hbusreq0 & v3754f2e | !hbusreq0 & v373031f;
assign v3a5d327 = hmaster0_p & v3746905 | !hmaster0_p & v3a555b3;
assign v374244e = hbusreq7 & v2acb5c8 | !hbusreq7 & v376c51e;
assign v374e032 = jx0_p & v373e679 | !jx0_p & v3a7135a;
assign v3765053 = hbusreq4 & v374fe1a | !hbusreq4 & v3a69487;
assign v3750c47 = hgrant2_p & v3a6cfe0 | !hgrant2_p & v376bf10;
assign v377fbbf = hmaster2_p & v3760d14 | !hmaster2_p & v376cfaa;
assign v375e04e = hbusreq7 & v377c2ff | !hbusreq7 & v35b774b;
assign v3a6f671 = hmaster2_p & v37379bb | !hmaster2_p & !v377957e;
assign v3777301 = hmaster2_p & v8455ab | !hmaster2_p & v3a697cc;
assign v3771ea7 = hbusreq6_p & v2aca977 | !hbusreq6_p & v3748900;
assign v3752f43 = hgrant5_p & v3730019 | !hgrant5_p & v3774f07;
assign v375d06a = hmaster2_p & v3a7097e | !hmaster2_p & v377d1dc;
assign v3a558ce = hbusreq7_p & v3760e78 | !hbusreq7_p & !v8455ab;
assign v377f1ff = hmaster0_p & v374a8db | !hmaster0_p & v377cccb;
assign v373276f = hbusreq0 & v360d048 | !hbusreq0 & v375559b;
assign v3a6fbd3 = hgrant5_p & v3777670 | !hgrant5_p & v3a60013;
assign v376ace2 = hbusreq6_p & v377b6fc | !hbusreq6_p & !v8455ab;
assign v3a67869 = hgrant4_p & v372493b | !hgrant4_p & v374affb;
assign v3a6d1a4 = hgrant0_p & v3759032 | !hgrant0_p & v3a6f415;
assign v3a70426 = hlock7 & v373b42d | !hlock7 & v37702e0;
assign v2092ab0 = hgrant3_p & v3727eca | !hgrant3_p & v3a5d923;
assign v373523c = hbusreq5_p & v377b24b | !hbusreq5_p & v3761b5e;
assign v377d21c = hmaster2_p & v8455ab | !hmaster2_p & v3735512;
assign v37264a3 = hlock8 & v3a5d4e9 | !hlock8 & v376dcf6;
assign v3a5cfbb = hbusreq5_p & c2e325 | !hbusreq5_p & v375b2af;
assign v3a6f275 = hmaster2_p & v374b3af | !hmaster2_p & v3729eeb;
assign v3a6f70a = hmaster2_p & v8455e7 | !hmaster2_p & v3a55456;
assign v3a6f95f = hgrant0_p & v3a5b71a | !hgrant0_p & !v376ca07;
assign v37473c5 = hmaster0_p & v3a5a510 | !hmaster0_p & v3a6f5a6;
assign v37560ff = hbusreq2_p & v3739336 | !hbusreq2_p & v8455bf;
assign v3a70848 = hgrant6_p & v8455ab | !hgrant6_p & v3808870;
assign v3775bd3 = hbusreq2_p & v3755d64 | !hbusreq2_p & v8455ab;
assign v376b6ba = hbusreq7_p & v3760da6 | !hbusreq7_p & v374d547;
assign v373ce6d = hmaster2_p & v3748ca3 | !hmaster2_p & v3a71350;
assign v3730930 = hmaster2_p & v23fe361 | !hmaster2_p & !v8455ab;
assign v375fe03 = hmaster2_p & v3748016 | !hmaster2_p & v373c2a2;
assign v3a6f327 = hmaster0_p & v3a70cc9 | !hmaster0_p & !v37665e1;
assign v37551b2 = hbusreq5 & v3772bb1 | !hbusreq5 & v3a63f9a;
assign v3768a37 = hgrant6_p & v3763ff7 | !hgrant6_p & !v3730e5d;
assign v3734e58 = hbusreq3_p & v373dfbe | !hbusreq3_p & !v377b3a8;
assign v374c693 = hbusreq1_p & v3a635ea | !hbusreq1_p & v373a7a6;
assign v374c02e = hmaster2_p & v3a5a807 | !hmaster2_p & !v3a6efe3;
assign v3727d95 = hbusreq6_p & v3776592 | !hbusreq6_p & v3806f24;
assign v3a6f0ee = hbusreq3_p & v3a6e438 | !hbusreq3_p & v3807107;
assign v372cb28 = hbusreq4 & v374b3cf | !hbusreq4 & v8455b3;
assign v374e6e3 = hlock0 & v373a341 | !hlock0 & v3a7136a;
assign v3755f22 = hbusreq8_p & v372cdec | !hbusreq8_p & v3750abf;
assign v373bfd9 = hgrant6_p & v3739f07 | !hgrant6_p & v3777cae;
assign v374edba = hmaster0_p & v372d727 | !hmaster0_p & v376d680;
assign b44720 = hlock7 & v37332eb | !hlock7 & v37399d4;
assign v374a36b = hmaster0_p & v3738c5f | !hmaster0_p & v3a6adff;
assign v374beb6 = hbusreq8_p & v376ae9f | !hbusreq8_p & v376ad73;
assign v377b8ee = hlock0_p & v8455b0 | !hlock0_p & v37485bd;
assign v374d7ec = hbusreq5 & v374f712 | !hbusreq5 & v37507dc;
assign v37344a0 = hgrant2_p & v8455ab | !hgrant2_p & v377e087;
assign v37550d4 = hbusreq6_p & v3a55526 | !hbusreq6_p & v3a647e2;
assign v376d774 = hmaster2_p & v3a653e4 | !hmaster2_p & !v3a6b873;
assign v3748bf9 = hgrant3_p & v8455ab | !hgrant3_p & v37273d7;
assign v3a62e99 = hbusreq8_p & v3759569 | !hbusreq8_p & v3776836;
assign v3a715fc = hmaster2_p & v8455ab | !hmaster2_p & v3723a00;
assign v3a61a37 = hlock8_p & v3733998 | !hlock8_p & v3762f2d;
assign v375e64d = hmaster1_p & v2aca977 | !hmaster1_p & v3773524;
assign v3a614d1 = hmaster0_p & v3775721 | !hmaster0_p & v3a70d93;
assign v3777da6 = hgrant4_p & v8455ab | !hgrant4_p & v374baac;
assign v3753093 = hmaster2_p & v3a705f2 | !hmaster2_p & v3a67905;
assign v3a617ad = hbusreq5_p & v3742649 | !hbusreq5_p & ca2eb2;
assign v3768364 = hgrant6_p & v8455ab | !hgrant6_p & v3762949;
assign v3a5877f = hbusreq5 & v374ab03 | !hbusreq5 & v3a7006d;
assign v374385c = hmaster0_p & v3761e62 | !hmaster0_p & !v3a6f6cf;
assign v372bebe = hlock7 & v3a2a106 | !hlock7 & v3a66bfa;
assign v37425a0 = hlock4_p & v3a61c41 | !hlock4_p & v8455b3;
assign v372e5fb = hmaster2_p & v3a6f27d | !hmaster2_p & v375b9c1;
assign v3751fa8 = locked_p & v377b24b | !locked_p & v3a6ffae;
assign v375c1d9 = hgrant4_p & v3729f6c | !hgrant4_p & !v377970b;
assign v3732d0f = hmaster2_p & v3a6fc66 | !hmaster2_p & v8455ab;
assign v37770df = hmaster1_p & v3a635ea | !hmaster1_p & v376502e;
assign v3747d68 = hgrant4_p & v2ff9314 | !hgrant4_p & v3727486;
assign v3742c9b = hmaster2_p & v3a71276 | !hmaster2_p & v376afdf;
assign v3778937 = hlock3_p & v3a6fa64 | !hlock3_p & v3760101;
assign v373cde5 = hmaster0_p & v3a5ec1a | !hmaster0_p & v8455ab;
assign v3a570cd = hbusreq7 & v3a6895d | !hbusreq7 & v3755d10;
assign v3736be5 = hmaster2_p & v3752536 | !hmaster2_p & !v3760700;
assign v375a8d6 = hbusreq5_p & v3a65552 | !hbusreq5_p & v373b4dc;
assign v3a69cd8 = hbusreq0 & v3752c04 | !hbusreq0 & !v3727ce4;
assign v37545ea = hbusreq4_p & v3809112 | !hbusreq4_p & v37328da;
assign v3a633b9 = hmaster2_p & v3747302 | !hmaster2_p & v373ae83;
assign v3745e71 = hbusreq8 & v373a6bf | !hbusreq8 & v376ea50;
assign v3a6727a = hbusreq5 & v3a71133 | !hbusreq5 & v373bf09;
assign v3756aa3 = hbusreq7_p & v3755549 | !hbusreq7_p & v372562a;
assign v37486c2 = hgrant3_p & v8455ab | !hgrant3_p & v375cc28;
assign v3729cfe = hbusreq4 & v3a66d0e | !hbusreq4 & v8455ab;
assign v376ec0d = hbusreq7 & v3a6895d | !hbusreq7 & v37448a7;
assign v3726cc1 = hlock0 & v377ae81 | !hlock0 & v3770ab1;
assign v3a6e21a = hbusreq6 & v3755665 | !hbusreq6 & v375b9c1;
assign v3743604 = hbusreq4 & v376992a | !hbusreq4 & v3a70a7f;
assign v3756dd8 = hmaster2_p & v375463e | !hmaster2_p & v3755b56;
assign v37377cf = hmaster0_p & v37693e7 | !hmaster0_p & v3731bb5;
assign v3806dda = hgrant4_p & v8455ab | !hgrant4_p & v373f0e6;
assign v3a6c0b7 = hlock8_p & v3725dbb | !hlock8_p & v3a61e79;
assign v3a64ef2 = hbusreq8 & v3772c08 | !hbusreq8 & v8455ab;
assign v3a7079a = hmaster0_p & v3774737 | !hmaster0_p & v3756820;
assign v372cdef = hmaster0_p & v3746496 | !hmaster0_p & v3a703b1;
assign v3a6e431 = start_p & v8455ab | !start_p & v845601;
assign v3775d6e = hmaster1_p & v8455ab | !hmaster1_p & v377f06c;
assign v374956a = hlock2 & v377542e | !hlock2 & v3725c68;
assign v3a584bf = hbusreq3 & v3730cda | !hbusreq3 & v8455ab;
assign v37402a4 = hlock7 & v3806465 | !hlock7 & v377cb3d;
assign v8455b2 = hbusreq0 & v8455ab | !hbusreq0 & !v8455ab;
assign v3759361 = hgrant6_p & v3779cf9 | !hgrant6_p & v3729561;
assign v374ace9 = hbusreq8 & v3746aa9 | !hbusreq8 & v3a59ddc;
assign v37328da = hbusreq0 & v3a71283 | !hbusreq0 & v372d967;
assign v377281c = hbusreq7 & v374771c | !hbusreq7 & v3a70e42;
assign v3a71213 = hbusreq0 & v376f7a0 | !hbusreq0 & v3729511;
assign v377b073 = hlock3 & v3a6fc64 | !hlock3 & v37481f3;
assign v3a59f9b = hbusreq4_p & v3a635ea | !hbusreq4_p & v375f370;
assign v3a59aa1 = hmaster2_p & v3a63621 | !hmaster2_p & v3a68d2e;
assign v37621e9 = hbusreq4 & v3763a20 | !hbusreq4 & v8455bf;
assign d99853 = hbusreq2_p & v373fe5e | !hbusreq2_p & v8455e7;
assign v3735d71 = hbusreq6_p & v3754fac | !hbusreq6_p & v377535a;
assign v3a700ac = hgrant6_p & v3736f2a | !hgrant6_p & v3a5d6a6;
assign v3761d47 = hmaster2_p & v37386c6 | !hmaster2_p & v372b881;
assign v3761d9f = hbusreq5 & v3808dd0 | !hbusreq5 & v372b27e;
assign v37399ef = hmaster1_p & v3a669c6 | !hmaster1_p & v376ee62;
assign v3765b88 = hbusreq0_p & v8455ab | !hbusreq0_p & v3379037;
assign v37378a3 = hbusreq8_p & v3723de9 | !hbusreq8_p & v373f418;
assign v3a701c4 = hgrant4_p & v375cc1b | !hgrant4_p & a90ef2;
assign v374742c = hlock4_p & v3728e1d | !hlock4_p & v372f071;
assign v3724bbf = jx1_p & v3749a29 | !jx1_p & v3a5657a;
assign v38073d4 = hmastlock_p & v37794be | !hmastlock_p & !v8455ab;
assign v374ed52 = hbusreq0 & v376a97b | !hbusreq0 & v3a5bac7;
assign v3a5f5db = hmaster1_p & v3a7010d | !hmaster1_p & v38064e3;
assign v374e800 = hmaster1_p & v374fb30 | !hmaster1_p & v376e441;
assign v3727713 = hlock6 & v3a6b15d | !hlock6 & v37565a5;
assign v3a6b1bf = hbusreq5 & v3a7022f | !hbusreq5 & v3a6d6fb;
assign v376c505 = hbusreq5_p & v3742a61 | !hbusreq5_p & v3a61094;
assign v374b8fe = hmaster1_p & v3a66110 | !hmaster1_p & v374fb02;
assign v3a5ee3a = hgrant2_p & v3a6d349 | !hgrant2_p & v37510ae;
assign v3749586 = hgrant2_p & v3a6fcc0 | !hgrant2_p & v377636a;
assign v3a6443f = jx1_p & v376dd80 | !jx1_p & v8455ab;
assign v3a6ec94 = stateG10_1_p & v3a6f436 | !stateG10_1_p & v376498a;
assign v374a296 = hmaster0_p & v3768ec7 | !hmaster0_p & v3a700a8;
assign v374c53a = hgrant6_p & v3a5c945 | !hgrant6_p & v373e748;
assign v377a942 = hbusreq4_p & v376aedb | !hbusreq4_p & v3a5f2c7;
assign v3762199 = hbusreq8 & v8fdd0d | !hbusreq8 & v3754d67;
assign v3724f54 = hbusreq1_p & v3a69de7 | !hbusreq1_p & v3a635ea;
assign v376cd84 = hmaster2_p & v3749356 | !hmaster2_p & v3a712bf;
assign v376a0f6 = hmaster2_p & v3a70147 | !hmaster2_p & v37769cc;
assign v374e7c5 = hbusreq4 & v376d9ad | !hbusreq4 & v8455e7;
assign v3a71542 = hlock0_p & a38ed7 | !hlock0_p & v37237bc;
assign v37788fc = hbusreq4_p & v3767650 | !hbusreq4_p & v375fdf5;
assign v372523e = hlock5_p & v3a55672 | !hlock5_p & v8455ab;
assign v3a5d20a = hbusreq7 & v37464f3 | !hbusreq7 & v3a712bb;
assign v3771232 = jx0_p & v3762d26 | !jx0_p & v37501e6;
assign v3759a00 = hgrant6_p & v377b6ce | !hgrant6_p & !v3a71354;
assign v372dc51 = hbusreq4_p & v32562a3 | !hbusreq4_p & v3a6bf63;
assign v3730097 = jx3_p & v3751fde | !jx3_p & v3a6b001;
assign v3a6f386 = hbusreq2 & v3a62a96 | !hbusreq2 & v375c1d1;
assign v3739d22 = hlock3 & v3a70dd0 | !hlock3 & v3762d80;
assign v3a6f8a0 = hbusreq4_p & v3a70e69 | !hbusreq4_p & v3a7139f;
assign v3808cf5 = hmaster3_p & v373ed37 | !hmaster3_p & v3730617;
assign v3a6f2a8 = hlock4_p & v8455e7 | !hlock4_p & !v8455ab;
assign v3a70606 = hbusreq5 & v3732558 | !hbusreq5 & v8455ab;
assign v3a6f134 = hmaster2_p & v3a6fb0c | !hmaster2_p & v3a6fa78;
assign v375c724 = hbusreq7_p & v377d850 | !hbusreq7_p & v3a703ab;
assign v3723be4 = hmaster2_p & v372386d | !hmaster2_p & v376d98d;
assign v374fd8a = hgrant6_p & v3a53f00 | !hgrant6_p & v3a605e2;
assign v3734081 = hbusreq5_p & v3a6cc93 | !hbusreq5_p & v3750ae0;
assign v377d891 = hmaster2_p & v3a70bf4 | !hmaster2_p & v37249cc;
assign v3a71344 = hbusreq2 & v37457fb | !hbusreq2 & v8455ab;
assign v37535bd = hgrant2_p & v8455ab | !hgrant2_p & v37273be;
assign v377af44 = hbusreq2_p & v8455ab | !hbusreq2_p & v3a6a939;
assign v3a62113 = hmaster2_p & v3a60a68 | !hmaster2_p & v374d0e3;
assign v373d6dd = hgrant5_p & v8455ab | !hgrant5_p & v373dff9;
assign v37679d9 = hbusreq4 & v377e1f6 | !hbusreq4 & v3727084;
assign v3a6f369 = hbusreq7 & v374771c | !hbusreq7 & v3a709f1;
assign v3747a53 = hbusreq6_p & v3a70a0e | !hbusreq6_p & v376fdb9;
assign v3a57de9 = hmaster0_p & v3a7002c | !hmaster0_p & v3a701e0;
assign v3a558c2 = hbusreq3 & v376430b | !hbusreq3 & v376653d;
assign v325b59f = hbusreq0 & v37778e2 | !hbusreq0 & v377f180;
assign v3a62f0f = hbusreq8_p & v376376a | !hbusreq8_p & v3a6f964;
assign v373d235 = hbusreq8 & cdcddf | !hbusreq8 & v3a576bd;
assign v3a702e5 = hbusreq2_p & v37495f2 | !hbusreq2_p & v8455ab;
assign v375ba66 = hbusreq5 & v3771882 | !hbusreq5 & v37363ae;
assign v3724c63 = hmaster0_p & v377167c | !hmaster0_p & v3731d67;
assign v994115 = hmaster1_p & v3a65b79 | !hmaster1_p & c4699e;
assign v37565c7 = hgrant6_p & v3771fb3 | !hgrant6_p & v3a6ff4c;
assign v375bf61 = hmaster2_p & v3771076 | !hmaster2_p & v3a70374;
assign v377b9a2 = hmaster0_p & v3a5fc34 | !hmaster0_p & v3a710f0;
assign v3a6a8d2 = hlock3_p & v3764261 | !hlock3_p & v8455b0;
assign v37434f4 = hbusreq2 & v3a5ad94 | !hbusreq2 & v3a5f5bb;
assign v3743cb5 = hlock2_p & v380971a | !hlock2_p & v8455b0;
assign v3a704c0 = hgrant0_p & v37773a9 | !hgrant0_p & ae6485;
assign v3770093 = hmaster2_p & v3a5e24e | !hmaster2_p & !v2092faa;
assign v376e833 = hbusreq2 & v3735809 | !hbusreq2 & v3a5b6de;
assign v373f56b = stateG10_1_p & v8455ab | !stateG10_1_p & !v37426ed;
assign b2d8a6 = hbusreq7 & v3a6a8b2 | !hbusreq7 & v3a67b58;
assign v375f86d = hlock7 & v3a630bc | !hlock7 & v3a55ab6;
assign v3a62a2d = hmaster1_p & v3a637dc | !hmaster1_p & v373d381;
assign v376fa80 = hgrant0_p & v37490cb | !hgrant0_p & v37417f6;
assign v3772f74 = hlock5 & v3a6b1bf | !hlock5 & v3a7022f;
assign v376f911 = hbusreq3 & v37796c6 | !hbusreq3 & v8455ab;
assign v3754fc6 = hlock8 & v37783d2 | !hlock8 & v3a701f7;
assign v3765dbe = hbusreq5_p & v3730370 | !hbusreq5_p & v3742950;
assign v3a71378 = hgrant0_p & v8455ab | !hgrant0_p & v3a5d448;
assign v3766d4b = hmaster0_p & v37377df | !hmaster0_p & v3729793;
assign v372422d = hgrant2_p & v3751d98 | !hgrant2_p & v3a6fd95;
assign v372ddbc = hmaster1_p & v375df71 | !hmaster1_p & v373fb22;
assign v376a4d3 = hgrant6_p & v37414b0 | !hgrant6_p & v3762db3;
assign v3754450 = hgrant6_p & v3729d65 | !hgrant6_p & v2aca977;
assign v3a7132d = hmaster1_p & v8455e7 | !hmaster1_p & v372e868;
assign v373b0a4 = hlock0_p & v376d793 | !hlock0_p & v3a707bb;
assign v3a6d33e = hmaster2_p & v1e382e7 | !hmaster2_p & !v1e38224;
assign v3753e3b = hbusreq7 & v37798bb | !hbusreq7 & v3737808;
assign v372bf1d = hgrant5_p & v8455ab | !hgrant5_p & v3a701ac;
assign v37774c7 = hlock0_p & v39a4e5f | !hlock0_p & v376773a;
assign v3a6c1d3 = hmaster2_p & v3a7101b | !hmaster2_p & v372cc25;
assign v37721fa = hmaster2_p & v376a6f1 | !hmaster2_p & !v8455ab;
assign v3773bd7 = jx2_p & v3763387 | !jx2_p & v3770359;
assign v375a8cf = hbusreq6 & v373a4e4 | !hbusreq6 & v3a70d99;
assign v3764109 = hmaster1_p & v37784d0 | !hmaster1_p & v3a70259;
assign v3a7113f = hbusreq8 & v3a6fd21 | !hbusreq8 & v8455ab;
assign v3760549 = hbusreq2 & v8455ab | !hbusreq2 & v3758233;
assign v37245a1 = hmaster0_p & v376c89f | !hmaster0_p & v948ef2;
assign v375c5cf = hbusreq3_p & v8455ab | !hbusreq3_p & v3a684af;
assign v3727c07 = hmaster0_p & v375abab | !hmaster0_p & v3a6fbd1;
assign v37241cc = hbusreq1_p & v35b70a0 | !hbusreq1_p & v8455ab;
assign v372b5b0 = hgrant0_p & v8455ab | !hgrant0_p & v375cea7;
assign v372c86a = hgrant6_p & v3a7138d | !hgrant6_p & v372f192;
assign v377a9b2 = hmaster1_p & v374a9d4 | !hmaster1_p & !v3768ae9;
assign v375b534 = hmaster2_p & v8455ab | !hmaster2_p & v374890e;
assign v376c76d = hgrant6_p & v3a70b92 | !hgrant6_p & v372c500;
assign v372de54 = hbusreq8_p & v3744990 | !hbusreq8_p & v3726d0c;
assign v3762363 = hgrant5_p & v8455ab | !hgrant5_p & v3724014;
assign v3a7139e = hlock3 & v377b292 | !hlock3 & v3807c0c;
assign v3751631 = hmaster2_p & v37325a2 | !hmaster2_p & v373de4b;
assign v3a6eb39 = hbusreq3_p & v3722e5c | !hbusreq3_p & v35772a6;
assign v3761f57 = jx1_p & v3a644ac | !jx1_p & v3a621e6;
assign afadd1 = hmaster0_p & v3740404 | !hmaster0_p & v3807670;
assign v376730a = hmaster2_p & v3a5bc2c | !hmaster2_p & v3a6f9c3;
assign v3a5a6cc = hbusreq5_p & v372fa9d | !hbusreq5_p & v377816f;
assign v3779709 = hgrant1_p & v3a70011 | !hgrant1_p & v39a537f;
assign v3a5bd12 = hbusreq8_p & v372953c | !hbusreq8_p & v8455ab;
assign v375ba6d = hbusreq5 & v3a71399 | !hbusreq5 & cc2999;
assign v3a6f7e4 = hbusreq7 & v375b247 | !hbusreq7 & v3767b70;
assign v3738ad8 = hbusreq0 & v3808dca | !hbusreq0 & v375a65f;
assign v3800ee4 = hgrant5_p & v3a711d5 | !hgrant5_p & v3a5551b;
assign v3806e5b = jx0_p & v3a6c849 | !jx0_p & v3a70989;
assign v37257e9 = hbusreq5 & v37354a9 | !hbusreq5 & v3742cd4;
assign b8cdcc = hgrant7_p & v8455ab | !hgrant7_p & v3736079;
assign v3764d6b = hmaster2_p & v1e382e7 | !hmaster2_p & !v3a5bf04;
assign v3a5d5e7 = hgrant6_p & v8455ca | !hgrant6_p & v3a55954;
assign v373fd94 = hmaster2_p & v3a635ea | !hmaster2_p & v376e041;
assign v3769160 = hgrant6_p & v3a57b60 | !hgrant6_p & v3a71302;
assign v3a6ebcc = hgrant2_p & v1e378b4 | !hgrant2_p & v376d7ee;
assign v37386f2 = start_p & v8455ab | !start_p & !v373aaca;
assign v3a71043 = hmaster1_p & v3736610 | !hmaster1_p & v375d9ad;
assign v37722a0 = hmaster2_p & v3a70a7f | !hmaster2_p & v3748d67;
assign v3736fc4 = hbusreq2_p & v373e877 | !hbusreq2_p & v3750178;
assign v375100c = hmaster2_p & v8455ab | !hmaster2_p & !v3748ca3;
assign v3752c99 = hgrant2_p & v8455ab | !hgrant2_p & v377dae6;
assign v3759c2e = hlock0_p & v376e914 | !hlock0_p & !v3a658bf;
assign bb97e8 = hgrant4_p & v8455ab | !hgrant4_p & v3a5a16a;
assign v3a691f2 = hbusreq4_p & v3726d1f | !hbusreq4_p & v3752cf6;
assign v3a6f3df = hgrant5_p & v375c07c | !hgrant5_p & !v8455ab;
assign v3779e1b = hgrant4_p & v3a7049a | !hgrant4_p & v3a7165d;
assign v3726ec0 = hgrant5_p & v8455ab | !hgrant5_p & v3a7047d;
assign v376c343 = hgrant0_p & v3735525 | !hgrant0_p & v375aae9;
assign v377cd9c = hbusreq7_p & v3762f2d | !hbusreq7_p & !v3725470;
assign v37711c3 = hgrant4_p & v374693f | !hgrant4_p & v3764809;
assign v376629a = hgrant4_p & v3769e94 | !hgrant4_p & v376cdf3;
assign v3a71083 = hbusreq5_p & bfe049 | !hbusreq5_p & v376cda5;
assign v372bdca = hgrant6_p & v37331af | !hgrant6_p & v377ee3c;
assign v375471b = hmaster0_p & v372e94f | !hmaster0_p & !v37712b7;
assign v3768c4c = hbusreq6 & v3a6beb6 | !hbusreq6 & v3a7011e;
assign v377108d = hmaster2_p & v3a6f4ba | !hmaster2_p & v3759387;
assign v3765ed6 = hbusreq8 & v37477b7 | !hbusreq8 & v374a565;
assign v3764099 = jx0_p & v3748251 | !jx0_p & v374e61c;
assign v360d0db = hbusreq3_p & v373c064 | !hbusreq3_p & v3a5bb64;
assign v3a54c2e = hready & v8455ab | !hready & v3a707c2;
assign v3769f60 = jx0_p & v37515e1 | !jx0_p & v8455ab;
assign v3732a31 = hlock7 & v377375f | !hlock7 & v3a700be;
assign v3a661cd = hbusreq7_p & v376740b | !hbusreq7_p & v377b3d5;
assign v3735485 = hmaster2_p & v1e37ca4 | !hmaster2_p & v3744ff3;
assign v3a6c7e8 = hmaster0_p & v3757d75 | !hmaster0_p & v3a70c91;
assign v3a7020b = hgrant6_p & v372bfa1 | !hgrant6_p & v3a62348;
assign v3746846 = hmaster2_p & v3a70f1c | !hmaster2_p & v3744a21;
assign v3727e69 = hmaster2_p & v3a635ea | !hmaster2_p & v37716ca;
assign v3a58907 = hbusreq0 & v3777342 | !hbusreq0 & v3743c22;
assign hmaster3 = v31c329f;
assign v23fd817 = hbusreq5 & v377d06b | !hbusreq5 & v3742efa;
assign v92acd8 = hlock6_p & v8455ab | !hlock6_p & !v376430b;
assign v3a70ee1 = hgrant2_p & v37314b5 | !hgrant2_p & v3a70b5d;
assign v3a68c0e = hbusreq0 & v374933f | !hbusreq0 & v373ab9e;
assign v3758f64 = hbusreq3_p & v3751e8d | !hbusreq3_p & !v377b3a8;
assign v3a6325a = hlock0_p & v375863a | !hlock0_p & v3a702a5;
assign v3a6f740 = hlock5_p & v3a7104e | !hlock5_p & v37511c6;
assign v374b0fb = hmaster2_p & v8455ab | !hmaster2_p & v375d3a2;
assign v372cbdb = hbusreq4 & v3a5e7fe | !hbusreq4 & v8455bb;
assign v3a62b11 = hbusreq4 & v3a6fd68 | !hbusreq4 & v8455ab;
assign v3a70c7f = hbusreq4 & v373b78b | !hbusreq4 & v3a6f044;
assign v376c7cc = hmaster0_p & v376f70a | !hmaster0_p & !v3a61c70;
assign v374c862 = hburst0 & v3745509 | !hburst0 & v8455ab;
assign v3a6f829 = hmaster0_p & v377b07a | !hmaster0_p & v3a6af83;
assign v3a6f2c6 = hbusreq5_p & v375016d | !hbusreq5_p & !v8455ab;
assign v3a6fb75 = hmaster1_p & v3727026 | !hmaster1_p & v376f2c8;
assign v376d793 = hlock1 & v374197c | !hlock1 & v3a70c94;
assign v375b031 = jx1_p & v377a4ef | !jx1_p & v37486d7;
assign v3a7119f = hbusreq4_p & v377876f | !hbusreq4_p & v8455ab;
assign v3a71437 = hgrant3_p & v8455ab | !hgrant3_p & !v37709c5;
assign v3743c51 = hlock6 & v3a70bff | !hlock6 & v373081f;
assign v3726f57 = hbusreq4_p & v3772a9b | !hbusreq4_p & v37331a1;
assign v3a6ae3e = hlock2 & v374172f | !hlock2 & v376d4ee;
assign v373fcc7 = hbusreq8_p & v3759569 | !hbusreq8_p & v3a6ef07;
assign v37474e1 = hbusreq5_p & v3728270 | !hbusreq5_p & v372b9d7;
assign d039bc = hlock4_p & v3a64f2d | !hlock4_p & v37395f5;
assign v3778ecc = hmaster2_p & v3736f61 | !hmaster2_p & v37386da;
assign v3737fe0 = hgrant1_p & v3a6d684 | !hgrant1_p & v3a70c07;
assign v3a71513 = hgrant6_p & v377f09a | !hgrant6_p & v3747f5d;
assign v373b938 = hbusreq7 & v3a65dad | !hbusreq7 & v374c28d;
assign v3750b71 = hgrant4_p & v3a704c7 | !hgrant4_p & !v37540df;
assign v3a5d11d = hmaster1_p & v3a67f5b | !hmaster1_p & !v372bc46;
assign v37405a3 = hbusreq8 & v3a66920 | !hbusreq8 & v374d409;
assign v376728e = hbusreq2_p & v374212c | !hbusreq2_p & !v8455ab;
assign v3743fba = hmaster2_p & v3a635ea | !hmaster2_p & v3a5f8a2;
assign v3762997 = hmaster2_p & v377accc | !hmaster2_p & v37745a0;
assign v3727e56 = hbusreq5_p & v374c288 | !hbusreq5_p & v3742cd5;
assign v374a84c = hgrant2_p & v8455b9 | !hgrant2_p & v3739062;
assign v372c08d = hmaster0_p & v3a6f6e2 | !hmaster0_p & v376305d;
assign v3751c73 = hmaster2_p & v3761719 | !hmaster2_p & v3777da6;
assign v3a63111 = hmaster2_p & v3725f77 | !hmaster2_p & !v3a6febd;
assign v373e2bc = jx1_p & v374b237 | !jx1_p & !v377c29b;
assign v3a57b88 = hbusreq4_p & v3a6ef00 | !hbusreq4_p & v3a6f902;
assign v3777853 = hbusreq5_p & v3749ab1 | !hbusreq5_p & v35ba1cf;
assign v37229c2 = hbusreq6_p & v3a5b5c4 | !hbusreq6_p & v8455bf;
assign v3a59529 = hmaster0_p & v3757ce3 | !hmaster0_p & !v3752b8f;
assign v3731c6f = hbusreq4_p & v372bd23 | !hbusreq4_p & v375265e;
assign v3775651 = hmaster0_p & v37582dc | !hmaster0_p & v3764683;
assign v3a6cb19 = hbusreq6 & v3a6fbd9 | !hbusreq6 & v3a6f3f9;
assign v3a6f619 = hgrant8_p & v8686c3 | !hgrant8_p & !v8455ab;
assign v37454c6 = hmaster0_p & v3a702c0 | !hmaster0_p & v3754d88;
assign v3a6275e = hbusreq5 & v374ad45 | !hbusreq5 & v3770aee;
assign v3a70be1 = hbusreq8 & v3768274 | !hbusreq8 & v3757bf1;
assign v375ea72 = hbusreq2_p & v376e093 | !hbusreq2_p & v8455ab;
assign v3a56cdb = hbusreq2_p & v376d45f | !hbusreq2_p & v3a5bf04;
assign v376ea88 = hbusreq7 & v3a5bc4f | !hbusreq7 & v376ae9f;
assign v377d9ab = jx0_p & v8455ab | !jx0_p & v3771b2a;
assign v39378d6 = hgrant3_p & v8455ab | !hgrant3_p & v8455bd;
assign v372704f = hbusreq8 & v3a6ed55 | !hbusreq8 & v8455c6;
assign v3a710f3 = hbusreq0 & v3732355 | !hbusreq0 & v3a70821;
assign v375c265 = hgrant2_p & v3a6f92f | !hgrant2_p & v3775642;
assign v374d173 = hbusreq2 & v3a5b213 | !hbusreq2 & v8455ab;
assign v377320f = hgrant3_p & v8455ab | !hgrant3_p & v3771720;
assign v39ebae8 = hmaster2_p & v8455ab | !hmaster2_p & !v3777deb;
assign v375c707 = stateG10_1_p & v3a5ce2d | !stateG10_1_p & v3758225;
assign v3777340 = hbusreq7_p & v374650b | !hbusreq7_p & v373478e;
assign v3a60131 = hgrant5_p & v3732849 | !hgrant5_p & v3a6540f;
assign v374b0bc = hgrant6_p & v3a69146 | !hgrant6_p & v3723549;
assign v3a6f1e4 = hbusreq0 & v373481c | !hbusreq0 & v375e973;
assign v3a70aa8 = hmaster3_p & v8455ab | !hmaster3_p & v3750da4;
assign v372a0bd = hgrant0_p & v3a6d18a | !hgrant0_p & v37772bf;
assign v3768f5f = hbusreq4_p & v3746259 | !hbusreq4_p & v3749a32;
assign v37728b9 = hmaster2_p & v3a6fe1a | !hmaster2_p & !v8455ab;
assign v375888e = hbusreq5 & b7dcc5 | !hbusreq5 & v8455ab;
assign v376a87b = hbusreq3 & v3a6430c | !hbusreq3 & v38072fd;
assign v37646ce = hlock8 & v3728840 | !hlock8 & v376cfc9;
assign v374d859 = hbusreq4_p & v373bf3c | !hbusreq4_p & v8455ab;
assign v3a61fcc = hbusreq6_p & v3742657 | !hbusreq6_p & v3744458;
assign v377b983 = hbusreq2_p & v373b8ff | !hbusreq2_p & v3a53f45;
assign v373a1f2 = hgrant0_p & v377b6ce | !hgrant0_p & v3a7044c;
assign v3a66632 = hmaster0_p & v377f5f2 | !hmaster0_p & v377b2f3;
assign v3a63831 = hbusreq5 & v3a701fa | !hbusreq5 & v3a6513d;
assign v3a69d06 = hbusreq3 & v376a8d5 | !hbusreq3 & v3a57309;
assign v3773e2a = hlock3_p & v3a71284 | !hlock3_p & v3a6f986;
assign v3a6d401 = hmaster1_p & v372455c | !hmaster1_p & v3722eee;
assign v373fcf4 = hbusreq2 & v3a5f0b2 | !hbusreq2 & v377b774;
assign v3a6b14a = hbusreq4_p & v3a7157e | !hbusreq4_p & v377b2d0;
assign v3a54853 = hlock6_p & v377ea86 | !hlock6_p & !v8455ab;
assign v37320ff = hbusreq4_p & v37786a6 | !hbusreq4_p & v376bb26;
assign v3a6c6d6 = hgrant6_p & v372919a | !hgrant6_p & v37315d5;
assign v374fa18 = hmaster1_p & v3a635ea | !hmaster1_p & v376dd64;
assign v374cad6 = hmaster3_p & v3a7166b | !hmaster3_p & v37348e5;
assign v3a565bc = hlock7_p & v3807008 | !hlock7_p & v3735fb2;
assign v373f8c8 = hlock8_p & v37308ae | !hlock8_p & v3a70b46;
assign v3a62cf3 = hgrant5_p & v3a56bb5 | !hgrant5_p & v3742d6c;
assign d6aeaf = hmaster2_p & v8455ab | !hmaster2_p & v377409c;
assign v3739815 = hbusreq0 & v3768202 | !hbusreq0 & !v373e814;
assign v3a6b285 = hmaster0_p & v3a6f443 | !hmaster0_p & v3a6ad0b;
assign v3a6fb00 = hmaster2_p & v8455e7 | !hmaster2_p & v373fe5e;
assign v3a70501 = hmaster0_p & v3779183 | !hmaster0_p & v3a6f736;
assign v3728346 = hbusreq2 & v3a66538 | !hbusreq2 & v3a5b614;
assign v3a68f04 = hbusreq0 & v3723aa8 | !hbusreq0 & v8455ab;
assign v3726abd = hburst1_p & v8455ab | !hburst1_p & v845605;
assign v3a5db41 = hbusreq4 & v3a6dc08 | !hbusreq4 & v8455b0;
assign v376c5af = hmaster0_p & v374cbc4 | !hmaster0_p & v376981e;
assign v37314d7 = hmaster1_p & v3a69267 | !hmaster1_p & v373bc2f;
assign v3a53e0e = hlock4_p & v3a70f29 | !hlock4_p & v8455ab;
assign v3a6f817 = hbusreq6_p & v8455ab | !hbusreq6_p & v3760b3d;
assign v3a6eb95 = hbusreq4_p & v3733fad | !hbusreq4_p & v3a70509;
assign v3a69b19 = hlock5 & v3a5b181 | !hlock5 & v377b6de;
assign v3745658 = hbusreq4_p & v37276f2 | !hbusreq4_p & v37480ec;
assign v3a6e438 = hgrant0_p & v3723430 | !hgrant0_p & v375863a;
assign v3a7099f = jx3_p & v3774af1 | !jx3_p & v9342d1;
assign v375e64c = hbusreq4 & v3a710c1 | !hbusreq4 & v2092abe;
assign v8db8b7 = hbusreq5_p & v376226e | !hbusreq5_p & v3733993;
assign v377957a = hmaster2_p & v8455ab | !hmaster2_p & !v3a690c2;
assign v374f860 = hbusreq2 & v3a6f8de | !hbusreq2 & v3a62a6d;
assign v375b8a2 = hbusreq5 & v374afa3 | !hbusreq5 & v3a704e3;
assign v3758c41 = hmaster0_p & v3a6eefb | !hmaster0_p & v3a59609;
assign v3a650a6 = hbusreq5 & v3722a46 | !hbusreq5 & v375d417;
assign v3733767 = hmaster2_p & v3a6854c | !hmaster2_p & v3a712af;
assign v374d3b3 = hbusreq6_p & v3a6e6c9 | !hbusreq6_p & v373a2f2;
assign v376a94e = hmaster0_p & v372ddf8 | !hmaster0_p & v3a706cb;
assign v3779879 = hbusreq8_p & v372e77b | !hbusreq8_p & v3a7142e;
assign v374bac7 = hbusreq5_p & v375b01e | !hbusreq5_p & v3a6f894;
assign v3a70461 = hlock7 & v3775b2f | !hlock7 & v375e29b;
assign v3a62bcf = hbusreq5 & v375a4ba | !hbusreq5 & v3a5e030;
assign v3a56b92 = hbusreq5_p & v3a6ebc9 | !hbusreq5_p & v8455ab;
assign v37662d3 = hbusreq6 & v376cad6 | !hbusreq6 & v3768ef1;
assign v374dddd = jx3_p & v3742ffc | !jx3_p & v37294f4;
assign v3776a3e = hmaster2_p & v3775303 | !hmaster2_p & v3749907;
assign v1e374d4 = hmaster0_p & v37731ce | !hmaster0_p & v3a5f3a1;
assign v376c72f = hbusreq3_p & v37487b0 | !hbusreq3_p & v373ad95;
assign v377ad9c = hbusreq4 & v374bf55 | !hbusreq4 & v8455ab;
assign v37716ca = hbusreq4_p & v375da10 | !hbusreq4_p & v376bb26;
assign v377a1d3 = hlock6 & v3a6ffab | !hlock6 & v374944b;
assign v3763afe = hmaster3_p & v37291f8 | !hmaster3_p & v37315fd;
assign v3760d14 = hbusreq4_p & v372eabb | !hbusreq4_p & !v8455ab;
assign v3a57d1f = hmaster2_p & v374282f | !hmaster2_p & !v3735b3e;
assign v3737d44 = hlock0_p & v39a537f | !hlock0_p & v3a702aa;
assign v377b030 = hgrant4_p & v37598ab | !hgrant4_p & v3740b8d;
assign v3723da9 = hbusreq0 & v39a5381 | !hbusreq0 & !v8455ab;
assign v3a6c5ee = hbusreq1_p & v37496fa | !hbusreq1_p & v3743b9e;
assign v375538e = hmaster1_p & v3a6f158 | !hmaster1_p & v23fd89c;
assign v3760ca3 = hbusreq8_p & v37303f0 | !hbusreq8_p & v3763502;
assign v3a70b66 = hgrant2_p & v375975b | !hgrant2_p & v3a6f119;
assign v3a6f4f4 = hbusreq2_p & v3a6fdf8 | !hbusreq2_p & v3a6eb5a;
assign v3765511 = hgrant4_p & v8455ab | !hgrant4_p & v2ff9291;
assign v3a70ad4 = hbusreq6 & v372ab46 | !hbusreq6 & v8455b3;
assign v3a53dbf = hgrant3_p & v8455be | !hgrant3_p & !v376dc58;
assign v3a594e8 = hbusreq8_p & v375d23b | !hbusreq8_p & v3a62a2d;
assign v3754603 = hgrant4_p & v8455ab | !hgrant4_p & v3a6ea3b;
assign v3a5bff1 = hgrant6_p & v8455ab | !hgrant6_p & v3770e43;
assign v3741b49 = hbusreq8 & b30936 | !hbusreq8 & v376ae9f;
assign v372567a = hmaster2_p & v3727943 | !hmaster2_p & v373ae83;
assign v3a6c4b3 = hmaster2_p & v3a6dc08 | !hmaster2_p & v373ee80;
assign v3a70a33 = hmaster2_p & v3a63ea7 | !hmaster2_p & v3753dab;
assign v3771533 = hgrant5_p & v376a77a | !hgrant5_p & v376b0cc;
assign v376644e = hbusreq5_p & v8455ab | !hbusreq5_p & v3722d5a;
assign v3a6fe35 = hbusreq4_p & v3a70725 | !hbusreq4_p & v37679d9;
assign v3730ca3 = stateG10_1_p & v37665bf | !stateG10_1_p & v3723aea;
assign v376b5f8 = hbusreq2_p & v37538f5 | !hbusreq2_p & v3742ce8;
assign v3741baf = hmaster2_p & v3a63e82 | !hmaster2_p & v3a56c66;
assign v3776479 = jx1_p & v374eec1 | !jx1_p & v37342ec;
assign v376306b = hbusreq2 & v37356f0 | !hbusreq2 & v8455ab;
assign v373619d = hgrant2_p & v3a71460 | !hgrant2_p & v373d62b;
assign v374704d = hlock6_p & v8455ab | !hlock6_p & !v3a6ac2a;
assign v94ea62 = hbusreq3_p & v377eaf2 | !hbusreq3_p & v3727aa3;
assign v3a634c9 = hgrant6_p & v3a5fb15 | !hgrant6_p & !v8455ab;
assign v372a460 = hbusreq5 & v9ae4c2 | !hbusreq5 & v3a635ea;
assign v3a5ab85 = hgrant6_p & v8455ab | !hgrant6_p & v373e031;
assign v37590d1 = hgrant4_p & v3723299 | !hgrant4_p & v3a702cc;
assign v1e3773a = hmaster2_p & v376a2c0 | !hmaster2_p & !v8455ab;
assign b0c091 = hbusreq1_p & v373fe5e | !hbusreq1_p & v8455e7;
assign v373a57d = hmaster0_p & v3a69de7 | !hmaster0_p & v376752b;
assign v3758a10 = hgrant6_p & v3743eae | !hgrant6_p & v37463a6;
assign v3736471 = hmaster0_p & v3a548c2 | !hmaster0_p & v3a658cf;
assign v3a623cb = hgrant6_p & v8455ab | !hgrant6_p & v3732d8f;
assign v3a6fa4d = hmaster2_p & v8455ab | !hmaster2_p & v3a6fffd;
assign v372a06a = hmaster1_p & v3a71588 | !hmaster1_p & v373c23c;
assign v3741609 = hbusreq4_p & v3722d9d | !hbusreq4_p & v3a60620;
assign v3a6a33a = hbusreq5_p & v3a715d6 | !hbusreq5_p & !v3736d97;
assign v375dab2 = hbusreq6_p & v8455ab | !hbusreq6_p & v375968a;
assign v3a6ffde = jx1_p & d03e23 | !jx1_p & v3a6bf00;
assign v37328a1 = stateG10_1_p & v3763961 | !stateG10_1_p & v373df14;
assign v372d24a = hbusreq5 & v3744bed | !hbusreq5 & v8455ab;
assign v372ab23 = hbusreq4_p & v3729186 | !hbusreq4_p & v8455ab;
assign v37443d6 = hgrant1_p & v3a6ebe7 | !hgrant1_p & v3a70d71;
assign v376fa50 = hmaster1_p & v3763c97 | !hmaster1_p & !v8455c3;
assign v377181f = hmaster2_p & v3767e76 | !hmaster2_p & !v3a7136e;
assign v3a709f7 = hmaster1_p & v3a67577 | !hmaster1_p & v3a59746;
assign v3723ee4 = hmaster0_p & v37245f8 | !hmaster0_p & bddd83;
assign v3a6f9e9 = hbusreq8 & v373158e | !hbusreq8 & v376b3d4;
assign v373e6cf = hbusreq4 & v3728d72 | !hbusreq4 & v3a70a88;
assign v3746e30 = hbusreq7_p & v372dc20 | !hbusreq7_p & v3768e37;
assign v3a5d6e3 = hmaster1_p & v37693fe | !hmaster1_p & v3a70365;
assign v377209b = hmaster1_p & v8455ab | !hmaster1_p & cceefd;
assign v372e74c = hmaster1_p & v375ba66 | !hmaster1_p & bfae74;
assign v376bd96 = hmaster1_p & v3a6ffb6 | !hmaster1_p & v3a683d9;
assign v377e345 = hmaster0_p & v372cacb | !hmaster0_p & v376a6f1;
assign v373f6cf = hmaster0_p & v3a635ea | !hmaster0_p & v374b285;
assign v3a6ef2e = hbusreq4 & v377d86e | !hbusreq4 & !v8455ab;
assign v375159d = hmaster2_p & v374b887 | !hmaster2_p & v3a54b46;
assign v372e8ed = hgrant1_p & v3747302 | !hgrant1_p & !v35772a5;
assign v3a6862e = hbusreq7 & v3755c3f | !hbusreq7 & v3774bad;
assign v372b2cb = hgrant8_p & v3a712a1 | !hgrant8_p & v373812a;
assign v3a6fff7 = hgrant3_p & v37331e7 | !hgrant3_p & v377ae65;
assign a2aef9 = hmaster0_p & v3a6f490 | !hmaster0_p & v374dfd5;
assign v375d23b = hmaster1_p & v3a637dc | !hmaster1_p & v37300ba;
assign v3764b0a = hbusreq0 & v3a7107a | !hbusreq0 & !v8455ab;
assign v377682b = hmaster0_p & v372bae3 | !hmaster0_p & v3a5f992;
assign v377e31d = hbusreq7 & v37499ac | !hbusreq7 & v375c8db;
assign v3a5e8ac = hbusreq8 & v3a67d7b | !hbusreq8 & v3a60276;
assign v3a6fe58 = hbusreq2_p & v3a5fc3c | !hbusreq2_p & v3763acf;
assign v3753d94 = hgrant4_p & v377bfc0 | !hgrant4_p & v373f3b5;
assign v3733249 = hbusreq7_p & v37264a3 | !hbusreq7_p & v3749e61;
assign v3577324 = hmaster0_p & v375725f | !hmaster0_p & !v8455ab;
assign v3a551f9 = hbusreq4 & v3759031 | !hbusreq4 & v8455ab;
assign v3a63fc5 = hbusreq4 & v3a649fd | !hbusreq4 & v3755abd;
assign v380a170 = hmaster0_p & v3778ecc | !hmaster0_p & v3a6ef24;
assign v3759ca5 = stateA1_p & v8455ab | !stateA1_p & v3739e55;
assign v3a69714 = hmaster1_p & v3751dd2 | !hmaster1_p & v3778aac;
assign v3a67b93 = hlock5_p & v3747192 | !hlock5_p & v3a70b15;
assign v37369e4 = hbusreq2_p & v3a5eeb4 | !hbusreq2_p & v377bb62;
assign v3a5ef0c = hburst0 & v35b9d52 | !hburst0 & v1e37a34;
assign v3a70fd6 = hmaster2_p & v8455ab | !hmaster2_p & v3745bc4;
assign v375f848 = hgrant5_p & v3727d4c | !hgrant5_p & !v8455ab;
assign v37445e2 = hmaster0_p & v3a61cd7 | !hmaster0_p & v3a6d48a;
assign v376634c = hmaster0_p & v3a650e9 | !hmaster0_p & v3732931;
assign v3a70f51 = hmaster0_p & v2aca977 | !hmaster0_p & v3a56a2c;
assign v3736779 = hlock8 & v3a715cb | !hlock8 & v374d246;
assign v3a67ff8 = hbusreq0 & v9aea50 | !hbusreq0 & v37654b9;
assign v3a6f018 = hburst1 & v3a6ab5f | !hburst1 & v377314f;
assign v3a70ecc = hbusreq8 & v3762116 | !hbusreq8 & v8455ab;
assign v3754a0d = hmaster1_p & v37666f6 | !hmaster1_p & v3770653;
assign ce8abd = hmaster1_p & v372b8a3 | !hmaster1_p & v377195f;
assign v3751a97 = hmaster2_p & v3a635ea | !hmaster2_p & v3a7024f;
assign v3a70a25 = hmaster0_p & v3a70ca8 | !hmaster0_p & v372bc50;
assign v3740541 = hmaster2_p & v375121b | !hmaster2_p & !v377d9aa;
assign v3a583f5 = hbusreq3 & v37735ec | !hbusreq3 & v3749b84;
assign v3a5a03f = hbusreq4_p & v374ebb0 | !hbusreq4_p & v3770116;
assign v2ff9397 = hmaster1_p & v3a5db7f | !hmaster1_p & v23fe052;
assign v376db27 = hmaster2_p & v3744b55 | !hmaster2_p & v374d057;
assign v37656c1 = hmaster2_p & v3771c59 | !hmaster2_p & !v373b5f0;
assign v3a71204 = hgrant5_p & v3a57139 | !hgrant5_p & v37426bf;
assign v372f100 = hgrant4_p & v3758166 | !hgrant4_p & v3735a7c;
assign v374d726 = hgrant5_p & v3758fc4 | !hgrant5_p & v3771ad8;
assign v35b70d2 = jx0_p & v3728389 | !jx0_p & v3725088;
assign v3a65245 = hgrant0_p & v8455ab | !hgrant0_p & v377f190;
assign v3740f89 = jx0_p & v3a675b9 | !jx0_p & v3770b33;
assign v360c3d7 = hlock6_p & v37282cf | !hlock6_p & v8455ab;
assign v376eea3 = hgrant4_p & v3a5ee62 | !hgrant4_p & v375e527;
assign v3778032 = hbusreq7_p & v3741759 | !hbusreq7_p & v3a71214;
assign v3a5690e = hbusreq4_p & v3741aca | !hbusreq4_p & v8455ab;
assign v37318cb = hbusreq8_p & v3a702f9 | !hbusreq8_p & v3a5fa09;
assign v37427d3 = hgrant0_p & v3a635ea | !hgrant0_p & a22759;
assign v3742ca7 = hmaster0_p & v3a66c5b | !hmaster0_p & v3767e71;
assign v376cfc9 = hbusreq8 & v376079d | !hbusreq8 & v3a6fcf5;
assign v372a831 = hgrant2_p & v3807f45 | !hgrant2_p & v3741e80;
assign v3a638f4 = hgrant5_p & v37535fd | !hgrant5_p & v37529f6;
assign v37464f0 = hgrant3_p & v3a653e4 | !hgrant3_p & !v37346be;
assign v373ee8b = hmaster3_p & v8455ab | !hmaster3_p & !v3739ddd;
assign v3a6c3ac = hmaster1_p & v376a4ec | !hmaster1_p & v3778c14;
assign v3a6f3b9 = hmaster2_p & v374465a | !hmaster2_p & v376be50;
assign v376b81b = hgrant4_p & v3a61603 | !hgrant4_p & v373d136;
assign v3a64f97 = hbusreq6_p & v3a6e0f2 | !hbusreq6_p & v373d848;
assign v3a707ff = jx1_p & v8455ab | !jx1_p & v375579f;
assign v380909e = hmaster2_p & v3747302 | !hmaster2_p & v3a6eb7b;
assign v3a6ef34 = hbusreq4 & v3744fc9 | !hbusreq4 & v8455ab;
assign v376eb57 = hmaster1_p & v37388aa | !hmaster1_p & v3753976;
assign v373d49c = hmaster1_p & v37570f8 | !hmaster1_p & v3748b15;
assign v87cef3 = hgrant6_p & v37414b0 | !hgrant6_p & v374815b;
assign v3749c91 = hgrant2_p & v3a6eb39 | !hgrant2_p & !v3a70ff9;
assign v37567c7 = hlock1 & v37722cc | !hlock1 & v3a706c0;
assign v3734b14 = hmaster0_p & v3a5e24e | !hmaster0_p & v3a6f8c9;
assign v375c917 = hbusreq0 & v3a6ff37 | !hbusreq0 & v375a0ec;
assign v377ecec = hlock7_p & v3765aa0 | !hlock7_p & v3a5c1e7;
assign v377109d = hgrant3_p & v3a6251b | !hgrant3_p & v37675e2;
assign v3a63fbc = hbusreq7 & v3765978 | !hbusreq7 & v3a715a4;
assign v3a59609 = hmaster2_p & v3a5fe2f | !hmaster2_p & v372ce98;
assign v3a568e8 = hmaster2_p & v3a6fd81 | !hmaster2_p & v3a621cb;
assign bb0568 = hlock5_p & v3a53ae0 | !hlock5_p & v3a7121a;
assign v3769981 = hgrant6_p & v8455ab | !hgrant6_p & v3735f02;
assign v374d9c0 = hmaster0_p & v8455ab | !hmaster0_p & v3740951;
assign v3769db7 = hbusreq7_p & v37723ed | !hbusreq7_p & !v3a62f72;
assign v37485df = hbusreq5 & v376af8c | !hbusreq5 & v8455ab;
assign v3733716 = hbusreq4 & v3a5b885 | !hbusreq4 & v3809ec3;
assign v37647ce = hbusreq0 & v373d032 | !hbusreq0 & v8455ab;
assign v35b8d36 = hbusreq2_p & v3a5891c | !hbusreq2_p & !v39a537f;
assign v377c9c3 = hbusreq8_p & v37387e6 | !hbusreq8_p & v3a6b22e;
assign v39a4e19 = hmaster1_p & v37757cb | !hmaster1_p & v373ba38;
assign v37797f4 = hmaster1_p & v3a6f563 | !hmaster1_p & !v3a5cf3c;
assign v37435eb = hmaster2_p & v37330dc | !hmaster2_p & v3a6eb7b;
assign v3a7018a = hlock0 & v372b5a3 | !hlock0 & v3a7151e;
assign v3769a60 = hbusreq5 & v3774937 | !hbusreq5 & v8455bb;
assign v3a5a4c0 = hbusreq8 & v3a70b62 | !hbusreq8 & v3760617;
assign v377b679 = jx1_p & v3763188 | !jx1_p & v3a5842b;
assign v373dfb8 = hbusreq3 & v376f332 | !hbusreq3 & v3735525;
assign v375049a = hmaster2_p & v3a635ea | !hmaster2_p & v374db6a;
assign v3738b8a = hmaster2_p & v8455ab | !hmaster2_p & v8455be;
assign v3771fbb = hbusreq4_p & v3774075 | !hbusreq4_p & v375c917;
assign v376d3f7 = hbusreq3_p & v375ad91 | !hbusreq3_p & v3768428;
assign v373006f = hready & v37386f2 | !hready & v3739bfa;
assign v97ea11 = hbusreq5_p & v376a87f | !hbusreq5_p & v375ac16;
assign v3a6706d = hgrant5_p & v8455b9 | !hgrant5_p & v3728a9f;
assign v372cae4 = hgrant5_p & v3765e47 | !hgrant5_p & v3747b74;
assign v3a5ddd4 = hgrant1_p & v3a5bf04 | !hgrant1_p & v1e38224;
assign v3751a4f = hgrant8_p & v8455c1 | !hgrant8_p & v3725872;
assign v3766dc8 = hmaster1_p & v3807aa1 | !hmaster1_p & v3a584fd;
assign v3a706f6 = hmaster0_p & v3769c47 | !hmaster0_p & v3759007;
assign v376a3fe = hgrant4_p & v3733170 | !hgrant4_p & v374a580;
assign v374e9d1 = hbusreq8 & v3732a31 | !hbusreq8 & v3773f27;
assign v3771e26 = hbusreq8 & v372f5ca | !hbusreq8 & v373b837;
assign v3779da3 = hbusreq5_p & v98068b | !hbusreq5_p & v373eadd;
assign v3a702a8 = hgrant6_p & v8455c9 | !hgrant6_p & v3762f98;
assign v373ebd2 = hmaster1_p & v376a31b | !hmaster1_p & v377da1e;
assign v3a70b9b = hmaster1_p & v372e967 | !hmaster1_p & v8455ab;
assign v376086c = hmaster0_p & v3743966 | !hmaster0_p & v376d21d;
assign v3750269 = hbusreq2_p & v372b790 | !hbusreq2_p & v372c503;
assign v372f5bd = hbusreq2_p & v3727ce4 | !hbusreq2_p & v23fe376;
assign v372a4c1 = hgrant6_p & v3771ea7 | !hgrant6_p & v2aca977;
assign v3806c41 = hlock2 & v3751c4b | !hlock2 & v373c01b;
assign b254e2 = hbusreq1_p & v360d1ca | !hbusreq1_p & v376f6d1;
assign v3742c68 = hmaster0_p & v3771076 | !hmaster0_p & v3a5a9e6;
assign v37712e5 = hmaster1_p & v374fac9 | !hmaster1_p & v375d1d4;
assign v3747ad5 = hbusreq4_p & v3739ea3 | !hbusreq4_p & v8455ab;
assign v3729f7b = hbusreq5 & v3a6a8c0 | !hbusreq5 & v3769740;
assign v3775fb0 = hbusreq6 & v377c38c | !hbusreq6 & v8455ab;
assign v3a6feaa = hbusreq2_p & v374047a | !hbusreq2_p & v3a6d156;
assign v3a68c87 = hbusreq7 & v373149a | !hbusreq7 & v374312f;
assign v376132a = hmaster2_p & v3a70230 | !hmaster2_p & v372f346;
assign v375e7aa = hbusreq6 & v3a6f431 | !hbusreq6 & v8455ab;
assign v35b91b6 = hbusreq0_p & v3757aa1 | !hbusreq0_p & v8455b5;
assign v1e37489 = hgrant4_p & v8455ab | !hgrant4_p & !v1e38241;
assign v376b4a8 = hgrant2_p & v376e04c | !hgrant2_p & v37c00b6;
assign v3743ecf = hlock5 & v376fc09 | !hlock5 & v3806def;
assign bca64b = hmaster1_p & v3a700d9 | !hmaster1_p & v3728dd0;
assign v3722b74 = hbusreq3 & v373997b | !hbusreq3 & v35b774b;
assign v3730b57 = hbusreq5 & v3a6ffca | !hbusreq5 & v8455ab;
assign v3759158 = hbusreq1_p & v375c3b0 | !hbusreq1_p & !v3a5bbed;
assign v3729113 = hbusreq8_p & v3763c1f | !hbusreq8_p & v376f583;
assign v3a6fcd1 = stateG10_1_p & v3733b65 | !stateG10_1_p & b33e26;
assign v3a56855 = hmaster1_p & v3806847 | !hmaster1_p & v375b320;
assign v3755731 = hmaster0_p & v3a61c1f | !hmaster0_p & v3a71202;
assign v3a6b73c = hmaster2_p & v372f151 | !hmaster2_p & v3a5d4d0;
assign v3a5a5c8 = hbusreq5_p & v3756bde | !hbusreq5_p & v3a6d9a6;
assign v375a0a1 = hbusreq6 & v3752e63 | !hbusreq6 & v3a70d99;
assign v377b170 = hmaster1_p & v8455ab | !hmaster1_p & v3753328;
assign v380731d = hbusreq7_p & v8455ab | !hbusreq7_p & v372cdde;
assign v3779f13 = hgrant2_p & v37320bb | !hgrant2_p & v372fc77;
assign v23fdbdc = hgrant0_p & v375a268 | !hgrant0_p & v3a65161;
assign v3723493 = hgrant2_p & v3723b00 | !hgrant2_p & v3a5e81d;
assign v3747a97 = hbusreq0 & v37343dc | !hbusreq0 & v8455ab;
assign v373b710 = hbusreq1_p & v3a70c73 | !hbusreq1_p & !v3a53cc3;
assign v372dde7 = hlock4 & v37487f7 | !hlock4 & v3a58674;
assign v376ae39 = hlock8_p & v3777474 | !hlock8_p & !v3735aa5;
assign v3726521 = hmaster0_p & v374f658 | !hmaster0_p & v3763a4a;
assign v3749ca6 = hmaster1_p & v373a327 | !hmaster1_p & v8455ab;
assign v3809de2 = hlock2 & v3a63a2a | !hlock2 & v3a5610f;
assign v3a67e97 = hbusreq5_p & v37509f2 | !hbusreq5_p & !v37796c3;
assign v8455e7 = locked_p & v8455ab | !locked_p & !v8455ab;
assign v3741dce = hbusreq3_p & v376b33c | !hbusreq3_p & v372a0bd;
assign v37773a2 = hlock3 & d2819e | !hlock3 & v3752bcc;
assign v3760989 = hmaster1_p & v8455ab | !hmaster1_p & v3a617ad;
assign v37404b3 = hgrant6_p & v3a53fa4 | !hgrant6_p & v375f98c;
assign v3739336 = hlock2_p & v3727eb8 | !hlock2_p & v8455bf;
assign v3741f39 = hgrant2_p & v3a62524 | !hgrant2_p & v3a56f66;
assign v37313b6 = hgrant3_p & v8455ab | !hgrant3_p & v376b0d6;
assign v3a697d2 = hmaster0_p & v376a907 | !hmaster0_p & v3a70574;
assign v39eb517 = hgrant0_p & v3a653e4 | !hgrant0_p & !v3750d06;
assign v37519ea = hgrant6_p & v3a708c2 | !hgrant6_p & v375de7f;
assign v376ea64 = hmaster2_p & v3a6935c | !hmaster2_p & v3730b6c;
assign v3a715e6 = hbusreq7_p & v3a53d2b | !hbusreq7_p & v3759232;
assign v373ed37 = jx0_p & v374a9cd | !jx0_p & v8455ab;
assign v3a70230 = hbusreq4_p & v3a67cff | !hbusreq4_p & v373b7c5;
assign v3a58016 = hbusreq5 & v375ff00 | !hbusreq5 & v3777c0c;
assign v3760860 = jx3_p & v3a59d00 | !jx3_p & v3a6ffb1;
assign v3760933 = hbusreq3 & v376495e | !hbusreq3 & v8455ab;
assign v3a6f1c6 = hlock1_p & v3a29803 | !hlock1_p & !v8455ab;
assign v3a6fb28 = hbusreq5_p & v3a66732 | !hbusreq5_p & v375caa0;
assign v2092f0f = hmaster2_p & v3a5f6d5 | !hmaster2_p & v3a66a01;
assign v372bbc7 = hmaster1_p & v3729189 | !hmaster1_p & v3740bf5;
assign v3a610f8 = hmaster2_p & v3a5cd4c | !hmaster2_p & v3a63bb7;
assign v3a5d08e = hbusreq0 & v3730c0a | !hbusreq0 & v3762e66;
assign v3a6fc0f = hmaster0_p & v37644ce | !hmaster0_p & v3379430;
assign v372aec7 = hmaster2_p & v3a635ea | !hmaster2_p & v3a70172;
assign v37398ac = hbusreq5 & v375f90e | !hbusreq5 & v3a59dd6;
assign v33790e7 = hgrant2_p & v8df61b | !hgrant2_p & v375d161;
assign v37470e6 = hmaster0_p & v377234d | !hmaster0_p & v8455e7;
assign v372935c = hbusreq1_p & v3a70c07 | !hbusreq1_p & v1e38224;
assign v37270dc = hlock5 & v3a6ab14 | !hlock5 & v37647fc;
assign v373b4dc = hbusreq5 & v37480b7 | !hbusreq5 & !v37358ab;
assign v372f770 = hmaster0_p & v3a5755b | !hmaster0_p & v3a710d0;
assign v3809542 = hmaster0_p & v376438f | !hmaster0_p & v3a7114b;
assign v37664b4 = hlock8 & v376f42c | !hlock8 & v376c8f2;
assign v3808d2f = hlock7_p & v3a5fdc8 | !hlock7_p & !v8455ab;
assign v3739cdb = hbusreq8_p & v373ab2b | !hbusreq8_p & v3777d70;
assign v374bd2c = hmaster2_p & v372647d | !hmaster2_p & v375bfdf;
assign v376c322 = hmaster1_p & v3731dc1 | !hmaster1_p & v376ca02;
assign v3a63408 = hgrant4_p & v374a99e | !hgrant4_p & v8455ab;
assign v3769559 = hmaster1_p & v37610ae | !hmaster1_p & v3757b39;
assign v23fdec8 = hbusreq5 & v3a70927 | !hbusreq5 & v3a700c8;
assign v373351d = hbusreq6_p & v376fdd6 | !hbusreq6_p & !v8455ab;
assign v376eed1 = hmaster0_p & v3a619c0 | !hmaster0_p & v3a70d3a;
assign v373f28d = hlock8 & v37680b5 | !hlock8 & v3a56570;
assign v3763a12 = hmaster1_p & v3a70cf1 | !hmaster1_p & v37412e9;
assign v3a6595f = hgrant4_p & v3a7133d | !hgrant4_p & v373bb50;
assign v372d691 = hlock8 & v376ae9f | !hlock8 & v377bd76;
assign v38073ff = hmaster1_p & v8455e7 | !hmaster1_p & bf6c15;
assign v377f0e7 = jx3_p & v377f7dd | !jx3_p & v3a7039c;
assign v3a614fe = hmaster0_p & v3807ae8 | !hmaster0_p & v3a6c605;
assign v3a70583 = hgrant8_p & v3a5ba5b | !hgrant8_p & v37646dc;
assign v3750d8e = hmaster0_p & v3746c51 | !hmaster0_p & v374a075;
assign v3757490 = hbusreq5_p & v3773201 | !hbusreq5_p & !v8455ab;
assign v3a69b74 = hgrant4_p & v8455ab | !hgrant4_p & v3a61ecf;
assign v374c6c5 = hbusreq8 & v3740663 | !hbusreq8 & !v3743b62;
assign v377834b = hbusreq3_p & v37694de | !hbusreq3_p & v8455ab;
assign v3a6aaa4 = hmaster1_p & v3a6961d | !hmaster1_p & v372fbb1;
assign v375380a = hbusreq4_p & v376cedc | !hbusreq4_p & !v8455ab;
assign v3766246 = hbusreq7_p & v3734279 | !hbusreq7_p & v373f28d;
assign v3a70485 = hbusreq7_p & v3730cb5 | !hbusreq7_p & !v8455ab;
assign v372ad1d = hbusreq2 & v374bf71 | !hbusreq2 & v8455ab;
assign v377f149 = hbusreq3 & v3a6c0b3 | !hbusreq3 & v3a7162d;
assign v373e8cb = hmaster0_p & v3733a1a | !hmaster0_p & v373a3c8;
assign v3734f04 = hgrant4_p & v376ab5d | !hgrant4_p & v376beaa;
assign v3a5a2e5 = hbusreq8 & v3a5509a | !hbusreq8 & v3736f6d;
assign v3a6e584 = hmaster2_p & v376c176 | !hmaster2_p & v8455e7;
assign v373261a = hgrant2_p & v373dbb0 | !hgrant2_p & !v3a61298;
assign v37468ea = hbusreq3_p & v3a635ea | !hbusreq3_p & v3a7139e;
assign v3757a13 = hgrant2_p & v3770559 | !hgrant2_p & v38063c7;
assign v3a6e2ce = jx1_p & v3a70aa8 | !jx1_p & v3774253;
assign v3a6a52c = hlock7 & v3732b30 | !hlock7 & v3761f69;
assign v1e3799d = hlock4 & v374e43a | !hlock4 & v3a61901;
assign v3a60fee = hbusreq5 & v3767797 | !hbusreq5 & v3a6f47a;
assign v37547ad = hlock6_p & v3a710c6 | !hlock6_p & v8455bb;
assign v3a711c8 = hgrant5_p & v372fef2 | !hgrant5_p & v3772612;
assign v3749412 = hgrant5_p & v8455ab | !hgrant5_p & !v8455f1;
assign v1e37407 = hmaster0_p & v375e944 | !hmaster0_p & v374e0f6;
assign v3763186 = hbusreq4 & v3768870 | !hbusreq4 & v38072fd;
assign v374b2c2 = hlock7_p & v373eeec | !hlock7_p & v3734810;
assign v37302a2 = hbusreq5_p & v377f3ae | !hbusreq5_p & v8455ab;
assign v374197c = hbusreq1 & v3a70c94 | !hbusreq1 & v3a635ea;
assign v3a57e1a = hbusreq8 & v3a695f1 | !hbusreq8 & v8455bf;
assign v3a6946d = hbusreq0_p & v37787ec | !hbusreq0_p & v374cc2a;
assign v3379037 = locked_p & v3a70a83 | !locked_p & v39a5381;
assign v3a59b5c = hbusreq3 & v3a715d2 | !hbusreq3 & v8455ab;
assign v3762ea7 = hbusreq0 & v373064e | !hbusreq0 & v8455ab;
assign v37383f6 = hgrant3_p & v3735809 | !hgrant3_p & v3a70b3a;
assign v373de1d = hbusreq8 & v3767be8 | !hbusreq8 & v3768734;
assign v3a62465 = hlock6 & v3733f37 | !hlock6 & v3a6eb8b;
assign v3a70168 = hlock0 & v3a6eb47 | !hlock0 & v3737d3f;
assign v3a6fac6 = hgrant6_p & v3a706b7 | !hgrant6_p & v3a70a05;
assign v374c2d6 = hmaster1_p & v373a4e4 | !hmaster1_p & v38070c7;
assign v3766ea9 = hgrant3_p & v3258d68 | !hgrant3_p & v37757e0;
assign v373d262 = hbusreq4 & v3a66a3b | !hbusreq4 & v8455ab;
assign v372f349 = hbusreq4_p & v373be25 | !hbusreq4_p & !v372935c;
assign v373e524 = hlock2_p & v3737e21 | !hlock2_p & v3731945;
assign v3740f78 = hmaster1_p & v3a6e31f | !hmaster1_p & v373ad86;
assign v373359b = hmaster2_p & v372fc81 | !hmaster2_p & !v376f2f8;
assign v374d741 = hmaster1_p & v3a67d66 | !hmaster1_p & v372dfc3;
assign v375fe5b = hbusreq6 & v37280b0 | !hbusreq6 & v3a6da8a;
assign v360d0fb = hmaster1_p & v37684b7 | !hmaster1_p & v374c8b8;
assign v3a70888 = hgrant0_p & v8455ab | !hgrant0_p & v37788ca;
assign v3777527 = hbusreq5_p & v372fa9d | !hbusreq5_p & v3758466;
assign v3762e16 = hmaster0_p & v3a70d99 | !hmaster0_p & v3775cb7;
assign v3722d9b = hgrant4_p & v8455ab | !hgrant4_p & v3a7164a;
assign v372c20d = hbusreq7 & v3a706ea | !hbusreq7 & v3a671f2;
assign v3809112 = hbusreq0 & v372fb60 | !hbusreq0 & v373e814;
assign v3a701cd = hgrant3_p & v372aacd | !hgrant3_p & !v3808d42;
assign v3a5c6d0 = hgrant4_p & v3775dbc | !hgrant4_p & v3a568e4;
assign v375caa2 = hmaster1_p & v3a70ccd | !hmaster1_p & v374e21e;
assign v3a7007e = hmaster2_p & v8455ab | !hmaster2_p & !v3a587f6;
assign v3a62041 = hgrant2_p & v37321b8 | !hgrant2_p & v3a68e39;
assign v38068c8 = hmaster2_p & v3a70b92 | !hmaster2_p & v3779cf9;
assign v3a5666f = hmaster1_p & v374851a | !hmaster1_p & v3a713da;
assign v372b4d7 = hbusreq2_p & v374c718 | !hbusreq2_p & v3766df9;
assign v3a6d6ff = hlock5_p & v375243f | !hlock5_p & v8455b7;
assign v37444d0 = stateG2_p & v8455ab | !stateG2_p & !v3759020;
assign v3a71286 = hmaster3_p & v3756fd9 | !hmaster3_p & v373714f;
assign v377cd7a = hbusreq3_p & v3763a20 | !hbusreq3_p & !v8455ab;
assign v3a5de50 = hbusreq2 & v377b8ee | !hbusreq2 & v8455ab;
assign v373bcea = hbusreq6 & v3742adb | !hbusreq6 & v8455ab;
assign v3a5a23b = hmaster1_p & v374729b | !hmaster1_p & v3761c19;
assign v377cc23 = hbusreq3 & v3a6abaa | !hbusreq3 & v37427d3;
assign v3757b55 = hgrant6_p & v3760e2e | !hgrant6_p & v3a6b710;
assign v3758b56 = hlock7 & v3773a96 | !hlock7 & v37655bf;
assign v37336f0 = hbusreq2 & v3a7036a | !hbusreq2 & v8455ab;
assign v3745e12 = hgrant5_p & v3755066 | !hgrant5_p & v3256555;
assign v3a62070 = hgrant6_p & v373b209 | !hgrant6_p & v3a70504;
assign v3773a3d = hmastlock_p & v3a648f2 | !hmastlock_p & !v8455ab;
assign v337904a = hbusreq8 & v37532a8 | !hbusreq8 & v376d9f3;
assign v1e37932 = hbusreq2 & v3a70641 | !hbusreq2 & v8455ab;
assign v3a6f974 = hbusreq5_p & v8455ab | !hbusreq5_p & v3743a77;
assign v3755db9 = jx0_p & v3a5f4ef | !jx0_p & v3a6f063;
assign v373ebf9 = hbusreq4_p & v372372d | !hbusreq4_p & v3a55b1d;
assign v3a6f8f7 = hbusreq4 & v3729e32 | !hbusreq4 & v37519ea;
assign v3a60247 = hbusreq5_p & v3a59529 | !hbusreq5_p & v3a6e986;
assign v37352a5 = hbusreq6 & v372e6f4 | !hbusreq6 & v3a6687c;
assign v3806507 = hlock1 & v37306bb | !hlock1 & v3a63621;
assign v3a6effc = hmaster2_p & v3747d68 | !hmaster2_p & v3767848;
assign v373015f = hgrant4_p & v374d6b2 | !hgrant4_p & v3766ddb;
assign v3a71214 = hgrant5_p & v376139f | !hgrant5_p & v3a70d19;
assign v37335ff = hmaster0_p & v374f31d | !hmaster0_p & v373c545;
assign v3a613f2 = hbusreq5_p & v3775610 | !hbusreq5_p & v3a701ce;
assign v3726e7b = hgrant5_p & v374248e | !hgrant5_p & v375bca7;
assign v376abcc = hbusreq7 & v2092b5f | !hbusreq7 & a0a219;
assign v3a69515 = hbusreq1_p & c60044 | !hbusreq1_p & !v8455ab;
assign v376ba63 = hmaster1_p & v3764f5c | !hmaster1_p & v373cc9a;
assign v3a60195 = hmaster2_p & v3a64d7c | !hmaster2_p & v3725578;
assign v372ff54 = hmaster2_p & v3769ecf | !hmaster2_p & v3748d67;
assign v3a698ed = hmaster0_p & v375c3f6 | !hmaster0_p & !v377de50;
assign v38097ae = hmaster0_p & v374729b | !hmaster0_p & v373c5dc;
assign v373a841 = hbusreq1_p & v8455ab | !hbusreq1_p & v37665bf;
assign v3a6ad93 = hmaster0_p & v3738253 | !hmaster0_p & ba83e3;
assign v373e16a = stateG10_1_p & v3a70ecf | !stateG10_1_p & v3a6eb77;
assign v372b1e8 = hbusreq7_p & v3749975 | !hbusreq7_p & !v3a56e45;
assign v95d97e = hburst1 & v372b0cd | !hburst1 & v372ef9b;
assign v3a6c68c = hbusreq4 & v374e35e | !hbusreq4 & v8455ab;
assign v3a70f5e = hbusreq4_p & v3766d10 | !hbusreq4_p & !v8455ab;
assign v376c6b3 = hlock7 & v372d28d | !hlock7 & v3742a4e;
assign v377e031 = hbusreq8 & v3a5e998 | !hbusreq8 & v8455ab;
assign v3a5459f = hmaster0_p & v3a6d574 | !hmaster0_p & !v372a696;
assign v372a27f = hbusreq5 & v3738279 | !hbusreq5 & v8455ab;
assign v372aadd = hbusreq6_p & v3768985 | !hbusreq6_p & v3727369;
assign v373554b = hgrant6_p & v3a53da1 | !hgrant6_p & !v3a6ef50;
assign v3a5788f = hbusreq2 & v8455ab | !hbusreq2 & v373a391;
assign v37c006d = hbusreq4 & v374d751 | !hbusreq4 & v3a6fdc7;
assign v3a70272 = hlock0_p & v3759032 | !hlock0_p & v372d943;
assign v3762a49 = hgrant4_p & v37300a5 | !hgrant4_p & v3a584f1;
assign v374059d = hlock0_p & v3a707de | !hlock0_p & v3736c94;
assign v3748d63 = hlock5 & v37551b2 | !hlock5 & v3772bb1;
assign v3738a70 = hmaster1_p & v3a65b79 | !hmaster1_p & v3757044;
assign v3a6519c = jx1_p & v8455d1 | !jx1_p & v3723fb3;
assign v375a513 = hmaster1_p & v374314f | !hmaster1_p & v3a7130b;
assign v374e663 = hbusreq5_p & v3a70f68 | !hbusreq5_p & v377f734;
assign v3807a26 = hmaster2_p & v377a002 | !hmaster2_p & bbcc5e;
assign v375070c = hbusreq2_p & v3746feb | !hbusreq2_p & v8455ab;
assign v377e9a4 = hlock2_p & v35772b3 | !hlock2_p & v35772a6;
assign v3770da3 = hmaster2_p & v3a712c4 | !hmaster2_p & v3754403;
assign v3a70f7f = hgrant4_p & v377e57f | !hgrant4_p & v37788fc;
assign v3a70596 = hmaster2_p & v3740171 | !hmaster2_p & v37395e6;
assign v372690e = hbusreq5_p & v3a71097 | !hbusreq5_p & !v8455ab;
assign v3a6c573 = hbusreq5_p & v3749993 | !hbusreq5_p & v360d0a9;
assign v3779955 = jx1_p & v37624a9 | !jx1_p & v373c15e;
assign v3a56d2d = hbusreq0 & v325b5df | !hbusreq0 & v37648f2;
assign c7ae7d = hmaster0_p & v375e993 | !hmaster0_p & v8455ab;
assign v3a6eac2 = hlock8_p & v3750ac3 | !hlock8_p & !v3a5a23b;
assign v3a70407 = hmaster2_p & v8455ab | !hmaster2_p & v373a841;
assign v3767650 = hbusreq0 & v373343b | !hbusreq0 & v376011a;
assign v3735436 = hbusreq3 & v3a6fdb4 | !hbusreq3 & v372cc25;
assign d54152 = hmaster2_p & v3a702a2 | !hmaster2_p & v3762502;
assign v2ff9229 = hbusreq5_p & v3a29850 | !hbusreq5_p & v3a71276;
assign v3a676d6 = locked_p & v3a5d74e | !locked_p & !v8455ab;
assign v3a5bc76 = hlock7 & v3762230 | !hlock7 & v374705f;
assign v373b9e9 = hbusreq8_p & v3a714b7 | !hbusreq8_p & c8ca6f;
assign v3724dfb = jx1_p & v8455ab | !jx1_p & v23fdbe6;
assign v3778f32 = hbusreq8_p & v375b676 | !hbusreq8_p & v373c7af;
assign v3a5724f = hbusreq8 & v376e6e2 | !hbusreq8 & v8455ab;
assign v3777c39 = hgrant3_p & v375917f | !hgrant3_p & v375a250;
assign v3773d96 = hbusreq5_p & v3778419 | !hbusreq5_p & v376021d;
assign v3a7046a = hmaster3_p & v3733c70 | !hmaster3_p & v37674f2;
assign v374a877 = hgrant4_p & v8455ab | !hgrant4_p & v37396de;
assign v3a69b5c = hgrant2_p & v37511c0 | !hgrant2_p & v3a6eeca;
assign v23fda6a = hbusreq2 & v37564e4 | !hbusreq2 & !v8455bd;
assign v3753fe3 = hbusreq7 & v37750a5 | !hbusreq7 & v3723025;
assign v374d246 = hlock7 & v3734279 | !hlock7 & v3a67715;
assign v3769f4a = hlock1 & v3748797 | !hlock1 & v3727507;
assign v377d8eb = hbusreq2_p & v374c718 | !hbusreq2_p & v375978a;
assign v376b438 = hmaster0_p & v3a713f2 | !hmaster0_p & v377b774;
assign v3772cf2 = hbusreq3 & v377ae65 | !hbusreq3 & v8455ab;
assign v372642b = hmaster1_p & v373823d | !hmaster1_p & v375993d;
assign v3727ec9 = hbusreq3 & v37299b3 | !hbusreq3 & v8455ab;
assign v3a6fd41 = hbusreq7 & v3a70577 | !hbusreq7 & v3a6fe04;
assign v3a6abcb = hmaster0_p & v3763175 | !hmaster0_p & v3764ec5;
assign v374e02b = jx0_p & v3734a96 | !jx0_p & v3a6a82d;
assign v375a463 = hbusreq4_p & v374f126 | !hbusreq4_p & v3a6f579;
assign v377b848 = hbusreq5_p & v375fcfa | !hbusreq5_p & v8455ab;
assign v374a3f3 = hbusreq6_p & v3742290 | !hbusreq6_p & v3a6687c;
assign v3764805 = hbusreq5_p & v3a70134 | !hbusreq5_p & v373c9c1;
assign v3a6c9c7 = hlock8_p & v37299ef | !hlock8_p & v8455ab;
assign v37231e5 = hmaster1_p & v374306c | !hmaster1_p & v37503bd;
assign v3a6f697 = hmaster1_p & v3a6eb67 | !hmaster1_p & v374e7fa;
assign v3a5cd50 = hbusreq3 & v3a59d9d | !hbusreq3 & v3762502;
assign v375145d = hmaster1_p & v3746487 | !hmaster1_p & v3a66335;
assign v3747c9f = hgrant7_p & v8455ce | !hgrant7_p & v372ad83;
assign v3a6094e = hmaster1_p & v3a6fe6f | !hmaster1_p & v374e21e;
assign v377a0e7 = hbusreq8_p & v3a7001c | !hbusreq8_p & v374fdc8;
assign v377ac0f = hmaster0_p & v3a619c0 | !hmaster0_p & v3a7031a;
assign v3a707d5 = hbusreq3 & v3a5952d | !hbusreq3 & v3a707c4;
assign v3a66606 = hbusreq6_p & v373d78b | !hbusreq6_p & v3a6fcb9;
assign v372b902 = hbusreq4_p & v3a701c7 | !hbusreq4_p & v375564e;
assign v3759fb9 = hbusreq5_p & v3765cd5 | !hbusreq5_p & v1e3737d;
assign v373ff40 = hbusreq7_p & v37249fe | !hbusreq7_p & v3758809;
assign v3725a38 = hlock7_p & v8455e7 | !hlock7_p & v374ac6d;
assign v3a707b9 = hbusreq5_p & v3750fee | !hbusreq5_p & v37512c1;
assign v3768739 = hlock5_p & v3a70ebc | !hlock5_p & v3a70077;
assign v3a6bf60 = hgrant2_p & v3809788 | !hgrant2_p & v37425a7;
assign v3722c80 = hgrant4_p & v3751081 | !hgrant4_p & v3733ae1;
assign v372b780 = hgrant4_p & v3744b1b | !hgrant4_p & v372b2ab;
assign v3a6f894 = hlock5 & v3736b4a | !hlock5 & v372ebd5;
assign v1e37c6e = hbusreq8_p & v3762cf7 | !hbusreq8_p & v3a59cde;
assign v373a0bf = locked_p & v374dd24 | !locked_p & !v8455ab;
assign v3728498 = hgrant2_p & v3a5b12c | !hgrant2_p & v375baed;
assign v3741bb2 = hlock0 & v3a67cff | !hlock0 & v3a63331;
assign v377d51d = hbusreq8_p & v37484e7 | !hbusreq8_p & v3a573ec;
assign v3759758 = hmaster1_p & v3727d4c | !hmaster1_p & v37617b9;
assign v3759dd9 = hlock3_p & v3737c0a | !hlock3_p & v377a4f1;
assign v3a68e0d = hbusreq8 & v8455ab | !hbusreq8 & v376e66e;
assign v37427e9 = hgrant4_p & v8455ab | !hgrant4_p & v3755420;
assign v3a70f2d = hlock5_p & v3a58182 | !hlock5_p & !v3728b31;
assign v375cb5e = hmaster2_p & v377b423 | !hmaster2_p & !v23fe339;
assign v375e566 = hbusreq7 & v3a5a01b | !hbusreq7 & v8455ab;
assign v37596de = hmaster0_p & v372dcfb | !hmaster0_p & v3a6230b;
assign v373f4fb = hbusreq4 & v3a6ab69 | !hbusreq4 & v374bc27;
assign v2acafaa = hmaster0_p & v3731fae | !hmaster0_p & v8455ab;
assign v374b9ee = hbusreq6_p & v3a6a489 | !hbusreq6_p & v3a6da8a;
assign v3a6f1e7 = hgrant4_p & v8455c1 | !hgrant4_p & v3776fb2;
assign v374bece = hmaster2_p & v374f9c6 | !hmaster2_p & v374db6a;
assign v377e568 = hbusreq8 & v3732f4d | !hbusreq8 & v8455ab;
assign v1e37d8e = hmaster2_p & v373c3e1 | !hmaster2_p & !v377b423;
assign v3a7022f = hmaster0_p & v3a635ea | !hmaster0_p & v37701af;
assign v372eada = hbusreq2 & v373d825 | !hbusreq2 & !v37507d0;
assign v3a708c6 = hbusreq4_p & v373aef5 | !hbusreq4_p & !v3a6f2b6;
assign v3754392 = hbusreq5 & v3a5a484 | !hbusreq5 & v8455ab;
assign v3a64f63 = hmaster0_p & v377c58e | !hmaster0_p & v3758ff0;
assign v3a6336e = hmaster2_p & v3a702c2 | !hmaster2_p & v3766202;
assign v37526a0 = hgrant3_p & v376f0c1 | !hgrant3_p & v375a613;
assign v3a7032b = hmaster1_p & v3a71203 | !hmaster1_p & v37698c3;
assign c63c1f = hbusreq5_p & v3752f9b | !hbusreq5_p & v377b429;
assign v377d9bb = hgrant6_p & v37285ad | !hgrant6_p & v3a6a051;
assign v372815e = hmaster0_p & v37640de | !hmaster0_p & !v375af99;
assign v3a67a41 = hgrant4_p & v377ddc1 | !hgrant4_p & !v3a5e96b;
assign v375ecf8 = hbusreq5 & v376a6f1 | !hbusreq5 & v3a5cc27;
assign v377a366 = hmaster2_p & v3738dac | !hmaster2_p & v8455ab;
assign v3a63f57 = hbusreq8_p & v3739e21 | !hbusreq8_p & v373046c;
assign v37471cb = hlock3_p & v3a71284 | !hlock3_p & v8455e7;
assign v373e209 = hbusreq2_p & v8455ab | !hbusreq2_p & v37665bf;
assign v3758fe4 = hbusreq6_p & v3a56338 | !hbusreq6_p & v2092b01;
assign v374d1b8 = hmaster1_p & v8455ab | !hmaster1_p & v3730526;
assign v37519d9 = hbusreq5_p & v374ff28 | !hbusreq5_p & v8455ab;
assign v3a6ee06 = hbusreq2 & v3a6dc08 | !hbusreq2 & v37406d2;
assign v3763d53 = hbusreq5 & v3a6826a | !hbusreq5 & v3a6edb5;
assign v374f7ec = hlock4 & v3765784 | !hlock4 & v3732797;
assign v3757fdd = hmaster3_p & v3778354 | !hmaster3_p & v3a70cd0;
assign v3a6cd4f = hbusreq7 & v37305e6 | !hbusreq7 & v375075b;
assign v3a6f30a = hmaster1_p & v3764219 | !hmaster1_p & v373823e;
assign v3726594 = hlock5_p & v3a5c945 | !hlock5_p & !v3777a8a;
assign v372da4f = hgrant3_p & v38099e8 | !hgrant3_p & v37609ac;
assign v3a70a57 = hbusreq5_p & v37280a0 | !hbusreq5_p & !v8455ab;
assign v37364bd = hlock5 & v375e767 | !hlock5 & v3a7086d;
assign v373cd41 = hlock4 & v376a464 | !hlock4 & v372e8cc;
assign v3a6eb01 = hgrant0_p & v3a56ccf | !hgrant0_p & v377c3fb;
assign v376e66e = hmaster1_p & v8455b0 | !hmaster1_p & v3a58c07;
assign v3733c7f = hbusreq8 & v3739915 | !hbusreq8 & v3a67beb;
assign v3729e5f = hbusreq6 & v375f317 | !hbusreq6 & v372781d;
assign v3a705d4 = hmaster0_p & v37282f7 | !hmaster0_p & v373a759;
assign v37621ff = hlock6 & v372495f | !hlock6 & v376d081;
assign v3769a1c = hmaster2_p & v375a94a | !hmaster2_p & v375bb92;
assign v375975b = hbusreq2_p & v8455ab | !hbusreq2_p & v3759512;
assign v37311de = hgrant2_p & v8455b9 | !hgrant2_p & v37265d6;
assign v376abd1 = jx3_p & v8455ab | !jx3_p & v3737ab4;
assign v375d067 = hbusreq4_p & v3a6d2df | !hbusreq4_p & v8455b0;
assign v3735a4f = hgrant2_p & v376cf8c | !hgrant2_p & v37240e8;
assign v372bc0c = hmaster0_p & be54b2 | !hmaster0_p & v3739774;
assign v374aa27 = hmaster0_p & v3739ab4 | !hmaster0_p & v3764d82;
assign v3757695 = hlock4 & v3743604 | !hlock4 & v3a6f751;
assign v3768622 = hbusreq4 & v375f98a | !hbusreq4 & v8455ab;
assign v373425d = hmaster0_p & v8455ab | !hmaster0_p & !v3a55454;
assign v37373ea = hbusreq3 & v3a54c77 | !hbusreq3 & v8455ab;
assign v3748665 = hlock3_p & v3a6b9e8 | !hlock3_p & v8455e7;
assign v372b679 = hmaster2_p & v374f307 | !hmaster2_p & v8455e7;
assign v3a54d59 = locked_p & v3a63043 | !locked_p & !v8455ab;
assign v3744752 = hbusreq3 & v376d9ad | !hbusreq3 & v8455e7;
assign v3a69329 = hmaster1_p & v3a6f224 | !hmaster1_p & v37558f2;
assign v3a70516 = hbusreq5_p & v3a55904 | !hbusreq5_p & v3752977;
assign v377e512 = hgrant6_p & v374510e | !hgrant6_p & v2889716;
assign v3723459 = hgrant5_p & v8455c6 | !hgrant5_p & b1fcb7;
assign v3a6ffa1 = hmaster0_p & v377d891 | !hmaster0_p & v3a5c026;
assign v3723fa6 = hbusreq7_p & v3a70c81 | !hbusreq7_p & v373c0b4;
assign v375783b = hmaster1_p & v3a6f7dd | !hmaster1_p & v38073b5;
assign v3a6f147 = hbusreq2 & v373014d | !hbusreq2 & v8455bf;
assign v375461f = hbusreq3_p & v3a5a41c | !hbusreq3_p & v8455ab;
assign v376fce9 = hmaster2_p & v1e382e7 | !hmaster2_p & v376d856;
assign v3a71018 = hgrant4_p & v3731c6f | !hgrant4_p & v3a6fcda;
assign v3733ba1 = hlock3 & v3724e67 | !hlock3 & v3a6fbfc;
assign v3756398 = hlock3 & v377cc23 | !hlock3 & v3a6abaa;
assign v3749e61 = hlock8 & v3a6e4b8 | !hlock8 & v3747587;
assign v3a6dcf5 = hmaster2_p & v37674f6 | !hmaster2_p & v3a711f9;
assign v37761cb = hbusreq6 & v37621ea | !hbusreq6 & v3760ff4;
assign v372b512 = hgrant2_p & v3732d55 | !hgrant2_p & v372b4d7;
assign v3a70c18 = jx0_p & cea42b | !jx0_p & v373fa33;
assign v3764530 = hmaster0_p & v373ee19 | !hmaster0_p & !v3a708a7;
assign v37288b6 = hbusreq3_p & v3a635ea | !hbusreq3_p & v3a5eafa;
assign v3771c6a = hbusreq8 & v3a6f92d | !hbusreq8 & v3768734;
assign v372deb9 = hbusreq7_p & v3754afa | !hbusreq7_p & v375145d;
assign v375b278 = hbusreq7 & v3737a21 | !hbusreq7 & !v37512f6;
assign v3a64032 = hbusreq5 & v3775c24 | !hbusreq5 & !v8455ab;
assign v3a70abe = hmaster2_p & v8455ab | !hmaster2_p & v3a70641;
assign v373191d = hmaster1_p & v3a65540 | !hmaster1_p & v3a69a50;
assign v3740a8a = hmaster1_p & v374306c | !hmaster1_p & v377de29;
assign v3774550 = hbusreq3_p & v3a705ad | !hbusreq3_p & !v37450cb;
assign v37637db = hgrant1_p & v3767abc | !hgrant1_p & v8455ab;
assign v3760a9d = stateG2_p & v8455ab | !stateG2_p & v3a70a28;
assign v3725269 = hmaster1_p & v3a6f173 | !hmaster1_p & v3763716;
assign v377429c = hmaster2_p & v3a70374 | !hmaster2_p & v377e889;
assign v3a7046c = hmaster0_p & v3a6fafe | !hmaster0_p & v3726991;
assign v377c32f = hbusreq6_p & v373fb30 | !hbusreq6_p & v3733dd3;
assign v3a64641 = hbusreq5_p & v376bfa7 | !hbusreq5_p & !v3a6f61c;
assign v3a5584b = hmaster0_p & v3a635ea | !hmaster0_p & v3769696;
assign v3a6f8fb = hbusreq4 & v3747994 | !hbusreq4 & v8455ab;
assign v374174c = hbusreq1 & v3a619c0 | !hbusreq1 & v8455ab;
assign v37470a5 = hbusreq8_p & v3a6ece9 | !hbusreq8_p & v377a5cc;
assign v3a56aae = hbusreq4_p & v3a56d78 | !hbusreq4_p & v3736c97;
assign v3a70859 = hbusreq5_p & v3758c13 | !hbusreq5_p & v3a66856;
assign v3737628 = hlock6 & v3a5de73 | !hlock6 & v3a6f2bf;
assign v3779002 = hlock4_p & v373eb4d | !hlock4_p & v3764c57;
assign v376f5b3 = hlock4 & v3744117 | !hlock4 & v3a6bf12;
assign v372feea = hbusreq5 & v3a66d47 | !hbusreq5 & v8455ab;
assign v374b080 = hmaster2_p & v3a635ea | !hmaster2_p & v37496fa;
assign v3752759 = hmaster1_p & v3a5e2a3 | !hmaster1_p & v3756981;
assign v37256d2 = hbusreq0 & v3739ac1 | !hbusreq0 & v8455ab;
assign b5394c = hgrant5_p & a80fe2 | !hgrant5_p & v37777d1;
assign v375eea5 = hbusreq8 & v3775932 | !hbusreq8 & v376ae94;
assign v37453d7 = hbusreq3_p & v37bfca2 | !hbusreq3_p & v8455ab;
assign v373a8b4 = hmaster2_p & v3a70d99 | !hmaster2_p & v3752fe6;
assign v377133f = hlock5 & v3a5ad17 | !hlock5 & v374cbe2;
assign v377dc65 = hmaster0_p & v37564a2 | !hmaster0_p & b2ea29;
assign v3a62cac = hbusreq5_p & v3a5ac8b | !hbusreq5_p & v8455ab;
assign v3a63930 = hmaster1_p & v375e21e | !hmaster1_p & v376cf96;
assign v3a5548b = hbusreq6_p & v3729531 | !hbusreq6_p & v3748797;
assign v3737bfe = hgrant5_p & v372e268 | !hgrant5_p & v3a6ac2c;
assign v3779d33 = hmaster2_p & v8455ab | !hmaster2_p & v3808eed;
assign v375930e = hmaster2_p & v3767561 | !hmaster2_p & v3a7084e;
assign v373ae4a = hmaster0_p & v37560b4 | !hmaster0_p & v373e2e5;
assign v3752248 = hmaster1_p & v3808ed2 | !hmaster1_p & v3a5958e;
assign v3a67bff = hbusreq2_p & v3a6f481 | !hbusreq2_p & v8455ab;
assign v3a5b51a = hgrant4_p & v373ae83 | !hgrant4_p & v374febd;
assign v3758a4b = hbusreq4_p & v3a6b860 | !hbusreq4_p & v3758a7b;
assign d3068c = hbusreq6 & v3730e7d | !hbusreq6 & v3a62a6d;
assign v3768036 = hbusreq7_p & v3777d51 | !hbusreq7_p & v3a66747;
assign v3739e25 = hbusreq0 & v372c86a | !hbusreq0 & v372984c;
assign v375dcd5 = hgrant4_p & v8455ab | !hgrant4_p & v37308a9;
assign v2093132 = hmaster0_p & v373b48c | !hmaster0_p & v3a6e8d9;
assign v3728cd0 = hgrant2_p & v8455ab | !hgrant2_p & v377df60;
assign v374a7b4 = hbusreq5_p & v3a561aa | !hbusreq5_p & !v8455ab;
assign v3758636 = hbusreq0 & v3a6fa86 | !hbusreq0 & v3750625;
assign v3759c96 = hmaster0_p & v375725f | !hmaster0_p & v8455ab;
assign v376e240 = hmaster1_p & v3a63777 | !hmaster1_p & v3a6f5e8;
assign v3735b64 = hmaster1_p & v9af7ec | !hmaster1_p & v374d59d;
assign v23fd7e1 = hmaster0_p & v374eb9e | !hmaster0_p & v3758c72;
assign v3a68c63 = hmaster1_p & v8455ab | !hmaster1_p & v3774200;
assign v39a4e7e = hbusreq7 & v374e3ab | !hbusreq7 & v3a6f703;
assign v377c0fe = hgrant2_p & v377b218 | !hgrant2_p & v374f12d;
assign v3a568ee = hmaster0_p & v376dcbe | !hmaster0_p & v375f145;
assign v37663a2 = hgrant1_p & v374b07b | !hgrant1_p & !v8455b6;
assign v372a61c = hbusreq0 & v3a6fc03 | !hbusreq0 & v8455ab;
assign v37632f8 = hbusreq6_p & v3759b2f | !hbusreq6_p & v3a6f43e;
assign v377c9bd = hbusreq6_p & v3a6efe1 | !hbusreq6_p & v8455ab;
assign v3a6fea0 = hmaster3_p & v37504f2 | !hmaster3_p & v372977b;
assign v374b992 = hbusreq0 & v374fe1a | !hbusreq0 & v8455ab;
assign v375c7b6 = stateA1_p & v37440c3 | !stateA1_p & v1e37481;
assign v3a715d0 = hlock8 & v3a6ae19 | !hlock8 & v373f6e7;
assign v374ff15 = hmaster0_p & v3749969 | !hmaster0_p & v3a63d22;
assign v3a711ee = hmaster0_p & v37447e9 | !hmaster0_p & v376aa3f;
assign v375a80c = hbusreq6 & v377bb66 | !hbusreq6 & v3a6d0a1;
assign v3a5e62b = hmaster2_p & v3a635ea | !hmaster2_p & v3a60a68;
assign cbc7dd = hbusreq5 & v3809542 | !hbusreq5 & v37333de;
assign v3a6f050 = hbusreq6 & v377e033 | !hbusreq6 & v372cc25;
assign v37240c0 = hgrant5_p & v8455ab | !hgrant5_p & v1e37b76;
assign a7afd8 = hlock2_p & v3747c3e | !hlock2_p & v8455ab;
assign v3a669bc = hmaster0_p & v3a57fb8 | !hmaster0_p & v8455e7;
assign v3754a4d = hbusreq4_p & v3a58907 | !hbusreq4_p & v3769945;
assign v3a5fb00 = hlock3 & v380733a | !hlock3 & v3768062;
assign v38075cd = hmaster0_p & v3769a1c | !hmaster0_p & v3a6f3a2;
assign v3793188 = hgrant4_p & v8455ab | !hgrant4_p & v8455c1;
assign v37678f8 = hmaster1_p & v3a639e7 | !hmaster1_p & !v375918d;
assign v373b71f = hmaster1_p & v373e553 | !hmaster1_p & v375993d;
assign v376c224 = hmaster2_p & v373c755 | !hmaster2_p & v8455ab;
assign v374f8b1 = hlock0_p & v376f665 | !hlock0_p & v8455ab;
assign v3a58640 = hmaster0_p & v3779060 | !hmaster0_p & v3a706f8;
assign v3731c79 = hbusreq6 & v376dcd0 | !hbusreq6 & !v3758e9e;
assign v3a70c90 = hgrant5_p & v3759fb9 | !hgrant5_p & v1e3737d;
assign v3777ce4 = hgrant6_p & v8455ab | !hgrant6_p & !v37395bc;
assign v3775aea = hbusreq3_p & v1e37ab9 | !hbusreq3_p & v376b734;
assign v3733cca = hgrant0_p & v8455ab | !hgrant0_p & v3a5ad13;
assign v3a5718e = hbusreq2_p & v3769628 | !hbusreq2_p & v8455ab;
assign v37625f2 = hmaster2_p & v377c7c0 | !hmaster2_p & v373aed4;
assign stateG10_8 = !v3a6521e;
assign v3763d10 = hbusreq4 & v3775303 | !hbusreq4 & v8455ab;
assign v3737d2f = hmaster2_p & v8455ab | !hmaster2_p & v37315da;
assign v374e18a = hbusreq8_p & v3a705cf | !hbusreq8_p & v372ee18;
assign v373fb30 = hgrant2_p & v3a6f6ba | !hgrant2_p & v374125a;
assign v3774901 = hbusreq5 & v3728d1d | !hbusreq5 & v8455ab;
assign v3a674e2 = hmaster1_p & v377aae4 | !hmaster1_p & v372a0a1;
assign v3a703fa = hmaster2_p & v8455ab | !hmaster2_p & v3a5b5ef;
assign v3752f21 = hlock0_p & v3748900 | !hlock0_p & v8455ab;
assign v377e04a = hmaster3_p & v37377f0 | !hmaster3_p & v3748004;
assign v375777d = hmaster0_p & v377d7bd | !hmaster0_p & v37445ff;
assign v3a705fc = hbusreq5 & v3a707a4 | !hbusreq5 & v374ab4b;
assign v376a77a = hmaster1_p & v3775651 | !hmaster1_p & v372ab0f;
assign v3755791 = hbusreq1 & v8455b0 | !hbusreq1 & v8455ab;
assign v37565ae = hgrant3_p & v3a710e9 | !hgrant3_p & v3a63197;
assign v3773434 = hlock0 & v373eaee | !hlock0 & v3740469;
assign v3739b38 = hmaster0_p & v3a6cccd | !hmaster0_p & !v373197c;
assign v37349ce = hlock6_p & v3724e8e | !hlock6_p & v3763a20;
assign v37433ff = hbusreq6 & v3a5e817 | !hbusreq6 & v37c0382;
assign v373abc5 = hmaster2_p & v380881d | !hmaster2_p & v3732359;
assign v373c183 = hbusreq7 & v3a6a413 | !hbusreq7 & v3a5e975;
assign v3730526 = hmaster0_p & v8455ab | !hmaster0_p & v376a0e3;
assign v3a6bd5a = hmaster3_p & v8455ab | !hmaster3_p & v3a6faab;
assign v3a664ba = hbusreq6_p & v8455ab | !hbusreq6_p & v3a5aee5;
assign v3a63866 = hmaster2_p & v3a5a01b | !hmaster2_p & v3747042;
assign v377dc0c = hbusreq0_p & v374f307 | !hbusreq0_p & v8455b0;
assign v3729c37 = hgrant0_p & v376e914 | !hgrant0_p & v374790d;
assign v3255a31 = hgrant0_p & v8455ab | !hgrant0_p & v3a66559;
assign v9c4c8d = hbusreq2 & v374732a | !hbusreq2 & v375b9c1;
assign v3a6f680 = hlock7_p & v3a71361 | !hlock7_p & v3a6d89d;
assign v3739b6a = hlock7 & v372b5c0 | !hlock7 & v375ff99;
assign v376fbcd = hbusreq2 & v376d9ad | !hbusreq2 & v8455e7;
assign v3a6cf75 = hmaster1_p & v376fbb5 | !hmaster1_p & v3724ced;
assign v374b24a = hmaster2_p & v372abac | !hmaster2_p & v3735272;
assign v376c9ee = locked_p & v376402f | !locked_p & v373d452;
assign v3766d0a = hmaster2_p & v3777da6 | !hmaster2_p & v37427e9;
assign v3750078 = hlock6_p & v3748ca3 | !hlock6_p & !v8455ab;
assign v373518a = hmaster1_p & v3a6fcb7 | !hmaster1_p & v8455ca;
assign v2619368 = decide_p & v3a6738f | !decide_p & v3a6fa4b;
assign v38094ca = hbusreq5_p & v375b6d4 | !hbusreq5_p & v3a65565;
assign v374bb9c = hgrant4_p & v8455ab | !hgrant4_p & v3a53e50;
assign v3a66db2 = hbusreq5 & v3a5b25b | !hbusreq5 & v8455e7;
assign v3a56f0b = hmaster0_p & v3a661fe | !hmaster0_p & v376db27;
assign v3743c89 = hbusreq4_p & v3a6fbe1 | !hbusreq4_p & v375a930;
assign v3a58dc1 = hlock6_p & v377de7b | !hlock6_p & v373f058;
assign v37356f0 = hlock3_p & v3763175 | !hlock3_p & !v8455ab;
assign v3737534 = hgrant2_p & v8455b9 | !hgrant2_p & v37607e8;
assign v3775da1 = hmaster3_p & v374e032 | !hmaster3_p & v3a6f8ce;
assign v373d661 = hbusreq5_p & v377de7f | !hbusreq5_p & v3766b6e;
assign v3746bdb = hburst0_p & v8455ab | !hburst0_p & v3769bf7;
assign v3a5e0e5 = hlock8 & v374e9d1 | !hlock8 & v376fddc;
assign v375d997 = hmaster1_p & v3a635ea | !hmaster1_p & v3a56e03;
assign v3a70e3a = hmastlock_p & v3760d59 | !hmastlock_p & v8455ab;
assign v3766c5c = hmaster2_p & v376e89b | !hmaster2_p & v3768685;
assign v375e854 = hbusreq0 & v3a54dfa | !hbusreq0 & v374ca4a;
assign v3808e9f = hmaster3_p & v3a714fe | !hmaster3_p & v376baad;
assign v374bd6a = hbusreq4_p & v3a6f365 | !hbusreq4_p & v3a70ee9;
assign v3a5bd05 = hlock4 & v38099a1 | !hlock4 & v3727b4a;
assign v3a70442 = hmaster1_p & v3769c6d | !hmaster1_p & v37735aa;
assign v3726e1f = hmaster2_p & v3763fdc | !hmaster2_p & v3732359;
assign v3a64d7c = hbusreq4_p & v3a61ce7 | !hbusreq4_p & v3a6c2a9;
assign v3725948 = hmaster1_p & v8455ab | !hmaster1_p & v374d9c0;
assign v3a69fde = hmaster0_p & v3754cb0 | !hmaster0_p & v3a6a9d7;
assign v3a6fa20 = hbusreq8 & v3a5faf0 | !hbusreq8 & v373c52e;
assign v3a70e4a = hlock7 & v3a6fe61 | !hlock7 & v3a702e3;
assign v3727b7f = hgrant5_p & v8455ab | !hgrant5_p & v3a70f68;
assign v3a6f796 = hmaster1_p & v372625f | !hmaster1_p & v3a5c7a2;
assign v37618ef = hbusreq4 & v3a6f7bf | !hbusreq4 & v8455e7;
assign v3765d05 = hlock8_p & v3734b5a | !hlock8_p & !v8455ab;
assign v3747569 = hbusreq2 & v373f622 | !hbusreq2 & v37731c3;
assign v3749139 = hbusreq5_p & v3757556 | !hbusreq5_p & v376dad4;
assign v9c1340 = hbusreq5_p & v37577cd | !hbusreq5_p & v3773eeb;
assign v3a6ed79 = hgrant2_p & v3748d67 | !hgrant2_p & v377002f;
assign v372f1a0 = hgrant2_p & v8455e7 | !hgrant2_p & !v374fd45;
assign v3729370 = hmaster1_p & v3a7166e | !hmaster1_p & v3744c88;
assign v376a040 = hbusreq6_p & v375a8cf | !hbusreq6_p & v3760658;
assign v3759aea = hbusreq8_p & v374fd0b | !hbusreq8_p & v377bc9f;
assign v375005c = hmaster1_p & v3a6220e | !hmaster1_p & v374ec57;
assign v3724475 = hbusreq6_p & v375937f | !hbusreq6_p & v3a53cfe;
assign v3762324 = hbusreq8_p & v372a1f6 | !hbusreq8_p & v374e620;
assign v3748c4c = jx3_p & v3751fde | !jx3_p & v376c3c2;
assign a15d51 = hbusreq5 & v3761472 | !hbusreq5 & v8455ab;
assign v3743ec6 = hmaster0_p & v3a64a9a | !hmaster0_p & v3a6fec4;
assign v3a6ec7a = hgrant3_p & v3a70626 | !hgrant3_p & v3a6ac26;
assign v3a71230 = hmaster0_p & v372b1dc | !hmaster0_p & v37471f0;
assign v3a6ca99 = hlock0_p & v380887a | !hlock0_p & v3736141;
assign v3a5bfc8 = hgrant4_p & v8455b5 | !hgrant4_p & v39a4e84;
assign v37558c7 = hmaster0_p & v3770957 | !hmaster0_p & v379318b;
assign v374e0f6 = hbusreq4_p & v8455ca | !hbusreq4_p & v3a640a0;
assign v377c6cf = hbusreq0 & v375b045 | !hbusreq0 & !v3765b09;
assign v376c863 = hlock4_p & v3772c12 | !hlock4_p & v375c845;
assign v3762cca = hgrant4_p & v39eb590 | !hgrant4_p & ce4c9b;
assign v2aca778 = hlock4 & v3738679 | !hlock4 & v3a6dfc9;
assign v3767aae = hgrant4_p & v8455ab | !hgrant4_p & v3737352;
assign v37545b7 = hmaster1_p & v8455e7 | !hmaster1_p & v374c120;
assign v3a6e0bf = jx1_p & v3a66039 | !jx1_p & v3a56aee;
assign v3767ff6 = hlock5 & v3a6eb5c | !hlock5 & v3735539;
assign v3a56f9f = hbusreq0 & v3a5bded | !hbusreq0 & v3a71138;
assign v373dc11 = hbusreq5 & v3a70209 | !hbusreq5 & !v8455ca;
assign v3a687ea = hbusreq2 & v3a5952d | !hbusreq2 & v3a707c4;
assign v3a6fc61 = hmaster1_p & v3a70276 | !hmaster1_p & v372895b;
assign v372fd4a = hmaster1_p & v3741869 | !hmaster1_p & v37611fb;
assign v3760629 = hbusreq2_p & v375c01d | !hbusreq2_p & v3a62122;
assign v1e37a26 = hgrant2_p & v3a653e4 | !hgrant2_p & !v209310e;
assign v373c8d0 = hlock4_p & v3a69515 | !hlock4_p & v3a6fe1a;
assign v3a5c8c9 = hbusreq5 & v3779680 | !hbusreq5 & v376cd02;
assign v372b686 = hmaster2_p & v3807aa1 | !hmaster2_p & !v3752536;
assign v374b25d = hlock3_p & v373ad95 | !hlock3_p & v8455ab;
assign v3767872 = hbusreq7_p & v3806ec9 | !hbusreq7_p & !v3378535;
assign v3731211 = hbusreq8_p & v376d542 | !hbusreq8_p & v3a647e7;
assign v37556fd = hbusreq6_p & v8455ab | !hbusreq6_p & v37665bf;
assign v3a71271 = hbusreq6_p & v374c33a | !hbusreq6_p & v374e26d;
assign v3a59d9d = hlock0_p & v3747302 | !hlock0_p & v37339f0;
assign v380989b = hbusreq0_p & v37682c6 | !hbusreq0_p & v377e928;
assign v3a67b58 = hgrant5_p & v3a671f2 | !hgrant5_p & v3722b10;
assign v3a2a770 = hgrant0_p & v8455ab | !hgrant0_p & v375356f;
assign v377b734 = hgrant6_p & v3a6ca4e | !hgrant6_p & v23fe10f;
assign v3a6f54d = hgrant4_p & v376935b | !hgrant4_p & !v3a70094;
assign v374abc9 = hgrant3_p & v376bb26 | !hgrant3_p & v3754e7b;
assign v37432d3 = hbusreq4_p & v37323a1 | !hbusreq4_p & v373d5dc;
assign v3732c0d = hmaster0_p & v374ea29 | !hmaster0_p & !v376df4c;
assign v37535c4 = hgrant4_p & v374a91e | !hgrant4_p & v3767adc;
assign v3a5f205 = hlock7 & v3759532 | !hlock7 & v3a63f7b;
assign v3a700af = hmaster0_p & v373b4e3 | !hmaster0_p & v3a6f3cd;
assign v3752b90 = hbusreq7_p & v3a710d3 | !hbusreq7_p & v3a5fa09;
assign v3740dc6 = hgrant4_p & v3769e94 | !hgrant4_p & v37503c9;
assign v3a6d156 = hgrant3_p & v374ef66 | !hgrant3_p & v360bcf2;
assign v3a57646 = hgrant7_p & v373a9db | !hgrant7_p & v3a70d76;
assign v3a571e5 = hbusreq7 & v37241a0 | !hbusreq7 & !v3744c88;
assign v3a70f44 = hmaster2_p & v3725bdc | !hmaster2_p & v8455ab;
assign v37574d3 = hgrant6_p & v37722e5 | !hgrant6_p & v372d9e0;
assign v3765d2b = hbusreq5_p & v8455ab | !hbusreq5_p & v376efcc;
assign v3a6fd95 = hbusreq2_p & v3772f4d | !hbusreq2_p & d0a27e;
assign v3754d47 = hbusreq5 & v3734502 | !hbusreq5 & v3a58c07;
assign v3764494 = hlock5 & v3734fba | !hlock5 & v3a63699;
assign v3a715e9 = hmaster1_p & v3a61149 | !hmaster1_p & v3a6efb9;
assign v373ce49 = hbusreq0 & v377f486 | !hbusreq0 & v8455ab;
assign v3763b94 = hmaster2_p & v3a5fabd | !hmaster2_p & v3a5f6d5;
assign v3748a0a = hbusreq7 & v3a69e59 | !hbusreq7 & v3734279;
assign v37609d6 = hbusreq4 & v325b5fd | !hbusreq4 & v3a68c23;
assign v3733132 = hbusreq6 & v374fe7b | !hbusreq6 & v375f9df;
assign v374fc6c = hgrant1_p & v374b07b | !hgrant1_p & !v8455ab;
assign v3a6bf00 = hmaster3_p & v375912e | !hmaster3_p & !v3a681f5;
assign v373f260 = hmaster1_p & v3a70225 | !hmaster1_p & v375a311;
assign v8a1014 = hmaster3_p & v3724579 | !hmaster3_p & v374e078;
assign v3a575e5 = hbusreq8 & v3a70878 | !hbusreq8 & !v8455c6;
assign v3757cd1 = hmaster0_p & v3776767 | !hmaster0_p & !v377e51b;
assign v3a714cc = hlock0 & v37763c2 | !hlock0 & v3a6f477;
assign v3774449 = hmaster0_p & v3731857 | !hmaster0_p & v374e8b4;
assign v3a6e8fa = hgrant3_p & v3779dae | !hgrant3_p & v374b383;
assign v373449c = hbusreq4 & v3a6b4ab | !hbusreq4 & v8455ab;
assign v373a452 = hlock6_p & v373fe5e | !hlock6_p & !v376430b;
assign v3776a2e = hmaster0_p & v375a10d | !hmaster0_p & v375e051;
assign v37386a9 = stateA1_p & v3a635ea | !stateA1_p & v8455ab;
assign v374c522 = hlock5 & v3751eb6 | !hlock5 & v377fc45;
assign v373c15d = hmaster0_p & v3a713f2 | !hmaster0_p & v37412f3;
assign v374809d = hbusreq2 & v372ca44 | !hbusreq2 & v3779cf9;
assign v374c1c3 = hbusreq1 & v373fe5e | !hbusreq1 & !v376653d;
assign v377d86e = hbusreq6_p & v39a537f | !hbusreq6_p & !v372d2ad;
assign v3754fcc = hmaster2_p & v3764dc0 | !hmaster2_p & v8455ab;
assign v3a6d5e2 = hmaster0_p & v3a70557 | !hmaster0_p & v3737a6e;
assign v3a6b4fb = hgrant1_p & v3a5b909 | !hgrant1_p & v376d327;
assign v373cdba = hmaster0_p & v3a5b289 | !hmaster0_p & v3a71288;
assign v37742d2 = hmaster1_p & v8455ab | !hmaster1_p & v3a56ffa;
assign v3807d59 = hlock4 & v37759b5 | !hlock4 & v3744b07;
assign v372c97c = hbusreq5 & v3a65b42 | !hbusreq5 & v375585a;
assign v375483e = hbusreq1 & v373d0b2 | !hbusreq1 & v3a7162d;
assign v3a53f45 = hgrant3_p & v372dcd4 | !hgrant3_p & v3a684ef;
assign v3767f36 = hmaster2_p & v39a537f | !hmaster2_p & v3728e09;
assign v3a57bd7 = hmaster2_p & v37583be | !hmaster2_p & !v3740df7;
assign v374df0b = hlock2_p & v37266b1 | !hlock2_p & v373e654;
assign v3761d7e = hbusreq8_p & v35b6dae | !hbusreq8_p & v3a6f737;
assign v376640a = hbusreq5_p & v3a71235 | !hbusreq5_p & v8455ab;
assign v372a79d = hmaster1_p & v3a71297 | !hmaster1_p & v3a706eb;
assign v372ac83 = hlock3_p & v3a6f052 | !hlock3_p & !v8455ab;
assign v3a59d65 = hlock0 & v3a67f97 | !hlock0 & v2ff8e9a;
assign v3766ef9 = hlock1 & v37722cc | !hlock1 & v373b288;
assign v372b34d = hbusreq8_p & v37250b5 | !hbusreq8_p & v3762720;
assign v3a5c066 = hmaster0_p & v3a62542 | !hmaster0_p & v3a595fe;
assign v3a61bac = hmaster2_p & v376b4e1 | !hmaster2_p & !v3759158;
assign v37731c3 = hgrant3_p & v8455ab | !hgrant3_p & v3a6c5fc;
assign v372ac49 = hlock3_p & v8455ab | !hlock3_p & v3a6ab5f;
assign v373833b = hmaster0_p & v375646d | !hmaster0_p & v3a6c892;
assign v372a3af = hbusreq0 & v3a6ff4f | !hbusreq0 & v373e814;
assign v3a6fc96 = hbusreq4_p & v372e562 | !hbusreq4_p & v8455ab;
assign v37449e7 = jx0_p & v376beca | !jx0_p & v8f4f53;
assign v3735580 = hgrant0_p & v8455ab | !hgrant0_p & !v3a70b0d;
assign v3752131 = hlock0 & v3a60a68 | !hlock0 & v3a6f908;
assign v3a6fe72 = hmaster2_p & v3733d6e | !hmaster2_p & v3a6a213;
assign v3a6f3d9 = hbusreq6_p & v3a6fb66 | !hbusreq6_p & v3a6fe9f;
assign v3a6fd67 = hmaster2_p & v373b589 | !hmaster2_p & v3776441;
assign v35b70ee = hmaster2_p & v375d616 | !hmaster2_p & v8455ab;
assign v3a714d8 = hmaster2_p & v39ea76e | !hmaster2_p & !v3735e39;
assign v3a55d7c = hbusreq6 & v8455b0 | !hbusreq6 & v3755791;
assign v3a710eb = hlock4 & v3a63da7 | !hlock4 & v376f23f;
assign v372b3b0 = hmaster2_p & v376501e | !hmaster2_p & !v3a6f081;
assign v3751ecb = hlock2_p & v3773250 | !hlock2_p & !v8455ab;
assign v3a6eab8 = hbusreq8_p & v3768a7b | !hbusreq8_p & v3a6ff56;
assign v3732b35 = hbusreq4_p & v3759032 | !hbusreq4_p & !v39a537f;
assign v3a71239 = hgrant5_p & v3a70746 | !hgrant5_p & v3a6f96b;
assign v3a69c73 = hready_p & v373578f | !hready_p & v3765ad4;
assign v3a6f72f = hmaster1_p & v3a56c60 | !hmaster1_p & v374bac7;
assign v3a70bba = hmaster2_p & v3764dc0 | !hmaster2_p & v372a1d6;
assign v373291c = hgrant3_p & v8455ab | !hgrant3_p & v33790da;
assign v3a71078 = hgrant2_p & v8455ab | !hgrant2_p & v3a7014e;
assign v3724b8c = hbusreq5 & v3a711cb | !hbusreq5 & v375d9df;
assign v3a7043e = hlock4_p & v8455ab | !hlock4_p & v8455e7;
assign ba7f1c = hmaster2_p & v8455ab | !hmaster2_p & v37433ef;
assign v3a67eec = hlock3 & v37408a3 | !hlock3 & v37416b5;
assign v373be21 = hbusreq6 & v3733383 | !hbusreq6 & v8455ab;
assign v3775b4d = hbusreq6_p & v3734e58 | !hbusreq6_p & v3758f64;
assign v373d943 = hlock5 & v3769cc4 | !hlock5 & v3809dfb;
assign v374e29a = hgrant2_p & v8455b9 | !hgrant2_p & v3a708e2;
assign v3a70112 = hlock4_p & v3a62072 | !hlock4_p & v3a615a2;
assign v3773343 = jx2_p & v3739246 | !jx2_p & v37fca9f;
assign v3775c51 = hmaster0_p & v3a66110 | !hmaster0_p & !v3760e51;
assign v32559c3 = hbusreq4 & v373aaa8 | !hbusreq4 & v8455ab;
assign v3a6ae04 = hlock5_p & v3764677 | !hlock5_p & v3a701f2;
assign v3a5ead2 = stateA1_p & v3743bc5 | !stateA1_p & v376a35c;
assign v3a71284 = hbusreq3 & v37665bf | !hbusreq3 & v8455ab;
assign v3759181 = hgrant3_p & v372493b | !hgrant3_p & v3758c46;
assign v3723211 = hgrant4_p & v37615c5 | !hgrant4_p & v3724d99;
assign v377beee = hbusreq8 & v37682dd | !hbusreq8 & v3a6f60c;
assign v3a56b4e = hlock0 & v373785d | !hlock0 & v3a6fab9;
assign v372814c = jx0_p & v373361a | !jx0_p & v3754e33;
assign v376d86d = hlock0 & v3753dd4 | !hlock0 & v3a63884;
assign v3a6ff0e = hmaster1_p & v3a635ea | !hmaster1_p & v3746473;
assign v3732dac = hbusreq0 & v373d78b | !hbusreq0 & v8455ab;
assign v3763c97 = hmaster0_p & v3a6f114 | !hmaster0_p & !v8455c3;
assign v3754a42 = hlock4 & v375a261 | !hlock4 & v372ea4b;
assign v373b1cb = hlock4_p & v373325b | !hlock4_p & v3a6fac6;
assign v3738eb6 = hbusreq1 & v39a5265 | !hbusreq1 & !v35b9d52;
assign v37613b3 = hmaster1_p & v3a70d99 | !hmaster1_p & v3762e16;
assign v3729555 = hmaster1_p & v377234d | !hmaster1_p & v3a7093d;
assign v3777b5b = hbusreq5 & v3763846 | !hbusreq5 & v357742d;
assign v3a56d01 = hbusreq6_p & v3a6a213 | !hbusreq6_p & !v373e8ad;
assign v373293c = hbusreq7_p & v372f03c | !hbusreq7_p & v3a6c555;
assign v374b05b = hbusreq0 & v3a7054a | !hbusreq0 & v37488fe;
assign v3771c3a = hgrant0_p & v3744693 | !hgrant0_p & !v3776a6e;
assign v3a6ed49 = hbusreq8 & v8455b0 | !hbusreq8 & v8455ab;
assign v3a62973 = hbusreq3 & v373a391 | !hbusreq3 & v8455ab;
assign v373e8df = hmaster2_p & v37469c4 | !hmaster2_p & dc5fea;
assign v372b5a3 = hgrant6_p & v3742ac7 | !hgrant6_p & v8455ab;
assign v377ef0b = hgrant5_p & v373e2aa | !hgrant5_p & v3725c60;
assign v37573a3 = hlock0 & v3765e79 | !hlock0 & v3a6f17b;
assign v3a5cc9d = hbusreq2_p & v377773f | !hbusreq2_p & v3757fcc;
assign v3a6f7f0 = hgrant0_p & v37384fa | !hgrant0_p & v374ab5b;
assign v39a4f17 = hbusreq4 & v3771c59 | !hbusreq4 & d1bf3b;
assign v37229f0 = hgrant4_p & v8455ab | !hgrant4_p & v3a7133b;
assign v3735fc0 = hlock6 & v373f953 | !hlock6 & v37248e4;
assign v3a62abc = hbusreq3_p & v3a67dc7 | !hbusreq3_p & !v8455ab;
assign v376296b = hmaster1_p & v3a5c57a | !hmaster1_p & v3a6988c;
assign v3756261 = hlock0_p & v377eaf2 | !hlock0_p & v377d33e;
assign v375c8db = hmaster1_p & v3a635ea | !hmaster1_p & v3758661;
assign v3737101 = hbusreq2_p & v374bb02 | !hbusreq2_p & v8455ab;
assign da7312 = hmaster1_p & v3757966 | !hmaster1_p & v3a6c610;
assign v37787ce = hmaster0_p & v375e217 | !hmaster0_p & !v3776f07;
assign v37373af = hgrant6_p & v3a637dc | !hgrant6_p & v3a70a92;
assign v3a61392 = hlock3_p & v3774a13 | !hlock3_p & !v1e379fe;
assign v3727981 = hmaster0_p & v372cd04 | !hmaster0_p & v23fe28c;
assign v3a6573d = hbusreq6_p & v8455bb | !hbusreq6_p & v3773ff0;
assign v376a006 = hgrant2_p & v8455ba | !hgrant2_p & v373e9a9;
assign v3a70b4b = hmaster0_p & v376025f | !hmaster0_p & v3756219;
assign v3a68e46 = hmaster0_p & v3759fd0 | !hmaster0_p & v376bad7;
assign v3a711f7 = hbusreq8_p & v3765583 | !hbusreq8_p & v3a58fe9;
assign v3a5cd4c = hbusreq4_p & v375808f | !hbusreq4_p & v3a5b855;
assign v377fb55 = hbusreq8 & v3724d8b | !hbusreq8 & v377a89f;
assign v3a6b691 = hlock3_p & v3776a5c | !hlock3_p & v372faf1;
assign v37389ba = hbusreq5 & v3a60924 | !hbusreq5 & v375b0ad;
assign v376740f = hmaster0_p & v8455ab | !hmaster0_p & !v37556ae;
assign v3a70b13 = hmaster1_p & v37666f6 | !hmaster1_p & v375aff8;
assign v380730d = hgrant2_p & v8455ab | !hgrant2_p & v3771e60;
assign v372cf62 = stateG2_p & v8455ab | !stateG2_p & v3a6446a;
assign v3a5bbec = hlock0 & v376e90a | !hlock0 & v3a69b93;
assign v3735f02 = hgrant2_p & v8455ab | !hgrant2_p & v375dbe0;
assign v3777e0a = hgrant6_p & v3a6f402 | !hgrant6_p & v3a60a40;
assign v3a6f187 = hmaster2_p & v20930c6 | !hmaster2_p & v3a6f1e7;
assign v3a711fd = hmaster1_p & v374a0b1 | !hmaster1_p & v374472d;
assign v3760509 = hgrant4_p & v2ff87b0 | !hgrant4_p & v3a70a70;
assign v3a64421 = hgrant4_p & v3a69de7 | !hgrant4_p & v3a635ea;
assign v3a5c4d5 = hgrant0_p & v37773a9 | !hgrant0_p & v3a5ae2f;
assign v37767e6 = hbusreq6_p & v3775179 | !hbusreq6_p & v8455ab;
assign v3768095 = hgrant1_p & v3766448 | !hgrant1_p & !v8455ab;
assign v3738cd4 = jx1_p & v3809dcb | !jx1_p & v3731edf;
assign v3a6528b = hbusreq3_p & v2092f90 | !hbusreq3_p & v8455b0;
assign v375035f = hbusreq7_p & v3809e77 | !hbusreq7_p & v375ea88;
assign v3a5e7be = hgrant5_p & v3728333 | !hgrant5_p & v3768c53;
assign v3742f0a = hgrant4_p & v372de1e | !hgrant4_p & v3807113;
assign v3a63eaf = hbusreq6_p & v8455e7 | !hbusreq6_p & v374f307;
assign v374674d = hmaster2_p & v3a54eae | !hmaster2_p & v373df13;
assign v3a70f06 = hmaster1_p & v3a5bf4c | !hmaster1_p & v3a29850;
assign v37641ad = hgrant4_p & v8455ab | !hgrant4_p & v372abf1;
assign v374d645 = hmaster0_p & v377bb3a | !hmaster0_p & v37545a0;
assign v374510e = hbusreq6_p & v375cfd7 | !hbusreq6_p & v377652b;
assign v3a70de3 = hmaster1_p & v374a36b | !hmaster1_p & v377e915;
assign v3a5ae6d = hbusreq1_p & v3a6fc6c | !hbusreq1_p & v3a70b73;
assign v3a708d6 = hbusreq5 & cd743d | !hbusreq5 & v3774bad;
assign v3a6fcbe = hbusreq5_p & v372e544 | !hbusreq5_p & v374aa1b;
assign v3733690 = hbusreq4 & v377c214 | !hbusreq4 & v3809ec3;
assign v3a7103a = hbusreq0 & v380a0c2 | !hbusreq0 & !v1e37cd6;
assign v3a70134 = hbusreq5 & v2092a9a | !hbusreq5 & v3a6f122;
assign v372d48d = hgrant2_p & v3a6cfe0 | !hgrant2_p & v3729e05;
assign v3746f89 = hbusreq8 & v37260fc | !hbusreq8 & v3a63f55;
assign v376ce6f = hbusreq5 & v372ca24 | !hbusreq5 & v374ed5a;
assign v3377b0f = hmaster0_p & v3a5e999 | !hmaster0_p & v3767b70;
assign v373ec8f = hmaster2_p & v377ef09 | !hmaster2_p & v374b8fa;
assign v3764a94 = hlock6_p & v3a5dd7f | !hlock6_p & v373006f;
assign v3a70753 = hbusreq4 & v3a6582b | !hbusreq4 & v3752cf6;
assign v375c2e2 = hmaster3_p & v377de72 | !hmaster3_p & v3a6764b;
assign v3a5b2fd = hgrant3_p & v3762502 | !hgrant3_p & v37427d3;
assign v3752397 = hbusreq2 & v373fda2 | !hbusreq2 & v3723efc;
assign v3774d04 = hgrant1_p & v373b288 | !hgrant1_p & v3a63621;
assign v3a709ed = hmaster2_p & v37718fb | !hmaster2_p & v3a63659;
assign v374ebe8 = hbusreq0 & v3764e52 | !hbusreq0 & v37742f1;
assign v37511c6 = hmaster0_p & v3a6d614 | !hmaster0_p & v3748179;
assign v374fcd2 = hbusreq6 & v3a70200 | !hbusreq6 & !v372870d;
assign v376eb68 = hmaster0_p & v3a7002c | !hmaster0_p & v375d263;
assign v377e453 = hmaster2_p & v377f526 | !hmaster2_p & v3732359;
assign v3a5f9d2 = hbusreq0 & v3a70629 | !hbusreq0 & v8455ab;
assign v376a06d = hmaster1_p & d7669b | !hmaster1_p & v3759cb9;
assign v3a6eb19 = hlock5_p & v3a5cff8 | !hlock5_p & v3a712e4;
assign v3a706ce = hlock4_p & v3a5614c | !hlock4_p & v3746fce;
assign v377a893 = jx0_p & v3772b42 | !jx0_p & v373d746;
assign v3757f6d = hmaster1_p & v3a6542a | !hmaster1_p & v9e6ddd;
assign v3771182 = hbusreq7_p & v3731d66 | !hbusreq7_p & v8455ab;
assign v376f237 = hmaster2_p & v373366b | !hmaster2_p & v37314fa;
assign v3a6ed4c = hbusreq4 & v376f0a0 | !hbusreq4 & v3731230;
assign v3a29842 = hgrant3_p & ae7027 | !hgrant3_p & v3740ee1;
assign v376c0d8 = hlock5_p & v3769a34 | !hlock5_p & v3a701f2;
assign v1e378da = hbusreq4 & v8455b0 | !hbusreq4 & v8455ab;
assign v376a21c = hlock0_p & v8455ab | !hlock0_p & v375401a;
assign v3a6f70f = hbusreq5 & v372954d | !hbusreq5 & v8455ab;
assign v3a67a06 = hlock1_p & v377dc87 | !hlock1_p & v3722dba;
assign v3a713e1 = locked_p & v3a6f71d | !locked_p & v8455ab;
assign v1e37cd7 = hmaster0_p & v375babe | !hmaster0_p & v3a6ee64;
assign v3a594ab = hmaster2_p & v3a620ef | !hmaster2_p & v373da95;
assign v37514e4 = hbusreq5 & v376d640 | !hbusreq5 & v37763b2;
assign v375eee3 = hgrant4_p & v8455ab | !hgrant4_p & v3747ad5;
assign v3a59391 = hgrant2_p & v8455ab | !hgrant2_p & b755d3;
assign v37667f7 = hbusreq4 & v3723fce | !hbusreq4 & v3a55641;
assign v3a7052a = hgrant3_p & v377dd3b | !hgrant3_p & v376d3f7;
assign v3745734 = hmaster0_p & v372a53e | !hmaster0_p & v3730d6c;
assign v3a704e0 = hbusreq8_p & v3767b77 | !hbusreq8_p & a13040;
assign v3754164 = hmaster2_p & v377c6ce | !hmaster2_p & v3a6a374;
assign v3a6e9a4 = stateG10_1_p & v8455e7 | !stateG10_1_p & !v3a60205;
assign v3726229 = hbusreq2_p & v375bdd4 | !hbusreq2_p & v8455e1;
assign v373d81e = jx1_p & v37528b8 | !jx1_p & v3a700d2;
assign v372f046 = hmaster2_p & v39a4ca8 | !hmaster2_p & !v3a55cd6;
assign v3a709c1 = hbusreq3_p & v3777d41 | !hbusreq3_p & v8455b0;
assign v3a70198 = hmaster2_p & v372935c | !hmaster2_p & !v3728e09;
assign v373a982 = hmaster1_p & v3775651 | !hmaster1_p & !v3a7124d;
assign v38087ba = hmaster2_p & v37535c4 | !hmaster2_p & v3775e2e;
assign v376983e = hbusreq4_p & v3754b79 | !hbusreq4_p & v3806798;
assign v374729b = hlock0_p & v3807bf8 | !hlock0_p & v3a5e357;
assign v23fdf76 = hbusreq0 & v374b3cf | !hbusreq0 & v8455ab;
assign v3a7137a = hgrant4_p & v376d285 | !hgrant4_p & !v37545a5;
assign v3a70f55 = hbusreq8_p & v3742c64 | !hbusreq8_p & v37c028d;
assign v3a55904 = hmaster0_p & v3772b14 | !hmaster0_p & v37243fe;
assign v377db88 = hgrant4_p & v37300a5 | !hgrant4_p & b6ae10;
assign v37246d9 = hlock5_p & v3768da7 | !hlock5_p & v3748a16;
assign v374d972 = hlock8_p & v8455ab | !hlock8_p & v3755e66;
assign v3a703c5 = hgrant4_p & v8455ab | !hgrant4_p & v3727420;
assign v374b3cf = hlock0_p & v3765e46 | !hlock0_p & !v8455ab;
assign v373e6d2 = hgrant4_p & v375cdee | !hgrant4_p & v374776e;
assign v3a6f668 = hbusreq3 & v8455ab | !hbusreq3 & v373a391;
assign v375c674 = hgrant6_p & v3744cfe | !hgrant6_p & v3a5b286;
assign v375feba = hgrant6_p & v3739a53 | !hgrant6_p & v2619ae8;
assign v37397c3 = hbusreq1_p & v37286bb | !hbusreq1_p & v374fef8;
assign v3770e35 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3746145;
assign v3a6f693 = hmaster2_p & v37356cc | !hmaster2_p & !v8455ab;
assign v3a6f15d = hbusreq7_p & v376fa86 | !hbusreq7_p & v3a296d3;
assign v3a6ccfe = hbusreq8 & v373b667 | !hbusreq8 & v374a98e;
assign v3754107 = hmaster1_p & v8455ab | !hmaster1_p & v3a714a6;
assign v3747d58 = hbusreq4 & v3808f45 | !hbusreq4 & v8455ab;
assign d24921 = hlock5 & v3731b28 | !hlock5 & v373d5b7;
assign v376c63d = hbusreq2 & v37637d6 | !hbusreq2 & v8455ab;
assign v37386f5 = hbusreq2_p & v3745158 | !hbusreq2_p & v8455ab;
assign v3a5ba97 = hlock2_p & v3769758 | !hlock2_p & v3a5e020;
assign v3753f59 = hmaster3_p & v374a601 | !hmaster3_p & v37408a1;
assign v3762434 = hbusreq1 & v3770f7a | !hbusreq1 & v3a635ea;
assign v23fdc13 = hgrant6_p & v8455ca | !hgrant6_p & v1e38239;
assign v377a606 = hbusreq4 & v376b88d | !hbusreq4 & v3a70d99;
assign v3733b84 = hbusreq8 & v23fe152 | !hbusreq8 & v376fff8;
assign v373c8db = hgrant5_p & v3a64bcf | !hgrant5_p & v3a64da2;
assign v3a7087c = hmaster1_p & v3730a34 | !hmaster1_p & v3734caf;
assign v3779931 = hbusreq5_p & v375b6c3 | !hbusreq5_p & !v376bc8c;
assign v37394b7 = hmaster0_p & v376d550 | !hmaster0_p & !v37654c4;
assign v37582e6 = hbusreq8_p & v37737d2 | !hbusreq8_p & b6057e;
assign v3a5eafa = hlock3 & v3726777 | !hlock3 & v3807c0c;
assign v3a2a107 = hmaster0_p & v8455ab | !hmaster0_p & v3a6fde0;
assign v3a5e9a3 = hlock1_p & v3a7103c | !hlock1_p & !v8455ab;
assign v3a6fe71 = hbusreq6 & v3a6dc08 | !hbusreq6 & v373f058;
assign v3a70ac9 = hbusreq4_p & v377d1cd | !hbusreq4_p & v8455b0;
assign v3739621 = hgrant5_p & v3a70938 | !hgrant5_p & v375e50f;
assign v3741dab = hgrant2_p & v3a70b17 | !hgrant2_p & v37313b6;
assign v374ae67 = jx0_p & v3a5d6f9 | !jx0_p & v3a6267a;
assign v377416d = hbusreq4 & v3a58924 | !hbusreq4 & v8455ab;
assign v3a70ba8 = hbusreq4_p & v3a6ac60 | !hbusreq4_p & v375cbdf;
assign v372cdd7 = hmaster2_p & v3a6bc65 | !hmaster2_p & !v3a71453;
assign v3a6f632 = hmaster0_p & v3763f95 | !hmaster0_p & v3a6fa7a;
assign v3762a76 = hmaster0_p & v3a7026c | !hmaster0_p & v37584e6;
assign c7885c = hmaster0_p & v374502e | !hmaster0_p & v3745c45;
assign v3a7086d = hmaster0_p & v3a6f60d | !hmaster0_p & v3735485;
assign v3809ebc = hbusreq3_p & v3764979 | !hbusreq3_p & v8455ab;
assign v917087 = hbusreq6 & v3a5a7fd | !hbusreq6 & v373d4ff;
assign v3767904 = hbusreq3_p & v3752ec0 | !hbusreq3_p & v374f318;
assign v3761d0c = hbusreq4_p & v377d377 | !hbusreq4_p & v376afc5;
assign v3775723 = hmaster1_p & v3a53e30 | !hmaster1_p & v377dd0d;
assign v3770b6c = hmaster0_p & v3738b8a | !hmaster0_p & v3a6f31f;
assign v3733383 = hready & v2619b26 | !hready & v8455e7;
assign v3a5795e = hlock2_p & v37399b4 | !hlock2_p & v3a6f147;
assign v3762de1 = hbusreq1 & v374cab9 | !hbusreq1 & v37674c1;
assign v3775932 = hmaster1_p & v377bb3a | !hmaster1_p & v3a6c016;
assign v3770161 = hbusreq4_p & v3a71213 | !hbusreq4_p & v3a71024;
assign v3a70e2a = hgrant2_p & v376e914 | !hgrant2_p & !v3a6f842;
assign v37711c5 = hgrant6_p & v3733e9e | !hgrant6_p & v3723ee7;
assign v3728d72 = hlock6 & v372a6c2 | !hlock6 & v3a5c700;
assign v374c256 = hbusreq8_p & v376ae9f | !hbusreq8_p & v3a68170;
assign v3a5fcc2 = hbusreq7_p & v3a5e5ec | !hbusreq7_p & v376e9e1;
assign v3a704c9 = hgrant2_p & v3730e2e | !hgrant2_p & v3809a76;
assign v3778993 = hbusreq3_p & v3a70641 | !hbusreq3_p & v8455e7;
assign v374d749 = hbusreq6 & v37338d8 | !hbusreq6 & v37443ab;
assign v3771758 = hbusreq4_p & v3a6f520 | !hbusreq4_p & !v8455ab;
assign v3a6f0f4 = hmaster2_p & v8455ab | !hmaster2_p & !v8455c1;
assign v3a6ec0f = hmaster1_p & v39eb550 | !hmaster1_p & v3a5f602;
assign v3746d75 = hgrant5_p & v3744f6f | !hgrant5_p & v372f0ee;
assign v3a67e67 = hbusreq4_p & v3a6fbe1 | !hbusreq4_p & v3751238;
assign v3a6126c = hgrant4_p & v374d011 | !hgrant4_p & v8455ab;
assign v3744131 = hbusreq6_p & v37560ff | !hbusreq6_p & v3a5beb5;
assign v325c960 = hbusreq6_p & v37416ea | !hbusreq6_p & !v8455ab;
assign v39a5293 = hgrant2_p & v372310a | !hgrant2_p & v3766a98;
assign v3752a6c = hgrant5_p & v3727d4c | !hgrant5_p & v3a5b51d;
assign v3a67eb2 = hmaster1_p & v377dacb | !hmaster1_p & v3a70ae8;
assign v3a70375 = hmaster2_p & v3a6df32 | !hmaster2_p & v3728d9c;
assign v375f55e = hlock5 & v3a64a14 | !hlock5 & v38072a2;
assign v3a62aef = hgrant4_p & v8455ab | !hgrant4_p & v38063a0;
assign v37385de = hlock2_p & v3a637dd | !hlock2_p & !v8455ab;
assign v3739b5c = hlock5_p & v377854f | !hlock5_p & v8455bb;
assign v3a6f832 = hgrant4_p & v8455ab | !hgrant4_p & v3809d45;
assign v37563ef = hbusreq7 & v3732b1d | !hbusreq7 & v377386a;
assign v372d925 = hmaster0_p & v373014d | !hmaster0_p & v3773ce0;
assign v3a683d2 = hgrant3_p & v3a6b873 | !hgrant3_p & v3759590;
assign v374c5b2 = hbusreq3_p & v372ac49 | !hbusreq3_p & v8455ab;
assign v377051a = hgrant1_p & v3747c3e | !hgrant1_p & v8455ab;
assign v3a64b90 = hlock4 & v3a5d6c6 | !hlock4 & d2e9f6;
assign v377da29 = hmaster1_p & v373e8cb | !hmaster1_p & v3779ac0;
assign v3a6f590 = hlock7_p & v374802b | !hlock7_p & v3a674c9;
assign v3a70dae = hlock4_p & v3768ac7 | !hlock4_p & v8455ab;
assign v3a709de = hmaster3_p & v3772c4d | !hmaster3_p & v2ff8e61;
assign v3a68232 = hlock5_p & v3a5d929 | !hlock5_p & v3a6b306;
assign v3a56789 = hbusreq5 & v3a70f62 | !hbusreq5 & v376fbb5;
assign v37519e5 = hmaster1_p & v3a6a2ab | !hmaster1_p & !v374a9eb;
assign v3a7055c = hbusreq5_p & v374f0ac | !hbusreq5_p & v372f4fe;
assign v3a5cb6f = hbusreq0 & v3723e5d | !hbusreq0 & v92a03a;
assign v377f67b = hgrant4_p & v3a6b873 | !hgrant4_p & v37259e6;
assign v3a70d42 = hgrant2_p & v3a6c580 | !hgrant2_p & v376ef36;
assign v3754445 = hbusreq8 & v376b4d4 | !hbusreq8 & v3a60276;
assign v373a196 = hlock4 & v3725bab | !hlock4 & v3a6a493;
assign v377380a = hbusreq5_p & v3a70cb2 | !hbusreq5_p & v3a6f3ac;
assign v3a6c4e4 = hbusreq6_p & v3a70214 | !hbusreq6_p & v8455ab;
assign v372ee4b = hmaster2_p & v377234d | !hmaster2_p & v3760a58;
assign v3a70a45 = hgrant0_p & v375dbeb | !hgrant0_p & v3753964;
assign v37681f3 = hbusreq4_p & v3a5f9d2 | !hbusreq4_p & v374ebc5;
assign v377586d = hmaster1_p & v3767b62 | !hmaster1_p & v3a5591a;
assign v375a33d = hmaster1_p & v377e018 | !hmaster1_p & a52d64;
assign v3a703a1 = hgrant0_p & v8b397d | !hgrant0_p & !v8455ab;
assign v3a59c73 = hmaster1_p & v3a706c2 | !hmaster1_p & v373e055;
assign v373c526 = hbusreq4_p & v380881d | !hbusreq4_p & v3a63bb7;
assign v3a7043d = hmaster1_p & v377b48b | !hmaster1_p & !v375b5eb;
assign v3808d0f = hmaster1_p & v8455ca | !hmaster1_p & v3756d53;
assign v3a65c29 = hlock1 & v38072fd | !hlock1 & v37748e5;
assign v3727db9 = hgrant2_p & v3743b9e | !hgrant2_p & v374b4a4;
assign v3a71275 = hbusreq4_p & v377edba | !hbusreq4_p & !v3a5c5f4;
assign v373794a = hmaster0_p & v3724703 | !hmaster0_p & v376f504;
assign v3a70f37 = hgrant3_p & v8455ab | !hgrant3_p & v3a6859a;
assign v3a6f2be = hmaster1_p & v3a6b8a0 | !hmaster1_p & v3a551d7;
assign v38073b0 = hbusreq6_p & v37796c6 | !hbusreq6_p & v372989d;
assign v3758a92 = hmaster2_p & v3a663b9 | !hmaster2_p & v377d58d;
assign v3726791 = hbusreq3 & v3a67e64 | !hbusreq3 & !v3746fce;
assign v3a627a7 = hgrant6_p & v3772404 | !hgrant6_p & v376646a;
assign v3a71377 = hgrant4_p & v3731320 | !hgrant4_p & v3757f01;
assign v3a7150f = hmaster1_p & v3a71110 | !hmaster1_p & v3a6b68e;
assign v372c335 = hmaster1_p & c03a6a | !hmaster1_p & !v3a67e97;
assign v3774aa2 = hbusreq6 & v3738d0b | !hbusreq6 & v375da10;
assign v37366fc = hbusreq6 & v3809788 | !hbusreq6 & v3779cf9;
assign v3772bb1 = hmaster0_p & v375469c | !hmaster0_p & v8455ab;
assign v3a704fe = hmaster1_p & v3a6e975 | !hmaster1_p & v374bb64;
assign v3737f8d = hmaster2_p & v3743c40 | !hmaster2_p & !v8455ab;
assign v3766f51 = hmaster1_p & v3a635ea | !hmaster1_p & v374f2d2;
assign b9d061 = hlock7 & v37563ef | !hlock7 & v3732b1d;
assign v3775e35 = hbusreq5_p & v377de7f | !hbusreq5_p & v375367c;
assign v3759b46 = hbusreq5_p & v373a9c4 | !hbusreq5_p & v3a71249;
assign v3a7144d = hmaster2_p & v3760513 | !hmaster2_p & v376d9c6;
assign v3a6f330 = hmaster1_p & v8455bd | !hmaster1_p & v3767e47;
assign v3a6eb21 = hbusreq5 & v3769edd | !hbusreq5 & v3774bad;
assign v3a6165b = hbusreq7 & v3769e10 | !hbusreq7 & a0a219;
assign v3770d70 = stateG10_1_p & v3751fa8 | !stateG10_1_p & v3726277;
assign v3a69118 = hgrant5_p & v3731003 | !hgrant5_p & v3a5aef6;
assign v3a7031d = hbusreq3 & v374362e | !hbusreq3 & !v3a568f7;
assign v3a6c243 = hgrant3_p & v3a5872a | !hgrant3_p & v375e6b3;
assign v372e367 = hbusreq4 & v3a7043e | !hbusreq4 & v8455ab;
assign v3774b25 = hready & v377ac6f | !hready & v8455ab;
assign v374974e = hmaster2_p & v3a71018 | !hmaster2_p & v3a6ebb3;
assign v3a6a19b = hmaster2_p & v8455ab | !hmaster2_p & v38072fd;
assign v3a6f550 = hmaster2_p & v373cf9c | !hmaster2_p & v3a6f4c7;
assign v375377b = hbusreq8_p & v3765763 | !hbusreq8_p & v37407ef;
assign v377e2e3 = hmaster0_p & v3724394 | !hmaster0_p & v3a6e118;
assign v3a70fad = hbusreq8 & v3762452 | !hbusreq8 & v3779075;
assign v37471c2 = hlock7_p & v3a6fc6b | !hlock7_p & v3a5e998;
assign v3750eb9 = hmaster2_p & v35b7092 | !hmaster2_p & v37697a3;
assign v3a62541 = hmaster1_p & v3a7006c | !hmaster1_p & v373a7a1;
assign v3728b28 = hmastlock_p & v865472 | !hmastlock_p & !v8455ab;
assign v374636c = hmaster2_p & v8455ab | !hmaster2_p & v37674c1;
assign v374a8bb = hmaster0_p & v3731c7b | !hmaster0_p & v3a5c3d3;
assign v3a5cd20 = hgrant0_p & v8455b3 | !hgrant0_p & v3776a6e;
assign v3a712d2 = hlock7_p & a36719 | !hlock7_p & v37586ed;
assign v373d53f = hbusreq6_p & v3a6f804 | !hbusreq6_p & v374569b;
assign v3767c3e = jx1_p & v375cce7 | !jx1_p & v8455ab;
assign v37316c9 = hgrant4_p & v8455ab | !hgrant4_p & v3a70db6;
assign v3a6a9cd = jx1_p & v374c048 | !jx1_p & v3a70392;
assign v3740a38 = hlock6 & v3a5f75a | !hlock6 & v3a67ec4;
assign v3a68b0a = hmaster2_p & v3a637dc | !hmaster2_p & v373ad95;
assign v374bf55 = hgrant6_p & v3726bff | !hgrant6_p & v3769e8c;
assign v376e1fb = hlock5 & v372a309 | !hlock5 & v37345de;
assign v3a62e91 = hmaster2_p & v3a6fd72 | !hmaster2_p & v3758fa8;
assign v2092f0a = start_p & v8455ab | !start_p & v375ab35;
assign v3744a60 = hbusreq6_p & v375af5d | !hbusreq6_p & v8455ab;
assign v374c837 = hmaster0_p & v3757993 | !hmaster0_p & v3a56002;
assign v3a5aac9 = hlock5_p & v3a5d2c5 | !hlock5_p & v3751022;
assign v37629e2 = hgrant3_p & v3a6f627 | !hgrant3_p & v377e9c4;
assign v375cdf4 = hbusreq4 & v3736c8d | !hbusreq4 & v3a70d64;
assign v3772464 = hlock5_p & v376e115 | !hlock5_p & v8455e7;
assign v377a808 = hbusreq5 & v3761c5e | !hbusreq5 & v377709a;
assign v377d839 = hmaster2_p & v3a635ea | !hmaster2_p & v373b288;
assign v374072b = hmaster1_p & v3757dee | !hmaster1_p & v3759ac1;
assign v3754e70 = hbusreq6_p & v3a712d6 | !hbusreq6_p & v3743b79;
assign v3763f6f = hlock4_p & v374b3bf | !hlock4_p & v37406d2;
assign v38079ff = hgrant0_p & v1e3791d | !hgrant0_p & v3a66559;
assign v373bf45 = hgrant6_p & v373313b | !hgrant6_p & v3a5bd48;
assign v37439a0 = hlock5_p & v3731866 | !hlock5_p & !v3a704af;
assign v37406e8 = hgrant4_p & v3a5aa3a | !hgrant4_p & v3a6f309;
assign v375a0af = hbusreq8 & v375d7d2 | !hbusreq8 & v3733483;
assign v3a71591 = hbusreq8 & v374bf93 | !hbusreq8 & v8455ab;
assign v3a6c98c = hbusreq6 & v376495e | !hbusreq6 & v8455ab;
assign v3a6fc57 = hmaster1_p & v3a6f942 | !hmaster1_p & v376c611;
assign v3a56243 = hmaster2_p & v37625a8 | !hmaster2_p & !v372493b;
assign v3742bc3 = hmaster0_p & v3a700b2 | !hmaster0_p & v3a6fcd2;
assign v374cab5 = hbusreq6_p & v376a96b | !hbusreq6_p & v3a5f485;
assign v377d6ba = hgrant6_p & v39eb4cb | !hgrant6_p & v3a6afe8;
assign v3761e59 = hmaster1_p & v376a3f7 | !hmaster1_p & v377de07;
assign v37490d7 = hbusreq8_p & v3763c1f | !hbusreq8_p & v37351ff;
assign v3741dee = hbusreq4_p & v372c17e | !hbusreq4_p & v8455ab;
assign v374c2e2 = hmaster1_p & v23fe361 | !hmaster1_p & v3a70381;
assign v3740bf7 = hmaster1_p & v374c5fc | !hmaster1_p & v23fda78;
assign v374bcb4 = hbusreq6 & v3747994 | !hbusreq6 & v8455ab;
assign v3743c35 = hmaster1_p & v209312a | !hmaster1_p & d2ccfa;
assign v37787ec = locked_p & v3a71137 | !locked_p & v8455ab;
assign v37377c8 = hmaster2_p & v3a61397 | !hmaster2_p & !v8455ab;
assign v375bc38 = hbusreq6_p & v3772e33 | !hbusreq6_p & v37413d5;
assign v374f16d = hbusreq7_p & v3775cc9 | !hbusreq7_p & v376e66e;
assign v373d91f = hbusreq6 & v3a70180 | !hbusreq6 & v3734db5;
assign v375eb1b = hmaster1_p & v37386c6 | !hmaster1_p & v3a6ec20;
assign v374044c = hgrant6_p & v3a669c2 | !hgrant6_p & v3757aa1;
assign v3778372 = hmaster0_p & v3762858 | !hmaster0_p & v3764683;
assign v3a702cc = hbusreq4_p & v3a68d49 | !hbusreq4_p & v360be60;
assign c7d127 = hbusreq4 & v37538ff | !hbusreq4 & v3763104;
assign v3a5cf3d = hbusreq2_p & v3772443 | !hbusreq2_p & v8455ab;
assign v3739be4 = hgrant4_p & v8455ab | !hgrant4_p & !v3a701d8;
assign v374fb2f = hgrant5_p & v3771162 | !hgrant5_p & v375b234;
assign v37526cd = hbusreq6 & v3a6dc08 | !hbusreq6 & v375d616;
assign v37482da = hmaster1_p & v3a5fabd | !hmaster1_p & v3a6f4e3;
assign v3a71189 = hmaster2_p & v3729421 | !hmaster2_p & !v37564e4;
assign c9c058 = hbusreq5 & v376a6f1 | !hbusreq5 & v38064e5;
assign v374c000 = hbusreq5_p & v3a6fd64 | !hbusreq5_p & !v8455ab;
assign v3a70891 = hgrant4_p & v3a65762 | !hgrant4_p & v3a6d1b9;
assign v3756bc2 = hbusreq3 & v8455b0 | !hbusreq3 & v3755791;
assign v37548f5 = hmaster0_p & v3739cfb | !hmaster0_p & v372efee;
assign v3744da3 = hmaster0_p & v3759031 | !hmaster0_p & v3742b9d;
assign v3733ea2 = hburst1 & v35b9d52 | !hburst1 & v3a5ef0c;
assign v3733103 = hbusreq6 & v3809259 | !hbusreq6 & v37372c9;
assign v374e985 = hmaster2_p & v3a5c562 | !hmaster2_p & v37711c3;
assign v8716e3 = hbusreq6 & v3a6e222 | !hbusreq6 & v372e83f;
assign v374294c = hmaster1_p & v3a708d4 | !hmaster1_p & v3746da7;
assign v3765a43 = hgrant0_p & v372b931 | !hgrant0_p & v37747fc;
assign v3751c1c = hmaster2_p & v3746d2a | !hmaster2_p & v3757c7f;
assign v3736afd = hbusreq0 & v376ba89 | !hbusreq0 & v37648cd;
assign v3a6f4dd = hmaster1_p & v376665a | !hmaster1_p & v3770fdb;
assign v374e6b1 = hmaster2_p & v3769950 | !hmaster2_p & v3778b60;
assign v3778ab7 = hbusreq5_p & v3a713e2 | !hbusreq5_p & v377ea3c;
assign v372dffe = hbusreq4_p & v3a5b0dd | !hbusreq4_p & v3736f61;
assign v3734d20 = hmaster1_p & v3a6edb5 | !hmaster1_p & v372c23b;
assign v37763bd = hbusreq5_p & v375e177 | !hbusreq5_p & v8455b0;
assign v376ecde = hbusreq5 & v3747b02 | !hbusreq5 & v8455ab;
assign v377209d = hbusreq7 & v3a7032b | !hbusreq7 & v3755a27;
assign d5959b = hbusreq0 & v3751291 | !hbusreq0 & v3a70b06;
assign v3a648c3 = hbusreq0_p & v3747302 | !hbusreq0_p & v3768062;
assign v3a623f2 = hgrant6_p & v3a653e4 | !hgrant6_p & !v3730f77;
assign v377d4dc = hgrant2_p & v3a70dc4 | !hgrant2_p & v3a62d54;
assign v37501a3 = hmaster3_p & v372bad7 | !hmaster3_p & v377180a;
assign v3a7112c = hbusreq4_p & v3a6efe8 | !hbusreq4_p & v373b381;
assign v375ff0d = hbusreq4 & v3737e04 | !hbusreq4 & v38072fd;
assign v375d00d = hmaster0_p & v372379e | !hmaster0_p & v3729173;
assign v37252c2 = hbusreq6_p & v373cb54 | !hbusreq6_p & v375975b;
assign v3753edb = hlock0_p & v3806db7 | !hlock0_p & v37536df;
assign v37414d1 = hbusreq6 & v37482f8 | !hbusreq6 & !v377b7ad;
assign v3a5a2c6 = hlock5_p & v374478f | !hlock5_p & v37647e3;
assign v3a66273 = hbusreq4 & v376ecc8 | !hbusreq4 & !v3a640a0;
assign v37771a8 = hgrant4_p & v8455ab | !hgrant4_p & v3763e76;
assign v377af0a = hbusreq2 & v374362e | !hbusreq2 & v3a676d6;
assign v373683d = hbusreq4 & v3a55bd0 | !hbusreq4 & v2092abe;
assign v377a13b = hbusreq5 & v372b10b | !hbusreq5 & v357742d;
assign v372b316 = hlock5_p & v3a63e68 | !hlock5_p & v374801c;
assign v3a6f119 = hbusreq2_p & v375dbe0 | !hbusreq2_p & v3761f39;
assign v3755a27 = hmaster1_p & v3746406 | !hmaster1_p & v3a70d99;
assign v3a70eee = hmaster3_p & v376f641 | !hmaster3_p & v3726bb7;
assign v3774058 = hmaster1_p & v3732b15 | !hmaster1_p & v372bd2b;
assign v3738726 = hmaster0_p & v3733dea | !hmaster0_p & v8455e7;
assign v376d3e2 = hmaster1_p & v39eb4e4 | !hmaster1_p & v3776923;
assign v3a708e2 = hbusreq2_p & v3a5fc3c | !hbusreq2_p & v373125c;
assign v3a67e25 = hbusreq5 & v3a6ae04 | !hbusreq5 & v8455ab;
assign v37450ff = hgrant2_p & v38072f4 | !hgrant2_p & !v373ed95;
assign v3a708b9 = hlock2 & v375b736 | !hlock2 & v372da4f;
assign v3a708fd = hlock0_p & v3a635ea | !hlock0_p & v3a70b5f;
assign v37541b4 = hmaster0_p & v39eaff9 | !hmaster0_p & v377b6b2;
assign v374f677 = hgrant6_p & v3a6eb2d | !hgrant6_p & v3748fba;
assign v3a5a2cd = hlock5_p & v3a6fa1c | !hlock5_p & !v8455ab;
assign v3a59a05 = hmaster2_p & v3771ddb | !hmaster2_p & v3a70809;
assign v37242f1 = hbusreq8_p & v3808943 | !hbusreq8_p & v3769a62;
assign v3a6f99b = hgrant4_p & a7adce | !hgrant4_p & v376575c;
assign v373fff3 = hgrant0_p & v8455ab | !hgrant0_p & !v37345e9;
assign v3a6eb63 = hgrant1_p & d44200 | !hgrant1_p & !v8455ab;
assign v89e294 = hmaster3_p & v3741edb | !hmaster3_p & v37347d9;
assign v3a69d8f = hmaster0_p & v8455e7 | !hmaster0_p & v3731741;
assign v375a338 = hgrant5_p & v3778b2a | !hgrant5_p & v374bd1f;
assign v3a70217 = hbusreq5_p & v3a540a1 | !hbusreq5_p & !v37474d6;
assign v3747462 = jx0_p & v8455bd | !jx0_p & !v8455b9;
assign v3723676 = hlock2_p & v3756206 | !hlock2_p & v3a63bdb;
assign v377d393 = hbusreq3 & v3767f33 | !hbusreq3 & v8455e7;
assign v374f609 = hgrant0_p & v8455ab | !hgrant0_p & !v8455b6;
assign v3a67f8e = hbusreq6 & v3a6ff0c | !hbusreq6 & v8455ab;
assign v3a680bd = hmaster2_p & ca01e4 | !hmaster2_p & v37522d3;
assign v3a6c8e4 = hbusreq5_p & v3730526 | !hbusreq5_p & v3736058;
assign v376c30a = hbusreq4 & v3a703bb | !hbusreq4 & v373f3b5;
assign v372ed79 = hmaster0_p & v3722e59 | !hmaster0_p & v3758cec;
assign v3a5bca4 = hbusreq2_p & v3a6f20d | !hbusreq2_p & v3748d67;
assign v3a71032 = hlock8 & v3756595 | !hlock8 & v376a946;
assign v374a7cd = hgrant0_p & v8455b5 | !hgrant0_p & v2678bee;
assign v374edb8 = hbusreq8 & v377faff | !hbusreq8 & v3a7118e;
assign v3a6190f = hbusreq6_p & v377476b | !hbusreq6_p & v3766e4a;
assign v3a70105 = hmaster0_p & v3a6df14 | !hmaster0_p & v3758ff0;
assign v374930c = hmaster0_p & v3a6f608 | !hmaster0_p & v3a71202;
assign v3a6eec3 = hbusreq5_p & v3a7075b | !hbusreq5_p & v377b416;
assign v3776386 = hbusreq6_p & v20d166d | !hbusreq6_p & v3725395;
assign v37571c8 = hmaster2_p & v3a6fc7f | !hmaster2_p & v374b526;
assign v3a65711 = hmaster0_p & v373318b | !hmaster0_p & v376e056;
assign v37772db = hbusreq6_p & v3a58ba8 | !hbusreq6_p & v3a63621;
assign v374063d = hbusreq0_p & v3a708ec | !hbusreq0_p & v8455ab;
assign v374d6b5 = jx1_p & v374b237 | !jx1_p & !v3774629;
assign v375043b = hbusreq7_p & v3a6680b | !hbusreq7_p & v3722d85;
assign v372bcf2 = hmaster1_p & v3735236 | !hmaster1_p & v3a64879;
assign v37647e3 = hmaster0_p & v3a65909 | !hmaster0_p & v3a69606;
assign v375d009 = hgrant3_p & v374212e | !hgrant3_p & cf6441;
assign v373a6f8 = hbusreq5 & v3a67965 | !hbusreq5 & v3a6ae2f;
assign v3a70743 = hmaster2_p & v3a55456 | !hmaster2_p & v8455e7;
assign v3754740 = jx1_p & v374ed80 | !jx1_p & v37602b1;
assign v3a5f4b1 = hlock4 & v376435f | !hlock4 & v373628e;
assign v376b870 = hmaster2_p & v8455b0 | !hmaster2_p & v35b7808;
assign v3751369 = hmaster2_p & v8455e7 | !hmaster2_p & v375571d;
assign v3a5d522 = hmaster0_p & v374e8b5 | !hmaster0_p & v3761719;
assign v376301d = hmaster2_p & v3741384 | !hmaster2_p & v373f2b6;
assign v3761950 = hbusreq5_p & v3742649 | !hbusreq5_p & v3747ef9;
assign v372d237 = hbusreq5_p & v3768b80 | !hbusreq5_p & v2aca81d;
assign v3a6f543 = hmaster3_p & v3758663 | !hmaster3_p & v3750e8a;
assign v3760bfa = hbusreq5 & v374bd23 | !hbusreq5 & v373de86;
assign v3a6d4f3 = hmaster0_p & v3a635ea | !hmaster0_p & v37670db;
assign v375c3f6 = hmaster2_p & v8455ab | !hmaster2_p & !v375efa4;
assign v3746cdc = hgrant2_p & v8455ab | !hgrant2_p & v3773b2f;
assign v375000b = hgrant2_p & v37435a0 | !hgrant2_p & v8455ab;
assign v3746cc5 = hgrant4_p & v8455ab | !hgrant4_p & v3a6eee4;
assign v376e5b6 = hmaster0_p & v8455ab | !hmaster0_p & v209325d;
assign v373c97a = hbusreq2 & v3777417 | !hbusreq2 & v8455ab;
assign v3a63f7b = hmaster1_p & v3a635ea | !hmaster1_p & v37484ac;
assign v3a7125f = hbusreq6 & v376289b | !hbusreq6 & v8455ab;
assign v37368df = hgrant1_p & v377eb2d | !hgrant1_p & v8455ab;
assign v3a6b51b = hlock4 & v3a6f105 | !hlock4 & v3a64056;
assign v377e9c1 = jx0_p & v377866b | !jx0_p & v3779486;
assign v37529d9 = hbusreq4 & v3a6fdd2 | !hbusreq4 & v8455ab;
assign v376e160 = hlock8 & v3a70e90 | !hlock8 & v3a64539;
assign v3a6eb7a = hmaster0_p & v372e443 | !hmaster0_p & v3750b8c;
assign v3a6ea2b = hbusreq5 & v37247b5 | !hbusreq5 & v3762642;
assign v373419f = hmaster1_p & v3a573af | !hmaster1_p & v3747514;
assign v3a63bde = hmaster0_p & v3a65c2a | !hmaster0_p & v3769f01;
assign v3a70725 = hbusreq4 & v3a6fe0e | !hbusreq4 & v3a63a66;
assign v325c90f = hmaster0_p & v372c41f | !hmaster0_p & v372f07d;
assign v3774369 = hmaster1_p & v377adf5 | !hmaster1_p & v3a70eac;
assign v3a5aef8 = hmaster1_p & v377234d | !hmaster1_p & v3a6fe7e;
assign v3a6b931 = hmaster0_p & v3a6de93 | !hmaster0_p & v3757765;
assign v3a6eb2f = hbusreq4_p & v3a7084e | !hbusreq4_p & v3a5c6f9;
assign v37674f2 = jx0_p & v376daac | !jx0_p & v373d0eb;
assign v3a6ffdc = hmaster0_p & v8455ab | !hmaster0_p & v3743486;
assign v3a64854 = hmaster2_p & v35772a6 | !hmaster2_p & v37580b3;
assign v3a55347 = hgrant0_p & v375297d | !hgrant0_p & ad2d05;
assign v3a69631 = hbusreq7 & v3725325 | !hbusreq7 & v8455c3;
assign v3a6fb49 = hbusreq8_p & v375faac | !hbusreq8_p & v3a6f5e6;
assign v3748acd = hmaster2_p & v3a5af28 | !hmaster2_p & v3771d4f;
assign v3770027 = hgrant4_p & v8455e7 | !hgrant4_p & !v3a7119f;
assign v3a6fa33 = hbusreq5_p & v375cc8b | !hbusreq5_p & !v8455ab;
assign v372bdef = hbusreq1_p & v377b690 | !hbusreq1_p & !v8455ab;
assign v3778e3f = hlock5 & v376b72d | !hlock5 & v373d66c;
assign v374afa4 = hbusreq4 & v3a63abb | !hbusreq4 & v8455ab;
assign v3a6fa2a = hmaster1_p & v376b036 | !hmaster1_p & c46b05;
assign v1e37dd9 = hbusreq2 & v37269f4 | !hbusreq2 & v3773ee6;
assign v3a6f5b8 = hlock7_p & d5e2c2 | !hlock7_p & !v3a6fd5d;
assign v3769d3e = hgrant3_p & v8455be | !hgrant3_p & v372b7e5;
assign v374834b = hmaster2_p & v35b774b | !hmaster2_p & v375e657;
assign v3a6f490 = hmaster2_p & v8455ab | !hmaster2_p & v373cc0f;
assign v37499ac = hmaster1_p & v3a635ea | !hmaster1_p & v375f9f1;
assign v209300b = hbusreq5_p & v37446d8 | !hbusreq5_p & v3a714c5;
assign v3749fd0 = hmaster0_p & v3a6c001 | !hmaster0_p & !v3a6fcab;
assign bdc0a1 = hgrant5_p & v377e319 | !hgrant5_p & ab4f60;
assign v3a6f425 = hbusreq3 & v372f85e | !hbusreq3 & v3807107;
assign v377974f = hmaster1_p & v3a71194 | !hmaster1_p & v3a70516;
assign v3a680e1 = hmaster2_p & v375e721 | !hmaster2_p & v376e35e;
assign a17325 = hlock2 & v372f6ce | !hlock2 & v3a587bc;
assign v376bbc5 = hmaster0_p & v373eba7 | !hmaster0_p & v3a5bd69;
assign v3777d41 = hlock3_p & v37502d9 | !hlock3_p & v377222b;
assign v3a705cf = hmaster1_p & v376e5b6 | !hmaster1_p & v8455ab;
assign v374f75e = hmaster2_p & v374f178 | !hmaster2_p & v3a5be6d;
assign v3a715ca = hbusreq4 & v3a5c6f9 | !hbusreq4 & v3727084;
assign v3a67904 = hgrant3_p & v376495e | !hgrant3_p & v3729ae4;
assign v3a6ad0b = hmaster2_p & v3a6f443 | !hmaster2_p & v3733e9e;
assign v3a712a5 = hmaster1_p & v3a7010b | !hmaster1_p & v3a67e97;
assign v3a70c83 = jx1_p & v3a70280 | !jx1_p & v3748443;
assign v3a70c8e = hmaster0_p & v3a675df | !hmaster0_p & v8455e7;
assign v3a64252 = hlock0_p & v2aca977 | !hlock0_p & v8455ab;
assign v372475e = hgrant2_p & v37699a0 | !hgrant2_p & v39a4db0;
assign v374bfa6 = hmaster2_p & v3a635ea | !hmaster2_p & v373a7a5;
assign v37593cb = hmaster2_p & v8455cb | !hmaster2_p & v37229c2;
assign v373187a = hbusreq4_p & v3726d1f | !hbusreq4_p & v3a7108f;
assign v3729724 = hbusreq1_p & v1e37d3f | !hbusreq1_p & v374648b;
assign v377b981 = hmaster2_p & v8455ab | !hmaster2_p & v3766487;
assign v3a5844c = hmaster0_p & v3748ded | !hmaster0_p & v3a68426;
assign v3761f13 = hmaster3_p & v3a68183 | !hmaster3_p & v3a70f6d;
assign v3a59c12 = hmaster0_p & v8455ab | !hmaster0_p & !v37525b0;
assign v3a5d1c9 = hlock8_p & v8c5d6a | !hlock8_p & v375a2ac;
assign a61f6b = hgrant2_p & v3a5c823 | !hgrant2_p & v37637d6;
assign v3758532 = hbusreq5 & v373c3e1 | !hbusreq5 & !v8455ab;
assign v37579f1 = hbusreq5_p & v3a57721 | !hbusreq5_p & v375a367;
assign v3a5e975 = hgrant5_p & b58331 | !hgrant5_p & v377bdd1;
assign v3767efa = hmaster0_p & v3a71678 | !hmaster0_p & v372a92a;
assign v3a663ef = hmaster0_p & v3a6f2c9 | !hmaster0_p & v3a6980b;
assign v3726739 = hlock0 & v3748797 | !hlock0 & v37233a7;
assign v3768918 = hbusreq5 & v3a63512 | !hbusreq5 & v3745bbe;
assign v3751141 = hbusreq7_p & v3a5666f | !hbusreq7_p & v3a60859;
assign v3a6f69f = hbusreq4 & v3731eff | !hbusreq4 & v3a635ea;
assign v3a614a0 = hlock5 & v3a705ae | !hlock5 & v3a70fc4;
assign v37319cd = hbusreq4_p & v3a5f69c | !hbusreq4_p & v37378e5;
assign v3a6f0be = hbusreq6 & v37314b5 | !hbusreq6 & v3a6c5ee;
assign v3749293 = jx2_p & v3737c52 | !jx2_p & v3a70473;
assign v37586e4 = hmaster0_p & v8455b0 | !hmaster0_p & v3a6d003;
assign v374df64 = hbusreq4 & v3a6e468 | !hbusreq4 & v8455ab;
assign v372ad5d = hmaster2_p & v8455ab | !hmaster2_p & v3a6c44c;
assign v3a61a75 = hlock5_p & v37694f9 | !hlock5_p & v37573f5;
assign v377928c = hbusreq2_p & v374da4a | !hbusreq2_p & v8455ab;
assign v3a6bbc6 = hmaster2_p & v8455ab | !hmaster2_p & v3a70cda;
assign v3a707bb = hbusreq0_p & v376d793 | !hbusreq0_p & v373b288;
assign v37497dd = hbusreq4_p & v3768c3c | !hbusreq4_p & !v374c7f4;
assign v3751e80 = hgrant6_p & v8455ab | !hgrant6_p & v37308b0;
assign v3769524 = hgrant8_p & v3a6f7b7 | !hgrant8_p & v377b4fa;
assign v3742ac7 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v374a637;
assign v3728455 = hmaster1_p & v3a635ea | !hmaster1_p & v374333e;
assign v3a61a2d = hmaster0_p & v373e474 | !hmaster0_p & v372e33d;
assign v3a6859a = hbusreq3_p & v1e37d2a | !hbusreq3_p & v8455ab;
assign v3744ca2 = hbusreq3_p & v3a6fc29 | !hbusreq3_p & !v37761b6;
assign v375cc11 = hbusreq0 & v3a6f962 | !hbusreq0 & v37578bd;
assign v3740490 = hmaster0_p & v37605e6 | !hmaster0_p & v3753097;
assign v37303f0 = hbusreq7_p & v3a6167d | !hbusreq7_p & v377d23d;
assign v3a70582 = hmaster0_p & v3a635ea | !hmaster0_p & v37729e0;
assign v3771204 = hbusreq5 & v3748ff3 | !hbusreq5 & v8455ab;
assign v373d07a = hmaster2_p & v3a57f59 | !hmaster2_p & v3a6d684;
assign v3732a75 = hbusreq5_p & v3735077 | !hbusreq5_p & v8455ab;
assign v374233c = hbusreq6_p & v3779cb7 | !hbusreq6_p & v376187f;
assign d95e20 = hmaster2_p & v3a63de8 | !hmaster2_p & !v8455ab;
assign v37559b4 = hmaster2_p & v3a6dfb2 | !hmaster2_p & v375e60f;
assign v209325d = hmaster2_p & v8455ab | !hmaster2_p & !v3755cb2;
assign v373070b = hgrant7_p & v373977e | !hgrant7_p & v3a6c42b;
assign v372f0e0 = hlock8 & v372cb36 | !hlock8 & v372b646;
assign v3741fe8 = hmaster1_p & v377e156 | !hmaster1_p & v377db66;
assign v3736cd2 = hbusreq8_p & v376ce17 | !hbusreq8_p & v3a70e73;
assign v3755820 = hbusreq6_p & v377caa3 | !hbusreq6_p & v37280b0;
assign v3a621be = hgrant2_p & v8455ab | !hgrant2_p & v3751905;
assign v37324bb = hmaster0_p & v374650c | !hmaster0_p & v373d40a;
assign v3a6cc5f = hbusreq7 & v3a5e388 | !hbusreq7 & !v3a5a954;
assign v3a715f2 = hbusreq4_p & v3a6a442 | !hbusreq4_p & v37235bd;
assign v3a6fb9b = hmaster0_p & v377adf5 | !hmaster0_p & v373739c;
assign v373330a = hbusreq4 & v3768685 | !hbusreq4 & v3a70d99;
assign v37556ec = hlock6 & v3a5f38a | !hlock6 & v3a70180;
assign v375d51e = hgrant3_p & v8455ab | !hgrant3_p & v37277c3;
assign v3760314 = hmaster0_p & v3a5b8a2 | !hmaster0_p & v3a6fe27;
assign v373f954 = hlock4_p & v3a6b5bc | !hlock4_p & v37395f5;
assign v375fed9 = hgrant6_p & v376a040 | !hgrant6_p & !v373e7c0;
assign v3767642 = locked_p & v8455ab | !locked_p & v3a70e49;
assign v9e2dd1 = hgrant6_p & v3771fb3 | !hgrant6_p & v3a71261;
assign v3a6f453 = hburst1_p & v3730383 | !hburst1_p & !v8455ab;
assign v3a6c0c5 = hgrant4_p & v3a7133d | !hgrant4_p & v3a59d07;
assign v3a6efe1 = hbusreq6 & v3749f78 | !hbusreq6 & v8455ab;
assign v373513a = hmastlock_p & v8455ff | !hmastlock_p & v8455ab;
assign v3a70c74 = hlock0_p & v374f35a | !hlock0_p & v374e16a;
assign v3a6f1a4 = hbusreq3 & v3a6fa39 | !hbusreq3 & v8455ab;
assign v3a6beb6 = hgrant2_p & v8455ab | !hgrant2_p & v3a708a8;
assign v3761da5 = hmaster1_p & v3a58017 | !hmaster1_p & v3762145;
assign v3a70967 = hmaster2_p & v8455ab | !hmaster2_p & v373f2b6;
assign v3a5d62d = hlock8 & v3726072 | !hlock8 & v37402a4;
assign v3750087 = hmaster1_p & v372673d | !hmaster1_p & v375e9a9;
assign v3a56abc = hmaster3_p & v3765322 | !hmaster3_p & !v3729caa;
assign v3a65605 = hgrant2_p & v3a5c823 | !hgrant2_p & v375cade;
assign v372408b = hbusreq0 & v3a63002 | !hbusreq0 & v3743332;
assign v3a6fec5 = hbusreq7 & v2ff8f77 | !hbusreq7 & v8455ab;
assign v380777c = hbusreq5_p & v3774e8d | !hbusreq5_p & v8455ab;
assign v372da2f = hmaster0_p & v372bd06 | !hmaster0_p & v373fdfb;
assign aebd68 = hbusreq2 & v373e296 | !hbusreq2 & v3a635ea;
assign v3a6fefa = hgrant3_p & v37496fa | !hgrant3_p & v372842d;
assign v37796c6 = hlock0_p & v3a6fa39 | !hlock0_p & !v8455ab;
assign v3a700fa = hmaster0_p & v3764276 | !hmaster0_p & v3727a4d;
assign v3779264 = hbusreq0_p & v3a635ea | !hbusreq0_p & v377857d;
assign v3a70624 = hbusreq2_p & v3a6613e | !hbusreq2_p & v37563fe;
assign v376b72d = hbusreq5 & v373d66c | !hbusreq5 & v374c5fc;
assign v3a703bb = hgrant6_p & v3a6fe44 | !hgrant6_p & v3741dac;
assign v376587d = hgrant5_p & v3765e47 | !hgrant5_p & v3731499;
assign v3752147 = hbusreq4_p & v3a635ea | !hbusreq4_p & v37592ca;
assign v3a7089f = hgrant2_p & v3a5a3c7 | !hgrant2_p & v37720ca;
assign v3738263 = hmaster1_p & v3726c8c | !hmaster1_p & v3728d9c;
assign v3750f1e = hbusreq8 & v3a5dab7 | !hbusreq8 & v8455ab;
assign v3806ff5 = hmaster2_p & v3747302 | !hmaster2_p & v376bb26;
assign v3730a93 = hbusreq4 & v380879c | !hbusreq4 & v38078ed;
assign v375d9b1 = hbusreq4_p & v373325f | !hbusreq4_p & v3a70025;
assign v37668cb = hbusreq6_p & v3723404 | !hbusreq6_p & v375d6ba;
assign v3737711 = hgrant5_p & v375f5c1 | !hgrant5_p & v3a70107;
assign v3a6f6eb = hmaster1_p & v3a58022 | !hmaster1_p & v37324bb;
assign v3a70195 = hmaster1_p & v8455ab | !hmaster1_p & v3749899;
assign v372c23b = hbusreq5_p & v3a6ff33 | !hbusreq5_p & v372620f;
assign v3a635ea = hmastlock_p & v3731d80 | !hmastlock_p & v8455ab;
assign v375018e = hbusreq3_p & v8455ab | !hbusreq3_p & v3a5cd20;
assign v373ac50 = hbusreq4 & v3733b37 | !hbusreq4 & v8455e7;
assign v3a69a50 = hbusreq5_p & v373cae5 | !hbusreq5_p & !v3a6fde5;
assign v3a5ce2d = hlock1 & v37764b1 | !hlock1 & v37386a9;
assign v3745131 = hgrant6_p & v37304b3 | !hgrant6_p & v377c723;
assign v377594d = hgrant6_p & v3a70ee7 | !hgrant6_p & v3a6ef23;
assign v372e708 = hbusreq4_p & v3748797 | !hbusreq4_p & v375c75c;
assign v3a5de1e = hmaster3_p & v3760337 | !hmaster3_p & !v3a681f5;
assign v3a70471 = hmaster3_p & v376f01b | !hmaster3_p & v377a893;
assign v374f5e0 = hgrant4_p & v375cdee | !hgrant4_p & v3a70d94;
assign v374df14 = hbusreq2_p & v3a6f8f5 | !hbusreq2_p & v3731487;
assign ab808e = hmaster0_p & v3740fe2 | !hmaster0_p & !v3a62dfa;
assign v372fd5d = hgrant4_p & v8455ab | !hgrant4_p & v3a585fd;
assign v3a6adb2 = hbusreq6_p & v376711c | !hbusreq6_p & v375d6ba;
assign v37604b3 = hbusreq6_p & v8455ab | !hbusreq6_p & v377803f;
assign v3a70476 = hmaster2_p & v8455ab | !hmaster2_p & v37438b9;
assign v3a5d156 = hgrant6_p & v8455ab | !hgrant6_p & v3a6fa06;
assign v875999 = hlock0_p & v372eaaf | !hlock0_p & !v8455ab;
assign v37583be = hburst1 & v1e38224 | !hburst1 & v373ed70;
assign v37694de = hbusreq3 & v3740171 | !hbusreq3 & v8455ab;
assign v3a6c97d = hbusreq2_p & v3a62826 | !hbusreq2_p & v35b774b;
assign v3a70952 = hgrant6_p & v375f2ec | !hgrant6_p & v3a591b4;
assign v374b5b6 = hgrant4_p & v9ed516 | !hgrant4_p & v3a70088;
assign v37680b5 = hbusreq8 & v3a56570 | !hbusreq8 & v3734279;
assign v376e0fa = hbusreq6_p & v3a6f9df | !hbusreq6_p & !v3a704c2;
assign v377e71d = hbusreq6 & v3772e46 | !hbusreq6 & v8455ab;
assign v377f785 = hbusreq0 & v8455ab | !hbusreq0 & !v377c31d;
assign v3743b11 = hbusreq7_p & v376ad33 | !hbusreq7_p & v376cd0a;
assign v377940a = hmaster2_p & v8455ab | !hmaster2_p & v3a60280;
assign v3a6f7ae = hmaster1_p & v3777bfc | !hmaster1_p & v3a70f10;
assign v3a70638 = hmaster1_p & v3a63777 | !hmaster1_p & v3772e8e;
assign v3758661 = hmaster0_p & v3a635ea | !hmaster0_p & v3a6d499;
assign v3748282 = hbusreq8_p & v3a712b5 | !hbusreq8_p & v96ab98;
assign v373fda2 = hbusreq3_p & v37583be | !hbusreq3_p & v3a6469c;
assign v3736184 = hmaster2_p & v3748cce | !hmaster2_p & v375f98a;
assign v3a5c30f = hgrant4_p & v8455ab | !hgrant4_p & v3733e62;
assign v3a70572 = hmaster0_p & v8455ab | !hmaster0_p & v376bbcc;
assign v3a70360 = hmaster1_p & v3a5cdf4 | !hmaster1_p & v8455ab;
assign v37555cb = hmaster3_p & v3a709db | !hmaster3_p & v377324f;
assign v3730217 = hbusreq6_p & v373cdb0 | !hbusreq6_p & v3747ec5;
assign v3769cff = hlock2_p & v3a704f3 | !hlock2_p & v37735a0;
assign v3723efc = hbusreq3_p & v376b4e1 | !hbusreq3_p & v1e37c3e;
assign v376b4a7 = hgrant6_p & v37c039c | !hgrant6_p & v375f53a;
assign v374cca4 = hready_p & v3a570c0 | !hready_p & v3a70291;
assign v3a6da33 = hlock3 & v376ff61 | !hlock3 & v373e5fb;
assign v3a6fdb7 = hmaster0_p & v375d70e | !hmaster0_p & v3774d9a;
assign v3a6fab1 = hbusreq5 & v376a47b | !hbusreq5 & v37494c3;
assign v3a5f4b8 = hmaster2_p & v3a6823d | !hmaster2_p & v3a615c8;
assign v376bb26 = hbusreq1_p & v3747302 | !hbusreq1_p & v3743b9e;
assign v375fcd6 = hmaster2_p & v35b774b | !hmaster2_p & !v3a69591;
assign v377eaa3 = hbusreq4 & v3a70791 | !hbusreq4 & v38073c9;
assign v3724be1 = hlock4_p & v3a60e7e | !hlock4_p & v8455cb;
assign v3a299cd = hbusreq5_p & v3a57ce9 | !hbusreq5_p & v374f691;
assign v373e11e = hmaster3_p & v377097e | !hmaster3_p & v8455ab;
assign v37531ff = hbusreq0_p & v3a70e52 | !hbusreq0_p & v8455b0;
assign v3749840 = hbusreq5 & v376747e | !hbusreq5 & v3806636;
assign v3a6af87 = hbusreq8 & v3a707e7 | !hbusreq8 & v3739f49;
assign v3a6f804 = hgrant2_p & v3a61a3d | !hgrant2_p & !v8455ab;
assign v3736d1d = hmaster1_p & v1e382e7 | !hmaster1_p & v373644e;
assign v3a5eecb = hmaster3_p & v37360c1 | !hmaster3_p & v3751c65;
assign v3a705b0 = hmaster3_p & v8455ab | !hmaster3_p & v3a70ad5;
assign v3378ef7 = hbusreq1_p & v2acb5a2 | !hbusreq1_p & !v8455ab;
assign v372f6a1 = stateA1_p & v3762fc4 | !stateA1_p & !v3723e5f;
assign v37527f2 = hmaster2_p & v3a5a01b | !hmaster2_p & v3a700c7;
assign v37447e1 = hlock4_p & v3806db7 | !hlock4_p & v8455b0;
assign v3a6f0f9 = hlock4_p & v373399e | !hlock4_p & !v8455ab;
assign v3731f7f = hmaster1_p & v3762ca2 | !hmaster1_p & v3730c86;
assign v35b70c9 = hmaster1_p & v3763175 | !hmaster1_p & v3738832;
assign v373b02e = hgrant4_p & v1e37b99 | !hgrant4_p & !v8455ab;
assign v37782ff = hgrant3_p & v8455ab | !hgrant3_p & v3a2a144;
assign v3a5927f = hbusreq2_p & v3a6feb9 | !hbusreq2_p & v3735c5d;
assign v3751bdd = hgrant5_p & v8455c6 | !hgrant5_p & v3730b67;
assign v3a6a261 = hbusreq3_p & v3a6ebbc | !hbusreq3_p & v8455b7;
assign v3724d93 = hgrant0_p & v8455e7 | !hgrant0_p & !v8455ab;
assign v37630ff = hbusreq5_p & v3733228 | !hbusreq5_p & v3770f17;
assign v3a63d83 = hmaster0_p & v375da36 | !hmaster0_p & !v8455ab;
assign v3746a62 = hmaster2_p & v373f911 | !hmaster2_p & v3a6603f;
assign v3a6eb88 = hlock7_p & v373ee66 | !hlock7_p & !v3a7137d;
assign v3a624e7 = hmaster2_p & v374bb76 | !hmaster2_p & v3a6eb7b;
assign v3a71250 = hgrant4_p & v3a6f1ab | !hgrant4_p & v37643af;
assign v2092abf = hmaster1_p & v8455ab | !hmaster1_p & !v37604d6;
assign v3a65da7 = hlock2_p & v3a6a939 | !hlock2_p & !v8455ab;
assign v375abab = hmaster2_p & v3a635ea | !hmaster2_p & v3a707ce;
assign v375c910 = hbusreq4 & v3a6fdc9 | !hbusreq4 & !v8455b5;
assign v37787f5 = hmaster2_p & v3a660af | !hmaster2_p & v3a6f83a;
assign v3a5ddea = hlock6_p & v37652a5 | !hlock6_p & v8455b3;
assign v3768c53 = hmaster1_p & v3a697a5 | !hmaster1_p & v3766de9;
assign v3735da3 = hmaster1_p & v8455ab | !hmaster1_p & v3a71604;
assign a9c905 = hgrant6_p & v374852b | !hgrant6_p & v3a6f10e;
assign v3a7014e = hlock2 & v3a71129 | !hlock2 & v372ae1b;
assign v3a5e3be = hlock4 & v3730052 | !hlock4 & v2acaeda;
assign v375e8aa = hmaster2_p & v37583be | !hmaster2_p & !v3759158;
assign v3a625eb = hmaster0_p & v3a5c369 | !hmaster0_p & v3a6fa45;
assign v376df4c = hmaster2_p & v3a6f55b | !hmaster2_p & v8455ab;
assign v377193a = hlock4_p & v374f87c | !hlock4_p & v8455b0;
assign v373f82c = hbusreq0 & v3a67cfe | !hbusreq0 & v8455ab;
assign v23fde6a = hmaster0_p & v3807aa1 | !hmaster0_p & v3748b83;
assign v373e806 = hbusreq5_p & v3767dc1 | !hbusreq5_p & v3a672e6;
assign bf6063 = hgrant3_p & v8455ab | !hgrant3_p & v3746ac7;
assign v3749fdc = hbusreq6 & v374ccb7 | !hbusreq6 & v8455ab;
assign v3a6b9e8 = hbusreq3 & v3a607af | !hbusreq3 & v8455ab;
assign v375982a = hbusreq7_p & v3771cac | !hbusreq7_p & v3a710cc;
assign v374828c = jx0_p & v3a70360 | !jx0_p & v375c861;
assign v3726a38 = hlock6_p & v3a568f7 | !hlock6_p & !v377395f;
assign v3736ea1 = hgrant6_p & v377e469 | !hgrant6_p & v3741e2a;
assign v3a60584 = hgrant1_p & v8455ab | !hgrant1_p & v376653d;
assign v373c372 = hmaster0_p & v3a62e91 | !hmaster0_p & v3a58b13;
assign v3a706de = hmaster1_p & v3a6fe18 | !hmaster1_p & v372d9e8;
assign b9675e = hbusreq5_p & v3a5e537 | !hbusreq5_p & v8455ab;
assign v375c6f5 = hmaster3_p & v3a6e943 | !hmaster3_p & v3a681f5;
assign b8006a = hlock0_p & v3a66140 | !hlock0_p & v37509af;
assign v37412e9 = hbusreq5_p & v3a6ff4b | !hbusreq5_p & v3a6fd84;
assign v377dc4a = hgrant5_p & v3772470 | !hgrant5_p & v3a61ce5;
assign v37281a4 = hmaster0_p & v8455ab | !hmaster0_p & v8455b2;
assign v3a56c1f = hbusreq5_p & v3765463 | !hbusreq5_p & v3a5c8c9;
assign v3a6f2e7 = hgrant3_p & v3764aea | !hgrant3_p & v375f462;
assign v3739916 = hmaster3_p & v3a6f508 | !hmaster3_p & v35b70d2;
assign v376e431 = hmaster2_p & v3a6f6a4 | !hmaster2_p & v3752dd0;
assign v3747020 = hlock8_p & v376ca61 | !hlock8_p & v377a9b2;
assign v376bded = jx1_p & v3738a45 | !jx1_p & v376a0d2;
assign v37626cc = hmaster0_p & v37689b5 | !hmaster0_p & !v3a6bbc6;
assign v380a188 = hbusreq6_p & v376e1c4 | !hbusreq6_p & v3a6da8a;
assign v3a6582b = hgrant6_p & v3a70cb1 | !hgrant6_p & v372b44a;
assign v3257354 = hbusreq8 & v3a6ba54 | !hbusreq8 & v3a6a95a;
assign v3737c13 = hlock3_p & v360cfe2 | !hlock3_p & v37509c7;
assign v3746e10 = hmaster0_p & v8455ab | !hmaster0_p & v374b6e8;
assign v375649a = hmaster2_p & a568f8 | !hmaster2_p & !v373ad2b;
assign v372f5ec = hbusreq4_p & v3764702 | !hbusreq4_p & v377e172;
assign v3a6fbf1 = hbusreq4_p & v3747a5f | !hbusreq4_p & !v8455ab;
assign v374a20f = jx0_p & v3a6f97f | !jx0_p & v3a6fefd;
assign v3741be8 = hgrant4_p & v8455ab | !hgrant4_p & v372e4e3;
assign v374c63d = jx0_p & v3a70455 | !jx0_p & !v8455ab;
assign v372cdb8 = hmaster2_p & v372988e | !hmaster2_p & v3735ecd;
assign v3a65f4c = hgrant3_p & v375c7b9 | !hgrant3_p & v377ee58;
assign v3a5d532 = locked_p & v8455ab | !locked_p & v3727345;
assign v3a57b57 = hlock5 & v3777bcf | !hlock5 & v3a7107e;
assign v3a5c1a5 = hlock0_p & v37674c1 | !hlock0_p & v8455ab;
assign v3a6f8e7 = hmaster1_p & v3809f73 | !hmaster1_p & v377936c;
assign v374d998 = hmaster3_p & v8455ab | !hmaster3_p & !v3a66c34;
assign v3764a1c = hgrant3_p & v3a70c36 | !hgrant3_p & v375d4fa;
assign v3a70b90 = hmaster1_p & v3a7002c | !hmaster1_p & v3a6d930;
assign v3759602 = hbusreq5_p & v3758ee1 | !hbusreq5_p & v3a70894;
assign v372301d = hmaster2_p & v8455ab | !hmaster2_p & v3a6f832;
assign v373e792 = hgrant5_p & v3778e2d | !hgrant5_p & v377a673;
assign v3a6f511 = hbusreq7_p & v37451c0 | !hbusreq7_p & v3753b93;
assign v3766877 = hlock3 & v3741694 | !hlock3 & v3767a7b;
assign v3757e4b = hgrant2_p & v3a6f99e | !hgrant2_p & v37369e4;
assign v2acafeb = hbusreq8 & v372791c | !hbusreq8 & v3727dab;
assign v37301f5 = hlock0_p & v3a68426 | !hlock0_p & v374e61f;
assign v3a69a42 = hmaster0_p & v3732e45 | !hmaster0_p & d4d3bb;
assign d26e1e = hmaster2_p & v374b1bc | !hmaster2_p & v376495e;
assign v376773b = hbusreq2 & v373f23c | !hbusreq2 & v8455ab;
assign v373e5d9 = hmaster2_p & v3a5c3a0 | !hmaster2_p & v37745c3;
assign v3743698 = hgrant3_p & v37669b4 | !hgrant3_p & v373dafc;
assign v3737ba0 = hmaster1_p & v3a700ee | !hmaster1_p & v3734081;
assign v2acaffd = hbusreq2 & v3757253 | !hbusreq2 & v3a70a7f;
assign v3a713a9 = hgrant5_p & v8455ab | !hgrant5_p & !v376e1ad;
assign v3a57139 = hmaster1_p & v3a29a44 | !hmaster1_p & v37415c3;
assign v374a058 = hmaster1_p & v374c34d | !hmaster1_p & v373f687;
assign v3a70521 = busreq_p & v37771a2 | !busreq_p & v8455e1;
assign v3767f06 = hlock4 & v372a39d | !hlock4 & v3a614cb;
assign v372fa7b = hbusreq6 & v3a6fe6a | !hbusreq6 & !v8455ab;
assign c587b2 = hbusreq8_p & v3a70c77 | !hbusreq8_p & v3a70e09;
assign v3763424 = hmaster2_p & v372988e | !hmaster2_p & v3a71308;
assign v37786a6 = hbusreq0 & v3729785 | !hbusreq0 & v3751a86;
assign v37745c3 = hgrant4_p & v3731d75 | !hgrant4_p & v3724fe7;
assign v373e32a = hgrant2_p & v8455ab | !hgrant2_p & v377d52e;
assign v372b7b1 = hgrant5_p & v8455ab | !hgrant5_p & !v3a5a825;
assign v3a58dce = hlock0 & v374e9c0 | !hlock0 & v2acae4c;
assign v3740bee = hbusreq5 & v377e9a5 | !hbusreq5 & v869938;
assign v3a6fd8a = hlock7_p & v3747465 | !hlock7_p & !v3a7068f;
assign v3a6ff75 = hmaster0_p & v8455ab | !hmaster0_p & v3a6eb26;
assign v37517f7 = hlock7 & v373b2da | !hlock7 & v3a58a3b;
assign v3a6f2ef = hbusreq1 & v3a7042b | !hbusreq1 & v8455ab;
assign v37529f6 = hmaster1_p & v3773eeb | !hmaster1_p & v375bcf7;
assign v373a181 = hgrant3_p & v3741669 | !hgrant3_p & v3a70c38;
assign v8455c7 = hlock5_p & v8455ab | !hlock5_p & !v8455ab;
assign v3a707f0 = hlock5 & v373623d | !hlock5 & v3766101;
assign v375f88a = hbusreq4_p & v374165f | !hbusreq4_p & v3a6ef22;
assign v3a6b306 = hmaster0_p & v3a53c63 | !hmaster0_p & v377de50;
assign v3735077 = hbusreq5 & v373a4ef | !hbusreq5 & v8455ab;
assign v3a704cb = hmaster0_p & v37710fb | !hmaster0_p & !v1e37cf9;
assign v374616d = hgrant6_p & v3723b00 | !hgrant6_p & v3723493;
assign v3741338 = hgrant6_p & v375811e | !hgrant6_p & v8455ab;
assign v3731d06 = hbusreq5 & v3a619c0 | !hbusreq5 & !v8455ab;
assign v373a305 = hlock0 & v3a70ad6 | !hlock0 & v373a196;
assign v377300f = hmaster0_p & v372cdd7 | !hmaster0_p & !v372fba0;
assign v3763b4d = hmaster1_p & v3a635ea | !hmaster1_p & v3748e0c;
assign v39a4e43 = hgrant2_p & v373397b | !hgrant2_p & v8455ab;
assign v3809d8e = hmaster1_p & v2093132 | !hmaster1_p & v37229e6;
assign v377378e = hbusreq0_p & v3a54c77 | !hbusreq0_p & v8455ab;
assign v377665f = hbusreq3 & v37438c9 | !hbusreq3 & v376bade;
assign v3771076 = hgrant4_p & v3a635ea | !hgrant4_p & v3a70749;
assign v375803d = hbusreq5 & v377ed18 | !hbusreq5 & v3a5b514;
assign v37735a0 = hbusreq2 & v3765e46 | !hbusreq2 & v8455ab;
assign v377c7ae = hgrant4_p & v3751389 | !hgrant4_p & v3727986;
assign v373cd68 = hlock6 & v3754777 | !hlock6 & v373081f;
assign v3a6a3ac = hbusreq0 & v3a5e2b2 | !hbusreq0 & v3a6ebaa;
assign v372fb3c = hmaster0_p & v372d905 | !hmaster0_p & v3a6f36d;
assign v3747a7b = hmaster2_p & v8455ab | !hmaster2_p & v3724940;
assign v376614e = hbusreq8_p & v3746fe7 | !hbusreq8_p & v3775498;
assign v3a71046 = hbusreq4 & v373f8d4 | !hbusreq4 & v3760d53;
assign v37536ae = hbusreq0 & v37583be | !hbusreq0 & !v8455ab;
assign v37719c6 = hgrant2_p & v3a5adfd | !hgrant2_p & dac346;
assign v373ea3f = hbusreq3_p & v3a635ea | !hbusreq3_p & v3a6fdef;
assign v3772f0f = hbusreq5 & v3a708c8 | !hbusreq5 & v3a681e8;
assign v376ba62 = hmaster2_p & v3a5d4d0 | !hmaster2_p & v3a70371;
assign v374db9d = hgrant0_p & v3a70070 | !hgrant0_p & !v3a709bf;
assign v373644e = hmaster0_p & v1e382e7 | !hmaster0_p & v3754bd4;
assign v3a69ca2 = hbusreq0 & v374270e | !hbusreq0 & v8455ab;
assign v375bc4b = hbusreq1 & v1e38224 | !hbusreq1 & !v8455ab;
assign v372da87 = hgrant0_p & v8455ab | !hgrant0_p & !v3a64dbd;
assign v3a6d6b8 = hmaster3_p & v373e491 | !hmaster3_p & v8455ab;
assign v3a6bce0 = hmaster2_p & v374b5a8 | !hmaster2_p & v3766202;
assign v377dc20 = hmaster1_p & v3a6ae45 | !hmaster1_p & v3a71083;
assign v377b32c = hgrant8_p & v37366df | !hgrant8_p & v3a6fbb8;
assign v3a6903e = hmaster0_p & v8455c1 | !hmaster0_p & !v3a6f0f4;
assign v3779cb1 = hlock0 & v375cf36 | !hlock0 & v3a6ff8f;
assign v376d559 = hmaster1_p & v3764f06 | !hmaster1_p & !v3a70bbe;
assign v374610d = hbusreq5_p & v3a636ce | !hbusreq5_p & v3726379;
assign v37761dd = hlock8 & v374deba | !hlock8 & v376c69d;
assign v375ab17 = hbusreq4 & v3a608b9 | !hbusreq4 & !v3a6ef42;
assign v3761e45 = hbusreq5 & v3a71196 | !hbusreq5 & v360bc74;
assign v377ad9a = hbusreq3 & v3a6f018 | !hbusreq3 & !v3a5db8a;
assign v3a63d63 = hgrant6_p & v3a62b8d | !hgrant6_p & v3a60882;
assign v37650b8 = hmaster2_p & v3a635ea | !hmaster2_p & v373b166;
assign v3a67d0d = jx0_p & v376d810 | !jx0_p & v375de72;
assign v3a5b539 = hgrant3_p & v373e642 | !hgrant3_p & v1e37e76;
assign v3a706c9 = hmaster0_p & v3a6e4ec | !hmaster0_p & v3a6adff;
assign v376b2f4 = hbusreq5_p & v375d00d | !hbusreq5_p & v37462ae;
assign v3a71476 = hgrant1_p & v8455ab | !hgrant1_p & !v8455b6;
assign v8fc6a0 = hgrant6_p & v375fac6 | !hgrant6_p & !v3760b7a;
assign v3a5bcfd = hmaster2_p & v3770415 | !hmaster2_p & v37522d3;
assign v375924f = hgrant6_p & v3735d71 | !hgrant6_p & v3a6ebd3;
assign v3755d23 = hmaster1_p & v3750746 | !hmaster1_p & v3a7079b;
assign v37320f4 = hbusreq5 & v377da10 | !hbusreq5 & v8455ab;
assign v3a5e2fa = jx0_p & v3774dcd | !jx0_p & v8455ab;
assign v37362fc = hbusreq3_p & v377934a | !hbusreq3_p & v8455b7;
assign v3774f38 = hbusreq6_p & v3807315 | !hbusreq6_p & !v8455ab;
assign v377dcf5 = hmaster0_p & v8455ab | !hmaster0_p & v37308bf;
assign aa8b86 = hmaster0_p & v377aa5d | !hmaster0_p & v375c76b;
assign v3a6ebfb = hgrant6_p & v8455ab | !hgrant6_p & v3745cea;
assign v3756ec2 = hgrant2_p & v3772c92 | !hgrant2_p & v374cc74;
assign v3a6fe8d = hmaster2_p & v3a56642 | !hmaster2_p & v8455ab;
assign v3a7104d = hbusreq4 & v3a6dc08 | !hbusreq4 & v3770769;
assign v376058c = hmaster2_p & v3a62968 | !hmaster2_p & v3a6fac0;
assign v3779749 = hmaster1_p & v37366d5 | !hmaster1_p & v8455ab;
assign v3806f24 = hbusreq6 & v3753dab | !hbusreq6 & v8455ab;
assign v35ba2cb = hgrant5_p & v3a6ef91 | !hgrant5_p & v3a70d2b;
assign v38074ac = hbusreq6_p & v376a166 | !hbusreq6_p & v8455ab;
assign v38078ed = hgrant6_p & v3a5b6de | !hgrant6_p & v372462b;
assign v3a714e4 = hbusreq4 & v3a6a075 | !hbusreq4 & v8455ab;
assign v37651b2 = hmaster0_p & v3724784 | !hmaster0_p & v3762d06;
assign v375d1e1 = hmaster3_p & v376766e | !hmaster3_p & v372da95;
assign v3a573cc = hbusreq4 & v373325f | !hbusreq4 & v8455ca;
assign v376c898 = hmaster2_p & v8455ab | !hmaster2_p & v3733c46;
assign v374e4c0 = hbusreq4 & v377d7dc | !hbusreq4 & !v8455ab;
assign v3a67a78 = hmaster3_p & v3742e95 | !hmaster3_p & v2ff8e61;
assign v3a5a52d = hmaster2_p & v373ca8d | !hmaster2_p & v377e9cd;
assign v377a551 = hgrant6_p & v3a60787 | !hgrant6_p & v3a69df1;
assign v3a7008b = hbusreq0_p & d44200 | !hbusreq0_p & !v3a7151d;
assign v3773881 = hmaster3_p & v376b03a | !hmaster3_p & v3727da5;
assign v3a5f12b = hmaster0_p & v3767e55 | !hmaster0_p & v3a71133;
assign v375a08b = hlock2_p & v372b75b | !hlock2_p & v3739bb2;
assign v3778a76 = hlock4 & v1e37e67 | !hlock4 & v375cfa5;
assign stateG10_3 = !v3937409;
assign v372567b = hbusreq4 & v3a70b51 | !hbusreq4 & v8455ab;
assign v3760f1e = hbusreq2 & v37675f4 | !hbusreq2 & v8455ab;
assign v37630f1 = hbusreq3_p & v3722ee2 | !hbusreq3_p & v8455ab;
assign v3743e4f = hmaster0_p & v3a6b924 | !hmaster0_p & v373d107;
assign v3744104 = hmaster2_p & v8455ab | !hmaster2_p & v375bf96;
assign v3a6f9fa = hmaster1_p & v37514f7 | !hmaster1_p & v37412e9;
assign v3765265 = hgrant4_p & v377cf67 | !hgrant4_p & v3a6a713;
assign v3731cc3 = hbusreq2_p & v377eaf2 | !hbusreq2_p & v374a637;
assign v373303f = hbusreq4 & v3747bea | !hbusreq4 & v3a67691;
assign v35b71cf = hgrant4_p & v8455ab | !hgrant4_p & v3a604bc;
assign v37289d4 = hbusreq3_p & v377eaf2 | !hbusreq3_p & a36a2a;
assign v3a70555 = hmaster1_p & v3a5fc34 | !hmaster1_p & v377f887;
assign v372f885 = hmaster2_p & v3a5f8a2 | !hmaster2_p & v3a68d2e;
assign v3a6f3a3 = hbusreq4_p & v375ab17 | !hbusreq4_p & !v8455ab;
assign v3a61120 = hgrant6_p & v8455ab | !hgrant6_p & v3806e88;
assign v374a60b = hgrant5_p & v3a71360 | !hgrant5_p & v3a60642;
assign v3a64ad6 = hbusreq0 & v3770bed | !hbusreq0 & v3775e82;
assign v3732aa6 = hbusreq0_p & v3729724 | !hbusreq0_p & v3a6f4fc;
assign v3a6603d = hlock0 & v3a635ea | !hlock0 & v3a70a18;
assign v3a60d11 = hmaster0_p & v3774829 | !hmaster0_p & v376df4c;
assign v3a71134 = hgrant4_p & v3a6f3c6 | !hgrant4_p & v3768751;
assign v372baf1 = hbusreq5 & c48c9d | !hbusreq5 & v376b374;
assign v3751b0e = hbusreq1_p & v3a67e2e | !hbusreq1_p & v3a63f05;
assign v3743c22 = hbusreq4 & v3a660b5 | !hbusreq4 & v8455ab;
assign v3a70d26 = hmaster0_p & v3a703f2 | !hmaster0_p & bb4062;
assign v377d770 = hbusreq2_p & v373edc8 | !hbusreq2_p & v377d2e7;
assign v372aff0 = hmaster1_p & v8455e7 | !hmaster1_p & v376d766;
assign v373557e = hmaster1_p & v3773336 | !hmaster1_p & !v375eb79;
assign v37550bd = hmaster1_p & v3a71175 | !hmaster1_p & v3767ff6;
assign v3747de2 = hmaster0_p & v372bcd0 | !hmaster0_p & v3a6c605;
assign v3a69539 = hmaster0_p & v37495ed | !hmaster0_p & v3769923;
assign v375c608 = hgrant6_p & v8455c9 | !hgrant6_p & v3a71271;
assign v947c98 = hbusreq4_p & v3755167 | !hbusreq4_p & v3a70c1a;
assign v3a6f09d = hlock7 & v3a6e231 | !hlock7 & v3765203;
assign v3a6614b = hmaster0_p & v3a5b27f | !hmaster0_p & v3a6ef24;
assign v377f171 = hbusreq4 & a9c905 | !hbusreq4 & v3a6b53f;
assign v3733a19 = hbusreq2_p & v377109d | !hbusreq2_p & v3755b54;
assign v3767704 = hbusreq8 & v3748efb | !hbusreq8 & v8455ab;
assign v32558c4 = hmaster1_p & v376df9f | !hmaster1_p & !v3a588e5;
assign v2ff8e3d = hbusreq8_p & v3a635ea | !hbusreq8_p & v3a5730e;
assign v3768888 = hmaster0_p & v3a606b7 | !hmaster0_p & v3a63033;
assign v373ea71 = hbusreq2_p & v3a63d7a | !hbusreq2_p & v8455ab;
assign v376847d = hbusreq6 & v37395e6 | !hbusreq6 & v8455e7;
assign v3a6f4d6 = hmaster2_p & v372e559 | !hmaster2_p & v8455ab;
assign v377b647 = hgrant5_p & v3743dce | !hgrant5_p & v3a70e5e;
assign v3a70ca1 = hmaster2_p & v3a5bf04 | !hmaster2_p & !v37521ed;
assign a19873 = hmaster0_p & v3a635ea | !hmaster0_p & v3a5e827;
assign v3a5e3d3 = hgrant1_p & v8455ab | !hgrant1_p & v377eaf2;
assign v37676c3 = hmaster0_p & v3a66d94 | !hmaster0_p & v377e8e4;
assign v37787dd = hbusreq5_p & v3736e12 | !hbusreq5_p & v3a5f891;
assign v3a63966 = hbusreq5 & v3a68848 | !hbusreq5 & v374e0a4;
assign v3762e8d = hbusreq5 & v376bbc5 | !hbusreq5 & v3a700eb;
assign v373dfcc = hbusreq3_p & v8455ab | !hbusreq3_p & v3729823;
assign v3a70028 = hgrant6_p & v3a6d30c | !hgrant6_p & v375f462;
assign v3a5b9cd = hmaster0_p & v3a715c1 | !hmaster0_p & v1e37af3;
assign v3a64b1e = hmaster1_p & v8455ab | !hmaster1_p & v374ea7d;
assign v3730cda = hgrant0_p & v8455ab | !hgrant0_p & v375803a;
assign v3a6f4a3 = hbusreq5 & v375129f | !hbusreq5 & v3a65ce7;
assign v3724da7 = hmaster2_p & v3a70957 | !hmaster2_p & v3a6fa8e;
assign v376d078 = hmaster2_p & v3a5971e | !hmaster2_p & v374448e;
assign v3744cea = hlock3 & v3a5a985 | !hlock3 & v373b0a4;
assign v3753b3f = hlock6 & v3a6fd63 | !hlock6 & v37383c0;
assign v373b1c8 = hlock7 & v3a715f9 | !hlock7 & v3a712bc;
assign v2619ad3 = hlock0_p & v377d5d7 | !hlock0_p & v3a6f373;
assign v3a685e1 = hgrant4_p & v373428e | !hgrant4_p & v37416c8;
assign ad2d05 = hbusreq1_p & v37570b7 | !hbusreq1_p & !v3a70056;
assign v374ac3f = hgrant3_p & v3a69c6f | !hgrant3_p & v375635b;
assign v37403cc = hbusreq5_p & v3a70cb2 | !hbusreq5_p & v37343e7;
assign v3a70ca3 = hbusreq4 & v3746d2a | !hbusreq4 & !v3a5b8b0;
assign v3763cfa = hbusreq4 & v3a6fe0d | !hbusreq4 & !v8455b5;
assign v377c34f = hgrant6_p & v377f09a | !hgrant6_p & v3761f22;
assign v37797d5 = hmaster2_p & v3a70d99 | !hmaster2_p & v3729f14;
assign v37508c2 = hlock0 & v377b946 | !hlock0 & v3a70e77;
assign v3735593 = hbusreq1 & v3745f76 | !hbusreq1 & !v8455ab;
assign v373c15e = hmaster3_p & v3a7026e | !hmaster3_p & v377d831;
assign v373822e = hbusreq5 & v3773c70 | !hbusreq5 & v3a63624;
assign v3772696 = hbusreq4_p & v8455cb | !hbusreq4_p & v375989b;
assign v3724121 = hbusreq3_p & v374b0a8 | !hbusreq3_p & v8455ab;
assign v3742b6a = hmaster2_p & v3a5a04c | !hmaster2_p & v3a67a41;
assign v377d19f = hmaster2_p & v3a66aa4 | !hmaster2_p & v372c3df;
assign v3733d02 = hmaster2_p & v372f95b | !hmaster2_p & v375f823;
assign v37246a5 = hgrant6_p & v3759379 | !hgrant6_p & v3764af3;
assign v376022e = hgrant6_p & v37711cc | !hgrant6_p & v2ff8f0a;
assign v3a6fd02 = hmaster2_p & v3725410 | !hmaster2_p & v3a68426;
assign v37590d5 = hmaster1_p & v1e382e7 | !hmaster1_p & v3746ab7;
assign v3765722 = hgrant2_p & v8455e1 | !hgrant2_p & !v3a65f4c;
assign v374c058 = jx1_p & v3a64103 | !jx1_p & v3739885;
assign v377da08 = hbusreq8_p & v3728cb3 | !hbusreq8_p & v373c56f;
assign v3741ccb = hlock4 & v37269f6 | !hlock4 & v373340d;
assign v374dce0 = hbusreq4 & v8455e1 | !hbusreq4 & !v8455ab;
assign v3a67b76 = hmaster0_p & v3a6452e | !hmaster0_p & v3767e71;
assign v373676d = hmaster0_p & v3a5a01b | !hmaster0_p & v37527f2;
assign v377f80c = hmaster1_p & v35b7168 | !hmaster1_p & v3a707c5;
assign v3742210 = hbusreq8 & v373b1c8 | !hbusreq8 & v3a6fb20;
assign v377a615 = hmaster2_p & v3a661fe | !hmaster2_p & v3a713df;
assign v37337e7 = hbusreq5 & v3a5ebbf | !hbusreq5 & v374a36b;
assign v3733862 = hbusreq6 & v372ee9a | !hbusreq6 & v3a6be44;
assign v3a6d9ac = hmaster2_p & v3a5a807 | !hmaster2_p & v1e3787a;
assign v3a6eb9d = hmaster1_p & v3a7066b | !hmaster1_p & v3a70641;
assign v372b858 = hlock4 & v373c7db | !hlock4 & v3729b6a;
assign c52384 = hmaster0_p & v3a5fee0 | !hmaster0_p & v3753b80;
assign v3777ff3 = hmastlock_p & v376bd2a | !hmastlock_p & v8455ab;
assign v3377af7 = hlock3 & v37518fa | !hlock3 & v3770af1;
assign v3729ae4 = hgrant0_p & v3a61b63 | !hgrant0_p & v37798c3;
assign v3731741 = hmaster2_p & v8455e7 | !hmaster2_p & !v372fc81;
assign be54b2 = hgrant4_p & v8455c2 | !hgrant4_p & v3a6ff08;
assign v372f9b4 = hbusreq5_p & v3769d07 | !hbusreq5_p & !v373b6ba;
assign v3a5def2 = hgrant6_p & v38064e4 | !hgrant6_p & d4de60;
assign v3a70b1e = hbusreq6 & v3a68cc4 | !hbusreq6 & v8455ab;
assign v3a695ec = hmaster3_p & v377c0fa | !hmaster3_p & v3a6879a;
assign v3758c3d = hbusreq5 & v3759263 | !hbusreq5 & v3a6ff33;
assign v3a6f842 = hbusreq2_p & v3738d68 | !hbusreq2_p & v35772a6;
assign v3a6eb72 = hmaster2_p & v3a635ea | !hmaster2_p & v376bb26;
assign v3a71082 = hmaster1_p & v37284f3 | !hmaster1_p & v373f691;
assign v3a65d4e = hbusreq2_p & v37765e1 | !hbusreq2_p & v37730bf;
assign v3a70c34 = hbusreq6 & v3a6fbd0 | !hbusreq6 & !v37238b1;
assign v37532f0 = hmaster1_p & v374a11d | !hmaster1_p & v3a6fd84;
assign v3a674fa = hmaster0_p & v376025f | !hmaster0_p & v374abee;
assign v3a6eaee = hbusreq7_p & v3733138 | !hbusreq7_p & !v8455ab;
assign v3a7055a = hmaster0_p & v3a6c4e4 | !hmaster0_p & v3a659b2;
assign v37368e1 = hbusreq4_p & v3763b0a | !hbusreq4_p & v3757a57;
assign v372ad4e = hbusreq4_p & v9773b9 | !hbusreq4_p & v8455ab;
assign v3740811 = hbusreq7_p & v3775806 | !hbusreq7_p & v37585c9;
assign v375787b = hmaster2_p & v8455ab | !hmaster2_p & v37326a1;
assign v3a6b77d = hgrant3_p & v3a696ed | !hgrant3_p & v3a57cb4;
assign v3a70f61 = hbusreq8 & v3a63b26 | !hbusreq8 & v377e30e;
assign v3739391 = hlock4 & v3723f2a | !hlock4 & v3765e6a;
assign v3754260 = hbusreq2_p & v3a70e65 | !hbusreq2_p & v377ab2c;
assign v373c8c3 = hbusreq8_p & v373f8c8 | !hbusreq8_p & v3a6f06a;
assign v3a70e0c = hgrant6_p & v8455ab | !hgrant6_p & v3a56d06;
assign v376bf04 = hbusreq1 & v1e38224 | !hbusreq1 & v8455ab;
assign v3a6f3da = hlock6 & v376f584 | !hlock6 & v3a70a50;
assign v37635f0 = hmaster2_p & v377adf5 | !hmaster2_p & v3736847;
assign v3744590 = hbusreq2 & v3a6143b | !hbusreq2 & !v8455b5;
assign v39a4e5f = hbusreq1_p & v3a635ea | !hbusreq1_p & !v3a6830c;
assign v3a7131d = hmaster1_p & v375a8d6 | !hmaster1_p & v3a705f1;
assign v3a5d8bc = hmaster2_p & v37570f8 | !hmaster2_p & v3724af9;
assign v3729516 = hbusreq5_p & v3764628 | !hbusreq5_p & v37523dd;
assign v373dc5a = hbusreq5 & v373a3e7 | !hbusreq5 & c79715;
assign v3a6ebd0 = hmaster1_p & v3753418 | !hmaster1_p & v377c35c;
assign dc6ea3 = hgrant0_p & v8455b0 | !hgrant0_p & v377c17f;
assign v375bfdf = hgrant4_p & v3a5bccf | !hgrant4_p & v3a60d86;
assign v3a53f53 = hbusreq4 & v3a58d22 | !hbusreq4 & !v8455ca;
assign v3a5b6de = hbusreq3_p & v3762502 | !hbusreq3_p & v3a5bb64;
assign v3733467 = hbusreq4_p & v372468b | !hbusreq4_p & v35772a6;
assign v3755596 = hbusreq7_p & v3723780 | !hbusreq7_p & v376ffa7;
assign v373a0e2 = hgrant5_p & v3a70f30 | !hgrant5_p & v3a6f30a;
assign v3a6913c = hbusreq5 & v3a62250 | !hbusreq5 & v3a70582;
assign v3739702 = hbusreq5_p & v373f042 | !hbusreq5_p & v8455e7;
assign v372c83a = hgrant5_p & v375f0d4 | !hgrant5_p & v374aa4f;
assign v3727fa7 = hmaster0_p & v373399e | !hmaster0_p & v3749e68;
assign v377d904 = hmaster1_p & v37644ff | !hmaster1_p & v3724798;
assign v3a5e660 = hgrant5_p & v8455c6 | !hgrant5_p & v3a655e9;
assign v3a2abd2 = hgrant6_p & v3a6f22e | !hgrant6_p & v3764462;
assign v3a54cd9 = hlock7_p & v3a6f1db | !hlock7_p & v3a70581;
assign v37778e2 = hgrant6_p & v3743cd6 | !hgrant6_p & v3a69e8c;
assign v373f785 = hgrant2_p & v8455e7 | !hgrant2_p & v35b70e6;
assign v3766d10 = hbusreq4 & v372fc81 | !hbusreq4 & !v8455ab;
assign v376352a = hbusreq4 & v377da37 | !hbusreq4 & v8455ab;
assign v3730169 = hmaster2_p & v3a5fe3c | !hmaster2_p & v1e3735b;
assign v3a6f4f1 = hgrant6_p & v375f2ec | !hgrant6_p & v3a59d47;
assign v377d142 = hbusreq0 & v375b429 | !hbusreq0 & v372ed51;
assign v374ab34 = hmaster0_p & v37667ed | !hmaster0_p & !v3758c58;
assign v9fecca = hbusreq7 & v3779b3a | !hbusreq7 & v3a6cf88;
assign v3a6fdf9 = hmaster1_p & v37445e2 | !hmaster1_p & v3a61cd7;
assign v3766d1b = hbusreq6 & v3755dcd | !hbusreq6 & !v8455bd;
assign v3a70ddd = hmaster2_p & v37476bd | !hmaster2_p & v23fd83f;
assign v376b5ac = hbusreq1 & v376d9ad | !hbusreq1 & v8455ab;
assign v3a70f5d = hgrant6_p & v375564e | !hgrant6_p & v376070d;
assign v3776767 = hmaster2_p & v8455ab | !hmaster2_p & !v373dfff;
assign v3a6fa55 = hbusreq4 & v374b320 | !hbusreq4 & v3a6bf41;
assign v3a70129 = hmaster1_p & v8455ab | !hmaster1_p & v37325eb;
assign v3a69591 = hbusreq1_p & v3a6667e | !hbusreq1_p & !v8455ab;
assign v3724488 = hmaster1_p & v3a701b7 | !hmaster1_p & v8455ab;
assign v3a6f378 = hbusreq4 & v3771607 | !hbusreq4 & v3737028;
assign v1e379fa = hbusreq5_p & v3a64931 | !hbusreq5_p & v3776abb;
assign v3731b41 = hgrant4_p & v8455ab | !hgrant4_p & v3a640ff;
assign v3a7049d = hmaster3_p & v2acaf9d | !hmaster3_p & v3a70766;
assign v3a70978 = hbusreq5_p & v37533c8 | !hbusreq5_p & v3a575dc;
assign v37281fb = hmaster2_p & v3768f0c | !hmaster2_p & v8455b3;
assign v3a69d9b = stateG10_1_p & v8455ab | !stateG10_1_p & v373602d;
assign v376b94a = jx0_p & v3a70ae5 | !jx0_p & v3a6f773;
assign v376fdbe = hbusreq5_p & v3a70f93 | !hbusreq5_p & v3a5fc48;
assign v3a7081e = hlock6_p & v3766ea9 | !hlock6_p & v8455b0;
assign v3a71243 = hmaster2_p & v3771c85 | !hmaster2_p & v374d52a;
assign v3a5f162 = hbusreq4_p & v3a6d5e9 | !hbusreq4_p & v376aa10;
assign v3750fc8 = busreq_p & v37386a9 | !busreq_p & v8455ab;
assign v377a9a1 = hgrant4_p & v8455ab | !hgrant4_p & v3750b0d;
assign v3a70642 = hbusreq5 & v39eb033 | !hbusreq5 & v3764a8a;
assign v377ed5e = hmaster2_p & v8455bb | !hmaster2_p & !v3a70e4f;
assign v3734ef4 = hgrant8_p & v372aeef | !hgrant8_p & v3a6fc95;
assign v3a6ffee = hlock5 & v3759c23 | !hlock5 & v3743f7a;
assign v3a6491d = hmaster0_p & v37548f4 | !hmaster0_p & !v373a246;
assign aa9893 = hmaster0_p & v3726f6b | !hmaster0_p & v3a6f53a;
assign v37c36c4 = hbusreq5_p & v375cf11 | !hbusreq5_p & v37626cc;
assign ae13ec = hgrant3_p & v8455e7 | !hgrant3_p & v3767d7c;
assign v37762b6 = hgrant2_p & v37346be | !hgrant2_p & !v37464f0;
assign v3a71645 = hmaster2_p & v37782c9 | !hmaster2_p & !v3a64349;
assign v3a70115 = hbusreq2_p & v3a60787 | !hbusreq2_p & !v377cfd9;
assign v377e31b = hgrant4_p & v8455ab | !hgrant4_p & v38097db;
assign v3a7138e = hlock5 & v3a6fd22 | !hlock5 & v373a6f8;
assign v3732b1d = hmaster1_p & v3a67c30 | !hmaster1_p & v374b0a3;
assign v372a4c3 = hgrant2_p & v3725f98 | !hgrant2_p & v3a6f557;
assign v3723f24 = hgrant3_p & v8455ab | !hgrant3_p & v3a7109d;
assign v372b7a5 = hmaster0_p & v373b98a | !hmaster0_p & v8455ab;
assign v3739892 = hbusreq4 & v377c38c | !hbusreq4 & v8455ab;
assign v374650b = hgrant5_p & v8455ab | !hgrant5_p & v3a6f4d5;
assign v3764caa = hlock5 & v377de7f | !hlock5 & v3769069;
assign v3a712c2 = hmaster2_p & v37784b9 | !hmaster2_p & v3a6c0c5;
assign v3765c85 = hbusreq2 & v3a6e3bb | !hbusreq2 & v3a5b2fd;
assign v37326a1 = hgrant4_p & v37346be | !hgrant4_p & v37500c2;
assign v3752ab6 = hmaster0_p & v2ff9190 | !hmaster0_p & v3a71502;
assign v3741b61 = hmaster1_p & v3a635ea | !hmaster1_p & v37759a7;
assign v1e37d2a = hlock3_p & v2acafff | !hlock3_p & v372538b;
assign v3a6f6a2 = hgrant6_p & v3723b0c | !hgrant6_p & v3754aa3;
assign v1e379b9 = hmaster0_p & v8455dd | !hmaster0_p & !v8455ab;
assign v375f370 = hbusreq0 & v3a5899d | !hbusreq0 & v37c0158;
assign v3a6ff69 = hbusreq5_p & v3735331 | !hbusreq5_p & v3a574d6;
assign v3765324 = jx0_p & v3747367 | !jx0_p & v37652ae;
assign v8455c3 = hlock4_p & v8455ab | !hlock4_p & !v8455ab;
assign v3a6f92d = hbusreq7 & v374c297 | !hbusreq7 & v3768734;
assign v3a70df1 = hgrant0_p & v3770559 | !hgrant0_p & !v3a7044c;
assign v375b9dc = hmaster1_p & v3762e13 | !hmaster1_p & v372d30b;
assign v3a652db = hlock8 & v3737808 | !hlock8 & v3a70719;
assign v390071e = hmaster2_p & v375144b | !hmaster2_p & v376629a;
assign v37725b5 = hmaster1_p & v3807a4a | !hmaster1_p & v3a6574d;
assign v377f5c9 = jx1_p & v3778f81 | !jx1_p & v3a649c2;
assign v3757adc = hbusreq4 & v3a61f9b | !hbusreq4 & v3737028;
assign v3a60181 = hlock4_p & v3766238 | !hlock4_p & v3768202;
assign v376b2a2 = hbusreq4 & v373abae | !hbusreq4 & v3a6efea;
assign v3a66140 = hbusreq1_p & v373df14 | !hbusreq1_p & v37328a1;
assign v3a6f948 = hmaster0_p & v3a6f94c | !hmaster0_p & v3747971;
assign v3a703de = hgrant2_p & v9da9d2 | !hgrant2_p & v3736ebd;
assign v3a55efa = hlock6 & v3725360 | !hlock6 & v373a568;
assign v3771ab9 = hlock6 & v373f953 | !hlock6 & v3a582d6;
assign v3a62826 = hbusreq1_p & v376045b | !hbusreq1_p & v8455ab;
assign v3a70c97 = hbusreq3 & v3807107 | !hbusreq3 & v8455ab;
assign v3a5cdc1 = hmaster2_p & v8455ab | !hmaster2_p & v37672aa;
assign v3743c90 = jx0_p & v377b6ce | !jx0_p & !v37691b8;
assign v374a7de = hmaster0_p & v8455ab | !hmaster0_p & v376fefa;
assign v3a68ee5 = hbusreq5 & v3a6f86b | !hbusreq5 & v375456e;
assign v377a2e4 = hburst1 & v3a299c1 | !hburst1 & v1e3746e;
assign v3773c57 = hgrant0_p & v3775b81 | !hgrant0_p & v8455ab;
assign v3768e52 = hmaster0_p & v3a6ebf7 | !hmaster0_p & v8455ab;
assign v3774399 = hbusreq5_p & v37510fb | !hbusreq5_p & v37591bc;
assign v377cb85 = hmaster1_p & v3730e7d | !hmaster1_p & v3774841;
assign v377873a = hgrant6_p & v377f09a | !hgrant6_p & !v3779f6b;
assign v3a5872b = hbusreq2_p & v3731b72 | !hbusreq2_p & !v8455ab;
assign v372d2d2 = hbusreq7_p & v3757506 | !hbusreq7_p & v372e6d0;
assign v3806cd2 = hbusreq6_p & v35b9d52 | !hbusreq6_p & v3733ea2;
assign v373d214 = hbusreq4_p & v3743de1 | !hbusreq4_p & v372cc0a;
assign v3a6fc6e = stateA1_p & v8455ab | !stateA1_p & v3a5a496;
assign v372c09a = hmaster1_p & v3777f05 | !hmaster1_p & v372d035;
assign v373281b = hmaster3_p & v373c8c3 | !hmaster3_p & v3a688f9;
assign v3747d0a = hbusreq7_p & v37249fe | !hbusreq7_p & v3a706a3;
assign v3a5514a = hmaster0_p & v373d0d3 | !hmaster0_p & v3a7062d;
assign v3a53b8b = hmaster0_p & v373e6d2 | !hmaster0_p & v372dcff;
assign v376a44f = hmaster2_p & v3747302 | !hmaster2_p & v375da10;
assign acc1e3 = hbusreq6_p & v375022e | !hbusreq6_p & v8455ab;
assign v3a64087 = hgrant2_p & v377182c | !hgrant2_p & v38065aa;
assign v3a580fb = hmaster2_p & v3a712dd | !hmaster2_p & v3a6f3e9;
assign v3765261 = hgrant2_p & v8455ab | !hgrant2_p & v3a5b614;
assign v3741797 = hgrant3_p & v8455ab | !hgrant3_p & v3722f88;
assign v37766d3 = jx0_p & v3756ce5 | !jx0_p & v3776d3e;
assign v3a61ce5 = hmaster1_p & v3a6f4d7 | !hmaster1_p & v3a6aac8;
assign v376f148 = hgrant0_p & v3744d52 | !hgrant0_p & v3a56417;
assign v3a6f244 = hgrant4_p & v3a6a22c | !hgrant4_p & v3a5fbad;
assign v3577306 = stateA1_p & v8455e1 | !stateA1_p & !v3a635ea;
assign v376da3f = hmaster2_p & v39a4ca8 | !hmaster2_p & !v8455ab;
assign v3a6e7d8 = hlock4 & v3a70481 | !hlock4 & v3a70cb1;
assign v3a58139 = hmaster0_p & v373ce86 | !hmaster0_p & v3733e77;
assign v37756ab = hbusreq4_p & v3775999 | !hbusreq4_p & v3a69c57;
assign v3a6f2ce = hmaster0_p & v377d1dc | !hmaster0_p & v23fd83c;
assign v37349e4 = hlock5 & v375e5ed | !hlock5 & v37357d0;
assign v373de66 = hlock2_p & v3735e39 | !hlock2_p & v376d856;
assign v373250a = hlock7_p & v375e5a6 | !hlock7_p & !v8455ab;
assign v3a704f8 = hbusreq2 & v39a537f | !hbusreq2 & !v8455ab;
assign v373380d = hmaster2_p & v3763f95 | !hmaster2_p & v3a70c39;
assign v3747d42 = hlock5 & v3728867 | !hlock5 & v3a66ca0;
assign v377ae81 = hlock4 & v3735444 | !hlock4 & v3a627a7;
assign v3a70dcb = hmaster0_p & v3a635ea | !hmaster0_p & v3a5b87f;
assign v3a58d5f = hmaster1_p & v3a6fcdc | !hmaster1_p & v374bac7;
assign v373f10d = hbusreq0 & v3a5948d | !hbusreq0 & v377a5df;
assign v3a5f80f = hmaster1_p & v3a635ea | !hmaster1_p & v3777142;
assign v3a61081 = hbusreq6_p & v372fa7b | !hbusreq6_p & !v8455ab;
assign v3748301 = hmaster1_p & v89a228 | !hmaster1_p & v3a62ad8;
assign v3a63d05 = hbusreq5_p & v39ebb2e | !hbusreq5_p & !v375a2ff;
assign v3a6fd64 = hlock5_p & v373f042 | !hlock5_p & !v8455ab;
assign v3a712fd = hbusreq0 & v3a65503 | !hbusreq0 & v376c5f5;
assign v374df3c = hgrant5_p & v372ab63 | !hgrant5_p & v3a53cf1;
assign v3765b08 = hbusreq3_p & v3736a92 | !hbusreq3_p & v3753fe0;
assign v3774deb = hmaster2_p & v37793e4 | !hmaster2_p & v3763a86;
assign v375b4cb = hmaster0_p & v3a70d99 | !hmaster0_p & v3724e7d;
assign v374ff28 = hlock5_p & v374a8da | !hlock5_p & v8455ab;
assign v3778648 = hbusreq4 & v3a6ff87 | !hbusreq4 & v8455ab;
assign v3a6eb76 = hbusreq6_p & v3737075 | !hbusreq6_p & v3a698c3;
assign v3a70455 = hgrant5_p & v3a6437e | !hgrant5_p & v375d2ee;
assign v3744039 = hmaster2_p & v35772a6 | !hmaster2_p & v3a66a01;
assign v377b0d8 = hmaster0_p & v3a635ea | !hmaster0_p & v3762d09;
assign v375d38f = hbusreq2_p & v374f860 | !hbusreq2_p & !v372fbf8;
assign v3751ad8 = hgrant3_p & v8455ab | !hgrant3_p & !v3a703a1;
assign v3752c04 = hlock0_p & v3a70385 | !hlock0_p & !v8455ab;
assign v3a70e93 = hlock0_p & v3735e39 | !hlock0_p & v374abf3;
assign v376442b = hlock3_p & v374bb56 | !hlock3_p & !v8455ab;
assign v3a5c5f4 = hbusreq2_p & v377cfd9 | !hbusreq2_p & !v372ee7e;
assign v3a59cae = hmaster2_p & v3a56531 | !hmaster2_p & v3752fbc;
assign v37744d9 = hmaster2_p & v8455ab | !hmaster2_p & v3a5bea0;
assign v374a4a0 = hbusreq6 & v3a6f5fb | !hbusreq6 & v8455ab;
assign v3779c8e = hbusreq5 & v37536fd | !hbusreq5 & v3a58fe2;
assign v3a706b1 = hbusreq3 & v3a6ffca | !hbusreq3 & v8455ab;
assign v3759b61 = hbusreq8_p & v373d6dd | !hbusreq8_p & v375c1fd;
assign v3a70298 = hbusreq5_p & v3760bfa | !hbusreq5_p & v3a70f8c;
assign v373f6b1 = hmaster1_p & v3807f45 | !hmaster1_p & v377c71e;
assign v3753b1b = hbusreq5 & v3724ff0 | !hbusreq5 & v8455ab;
assign v376b397 = hgrant4_p & v38072fd | !hgrant4_p & v8455ab;
assign v3a7094b = hmaster0_p & v8455ab | !hmaster0_p & v377b311;
assign v3741020 = hbusreq6_p & v3a56898 | !hbusreq6_p & v3a71219;
assign v3a6a95e = hbusreq6_p & v3766218 | !hbusreq6_p & v3a703d3;
assign v3a6fd35 = jx1_p & v3a54789 | !jx1_p & v3747cfc;
assign v3737028 = hlock4_p & v3773ee6 | !hlock4_p & v8455b3;
assign v3772185 = hgrant4_p & v3739896 | !hgrant4_p & v373ccc7;
assign v374c6e1 = hgrant6_p & v3760e2e | !hgrant6_p & v375208a;
assign v3a6d2e2 = hbusreq7 & v3743c84 | !hbusreq7 & v372d827;
assign v3762892 = hbusreq7 & v3724d8c | !hbusreq7 & v37786c6;
assign v39a4dd7 = hgrant0_p & v3a6eeb5 | !hgrant0_p & v375b80e;
assign v37750e4 = hbusreq5_p & v374930c | !hbusreq5_p & v3a62f50;
assign v3730bb7 = stateG10_1_p & v8455ab | !stateG10_1_p & v3744c95;
assign v3a7011e = hgrant2_p & v8455ab | !hgrant2_p & v3a6a82a;
assign v3a714c7 = hmaster2_p & v3a6206d | !hmaster2_p & !v8455ab;
assign v375bfc4 = hgrant5_p & v3a6f6e0 | !hgrant5_p & v3806ed4;
assign v375b4a7 = hbusreq2_p & v377ac7e | !hbusreq2_p & v37686c1;
assign v3722af7 = hbusreq7 & v3766607 | !hbusreq7 & v3774bad;
assign v23fe312 = hlock7 & v3a71048 | !hlock7 & v37305c2;
assign v372b8a3 = hbusreq5_p & v3a706bd | !hbusreq5_p & !v8455ab;
assign v3a6f195 = hmaster2_p & v209312a | !hmaster2_p & v372cac6;
assign v3a66778 = hmaster2_p & v1e37370 | !hmaster2_p & v3a6b1d4;
assign v2acae68 = hbusreq3_p & v3a70aa2 | !hbusreq3_p & v377bdd6;
assign v3723dac = hlock0 & v375aea6 | !hlock0 & v372af57;
assign v3a60026 = hmaster1_p & v3a694b9 | !hmaster1_p & !v377b8fb;
assign v373a3dd = hbusreq3_p & v3725cbf | !hbusreq3_p & v376905f;
assign v3730749 = hgrant4_p & v3747c4c | !hgrant4_p & v3740f3d;
assign v3a5733c = hbusreq5_p & v3768739 | !hbusreq5_p & !v37766cf;
assign v3a6a934 = hgrant6_p & v8455ab | !hgrant6_p & v3a5ee6e;
assign v376cd19 = hbusreq7 & v372e8ae | !hbusreq7 & v37431a0;
assign v38067bb = hbusreq7 & v375be57 | !hbusreq7 & v3808f75;
assign bc8871 = hmaster0_p & v8455e7 | !hmaster0_p & v374e692;
assign v3a6d1a5 = hmaster2_p & v376dc26 | !hmaster2_p & v37287d8;
assign v3735afb = hbusreq4_p & v8455bf | !hbusreq4_p & v375590f;
assign v376ee20 = hmaster2_p & v3a70f68 | !hmaster2_p & v3a6f8e6;
assign v3759c80 = hbusreq5_p & v3723f71 | !hbusreq5_p & !v8455ab;
assign v37798c3 = hlock0_p & v3766e3a | !hlock0_p & v3a713d8;
assign v3a6ffff = hlock6 & v3a7118a | !hlock6 & v3a703d0;
assign v3a5d079 = hgrant4_p & v37c3782 | !hgrant4_p & v373855c;
assign v3a556c2 = hmaster3_p & v376a054 | !hmaster3_p & v8455ab;
assign v3a58b9f = hmaster2_p & v3a5d9e7 | !hmaster2_p & v37395e8;
assign v377de07 = hmaster0_p & v3768589 | !hmaster0_p & v3750b22;
assign v375d17d = hbusreq7_p & v37260af | !hbusreq7_p & v377546d;
assign ca1199 = hbusreq6 & v37457fb | !hbusreq6 & v8455e7;
assign v3a693af = hgrant0_p & v8455ab | !hgrant0_p & v3723ac5;
assign v3a70280 = hmaster3_p & v3a6fb53 | !hmaster3_p & v3a6b213;
assign v377a337 = hmaster0_p & v3a6ffca | !hmaster0_p & v3a6dc57;
assign v3a7057b = locked_p & v8455ab | !locked_p & !v377ec9b;
assign v3758809 = hmaster1_p & v3a61516 | !hmaster1_p & v8455ab;
assign v3a70e4f = hlock2_p & v373ad95 | !hlock2_p & v8455ab;
assign v372f1b8 = hlock4 & v37752c8 | !hlock4 & v3a711e2;
assign v37761fe = hbusreq4 & v3a6ecf6 | !hbusreq4 & v377e698;
assign v3728506 = hbusreq3_p & v23fe379 | !hbusreq3_p & v374f609;
assign v372a954 = hbusreq4 & v375e682 | !hbusreq4 & v8455ab;
assign v3a704c2 = hbusreq6 & v374cab9 | !hbusreq6 & v37674c1;
assign v37334c5 = hmaster2_p & v3740171 | !hmaster2_p & v3a6f7bf;
assign v3a6d0af = hmaster0_p & v3a635ea | !hmaster0_p & v3a5b912;
assign v3750deb = hbusreq1_p & v3773091 | !hbusreq1_p & v3754586;
assign v3a6eef0 = hbusreq7_p & v37681ec | !hbusreq7_p & v3732a95;
assign v3a70728 = hbusreq4 & v376dc16 | !hbusreq4 & v373abde;
assign v37609ac = hlock3 & v3769404 | !hlock3 & v3738397;
assign v9a3ffa = hmaster0_p & v3a5bd76 | !hmaster0_p & v3726983;
assign v373d42f = hmaster0_p & v3755000 | !hmaster0_p & v3731c2f;
assign v3a6f3e9 = hgrant4_p & v1e37b99 | !hgrant4_p & !v372516b;
assign v376e1b7 = hbusreq2_p & v374f0c1 | !hbusreq2_p & v3a669ac;
assign v3a70b3c = hmaster0_p & v3a6ffca | !hmaster0_p & v3732772;
assign v3a6ffc3 = hmaster1_p & v3a71110 | !hmaster1_p & v372993f;
assign v3a6fdc7 = hlock4_p & v3a5980d | !hlock4_p & v8455b7;
assign v37274be = hbusreq2 & v375911a | !hbusreq2 & v3a69487;
assign v3a70a97 = hmaster1_p & v3775dbc | !hmaster1_p & v3774391;
assign v3a6c605 = hbusreq4_p & v37406d2 | !hbusreq4_p & v3753dab;
assign v374bf71 = hgrant3_p & v3723430 | !hgrant3_p & v3a6e438;
assign v3748990 = hmaster0_p & v3763f38 | !hmaster0_p & v377b774;
assign v3759506 = hgrant4_p & v3a53eeb | !hgrant4_p & v3a70c9a;
assign v373d5dc = hbusreq0 & v3734247 | !hbusreq0 & v3a60aca;
assign v3724270 = hbusreq4_p & v3a58b5a | !hbusreq4_p & v8455ab;
assign v3775a92 = hgrant6_p & v3809752 | !hgrant6_p & v8455ab;
assign v3a563aa = hready_p & v3a6307d | !hready_p & !v37771cc;
assign v37724fc = hlock5 & v375803d | !hlock5 & v373dac4;
assign v377246b = hmaster0_p & v3741baf | !hmaster0_p & v3a702e9;
assign v3a64e91 = hbusreq3_p & v375bc6e | !hbusreq3_p & v374fa0a;
assign v3749e68 = hmaster2_p & v3a70530 | !hmaster2_p & v377af44;
assign v376ce17 = hmaster1_p & v8455ab | !hmaster1_p & v375a2a3;
assign v3730c49 = hgrant5_p & v8455ab | !hgrant5_p & v3752d9f;
assign v3a6fa72 = hbusreq6_p & v3a5846c | !hbusreq6_p & b72b90;
assign v37349f9 = hbusreq5 & v37560ef | !hbusreq5 & v375b0ad;
assign v37650d7 = hbusreq5_p & v3762873 | !hbusreq5_p & v37738be;
assign v3765f9e = hmastlock_p & v3778565 | !hmastlock_p & v8455ab;
assign v3a5c16e = hmaster2_p & v3a7066c | !hmaster2_p & v37793a4;
assign v3724002 = hbusreq2_p & v3a6f1b2 | !hbusreq2_p & v3a605bd;
assign v3a58723 = hmaster1_p & v3a70484 | !hmaster1_p & v8f1dd1;
assign v37712c2 = hlock8 & v3773b66 | !hlock8 & v37734d2;
assign v372d8ff = hbusreq5_p & v3a6efe8 | !hbusreq5_p & v3a7112c;
assign v3773fc7 = hgrant4_p & v8455ab | !hgrant4_p & v3751e80;
assign v374d695 = hbusreq5 & v3a6fc38 | !hbusreq5 & v3738844;
assign v3a618ea = hgrant5_p & v3744f6f | !hgrant5_p & v373ac65;
assign v374cb86 = hbusreq8_p & v3a57ef6 | !hbusreq8_p & v3a616aa;
assign v373112c = hmaster0_p & v3a70a7e | !hmaster0_p & !v3a6607f;
assign v3a711e0 = hgrant6_p & v3750c38 | !hgrant6_p & v3a5a397;
assign v375ae53 = hlock7_p & v3a70017 | !hlock7_p & !v8455ab;
assign v377972c = hmaster2_p & v377b92f | !hmaster2_p & v3a6feee;
assign v3768723 = hbusreq4 & v374d0f9 | !hbusreq4 & v374f35a;
assign v37475f4 = hgrant5_p & v3743831 | !hgrant5_p & v3a7166a;
assign v3a6a82a = hgrant3_p & v8455ab | !hgrant3_p & v3a70452;
assign v3776ae5 = hmaster0_p & v375afe9 | !hmaster0_p & v3a71518;
assign v3a6f625 = hbusreq7_p & v37343f6 | !hbusreq7_p & v37664b4;
assign c98bc3 = hbusreq5_p & v3756b5c | !hbusreq5_p & v3a70932;
assign v3773092 = stateA1_p & v3757c6f | !stateA1_p & a81487;
assign v375c01e = hlock5 & v3a656be | !hlock5 & v3a60fee;
assign v380854b = hgrant3_p & v35b7299 | !hgrant3_p & !v3772ab1;
assign v377818c = hbusreq4 & v373e2c3 | !hbusreq4 & v8455ab;
assign v3a702f8 = hbusreq2_p & v38072fd | !hbusreq2_p & v3a6fb9d;
assign v377a525 = hlock8 & v3779ba9 | !hlock8 & v374148a;
assign v3a65104 = hbusreq4_p & v37425c6 | !hbusreq4_p & v3a702c2;
assign v3a6900b = hgrant3_p & v3a6251b | !hgrant3_p & v3736a92;
assign v3733599 = hbusreq0 & v3754f0f | !hbusreq0 & v373de53;
assign v37424df = hmaster2_p & v3739b80 | !hmaster2_p & !v3766ff7;
assign v3a6fbe1 = hbusreq4 & v8455ab | !hbusreq4 & !v38097d8;
assign v23fe0c2 = hbusreq4_p & v375d149 | !hbusreq4_p & v3a635ea;
assign v3a6094b = hbusreq5 & v3a6fec1 | !hbusreq5 & v3771e69;
assign v377af34 = hbusreq6_p & v375a766 | !hbusreq6_p & v8455ab;
assign v3a71162 = hgrant4_p & v3a71267 | !hgrant4_p & v37512f3;
assign v3728dc7 = hgrant4_p & v3770559 | !hgrant4_p & v374ad82;
assign v3756a6a = hmaster2_p & v9b03cc | !hmaster2_p & v23fd83f;
assign v3763fec = hmaster2_p & v373dd77 | !hmaster2_p & v3731e7b;
assign v3a710e4 = hbusreq2_p & v3a70f74 | !hbusreq2_p & v376bb26;
assign v3727976 = hbusreq3_p & v375bd16 | !hbusreq3_p & !v8455ab;
assign v3740777 = hmaster1_p & v373b5c1 | !hmaster1_p & !v3762145;
assign v3a62c11 = hmaster2_p & v3769ecf | !hmaster2_p & v3771d4f;
assign v3753a3f = hbusreq1 & v3778528 | !hbusreq1 & v3a7162d;
assign v3748a4f = hbusreq6_p & v3a70e86 | !hbusreq6_p & v37571a9;
assign v3a6f810 = hmaster0_p & v8455b0 | !hmaster0_p & v3a5aaf9;
assign v377c8d1 = hmaster2_p & v3a62542 | !hmaster2_p & v3a6fa93;
assign v377b460 = hmaster2_p & v372f309 | !hmaster2_p & v3a6a3e6;
assign v3a56b72 = hbusreq5 & v976f99 | !hbusreq5 & v8455ab;
assign v3756546 = hmaster1_p & v37430c6 | !hmaster1_p & v3a63bd4;
assign v2ff91fe = hbusreq0 & v8cdbc1 | !hbusreq0 & v23fd804;
assign v3a664b8 = hlock0_p & v3776670 | !hlock0_p & v3a70bb2;
assign v3727c62 = hlock4 & v373471f | !hlock4 & v377d10c;
assign v3a5a825 = hmaster1_p & v374beee | !hmaster1_p & v3729830;
assign v3a68c26 = hmaster0_p & v3a702ee | !hmaster0_p & v3a67cf0;
assign v3a61100 = hbusreq8_p & v3a6dea6 | !hbusreq8_p & v3a70e09;
assign v3a6efa4 = hbusreq6_p & v3a6b6dc | !hbusreq6_p & v8455ab;
assign v3a5d448 = hgrant1_p & v8455ab | !hgrant1_p & v3724581;
assign v376e115 = hmaster0_p & v3a70596 | !hmaster0_p & v3a6fd67;
assign v3778333 = hmaster0_p & v373e474 | !hmaster0_p & v3a6497b;
assign v23fdeaf = hbusreq0 & v3a63abb | !hbusreq0 & !v3724a6e;
assign v372c257 = hgrant4_p & v8455ab | !hgrant4_p & v3a70e6b;
assign v376d3e1 = hbusreq4_p & v375ce35 | !hbusreq4_p & v3739cda;
assign v3808e2e = hmaster2_p & v8455ab | !hmaster2_p & v37579ab;
assign v3a6f7fa = hbusreq7_p & v3769199 | !hbusreq7_p & v8455ab;
assign v375a475 = hbusreq7 & v377c22b | !hbusreq7 & v8455ab;
assign v3806e0e = hgrant2_p & v3a2a348 | !hgrant2_p & v3764a16;
assign v3a6fee3 = jx0_p & v3a60628 | !jx0_p & v3779d91;
assign v374a4ea = hbusreq2 & v3a55cd6 | !hbusreq2 & !v8455b5;
assign bf6c15 = hmaster0_p & v8455e7 | !hmaster0_p & v3a6842c;
assign v3a71129 = hbusreq2 & v372ae1b | !hbusreq2 & bf3e2b;
assign v376b082 = hbusreq6 & v3a702bc | !hbusreq6 & v3a6fa2c;
assign v373b317 = hgrant3_p & v8455bd | !hgrant3_p & v373a803;
assign v377d67a = hbusreq2_p & v35b70e6 | !hbusreq2_p & v3761be0;
assign v375e8a2 = hbusreq2 & v3a5e817 | !hbusreq2 & v37c0382;
assign v3a62e1b = hbusreq2_p & v377eaf2 | !hbusreq2_p & v3a7162d;
assign v374fa4f = hbusreq0 & v375d3bc | !hbusreq0 & v8455ab;
assign v3755e4e = hbusreq6_p & v3778b51 | !hbusreq6_p & v35772a6;
assign v3760c32 = hbusreq5_p & v3a603b6 | !hbusreq5_p & !v372f441;
assign v3739e05 = hmaster1_p & a2aef9 | !hmaster1_p & v372e499;
assign v374a6ce = hmaster2_p & v376d268 | !hmaster2_p & v3723a00;
assign v3a6df14 = hmaster2_p & v3a5a807 | !hmaster2_p & v3a71016;
assign v3a6f87e = hmaster0_p & v8455b0 | !hmaster0_p & v372a20b;
assign v37399f7 = hmaster1_p & v3a587d6 | !hmaster1_p & v3769b3f;
assign v376efcf = hlock3 & v38072fd | !hlock3 & v3a6f588;
assign v3a6fbf8 = hbusreq4 & v374db8d | !hbusreq4 & !v8455ab;
assign v3726262 = hmaster2_p & v3a6c20e | !hmaster2_p & v3a6fae9;
assign v3a70c78 = hbusreq7_p & v3a7007c | !hbusreq7_p & v3770ffb;
assign v376218c = hbusreq2_p & v372af46 | !hbusreq2_p & v375f3bd;
assign c3f48e = hmaster2_p & v377adf0 | !hmaster2_p & v37299dd;
assign v3a602cd = hlock5_p & v3a6e8bc | !hlock5_p & !v1e37e4f;
assign v372ca6e = hmaster0_p & v375cec2 | !hmaster0_p & v3a7163a;
assign v3a63039 = hmaster0_p & v373a3b9 | !hmaster0_p & v3a715c5;
assign v3768486 = hbusreq2_p & v375dd60 | !hbusreq2_p & v373c5f5;
assign v373cdbf = hbusreq3_p & v3779060 | !hbusreq3_p & !v3a6dfb2;
assign v23fd8a7 = hbusreq5_p & v3734d60 | !hbusreq5_p & v372e4e1;
assign v3723f33 = hmaster1_p & v376d66b | !hmaster1_p & v35b77ab;
assign v3769945 = hbusreq0 & v3a70848 | !hbusreq0 & v8e4749;
assign v3a67241 = hmastlock_p & v3a70a83 | !hmastlock_p & !v8455ab;
assign v3774a77 = hgrant4_p & v8455ab | !hgrant4_p & v39a4ed6;
assign v373d72e = hgrant6_p & v3733d6e | !hgrant6_p & v377bb21;
assign v373abbe = hbusreq3_p & v3743f94 | !hbusreq3_p & v8455ab;
assign v3a57540 = hlock8_p & v3808db4 | !hlock8_p & v372dbe7;
assign v3a5a01a = hbusreq2 & v3733b37 | !hbusreq2 & v8455e7;
assign v3a660e6 = hbusreq5_p & v37678e2 | !hbusreq5_p & v376e029;
assign v3808d42 = hgrant0_p & v3a653e4 | !hgrant0_p & !v376a21c;
assign v374a277 = hmaster2_p & v3724a4b | !hmaster2_p & v3a6f0f6;
assign v3a6fb95 = hmaster2_p & v3738510 | !hmaster2_p & v3a5cfac;
assign v3a706e4 = hgrant4_p & v3a6eaf3 | !hgrant4_p & v3763aec;
assign v3a65e71 = hmaster2_p & v8455ab | !hmaster2_p & v3a55198;
assign v3749c22 = hgrant1_p & v8455e7 | !hgrant1_p & v3764463;
assign v37635a4 = hbusreq7 & v376ef3d | !hbusreq7 & v3a701cb;
assign v3750fbb = hbusreq4 & v3a61cb2 | !hbusreq4 & v3a6f43a;
assign v3a6b393 = hbusreq6 & v3a65827 | !hbusreq6 & v3a70b92;
assign v3a711ed = hgrant4_p & v8455ab | !hgrant4_p & v3740546;
assign v3a70850 = hbusreq4_p & v3a70373 | !hbusreq4_p & v8455ab;
assign v375685c = hmaster2_p & v37306c2 | !hmaster2_p & v3766ce0;
assign v3728464 = hmaster1_p & v3727bc6 | !hmaster1_p & v3736ded;
assign v375c48c = hmaster0_p & v3a710bd | !hmaster0_p & v88d9b8;
assign v3a5cd5c = hbusreq0 & v37543a0 | !hbusreq0 & v373d9d3;
assign v3766232 = hbusreq7 & v3a70739 | !hbusreq7 & v373a005;
assign v3a7044d = hlock0_p & v2ff9190 | !hlock0_p & v8455ab;
assign v3735c5d = hgrant3_p & v35b7299 | !hgrant3_p & !v1e37a69;
assign v373fa89 = hgrant4_p & v375e752 | !hgrant4_p & v376acee;
assign v3a7156d = hbusreq3_p & v8455e7 | !hbusreq3_p & v374f307;
assign v3a53b85 = hmaster2_p & v9bf1d8 | !hmaster2_p & v374eedb;
assign v372aed1 = hgrant4_p & v3768857 | !hgrant4_p & v3a7163e;
assign v376c477 = hmaster1_p & v8455ab | !hmaster1_p & v37231c2;
assign v37259bc = hlock2 & v3722e4c | !hlock2 & v3a6741a;
assign v3a710f0 = hmaster2_p & v3a5fc34 | !hmaster2_p & v3a6f42e;
assign v3a6a609 = hbusreq3_p & v3a59f74 | !hbusreq3_p & v372e59e;
assign v3763387 = hgrant8_p & v3a6443f | !hgrant8_p & v376634b;
assign v3a706da = hmaster0_p & v8455ab | !hmaster0_p & v374c88d;
assign v3a6603f = hgrant4_p & v8455ab | !hgrant4_p & v3a71247;
assign v3774b71 = hmaster1_p & v3a6f3ae | !hmaster1_p & !v3779613;
assign v37560b0 = hbusreq5_p & v3a60f9b | !hbusreq5_p & v8455ab;
assign v3a66667 = hmaster0_p & v3728d9c | !hmaster0_p & v37504fd;
assign v37571f1 = hbusreq6 & v375185f | !hbusreq6 & v3a5edcb;
assign v374efb3 = hlock5_p & v377be84 | !hlock5_p & v373520f;
assign v376ff89 = hgrant6_p & v3771b2c | !hgrant6_p & v373d3dd;
assign v3765626 = hbusreq2_p & v3a700ad | !hbusreq2_p & v3a713e3;
assign v376a3ca = hbusreq6_p & v3757ec8 | !hbusreq6_p & v3a6b405;
assign v3a70c61 = hgrant1_p & v8455b7 | !hgrant1_p & v3a70293;
assign v377cc72 = hbusreq7_p & v37547f7 | !hbusreq7_p & v8455ab;
assign v3761ad8 = hbusreq3_p & v3729e65 | !hbusreq3_p & !v35772a6;
assign v3769069 = hbusreq5 & v376ed63 | !hbusreq5 & v377de7f;
assign v3a6efdf = jx0_p & v3a6eb7f | !jx0_p & v3752535;
assign v376848c = hbusreq7 & v372bb82 | !hbusreq7 & v372bf1d;
assign v377ab2c = hgrant3_p & v375c1d1 | !hgrant3_p & v8455ab;
assign v3a6fedc = hgrant6_p & v3a5cfac | !hgrant6_p & v374b429;
assign v3a59e5e = hbusreq4 & v37639c3 | !hbusreq4 & v8455ab;
assign v375e5a6 = hmaster1_p & v3733168 | !hmaster1_p & !v8455ab;
assign v37300b7 = hgrant3_p & v3a6251b | !hgrant3_p & v374a891;
assign v3753fe0 = hgrant0_p & v37773a9 | !hgrant0_p & v376e611;
assign v375c90b = hbusreq6_p & v3a6a1fd | !hbusreq6_p & v373c95b;
assign v3771319 = hmaster1_p & v376f9be | !hmaster1_p & v37258e7;
assign v97ecca = hlock0_p & v377eaf2 | !hlock0_p & v3a70bd2;
assign v374b160 = hmaster2_p & v3a716a0 | !hmaster2_p & v3a7153c;
assign v3729180 = hmaster1_p & a94d63 | !hmaster1_p & v8455ab;
assign v3a69043 = hlock3 & v375b7dc | !hlock3 & v3a70a45;
assign v3a6fba1 = hlock6 & v3a6767d | !hlock6 & v376c351;
assign v372fba0 = hmaster2_p & v3737d02 | !hmaster2_p & v374e64f;
assign v864fe4 = hbusreq5_p & v3765f99 | !hbusreq5_p & v3a709fc;
assign v3a70a6f = hbusreq3 & v376a14f | !hbusreq3 & v8455ab;
assign v374503d = hbusreq0 & v3a56494 | !hbusreq0 & v373bd6c;
assign v3734c47 = hbusreq5 & v374f077 | !hbusreq5 & v374c6b8;
assign v3a6f24c = hlock4_p & v3a5d08a | !hlock4_p & v3a6ef6d;
assign v37669b4 = hbusreq3_p & v375928d | !hbusreq3_p & v3725994;
assign v3a6f37f = hbusreq2_p & v3a554b9 | !hbusreq2_p & !v3a68591;
assign v377cd5b = hbusreq6 & v37484df | !hbusreq6 & v372914b;
assign v3a6fce0 = hmaster0_p & v3a6f591 | !hmaster0_p & v3a6f4f5;
assign v3729823 = hgrant0_p & v8455ab | !hgrant0_p & v3a7168a;
assign v3735bf3 = hbusreq7_p & v373a0f4 | !hbusreq7_p & v8455ab;
assign v3763d52 = hbusreq0 & v3a5a0e2 | !hbusreq0 & v3a67519;
assign v3a6f483 = hgrant0_p & v8455ab | !hgrant0_p & v3744b38;
assign v3809865 = hbusreq3 & v3750e9a | !hbusreq3 & v377ad8f;
assign v3735a94 = hmaster2_p & v8455ab | !hmaster2_p & !v3770ccf;
assign v376fb37 = hgrant5_p & v8455ab | !hgrant5_p & v23fde6d;
assign v37615c5 = hbusreq4_p & v3759886 | !hbusreq4_p & !v8455c2;
assign v373b36c = hgrant6_p & v377f21b | !hgrant6_p & v377657c;
assign v373f364 = hbusreq8_p & v376209f | !hbusreq8_p & v3a5d6b7;
assign v3a5e070 = hgrant4_p & v3a656d0 | !hgrant4_p & v3751338;
assign v376064b = hbusreq2_p & v337901e | !hbusreq2_p & v8455ab;
assign v375ff11 = hbusreq5_p & v3a6f7d0 | !hbusreq5_p & v3758f89;
assign v377e056 = hmaster0_p & v37774ca | !hmaster0_p & v37458ca;
assign v3a71461 = jx1_p & v3764f01 | !jx1_p & v37274a1;
assign v3a65402 = hmaster0_p & v3a6f84a | !hmaster0_p & v3a6ebac;
assign v3809464 = hmaster1_p & v374f432 | !hmaster1_p & v3773d96;
assign v375178a = hbusreq8_p & v373635b | !hbusreq8_p & v3a70e53;
assign v3a68525 = hmaster0_p & v37763d1 | !hmaster0_p & v372cde4;
assign v3750735 = hbusreq5_p & v375c6c1 | !hbusreq5_p & v377b429;
assign v373e12e = hbusreq3_p & v373588a | !hbusreq3_p & !v3a6ff7d;
assign v373dad7 = hmaster2_p & v8455e1 | !hmaster2_p & !v3738877;
assign v3a7113c = hmaster2_p & v8455ab | !hmaster2_p & v372414d;
assign v3761181 = hbusreq3 & v35772c9 | !hbusreq3 & v8455ab;
assign v3a6fb8a = hgrant5_p & v3808d74 | !hgrant5_p & v3808cbf;
assign v3739ed3 = hmaster1_p & v8455ab | !hmaster1_p & v372ed93;
assign v374c5c6 = hmaster2_p & v37640e9 | !hmaster2_p & v374d4e6;
assign v39a4f09 = hlock4_p & v37624a2 | !hlock4_p & v8455b0;
assign v3a6802b = hgrant2_p & v375c55a | !hgrant2_p & v37299e2;
assign v37786f9 = hmaster1_p & v377a3bd | !hmaster1_p & v3778419;
assign v372c0cc = hbusreq5_p & v3a68dcb | !hbusreq5_p & v8455ab;
assign v3731725 = hlock5 & v37251c9 | !hlock5 & v3732f19;
assign v377e1d0 = hbusreq6_p & v3a6f696 | !hbusreq6_p & v37603b3;
assign v3a71020 = hmaster1_p & v38094ca | !hmaster1_p & v3768774;
assign v3762158 = hmaster2_p & v8455ab | !hmaster2_p & v3a5915c;
assign v3758892 = hlock7 & v3772e44 | !hlock7 & v37690e7;
assign v372cdf6 = hbusreq4 & v37348ee | !hbusreq4 & v3a69487;
assign v3a6f814 = hlock1_p & v1e38275 | !hlock1_p & v39a537f;
assign hgrant4 = !v39e9ca4;
assign v3742ce8 = hbusreq2 & v3a6dc08 | !hbusreq2 & v8455b0;
assign v377de6f = hmaster2_p & v375a268 | !hmaster2_p & !v376e914;
assign v3a6f11e = hbusreq5 & v376e9fd | !hbusreq5 & v3a70894;
assign v3776691 = hbusreq7_p & a0a219 | !hbusreq7_p & v374373c;
assign v37522ff = hlock4 & v373e450 | !hlock4 & v3809e93;
assign v372a704 = hmaster1_p & v3736d47 | !hmaster1_p & v374d86e;
assign v376a59f = hbusreq7_p & a0a219 | !hbusreq7_p & v373a7dc;
assign v37574d2 = hlock2 & v374d480 | !hlock2 & v3751dc9;
assign v372aa71 = hmaster0_p & v373dd7f | !hmaster0_p & v374f397;
assign v3a6c001 = hmaster2_p & v372fc81 | !hmaster2_p & !v3a696ed;
assign v3a703b8 = hmaster3_p & v377435d | !hmaster3_p & v3a59b42;
assign v3a54dd4 = hmaster0_p & v3a7066c | !hmaster0_p & v3a71340;
assign v3732949 = hlock2_p & v37463bc | !hlock2_p & !v8455ab;
assign v37716e1 = hlock8 & v3a59d6b | !hlock8 & v3725e9a;
assign v3a6fdb3 = hbusreq5_p & v376fe45 | !hbusreq5_p & v3767080;
assign v373197e = hbusreq3_p & v376dbdf | !hbusreq3_p & !v372fc81;
assign v374a2f3 = hbusreq0 & v8455b3 | !hbusreq0 & v373e814;
assign v37702e0 = hgrant5_p & v377c8ca | !hgrant5_p & v3a6c0c1;
assign hgrant7 = !v39a4f35;
assign v3723b00 = hbusreq1_p & v8455e7 | !hbusreq1_p & v374f307;
assign v3a63f6d = hlock7_p & v3735ae4 | !hlock7_p & !v8455ab;
assign v37600af = hlock0_p & v3a660f2 | !hlock0_p & v3a6fa39;
assign v3757598 = hgrant3_p & v3a7000e | !hgrant3_p & v8455ab;
assign v3a611b0 = hbusreq0 & v377dfec | !hbusreq0 & !v8455ab;
assign v3771dda = hbusreq0 & v3a612a3 | !hbusreq0 & v3777642;
assign v37682dd = hmaster1_p & v374502e | !hmaster1_p & v374ca8a;
assign v3a55861 = hmaster1_p & v8455ab | !hmaster1_p & v3a6f66a;
assign v37297f9 = hbusreq7 & v3a6eedf | !hbusreq7 & a0a219;
assign v37760b8 = jx0_p & v37414cd | !jx0_p & v376930a;
assign v3a6fc93 = hbusreq7_p & v3740a1e | !hbusreq7_p & v3a6fe81;
assign v373ce36 = hmaster1_p & v37485cb | !hmaster1_p & v375ed37;
assign v373d67c = hmaster2_p & v126f91f | !hmaster2_p & v8455ab;
assign v3728fd2 = hbusreq5 & v377ad63 | !hbusreq5 & v3772231;
assign v3727af8 = hmaster2_p & v37566b2 | !hmaster2_p & v39a537f;
assign v3a5bf4c = hmaster0_p & v380a1f3 | !hmaster0_p & v37686ea;
assign v376d312 = hmaster2_p & v3770754 | !hmaster2_p & v3a5d36a;
assign v3a6a4e6 = hmaster2_p & v3a703fc | !hmaster2_p & !v8455ab;
assign v3738cfc = start_p & v3776483 | !start_p & v3a7111f;
assign v3a70650 = hmaster0_p & v3738b0b | !hmaster0_p & v37585d8;
assign v373373d = hmaster0_p & v8455bf | !hmaster0_p & v37374a1;
assign v3a6f958 = hburst1 & v3a70cd5 | !hburst1 & v376b4d7;
assign v3751968 = hbusreq4_p & v3a70ca3 | !hbusreq4_p & !v3748a87;
assign v3a6210a = hbusreq4 & v37697ba | !hbusreq4 & v373d4ff;
assign v3a6fed7 = hmaster0_p & v3750a45 | !hmaster0_p & v376db34;
assign v37470c7 = hgrant4_p & v377aa81 | !hgrant4_p & v2925ca9;
assign v373918a = hgrant1_p & v3807bf8 | !hgrant1_p & v372c11d;
assign v3724596 = hmaster2_p & v3774647 | !hmaster2_p & v373b779;
assign v376ab72 = hlock3 & v3769616 | !hlock3 & v374ace7;
assign v3a700e2 = hgrant4_p & v8455b0 | !hgrant4_p & v3722e7a;
assign v3757c91 = hbusreq2_p & v37749bf | !hbusreq2_p & v3a70b6e;
assign v37353b5 = hlock6_p & v373f63e | !hlock6_p & v3a6dfc6;
assign v373aea0 = hbusreq3 & v372c3df | !hbusreq3 & !v3a69515;
assign v37570eb = hbusreq5_p & v3760bfa | !hbusreq5_p & v3753994;
assign v3a6ee64 = hmaster2_p & v3729a2a | !hmaster2_p & v377960b;
assign v3739120 = hlock5_p & v3778372 | !hlock5_p & v35772a6;
assign v3a6f97d = hbusreq4 & v3739aa6 | !hbusreq4 & v8455ab;
assign v3a707ef = hmaster1_p & v8455ab | !hmaster1_p & v3745717;
assign v23fdac1 = hmaster0_p & v37719a1 | !hmaster0_p & v37382eb;
assign v376bbcc = hmaster2_p & v8455ab | !hmaster2_p & v372342b;
assign v3a6ec76 = hbusreq4 & v375153e | !hbusreq4 & v3777460;
assign v3756206 = hbusreq2 & v3a617b4 | !hbusreq2 & v3773ee6;
assign v3a5f622 = hmaster1_p & v377766c | !hmaster1_p & v376a915;
assign v375aff8 = hmaster0_p & v37666f6 | !hmaster0_p & v3a6d531;
assign v3759623 = hgrant2_p & v37321b8 | !hgrant2_p & v374189b;
assign v3a5e6f6 = hbusreq2_p & v37765e1 | !hbusreq2_p & v374b4a4;
assign v37391e8 = hgrant6_p & v377b6ce | !hgrant6_p & v372fd45;
assign v376db9c = hmaster2_p & v3769be7 | !hmaster2_p & v377ef4a;
assign v35b77ec = hmaster2_p & v3766a8d | !hmaster2_p & v375bb92;
assign v3755691 = hmaster0_p & v3767d57 | !hmaster0_p & v8455ab;
assign v3a70e77 = hlock4 & v377e85a | !hlock4 & v3a53d12;
assign v372eafa = hbusreq4 & v3740171 | !hbusreq4 & v8455e7;
assign v3779069 = hmaster2_p & v374314f | !hmaster2_p & v3758133;
assign v3755b54 = hgrant3_p & v3a710e9 | !hgrant3_p & v3a70d90;
assign v3a5f20d = hgrant6_p & v3a702bb | !hgrant6_p & v3a5a52a;
assign b79c3c = hmaster1_p & v8455ab | !hmaster1_p & v3a7097f;
assign v3766a37 = hbusreq7 & v3a5f447 | !hbusreq7 & v3a6ef56;
assign v37651b4 = hgrant4_p & v3a53eeb | !hgrant4_p & v37659f8;
assign v37499a9 = hmaster0_p & v3a6efe8 | !hmaster0_p & v375dd80;
assign v3752f78 = stateA1_p & v8455ab | !stateA1_p & v3777ff3;
assign v3a58b1f = hbusreq4_p & v337900b | !hbusreq4_p & v37451ad;
assign v3a296dc = hbusreq4_p & v372fd0a | !hbusreq4_p & !v8455ab;
assign v3749e5a = hgrant6_p & v3a62b8d | !hgrant6_p & v3a6eb94;
assign v3723a2c = hbusreq8 & v376aa62 | !hbusreq8 & v373c433;
assign v37721df = hlock4_p & v3379037 | !hlock4_p & !v8455ab;
assign v377e5e1 = hmaster0_p & v2092b0b | !hmaster0_p & !v8455ab;
assign v3752fb7 = hbusreq2 & v3a603bb | !hbusreq2 & v376e041;
assign v37496fa = locked_p & v8455ab | !locked_p & v3a635ea;
assign v372b59d = hbusreq6 & v3723b00 | !hbusreq6 & v8455ab;
assign v373357d = hmaster1_p & v377ea20 | !hmaster1_p & v37627ec;
assign d90332 = hbusreq0 & v3a67f60 | !hbusreq0 & v3733f28;
assign v375b713 = hbusreq2_p & v3a70e65 | !hbusreq2_p & v3a6fcef;
assign v3809e90 = hbusreq5_p & v373ed5c | !hbusreq5_p & v3a661c2;
assign v3752a45 = hlock1_p & v37686af | !hlock1_p & v37547c9;
assign v37608ba = hmaster2_p & v377eb2d | !hmaster2_p & v8455ab;
assign v3a70bf5 = hbusreq6_p & v3a53c9d | !hbusreq6_p & v3a708f0;
assign v3a6fefc = hlock4 & v3726054 | !hlock4 & v3a70f3d;
assign v3a5b855 = hbusreq0 & v3769cd3 | !hbusreq0 & v8455ab;
assign d2dc90 = hbusreq0 & v3a6fabe | !hbusreq0 & v1e37cd6;
assign v374e4fa = hmaster0_p & v374d43f | !hmaster0_p & v376132a;
assign v3733d60 = hmaster0_p & v3a7071a | !hmaster0_p & v88d9b8;
assign v3738f5a = hbusreq6 & v3750dd3 | !hbusreq6 & v8455bb;
assign v375ff00 = hmaster0_p & v37349cc | !hmaster0_p & v372acd0;
assign v3a62ad5 = hbusreq0 & v3748cce | !hbusreq0 & v8455ab;
assign v374b690 = hgrant3_p & v8455ab | !hgrant3_p & v3a70e9f;
assign v3a55b61 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a70a7f;
assign v3759d52 = hbusreq6_p & v37439c2 | !hbusreq6_p & v8455ab;
assign v3763004 = hgrant2_p & v374ca41 | !hgrant2_p & cd3a92;
assign v3a6efc9 = hmastlock_p & v3745b52 | !hmastlock_p & v8455ab;
assign v3758f89 = hbusreq5 & v376ee43 | !hbusreq5 & v3a71506;
assign v3a711de = hlock4 & v3a6fba9 | !hlock4 & v3a6eb1e;
assign v3a713bf = hmaster1_p & v3a564d9 | !hmaster1_p & v3a70217;
assign v3750012 = hready_p & v3a6f337 | !hready_p & c8f3d0;
assign v37494da = hbusreq7_p & v3a704a7 | !hbusreq7_p & v3a575a5;
assign v376ac56 = hmaster0_p & v3a661fe | !hmaster0_p & v3a711db;
assign v37718cc = hgrant4_p & v8455ab | !hgrant4_p & !v3a6d0ec;
assign v3730755 = hbusreq6_p & v39a537f | !hbusreq6_p & !v39a5381;
assign v377c2d9 = hmaster2_p & v3a70c3e | !hmaster2_p & v3a7119c;
assign v374caf9 = hlock5 & v375970d | !hlock5 & v376256c;
assign v3a5f60f = hmaster3_p & v372d1b1 | !hmaster3_p & v3a71398;
assign v374216a = hmaster2_p & v3a6cc65 | !hmaster2_p & v8455ab;
assign v3754c86 = hlock6_p & v373a841 | !hlock6_p & v3765e46;
assign v375fed2 = stateA1_p & v3a5b585 | !stateA1_p & v3a6f682;
assign v3a7024a = hmaster1_p & v3775303 | !hmaster1_p & v37651cc;
assign v3733a5f = hbusreq0 & v376c1e4 | !hbusreq0 & v3729280;
assign v3a58b4c = hlock6_p & v3a687be | !hlock6_p & v373f058;
assign v3806b78 = hbusreq4_p & v37656b8 | !hbusreq4_p & v37643e5;
assign v3a6fef2 = hmaster1_p & v3a6fc5e | !hmaster1_p & v3768196;
assign v377a3af = hmaster1_p & v3a70c92 | !hmaster1_p & v8455ab;
assign v37289bc = hmaster1_p & v373013d | !hmaster1_p & v377eb8b;
assign v3a6f884 = hbusreq3_p & v374b0a8 | !hbusreq3_p & v3a5cd20;
assign v37429a7 = hmaster1_p & v3a6fc19 | !hmaster1_p & v3779678;
assign v376d550 = hmaster2_p & v374c7f4 | !hmaster2_p & v3a627cc;
assign v37370f0 = hmaster2_p & v3a70ff5 | !hmaster2_p & v3a6a8ee;
assign v3735ad7 = hbusreq8 & v3731974 | !hbusreq8 & v8455ab;
assign v89fdcf = hbusreq5 & v374db73 | !hbusreq5 & v377234d;
assign v3a70675 = hmaster0_p & v373abc5 | !hmaster0_p & v3728fda;
assign v3a5509a = hmaster1_p & v377bb3a | !hmaster1_p & v8ebe6e;
assign v3a6ff85 = hlock6_p & v3746063 | !hlock6_p & v8455b0;
assign v3726ae2 = hbusreq0 & v3a70006 | !hbusreq0 & v1e37cd6;
assign v376693b = hbusreq2_p & bf3e2b | !hbusreq2_p & v373fbc7;
assign v3a6826a = hmaster0_p & v377b2e1 | !hmaster0_p & v3764a7d;
assign v3a5c1a1 = hbusreq7_p & v8fa780 | !hbusreq7_p & !v374d7fc;
assign v3a5ba93 = hmaster0_p & v3a635ea | !hmaster0_p & v377d839;
assign v3a689bb = hmaster2_p & v3a635ea | !hmaster2_p & v374f35a;
assign v3a6d2eb = hmaster1_p & v372da2f | !hmaster1_p & v3a6db03;
assign v3770c1a = hmaster0_p & v3a5e665 | !hmaster0_p & v3754727;
assign v3740ee1 = hgrant0_p & v372beb8 | !hgrant0_p & v3a68426;
assign v372e2cd = hmaster0_p & v377accc | !hmaster0_p & v3762997;
assign v3744d36 = hbusreq6 & v3a702b5 | !hbusreq6 & v3a635ea;
assign v375654b = hlock8_p & v37261b2 | !hlock8_p & v8455cb;
assign v375986d = hgrant5_p & v3a6924e | !hgrant5_p & v3a600a8;
assign v373ce84 = hbusreq6 & v37436a8 | !hbusreq6 & v3a7011e;
assign v37412f3 = hmaster2_p & v3a707b7 | !hmaster2_p & v372a00b;
assign v3771e18 = hlock3_p & v377bb86 | !hlock3_p & v377a4f1;
assign v372d8c9 = hgrant6_p & v3a71164 | !hgrant6_p & v3a6f547;
assign v373b5f5 = hlock2_p & v372af30 | !hlock2_p & !v8455ba;
assign v37707d5 = hgrant6_p & v37728a5 | !hgrant6_p & v3a70988;
assign v3752cf6 = hgrant6_p & v3a6c5ee | !hgrant6_p & v373fc8a;
assign v3769a1e = hgrant6_p & v8455ab | !hgrant6_p & v3742aae;
assign v3778aa0 = hmaster0_p & v3a5b8b9 | !hmaster0_p & v3a64fb4;
assign v372aeef = jx1_p & v3747db9 | !jx1_p & v3a6c73d;
assign v3a56929 = hbusreq8 & v374294f | !hbusreq8 & v3a62ba4;
assign v3a6f056 = hburst1_p & v3a7111f | !hburst1_p & !v8455ab;
assign v3a6f03d = hmaster0_p & v377574b | !hmaster0_p & v376d1cb;
assign v3a67d66 = hbusreq2_p & v3764c4c | !hbusreq2_p & v8455ab;
assign v376eaed = hgrant5_p & v373c1ed | !hgrant5_p & v3a62ee2;
assign v3a70089 = hmaster1_p & v8455ab | !hmaster1_p & v37264a2;
assign v376acd9 = hmaster0_p & v3a6fe31 | !hmaster0_p & !v3726434;
assign v376b1bf = hgrant2_p & v3a632f4 | !hgrant2_p & v375b269;
assign v866387 = hmaster3_p & v37361ad | !hmaster3_p & v8455d1;
assign v372e889 = hmaster2_p & v3730b98 | !hmaster2_p & v3a7089d;
assign v3750c52 = hgrant6_p & v3a62a6d | !hgrant6_p & v3a708f0;
assign v376dc21 = hgrant1_p & v37416b5 | !hgrant1_p & v376d327;
assign v372ad29 = hmaster3_p & v39eb418 | !hmaster3_p & v372e3db;
assign v3a6b6dc = hlock6_p & v3775b81 | !hlock6_p & v8455ab;
assign v3723af9 = hgrant2_p & v376b087 | !hgrant2_p & v3736785;
assign v3a57887 = jx3_p & v377d6c5 | !jx3_p & v373cb13;
assign b30936 = hlock7 & v3a705aa | !hlock7 & v373f2d2;
assign v3a6ebed = hbusreq4_p & v377a99d | !hbusreq4_p & v374bbcc;
assign v377e896 = hgrant7_p & v8455ab | !hgrant7_p & v3a6f626;
assign v37706fd = hbusreq4 & ade0d8 | !hbusreq4 & v377b2d0;
assign v375f2e8 = hmaster1_p & v375d364 | !hmaster1_p & v376314e;
assign v28896da = hbusreq2_p & v3a6d642 | !hbusreq2_p & v8455ab;
assign v376c1cc = hbusreq3_p & v37741bc | !hbusreq3_p & v3a6f7f9;
assign v37759ff = hmaster2_p & v3a5fe3c | !hmaster2_p & v3a70ecb;
assign v3a54059 = hbusreq8 & v37500db | !hbusreq8 & v3a6194e;
assign v37266d1 = hmaster0_p & v3a6efe8 | !hmaster0_p & v377041c;
assign v3769f2f = hgrant2_p & v3a6f02f | !hgrant2_p & v3a6ef6e;
assign v3a6bff5 = hbusreq5 & v377997f | !hbusreq5 & v3a6fe59;
assign v3756c5d = hgrant4_p & v373ee17 | !hgrant4_p & v3773bb0;
assign v374ca4a = hlock0 & v376bade | !hlock0 & v3a54dfa;
assign v373e91a = hbusreq5_p & v3769ae2 | !hbusreq5_p & v376999f;
assign v3a5bb85 = hmaster0_p & v3a6aaea | !hmaster0_p & v3742abe;
assign v3762f27 = hmaster0_p & v3a5fe00 | !hmaster0_p & v3a6f291;
assign v3730b3a = hbusreq8_p & v3759569 | !hbusreq8_p & v3a65130;
assign v37700ee = hbusreq0_p & v8455ab | !hbusreq0_p & v3a6a939;
assign v3745a3b = hmaster0_p & v3a58cfc | !hmaster0_p & v372d149;
assign v372b006 = hbusreq5_p & v374b497 | !hbusreq5_p & v373c58c;
assign a9ca33 = hmaster0_p & v37320bf | !hmaster0_p & v376669c;
assign v3a61c73 = hlock7 & v94335e | !hlock7 & v3a5d25d;
assign v3725556 = hbusreq2_p & v3a635ea | !hbusreq2_p & v372e132;
assign v3a6f1a6 = hmaster0_p & v3772962 | !hmaster0_p & v3723be4;
assign v3a58d63 = hbusreq0 & v3724c35 | !hbusreq0 & v3a6b8d8;
assign v37245d9 = hbusreq1_p & v3a5ce2f | !hbusreq1_p & !v375d651;
assign v3a6e127 = hmaster0_p & v3a6fe0d | !hmaster0_p & v3756de7;
assign v37229ba = hmaster0_p & v3a54aa0 | !hmaster0_p & v3a710f7;
assign v372554a = hbusreq2 & v8455b0 | !hbusreq2 & adf78a;
assign v373a41e = hbusreq7_p & v3a6f680 | !hbusreq7_p & v3a5f5dd;
assign v374eb6a = hbusreq6 & d44200 | !hbusreq6 & v374e35e;
assign v374916a = hgrant4_p & v3a61acf | !hgrant4_p & v3a6fb86;
assign v374b03c = hmaster2_p & v37416c6 | !hmaster2_p & v374693f;
assign v3a702b4 = hbusreq2_p & v3761c68 | !hbusreq2_p & v3a710b7;
assign v377de0d = hbusreq2 & v3a67904 | !hbusreq2 & v8455ab;
assign v3a7042c = hgrant5_p & v8455ab | !hgrant5_p & v374f31c;
assign v3770b26 = hgrant4_p & v8455ab | !hgrant4_p & v372c84a;
assign v3a6219d = hbusreq2 & v372d203 | !hbusreq2 & v376de4e;
assign v3a6f931 = hbusreq7_p & v376e160 | !hbusreq7_p & v3a5dc5c;
assign v374551a = hbusreq3_p & v37bfcae | !hbusreq3_p & v3756bc2;
assign v375d20f = hbusreq7_p & v373d09a | !hbusreq7_p & !v3748984;
assign v9015e2 = hlock6_p & v2ff9190 | !hlock6_p & v8455ab;
assign v3761954 = hmaster0_p & v3a5a6e6 | !hmaster0_p & v3a6f4f0;
assign v3a709f1 = hmaster1_p & v3a63bde | !hmaster1_p & v37330ca;
assign v3768202 = hlock0_p & v373ad95 | !hlock0_p & v8455ab;
assign v3744dda = hmaster3_p & v3737808 | !hmaster3_p & v8455ab;
assign v3761587 = hgrant6_p & v8455ab | !hgrant6_p & v3a6fa36;
assign v3a603e0 = hlock3 & v3748797 | !hlock3 & v3a61668;
assign v3760101 = hbusreq3 & v3a693af | !hbusreq3 & v8455ab;
assign v3722b6f = jx0_p & v374e5e9 | !jx0_p & v3736af1;
assign v3a5cf0b = start_p & v3730a0f | !start_p & v3730383;
assign v377437f = hgrant3_p & v3a70710 | !hgrant3_p & v373b2ce;
assign v375a5e3 = hmaster0_p & v372ff6d | !hmaster0_p & v37691e2;
assign v3a60628 = hbusreq7_p & v3734279 | !hbusreq7_p & v377ece3;
assign v377f01a = hbusreq3 & v3806db7 | !hbusreq3 & v8455ab;
assign v373977e = jx1_p & v376fddd | !jx1_p & v377f7dd;
assign v3a29da0 = hmaster2_p & v3746d2a | !hmaster2_p & v376a056;
assign v3731312 = hmaster1_p & v3754e8e | !hmaster1_p & v3a70f68;
assign v3768538 = hgrant6_p & v8455ab | !hgrant6_p & v375add8;
assign v373d78b = hlock0_p & v3a70641 | !hlock0_p & v3742259;
assign v3a6eb28 = hmaster1_p & v3744c88 | !hmaster1_p & v376b87b;
assign v375be64 = hbusreq3 & v3a5f265 | !hbusreq3 & v3a59d9d;
assign v3757f01 = hbusreq0 & v3a6f70c | !hbusreq0 & v8455ab;
assign v3a6731d = hbusreq8_p & v372dc77 | !hbusreq8_p & v3a6fc76;
assign v3778430 = hlock4 & v3767892 | !hlock4 & v3a54919;
assign v3a70766 = hbusreq8_p & v3a5c1a1 | !hbusreq8_p & v8455ab;
assign v3a6fe6c = hmaster2_p & v8455ab | !hmaster2_p & v3747c3e;
assign v1e37ebb = hbusreq4_p & v3a6f801 | !hbusreq4_p & v3750c52;
assign v3769245 = hlock5_p & v372771e | !hlock5_p & v3a67f0c;
assign v3a576c0 = hmaster2_p & v8455ab | !hmaster2_p & !v37681fa;
assign v3771c38 = hbusreq5 & b8f5a8 | !hbusreq5 & v3a6d4f3;
assign v372b5a8 = hbusreq2_p & v3a70799 | !hbusreq2_p & v37400bc;
assign v3a7159c = hgrant6_p & v3a64045 | !hgrant6_p & v3a652a6;
assign v376e854 = hbusreq0 & v376b21a | !hbusreq0 & v8455ab;
assign v3a544de = hlock6_p & v8455ab | !hlock6_p & v360d080;
assign v3744657 = hgrant5_p & v3a6f851 | !hgrant5_p & v372ce4a;
assign v376c22c = hmaster2_p & v8455ab | !hmaster2_p & v373c665;
assign v3a6f850 = jx0_p & v37512d2 | !jx0_p & v3a7046f;
assign v3a70989 = hbusreq8_p & v3728fee | !hbusreq8_p & v3a6877a;
assign v375ab92 = hgrant5_p & v37621c1 | !hgrant5_p & v3728a6d;
assign v3770edc = hmaster1_p & v374decf | !hmaster1_p & v3735d84;
assign v3a6fac3 = hbusreq5_p & v3a70b9f | !hbusreq5_p & !v8455ab;
assign v3761ff9 = hmaster1_p & v8455ab | !hmaster1_p & v3760646;
assign v374d163 = hmaster1_p & v3731839 | !hmaster1_p & v8455ab;
assign v3a63dba = hbusreq5_p & v3779bde | !hbusreq5_p & v3a61d1f;
assign d38ecb = hlock5 & v3a6c905 | !hlock5 & v3a66c9a;
assign v373f461 = hmaster1_p & v3729263 | !hmaster1_p & v3a5e7f7;
assign v373287a = hgrant5_p & v8455ab | !hgrant5_p & v3730a7b;
assign v377b73b = hlock8 & v3a5f358 | !hlock8 & v37529d6;
assign v3a64355 = hmaster0_p & v3a6fd02 | !hmaster0_p & v3a68426;
assign v376462a = hbusreq4_p & v3740df7 | !hbusreq4_p & v3759158;
assign v3738679 = hbusreq4 & v3a6f3da | !hbusreq4 & v3a70b92;
assign v8bc7a8 = hmaster2_p & v8455ab | !hmaster2_p & v3754450;
assign v3a70fde = hbusreq8_p & v3a68e0d | !hbusreq8_p & v376e66e;
assign v35b724a = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3778528;
assign v374c062 = hgrant1_p & v3a6f10f | !hgrant1_p & v377989c;
assign v3768933 = hbusreq3_p & v3766996 | !hbusreq3_p & v8455ab;
assign v3777deb = hbusreq6_p & c29340 | !hbusreq6_p & v372cc25;
assign v372672f = hbusreq6_p & v374a3c5 | !hbusreq6_p & v8455b0;
assign v376c176 = hbusreq6_p & v373fe5e | !hbusreq6_p & v8455e7;
assign v37729e0 = hmaster2_p & v3a635ea | !hmaster2_p & v3765e79;
assign v377d9aa = hbusreq4 & v374cab9 | !hbusreq4 & !v8455ab;
assign v375b5d3 = hmaster2_p & v374306c | !hmaster2_p & v35772a6;
assign v372aacd = hlock0_p & v8455ab | !hlock0_p & v3775107;
assign v377027e = hmaster2_p & v39a5381 | !hmaster2_p & !v3751734;
assign v372d4de = hbusreq6 & v3a6f20d | !hbusreq6 & v376e041;
assign v375edd8 = jx0_p & v37523b5 | !jx0_p & v3779c8d;
assign v3a70486 = hbusreq3 & v3723247 | !hbusreq3 & v376c343;
assign v376aaf5 = hlock8 & v37465d4 | !hlock8 & v37586d1;
assign v372c6c4 = hlock5_p & v8455e7 | !hlock5_p & !v8455ab;
assign v3a70a50 = hlock2 & v3806a6f | !hlock2 & v37645a8;
assign v374ae3d = hbusreq3 & v37718fb | !hbusreq3 & v8455ab;
assign v3a715ce = hbusreq8 & v3a70426 | !hbusreq8 & v3768734;
assign v3a7133f = hbusreq2_p & v3a65a33 | !hbusreq2_p & v2619ac3;
assign v3731381 = hmaster0_p & v37770f5 | !hmaster0_p & v3a71614;
assign v3a5f5dd = hgrant5_p & v3a661f8 | !hgrant5_p & v3a70695;
assign v3a5c58f = hbusreq4_p & v3748797 | !hbusreq4_p & v3a6d6be;
assign v3a6f873 = hgrant5_p & v376e240 | !hgrant5_p & v9aa32c;
assign v3767919 = hmaster1_p & v3728916 | !hmaster1_p & v37424a9;
assign v3757ecc = hgrant6_p & v377e13b | !hgrant6_p & !v37474c2;
assign v3809752 = hbusreq6_p & v3748797 | !hbusreq6_p & v374ed0a;
assign v375f823 = hgrant4_p & v3a71025 | !hgrant4_p & v3746202;
assign v3a6fca0 = hbusreq8_p & v3765d05 | !hbusreq8_p & !v8455ab;
assign v3a6fa69 = hmaster2_p & v37267d6 | !hmaster2_p & v3a65762;
assign v3a606e8 = hgrant3_p & v8455ab | !hgrant3_p & !v2ff9287;
assign v3a6f5a1 = hbusreq0 & v377d2bc | !hbusreq0 & v3a6b102;
assign v3a70353 = hgrant6_p & v3761fb5 | !hgrant6_p & v377a478;
assign v3758988 = hgrant2_p & v3a2a348 | !hgrant2_p & v3a714ac;
assign v373127a = hmaster1_p & v3a64fce | !hmaster1_p & v3757996;
assign v372abd2 = hmaster0_p & v3a5ba7f | !hmaster0_p & v372e8ff;
assign v3740da1 = hbusreq8 & v3a583cd | !hbusreq8 & v3728f66;
assign v3774359 = hbusreq5_p & v372c08d | !hbusreq5_p & v37541c6;
assign v3a61ecf = hbusreq0 & v3a6f8d7 | !hbusreq0 & v3a5741c;
assign v3a6b873 = hbusreq1_p & v8455ab | !hbusreq1_p & !v3a637dd;
assign v3a6caab = hbusreq8 & v3727195 | !hbusreq8 & v3737411;
assign v3a7109d = hbusreq3_p & v372a414 | !hbusreq3_p & v8455ab;
assign v375eba9 = hbusreq5_p & bf5753 | !hbusreq5_p & v3a6f388;
assign v3807b28 = hmaster2_p & v3a61a7f | !hmaster2_p & v37590a2;
assign v377b5f6 = hgrant4_p & v375d067 | !hgrant4_p & v3767650;
assign v3a55785 = hbusreq0 & v3a62a51 | !hbusreq0 & v377e698;
assign v3763ad3 = stateA1_p & v8455ab | !stateA1_p & !v3807071;
assign v3a70af5 = hbusreq4 & v3739b80 | !hbusreq4 & v3a5b7c2;
assign v3a57e40 = hgrant0_p & v8455b3 | !hgrant0_p & v377e142;
assign v3a607ba = hbusreq7 & v3741e9f | !hbusreq7 & v377a89f;
assign v37247c8 = hbusreq7_p & v37586cd | !hbusreq7_p & !v375a30e;
assign v3724368 = hbusreq0 & v3a621ea | !hbusreq0 & c7355c;
assign v3a6243f = hlock4 & v3a61c45 | !hlock4 & v3764141;
assign v3a5bc5d = hmaster1_p & v3775dbc | !hmaster1_p & v3a5b1ca;
assign v3a5c2ff = hlock8 & v375a0af | !hlock8 & v375d7d2;
assign v3723012 = hbusreq6 & v375da95 | !hbusreq6 & v37386c5;
assign v3770322 = hbusreq5 & v3a7136b | !hbusreq5 & v377077a;
assign v376e040 = hlock0_p & v37401f0 | !hlock0_p & v377374f;
assign v37500e2 = hgrant7_p & v3767dac | !hgrant7_p & v3a6dea7;
assign v376293f = hmaster0_p & v377d107 | !hmaster0_p & v23fdd8d;
assign v3727581 = hmaster2_p & v3767cc9 | !hmaster2_p & v372346b;
assign v37642fa = hbusreq7_p & v37362fd | !hbusreq7_p & v377435f;
assign v37526d6 = hlock2 & v3a590fb | !hlock2 & v3377af7;
assign v3a7097e = hgrant4_p & v3a67c36 | !hgrant4_p & !v8455ab;
assign v377041c = hmaster2_p & v3a6efe8 | !hmaster2_p & v3723af9;
assign v374dc1b = hmaster1_p & v3a6fa8f | !hmaster1_p & v3a6fdb6;
assign v375121b = hbusreq4 & v37566b2 | !hbusreq4 & v8455ab;
assign v3727ee9 = hbusreq5 & v374b2f5 | !hbusreq5 & v3a6fc70;
assign v3a71416 = hbusreq2_p & v3a6eb2a | !hbusreq2_p & v8455ab;
assign v37739af = hgrant5_p & v3778595 | !hgrant5_p & v3a55b16;
assign v3a58353 = hlock6_p & v1e38224 | !hlock6_p & v8455ab;
assign v37467da = hgrant6_p & v37c039c | !hgrant6_p & v3743702;
assign v37670b6 = jx0_p & v3a5d90d | !jx0_p & v3777c6f;
assign v3a6efe2 = hlock0 & v3a552c9 | !hlock0 & v3737d3f;
assign v37315e2 = hgrant4_p & v375805a | !hgrant4_p & !v8455ab;
assign v37457b1 = hbusreq3_p & v375aca9 | !hbusreq3_p & v8455ab;
assign v3a6d3f2 = hmaster0_p & v373ce6d | !hmaster0_p & v3a5ef76;
assign v3a58c2f = hlock0 & v3a7162d | !hlock0 & v37269de;
assign v3a715e3 = hbusreq6 & v372992f | !hbusreq6 & v8455ab;
assign v37370a1 = hbusreq7_p & v3763c0d | !hbusreq7_p & v3a70fcd;
assign v373e10f = hbusreq6_p & v3806e0e | !hbusreq6_p & v3a6a1fd;
assign v3a6f225 = hmaster1_p & v37737aa | !hmaster1_p & v3a6396b;
assign v375c648 = hbusreq8 & v3807472 | !hbusreq8 & v8455ab;
assign v899d31 = hbusreq4 & v372bdca | !hbusreq4 & v375d1d9;
assign v3727d77 = hmaster1_p & v373a4ef | !hmaster1_p & v3a60b37;
assign v37723ed = hlock7_p & v37368bb | !hlock7_p & v374d3b0;
assign v3742e95 = hbusreq8_p & v375f2ab | !hbusreq8_p & !v3a70428;
assign v3722d81 = hbusreq6 & v3a570f5 | !hbusreq6 & v8455ab;
assign v35b77ab = hbusreq5_p & v3a58c15 | !hbusreq5_p & v3a5c576;
assign v3a6f9e3 = hbusreq6 & v373498b | !hbusreq6 & v8455ab;
assign v3a5fae4 = hlock7_p & v377a522 | !hlock7_p & !v3a67d49;
assign v3a70f70 = hbusreq8 & v376f271 | !hbusreq8 & v3768048;
assign v3a6d92f = hmaster2_p & v3758cec | !hmaster2_p & v3a7116b;
assign v377ab40 = hbusreq8 & v374e58f | !hbusreq8 & v3779c26;
assign v3725496 = hmaster2_p & v3807a47 | !hmaster2_p & v376f2a5;
assign v3740409 = hlock3_p & v376eca3 | !hlock3_p & v3a70219;
assign v3a6abdc = hlock6 & v3a6f62c | !hlock6 & v3a6d10a;
assign v3772e8e = hmaster0_p & v3a63777 | !hmaster0_p & v3a709b4;
assign v3750ad1 = hmaster2_p & v3a635ea | !hmaster2_p & v37270bc;
assign v377d01e = hbusreq4_p & v377057c | !hbusreq4_p & v35772a6;
assign v373a005 = hmaster1_p & v3a5cb2c | !hmaster1_p & v8455ab;
assign v373f24b = hgrant4_p & v8455ab | !hgrant4_p & v373cd0a;
assign v3a5e696 = hgrant4_p & v8455ab | !hgrant4_p & v3734aef;
assign v3a6f463 = hmaster2_p & v376d856 | !hmaster2_p & v37521ed;
assign v3a70e5e = hmaster1_p & v37386c6 | !hmaster1_p & v37319c5;
assign v376e9e2 = hgrant0_p & v3764276 | !hgrant0_p & v374053e;
assign v3a5bded = hgrant6_p & v3759b6f | !hgrant6_p & v3724ee0;
assign v373285d = hmaster0_p & v3735974 | !hmaster0_p & v375c621;
assign v376ef9f = hmaster2_p & v3a6f17f | !hmaster2_p & v23fda38;
assign v3777d29 = hbusreq4_p & v376d285 | !hbusreq4_p & !v372c007;
assign v3756716 = hlock2_p & v3750714 | !hlock2_p & v3a59545;
assign v3a6f102 = hgrant6_p & v3760e2e | !hgrant6_p & v3a70ac0;
assign v3a5d678 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a6f8ee;
assign v3a6fd7b = hbusreq4_p & v3a70ee5 | !hbusreq4_p & v8455b0;
assign v372ee70 = hbusreq2 & v3a61f82 | !hbusreq2 & v3a6a82a;
assign v1e382a5 = hbusreq6_p & v3a62a71 | !hbusreq6_p & v3a6f81d;
assign v37368b3 = hlock6 & v3a6f0b8 | !hlock6 & v3a676a9;
assign v3740f92 = hlock6 & v3a6d9fa | !hlock6 & v3806ec4;
assign v3a69d81 = hgrant3_p & v3739018 | !hgrant3_p & v377b68c;
assign v3738ab6 = hbusreq5 & v3a70421 | !hbusreq5 & v8455ab;
assign v3a65847 = hlock5 & v37385c6 | !hlock5 & v3775fa5;
assign v3a6ebf7 = hmaster2_p & v8455ab | !hmaster2_p & !v8455be;
assign v377e26b = hlock2 & v35b708f | !hlock2 & v3a6f02e;
assign v37788d5 = hmaster2_p & v8455e7 | !hmaster2_p & !v376430b;
assign v374f345 = hmaster0_p & v3731f9a | !hmaster0_p & v373931a;
assign v37541a7 = hbusreq4 & v3378c57 | !hbusreq4 & v8455ab;
assign v3723ec6 = hmaster0_p & v373195f | !hmaster0_p & v3756e20;
assign v3a6eaea = jx1_p & v380a20c | !jx1_p & v372dd14;
assign v3732510 = hmaster0_p & v376c224 | !hmaster0_p & !v8455e7;
assign v37266a0 = hbusreq5_p & v3a5d438 | !hbusreq5_p & v37247b2;
assign v3744deb = jx0_p & v376d06c | !jx0_p & v8455ab;
assign v3748e82 = hbusreq7_p & v3a6ff88 | !hbusreq7_p & v3a708a1;
assign v3a6fe80 = hbusreq0_p & v37775c4 | !hbusreq0_p & b27f78;
assign v372e751 = hgrant3_p & v377dd3b | !hgrant3_p & v375f52b;
assign v374ea10 = hgrant7_p & v3a6e2ce | !hgrant7_p & v372ab42;
assign v377073f = hbusreq7_p & v376198e | !hbusreq7_p & v375dd4c;
assign v3765385 = hmaster2_p & v3a6fb30 | !hmaster2_p & v8455ab;
assign v3a70ce6 = hbusreq6_p & v3a5ce1e | !hbusreq6_p & v374765b;
assign v37232a3 = hmaster0_p & v3a5af94 | !hmaster0_p & v3728045;
assign v3a66a3a = hbusreq5_p & v3a70ea2 | !hbusreq5_p & !v374e168;
assign v3740060 = hbusreq3_p & v39eb4de | !hbusreq3_p & v377437a;
assign v3806db2 = hbusreq8 & v37679b0 | !hbusreq8 & v3a6051e;
assign v376d7d5 = hmaster1_p & v37730d2 | !hmaster1_p & v37546a9;
assign v20930ad = hbusreq2_p & v375783c | !hbusreq2_p & v37401ce;
assign v376d007 = hmaster1_p & v377703d | !hmaster1_p & v8455e7;
assign v375411b = hgrant4_p & v8455ab | !hgrant4_p & v3a66f35;
assign v373c49e = hbusreq2 & v3a54a76 | !hbusreq2 & v8455ab;
assign v374e55f = jx0_p & v3731ab1 | !jx0_p & v8455ab;
assign v374eaf4 = hmaster2_p & bbeeaf | !hmaster2_p & v3750dd3;
assign v3a6ba6a = hbusreq6_p & v3a70649 | !hbusreq6_p & v3a704f1;
assign v3725f24 = hbusreq2 & v3742d54 | !hbusreq2 & v372da76;
assign v376ab53 = hbusreq5_p & v376ff46 | !hbusreq5_p & v3a666bb;
assign v3a5664b = hbusreq7 & v3723f33 | !hbusreq7 & v8455ab;
assign v3806b0b = hbusreq7 & d52046 | !hbusreq7 & v373216d;
assign v2aca978 = hlock2_p & v3760549 | !hlock2_p & v8455ab;
assign v3a6eb3f = hlock0_p & v1e38275 | !hlock0_p & v3a7011c;
assign v2619b43 = hbusreq2_p & v3a5b289 | !hbusreq2_p & !v8455ab;
assign v3a713da = hbusreq5_p & v3a6e7ed | !hbusreq5_p & v3a5b514;
assign v3a70cee = hgrant4_p & v8455ab | !hgrant4_p & v3757009;
assign v3a6dea6 = hlock8_p & v3777b18 | !hlock8_p & v8455c7;
assign v3a6fbc4 = hmaster1_p & v3a70d99 | !hmaster1_p & v39eb4a5;
assign v3733483 = hgrant5_p & v373ab60 | !hgrant5_p & v3a70433;
assign v372ce4a = hmaster1_p & v373dc55 | !hmaster1_p & v377dc60;
assign aeff0f = hmaster0_p & v372b390 | !hmaster0_p & a97cd0;
assign v3a715a8 = hlock4 & v3739a3b | !hlock4 & v377cdf0;
assign v372bc50 = hmaster2_p & v3a70ca8 | !hmaster2_p & v372adb5;
assign v3a70e5c = hbusreq8 & v3772c8e | !hbusreq8 & !v3a70700;
assign v3733955 = jx0_p & v376beea | !jx0_p & v377c9c3;
assign v375dd2b = hgrant6_p & v8455ab | !hgrant6_p & v37613d3;
assign v372745b = hgrant4_p & v37300a5 | !hgrant4_p & v3a6a435;
assign v37362dc = hbusreq7_p & v3734279 | !hbusreq7_p & v3740be8;
assign v86d3dc = hgrant3_p & v3a61cbf | !hgrant3_p & v3a6fac4;
assign v375e4a0 = hlock2 & v3806ff0 | !hlock2 & v375df25;
assign v3a627d8 = hgrant0_p & v377714d | !hgrant0_p & !v3776a6e;
assign v3761362 = hlock6_p & v3a7094d | !hlock6_p & v3759daf;
assign v3a6762b = hbusreq4 & v3730e7d | !hbusreq4 & v3a62a6d;
assign v3a2a2ee = hbusreq2 & v3a299d4 | !hbusreq2 & v8455ab;
assign v372f649 = hmaster1_p & v3728419 | !hmaster1_p & v376dce5;
assign v3807ae8 = hmaster2_p & v3753dab | !hmaster2_p & v37796c6;
assign v372c85e = hmaster0_p & v3779680 | !hmaster0_p & v3a5c983;
assign v373dbc5 = hgrant2_p & v3a6c33a | !hgrant2_p & !v3730b77;
assign v3769fe3 = hbusreq7_p & v3769dcb | !hbusreq7_p & v3a70919;
assign v376592b = hmaster1_p & v37363ae | !hmaster1_p & v3a5f869;
assign v37698c3 = hbusreq5_p & v3a5f711 | !hbusreq5_p & v3737ce3;
assign v3749674 = hlock6 & v375b90a | !hlock6 & v3a5bc77;
assign v3a6fd79 = hburst1 & v2aca977 | !hburst1 & v373d357;
assign v373d5b7 = hbusreq5 & v377aed1 | !hbusreq5 & v3a5ef9d;
assign v3747c23 = hmaster2_p & v374f307 | !hmaster2_p & v3723b00;
assign v372a94e = hgrant6_p & v3a55efa | !hgrant6_p & v3577338;
assign v37685bb = hbusreq1_p & v375d5f3 | !hbusreq1_p & v8455b0;
assign v3739f29 = hbusreq4_p & v3755420 | !hbusreq4_p & v374673a;
assign v3a66387 = hgrant4_p & v3a5e63b | !hgrant4_p & v3a68d49;
assign v372e712 = hmaster2_p & v3740890 | !hmaster2_p & !v377957e;
assign v3778419 = hmaster0_p & v377a3bd | !hmaster0_p & v373d9a2;
assign v3a6f60c = hmaster1_p & v374502e | !hmaster1_p & v3a5f1e8;
assign v3a6a713 = hbusreq4_p & v373fad7 | !hbusreq4_p & v3a57156;
assign v3a2a14e = hbusreq0 & v375e03c | !hbusreq0 & v37777ba;
assign v373a1d7 = hmaster2_p & v37457b1 | !hmaster2_p & v8455ab;
assign v374b204 = hmaster2_p & v373a27c | !hmaster2_p & v374362e;
assign v37528fd = hbusreq4_p & v377eaf2 | !hbusreq4_p & v374a637;
assign v377c2e6 = hmastlock_p & v377f108 | !hmastlock_p & v8455ab;
assign v376d902 = hlock4 & v3730451 | !hlock4 & v375f302;
assign v3a70cc9 = hmaster2_p & b66740 | !hmaster2_p & !v3a6f312;
assign v3a6cd48 = hlock8 & v3a71492 | !hlock8 & v3758b56;
assign v3a702d0 = hmaster1_p & v3a6e124 | !hmaster1_p & v3a6bb65;
assign v3a6ddc7 = hbusreq7 & v3808e88 | !hbusreq7 & v372aaf8;
assign v37736a6 = hbusreq0_p & v376ef42 | !hbusreq0_p & v3733e9e;
assign hgrant0 = !v3a6c363;
assign v3779060 = hbusreq1_p & v3a68c1f | !hbusreq1_p & v3a57f59;
assign v3731370 = hbusreq8 & v3769ce7 | !hbusreq8 & v37582e0;
assign v3a29706 = hgrant3_p & v8455be | !hgrant3_p & v376b8e9;
assign v3767744 = hmaster0_p & v377dedb | !hmaster0_p & !v2ff9391;
assign v3a6f52c = hlock4 & v3a646ae | !hlock4 & v3a6582b;
assign v373b6dd = hbusreq8_p & v3a65b00 | !hbusreq8_p & v3a70254;
assign v37464f3 = hmaster1_p & v375c48c | !hmaster1_p & v38064e3;
assign v375cfd9 = hlock7 & v3a675eb | !hlock7 & v3a5f80f;
assign v3a6f6f4 = hgrant3_p & v3774c1b | !hgrant3_p & !v3a6494a;
assign v37265f6 = hgrant2_p & v3a6c33a | !hgrant2_p & !v3752201;
assign v3752348 = hbusreq7 & v372a79d | !hbusreq7 & v377c620;
assign v377053a = hbusreq8_p & b1f7c8 | !hbusreq8_p & v37571fc;
assign v37651fe = hbusreq7 & v374bbaf | !hbusreq7 & v3a62a6d;
assign v3a70dfb = hbusreq0_p & v37317a9 | !hbusreq0_p & v3a68d2e;
assign v372d51c = hmaster2_p & v375f452 | !hmaster2_p & v37572c1;
assign v3a7164a = hgrant6_p & v8455ab | !hgrant6_p & v3a6adb2;
assign v373b548 = hbusreq4 & v37678fc | !hbusreq4 & v8455b3;
assign v3a645d7 = hlock2_p & v373e046 | !hlock2_p & v8455b0;
assign v3a70a28 = start_p & v8455ab | !start_p & v3766cf9;
assign v372b74c = hgrant0_p & v3723cff | !hgrant0_p & v8455ab;
assign v37441b5 = hgrant0_p & v9ed516 | !hgrant0_p & v3a65934;
assign v3a6ff4c = hgrant2_p & v375ca6c | !hgrant2_p & v3a54a76;
assign v375f1db = jx0_p & v3764a58 | !jx0_p & v37559d6;
assign v373c23e = hbusreq6 & v3731991 | !hbusreq6 & v3a62a6d;
assign v37316d9 = hbusreq2_p & v3a554b9 | !hbusreq2_p & !v3752397;
assign v1e379ef = hbusreq4 & v377a5a9 | !hbusreq4 & v374a637;
assign v37451b8 = hmaster2_p & v3a702c2 | !hmaster2_p & v376d374;
assign v37573c5 = hbusreq7_p & v3734279 | !hbusreq7_p & v3a544c4;
assign v3a70d8a = hgrant6_p & v3a6c7fe | !hgrant6_p & v3a5919f;
assign v35b7174 = hbusreq8 & v3a6fb3f | !hbusreq8 & v3764e55;
assign v374ea19 = hbusreq5 & v3a663ef | !hbusreq5 & v3a67471;
assign v376dce5 = hbusreq5_p & v3741280 | !hbusreq5_p & v374c870;
assign v3729b2e = hbusreq4 & v375139d | !hbusreq4 & !v374742c;
assign v3a71693 = hmaster1_p & v3a6ff12 | !hmaster1_p & v375b0ad;
assign v374ca62 = hgrant4_p & v8455ab | !hgrant4_p & v3a6403e;
assign v374021a = hlock4 & v373b51b | !hlock4 & v3a704b0;
assign v3a713d2 = hmaster1_p & v373a4e4 | !hmaster1_p & v376f182;
assign v3746a04 = hlock0_p & v377b24b | !hlock0_p & v3768add;
assign v3744ea3 = hbusreq4_p & v3a6ff80 | !hbusreq4_p & !v3725f77;
assign v37314fa = hgrant4_p & v376f2f8 | !hgrant4_p & v3a6fd37;
assign v377a468 = hmaster1_p & v3743677 | !hmaster1_p & !v377559f;
assign v373c58c = hmaster0_p & v37358ab | !hmaster0_p & v3a5d7ba;
assign v3747141 = hmaster1_p & v3a5e000 | !hmaster1_p & !v3a67e97;
assign v3a6f909 = hburst0 & v8455ab | !hburst0 & v3a70cd5;
assign v3a6440f = hgrant3_p & v373e521 | !hgrant3_p & v3733ba1;
assign v373a265 = hbusreq5_p & v3a2abf4 | !hbusreq5_p & v8455ab;
assign v3a57506 = hlock4_p & v3748ca3 | !hlock4_p & !v8455ab;
assign v374eda5 = hgrant6_p & v37418ac | !hgrant6_p & v375aaf3;
assign v375f2ab = hlock8_p & v3a6f7b8 | !hlock8_p & !v372428a;
assign v375e6a0 = hmaster2_p & v3a63bb7 | !hmaster2_p & v3a5a8ce;
assign v37386c6 = hgrant4_p & v3a635ea | !hgrant4_p & v376ca86;
assign v3a6be9f = hbusreq7_p & v3764448 | !hbusreq7_p & v3722d8b;
assign v372509d = hbusreq8_p & v3762729 | !hbusreq8_p & v37482f5;
assign v3748353 = hlock6 & v3760e46 | !hlock6 & v3a7062b;
assign v3a6d810 = hbusreq3_p & v3a635ea | !hbusreq3_p & v37744c1;
assign v3a6514f = hbusreq8_p & v3755549 | !hbusreq8_p & v3756aa3;
assign v3744f35 = hlock0_p & v8455e1 | !hlock0_p & v8455ab;
assign v3a70ed4 = hbusreq5 & v3a6f321 | !hbusreq5 & v8455ab;
assign v3734ec1 = hlock4_p & v3a7136f | !hlock4_p & !v8455ab;
assign v37685c3 = hmaster2_p & v3727943 | !hmaster2_p & v376d1bb;
assign v3724e30 = hbusreq6_p & v3a6c98c | !hbusreq6_p & v8455ab;
assign v372e48a = hbusreq3_p & v3a7150d | !hbusreq3_p & !v376d45f;
assign v3724784 = hmaster2_p & v37600c0 | !hmaster2_p & v3a67fea;
assign v3a62d5d = hmaster0_p & v3a635ea | !hmaster0_p & v3737202;
assign v3740742 = hbusreq7_p & v372641e | !hbusreq7_p & v3a6bce9;
assign v3a67d2e = hgrant1_p & v8455ab | !hgrant1_p & !v37271f9;
assign v3a707e1 = hbusreq7 & v373bbe6 | !hbusreq7 & v3a6abfe;
assign v3a65b53 = hgrant6_p & v3a6f17e | !hgrant6_p & v37288db;
assign v37662f4 = hgrant8_p & v1e37c79 | !hgrant8_p & v3a70968;
assign v3a6602d = hmaster1_p & v3a661fe | !hmaster1_p & v3727c3c;
assign v376746b = hgrant5_p & v3a71285 | !hgrant5_p & v3a5c2d6;
assign v3809ee9 = hbusreq2_p & v3734100 | !hbusreq2_p & v3a5bb64;
assign v376d89f = hmaster0_p & v3a5bf28 | !hmaster0_p & v23fd7a9;
assign v3a70a82 = hmaster0_p & v373bc28 | !hmaster0_p & v3722caa;
assign v3a5d646 = hlock8 & v376d258 | !hlock8 & v37644ee;
assign v380776b = hmaster1_p & v373695f | !hmaster1_p & v3a56323;
assign v374bb64 = hbusreq5_p & v3778ca0 | !hbusreq5_p & v8455ab;
assign v376e7c1 = hlock8 & v376ae9f | !hlock8 & v372cdd4;
assign v373a6ba = hmaster2_p & v3775dbc | !hmaster2_p & v3a5a807;
assign v372b6c4 = hgrant0_p & v8455ab | !hgrant0_p & v1e37bdd;
assign v3773c5d = hbusreq5_p & v373a327 | !hbusreq5_p & v373b7b5;
assign v376f9a1 = hmaster0_p & v372455c | !hmaster0_p & v3a59ed6;
assign v3752cac = hmaster0_p & v9de657 | !hmaster0_p & v3736184;
assign v37648fb = hmaster1_p & v3772c0a | !hmaster1_p & v8455e7;
assign v373c545 = hmaster2_p & v372ad6d | !hmaster2_p & v3a5a01b;
assign v376c4c9 = hbusreq5_p & v93c94e | !hbusreq5_p & v376c652;
assign v3a6ca1d = hbusreq3_p & v3a6acbb | !hbusreq3_p & a21c18;
assign v3743d23 = hbusreq6 & v37482f8 | !hbusreq6 & v8455ab;
assign v373c074 = hmaster1_p & v377c15d | !hmaster1_p & v372b077;
assign v377a4c1 = hgrant6_p & v8455ab | !hgrant6_p & v375bd53;
assign v39eb4a7 = hgrant2_p & v3a5eadd | !hgrant2_p & v377c039;
assign v375ab99 = hlock0 & v373abde | !hlock0 & v3a63a46;
assign v37c03ad = hmaster2_p & v3a635ea | !hmaster2_p & v375d800;
assign v3747212 = hmaster2_p & v3754ec1 | !hmaster2_p & v3a55cd6;
assign v372ef40 = hgrant2_p & v3a70326 | !hgrant2_p & v377d4ab;
assign v377bd97 = hbusreq2 & v37738fc | !hbusreq2 & v35b774b;
assign v3a6eb7b = hbusreq4_p & v3a6f4c7 | !hbusreq4_p & v3748d67;
assign v37494ed = hbusreq5 & v376c0d8 | !hbusreq5 & v8455ab;
assign v37664a1 = hlock0 & v373f3b5 | !hlock0 & v3767385;
assign v374637b = hbusreq7_p & v3771303 | !hbusreq7_p & v376749b;
assign v37440e4 = hbusreq5_p & v37375e2 | !hbusreq5_p & v8455ab;
assign v372700a = hmaster2_p & v8455ab | !hmaster2_p & v375b5b4;
assign v375025f = hmaster0_p & v8455c9 | !hmaster0_p & !v3903ee2;
assign v375b234 = hmaster1_p & v374d4e6 | !hmaster1_p & v373cfd0;
assign v3731caa = hgrant4_p & v37311d8 | !hgrant4_p & v3a70d7f;
assign v375a6d3 = hgrant4_p & v8455ab | !hgrant4_p & v372452c;
assign v375a510 = hbusreq5_p & v3774bad | !hbusreq5_p & v380760a;
assign v37484b6 = hbusreq7 & v3a7079c | !hbusreq7 & v3734279;
assign v37509a9 = hmaster2_p & v3758cf5 | !hmaster2_p & acc1e3;
assign v3a699d3 = hbusreq2 & v3753dab | !hbusreq2 & v8455ab;
assign v3a6f9e7 = hmaster0_p & v3724394 | !hmaster0_p & v3748b43;
assign v3778211 = hmaster1_p & v8455ab | !hmaster1_p & !v37356a7;
assign v372a5c8 = hgrant2_p & v3a6c80b | !hgrant2_p & v37273c2;
assign v3a6f8ec = hmaster2_p & v8455ab | !hmaster2_p & v3767f33;
assign v3778baf = hbusreq8 & v3a6fb24 | !hbusreq8 & v37302b7;
assign v23fe1ad = hmaster0_p & v377982c | !hmaster0_p & v337902c;
assign v3764fd7 = hmaster1_p & v3770b6c | !hmaster1_p & v377559f;
assign v376f569 = hbusreq0 & v3a6f586 | !hbusreq0 & v8455ab;
assign v3769a8e = hbusreq4_p & v3a70ad6 | !hbusreq4_p & v37562a5;
assign v3a68b7d = hmaster2_p & v373561e | !hmaster2_p & v3731b41;
assign v373edd6 = hbusreq5 & v37281ca | !hbusreq5 & v8455ab;
assign v3257687 = hbusreq8 & v373f3e4 | !hbusreq8 & v376195b;
assign v3729178 = hmaster2_p & v375a1ab | !hmaster2_p & v372d2dc;
assign v3776eff = hgrant4_p & v8455bd | !hgrant4_p & v375c50a;
assign v373a803 = hbusreq3_p & v3a6b691 | !hbusreq3_p & v3a5cd20;
assign v3728823 = hlock4 & v374a4ca | !hlock4 & v3756483;
assign v372da78 = hmaster2_p & v375b2e2 | !hmaster2_p & v374355e;
assign v3749628 = hmaster0_p & v3a6ff61 | !hmaster0_p & v3758ff0;
assign v39eaff9 = hmaster2_p & v376fe6e | !hmaster2_p & v3778b19;
assign v3a64bc4 = hmaster2_p & c6a502 | !hmaster2_p & v3a6ef4a;
assign v372edd9 = hgrant4_p & v3a6f4de | !hgrant4_p & v3733599;
assign v37369df = hmaster1_p & v3a6e7b3 | !hmaster1_p & v376537c;
assign v37461d9 = hmaster2_p & v3a635ea | !hmaster2_p & v37356b4;
assign v377e30e = hgrant5_p & v3a57037 | !hgrant5_p & v376cddf;
assign v373a25b = hbusreq2_p & v377fb84 | !hbusreq2_p & bb611d;
assign v3757091 = hbusreq4 & v3753d51 | !hbusreq4 & v374165f;
assign v3744417 = hbusreq4_p & v3a70cc0 | !hbusreq4_p & v3a56864;
assign v3748efb = hmaster1_p & v37738ae | !hmaster1_p & v3a6a73a;
assign v376362f = hlock0 & v37496fa | !hlock0 & v375a8ad;
assign v3a6eb66 = hbusreq0_p & v376f9a8 | !hbusreq0_p & v376d856;
assign v376b57f = hgrant6_p & v8455ab | !hgrant6_p & v3779746;
assign v3727507 = hbusreq1 & v374e2a1 | !hbusreq1 & v3748797;
assign v376cab5 = hbusreq7_p & v3732853 | !hbusreq7_p & v376a74a;
assign v3a6f8a8 = hbusreq5 & v3763175 | !hbusreq5 & v8455ab;
assign v377d766 = hmaster2_p & v2ff9190 | !hmaster2_p & v373f72a;
assign v3744d52 = hlock0_p & v35772c9 | !hlock0_p & !v8455ab;
assign v3770be3 = hgrant3_p & v8455ab | !hgrant3_p & v3749e33;
assign v3738491 = hbusreq4_p & v3a67ecb | !hbusreq4_p & v3a5741c;
assign v376702a = hmaster0_p & v3a59819 | !hmaster0_p & v375f014;
assign v3a6427b = hbusreq7 & v375a76e | !hbusreq7 & v377b774;
assign v375c50a = hgrant6_p & v8455bd | !hgrant6_p & v3a58b3f;
assign v3773982 = hbusreq2 & v375fa8b | !hbusreq2 & v377efdc;
assign v3a645b4 = hlock4 & v374aa90 | !hlock4 & v3762388;
assign v375dc01 = hgrant4_p & v3a6c21d | !hgrant4_p & v3a62cff;
assign v3769d19 = hgrant1_p & v3a57445 | !hgrant1_p & v375003c;
assign v3a6efac = hbusreq6 & v3766a74 | !hbusreq6 & v3767690;
assign v37281d0 = hbusreq3 & v3733471 | !hbusreq3 & v8455ab;
assign v375d8af = hmaster1_p & v3a70a65 | !hmaster1_p & v3a69ad9;
assign v376a5c1 = hmaster1_p & v3779183 | !hmaster1_p & v3a59f8c;
assign v373e01f = hbusreq5_p & v3a70423 | !hbusreq5_p & v3a60d50;
assign v3749ab1 = hbusreq5 & v3a67996 | !hbusreq5 & v8455ab;
assign v377b461 = hgrant4_p & v377498e | !hgrant4_p & v375e6b2;
assign v3a6f7fe = hbusreq7_p & v37290fa | !hbusreq7_p & !v3766a37;
assign v3809adf = stateA1_p & v8455ab | !stateA1_p & !v3a708aa;
assign v3a6f32f = hbusreq1_p & v37773c4 | !hbusreq1_p & v8455ab;
assign v373d746 = hbusreq8_p & v1e38301 | !hbusreq8_p & v372ff75;
assign v37474c2 = hgrant2_p & v8455e7 | !hgrant2_p & !v3a6d219;
assign v3749649 = hmaster2_p & d44200 | !hmaster2_p & v3a7156d;
assign v376d6f9 = hbusreq2 & v3731487 | !hbusreq2 & v375c1d1;
assign v3725475 = hbusreq2_p & v3733e9e | !hbusreq2_p & v1e38224;
assign v376e87e = hmaster2_p & v3723b5b | !hmaster2_p & v3756304;
assign v3a71227 = hbusreq8_p & v3a635ea | !hbusreq8_p & v37712c2;
assign v3734e23 = hlock7 & a0a219 | !hlock7 & v375bf36;
assign v3a645ca = hbusreq3_p & v3a69487 | !hbusreq3_p & v375d288;
assign v3769ed3 = hbusreq4_p & v37432c6 | !hbusreq4_p & !v37521ed;
assign v3a63b26 = hlock7 & v3a6c4bb | !hlock7 & v375973d;
assign v37460de = hbusreq5 & v3a6fd64 | !hbusreq5 & !v3a6f826;
assign v37291e7 = hmaster2_p & v3a7039a | !hmaster2_p & v3a6f1e4;
assign v3761472 = hmaster0_p & v3a6ffca | !hmaster0_p & v377ee74;
assign v3748481 = hbusreq0_p & v3747302 | !hbusreq0_p & v23fe0bb;
assign v3763344 = hlock2_p & v2ff9190 | !hlock2_p & v8455ab;
assign v3a70125 = hbusreq6 & v376c351 | !hbusreq6 & v3767266;
assign v372414d = hgrant4_p & v8455ab | !hgrant4_p & v3a5f9e6;
assign v374fab7 = hmaster0_p & v3a70899 | !hmaster0_p & v8455ab;
assign v2619b54 = hbusreq6_p & v3741f39 | !hbusreq6_p & v325b5e0;
assign v376e500 = hbusreq3_p & v3a68c1f | !hbusreq3_p & !v3807bf8;
assign v37621b5 = hlock6_p & v3769cc2 | !hlock6_p & v8455ab;
assign v3a6f4da = hbusreq5_p & v3742ca7 | !hbusreq5_p & v3a67b76;
assign baf7ba = hlock2 & v3727ffa | !hlock2 & v37275ef;
assign v3a66d14 = hmaster2_p & v3a5a807 | !hmaster2_p & !v3a703c3;
assign v3a55173 = hlock6_p & v374caab | !hlock6_p & v373399e;
assign v37646e1 = hgrant4_p & v8455ab | !hgrant4_p & v372ab23;
assign v3a59b9e = hbusreq6_p & v376e9c5 | !hbusreq6_p & v3751f46;
assign v3764bf2 = hmaster2_p & v3a635ea | !hmaster2_p & v3a70b92;
assign v3a6ff5b = hgrant4_p & v376a6f1 | !hgrant4_p & v37388a7;
assign v374fe1a = hbusreq6_p & v376d1e2 | !hbusreq6_p & v37348ee;
assign cee4af = hbusreq3_p & v37796c6 | !hbusreq3_p & v3a6fa39;
assign v3a70fe8 = hbusreq0 & v3a62070 | !hbusreq0 & v3a568e4;
assign a708cc = hbusreq4 & v3a68e5d | !hbusreq4 & v8455ab;
assign v3760b7a = hbusreq6_p & v3a6ef49 | !hbusreq6_p & v375b34f;
assign v3a6e78d = start_p & v3776483 | !start_p & v3a6b463;
assign b8f5a8 = hmaster0_p & v3a635ea | !hmaster0_p & v3a70665;
assign v3747f81 = hbusreq0 & v3a5b079 | !hbusreq0 & v373f950;
assign v3a6fad2 = hgrant4_p & v8455ab | !hgrant4_p & v37bfc4d;
assign v3736cb3 = hbusreq4_p & v37522d3 | !hbusreq4_p & v3a5be57;
assign a96343 = hgrant4_p & v3723b5b | !hgrant4_p & b65b94;
assign v37315c8 = hgrant6_p & v8455ab | !hgrant6_p & v377c923;
assign v375f3bd = hbusreq2 & v37521ed | !hbusreq2 & !v8455ab;
assign v376bc5b = hbusreq8_p & v374d1d7 | !hbusreq8_p & v3745e71;
assign v375ac88 = hbusreq7 & v1e373d9 | !hbusreq7 & v3768734;
assign v3765784 = hbusreq4 & v3732797 | !hbusreq4 & v1e37bf6;
assign v376277f = hmaster1_p & v3768dbc | !hmaster1_p & v3a66210;
assign v3a70c73 = hgrant1_p & v3a68c1f | !hgrant1_p & !v372c11d;
assign v3a715b7 = hmaster2_p & v3a70374 | !hmaster2_p & v3a6fac0;
assign v20930b8 = hlock6 & v374af2f | !hlock6 & v3a6e8d4;
assign v3778bb4 = hmaster0_p & v8455ab | !hmaster0_p & v3a6ec30;
assign v372873a = hmaster0_p & v3a5a24b | !hmaster0_p & v1e37b47;
assign v3768a9c = hbusreq4_p & v3747302 | !hbusreq4_p & v3a70a88;
assign v37647e7 = hbusreq3_p & v3757dad | !hbusreq3_p & v8455b0;
assign v372e6f4 = hgrant2_p & v37609e7 | !hgrant2_p & v8455ab;
assign v3a5e035 = hmaster1_p & v3a6f8bd | !hmaster1_p & v3a5b6b0;
assign v373dcdd = hmaster0_p & v3736969 | !hmaster0_p & v375fb03;
assign v3a65383 = jx3_p & v37769d5 | !jx3_p & v3a610f7;
assign v374944b = hlock2 & v37551e3 | !hlock2 & v372f76a;
assign v2925c39 = stateA1_p & v376faea | !stateA1_p & !v3739e55;
assign v37745e9 = hmaster1_p & v37272ca | !hmaster1_p & v3a6fd9b;
assign v375a771 = hgrant6_p & v37332c8 | !hgrant6_p & v3a7057f;
assign v377dca9 = hbusreq5 & v3a5948f | !hbusreq5 & v8455ab;
assign v375fd8d = hbusreq0 & v3a71527 | !hbusreq0 & v1e37cd6;
assign v37375e2 = hbusreq5 & v37233f1 | !hbusreq5 & v8455ab;
assign a4a7a5 = stateG10_1_p & v35772a5 | !stateG10_1_p & !v375aa47;
assign v376e677 = hgrant3_p & v8455ab | !hgrant3_p & v37257f8;
assign v3a707de = hbusreq1_p & v3732817 | !hbusreq1_p & v3741d00;
assign v3a60faf = hgrant2_p & v3a61a7f | !hgrant2_p & v373dd9b;
assign v37638f9 = hbusreq8_p & v3a71386 | !hbusreq8_p & v1e37776;
assign v372d780 = jx0_p & v372779c | !jx0_p & v372de54;
assign v35b7d97 = jx0_p & v3a6fe8c | !jx0_p & v3a70ad1;
assign v375fdb5 = hmaster0_p & v37328b0 | !hmaster0_p & v377a985;
assign v375c939 = hlock3_p & v3a5acd9 | !hlock3_p & v3a6958b;
assign v3a7059b = hgrant4_p & v3758d3f | !hgrant4_p & v373d214;
assign v377bf7b = hmaster1_p & v376ae7f | !hmaster1_p & v37558f2;
assign v3a6fd75 = hbusreq5 & v38099a4 | !hbusreq5 & v3a60d11;
assign v3742c52 = hbusreq2_p & v375d40b | !hbusreq2_p & v3a6f37c;
assign v37241a0 = hmaster1_p & v3756cf2 | !hmaster1_p & v372e8f2;
assign v3a5f9f2 = hbusreq3_p & v3722b74 | !hbusreq3_p & v39a536d;
assign v377a2f3 = hlock5_p & v3a674b3 | !hlock5_p & v3758466;
assign v373e924 = hmaster1_p & v8455b5 | !hmaster1_p & v3a6a6c6;
assign v37280b2 = hmaster0_p & v3a7071a | !hmaster0_p & v374d339;
assign v373fdce = hbusreq8 & v8455b0 | !hbusreq8 & v3750fa9;
assign v375fb9d = hmaster0_p & v377bf88 | !hmaster0_p & v3a6abf7;
assign v377ec59 = hbusreq4_p & v3a70725 | !hbusreq4_p & v2092f41;
assign v377b84e = hlock2 & v3753b5e | !hlock2 & v3770ae6;
assign v3a6fb7c = hbusreq6_p & v372cda0 | !hbusreq6_p & v8455ab;
assign v3a715d1 = hmaster0_p & v376d774 | !hmaster0_p & !v374514c;
assign v3763a4a = hmaster2_p & v374f658 | !hmaster2_p & v372424e;
assign v373635b = hbusreq7_p & v37651fe | !hbusreq7_p & v3740dcc;
assign v3732b92 = hbusreq5 & v1e37cba | !hbusreq5 & v3765bf4;
assign v3809380 = hmaster1_p & v377e4d8 | !hmaster1_p & v3734d9a;
assign v372cb06 = hbusreq5_p & v37699c7 | !hbusreq5_p & !v3a70d09;
assign v3758aec = hbusreq4_p & v3a5a510 | !hbusreq4_p & !v1e382e7;
assign v3a61ad3 = hgrant7_p & v372766c | !hgrant7_p & v380877d;
assign v3761f69 = hbusreq7 & v376d795 | !hbusreq7 & v3753b70;
assign v3a59905 = hmaster2_p & v3756203 | !hmaster2_p & v3760740;
assign v372d630 = hgrant2_p & v3a6c80b | !hgrant2_p & v377109d;
assign v3a71050 = hbusreq5_p & v373d5e7 | !hbusreq5_p & v3a5455e;
assign v375981e = hbusreq0 & v3a6c60e | !hbusreq0 & v8455ab;
assign v126f91f = hbusreq6_p & v3736ded | !hbusreq6_p & v377169f;
assign v377bac2 = hbusreq5_p & v3a712c6 | !hbusreq5_p & v8455ab;
assign v3a6f868 = hmaster0_p & v8455ab | !hmaster0_p & v3a70ac2;
assign v3a710aa = hbusreq4 & v375c44b | !hbusreq4 & v8455ab;
assign v373158e = hmaster1_p & v3761bd1 | !hmaster1_p & v373c23c;
assign v373e9a9 = hgrant3_p & v8455be | !hgrant3_p & v3a7066e;
assign v3a70fa7 = hbusreq6_p & v3a60787 | !hbusreq6_p & !v377cfd9;
assign v3a70b5e = hbusreq4_p & v38072fd | !hbusreq4_p & v3756205;
assign v3a62251 = start_p & v3746c8d | !start_p & v3730383;
assign v375b400 = hbusreq5_p & v3766b26 | !hbusreq5_p & v3779c8e;
assign v377e7ac = hmaster0_p & v3765466 | !hmaster0_p & v37665e1;
assign v3747fdb = hmaster2_p & v376bade | !hmaster2_p & v3a57959;
assign v373827a = hbusreq8_p & v377cd7f | !hbusreq8_p & v373dbbb;
assign v3a61e9a = hbusreq4_p & v3726d1f | !hbusreq4_p & v373eaee;
assign v377dd4e = hbusreq4_p & v376b1f6 | !hbusreq4_p & v8455ab;
assign v374f329 = hgrant4_p & v377edba | !hgrant4_p & v374ae4a;
assign v377c56c = hlock8_p & v3733e5a | !hlock8_p & !v377bcfc;
assign v3763f3f = hmaster3_p & v3a575d5 | !hmaster3_p & v3737e97;
assign v37259cc = hbusreq4 & v8455e1 | !hbusreq4 & v8455ab;
assign v373b600 = hgrant6_p & v377b6ce | !hgrant6_p & v377e158;
assign v375bfe5 = hmaster2_p & v3a6dc83 | !hmaster2_p & v376926f;
assign v3a5e7c0 = hbusreq6_p & v3a57bb0 | !hbusreq6_p & v376730e;
assign v374e64f = hbusreq2_p & v3a6ca24 | !hbusreq2_p & v8455ab;
assign v3a55630 = hgrant2_p & v3728eef | !hgrant2_p & v374f1c3;
assign v3a7060c = hbusreq5_p & v38076cf | !hbusreq5_p & v3a6fce0;
assign v373a3e4 = hbusreq3 & aab2b0 | !hbusreq3 & v8455e7;
assign v3742d54 = hlock3 & v3731399 | !hlock3 & v3779fec;
assign v9cbad6 = hbusreq6 & v3a6f4d0 | !hbusreq6 & v8455ab;
assign v3a71610 = hbusreq7 & v374bd7d | !hbusreq7 & v376e66e;
assign v373b732 = hlock5_p & v375b48b | !hlock5_p & !v8455ab;
assign v37788a6 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f12a;
assign v3a652a2 = hmaster0_p & v3773b30 | !hmaster0_p & v3a6ab7f;
assign v375d1a1 = hmaster2_p & v374fb58 | !hmaster2_p & v37648af;
assign v3724c8c = hmaster1_p & v3a5b289 | !hmaster1_p & v374801c;
assign v3a71180 = hmaster2_p & v3a635ea | !hmaster2_p & v3a57959;
assign v37290a1 = hgrant6_p & v372ffaa | !hgrant6_p & v37425a1;
assign v373c050 = hmaster0_p & v8455ca | !hmaster0_p & !v3a5a807;
assign v3a71667 = hmaster2_p & v3a66ade | !hmaster2_p & v3732e59;
assign v3a5c0f8 = hmaster3_p & v3736fb1 | !hmaster3_p & !v3a681f5;
assign v3a6f806 = hbusreq3_p & v3a5495d | !hbusreq3_p & v8455ab;
assign v373100d = hlock5 & v3a650a6 | !hlock5 & v3722a46;
assign v3a6d31d = hbusreq5_p & v373195f | !hbusreq5_p & v3774647;
assign v372fe8b = hbusreq4_p & v3a70a70 | !hbusreq4_p & v3a582d8;
assign v375b990 = hburst0 & v3745b85 | !hburst0 & !v8455ab;
assign v3723e64 = hgrant6_p & v376495e | !hgrant6_p & v3751215;
assign v3736af1 = hbusreq8_p & v3a635ea | !hbusreq8_p & v375aa99;
assign v3765c6d = hbusreq4 & v376f2f8 | !hbusreq4 & v8455ab;
assign v3a716a2 = hbusreq8 & v3773c13 | !hbusreq8 & v3767b5a;
assign v3a70879 = hmaster1_p & v3743ecf | !hmaster1_p & v8455ab;
assign v3a5b1ea = hbusreq4_p & v3747302 | !hbusreq4_p & v3a70b92;
assign v373ce66 = hbusreq8_p & v37299d5 | !hbusreq8_p & v1e37c44;
assign v377a6bf = hmaster0_p & v373c721 | !hmaster0_p & v3a64bc4;
assign v3760c1b = hmaster2_p & v3771ce2 | !hmaster2_p & v3a6ab5f;
assign v3772080 = hmaster0_p & v375121b | !hmaster0_p & v3740541;
assign v3a62eee = hmaster2_p & v3760881 | !hmaster2_p & v3a65762;
assign v3a699a1 = hbusreq6 & v3379037 | !hbusreq6 & v8455ab;
assign v37447df = hmaster2_p & v3a64349 | !hmaster2_p & !v374693f;
assign v375c4b0 = hbusreq5 & v35b9d58 | !hbusreq5 & v375b0ad;
assign v373c668 = hgrant0_p & v3808553 | !hgrant0_p & v3a65934;
assign v37495f2 = hlock2_p & v3731df6 | !hlock2_p & v374d173;
assign v37723a2 = hbusreq6_p & v37496b5 | !hbusreq6_p & !v8455ab;
assign v3a6a233 = hbusreq2 & v3a5a158 | !hbusreq2 & v3a62a6d;
assign v3a690ec = locked_p & v3a56346 | !locked_p & v8455ab;
assign v372a161 = hmaster2_p & v3a635ea | !hmaster2_p & v3a6efad;
assign v3a5397f = jx3_p & v3732ef8 | !jx3_p & v3a71392;
assign v3a713d8 = hbusreq0_p & v3766e3a | !hbusreq0_p & v3a70e52;
assign v376fc7f = hmaster1_p & v337905c | !hmaster1_p & v3a6fb0e;
assign v3a70040 = hmaster1_p & v3764761 | !hmaster1_p & v373aa0e;
assign v3a69547 = hmaster0_p & v375808f | !hmaster0_p & v3732d3e;
assign v374dd5f = hbusreq7_p & v3758c4d | !hbusreq7_p & !v3a704b8;
assign v3776633 = hmaster2_p & v3763a20 | !hmaster2_p & v3a6f8f5;
assign v3731be2 = hbusreq7 & v3a587dd | !hbusreq7 & v3a6f0c6;
assign v3750e4f = hbusreq7_p & v3771901 | !hbusreq7_p & !v3761916;
assign v3760b79 = hlock0 & v375da10 | !hlock0 & v375c0c4;
assign v3a672e6 = hmaster0_p & v3738a50 | !hmaster0_p & !v8455ab;
assign v3a7157b = hmaster2_p & v3a70641 | !hmaster2_p & v35772c9;
assign v37514f1 = hbusreq7 & v33790a4 | !hbusreq7 & v3732c96;
assign v37627bf = hbusreq6_p & v3a652a6 | !hbusreq6_p & v373e2db;
assign v3735331 = hbusreq5 & v37520d9 | !hbusreq5 & v8455ab;
assign v1e37b47 = hmaster2_p & v3a5a24b | !hmaster2_p & !v2ff8cfd;
assign v37777d5 = hmaster2_p & v3a61a7f | !hmaster2_p & v35b7092;
assign v3a70e25 = hmaster0_p & v1e382e7 | !hmaster0_p & v376fce9;
assign v372d417 = hmaster3_p & v377d9ab | !hmaster3_p & v3a6efdf;
assign v377d7bd = hmaster2_p & v3a6f781 | !hmaster2_p & v3775e81;
assign v376f576 = hmaster2_p & v3a703c3 | !hmaster2_p & !v37466cb;
assign v3a67b62 = hbusreq5_p & v3a6f051 | !hbusreq5_p & v3a5e000;
assign v3750613 = hlock6_p & v375d9f8 | !hlock6_p & v8455b3;
assign v377dee0 = hbusreq4_p & v3a707e9 | !hbusreq4_p & v373173e;
assign v375b258 = hmastlock_p & v2092f0a | !hmastlock_p & v8455ab;
assign v3755090 = hlock0 & v3a5741c | !hlock0 & v3a70a8f;
assign v3a6f2bb = hbusreq7_p & v375967d | !hbusreq7_p & v3733480;
assign v3768c19 = jx0_p & v373531a | !jx0_p & v3a7036b;
assign v377b0f7 = hbusreq0 & v3a70315 | !hbusreq0 & v372fa70;
assign v3743256 = hbusreq3_p & v376f860 | !hbusreq3_p & !v8455ab;
assign v3a6f335 = hmaster0_p & v3a6fad6 | !hmaster0_p & !v3725496;
assign v373ac12 = hlock4 & v377564e | !hlock4 & c2c2bc;
assign v3a671f4 = hburst0 & v3a5f308 | !hburst0 & v372f6a1;
assign v3774ccf = hmaster2_p & v377e089 | !hmaster2_p & !v372ee9a;
assign v3a6f6a9 = hmaster2_p & v3736d47 | !hmaster2_p & v3a70374;
assign v3728739 = hmaster2_p & v374b10b | !hmaster2_p & !v372c1a7;
assign v3766d0d = hbusreq2_p & v3a62986 | !hbusreq2_p & v3779e66;
assign v3a62229 = hmaster1_p & v3764494 | !hmaster1_p & v8455ab;
assign v3741dea = hmaster2_p & v3a6c8cc | !hmaster2_p & v3738251;
assign v3a681e8 = hmaster0_p & v3a7149d | !hmaster0_p & v2ff8c74;
assign v374952b = hbusreq8 & v3809ab5 | !hbusreq8 & v3a60276;
assign v3a6d806 = hgrant4_p & v3746806 | !hgrant4_p & !v3a623f2;
assign v37374e5 = hbusreq8 & v2acb0ef | !hbusreq8 & !v3773536;
assign v377b67d = hlock6 & v3a69efa | !hlock6 & v375b044;
assign v37635d6 = hlock8_p & v372f5e5 | !hlock8_p & v3a71096;
assign v375d92e = hmaster2_p & v8455bf | !hmaster2_p & v3a6f8f5;
assign v377497c = hgrant6_p & v3807f45 | !hgrant6_p & v372a831;
assign v3807abe = hmaster1_p & v3a5e24e | !hmaster1_p & v3734b14;
assign v3762c7c = hmaster0_p & v372a3de | !hmaster0_p & v3732931;
assign v3a6b31c = hgrant5_p & v3734ab5 | !hgrant5_p & v3a5a637;
assign v376653d = locked_p & v3762fc4 | !locked_p & v8455ab;
assign v373a0db = hbusreq5_p & v3a57ce9 | !hbusreq5_p & v3741627;
assign v3a71372 = hmaster0_p & v3a5f41b | !hmaster0_p & v372a2ae;
assign v372ab45 = jx0_p & v3731e5c | !jx0_p & v372bf72;
assign v37774ca = hmaster2_p & v3743b9e | !hmaster2_p & v3748d67;
assign v3a5fc9c = hbusreq8_p & v373fecb | !hbusreq8_p & v3a7042d;
assign v3a5b7b9 = hlock6 & v8716e3 | !hlock6 & v3a6e222;
assign v377672d = hmaster0_p & v8455ca | !hmaster0_p & v37327c5;
assign v373ff1c = hbusreq4 & v3a7024c | !hbusreq4 & v37450b8;
assign v3738832 = hmaster0_p & v3763175 | !hmaster0_p & v3a62841;
assign v375ce2d = hbusreq8_p & v3723698 | !hbusreq8_p & v37345a4;
assign v3744081 = hmaster0_p & v3742c9b | !hmaster0_p & v3a70bf8;
assign v3753f36 = jx0_p & v8455cd | !jx0_p & !v8455c9;
assign v9fa0b5 = hlock4 & v372fc07 | !hlock4 & v3a6fdb0;
assign v3730c3c = hmaster0_p & v3a71195 | !hmaster0_p & v372f151;
assign v377ec08 = hbusreq3 & v3a71452 | !hbusreq3 & v37496fa;
assign v3a6a758 = hbusreq5_p & v3740f7e | !hbusreq5_p & !v3a58cfc;
assign v373abdb = hbusreq6 & v3722f16 | !hbusreq6 & v375db62;
assign v3754eca = hmaster1_p & v3a6e581 | !hmaster1_p & v3a5ad83;
assign v377f66c = hbusreq7_p & v3765268 | !hbusreq7_p & v377074b;
assign v3a67ab9 = hbusreq3_p & v3750c92 | !hbusreq3_p & v8455ab;
assign v374693f = hbusreq0 & v3a645ca | !hbusreq0 & v8455ab;
assign v3a712a8 = hbusreq2 & v3776fa4 | !hbusreq2 & !v8455ab;
assign v3a709e1 = hbusreq4 & v8455ab | !hbusreq4 & v3737a76;
assign v3737ad2 = hgrant3_p & v8455bd | !hgrant3_p & v3725ccb;
assign v3736e19 = hmaster2_p & v3740161 | !hmaster2_p & v3727ad4;
assign v3a6fa58 = hmaster1_p & v37659c5 | !hmaster1_p & !v3a70f1e;
assign v3a713dd = hgrant6_p & v3778ed4 | !hgrant6_p & !v8455ab;
assign v376e717 = hgrant4_p & v377097a | !hgrant4_p & v3a6f801;
assign v3762ca6 = hmaster1_p & v3771076 | !hmaster1_p & v3a6fa2d;
assign v3758472 = hbusreq2_p & v8455e7 | !hbusreq2_p & !v8455ab;
assign v3734465 = hgrant3_p & v377dd3b | !hgrant3_p & v372faf1;
assign v375133a = hmaster1_p & v376b7e1 | !hmaster1_p & v373d245;
assign v3750e83 = hbusreq2 & v3a5f8d0 | !hbusreq2 & v8455ab;
assign v37572df = hbusreq6_p & v3733d6e | !hbusreq6_p & v372ee7e;
assign v3a5b0ea = hlock7_p & v3748f40 | !hlock7_p & v37788d6;
assign v3a5ad26 = hmaster2_p & v3747302 | !hmaster2_p & v3759f09;
assign v3a5ffac = hlock0 & v373bde3 | !hlock0 & v38078e5;
assign v376dfc9 = hmaster1_p & v3806a7b | !hmaster1_p & v3754e8c;
assign v3731fae = hmaster2_p & v374a343 | !hmaster2_p & v8455ab;
assign v3a7054a = hgrant6_p & v3a6f61e | !hgrant6_p & !v3a544db;
assign v374000d = hmaster2_p & v3a6297f | !hmaster2_p & v8b51d2;
assign v3a5dd60 = hmaster0_p & v3a5e24e | !hmaster0_p & v3752ee5;
assign v3809516 = hlock3 & v3a5cb68 | !hlock3 & v3809093;
assign v3741cc4 = hlock7 & v3a6ccc6 | !hlock7 & v3744657;
assign v3a6feb8 = hlock5_p & v374306c | !hlock5_p & v3a6ffae;
assign v37282c1 = hgrant6_p & v37484e0 | !hgrant6_p & v3748870;
assign v3744a0c = hgrant4_p & v37648af | !hgrant4_p & v373ce74;
assign v372d4d4 = hlock5_p & v3a5e3f1 | !hlock5_p & !v8455ab;
assign v3a65eba = hbusreq6_p & v3a70bb8 | !hbusreq6_p & v3734abe;
assign v3727ffa = hbusreq2 & v37275ef | !hbusreq2 & v3a5ab6e;
assign v3733170 = hbusreq4_p & v373512b | !hbusreq4_p & v3a658bf;
assign v3767578 = hgrant2_p & v3a709df | !hgrant2_p & v3739f1f;
assign v374b362 = hbusreq5 & v3a6eff8 | !hbusreq5 & v3754bc9;
assign v374bd7d = hgrant5_p & v374f307 | !hgrant5_p & v374314f;
assign v376ac47 = jx0_p & v3a65dbb | !jx0_p & v3a6fca0;
assign v374ab4f = hbusreq0 & v373e21a | !hbusreq0 & !v1e379fe;
assign v3730f34 = hbusreq7 & v37435b7 | !hbusreq7 & v8455b3;
assign v372eaaf = locked_p & v3a6c088 | !locked_p & !v8455ab;
assign v3a5ec1a = hmaster2_p & v37271e7 | !hmaster2_p & v8455ab;
assign v3a70dd8 = hmaster0_p & v3a57f59 | !hmaster0_p & v373d07a;
assign v3a59c87 = hbusreq6_p & v372c713 | !hbusreq6_p & v3a6f0d9;
assign v3a5ce0f = hmaster0_p & v3763f95 | !hmaster0_p & v373380d;
assign v38090e9 = hlock4_p & v8455ab | !hlock4_p & v3771ce2;
assign d9e97c = hbusreq5_p & v37494ed | !hbusreq5_p & v8455ab;
assign v372ff37 = hbusreq7_p & v37583ea | !hbusreq7_p & v3a71204;
assign v3737681 = hbusreq4 & v377221f | !hbusreq4 & v3755a05;
assign v3a675d9 = hmaster0_p & v3a5b28d | !hmaster0_p & v3a62e42;
assign v37bfc8a = hbusreq7 & v3779177 | !hbusreq7 & v377234d;
assign v3771cf0 = hbusreq4 & v3749907 | !hbusreq4 & v8455ab;
assign v377ba7d = hlock5_p & v3a57f59 | !hlock5_p & !v3a70c59;
assign v3726fff = hlock8_p & v3a663d6 | !hlock8_p & v3a6eb4e;
assign v372aafa = hlock8_p & v3a6e9fc | !hlock8_p & !v8455ab;
assign v3747704 = hgrant3_p & v3754877 | !hgrant3_p & v37485e0;
assign v3734579 = hmaster1_p & v3a5a510 | !hmaster1_p & v3a5ada9;
assign v375eeaf = hmaster1_p & v3a5b8b9 | !hmaster1_p & v3a70eeb;
assign v3774f45 = hbusreq1 & v376d9ad | !hbusreq1 & v8455e7;
assign v376b8e1 = hready_p & v3776225 | !hready_p & v3a70ca6;
assign v373ff8d = hready_p & v3742584 | !hready_p & !v8455ab;
assign v3a55844 = hbusreq2 & v37360b3 | !hbusreq2 & v8455ab;
assign v375f42e = jx0_p & v374eb9c | !jx0_p & v3a5dd98;
assign v372ce98 = hgrant4_p & v8455c1 | !hgrant4_p & v3725149;
assign v3743c45 = hmaster2_p & v8455e7 | !hmaster2_p & b0c091;
assign v3737808 = hmaster1_p & v8455ab | !hmaster1_p & v3a2a107;
assign v376bb9f = hgrant2_p & v8455ab | !hgrant2_p & !v3a71409;
assign v3a593e0 = stateG10_1_p & v3723430 | !stateG10_1_p & !v37598e6;
assign v3a6b53f = hgrant6_p & v3a6eb47 | !hgrant6_p & v3726f2e;
assign v3734a80 = hmaster1_p & v3a584d6 | !hmaster1_p & v372dd4b;
assign v33789d0 = hbusreq7 & v3723b33 | !hbusreq7 & v3743a4c;
assign v377a376 = hbusreq6_p & v3a5b7c2 | !hbusreq6_p & !v8455ab;
assign v3735749 = hmaster1_p & v373d703 | !hmaster1_p & v3748929;
assign v374e745 = hmaster0_p & v8455ab | !hmaster0_p & v8455e7;
assign v37402ee = hbusreq5_p & v3751887 | !hbusreq5_p & v3a709ae;
assign v375984e = hbusreq1 & v374e35e | !hbusreq1 & v8455ab;
assign v3a61ff4 = hmaster1_p & v3807754 | !hmaster1_p & v3a708c1;
assign v3744ada = hgrant4_p & v3746351 | !hgrant4_p & v3a6fd11;
assign v372e6d3 = hbusreq5 & v3a713a3 | !hbusreq5 & v39eb44a;
assign v3732bc0 = hbusreq2_p & v380749d | !hbusreq2_p & v372d59e;
assign v3779239 = hbusreq7_p & v3a5cb9d | !hbusreq7_p & !v372a1a9;
assign v380700f = hmaster3_p & v8455ab | !hmaster3_p & v3a715a2;
assign v3a62efa = hmaster2_p & v3a696a7 | !hmaster2_p & !v8455ab;
assign v3773df0 = hbusreq1 & v37757e0 | !hbusreq1 & v8455ab;
assign v37395bc = hgrant2_p & v3a5f50e | !hgrant2_p & !v8455ab;
assign v372d48a = hlock0 & v3809ec3 | !hlock0 & v37321c2;
assign v3760e6e = hmaster0_p & v3a57f59 | !hmaster0_p & v372ced7;
assign v3760a55 = hlock6 & v3753456 | !hlock6 & v3769bcb;
assign v3a691ea = hgrant5_p & v3a5cb95 | !hgrant5_p & v3378c5b;
assign v3772dd1 = hbusreq0_p & v3a670a1 | !hbusreq0_p & v3744265;
assign v3a5bb42 = hgrant4_p & v8455ab | !hgrant4_p & v3a70c95;
assign v373b286 = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a6fa72;
assign v373893a = hgrant4_p & v3752a0d | !hgrant4_p & v374572e;
assign v3774c25 = hmaster0_p & v3a661fe | !hmaster0_p & v3a70aae;
assign v3a70080 = hbusreq7 & v3a6edf6 | !hbusreq7 & cb8cbb;
assign v3731599 = hbusreq6 & v375301b | !hbusreq6 & v8455ab;
assign v3779324 = hbusreq1_p & v3a5c5ae | !hbusreq1_p & !v3a6368a;
assign v9e52e0 = hmaster2_p & v3a65b4a | !hmaster2_p & v8455ab;
assign v377c6ce = hbusreq0 & v3746ef3 | !hbusreq0 & v3760464;
assign v3a70336 = hlock4 & v3a6b70e | !hlock4 & v37659e2;
assign v37613bf = hmaster0_p & v3a58bb0 | !hmaster0_p & v3a6f541;
assign v39372da = hgrant5_p & v8455ab | !hgrant5_p & v372463a;
assign v3a6f08c = hbusreq5_p & v372a77f | !hbusreq5_p & v3a707a7;
assign v3750b5b = hmaster0_p & v375ad9f | !hmaster0_p & v3770a68;
assign v3a5a80c = hlock0_p & v372c3d4 | !hlock0_p & v3778f83;
assign v3a705d0 = jx0_p & af345a | !jx0_p & v3734632;
assign v3a70a3b = hbusreq0 & v37354b5 | !hbusreq0 & v3723400;
assign v3a645ac = hmaster0_p & v3a63ea7 | !hmaster0_p & v372ef80;
assign a6c8aa = hmaster1_p & v376ff3d | !hmaster1_p & v372661f;
assign v376ff64 = hmaster2_p & v3a5b1ea | !hmaster2_p & v3a5b6de;
assign v3a6f99d = hlock2_p & v3a6c1ac | !hlock2_p & v376430b;
assign v3751510 = hbusreq0 & v3a70aa2 | !hbusreq0 & v8455ab;
assign v37745b8 = hbusreq2_p & v3755a0f | !hbusreq2_p & v3743b9e;
assign v376eaf2 = hmaster2_p & v3a6f443 | !hmaster2_p & v3759032;
assign v3a6e8bc = hmaster0_p & v3a5bc35 | !hmaster0_p & v3750403;
assign v3a71602 = hmaster0_p & v374a277 | !hmaster0_p & v374e758;
assign d57388 = hlock6 & v3744d36 | !hlock6 & v3a702b5;
assign v3a653d5 = hbusreq8_p & v3745b5b | !hbusreq8_p & v376a6ae;
assign v3759c23 = hbusreq5 & v3743f7a | !hbusreq5 & v3a6f3f0;
assign v3764ec5 = hmaster2_p & v376a14f | !hmaster2_p & v3a70641;
assign v3a71356 = hmaster2_p & v8455ab | !hmaster2_p & v376c4f9;
assign v3a6fbe8 = hmaster0_p & v3a6dfb2 | !hmaster0_p & !v3779060;
assign v3a70512 = hgrant6_p & v91cdff | !hgrant6_p & v376b1bf;
assign v3777e69 = hgrant6_p & v3a62b8d | !hgrant6_p & v375f0ba;
assign v3a53da1 = hbusreq6_p & v37560f7 | !hbusreq6_p & v373ad95;
assign v37297ac = hmaster1_p & v3a7110d | !hmaster1_p & v8455ab;
assign v3a711bd = hmaster0_p & v37571c5 | !hmaster0_p & !v37c0294;
assign v3a71270 = hbusreq3_p & v376e41a | !hbusreq3_p & v374dfd9;
assign v37244a0 = hgrant2_p & v8455ab | !hgrant2_p & !v3729ffd;
assign v3a6de95 = hbusreq4 & v374cda0 | !hbusreq4 & v373bd6c;
assign v3a5d2f0 = hmaster2_p & v3746641 | !hmaster2_p & v3735ecd;
assign v373f911 = hgrant4_p & v8455ab | !hgrant4_p & v3a5dde7;
assign v3a6fcc8 = hlock6_p & v8455ab | !hlock6_p & !v1e379fe;
assign v3a7136b = hmaster0_p & v8455ab | !hmaster0_p & v3a71579;
assign v3766ff1 = hbusreq4_p & v375b9b2 | !hbusreq4_p & v375f3f4;
assign v3746bce = hmaster0_p & v3756ef4 | !hmaster0_p & v3746a7e;
assign v37353be = hgrant8_p & v3761f57 | !hgrant8_p & v3a6e733;
assign v377c3fb = hbusreq1_p & v360c6f5 | !hbusreq1_p & v3759c9c;
assign v375a10d = hbusreq4_p & v3a58218 | !hbusreq4_p & v3769cd3;
assign v3a5acd9 = hbusreq3 & v37482f8 | !hbusreq3 & !v3a709ea;
assign v39a4dc7 = hbusreq7 & v375ec51 | !hbusreq7 & v3a700d4;
assign v3761702 = hlock7_p & v374237b | !hlock7_p & v3777c7f;
assign v3a591b4 = hbusreq6_p & v3a70832 | !hbusreq6_p & v376a220;
assign v3728a4a = hbusreq8_p & v3763c1f | !hbusreq8_p & v37c36b9;
assign v3777386 = hgrant2_p & v3a6b873 | !hgrant2_p & v3a683d2;
assign v37751b4 = hlock7 & v3a70b10 | !hlock7 & v3731f35;
assign v3a70f26 = hgrant2_p & v37280c8 | !hgrant2_p & v374cf20;
assign v3a7022e = hgrant6_p & v8455ab | !hgrant6_p & v37520a9;
assign v377e864 = hbusreq4 & v3745f76 | !hbusreq4 & !v8455ab;
assign v3a6f54e = hmaster0_p & v3a66110 | !hmaster0_p & v3725d79;
assign v3730c26 = hgrant6_p & v8455ab | !hgrant6_p & v37602cf;
assign v374a86a = hbusreq6_p & v3732c72 | !hbusreq6_p & v3a6f90a;
assign v375d36b = hbusreq7_p & v3767d4a | !hbusreq7_p & v8455cb;
assign v3a6e222 = hlock2 & v3740dcd | !hlock2 & v37468ea;
assign v3746d2a = hbusreq6_p & v374249f | !hbusreq6_p & v8455ab;
assign v3a713f4 = hgrant2_p & v8455ab | !hgrant2_p & v3777d1f;
assign v376d892 = hgrant5_p & v3a7072e | !hgrant5_p & v3737ba0;
assign v374f028 = hbusreq0 & v374922a | !hbusreq0 & v1e37cd6;
assign v3a6fd54 = jx2_p & v3a60c59 | !jx2_p & v3a68f05;
assign v37332b8 = hbusreq8_p & v3a71294 | !hbusreq8_p & v3a5fcc2;
assign v376975e = hbusreq6_p & v377c7cf | !hbusreq6_p & v3766315;
assign v374801f = hmaster1_p & v3779183 | !hmaster1_p & v3a70501;
assign v3765d84 = hlock1_p & v3726aa5 | !hlock1_p & v3a63bb0;
assign v3763c39 = hmaster2_p & v3a7162d | !hmaster2_p & v8455ab;
assign v374fbca = hbusreq3 & v375f462 | !hbusreq3 & !v8455ab;
assign v3a71567 = hbusreq2 & v3763175 | !hbusreq2 & v8455ab;
assign v373bcdd = hlock5_p & v375bab8 | !hlock5_p & v8455ab;
assign v374b394 = busreq_p & v3577306 | !busreq_p & !v3a635ea;
assign v375408a = hlock2 & aebd68 | !hlock2 & v373413c;
assign v37498bd = hmaster2_p & v3739b80 | !hmaster2_p & !v3752fbc;
assign v3734312 = hbusreq1_p & v38071c1 | !hbusreq1_p & !v3a6f351;
assign v3741669 = hbusreq3_p & v37665ea | !hbusreq3_p & v35772a6;
assign v3a6f8d7 = hlock4 & v3a7138a | !hlock4 & v3a6af1d;
assign v3a5bc27 = hmaster1_p & v3755002 | !hmaster1_p & v3a6eb0e;
assign v3a552d4 = hbusreq2_p & v375b506 | !hbusreq2_p & v3740473;
assign v375d1d4 = hbusreq5_p & v3739938 | !hbusreq5_p & v374385c;
assign v3762f1a = hgrant6_p & v8455ab | !hgrant6_p & v3a714e8;
assign v3a712af = hbusreq0 & v37291ce | !hbusreq0 & !v3a6f744;
assign v3766e31 = hmaster0_p & d58c24 | !hmaster0_p & v3731bb5;
assign v3771c85 = hgrant4_p & v3736f61 | !hgrant4_p & v374a2f3;
assign v372e30c = hgrant6_p & v3a70f14 | !hgrant6_p & v3a64252;
assign v3771ee8 = hlock1_p & v3a5a0b3 | !hlock1_p & v374c4e1;
assign v3a67851 = stateA1_p & v8455e1 | !stateA1_p & v3768180;
assign v3a63da7 = hbusreq4 & v3777eed | !hbusreq4 & v372348c;
assign v376dc03 = hbusreq8 & v3a60815 | !hbusreq8 & v8455ab;
assign v3763b09 = hgrant7_p & v3a55fc1 | !hgrant7_p & v3751c00;
assign v3747d82 = hbusreq5 & v377c79a | !hbusreq5 & v375355c;
assign v3758d37 = hbusreq2_p & v37796f6 | !hbusreq2_p & v377002f;
assign a39369 = hgrant4_p & v8455ab | !hgrant4_p & v37515a6;
assign v3a6b368 = jx1_p & v3773881 | !jx1_p & !v372a478;
assign v377115c = hmaster3_p & v374fe65 | !hmaster3_p & v90a475;
assign v373fde1 = hmaster1_p & v3a5a6e6 | !hmaster1_p & v375f77f;
assign v3a630ba = stateG10_1_p & v3777ff7 | !stateG10_1_p & v374089e;
assign v372ac5c = hbusreq1_p & b4fa3c | !hbusreq1_p & v3807ddf;
assign v3a55bfa = hlock7 & v373b733 | !hlock7 & v37668b8;
assign v3a5edfe = hmaster1_p & v38074a8 | !hmaster1_p & !v375c7b9;
assign v3a69f0e = hmaster0_p & v3a70ec7 | !hmaster0_p & v3a6bc9a;
assign v3a58261 = hbusreq6_p & v39a5265 | !hbusreq6_p & v8455e1;
assign v3737d02 = hbusreq4_p & v3a71416 | !hbusreq4_p & !v3a6bc65;
assign v3751a9f = hbusreq4_p & v3726d1f | !hbusreq4_p & v3a6bb84;
assign v3773ff0 = hbusreq2_p & v8455bb | !hbusreq2_p & v8455b3;
assign v3a714e9 = hgrant2_p & v8455ab | !hgrant2_p & v3a5cc9d;
assign v3764910 = hmaster0_p & v3a635ea | !hmaster0_p & v3731dfe;
assign c6a502 = hgrant4_p & v37632f8 | !hgrant4_p & !v37243dc;
assign v3a573a7 = hmaster0_p & v375a10d | !hmaster0_p & v3727acb;
assign v372936a = hgrant6_p & v3a60576 | !hgrant6_p & v3a6f0e7;
assign a11f42 = hlock3_p & v372dbf1 | !hlock3_p & v23fdbca;
assign v373741d = hbusreq8 & v3773afc | !hbusreq8 & v3a6fb21;
assign v373b003 = stateA1_p & v3773a3d | !stateA1_p & v8455ab;
assign v3a661f3 = hbusreq5_p & v375897d | !hbusreq5_p & v3a5912f;
assign v373ba38 = hbusreq5_p & v3a66db2 | !hbusreq5_p & v3747ec9;
assign v955d7b = hmaster1_p & v3a6fa7a | !hmaster1_p & v37640e2;
assign v3a6f5e9 = hgrant5_p & v3a67af1 | !hgrant5_p & c0d797;
assign v377c6e8 = hbusreq2 & v37660d2 | !hbusreq2 & v3a635ea;
assign v376f501 = hgrant2_p & v3806c41 | !hgrant2_p & v3737209;
assign bd3213 = hbusreq3_p & v3748ae2 | !hbusreq3_p & v8455ab;
assign v3746e4e = hlock2_p & v8455ab | !hlock2_p & v35b70e6;
assign v38076a8 = hbusreq2_p & v3772020 | !hbusreq2_p & v37780f6;
assign v377baa6 = stateG10_1_p & v372c11d | !stateG10_1_p & !v3726570;
assign v374fefc = hmaster0_p & v373a822 | !hmaster0_p & v3738ed8;
assign v377225c = hbusreq7_p & v372b9a2 | !hbusreq7_p & v8455ab;
assign v37678e2 = hbusreq5 & v3a5af26 | !hbusreq5 & v3a5fc34;
assign v374dd24 = stateA1_p & v373f392 | !stateA1_p & !v3a7147e;
assign v372a04c = hbusreq4 & v3a5548b | !hbusreq4 & v3748797;
assign v372ba45 = hgrant6_p & v3a66e4c | !hgrant6_p & v3a5a211;
assign v380974c = hlock0_p & v3737554 | !hlock0_p & !v8455ab;
assign v375c70a = hbusreq5_p & v3a5b45b | !hbusreq5_p & v3770b26;
assign v3744640 = hbusreq6 & v376c2da | !hbusreq6 & v8455ab;
assign v375cb83 = hgrant6_p & v3a5cb45 | !hgrant6_p & v3737511;
assign v3748004 = jx0_p & v375dbb6 | !jx0_p & v373617a;
assign v3a5af28 = hbusreq0 & v3759f23 | !hbusreq0 & v3730d34;
assign v377e905 = hbusreq7 & v375cfaa | !hbusreq7 & !v3a6ff6e;
assign v3a6f1f2 = hbusreq6_p & v9cbad6 | !hbusreq6_p & v8455ab;
assign v3742033 = hbusreq2_p & v3743e29 | !hbusreq2_p & v8455b0;
assign v357732f = hbusreq1 & v3a70a12 | !hbusreq1 & v3a635ea;
assign ca2eb2 = hlock5 & v3761dda | !hlock5 & v376fbe3;
assign v3751861 = hmaster2_p & v3734967 | !hmaster2_p & v2092faa;
assign v1e37561 = hbusreq5_p & v3a6513d | !hbusreq5_p & v2925d06;
assign v376f09b = hlock5 & v372cd65 | !hlock5 & v3a57ebf;
assign v3a610e9 = hgrant1_p & v3a6ffae | !hgrant1_p & v3751fa8;
assign v3a68f4f = hbusreq6 & v3a710a2 | !hbusreq6 & v3a708c2;
assign v37629fc = hlock7 & v3734279 | !hlock7 & v377081e;
assign v3a70293 = hlock1_p & v37328bf | !hlock1_p & !v8455ab;
assign v37649a5 = hbusreq7 & v37273f4 | !hbusreq7 & v3a71167;
assign v376c5b4 = hmaster2_p & v3a70374 | !hmaster2_p & v3a71526;
assign v3774e8d = hbusreq5 & v3761a32 | !hbusreq5 & v8455ab;
assign v3a704e1 = hbusreq7_p & v37596f3 | !hbusreq7_p & v375e813;
assign v3a70a24 = hbusreq1 & v3748ca3 | !hbusreq1 & v373006f;
assign v3a6eb5c = hbusreq5 & v3735539 | !hbusreq5 & v3a5e030;
assign v37684c3 = hmaster2_p & v3a6e123 | !hmaster2_p & v3733471;
assign v3764ad1 = hbusreq4 & v376d2f4 | !hbusreq4 & v3737028;
assign v376eeea = hlock4_p & v8455ab | !hlock4_p & v373e21a;
assign v377bcfc = hmaster1_p & v3731d87 | !hmaster1_p & v376ca02;
assign v37277a5 = hgrant4_p & v37777ad | !hgrant4_p & v3a7092a;
assign v3a7065a = hgrant0_p & v8455ab | !hgrant0_p & !v3753233;
assign v3748ba4 = hlock4 & v374641d | !hlock4 & v3a70e5b;
assign v373cb58 = hbusreq6 & v3a71078 | !hbusreq6 & v37686f6;
assign v376dc15 = hbusreq2_p & v376cc8d | !hbusreq2_p & v3a5f5bb;
assign v37241db = hbusreq5_p & v37247b3 | !hbusreq5_p & v39eb5b0;
assign v37305cc = hgrant3_p & v3759512 | !hgrant3_p & !v3768264;
assign v3a70a7d = hbusreq0 & v3731b02 | !hbusreq0 & v8455ab;
assign v3a5d259 = hmaster2_p & v374d8ac | !hmaster2_p & v37287d8;
assign v372a0ed = hmaster0_p & v3747212 | !hmaster0_p & v3a6bc9a;
assign v372af06 = hbusreq5_p & v3774bad | !hbusreq5_p & v3a711e6;
assign v3a70ff1 = hlock4 & v37473ca | !hlock4 & v376a21e;
assign v3a70540 = hmaster0_p & v3a5d4ac | !hmaster0_p & v373c526;
assign v38069e7 = hmaster1_p & v3a64032 | !hmaster1_p & v8455c6;
assign v3774911 = hbusreq1 & v377989c | !hbusreq1 & v8455ab;
assign v375ceb9 = hgrant5_p & v3808e88 | !hgrant5_p & v3731e55;
assign v3a6a9d7 = hmaster2_p & v377489e | !hmaster2_p & v3257acb;
assign v3a62841 = hmaster2_p & v3763175 | !hmaster2_p & v3a6dc08;
assign v3a2ad1b = hbusreq4_p & v3755312 | !hbusreq4_p & v3743ef0;
assign v372a51d = hbusreq6_p & a3cddb | !hbusreq6_p & v3a5ffbf;
assign v37302fa = hmaster0_p & v8455ab | !hmaster0_p & v3a67d3d;
assign v3740c13 = hbusreq5_p & v3739589 | !hbusreq5_p & v37724b9;
assign v376f14f = hmaster1_p & v37255a1 | !hmaster1_p & !v8455ab;
assign v37629b0 = hbusreq5_p & v3725882 | !hbusreq5_p & v37315a3;
assign v372b9a2 = hlock7_p & v3a68825 | !hlock7_p & v3a6fb17;
assign v37543a0 = hbusreq4 & v3a61220 | !hbusreq4 & v3a6fee1;
assign v3a70efb = hlock8_p & v376230d | !hlock8_p & v8455ab;
assign v3764dc0 = hgrant4_p & v9ed516 | !hgrant4_p & v3a702e1;
assign v3a70f83 = hlock1_p & v373dd82 | !hlock1_p & v8455b0;
assign v3a6e66e = hgrant1_p & v8455ab | !hgrant1_p & !v3778ed4;
assign v3736c8c = hmaster1_p & v3577484 | !hmaster1_p & v3748929;
assign v372fff7 = hlock8_p & v37795eb | !hlock8_p & !v8455ab;
assign v3750b64 = hmaster1_p & v8455ab | !hmaster1_p & v3a7161c;
assign v3a70ab8 = hbusreq8_p & v3a708d8 | !hbusreq8_p & v375abaa;
assign v372c0de = hmaster1_p & c6fb51 | !hmaster1_p & v37793d4;
assign v372451b = hbusreq4_p & v373330f | !hbusreq4_p & v3757a57;
assign v3740ff7 = hbusreq8 & v3a6a367 | !hbusreq8 & v3a60276;
assign v3739646 = hmaster0_p & v3763f95 | !hmaster0_p & v37362e9;
assign v3748544 = hmaster0_p & v3a7147c | !hmaster0_p & v37243fe;
assign v37585d8 = hmaster2_p & v377c6dc | !hmaster2_p & v8455ab;
assign v3a7040e = hmaster0_p & v3758a92 | !hmaster0_p & v3a7090f;
assign v3a707e8 = hmaster1_p & v3758c15 | !hmaster1_p & v37258e7;
assign v376753a = hbusreq7_p & v3734200 | !hbusreq7_p & v374835b;
assign v3779910 = jx0_p & v374410c | !jx0_p & v39eb30a;
assign v3a70b7d = hmaster2_p & v8455ab | !hmaster2_p & v377e0b8;
assign v3756c19 = hbusreq8 & v377cb05 | !hbusreq8 & v3a715f8;
assign v3a7053b = hgrant6_p & v3a6b89e | !hgrant6_p & v3761224;
assign v3a5ebc8 = hmaster1_p & v3a6ffd3 | !hmaster1_p & v3a6f7b5;
assign v3a6bab9 = hgrant6_p & v8455ab | !hgrant6_p & v376a867;
assign v377a4ef = hmaster3_p & v375f106 | !hmaster3_p & v372814c;
assign v376a6f1 = hbusreq4_p & v8455ab | !hbusreq4_p & v1e37cd6;
assign v375a65f = hgrant6_p & v3a6f18f | !hgrant6_p & v372475e;
assign v3a6ff9e = hgrant4_p & v3a7133d | !hgrant4_p & v3a70204;
assign v376f536 = hbusreq7 & v374a0ab | !hbusreq7 & v3779f1e;
assign v3a6f847 = hbusreq7 & v3726e7b | !hbusreq7 & v3a7015b;
assign v3770fa1 = hmaster2_p & v375cde6 | !hmaster2_p & v3a70507;
assign v3758d7e = hbusreq0 & v374586b | !hbusreq0 & v3a6abcc;
assign v374b2f5 = hmaster0_p & v3a6f7dd | !hmaster0_p & v3a70941;
assign v377815b = hbusreq6_p & v373e748 | !hbusreq6_p & v3757b0e;
assign v3a70788 = hgrant2_p & v376ddfb | !hgrant2_p & v374047a;
assign v3a6ff9c = jx0_p & v37798bd | !jx0_p & v375043b;
assign v3a6c5fc = hgrant0_p & v38072fd | !hgrant0_p & v8455ab;
assign v376b1ad = hmaster0_p & v8455ab | !hmaster0_p & v37609a8;
assign v3a7145a = hgrant6_p & v3741f22 | !hgrant6_p & v3776a27;
assign v3756559 = hbusreq2_p & v374b724 | !hbusreq2_p & v8455ab;
assign v3a61be2 = hmaster2_p & v8455ab | !hmaster2_p & !v8455e1;
assign v3a5f371 = hbusreq6_p & v3a63545 | !hbusreq6_p & v8455ab;
assign v3a70c02 = hgrant2_p & v3758472 | !hgrant2_p & !v3a5eaa1;
assign v376fdb9 = hbusreq6 & v3777009 | !hbusreq6 & v37443ab;
assign v374b724 = hlock2_p & v3a70c96 | !hlock2_p & v3723f1a;
assign v3725673 = hmaster2_p & v3770e95 | !hmaster2_p & v3748d67;
assign v376f87a = hbusreq4 & v3730c26 | !hbusreq4 & v3a7164a;
assign v3735012 = hmaster2_p & v3a70209 | !hmaster2_p & v37771e3;
assign v37775f9 = hbusreq6_p & v3a635ea | !hbusreq6_p & v373cd68;
assign v3769ba9 = hbusreq4_p & v3a65bad | !hbusreq4_p & v3a6f817;
assign v372f235 = hmaster0_p & v3a6d81e | !hmaster0_p & v3732208;
assign v373031f = hgrant6_p & v38072fd | !hgrant6_p & v8455ab;
assign v375ff1e = jx0_p & v37702e6 | !jx0_p & !v8455ab;
assign v3723048 = hgrant6_p & v3a6dae2 | !hgrant6_p & v3a6f1ee;
assign v3a5b68a = hlock0_p & v39a537f | !hlock0_p & v3a7011c;
assign v3744794 = hlock2_p & v373c49e | !hlock2_p & v373929f;
assign v3a71340 = hmaster2_p & v3a7066c | !hmaster2_p & v35772a6;
assign v3a6ba08 = hbusreq5_p & v373ea09 | !hbusreq5_p & v373e873;
assign v3a6604e = hmaster2_p & v8455ab | !hmaster2_p & !v8455b6;
assign v3a5e60c = hmaster2_p & v37482f8 | !hmaster2_p & v3740df7;
assign v3752321 = hmaster0_p & v3a60229 | !hmaster0_p & v377ce5e;
assign v3a619c0 = busreq_p & v39a537f | !busreq_p & !v3a71084;
assign v377c35c = hmaster0_p & v3753418 | !hmaster0_p & v375fbae;
assign v3755026 = hbusreq2 & v3750859 | !hbusreq2 & v3a6ef1f;
assign v379318f = decide_p & v372cd7e | !decide_p & v3751a4f;
assign v377cb3d = hmaster1_p & v3a635ea | !hmaster1_p & v3a68315;
assign v3759cad = hmaster1_p & v3a6eb46 | !hmaster1_p & v3a6efb9;
assign v3a64af7 = hgrant6_p & v8455ab | !hgrant6_p & v380730d;
assign v374704e = hbusreq7 & v374ad23 | !hbusreq7 & v8455ab;
assign v3755dfa = hmaster3_p & v8455ab | !hmaster3_p & v375facd;
assign v3a647e7 = hlock8 & v372c345 | !hlock8 & v3a70f35;
assign v373c4e4 = hbusreq1 & v374362e | !hbusreq1 & v3a676d6;
assign v3743de1 = hgrant6_p & v3a62826 | !hgrant6_p & v3a6e699;
assign v3a5e2eb = hmaster0_p & v376c5b4 | !hmaster0_p & v3a70c2c;
assign v377c965 = hbusreq7 & v377981a | !hbusreq7 & v375bfc4;
assign v377911e = hgrant3_p & v9f7a48 | !hgrant3_p & !v375b203;
assign v3775d26 = hmaster2_p & v3a6f59d | !hmaster2_p & !v3777a00;
assign v375a9c1 = hmaster0_p & v8455ab | !hmaster0_p & !v3a6ab7f;
assign v3a6f88a = hbusreq7_p & v3a5dfa3 | !hbusreq7_p & v37240c0;
assign v3733a1a = hmaster2_p & v374a00a | !hmaster2_p & v3a7136e;
assign v3a53e45 = hmaster0_p & v380974c | !hmaster0_p & v3a6faf3;
assign v3a6ef91 = hmaster1_p & v3a70592 | !hmaster1_p & !v376acd9;
assign v376cc0e = hbusreq8_p & v3a7156b | !hbusreq8_p & v3a70646;
assign v38064a1 = hmaster3_p & v3a712b5 | !hmaster3_p & v3a5971d;
assign c98f7c = hgrant2_p & v3a5f50e | !hgrant2_p & v2acaf6f;
assign v3a6eb4e = hbusreq8 & v374e74c | !hbusreq8 & v3753838;
assign v37483db = hgrant3_p & v3a5b5d3 | !hgrant3_p & v37345f3;
assign v3722d9d = hbusreq4 & v37438b9 | !hbusreq4 & v3a5a807;
assign v37652cb = hbusreq0 & v3a7168b | !hbusreq0 & v3777da2;
assign v3a6fa9f = hgrant0_p & v3a6d6fe | !hgrant0_p & !v8455ab;
assign v3a6f5cd = hmaster0_p & v3a554d8 | !hmaster0_p & v374514c;
assign v374c9f0 = hbusreq2 & v3a67aaa | !hbusreq2 & v374f35a;
assign v3757e0b = hbusreq3 & v3726845 | !hbusreq3 & !v8455ab;
assign v37723b7 = hlock5 & v3762e54 | !hlock5 & v3a61724;
assign v3768e15 = hbusreq7_p & v3750d6d | !hbusreq7_p & v37703cb;
assign v9b63b0 = hmaster2_p & v3a637dd | !hmaster2_p & !v377f67b;
assign v3a6b27d = hlock5 & v3a70f09 | !hlock5 & v3a7161b;
assign v3a66cd7 = hmaster2_p & v37731ce | !hmaster2_p & v375a1ab;
assign v373cedb = jx1_p & v3a6f3b5 | !jx1_p & v3775da1;
assign v3a5be74 = hbusreq4_p & v3779283 | !hbusreq4_p & v8455ab;
assign v375dbb6 = hbusreq8_p & v3a63b69 | !hbusreq8_p & v3a70ed0;
assign v372abb9 = hmaster0_p & v3754a41 | !hmaster0_p & !v3a5c3d3;
assign v3764370 = hgrant6_p & v3772b34 | !hgrant6_p & !v3a57c2a;
assign v3a70c6c = hlock5 & v37596df | !hlock5 & v377d6fc;
assign v3a58102 = hgrant2_p & v8455ab | !hgrant2_p & v37731c3;
assign v373c703 = hgrant0_p & v3a70070 | !hgrant0_p & !v376ad4e;
assign v3a693b7 = hmaster2_p & v3a71026 | !hmaster2_p & v3a5bdd2;
assign v376f978 = stateA1_p & v8455ab | !stateA1_p & v3777a07;
assign v374a89b = hlock8 & v94b9e7 | !hlock8 & v37667d3;
assign v3a658d5 = hbusreq7_p & v3743def | !hbusreq7_p & v3a6724f;
assign v372ed5f = hmaster2_p & v374284d | !hmaster2_p & v8455ab;
assign v3758615 = locked_p & v375fed2 | !locked_p & v8455ab;
assign v376198e = hbusreq8 & v3774eec | !hbusreq8 & v3756a20;
assign v3a7014f = hbusreq8_p & v3737808 | !hbusreq8_p & v376f3ae;
assign v3a6f41c = hbusreq3_p & v3a70794 | !hbusreq3_p & v37447bf;
assign v3a714b7 = hmaster1_p & v3a5c945 | !hmaster1_p & v374d525;
assign v3758983 = hgrant2_p & v8455ab | !hgrant2_p & v3a6f6c6;
assign v376c1c3 = hbusreq5_p & v374a3b7 | !hbusreq5_p & v374d695;
assign v3727ff7 = hbusreq6_p & v374faa9 | !hbusreq6_p & v372f87c;
assign v3771931 = hmaster2_p & v3a703df | !hmaster2_p & !v3759158;
assign v3753404 = hlock7 & v374c9d9 | !hlock7 & v3a5c5e1;
assign v373f924 = hgrant6_p & v8455ca | !hgrant6_p & v3738c45;
assign v375c1d1 = hbusreq3_p & v8455bf | !hbusreq3_p & !v8455ab;
assign v3754a25 = hbusreq5_p & v8455c2 | !hbusreq5_p & v37358ab;
assign v375c6cc = jx1_p & v3755dfa | !jx1_p & v3a6d3c9;
assign v3a69584 = hlock4_p & v374306c | !hlock4_p & v3a6ffae;
assign v374b72f = hbusreq2_p & v3a5d28b | !hbusreq2_p & !v8455ab;
assign v3a711a8 = hmaster0_p & v37433e6 | !hmaster0_p & v8455ab;
assign v37676b8 = hbusreq2_p & v377286e | !hbusreq2_p & v8455b3;
assign v372c863 = hbusreq5 & v3a5ddaa | !hbusreq5 & v374ff15;
assign v3773666 = hmaster2_p & v3747302 | !hmaster2_p & v3745f9b;
assign v375987e = hbusreq6_p & v38072fd | !hbusreq6_p & v3746696;
assign beaea1 = hmaster2_p & v37c3782 | !hmaster2_p & v377d58d;
assign v3a71208 = stateG10_1_p & v377989c | !stateG10_1_p & v374c062;
assign v3a6fab6 = hmaster2_p & v1e3735b | !hmaster2_p & v8455ab;
assign v3744d54 = hmaster2_p & v3a62caa | !hmaster2_p & v3a709f2;
assign v3726339 = hmaster0_p & v372b9e9 | !hmaster0_p & v3774878;
assign v377af09 = hbusreq6_p & v3a5e7fe | !hbusreq6_p & v325b591;
assign v3a5b0b3 = hbusreq8 & v376c592 | !hbusreq8 & v3a6fa63;
assign v372438e = hbusreq5 & v3a67862 | !hbusreq5 & v3774bad;
assign v3a61b9d = hmaster1_p & v3a5e24e | !hmaster1_p & v374fdc9;
assign v3766462 = hmaster2_p & v375e854 | !hmaster2_p & v376bb26;
assign v3769093 = hbusreq4_p & v3a6589b | !hbusreq4_p & v8455ab;
assign v3a6836a = hbusreq5_p & v37384a9 | !hbusreq5_p & v374aa27;
assign v372b077 = hbusreq5_p & v376824b | !hbusreq5_p & v3778333;
assign v37556cb = hgrant0_p & v8455ab | !hgrant0_p & v37263bc;
assign v372846c = hbusreq3_p & v37361aa | !hbusreq3_p & v3a6816a;
assign v288971d = decide_p & v373ff8d | !decide_p & v372a7c2;
assign v37654bc = hbusreq8 & v3747280 | !hbusreq8 & v3a5e7bf;
assign v3a53e5c = hbusreq8 & v374fe7f | !hbusreq8 & v376f718;
assign v377ee33 = hbusreq2_p & v3779227 | !hbusreq2_p & v374d218;
assign v377d5d7 = hbusreq1_p & v37551f2 | !hbusreq1_p & bd3fa8;
assign v3735bdc = hgrant2_p & v3a682b1 | !hgrant2_p & v3a5a1ff;
assign v376219d = hmaster1_p & v3a70978 | !hmaster1_p & v3a6e0cc;
assign v23fd967 = hgrant2_p & v3a635ea | !hgrant2_p & v372d741;
assign v374096a = hgrant6_p & v3a71411 | !hgrant6_p & v3a5f5b3;
assign v3765f5c = hbusreq5 & v3758abd | !hbusreq5 & v3a57cc8;
assign v374fe7f = hmaster1_p & v8455e7 | !hmaster1_p & v3727f67;
assign v37238b1 = hlock6_p & v2acb5a2 | !hlock6_p & v8455ab;
assign v377744b = hbusreq0_p & v35772a5 | !hbusreq0_p & !v3a63621;
assign v3a67f13 = hmaster0_p & v3754685 | !hmaster0_p & v373c526;
assign v3754df4 = hbusreq0 & v3a5aaee | !hbusreq0 & v37298f1;
assign v375d889 = hmaster0_p & v3a70641 | !hmaster0_p & v376b86f;
assign v375ac6a = stateG10_1_p & v3806507 | !stateG10_1_p & v375a842;
assign v3760512 = hmaster2_p & v373997b | !hmaster2_p & v3a6773a;
assign v3a58a16 = hgrant3_p & v374383b | !hgrant3_p & v37584fe;
assign v374aca8 = hgrant2_p & v3a59bb4 | !hgrant2_p & v3a6f6fa;
assign v3739c66 = hmaster0_p & v37403fe | !hmaster0_p & v3747bfe;
assign v3770a1c = jx0_p & v373eea8 | !jx0_p & v37664aa;
assign d1f2e2 = hbusreq2_p & v37538e4 | !hbusreq2_p & v3743f47;
assign v3a6d1ea = hmaster0_p & v37536bf | !hmaster0_p & v3763e55;
assign v372ab8f = hbusreq4_p & v3a70f11 | !hbusreq4_p & v3a5c6e9;
assign v3a59dd6 = hmaster0_p & v3735b31 | !hmaster0_p & a97cd0;
assign v3a6f9d7 = hbusreq0 & v3741ccb | !hbusreq0 & v376efb6;
assign v3a64ad2 = hbusreq4 & v372a536 | !hbusreq4 & v8455ab;
assign v3a7006b = hgrant3_p & v3a56fcd | !hgrant3_p & !v3a6f342;
assign v37632c3 = jx1_p & a56488 | !jx1_p & v3808e9f;
assign v377d202 = hbusreq5_p & v377f78c | !hbusreq5_p & !v376b654;
assign v376b4d7 = hburst0 & v3a70cd5 | !hburst0 & v8455ab;
assign v377e4b4 = hmaster0_p & v376e431 | !hmaster0_p & v37341d3;
assign v372771e = hmaster0_p & v8455ab | !hmaster0_p & v37322a9;
assign v3773c62 = hlock4_p & v373fe5e | !hlock4_p & !v376430b;
assign v3a6f158 = hmaster0_p & v374fac7 | !hmaster0_p & v1e37cc1;
assign v372f95b = hgrant4_p & v3a6f65c | !hgrant4_p & v3a65856;
assign v3a6338d = hbusreq8_p & v375efe0 | !hbusreq8_p & v375a159;
assign v3a55eda = hmaster0_p & v375c791 | !hmaster0_p & v3a685db;
assign v3a6fcd2 = hmaster2_p & v3744b55 | !hmaster2_p & v3a5be93;
assign v3a6ca82 = hgrant3_p & v377dd3b | !hgrant3_p & v3a68a30;
assign v3a62403 = hbusreq5 & v3763364 | !hbusreq5 & v3730c96;
assign v376045b = hbusreq1 & v3723430 | !hbusreq1 & v8455ab;
assign v360d144 = hgrant5_p & v8455ab | !hgrant5_p & v373f684;
assign v3764955 = hbusreq8 & v3779c09 | !hbusreq8 & v1e37943;
assign v3a640d1 = hmaster0_p & v374f31d | !hmaster0_p & v3a715c5;
assign v3a5cccf = hbusreq4_p & v3a5ad1d | !hbusreq4_p & v3a5d841;
assign v374ac2c = hbusreq3_p & v3724d93 | !hbusreq3_p & v3a5903a;
assign v3a5f869 = hbusreq5_p & v3a6513d | !hbusreq5_p & v37554cd;
assign v372c92c = hbusreq5_p & v3a6de06 | !hbusreq5_p & v372c8d0;
assign v3a70b20 = hgrant5_p & v3a70955 | !hgrant5_p & v3736011;
assign v3738937 = hlock4 & v3a625c9 | !hlock4 & v3a5cb14;
assign v37724b9 = hmaster0_p & v3a53c18 | !hmaster0_p & v39eb565;
assign v3a70f66 = hmaster2_p & v3a64421 | !hmaster2_p & v3a70374;
assign v376acd5 = hgrant4_p & v8455ab | !hgrant4_p & v3a70bde;
assign v3a612fa = hmaster1_p & v3a606a0 | !hmaster1_p & v3a563c1;
assign v3a706a0 = hbusreq4_p & v37256d2 | !hbusreq4_p & v3761136;
assign v3a711cf = hbusreq7 & v3759c48 | !hbusreq7 & v3a6fe04;
assign v3a702c0 = hmaster2_p & v3744835 | !hmaster2_p & v3a6f99c;
assign v3735b31 = hmaster2_p & v3775eee | !hmaster2_p & v3747a41;
assign v373f2d8 = hgrant6_p & v3731e91 | !hgrant6_p & v3a6f8f9;
assign v373b1ae = hmaster2_p & v3738d63 | !hmaster2_p & v8455ab;
assign v372d744 = hbusreq4_p & v374ebe8 | !hbusreq4_p & v8455ab;
assign v3a6fec8 = hmaster2_p & v37640e9 | !hmaster2_p & v3a7142f;
assign v3729b75 = hmaster2_p & v3767cc9 | !hmaster2_p & v372d8f9;
assign v3755967 = hlock7_p & v374cc43 | !hlock7_p & v3a6199f;
assign v376563d = hbusreq1 & v3a619c0 | !hbusreq1 & !v8455ab;
assign v373b5f0 = hgrant2_p & v3a70823 | !hgrant2_p & v3730818;
assign v8cd321 = hlock5 & v3766b5a | !hlock5 & v3727981;
assign v3770db8 = hbusreq1 & v373b288 | !hbusreq1 & v3a635ea;
assign v375f98c = hgrant2_p & v3742033 | !hgrant2_p & v375d4f9;
assign v3747b78 = hbusreq8 & v3985142 | !hbusreq8 & v3734d58;
assign v3740a1e = hgrant5_p & v8455c6 | !hgrant5_p & v372f6ec;
assign v3741aa1 = hgrant2_p & v35b774b | !hgrant2_p & v375b974;
assign v377b9ab = hlock6_p & v3767f33 | !hlock6_p & v8455e7;
assign v3a70a04 = hgrant4_p & v3a6a0aa | !hgrant4_p & !v37584c6;
assign v3761cbb = hbusreq2_p & v37765e1 | !hbusreq2_p & v374d273;
assign v3a6f9a8 = hbusreq3 & v37453d8 | !hbusreq3 & v3773ee6;
assign v3a6f601 = hbusreq5_p & v377dca9 | !hbusreq5_p & v8455ab;
assign v374e828 = hbusreq7 & v376f7d1 | !hbusreq7 & v3768734;
assign v3a6dbaa = hbusreq0 & v380922b | !hbusreq0 & v3a71046;
assign v377bbd9 = hgrant4_p & v3779cf9 | !hgrant4_p & v3759361;
assign v374089d = hmaster2_p & v372a4c1 | !hmaster2_p & !v373dfff;
assign v373d7e9 = hmaster2_p & v375c791 | !hmaster2_p & v3a70374;
assign v3a6879a = jx0_p & v8455ab | !jx0_p & v373f364;
assign v3a6f7e9 = hmaster2_p & v376aa76 | !hmaster2_p & v373ae83;
assign v3a600b8 = hbusreq2 & v3746063 | !hbusreq2 & v374b3bf;
assign v374145b = hbusreq4 & v3a70bb7 | !hbusreq4 & v374165f;
assign v3a6fb6d = hmaster2_p & v376ac08 | !hmaster2_p & v37466cb;
assign a012c1 = hmaster2_p & v8455ab | !hmaster2_p & v3754d21;
assign v3a70769 = hmaster1_p & v374d6de | !hmaster1_p & v37246b5;
assign v3a70e68 = hgrant5_p & v3769323 | !hgrant5_p & v372351f;
assign d7cff8 = hmaster0_p & v8455ab | !hmaster0_p & v377f71d;
assign v372d0de = hbusreq6_p & v3a5ee3a | !hbusreq6_p & v372a4c3;
assign d7f8bb = hbusreq4 & v3746c51 | !hbusreq4 & v8455ab;
assign v3a701f3 = hbusreq8_p & v375035f | !hbusreq8_p & v37268b6;
assign v39eb550 = hbusreq5_p & v3a635ea | !hbusreq5_p & v377b3df;
assign v3742d60 = hlock1_p & v3775b81 | !hlock1_p & v8455ab;
assign v375c8c8 = hlock5 & v3a6678b | !hlock5 & v3740c5f;
assign v3a60c05 = hbusreq6_p & v3a6a78c | !hbusreq6_p & v3737534;
assign v3a70b72 = hbusreq0_p & v377217c | !hbusreq0_p & v3a6d8ce;
assign v3a70688 = hgrant3_p & v3735525 | !hgrant3_p & v376c343;
assign v3a70bea = hgrant6_p & v3a70dbe | !hgrant6_p & v376ab4e;
assign v376dcf6 = hlock7 & v3767b2e | !hlock7 & v375dd92;
assign v37371b2 = hbusreq4 & v376bea3 | !hbusreq4 & v3a641d5;
assign v376b11e = hbusreq0 & v3765219 | !hbusreq0 & v8fffa6;
assign v374ce71 = hbusreq0 & v3a7046b | !hbusreq0 & v373abde;
assign v37606f4 = hmaster0_p & v3753298 | !hmaster0_p & v3a705e6;
assign v3756ead = hbusreq5 & v373ebcf | !hbusreq5 & v37245a1;
assign v3a6f975 = hlock2_p & v377e2e2 | !hlock2_p & v3a66027;
assign v3766572 = hbusreq3_p & v3a70bd0 | !hbusreq3_p & v8455ab;
assign v3724882 = hmaster0_p & v3a62a6d | !hmaster0_p & v376e370;
assign v37769cc = hgrant4_p & v8455ab | !hgrant4_p & v3a577fe;
assign v3806d42 = hbusreq3 & v3723430 | !hbusreq3 & v8455ab;
assign v3753a65 = hmaster2_p & v376bcaa | !hmaster2_p & aab2b0;
assign v3a640ab = hbusreq6 & v3a70e10 | !hbusreq6 & v38072fd;
assign v376faf9 = jx1_p & v3a667ea | !jx1_p & v3779e21;
assign v37720ce = hmaster2_p & v372ae9d | !hmaster2_p & !v374e542;
assign v3a6fc3a = hmaster2_p & v372ee9a | !hmaster2_p & !v8455ab;
assign v376a27b = hgrant8_p & v8455ab | !hgrant8_p & v37274a2;
assign v372c221 = hgrant4_p & v3807f45 | !hgrant4_p & v377497c;
assign v373a391 = hburst1 & v372b0cd | !hburst1 & v3774074;
assign v3751dd2 = hbusreq5_p & v3749e4b | !hbusreq5_p & v372438e;
assign v3a6f6e2 = hmaster2_p & v3a635ea | !hmaster2_p & v3a68d2e;
assign v3a5bc35 = hmaster2_p & v3a637dd | !hmaster2_p & v2678c40;
assign v373edb9 = hmaster1_p & v375e50c | !hmaster1_p & v3775cca;
assign v373fa48 = hmaster0_p & v37681cc | !hmaster0_p & v8455ab;
assign v3a6fadc = hbusreq0 & v377349f | !hbusreq0 & v3769981;
assign v3a5f586 = hlock8 & v376ae9f | !hlock8 & v3763e46;
assign v3a70e49 = hmastlock_p & v37688a5 | !hmastlock_p & v8455ab;
assign v3771dc9 = hbusreq7_p & v3727a82 | !hbusreq7_p & !v8455ab;
assign v3a6f634 = hgrant5_p & v373b077 | !hgrant5_p & v375b9dc;
assign v3775a84 = hgrant0_p & v375f74a | !hgrant0_p & !v3757082;
assign v37758d0 = hmaster2_p & v8455ab | !hmaster2_p & !v3a715b0;
assign v3a5e90f = hgrant6_p & v8455ab | !hgrant6_p & v377433b;
assign v37794be = hburst0_p & v8455ab | !hburst0_p & v377f3af;
assign v376d33b = hmaster0_p & v3743ff2 | !hmaster0_p & v3a6f008;
assign v372ef62 = jx1_p & v380a20c | !jx1_p & v377b5aa;
assign v3a710d2 = hbusreq2 & v37406d2 | !hbusreq2 & v8455ab;
assign v376afc5 = hbusreq0 & v3744aed | !hbusreq0 & v375fed9;
assign v3731349 = hbusreq5_p & v372e36d | !hbusreq5_p & v3a70d63;
assign v374eac6 = hlock6 & v375b980 | !hlock6 & v375733e;
assign v3a5b91d = hgrant2_p & v8455ba | !hgrant2_p & v37749bf;
assign v3a678f9 = jx1_p & v3a5b78f | !jx1_p & v372ad29;
assign v3773100 = hbusreq1_p & v3a6fcc1 | !hbusreq1_p & !v3a70a60;
assign v3a5cd88 = hbusreq6 & v325b591 | !hbusreq6 & v37443ab;
assign v3a6f897 = hbusreq6 & v374282f | !hbusreq6 & v376fcc3;
assign v373e365 = hbusreq7_p & v37249fe | !hbusreq7_p & v3729520;
assign v376a3bb = hbusreq4 & v3a649fd | !hbusreq4 & v3a6a934;
assign v37464c8 = start_p & v3776483 | !start_p & v3730383;
assign v3a5f4e1 = hgrant2_p & v3757568 | !hgrant2_p & v3a5bead;
assign v374733b = hlock4 & v3730f35 | !hlock4 & v23fe101;
assign v374a99e = hbusreq4 & v3741022 | !hbusreq4 & v37c2b31;
assign v377b515 = hbusreq3 & v39a5350 | !hbusreq3 & v377ad8f;
assign v3756f06 = hbusreq4 & v373ee17 | !hbusreq4 & v8455ab;
assign v3a70c31 = hbusreq8_p & v3751849 | !hbusreq8_p & !v376dd7a;
assign v3a5bbed = stateG10_1_p & v375c196 | !stateG10_1_p & v372e6ad;
assign v37386d3 = hbusreq7_p & v3771533 | !hbusreq7_p & v3a5c842;
assign v3763076 = hmaster0_p & v3777301 | !hmaster0_p & v375daac;
assign v3760ba7 = hbusreq8 & v375580b | !hbusreq8 & v3a715f8;
assign v2ff8e1f = hlock0_p & v3a63e82 | !hlock0_p & !v35772a6;
assign v376fb07 = hlock7 & v3734279 | !hlock7 & v376ac10;
assign v377975f = hmaster0_p & v374306c | !hmaster0_p & c118e3;
assign v3a70342 = hgrant5_p & v3755066 | !hgrant5_p & v377af5d;
assign v3755f9a = hgrant6_p & v3747a53 | !hgrant6_p & v374a2be;
assign v3a70d01 = hbusreq0 & v3734bf8 | !hbusreq0 & v8455ab;
assign v372e1bc = hbusreq7_p & v375f2ab | !hbusreq7_p & v376ae39;
assign v3736f3b = hgrant2_p & v9ed516 | !hgrant2_p & v372e27f;
assign v3a6ff70 = hmaster1_p & v3a635ea | !hmaster1_p & v374c720;
assign v373dfbe = hbusreq3 & v37482f8 | !hbusreq3 & !v3a6fe6a;
assign v374fac6 = hgrant2_p & v3758fa7 | !hgrant2_p & v3766df9;
assign v3a5f21c = hbusreq4 & v8455c3 | !hbusreq4 & !v8455ab;
assign v3a71297 = hmaster0_p & v372b1b5 | !hmaster0_p & v374fe44;
assign v1e37846 = hbusreq4 & v37395e6 | !hbusreq4 & v8455e7;
assign v373b80b = hlock1_p & v374174c | !hlock1_p & !v8455ab;
assign v3a70c38 = hgrant0_p & v373b414 | !hgrant0_p & v3737462;
assign v3a6f551 = hbusreq8 & v3a595fd | !hbusreq8 & v3a6ec01;
assign v3a70497 = hbusreq8_p & v372a652 | !hbusreq8_p & v377329f;
assign v3a70d63 = hmaster0_p & v373505c | !hmaster0_p & v37509a9;
assign v374b4a4 = hgrant3_p & v3743b9e | !hgrant3_p & v37366d2;
assign v3a68591 = hbusreq2 & v37583be | !hbusreq2 & v376b4e1;
assign v3a5ce6f = hbusreq2_p & v3a6eb6b | !hbusreq2_p & v3761efb;
assign v377d652 = hmaster2_p & v8455ab | !hmaster2_p & v3739395;
assign v3a6d7f2 = hbusreq5_p & v3729f7b | !hbusreq5_p & v3a57046;
assign v3a7142a = hmaster0_p & v3a54c2e | !hmaster0_p & v3a59e1c;
assign v375e400 = hbusreq4_p & v3a6f856 | !hbusreq4_p & !v8455ab;
assign v3a6831c = hbusreq3_p & v3740409 | !hbusreq3_p & v8455ab;
assign v3807a32 = hbusreq4 & v374362e | !hbusreq4 & v3a676d6;
assign v3a6f4eb = hbusreq0 & v372c3a4 | !hbusreq0 & !v377d8b7;
assign v376501e = hbusreq4_p & v3741069 | !hbusreq4_p & v8455b0;
assign v37665ea = hlock3_p & v3722e5c | !hlock3_p & v35772a6;
assign v375ed63 = hbusreq0 & v372d366 | !hbusreq0 & v3727662;
assign v3774bed = hmaster1_p & v3769093 | !hmaster1_p & v375f41f;
assign d390f8 = hmaster0_p & v3a5865e | !hmaster0_p & v3a6fe27;
assign v3727bca = hbusreq6 & v3750613 | !hbusreq6 & v3a61445;
assign v3774494 = stateG10_1_p & v3a635ea | !stateG10_1_p & v376dc2e;
assign v3378c5b = hmaster1_p & v37432cd | !hmaster1_p & v3a5b20c;
assign v3a71387 = hlock0_p & v377eb2d | !hlock0_p & v8455b0;
assign v3a71249 = hbusreq5 & v37573f5 | !hbusreq5 & v3a6faae;
assign d70af8 = hlock0_p & v3748797 | !hlock0_p & v3a6212a;
assign v373bb90 = hbusreq0 & v373f058 | !hbusreq0 & v375d616;
assign v37237bc = hbusreq0_p & a38ed7 | !hbusreq0_p & v377b673;
assign v37380c4 = hgrant4_p & v37432c6 | !hgrant4_p & v372b1c8;
assign v31c3043 = hgrant5_p & v3770f97 | !hgrant5_p & v2ff9189;
assign v3a6f574 = hbusreq1 & v373c755 | !hbusreq1 & !v8455ab;
assign v37675e2 = hgrant0_p & v37773a9 | !hgrant0_p & v37376c8;
assign v3a689b8 = hgrant5_p & v8455ab | !hgrant5_p & v376ad46;
assign v373464d = hmaster2_p & v3a70374 | !hmaster2_p & v3746540;
assign v373b610 = hbusreq0 & v38073b0 | !hbusreq0 & v8455ab;
assign v3a67269 = hmaster0_p & v373418b | !hmaster0_p & v37628cd;
assign v3a667ea = hmaster3_p & v373ca17 | !hmaster3_p & v375edd8;
assign v3a6b0c7 = hbusreq3_p & v373be25 | !hbusreq3_p & !v372935c;
assign v3a56582 = hbusreq6 & v3a70e2e | !hbusreq6 & !v3a55033;
assign v3a71197 = hbusreq4 & v3742b84 | !hbusreq4 & v3748797;
assign v3777239 = hbusreq8 & v3774e48 | !hbusreq8 & v377c4d7;
assign v1e37c22 = hlock5_p & v3749f94 | !hlock5_p & v3a6546b;
assign v373ae27 = jx0_p & v374e207 | !jx0_p & v2092abf;
assign v376142c = hmaster2_p & v3739d88 | !hmaster2_p & v376a056;
assign v3755bb0 = hbusreq4 & v3731e7b | !hbusreq4 & v8455ab;
assign v3758f58 = hbusreq2 & v8455b0 | !hbusreq2 & v376648d;
assign v3759eb6 = hbusreq0 & v3765ef0 | !hbusreq0 & !v8455ab;
assign v922f0a = hgrant6_p & v8455ab | !hgrant6_p & !v3a6fb45;
assign v374a664 = hbusreq6_p & v8455e7 | !hbusreq6_p & !v8455ab;
assign v3734100 = hlock2 & v3767cfb | !hlock2 & v3742f4c;
assign v3a70cf0 = hbusreq6 & v37349ce | !hbusreq6 & v3a56e79;
assign v3a6fb52 = hmaster2_p & v373b7c5 | !hmaster2_p & v374ed52;
assign v375ee73 = hbusreq4_p & v3a59e5e | !hbusreq4_p & v8455ab;
assign v373d35d = hmaster0_p & v377ba41 | !hmaster0_p & v376a6f1;
assign v3a637ca = hgrant2_p & v8455ab | !hgrant2_p & v3a715e1;
assign v3736358 = hbusreq5_p & v23fde61 | !hbusreq5_p & v3a69a4c;
assign v37610ae = hbusreq5_p & v3765463 | !hbusreq5_p & v3a64612;
assign v3737415 = hmaster0_p & v360d036 | !hmaster0_p & v2925ce0;
assign v37390ba = hbusreq3 & v3a6eb01 | !hbusreq3 & v8455ab;
assign v37470fc = hmaster1_p & v3763f95 | !hmaster1_p & v3a5ce0f;
assign v3a6f462 = hmaster0_p & v3766da7 | !hmaster0_p & v372b7a3;
assign v37331c0 = hgrant6_p & v3a71164 | !hgrant6_p & v372d3e5;
assign v3a6c2b6 = hbusreq3_p & v8455ab | !hbusreq3_p & v8455b3;
assign v377bf2d = hbusreq6_p & v374faa9 | !hbusreq6_p & v372c500;
assign v3a6b9d9 = hlock8 & v3a611d8 | !hlock8 & v374c5f6;
assign v3a685cd = hready & v3a6bfea | !hready & v377eaf2;
assign v3725a73 = hmaster0_p & v3776d6e | !hmaster0_p & v374e288;
assign v3779b3a = hgrant5_p & v3a6e927 | !hgrant5_p & v377241f;
assign v374fba1 = hlock5 & v975066 | !hlock5 & v3759aca;
assign v3a715cb = hbusreq8 & v374d246 | !hbusreq8 & v3734279;
assign ce82b0 = hgrant2_p & v374a6fc | !hgrant2_p & v374056e;
assign v3a705a2 = hbusreq5_p & v3a672de | !hbusreq5_p & v3a672e6;
assign v376321e = hlock8 & v3a715ce | !hlock8 & v3a70426;
assign v3a64f96 = hlock7 & v377b205 | !hlock7 & v373e07e;
assign v3730f77 = hbusreq6_p & v8455ab | !hbusreq6_p & v375fd38;
assign v3724aaf = hlock6_p & v3a700ec | !hlock6_p & v3763668;
assign v376faf0 = hbusreq8 & v3a5fa45 | !hbusreq8 & v3a6e721;
assign v377b7ad = hlock6_p & v372b24d | !hlock6_p & v3a70131;
assign v3a6f7de = hgrant1_p & v377e8be | !hgrant1_p & !v35772a6;
assign v3a2a106 = hbusreq7 & v3a66bfa | !hbusreq7 & v3a635ea;
assign v3750b22 = hmaster2_p & v372abac | !hmaster2_p & v37647d8;
assign v3a6fe3d = hmaster0_p & v377348f | !hmaster0_p & v372700a;
assign v3769dcb = hgrant5_p & v8455c6 | !hgrant5_p & v3a6a7e8;
assign v3a6fcfd = hmaster2_p & v3a635ea | !hmaster2_p & v33789b9;
assign v376ab4e = hlock6 & v3a6c02f | !hlock6 & v3a583ee;
assign v3742b0e = hmastlock_p & v3722f37 | !hmastlock_p & !v8455ab;
assign v375f9df = hbusreq2_p & v3a635ea | !hbusreq2_p & v375cf36;
assign v374d260 = hbusreq1 & v3764463 | !hbusreq1 & v8455ab;
assign v3757537 = hbusreq5 & v3a53ed2 | !hbusreq5 & v380925f;
assign v377f384 = hburst0_p & v8455ab | !hburst0_p & v373db51;
assign v39eb4de = hbusreq3 & v376e568 | !hbusreq3 & v377437a;
assign v38063c7 = hgrant3_p & v3770559 | !hgrant3_p & v3775abc;
assign v3a60ef2 = hmaster3_p & v3734dc5 | !hmaster3_p & !v376b1ee;
assign v3771d77 = hlock3 & v372f8c1 | !hlock3 & v3a5f265;
assign v3739761 = hbusreq6_p & v377a9e7 | !hbusreq6_p & !v3747623;
assign v3734b6e = jx0_p & v2aca83b | !jx0_p & v8455ab;
assign v372bef3 = hbusreq5_p & v377a1dd | !hbusreq5_p & v3a6fb5a;
assign v3a6fd70 = hmaster1_p & v3a7159b | !hmaster1_p & !v377b6ce;
assign v9bf1d8 = hgrant4_p & v3a5fc34 | !hgrant4_p & v3a626e4;
assign v37294d3 = hbusreq0 & v39a537f | !hbusreq0 & v8455ab;
assign v3737075 = hgrant2_p & v8455ba | !hgrant2_p & v3a6106c;
assign v377f71d = hmaster2_p & v8455ab | !hmaster2_p & !v3a58261;
assign v3a587dd = hmaster1_p & v375d886 | !hmaster1_p & v3a66811;
assign v3763c59 = hmaster3_p & v3a68183 | !hmaster3_p & v3a60276;
assign v3a6eae9 = hmaster2_p & v3744b55 | !hmaster2_p & v3a65104;
assign v3739cfb = hmaster2_p & v3a635ea | !hmaster2_p & v3a6a374;
assign v3a70459 = hready & v3a63621 | !hready & v373b288;
assign v37646c7 = hbusreq2_p & v3748ca5 | !hbusreq2_p & v3752e65;
assign v376ffa7 = hgrant5_p & v372f4ce | !hgrant5_p & v3762640;
assign v3a539ae = hgrant4_p & v3a7018e | !hgrant4_p & v3a6f3ee;
assign v3a2978d = hbusreq6 & v372dd09 | !hbusreq6 & v8455ab;
assign v3740a9c = jx1_p & v376e966 | !jx1_p & v37683f8;
assign v3727dab = hmaster1_p & v3a7152b | !hmaster1_p & v3a70d30;
assign v372fe3d = hmaster1_p & v375025f | !hmaster1_p & v8455c9;
assign v37653a2 = hmaster0_p & v3747b29 | !hmaster0_p & v373e267;
assign v3a709c4 = hgrant3_p & v373efc2 | !hgrant3_p & v376c4fe;
assign v375d57e = jx1_p & v3a70e6e | !jx1_p & v2aca76c;
assign v3a6230b = hmaster2_p & v375b05e | !hmaster2_p & v3a6ff23;
assign v3732aca = hbusreq3 & v373aaa8 | !hbusreq3 & v8455ab;
assign v3a638aa = hmaster0_p & v98083e | !hmaster0_p & a7394c;
assign v377af11 = hlock5 & v374882c | !hlock5 & v3a5d678;
assign v377763c = hlock0 & v38078ed | !hlock0 & v3735c5a;
assign v375f99c = jx3_p & v3a549f5 | !jx3_p & v3a68d26;
assign v3a6ffc7 = hgrant4_p & v8455ab | !hgrant4_p & v1e37bf6;
assign v3727385 = hbusreq5 & v376fd32 | !hbusreq5 & v8455ab;
assign v3758233 = hgrant3_p & v374c937 | !hgrant3_p & v95d97e;
assign v3577354 = hgrant6_p & v8455ab | !hgrant6_p & v3a71393;
assign v3730f98 = hbusreq1_p & v3a6eb63 | !hbusreq1_p & !v373a2fc;
assign v3a5d929 = hmaster0_p & d0c237 | !hmaster0_p & v3752281;
assign v3a6106c = hgrant3_p & v8455be | !hgrant3_p & !c511c2;
assign v377cd6c = hlock4_p & v3a70327 | !hlock4_p & v374d402;
assign v374fd8d = hlock2_p & v3a70621 | !hlock2_p & v3a6ef74;
assign v373abd0 = hmaster0_p & v3a63ea7 | !hmaster0_p & v3773729;
assign v3a6fbb5 = hgrant5_p & v3a7131d | !hgrant5_p & !v3762f5b;
assign v3a6f1ea = hmaster0_p & v373c5a6 | !hmaster0_p & v374000d;
assign v376bcad = stateG2_p & v8455ab | !stateG2_p & v3751860;
assign v3745451 = hbusreq2 & v1e3755f | !hbusreq2 & v8455ab;
assign v3735809 = hbusreq3_p & v3771d77 | !hbusreq3_p & v3a5bb64;
assign v3772c7d = hbusreq4 & v373f058 | !hbusreq4 & v8455ab;
assign v3a5a41c = hlock3_p & v374b07a | !hlock3_p & v3a6fafa;
assign v9cc76d = hbusreq6_p & v3a70272 | !hbusreq6_p & !v3a5b68a;
assign v3a6d614 = hmaster2_p & v8455bf | !hmaster2_p & v3a6ac60;
assign v3a5c559 = stateG10_1_p & v3a539ee | !stateG10_1_p & v37526e0;
assign v374ba04 = hbusreq6 & v37719f2 | !hbusreq6 & v375cf36;
assign v373eeed = hbusreq7_p & v3a714b7 | !hbusreq7_p & v3a5b01c;
assign v3774653 = hbusreq4_p & v3a5bc04 | !hbusreq4_p & v35b724d;
assign v3a6ee50 = hmaster0_p & v375b429 | !hmaster0_p & v3a6f888;
assign v3a6f62c = hbusreq6 & v3a6d10a | !hbusreq6 & v391331d;
assign v3777c6d = hbusreq7_p & v3a56d3a | !hbusreq7_p & !v3746f4c;
assign v373b7b5 = hmaster0_p & v3740627 | !hmaster0_p & v8455ab;
assign v37310c2 = hgrant4_p & v377b6ce | !hgrant4_p & v37391e8;
assign v37658d7 = hbusreq6_p & v3764ac0 | !hbusreq6_p & v375492b;
assign v3a6f75e = hgrant6_p & v8455ca | !hgrant6_p & v37463ae;
assign v380987d = hmaster1_p & v3a71159 | !hmaster1_p & v3774399;
assign v372a2ff = hbusreq7 & v3a700ef | !hbusreq7 & v373abcf;
assign v376d66b = hmaster0_p & v3729a7a | !hmaster0_p & v2092ec6;
assign v3761adc = hgrant4_p & v3a71275 | !hgrant4_p & v35b7044;
assign v375aa99 = hlock8 & v3a716a2 | !hlock8 & v377c798;
assign v3773040 = hbusreq7_p & v8455cb | !hbusreq7_p & v3a6e675;
assign v3a707b1 = hmaster0_p & v8455b5 | !hmaster0_p & v3728202;
assign v3a700cd = hbusreq6 & v3a70200 | !hbusreq6 & !v3a5f89e;
assign v3a6adb8 = hlock8_p & v375722a | !hlock8_p & !v8455ab;
assign v3733c39 = hgrant0_p & v375da10 | !hgrant0_p & v374f35a;
assign v373f647 = hbusreq6_p & v3731eb5 | !hbusreq6_p & !v8455ab;
assign v376bf8a = hbusreq8_p & v3a70578 | !hbusreq8_p & v37274e6;
assign v3a5b0a6 = hbusreq5_p & v3742649 | !hbusreq5_p & v3a5cb2c;
assign v3736be1 = hbusreq4_p & v37294d3 | !hbusreq4_p & !v3723da9;
assign v3772608 = hgrant4_p & v8455ab | !hgrant4_p & v3a59548;
assign v37544cb = hlock4 & v373471f | !hlock4 & v2925d19;
assign v3a62329 = hbusreq2 & v373a27c | !hbusreq2 & v8455e7;
assign v376ca13 = hbusreq0 & v3378302 | !hbusreq0 & v377261b;
assign v3723b0c = hbusreq6_p & v3754aa3 | !hbusreq6_p & v375aaca;
assign v372c298 = hbusreq8 & v3a69ba1 | !hbusreq8 & v8455ab;
assign v3a6fbef = hbusreq2 & v374cab9 | !hbusreq2 & !v8455ab;
assign v3743f4d = hlock5_p & v3a6fb56 | !hlock5_p & v3750e0b;
assign v374e06f = hlock1 & v3a6d5b3 | !hlock1 & v37386a9;
assign v3a66822 = hbusreq0 & v3744a60 | !hbusreq0 & v373055c;
assign v3a6c022 = hgrant8_p & v3a6f548 | !hgrant8_p & v3a67c41;
assign v3a69ada = hgrant2_p & v3771137 | !hgrant2_p & v3751f28;
assign stateG3_2 = !v3a60ce2;
assign c4699e = hbusreq5_p & v37531fd | !hbusreq5_p & v3a70c04;
assign v3774a7d = hmaster0_p & v3a6672b | !hmaster0_p & v3a64bc8;
assign v37584e6 = hmaster2_p & v372bbd2 | !hmaster2_p & v3a6f329;
assign v375b233 = hlock4_p & v3a7153a | !hlock4_p & v373cc68;
assign v3a664e6 = hmaster1_p & v375ff00 | !hmaster1_p & v37698c3;
assign v3a64ba3 = hgrant5_p & v3a6e82d | !hgrant5_p & v372bbc7;
assign v3730c0a = hlock4 & v3a6f7ed | !hlock4 & v374829e;
assign v376ee82 = hmaster0_p & v3a71497 | !hmaster0_p & !v3739ea5;
assign v375d774 = hbusreq2 & v377109d | !hbusreq2 & v8455ab;
assign v3747c10 = hgrant6_p & v3735461 | !hgrant6_p & !v8455ab;
assign v37331b5 = hbusreq3 & v377af98 | !hbusreq3 & v8455ab;
assign v373db07 = hlock8_p & v3736ecc | !hlock8_p & v37758d3;
assign v376db9b = hmaster2_p & v375e60f | !hmaster2_p & v3728e09;
assign v3776445 = hbusreq7 & v3750700 | !hbusreq7 & v8455ab;
assign v375fd38 = hgrant2_p & v374fb58 | !hgrant2_p & v37758ce;
assign v3763191 = hlock0_p & v373997b | !hlock0_p & d3af9c;
assign v3a71057 = hmaster1_p & v37640e9 | !hmaster1_p & v377ea64;
assign v372ff96 = jx0_p & v374bfd6 | !jx0_p & v376e0cb;
assign v360d195 = hbusreq5 & v37522a0 | !hbusreq5 & v3a2a107;
assign v3753cf6 = hmaster0_p & v37782c9 | !hmaster0_p & v37396f7;
assign v2925d06 = hmaster0_p & v3a6fc3f | !hmaster0_p & v3a6f187;
assign aac06c = hmaster0_p & v8455ab | !hmaster0_p & v3a6f209;
assign v3a605e8 = hgrant0_p & v8455ab | !hgrant0_p & v3747dd0;
assign v375bd16 = hbusreq3 & v3a7151d | !hbusreq3 & !v8455ab;
assign v3725c63 = hbusreq6_p & v3768c3c | !hbusreq6_p & v3a70326;
assign v3738b70 = hmaster0_p & v3a6eb7e | !hmaster0_p & v37697ed;
assign v376a70f = hmaster3_p & v3a70ae5 | !hmaster3_p & v375d3da;
assign v3a70008 = jx1_p & v3a705b0 | !jx1_p & v376f98e;
assign v37339c8 = hbusreq4 & v3766025 | !hbusreq4 & v8455ab;
assign v3a60a2b = hmaster0_p & v8455ab | !hmaster0_p & !v3757740;
assign v3a6ebf6 = hlock0_p & v37416b5 | !hlock0_p & v3a70eff;
assign v3a6f547 = hgrant2_p & v3a71164 | !hgrant2_p & v376a898;
assign v3729e17 = hmaster0_p & v37656c1 | !hmaster0_p & !v374b1a4;
assign v3766f2e = hbusreq6_p & v3806e0e | !hbusreq6_p & v373c95b;
assign v377ae9c = hlock0_p & v373e67e | !hlock0_p & v3765cfd;
assign v3a7169e = hbusreq4 & v3765e46 | !hbusreq4 & v8455ab;
assign v3a7115d = hmaster0_p & v1e382e7 | !hmaster0_p & v3a6d33e;
assign v376c62d = hbusreq6 & v374d5c0 | !hbusreq6 & v8455ab;
assign v372eecf = hgrant3_p & v3779dae | !hgrant3_p & v377dfe2;
assign v3a55e3c = hmaster1_p & v376b438 | !hmaster1_p & v377b774;
assign v376648d = hbusreq3_p & v37406d2 | !hbusreq3_p & v8455b0;
assign v3764cea = hbusreq0 & v3a5f580 | !hbusreq0 & v3747ad6;
assign v37504eb = hbusreq4 & v3a676d6 | !hbusreq4 & v8455ab;
assign v3768c3e = hbusreq6_p & ae317f | !hbusreq6_p & !v8455ab;
assign v372ae0b = hgrant0_p & v37600af | !hgrant0_p & v3a70a68;
assign v3a6ae23 = hbusreq5 & v3a6b768 | !hbusreq5 & v3a5cb2c;
assign v3a6fd89 = hlock0 & v3749bf0 | !hlock0 & v3a6cc67;
assign v3a6c21d = hbusreq4_p & v376dbdf | !hbusreq4_p & !v372fc81;
assign v374af2f = hbusreq6 & v3a6e8d4 | !hbusreq6 & v373f492;
assign v37240c8 = hbusreq8_p & v372a8fd | !hbusreq8_p & v372db12;
assign v372ae1b = hgrant3_p & v8455ab | !hgrant3_p & v377b073;
assign v3745589 = hmaster2_p & v377d1dc | !hmaster2_p & v37763d1;
assign v37579ab = hbusreq4_p & v376f9eb | !hbusreq4_p & v8455ab;
assign v3a5c369 = hmaster2_p & v1e3735b | !hmaster2_p & v3770f75;
assign v3a5e3e2 = jx1_p & v3a7140d | !jx1_p & v3729f3c;
assign v377d4e1 = hbusreq5 & v3762a76 | !hbusreq5 & v377ee7c;
assign v3a71231 = hbusreq2_p & v3772117 | !hbusreq2_p & v3730b62;
assign v3770173 = hbusreq6_p & v3a70113 | !hbusreq6_p & v8455ab;
assign v3a67182 = hlock7_p & v3a6f7e4 | !hlock7_p & v3a5aff3;
assign v3746069 = hbusreq5_p & v3754d47 | !hbusreq5_p & v3a58c07;
assign v3a7019a = hbusreq4 & v375cf55 | !hbusreq4 & v38072fd;
assign v374ef97 = hbusreq8_p & v3762fd0 | !hbusreq8_p & v8455ab;
assign cfe9c3 = hbusreq6_p & v3743c51 | !hbusreq6_p & v3a63621;
assign v37229db = hmaster2_p & v3a6c23b | !hmaster2_p & v3749907;
assign v3a707c7 = hbusreq2_p & c58ea1 | !hbusreq2_p & v375bb6b;
assign v3a55162 = hmaster1_p & v3a711ee | !hmaster1_p & v37447e9;
assign v3a5cd6c = hlock6 & v3748797 | !hlock6 & v3729531;
assign v2ff918d = hmaster0_p & v376e2bb | !hmaster0_p & v8455ab;
assign v373384b = hgrant4_p & v3771697 | !hgrant4_p & v3a6a680;
assign v375b912 = hbusreq6_p & v3a70065 | !hbusreq6_p & v375d8ea;
assign v375abc2 = hmaster0_p & v3770f96 | !hmaster0_p & v3761c1a;
assign v3777d1f = hbusreq2_p & v372a960 | !hbusreq2_p & v3771e60;
assign v376e1ad = hmaster1_p & v37709d8 | !hmaster1_p & v376b27a;
assign v3a712ed = hmaster0_p & v3a70209 | !hmaster0_p & v3735012;
assign v3a7159b = hmaster0_p & v37750bb | !hmaster0_p & !v377b6ce;
assign v3a68b8a = hmaster0_p & v376501e | !hmaster0_p & v37273b1;
assign v3a66f07 = hgrant6_p & v3a645b0 | !hgrant6_p & v375c90b;
assign v3a56049 = hlock4_p & v3a6eb2b | !hlock4_p & v8455bf;
assign v372d28d = hbusreq7 & v3a5eefd | !hbusreq7 & v372d5e5;
assign v3a58d6b = hlock8 & v3a670e9 | !hlock8 & v373804d;
assign v376ff3d = hbusreq5_p & v373e12b | !hbusreq5_p & !v8455ab;
assign v377dae6 = hgrant3_p & v8455ab | !hgrant3_p & v3a647f3;
assign v3a6cad7 = hbusreq8_p & v3742fc4 | !hbusreq8_p & v377cd9c;
assign v3734b35 = hbusreq6 & v376d9ad | !hbusreq6 & v8455e7;
assign v3a6f477 = hlock4 & v374d965 | !hlock4 & v3725494;
assign v3772e46 = hlock6_p & v373ec0f | !hlock6_p & v3a6f5d1;
assign v3a70c1f = hbusreq4_p & v37250fa | !hbusreq4_p & v3a29810;
assign b0015f = hgrant5_p & v3a53d04 | !hgrant5_p & v376b220;
assign v376079f = hbusreq0 & v372d60f | !hbusreq0 & !v8455ab;
assign v3a549f0 = hbusreq7 & v3747b55 | !hbusreq7 & v37399ef;
assign v37288bc = hmaster2_p & v377ba59 | !hmaster2_p & v3a70e28;
assign v3744981 = hbusreq4_p & v39a537f | !hbusreq4_p & !v1e38224;
assign v3773c36 = hbusreq6_p & v373da8d | !hbusreq6_p & !v8455ab;
assign v3743d03 = hbusreq8 & v375a6d8 | !hbusreq8 & v8455ab;
assign v3a6d349 = hbusreq2_p & v3a6ff9b | !hbusreq2_p & !v3728eeb;
assign v3775c03 = hmaster2_p & v377b24b | !hmaster2_p & v35772b3;
assign v372b971 = hlock5_p & v3733384 | !hlock5_p & v8455ab;
assign v37232a6 = hlock4 & v3767c46 | !hlock4 & v3a6f567;
assign v372f6ce = hbusreq2 & v3a587bc | !hbusreq2 & v3771e60;
assign v3726f6b = hmaster2_p & v3a68084 | !hmaster2_p & !v8455ab;
assign v37291d1 = hbusreq2 & v373bff4 | !hbusreq2 & v377bb62;
assign v377d850 = hlock7_p & v3a542c0 | !hlock7_p & v3748301;
assign v3a70cfb = hbusreq3 & v3751734 | !hbusreq3 & v8455ab;
assign v3760765 = hmaster0_p & v3a703f2 | !hmaster0_p & v375d263;
assign v374586b = hlock4 & v3730052 | !hlock4 & v3a2a33d;
assign v3a56a79 = hbusreq5 & v3774103 | !hbusreq5 & v3776c87;
assign v37523ef = hbusreq5 & v372cdb0 | !hbusreq5 & v380925f;
assign v3a6380f = hmaster2_p & v376b4e1 | !hmaster2_p & !v3740df7;
assign v3a5a4ce = hbusreq7 & v37695e0 | !hbusreq7 & v8455ab;
assign v3730094 = hmaster1_p & v3a54466 | !hmaster1_p & v3a702fc;
assign v3751215 = hgrant2_p & v376495e | !hgrant2_p & v3a67904;
assign v376bfe6 = hmaster1_p & v3a67d66 | !hmaster1_p & v3778998;
assign v3a5c7a6 = hmaster0_p & v377bb3a | !hmaster0_p & v376dad7;
assign v3742ffc = hgrant7_p & v3a6fd35 | !hgrant7_p & !v3746cdd;
assign v373739c = hmaster2_p & v377adf5 | !hmaster2_p & !v3766bc8;
assign v3a63b57 = hbusreq4 & v35772a2 | !hbusreq4 & v8455ab;
assign v3749b46 = hgrant3_p & v8455ab | !hgrant3_p & v373f6c9;
assign v374a192 = hbusreq6 & v373997b | !hbusreq6 & v35b774b;
assign v3a656be = hbusreq5 & v3767797 | !hbusreq5 & v3a635ea;
assign v3a6ebea = hgrant5_p & v3a5fc34 | !hgrant5_p & v3a6f7e1;
assign v373621d = hgrant2_p & v374e5ac | !hgrant2_p & v372923a;
assign v37767cd = hbusreq4 & v372c007 | !hbusreq4 & !v8455ab;
assign v37513b7 = hgrant6_p & v377938d | !hgrant6_p & v3a64087;
assign v3a6f3ec = hmaster2_p & v8455ab | !hmaster2_p & !v3756925;
assign v3776fb2 = hbusreq4_p & v374304d | !hbusreq4_p & v372d967;
assign v3756971 = hgrant1_p & v3a7162d | !hgrant1_p & v8455ab;
assign v3a657bf = hbusreq6 & v3751734 | !hbusreq6 & !v8455ab;
assign v374ed4f = hgrant3_p & v3a71548 | !hgrant3_p & v3a5d04e;
assign v3a59bf7 = hbusreq8_p & v372bef4 | !hbusreq8_p & v375c4ef;
assign v3747c4c = hbusreq4_p & v3740f3d | !hbusreq4_p & v3a5db8a;
assign d60033 = hbusreq8_p & v375c7cb | !hbusreq8_p & v3777c6d;
assign v37758ad = hbusreq4_p & v3a7165b | !hbusreq4_p & v3758a02;
assign v3a5ee73 = hbusreq4_p & v3759b2f | !hbusreq4_p & v3a6f43e;
assign v375a2ff = hmaster0_p & v3a5acc7 | !hmaster0_p & !v3a713b7;
assign v3a714f5 = hlock0_p & v3a71452 | !hlock0_p & v3a5a647;
assign v373c059 = stateG10_1_p & v8455ab | !stateG10_1_p & v377e124;
assign v375cc1b = hbusreq4_p & v3a63a66 | !hbusreq4_p & v8455bb;
assign v3a6e8d4 = hgrant2_p & v8455ab | !hgrant2_p & v374a48c;
assign v3771555 = hmaster0_p & v3a6ff25 | !hmaster0_p & v375941a;
assign v3a70bd2 = hbusreq0_p & v37787ec | !hbusreq0_p & v3735512;
assign v376604d = hbusreq8 & v3734a93 | !hbusreq8 & v3a549f0;
assign v3a581e4 = hgrant6_p & v8455ca | !hgrant6_p & v3a6a2b5;
assign v3a7101d = hmaster0_p & v372757f | !hmaster0_p & v3a539bf;
assign v373ee3e = hmaster0_p & v3a712e2 | !hmaster0_p & v3a62092;
assign v3a70823 = hbusreq2_p & v3730818 | !hbusreq2_p & v3758e3c;
assign v376b1be = hgrant6_p & v377f397 | !hgrant6_p & v372bfbb;
assign v37235b8 = hmaster0_p & v377d1dc | !hmaster0_p & v3755289;
assign v3769921 = hgrant4_p & v3a70e7b | !hgrant4_p & !v8455ab;
assign v377d310 = hbusreq6 & v3a63ea7 | !hbusreq6 & v8455ab;
assign v3774b98 = hbusreq0 & v372cfd5 | !hbusreq0 & v3729b9f;
assign v3a54eae = hbusreq0 & v3a6ff8f | !hbusreq0 & v3779cb1;
assign v3730876 = hmaster2_p & v3a6e31f | !hmaster2_p & v3733e9e;
assign v3729f25 = hlock4_p & v3765e46 | !hlock4_p & !v8455ab;
assign v373ea7f = hmaster2_p & v8455b9 | !hmaster2_p & v376728e;
assign v3a7012a = hbusreq5_p & v374bace | !hbusreq5_p & v8455ab;
assign v3746211 = hmaster2_p & v8455ab | !hmaster2_p & v372fba5;
assign v372d92b = hmaster0_p & v3a6336e | !hmaster0_p & b2ea29;
assign v2092eaf = hlock2_p & v377e288 | !hlock2_p & v375eff3;
assign v3a5f47b = hbusreq8 & v3757ab6 | !hbusreq8 & v3a6ffb2;
assign v375b9c3 = hgrant3_p & v360d1cb | !hgrant3_p & v3725c02;
assign v3734a93 = hmaster1_p & v3a6e5f0 | !hmaster1_p & v3a70016;
assign v3a61e79 = hbusreq8 & v3a70daf | !hbusreq8 & v3778211;
assign v377ab6b = hmaster1_p & v9af7ec | !hmaster1_p & v3a70796;
assign v380956d = hbusreq0 & v3a6f378 | !hbusreq0 & v8455ab;
assign v3774608 = hmaster1_p & v8455bf | !hmaster1_p & v3a6fd1b;
assign b4f73f = hgrant2_p & v37672a5 | !hgrant2_p & v376a2bf;
assign v3a5ce54 = hmaster2_p & v3759031 | !hmaster2_p & v35772a2;
assign v3a675dc = hbusreq5 & v3a53b76 | !hbusreq5 & v8455ab;
assign v37249cc = hgrant4_p & v3729f14 | !hgrant4_p & v3764703;
assign v376ca9f = hmaster0_p & v3a58615 | !hmaster0_p & !v372fba0;
assign v3a63989 = hmaster2_p & v3a6dfb2 | !hmaster2_p & !v3a672c9;
assign v3a6ef77 = hbusreq8_p & v3a65587 | !hbusreq8_p & v376cf03;
assign v3a68289 = hbusreq5_p & v376d89f | !hbusreq5_p & v3a6dd1a;
assign v3778fec = hlock2 & v3767cfb | !hlock2 & v3771d77;
assign v37517f4 = hmaster2_p & v3a6890e | !hmaster2_p & v37425a5;
assign v3a55392 = hmaster2_p & v373014d | !hmaster2_p & v8455bf;
assign v374c0a4 = hmaster0_p & v375b429 | !hmaster0_p & v3a62d82;
assign v3a713c8 = hgrant6_p & v37445b9 | !hgrant6_p & v8455ab;
assign v3734d58 = hbusreq7 & v3a7157c | !hbusreq7 & v3a6a73d;
assign v3750674 = hlock6_p & v3a70bfa | !hlock6_p & v3773a45;
assign v375b261 = hbusreq2 & v29256bb | !hbusreq2 & v377c6b3;
assign v377a0a1 = hlock8_p & v376cff4 | !hlock8_p & v3747141;
assign v3a659b2 = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v3764881;
assign v3722bcf = hbusreq2_p & v3a6ff59 | !hbusreq2_p & v37313b6;
assign v3a71525 = hbusreq5 & v3748d2f | !hbusreq5 & v3a7107f;
assign dac24d = hmaster0_p & v3a60c38 | !hmaster0_p & v3779df7;
assign v3a2a33d = hgrant6_p & v8455ab | !hgrant6_p & v20930b8;
assign v3a70005 = hmaster1_p & v3734c40 | !hmaster1_p & v37568c9;
assign v3a708d4 = hbusreq5_p & v3a5aa5c | !hbusreq5_p & v3764dac;
assign v3725f77 = hlock0_p & v376d45f | !hlock0_p & v96020f;
assign v3a6da41 = hbusreq5_p & v3a5f6c3 | !hbusreq5_p & v3a7122f;
assign v3a6c555 = hbusreq8 & v3a6862e | !hbusreq8 & v3722af7;
assign v375c144 = hbusreq7 & v3808e88 | !hbusreq7 & a80fe2;
assign v3a64200 = hmaster1_p & v3a635ea | !hmaster1_p & v3761cd2;
assign v3775b82 = hgrant4_p & v372aacd | !hgrant4_p & v3a6f0ed;
assign v373bb89 = hbusreq8_p & v3a6adb8 | !hbusreq8_p & !v8455ab;
assign v376b1b7 = hmaster1_p & v377011b | !hmaster1_p & v3a704e3;
assign b85e8b = hbusreq7_p & v3723a2c | !hbusreq7_p & v376a74a;
assign v37365ce = hmaster2_p & v3737e2d | !hmaster2_p & v377f32e;
assign v372cf70 = hmaster0_p & v9f45ca | !hmaster0_p & v8455ab;
assign v374b5c5 = hgrant4_p & v3738636 | !hgrant4_p & v372367c;
assign v3a62a6d = hbusreq3_p & v375ea58 | !hbusreq3_p & v8455ab;
assign v376fa94 = hgrant6_p & v377f21b | !hgrant6_p & v372bcb0;
assign v3a7096d = hbusreq5 & v3809cc0 | !hbusreq5 & v8455ab;
assign v3807029 = hbusreq8 & v3a67d4f | !hbusreq8 & cb8cbb;
assign v3a5df94 = hbusreq0_p & v373f503 | !hbusreq0_p & v8455ab;
assign v3760912 = hgrant7_p & v3a62ef1 | !hgrant7_p & v3a710d1;
assign v3a692f6 = hmaster2_p & v23fe061 | !hmaster2_p & v35772a6;
assign v372d83d = hbusreq6 & v372d411 | !hbusreq6 & v3774175;
assign v3a5af5c = hbusreq4_p & v3a64ad6 | !hbusreq4_p & v8455ab;
assign v376f2fc = hbusreq5_p & v8455ab | !hbusreq5_p & v373f90a;
assign v3a70142 = hbusreq3_p & v375833e | !hbusreq3_p & v8455ab;
assign v37473af = hmaster2_p & v374362e | !hmaster2_p & v37395e6;
assign v3a5fe51 = hbusreq5_p & v3a5d438 | !hbusreq5_p & v3762079;
assign v37348ee = hbusreq0_p & v37457fb | !hbusreq0_p & v8455ab;
assign v3724543 = hbusreq6 & v37284f8 | !hbusreq6 & v8455ab;
assign v3776340 = hmaster2_p & v3a59c65 | !hmaster2_p & v37528d5;
assign v37709c5 = hgrant0_p & v3779647 | !hgrant0_p & !v8455ab;
assign v37790ef = hbusreq3_p & v375a4b3 | !hbusreq3_p & !v377b3a8;
assign v3736518 = hgrant8_p & v8455ab | !hgrant8_p & v3a6fca7;
assign v3a6eddd = hgrant6_p & v3763fb5 | !hgrant6_p & v374ed99;
assign v376e79d = hmaster0_p & v3a6f942 | !hmaster0_p & v3a6f073;
assign v3728625 = hbusreq4_p & v373506a | !hbusreq4_p & v3a6bb84;
assign v3766cf9 = stateG3_2_p & v8455ab | !stateG3_2_p & !v845603;
assign v37604fe = hbusreq5 & v3769982 | !hbusreq5 & v3a70cc8;
assign v3a6bba4 = hbusreq7 & v3a6fdf5 | !hbusreq7 & v3769a6c;
assign v3a62f05 = hgrant5_p & v8455ab | !hgrant5_p & v3a713b0;
assign v372cc01 = hmaster2_p & v373c3e1 | !hmaster2_p & !v3778e28;
assign v375b3b9 = jx0_p & v37c0339 | !jx0_p & v377b170;
assign v3a576d3 = hbusreq0 & v3755a84 | !hbusreq0 & v376b4a7;
assign v37559c4 = hmaster2_p & v373ee52 | !hmaster2_p & v377ad76;
assign v374ab4b = hmaster0_p & v373924d | !hmaster0_p & v37420bb;
assign v374d2dd = hgrant3_p & v3a6ffb6 | !hgrant3_p & v373ccb9;
assign v3766d11 = hgrant0_p & v37773a9 | !hgrant0_p & v3a6f1de;
assign v3a6980b = hmaster2_p & v3746b4f | !hmaster2_p & v373e2c3;
assign v374cc74 = hbusreq2_p & v374125a | !hbusreq2_p & v2092bae;
assign v376baef = hgrant2_p & v8455b9 | !hgrant2_p & v37272a8;
assign v37481e4 = hbusreq6_p & v375640f | !hbusreq6_p & !v372df2a;
assign v3768b2d = jx1_p & v376013c | !jx1_p & v372a7e7;
assign v374ca41 = hbusreq2_p & v3761c68 | !hbusreq2_p & v374ff44;
assign v376ae9c = hgrant6_p & v8455ab | !hgrant6_p & v3762c44;
assign v3a5f5bb = hgrant3_p & v3748797 | !hgrant3_p & v8455ab;
assign v374431a = hbusreq8_p & v3a696ee | !hbusreq8_p & v37628f6;
assign v3a67691 = hgrant6_p & v3a68f98 | !hgrant6_p & v3a70fd1;
assign v37568c8 = hlock1_p & v3769df4 | !hlock1_p & !v8455ab;
assign v377f70a = hbusreq4 & v3a6134b | !hbusreq4 & v3757009;
assign v377b24b = busreq_p & v3729480 | !busreq_p & v3724b72;
assign v1e38301 = hgrant5_p & v8455ab | !hgrant5_p & v3a6eb40;
assign v3768428 = hgrant0_p & v37773a9 | !hgrant0_p & v37457d1;
assign v374e849 = hbusreq4_p & v375b26a | !hbusreq4_p & v375a345;
assign v377d206 = hmaster2_p & v3577306 | !hmaster2_p & !v377b6ce;
assign v3773044 = hbusreq6_p & v3a6f92f | !hbusreq6_p & !v377adf5;
assign v3a5e030 = hmaster0_p & v374b0fb | !hmaster0_p & v3a66ab2;
assign v3736ae5 = hmaster1_p & v3753a34 | !hmaster1_p & v3a70cc7;
assign v3765f12 = hlock7 & b2d8a6 | !hlock7 & v3a6a8b2;
assign v3a6cc65 = hbusreq4_p & v3731b60 | !hbusreq4_p & !v8455ab;
assign v3a7152d = hmaster2_p & v3a68d0e | !hmaster2_p & v3a61cd7;
assign v3a627a1 = hmaster1_p & v8455ab | !hmaster1_p & v37431d8;
assign v3730766 = jx0_p & v3779e21 | !jx0_p & v3771dc9;
assign v3774063 = hmaster1_p & v2ff87a0 | !hmaster1_p & v3778628;
assign v375068a = hbusreq6 & v3a6bf60 | !hbusreq6 & v3729561;
assign v3a648a6 = hbusreq8 & v3a5b7e3 | !hbusreq8 & v3a635ea;
assign v377a9e2 = hbusreq5 & v3a70cf2 | !hbusreq5 & !v8455ab;
assign v37540dd = hmaster0_p & v3a7162f | !hmaster0_p & v3a59bbd;
assign v3a6f2cb = hbusreq0 & v3a5c25e | !hbusreq0 & v3a7137f;
assign v373ec0f = hgrant2_p & v3a5ff76 | !hgrant2_p & v3755b54;
assign v3771cf7 = hlock5 & v3734c47 | !hlock5 & v3a6f758;
assign v3a70e06 = hbusreq1 & v373fe5e | !hbusreq1 & v8455ab;
assign v37709d8 = hmaster0_p & v377d1dc | !hmaster0_p & v98083e;
assign v373fe10 = hbusreq0 & v3773a84 | !hbusreq0 & v8455ab;
assign v3a5dd86 = hbusreq4_p & v3748797 | !hbusreq4_p & v374bce0;
assign v37386c5 = hlock6_p & v3724940 | !hlock6_p & !v8455ab;
assign v374de73 = hmaster0_p & v3a6ff5b | !hmaster0_p & v3a71518;
assign v374355e = hbusreq0 & v3a5d469 | !hbusreq0 & v8455ab;
assign v3722b17 = hbusreq5_p & v37695c7 | !hbusreq5_p & v3a61336;
assign v37753e0 = hgrant6_p & v3757568 | !hgrant6_p & v3a5f4e1;
assign v376f53e = hmaster2_p & v3736847 | !hmaster2_p & v3732569;
assign v3773201 = hlock5_p & v37293c3 | !hlock5_p & !v8455ab;
assign v373540f = hmaster1_p & v3727d45 | !hmaster1_p & v37615d0;
assign v376725e = hbusreq4_p & v3a6fadc | !hbusreq4_p & v37666dd;
assign v3a70fc9 = hbusreq4 & v3a6fe44 | !hbusreq4 & v377bfc0;
assign v373185b = hmaster2_p & v37692c1 | !hmaster2_p & v3770719;
assign v376dbdf = hready & v373ff99 | !hready & v8455ab;
assign v3a6ad19 = hbusreq3 & v376129a | !hbusreq3 & v377ad8f;
assign v373fe61 = hgrant5_p & v8455ab | !hgrant5_p & v3735fd1;
assign v3807d51 = hbusreq7_p & v3a606b9 | !hbusreq7_p & v3a62cda;
assign v3a62037 = hbusreq3_p & v3a5ee99 | !hbusreq3_p & v3758c62;
assign v3745ee1 = hbusreq8 & v3a710f8 | !hbusreq8 & v37557c6;
assign v3a69ad1 = hmastlock_p & v37643ee | !hmastlock_p & !v8455ab;
assign v3a6f224 = hlock5 & v3748cd9 | !hlock5 & v3769f4e;
assign v38092f5 = hmaster1_p & v3738253 | !hmaster1_p & v377a2e1;
assign v8b32e5 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3743f9a;
assign v377d33e = hbusreq0_p & v37787ec | !hbusreq0_p & v3a6c0b3;
assign v373951e = hlock8_p & v3742e25 | !hlock8_p & v8455ab;
assign v3777149 = hmaster2_p & v3a672c9 | !hmaster2_p & !v3728e09;
assign v377297e = hbusreq6_p & v3777ee9 | !hbusreq6_p & !v8455ab;
assign v3a70e6e = hmaster3_p & v3a5b40f | !hmaster3_p & v3806e5b;
assign v376480b = hmaster0_p & v3a6b07b | !hmaster0_p & !v37628cd;
assign v375f462 = hlock0_p & v3a6fe6a | !hlock0_p & v375ecc7;
assign v3742ed3 = hgrant8_p & v8455c5 | !hgrant8_p & v376e5ef;
assign v376752b = hmaster2_p & v3a69de7 | !hmaster2_p & v3747302;
assign v3a70909 = hmaster2_p & v3753418 | !hmaster2_p & v3a705f2;
assign v3146177 = hgrant2_p & v8455ab | !hgrant2_p & v8455b9;
assign v376856b = hbusreq0 & v372c91d | !hbusreq0 & v8455ab;
assign v3a563cf = hlock5 & v37790a6 | !hlock5 & v372f0bc;
assign v38093a8 = hlock5_p & v3768695 | !hlock5_p & v8455ab;
assign v375d1ae = hbusreq4 & v3771ab9 | !hbusreq4 & v3a68f98;
assign v3737511 = hbusreq6_p & v373e09c | !hbusreq6_p & v94e000;
assign adf78a = hlock3_p & v8455b0 | !hlock3_p & !v8455ab;
assign v373c3a0 = hmaster2_p & v37690f3 | !hmaster2_p & v374243d;
assign v3a55959 = hgrant4_p & v8455ab | !hgrant4_p & v3765eee;
assign v374d8ea = hmaster2_p & v3a6ef5a | !hmaster2_p & v37447e9;
assign v3a6ff31 = hmaster0_p & v3736104 | !hmaster0_p & v3a61c70;
assign v37234d1 = hmaster2_p & v377adf5 | !hmaster2_p & !v3a56cdb;
assign v3257acb = hbusreq0 & v3a61580 | !hbusreq0 & v376a0fc;
assign v374c900 = hgrant4_p & v8455ab | !hgrant4_p & v374503d;
assign c45930 = hmaster0_p & v3724394 | !hmaster0_p & v375e099;
assign v3743038 = jx1_p & v372e49a | !jx1_p & v3763c59;
assign v3a6f8f9 = hbusreq3_p & v37367da | !hbusreq3_p & !v8455ab;
assign v3764f48 = hmaster2_p & v3a62a6d | !hmaster2_p & v3a5e544;
assign v375f689 = hmaster1_p & v3a63de8 | !hmaster1_p & v3a6fc50;
assign v3a70ac2 = hmaster2_p & v8455ab | !hmaster2_p & !v3a6f742;
assign v3770ab9 = hbusreq6_p & v377c3ea | !hbusreq6_p & v3a6fe8e;
assign v3a6fa28 = hgrant2_p & v3a5eadd | !hgrant2_p & v376d82f;
assign v3760ef5 = stateG2_p & v8455ab | !stateG2_p & v3a5fcfc;
assign v3a70c98 = hmaster2_p & v20d166d | !hmaster2_p & v8455ab;
assign v373ed57 = hbusreq5_p & v3a6d2ed | !hbusreq5_p & v3a55ea1;
assign v3746feb = hlock2_p & v376725a | !hlock2_p & v3748645;
assign v3731579 = hbusreq8 & v375d5e1 | !hbusreq8 & v3741b61;
assign v377af48 = hbusreq8_p & v3a5d834 | !hbusreq8_p & v3a5dcd4;
assign v377fc51 = hbusreq5 & v374e843 | !hbusreq5 & v376072e;
assign v3773a9d = hbusreq1_p & v3a711f0 | !hbusreq1_p & !v8455ab;
assign v3753231 = hmaster1_p & v375d434 | !hmaster1_p & v3757a04;
assign v3722ba9 = hbusreq8_p & v3a716a4 | !hbusreq8_p & v3a53709;
assign v3a703db = hmaster2_p & v3a5c945 | !hmaster2_p & v3733e9e;
assign v3730b6c = hgrant4_p & v8455ab | !hgrant4_p & v3728a77;
assign v3a6fe5e = hmaster2_p & v3745181 | !hmaster2_p & v3740f5d;
assign v3754ec0 = hbusreq6 & v3768ef1 | !hbusreq6 & v376bade;
assign v372c11d = locked_p & v3a5e24e | !locked_p & v3807bf8;
assign v3728a76 = hlock0 & v38073c9 | !hlock0 & v3a70532;
assign v3767d14 = hlock0 & v375f9df | !hlock0 & v3736bcd;
assign v23fdbce = hlock7_p & v3a66e63 | !hlock7_p & !v8455ab;
assign v3a7032d = hbusreq3 & v3a5f8d0 | !hbusreq3 & v8455ab;
assign v37451c0 = hlock8_p & v3a66d74 | !hlock8_p & v376b829;
assign v3777da5 = hmaster2_p & v37590d1 | !hmaster2_p & v3a6d622;
assign v374a580 = hbusreq4_p & v3a5794d | !hbusreq4_p & v35772a6;
assign v3a5f447 = hgrant5_p & v3a70c1d | !hgrant5_p & v375b99c;
assign v3735e89 = hlock4 & v376ee80 | !hlock4 & v376ebbf;
assign v373bee7 = hbusreq5_p & v374743d | !hbusreq5_p & v372707d;
assign v3a5ad17 = hbusreq5 & v374cbe2 | !hbusreq5 & v373790d;
assign v3a66671 = hbusreq2_p & v3765b28 | !hbusreq2_p & !v375e8a2;
assign v377c31d = hgrant6_p & v8455ab | !hgrant6_p & v3a55349;
assign v3729280 = hlock0 & v377e8da | !hlock0 & v376c1e4;
assign v372ad52 = hgrant2_p & v38095ed | !hgrant2_p & v37424b5;
assign v3731eb8 = hbusreq3 & v374e35e | !hbusreq3 & v8455ab;
assign v375e33e = hgrant5_p & v3a57733 | !hgrant5_p & v3a6fcb5;
assign v3a5faaa = hbusreq6_p & v373261a | !hbusreq6_p & v3a6b80e;
assign v3770c96 = hbusreq4 & v8455b0 | !hbusreq4 & v3730ffe;
assign v3747035 = hgrant3_p & v377b6ce | !hgrant3_p & v3729c37;
assign v3a63e82 = stateA1_p & v375956a | !stateA1_p & !v3732170;
assign v3732849 = hmaster1_p & v3a70298 | !hmaster1_p & v373a3c3;
assign v3778901 = hgrant5_p & v8455ab | !hgrant5_p & v3a7027a;
assign v375ea88 = hgrant5_p & v8455ab | !hgrant5_p & v3777da6;
assign v372a1d6 = hgrant4_p & v3730e2a | !hgrant4_p & v3731d89;
assign v3742abe = hmaster2_p & v372433d | !hmaster2_p & v3a6f7a2;
assign v375a5f9 = hmaster0_p & v372d8e8 | !hmaster0_p & a3d29c;
assign v373c65b = hgrant6_p & v8455ca | !hgrant6_p & v376c630;
assign v375d17c = hmaster0_p & v373f42d | !hmaster0_p & v3757966;
assign v3a5ab08 = hbusreq5_p & v37480b3 | !hbusreq5_p & v3a6ef2c;
assign v373da59 = hmaster2_p & v3750c50 | !hmaster2_p & v8455ab;
assign v372416d = hbusreq5 & v38069c8 | !hbusreq5 & v3736a50;
assign v37413d5 = hgrant2_p & v37320bb | !hgrant2_p & v3a62654;
assign v37436a8 = hgrant2_p & v8455ab | !hgrant2_p & v3a703b9;
assign v375afc1 = hbusreq2_p & v3748797 | !hbusreq2_p & v3a64f05;
assign v372debd = hgrant7_p & v8455c9 | !hgrant7_p & v37530d1;
assign v3724579 = hgrant5_p & v8455ab | !hgrant5_p & v3757966;
assign v3a6f945 = hmaster1_p & v376b662 | !hmaster1_p & v37469ba;
assign v3a6f989 = hgrant3_p & v3759032 | !hgrant3_p & v3747eef;
assign v3a70613 = hbusreq5 & v3a6fb7f | !hbusreq5 & v3772e85;
assign v3a66529 = hgrant5_p & v3a6b078 | !hgrant5_p & v3809464;
assign v3a53e30 = hbusreq5_p & v374b393 | !hbusreq5_p & v8455ab;
assign v3738e62 = hbusreq5 & a0715f | !hbusreq5 & !v8455ab;
assign v3760bdd = hbusreq4_p & v3a59b8a | !hbusreq4_p & v3728399;
assign v376c644 = hgrant4_p & v8455ab | !hgrant4_p & v3a711e7;
assign v373f058 = hlock2_p & v8455b0 | !hlock2_p & !v8455ab;
assign v377b218 = hbusreq2_p & v374f12d | !hbusreq2_p & v376aa6d;
assign v3775831 = hlock4 & v3775144 | !hlock4 & v3730bf9;
assign v3773cda = hmaster0_p & v3750b9d | !hmaster0_p & v37584e6;
assign v376b70a = hgrant5_p & v8455ab | !hgrant5_p & !v3a70b57;
assign v3a563d3 = hbusreq6 & v37677a3 | !hbusreq6 & v8455ab;
assign v1e37e1f = hbusreq7_p & v3740766 | !hbusreq7_p & !v3767e03;
assign v373867a = hlock8 & v3a6fb6a | !hlock8 & v3a6f0f3;
assign v374650c = hmaster2_p & v8455ab | !hmaster2_p & v377d0fc;
assign v3768a43 = hbusreq7 & v376ed58 | !hbusreq7 & v374312f;
assign v39a4ca6 = hmaster1_p & v3766d4b | !hmaster1_p & v3734d9a;
assign v3a6d32c = hgrant6_p & v373351d | !hgrant6_p & !v8455ab;
assign v3768304 = hlock0 & v3a70a7f | !hlock0 & v3757695;
assign v3a6f407 = hmaster3_p & v376ae9f | !hmaster3_p & v8455ab;
assign v3a6ebcd = hgrant4_p & v3739896 | !hgrant4_p & v374f677;
assign v37784a9 = hlock8_p & v3a6fc5c | !hlock8_p & v3a70623;
assign v372dcfb = hmaster2_p & v376dc26 | !hmaster2_p & v3a7058a;
assign v3a6f328 = hgrant6_p & v374a664 | !hgrant6_p & v3a5b4c1;
assign v3751161 = hbusreq3 & v3777baa | !hbusreq3 & v8455ab;
assign v3a70b4c = hmaster3_p & v376130f | !hmaster3_p & v3a5edfe;
assign v3a70176 = hlock8_p & v3725ca4 | !hlock8_p & v3a63f6d;
assign v373d3ec = hlock5_p & v3756263 | !hlock5_p & v377bae8;
assign v3744710 = hbusreq0_p & v8455ab | !hbusreq0_p & v8455b5;
assign v376d268 = hgrant4_p & c8ab71 | !hgrant4_p & v3739e25;
assign v3758a9c = hbusreq4 & v372e4de | !hbusreq4 & v38073c9;
assign v372842d = hgrant0_p & v37496fa | !hgrant0_p & v375fbd7;
assign v3723c0d = hlock3 & v376d34b | !hlock3 & v372e169;
assign v37294c5 = hmaster1_p & v3a56b92 | !hmaster1_p & v375b9b0;
assign v375c999 = hbusreq7_p & v375f3cf | !hbusreq7_p & v3733664;
assign v375d2cf = hlock8_p & v3a705bd | !hlock8_p & v377444f;
assign v374c9ee = hbusreq0_p & v8455ab | !hbusreq0_p & !v373ad95;
assign v377419d = hlock2_p & v8455ab | !hlock2_p & v8455e7;
assign v377800b = hmaster1_p & v3750fc9 | !hmaster1_p & c46b05;
assign v3a6fdec = hmaster1_p & v3a637dc | !hmaster1_p & v2ff87c6;
assign v374de0d = hmaster2_p & v375b2e2 | !hmaster2_p & v37514c7;
assign v3a55198 = hbusreq0 & v374021a | !hbusreq0 & v3743adf;
assign v3a713fb = hlock0_p & v3a5b5d3 | !hlock0_p & v3a658bf;
assign v3751dba = hmaster2_p & v3a635ea | !hmaster2_p & v3a70410;
assign v372f5c5 = hbusreq7 & v37385d3 | !hbusreq7 & v374c790;
assign v372c1a7 = hgrant4_p & v375c7b9 | !hgrant4_p & v372f12d;
assign v372b7a8 = hmaster2_p & v3a696a7 | !hmaster2_p & v3a637dd;
assign v3a5da8f = hmaster2_p & v3a5a807 | !hmaster2_p & v376ac08;
assign v37387ed = hbusreq6 & v3a6ffca | !hbusreq6 & v8455ab;
assign v3a6f36e = hbusreq3_p & v375bc6e | !hbusreq3_p & v3728ca9;
assign v3a6f93a = hgrant4_p & v37300a5 | !hgrant4_p & v3746dc9;
assign v374764e = hmaster0_p & v3a7066c | !hmaster0_p & v3a5c16e;
assign v3a70607 = hgrant1_p & v8455ab | !hgrant1_p & v37547c9;
assign v3a63383 = hbusreq8_p & cc70ad | !hbusreq8_p & v377c348;
assign v3761953 = hbusreq7 & v3a7088a | !hbusreq7 & v3a70b3f;
assign v376b141 = hlock2_p & v377b774 | !hlock2_p & v8455bf;
assign v37480fe = hgrant6_p & v3a7083b | !hgrant6_p & v374429f;
assign v9af7ec = hbusreq4_p & v374db8d | !hbusreq4_p & !v8455ab;
assign v3a6a693 = hmaster0_p & v3a713c3 | !hmaster0_p & v3758c72;
assign v3a65b42 = hmaster0_p & v376b044 | !hmaster0_p & v3a7090f;
assign v374af92 = hlock4_p & v374d057 | !hlock4_p & v3a702c2;
assign v3a71333 = hmaster1_p & v3724f4f | !hmaster1_p & v3577318;
assign v3a6ec30 = hmaster2_p & v8455ab | !hmaster2_p & v8455b0;
assign v3a6f6f1 = hmaster1_p & v3a70fd5 | !hmaster1_p & d3ed45;
assign v3a563af = hgrant4_p & v3751d73 | !hgrant4_p & v3a7105c;
assign v3a5d99f = hlock7 & v3a70bc4 | !hlock7 & v37735ba;
assign v3a66151 = hbusreq1_p & v3a69a06 | !hbusreq1_p & v373d0e1;
assign v3a563ba = hlock2_p & v377362f | !hlock2_p & !v8455ab;
assign v3a6f316 = hgrant1_p & v8455ab | !hgrant1_p & v3775b81;
assign v3776f8c = hbusreq6_p & v3a6324b | !hbusreq6_p & v37443ab;
assign v3755cf7 = hbusreq5 & v372c483 | !hbusreq5 & v3a62a6d;
assign v373cd03 = hmaster2_p & v3a70374 | !hmaster2_p & v3730986;
assign b3b89e = hmaster1_p & v37289f0 | !hmaster1_p & v3a708f4;
assign v376f641 = jx0_p & v376bf8a | !jx0_p & v3757a61;
assign v3a70070 = hlock0_p & v3735e39 | !hlock0_p & v3a70964;
assign d5ffe1 = hlock4 & v3a71615 | !hlock4 & v3748de3;
assign v376f920 = hlock5_p & v3768da7 | !hlock5_p & v373eadd;
assign c80162 = hgrant5_p & v37621c1 | !hgrant5_p & v3a70b90;
assign v37476c2 = hlock5 & v2ff8e74 | !hlock5 & v3745202;
assign v3754a39 = hmaster0_p & v3728164 | !hmaster0_p & v8455ab;
assign v3a70c2e = hbusreq0 & v3765f13 | !hbusreq0 & v3809ec3;
assign v3a5c858 = hbusreq6_p & v3735f02 | !hbusreq6_p & v3a70b66;
assign v37621ea = hbusreq2_p & v3a635ea | !hbusreq2_p & v376eaca;
assign v374dabc = hlock7 & v3a6f25b | !hlock7 & v3a7159f;
assign v3776bdf = hmaster0_p & v377504a | !hmaster0_p & v373d076;
assign v374dcbd = hmaster0_p & v3a70ded | !hmaster0_p & v3731079;
assign v3a70077 = hmaster0_p & v376db9b | !hmaster0_p & !v37243fe;
assign v374bfc8 = hbusreq2_p & v377144d | !hbusreq2_p & v3758f58;
assign v376a2d6 = hmaster2_p & v3767437 | !hmaster2_p & v374b3cf;
assign v3733e04 = hbusreq8 & v3736d3a | !hbusreq8 & v3735f30;
assign v3a5f1e8 = hmaster0_p & v374502e | !hmaster0_p & v374908e;
assign v3a6830c = stateG10_1_p & v35772a5 | !stateG10_1_p & !v3806507;
assign v37535fd = hmaster1_p & v37790c8 | !hmaster1_p & v3a70859;
assign v373c379 = hmaster0_p & v377adf5 | !hmaster0_p & !v99aa13;
assign v3767ed6 = hbusreq3 & v3a5600a | !hbusreq3 & v37757e0;
assign v9204d4 = hmaster0_p & v3736d47 | !hmaster0_p & v3747edc;
assign v3750295 = hready_p & v3a6fd54 | !hready_p & v2093068;
assign v375a9d0 = hgrant4_p & v374a950 | !hgrant4_p & v3a56318;
assign v3742d6c = hmaster1_p & v37737aa | !hmaster1_p & v377cf20;
assign v3a69dd2 = hbusreq8_p & v372b1e8 | !hbusreq8_p & v3736382;
assign v37652d7 = hlock8_p & v377974f | !hlock8_p & v3a5e74c;
assign v3778ac2 = hmaster0_p & v3a6fb6d | !hmaster0_p & v374c164;
assign v3a6f0c6 = hmaster1_p & v3753f1d | !hmaster1_p & v372c28d;
assign v3765433 = hlock7 & v372d3f1 | !hlock7 & v3a6ff70;
assign v373568b = hmaster0_p & v376db9c | !hmaster0_p & v374d339;
assign v3a705e2 = hmaster2_p & v373e6d2 | !hmaster2_p & v374f5e0;
assign v3a5eae2 = hmaster0_p & v3757f54 | !hmaster0_p & v3a59bbd;
assign v3759b09 = hlock5_p & v3a6810b | !hlock5_p & v3738726;
assign v3775782 = hmaster2_p & v3a62a6d | !hmaster2_p & v37453d7;
assign v3a6f20f = hbusreq6_p & v376d9aa | !hbusreq6_p & v373b288;
assign v375cf55 = hbusreq6_p & v373f7b7 | !hbusreq6_p & v38072fd;
assign a26fed = hmaster2_p & v374b5a8 | !hmaster2_p & v376d374;
assign v3a5e65e = hmaster3_p & v3a5f0f0 | !hmaster3_p & v8455ab;
assign v23fe175 = hlock4 & v3731685 | !hlock4 & v376c87d;
assign v3767261 = hmaster1_p & v3a6fdc0 | !hmaster1_p & v8455ab;
assign v3a66f83 = hbusreq3_p & d44200 | !hbusreq3_p & !v3a7151d;
assign v3734965 = hmaster3_p & v3a6843e | !hmaster3_p & v376a7bf;
assign v374710b = hbusreq1_p & v375104f | !hbusreq1_p & v3745dba;
assign v374b274 = hlock4 & v3745c75 | !hlock4 & v376dcca;
assign v37c2b31 = hlock4_p & v3724940 | !hlock4_p & !v8455ab;
assign v375e1f6 = jx1_p & v374b237 | !jx1_p & !v3725be8;
assign v3a6f81d = hgrant2_p & v3758472 | !hgrant2_p & !v3a5cf3d;
assign v372989c = hgrant3_p & v377a42f | !hgrant3_p & v372b6c4;
assign v3a5a225 = stateG2_p & v8455ab | !stateG2_p & !v373e80b;
assign v376e441 = hbusreq5_p & v3746818 | !hbusreq5_p & v38072fe;
assign v3807a7d = hbusreq8 & v3736a59 | !hbusreq8 & v3a704ef;
assign v377a0f2 = hbusreq8_p & v3a713bb | !hbusreq8_p & v3a56f2d;
assign v376fb6b = hgrant6_p & v3737571 | !hgrant6_p & v376b3bc;
assign v374581a = hmaster2_p & v3a64421 | !hmaster2_p & v3a6fc7f;
assign v377aa23 = hlock2 & v3749b37 | !hlock2 & v3731ffc;
assign c60044 = hlock1_p & v3a63af6 | !hlock1_p & !v377c2ac;
assign v37637d4 = hmaster0_p & v8455ab | !hmaster0_p & v3a6e91e;
assign v3750ea5 = hmaster2_p & v8455ab | !hmaster2_p & v37648af;
assign v37c039c = hbusreq6_p & v3a636d9 | !hbusreq6_p & v3731172;
assign v3a6f7a6 = hlock8_p & v3a5724f | !hlock8_p & !v8455d2;
assign v3a56593 = hgrant2_p & v377a42f | !hgrant2_p & v372989c;
assign v3776fc5 = hbusreq5 & v3746dbf | !hbusreq5 & v3771c85;
assign v377e419 = hgrant4_p & v8455ab | !hgrant4_p & v375e262;
assign v3a706e3 = hmaster2_p & v374e531 | !hmaster2_p & v3a609bb;
assign v3734d12 = hgrant6_p & v8455ca | !hgrant6_p & v3723ded;
assign v3a6d7a0 = hmaster1_p & v3725de9 | !hmaster1_p & v3a70516;
assign v373ade9 = hbusreq4_p & v3758166 | !hbusreq4_p & !v3a56e63;
assign v3a65afd = hmaster1_p & v3a57801 | !hmaster1_p & v3a70cc7;
assign v373badc = hbusreq4_p & v373997b | !hbusreq4_p & v37738fc;
assign v2ff8bbc = hbusreq4_p & v3723fcc | !hbusreq4_p & v373b288;
assign v377c079 = hlock4 & v3762656 | !hlock4 & v376f23f;
assign v3731684 = hbusreq5_p & v3a6f4e3 | !hbusreq5_p & v3775e7e;
assign v37467e9 = hmaster1_p & v375e50c | !hmaster1_p & c98bc3;
assign v3a71405 = hmaster0_p & v3807f45 | !hmaster0_p & v3727e33;
assign v3a68821 = hbusreq5_p & v372ec65 | !hbusreq5_p & v3a66bc6;
assign v373d219 = hgrant4_p & v3746cc0 | !hgrant4_p & v8455ab;
assign v37712b7 = hmaster2_p & v376460f | !hmaster2_p & !v380951e;
assign v377360d = hbusreq7_p & v3a6ef3e | !hbusreq7_p & !v8455ab;
assign v3767e6a = jx0_p & v3a621d5 | !jx0_p & v3a6277d;
assign v374fbb6 = hmaster2_p & v3a6bc65 | !hmaster2_p & !v3775bd3;
assign v372e468 = hgrant6_p & v8455ab | !hgrant6_p & v3a5706c;
assign v37666f6 = hgrant4_p & v8455ab | !hgrant4_p & v3760fb0;
assign v375fa8b = hbusreq3_p & v3760ab8 | !hbusreq3_p & !v8455ab;
assign v3a6fcc3 = hgrant4_p & v3a6eaf4 | !hgrant4_p & v3a5db8b;
assign v360d1b0 = hmaster2_p & v8455ab | !hmaster2_p & v3a6595f;
assign v3a5f648 = hmaster0_p & v3a62ad0 | !hmaster0_p & v3a6be79;
assign v3a6eff6 = hbusreq7_p & v37249fe | !hbusreq7_p & v3a672b6;
assign v3a2951d = hmaster1_p & v3769e01 | !hmaster1_p & v3a6acd3;
assign v375ba37 = hgrant6_p & v37245f8 | !hgrant6_p & v3a62a53;
assign v373ca8d = hgrant4_p & v373bf6a | !hgrant4_p & v8455ab;
assign v3a544db = hbusreq6_p & v37485ec | !hbusreq6_p & v3a6fe06;
assign v3a6fe4a = hbusreq5 & v8455e7 | !hbusreq5 & v8455ab;
assign c39ea5 = hbusreq7_p & v372a7c1 | !hbusreq7_p & !v373b785;
assign v3753dab = hready & v3735ed0 | !hready & !v8455ab;
assign v37249c7 = hmaster0_p & v3a68c94 | !hmaster0_p & v3a6cf7f;
assign v3a7071a = hmaster2_p & v3a63805 | !hmaster2_p & v377ef4a;
assign v37697e2 = hlock3_p & v3735436 | !hlock3_p & v3761224;
assign v376c017 = hbusreq2 & v37270d9 | !hbusreq2 & v8455e7;
assign v3a56864 = hbusreq3_p & v377ddae | !hbusreq3_p & !v8455ab;
assign v3a58a90 = hlock4_p & v373006f | !hlock4_p & !v8455ab;
assign v372efc8 = hbusreq5 & v3a70b3c | !hbusreq5 & v373af6f;
assign v3762a2a = hgrant6_p & v8455ab | !hgrant6_p & v376adaf;
assign v3725de9 = hmaster0_p & v374f92e | !hmaster0_p & v3a6cf7f;
assign v3736b43 = hmaster0_p & v372404f | !hmaster0_p & v3753097;
assign v377fb43 = hbusreq4_p & v373b4e6 | !hbusreq4_p & v373f647;
assign v373f394 = hmaster2_p & v3725198 | !hmaster2_p & v377169f;
assign v3a5f4c6 = hmaster0_p & v3a635ea | !hmaster0_p & v376a3c2;
assign v376a65a = hgrant6_p & v8455ab | !hgrant6_p & v3a6fd15;
assign v8455ca = hbusreq6 & v8455ab | !hbusreq6 & !v8455ab;
assign v377dc87 = hbusreq1 & v372fba5 | !hbusreq1 & v8455ab;
assign v3732c52 = hbusreq0_p & v376f9a8 | !hbusreq0_p & !v376d45f;
assign v3a69df3 = hmaster1_p & v3a619c0 | !hmaster1_p & v376eed1;
assign v3744af7 = hbusreq8 & v377b8c5 | !hbusreq8 & v8455ab;
assign v3759379 = hbusreq2_p & v37598a3 | !hbusreq2_p & v8455ab;
assign v3730afc = hgrant6_p & v374bc10 | !hgrant6_p & v3a70e07;
assign v376ad33 = hmaster1_p & v8455ab | !hmaster1_p & v3725036;
assign v3a70b2f = hbusreq5 & v3737dee | !hbusreq5 & v8455ab;
assign v3a5fc34 = hbusreq0 & v3a69487 | !hbusreq0 & v8455ab;
assign v373c164 = jx1_p & v3a70a64 | !jx1_p & v3a5f60f;
assign v374eab4 = hbusreq6_p & a75a41 | !hbusreq6_p & v8455ab;
assign v3764677 = hmaster0_p & v376111d | !hmaster0_p & v37432e2;
assign ab0224 = hmaster2_p & v3a635ea | !hmaster2_p & v3771d4f;
assign v3751606 = hbusreq5_p & v3757d5b | !hbusreq5_p & v37674d1;
assign v377d6c5 = jx1_p & v3a6f657 | !jx1_p & v3762f14;
assign v3764e58 = hmaster0_p & v3a63c47 | !hmaster0_p & v374077c;
assign v377e52f = hbusreq2_p & v38099ce | !hbusreq2_p & v3730b62;
assign v374a19d = hgrant6_p & v3a6ecd9 | !hgrant6_p & v375e948;
assign v3a6e6c9 = hbusreq6 & v3a5c00e | !hbusreq6 & v8455ab;
assign v376858c = hgrant7_p & v8455bd | !hgrant7_p & v3730a6a;
assign v3745928 = hmaster1_p & v3a59c12 | !hmaster1_p & v8455ab;
assign v3a6487f = hbusreq4 & v3a6f24c | !hbusreq4 & v8455ab;
assign v3767885 = hbusreq3 & v3735580 | !hbusreq3 & v372c6fb;
assign v376b7e1 = hbusreq5_p & v3a63c12 | !hbusreq5_p & v37796e9;
assign v374f0bb = hgrant8_p & v8455ab | !hgrant8_p & v374f4ae;
assign v3a6f3b1 = hbusreq2 & v3725230 | !hbusreq2 & v8455ab;
assign v37672a5 = hlock2 & v373c9b1 | !hlock2 & v3a6f4ac;
assign v375df95 = hgrant6_p & v8455ab | !hgrant6_p & v3761ac7;
assign v377cc69 = hmaster2_p & v377234d | !hmaster2_p & v375f61e;
assign v3a70ed7 = hgrant4_p & v377dd4e | !hgrant4_p & v8455ab;
assign v372c762 = hbusreq5_p & v376f9ca | !hbusreq5_p & !v8455ab;
assign v37681fa = hbusreq1_p & v3744982 | !hbusreq1_p & !v8455ab;
assign v3749f3b = hgrant5_p & v3773f27 | !hgrant5_p & v3a63f6b;
assign v3a5a1ba = hgrant3_p & v3a6f627 | !hgrant3_p & v3a65436;
assign v374bd1f = hmaster1_p & v377a3bd | !hmaster1_p & v3a6a57c;
assign v3739a33 = hmaster3_p & v3738f36 | !hmaster3_p & v3741bd4;
assign v3728650 = hmaster0_p & v3771ce2 | !hmaster0_p & v39a52b7;
assign v3a5950d = hmaster2_p & v374a08a | !hmaster2_p & v37364cf;
assign v3742e6b = hgrant4_p & v8455ab | !hgrant4_p & v377d651;
assign v37795d3 = hgrant4_p & v3758aec | !hgrant4_p & v374b32b;
assign v3a6c363 = decide_p & v3750295 | !decide_p & v3a5946d;
assign v3769c4c = hmaster1_p & v3773103 | !hmaster1_p & v373a0dc;
assign v3749bc0 = hbusreq5 & v376d8fd | !hbusreq5 & !v3a56f9d;
assign v372a95a = hbusreq7_p & v3a709cd | !hbusreq7_p & v3747020;
assign v372f3e8 = hgrant4_p & v8455ab | !hgrant4_p & v3756eca;
assign v37c03ff = hbusreq8_p & v376740b | !hbusreq8_p & v3a661cd;
assign v373643b = hlock7 & v3731517 | !hlock7 & v373aa47;
assign v3739d2a = hbusreq5 & v374c0a4 | !hbusreq5 & v3770700;
assign v3778083 = hmaster2_p & v8455ab | !hmaster2_p & v37494a9;
assign v3a595b8 = hbusreq0 & v372339a | !hbusreq0 & v3a59d59;
assign v3a70526 = hbusreq2 & v39a5265 | !hbusreq2 & !v2acb5a2;
assign v373f200 = hgrant6_p & v8455ab | !hgrant6_p & v376bb9f;
assign v377b4fb = hlock3 & v373c3e4 | !hlock3 & v3a6500c;
assign v3749356 = hgrant4_p & v37692c1 | !hgrant4_p & v376a9ee;
assign v37356a7 = hbusreq5_p & v373dc5a | !hbusreq5_p & !v8455ab;
assign v375e232 = hgrant3_p & v377b6ce | !hgrant3_p & v372b445;
assign v3a6ef47 = hmaster0_p & v3a659e5 | !hmaster0_p & v37420bb;
assign v377be84 = hmaster0_p & v376111d | !hmaster0_p & v375647b;
assign v3a6c127 = hbusreq8 & v3a6b0a1 | !hbusreq8 & v37258d0;
assign v372fc9d = hlock0_p & v3806db7 | !hlock0_p & v8455b0;
assign v38069c0 = hbusreq8 & v376af8e | !hbusreq8 & a0a219;
assign v3735324 = hgrant4_p & v8455ab | !hgrant4_p & v3a6b3d4;
assign v3769a6c = hmaster1_p & v3754a74 | !hmaster1_p & v373aa0e;
assign v3a6680b = hmaster1_p & v3a7046c | !hmaster1_p & v3738826;
assign v3a70157 = hmaster1_p & v8455ab | !hmaster1_p & v3768695;
assign v3766d07 = hbusreq4_p & v3a6d625 | !hbusreq4_p & v3809240;
assign v3a69913 = hbusreq5_p & d24921 | !hbusreq5_p & v3a713ad;
assign v3a6fa1d = hlock7 & v3768a43 | !hlock7 & v376ed58;
assign v3740d3b = hgrant4_p & v37496fa | !hgrant4_p & v3749bf0;
assign v3777586 = hgrant5_p & v3a702d0 | !hgrant5_p & v3725ad3;
assign v3770116 = hbusreq3_p & v375b012 | !hbusreq3_p & v8455b0;
assign v3a71547 = hgrant3_p & v377abd1 | !hgrant3_p & v372538e;
assign v376b8c2 = hmaster0_p & v3a6b60d | !hmaster0_p & v39eb431;
assign v37398a1 = hmaster1_p & v3a70221 | !hmaster1_p & v3a5c9df;
assign v3759265 = hmaster0_p & v8455ab | !hmaster0_p & !v372e466;
assign v3a6fc1a = hmaster3_p & v3726a8d | !hmaster3_p & v3756960;
assign v3733480 = hlock8 & v376cd8f | !hlock8 & v3762712;
assign v3a70d22 = hbusreq3_p & v3774e8c | !hbusreq3_p & v3736fdd;
assign v3725f3e = hbusreq6_p & v3773a5b | !hbusreq6_p & v3765261;
assign v376fbfe = hgrant4_p & v8455ab | !hgrant4_p & v3a623cb;
assign v374e16a = hbusreq0_p & v374f35a | !hbusreq0_p & v3a68d2e;
assign v3739a05 = hbusreq5 & v3a67b93 | !hbusreq5 & v8455ab;
assign v372d490 = hbusreq2 & v375ac23 | !hbusreq2 & v8455ab;
assign v3a70264 = hbusreq5 & v3a6fb40 | !hbusreq5 & v3768343;
assign v3a55641 = hgrant6_p & v8455ab | !hgrant6_p & v373d293;
assign v372bda4 = hmaster1_p & v360d2c6 | !hmaster1_p & !v8455ab;
assign v2092ac3 = hmaster0_p & v375cbe2 | !hmaster0_p & !v1e37cf9;
assign v3a6b798 = hmaster1_p & v8455ab | !hmaster1_p & v377dcf5;
assign v374933f = hgrant6_p & v3a57b60 | !hgrant6_p & v377b779;
assign v376e5ab = hmaster2_p & v3a635ea | !hmaster2_p & v3a709f2;
assign v374189b = hbusreq2_p & v3a68e39 | !hbusreq2_p & v37344c6;
assign v374ebb0 = hbusreq3_p & v373fa07 | !hbusreq3_p & v8455b0;
assign v3724b93 = hgrant3_p & v3775b81 | !hgrant3_p & v8455ab;
assign v374bbbf = hgrant1_p & v376563d | !hgrant1_p & v375f077;
assign v376fd9a = hmaster2_p & v3a6f9b3 | !hmaster2_p & v3738cab;
assign v37592a3 = hbusreq4_p & v3748858 | !hbusreq4_p & v3a70d94;
assign v3a70bbc = stateG10_1_p & v375f077 | !stateG10_1_p & v374bbbf;
assign v3760707 = hlock6_p & v37716c3 | !hlock6_p & v3a7084e;
assign v3a6f608 = hmaster2_p & v3a635ea | !hmaster2_p & v374d0e3;
assign v3741d51 = hgrant3_p & v8455ab | !hgrant3_p & v375c8b0;
assign v37499c4 = jx1_p & v377260b | !jx1_p & v8f2b25;
assign v373df3d = hgrant3_p & v3a712f0 | !hgrant3_p & v37667f9;
assign v3726634 = hbusreq5 & v377db89 | !hbusreq5 & v8455ab;
assign v3a5b404 = hmaster2_p & v8455ab | !hmaster2_p & !v3a6ffe1;
assign v37748e5 = hbusreq1 & v3a6f428 | !hbusreq1 & v38072fd;
assign v373e814 = hgrant6_p & v8455ab | !hgrant6_p & v373a2f2;
assign v3a65aeb = hbusreq4 & v3a6fa84 | !hbusreq4 & !v372acab;
assign v3a707f9 = hmaster2_p & v374d4e6 | !hmaster2_p & v3a70bf4;
assign v373f8d4 = hlock4_p & v3a68838 | !hlock4_p & v8455b0;
assign v3a55e7f = hgrant3_p & v8455be | !hgrant3_p & !v373d9aa;
assign v3a5907f = hgrant5_p & v37781fe | !hgrant5_p & v3a6f487;
assign v3a63306 = hmaster0_p & v3743522 | !hmaster0_p & !v3735f79;
assign v3a5b071 = hmaster2_p & v372d299 | !hmaster2_p & v37762bd;
assign v3768fe7 = hgrant4_p & v3a6eeef | !hgrant4_p & v3a702b6;
assign v3a6fa19 = hbusreq6_p & v376041f | !hbusreq6_p & !v8455ab;
assign v3a61895 = hgrant6_p & v3739884 | !hgrant6_p & v376d328;
assign v3a712f2 = hbusreq0 & v337900b | !hbusreq0 & v3a6ec76;
assign v3a70b98 = hmaster2_p & v372580e | !hmaster2_p & v8455ab;
assign v3a5dc67 = hbusreq5 & v37548f5 | !hbusreq5 & v3728903;
assign v374e684 = hmaster1_p & v3756e39 | !hmaster1_p & v373a973;
assign v3772715 = hgrant4_p & v8455ab | !hgrant4_p & v2ff8e9c;
assign v3756219 = hmaster2_p & v376025f | !hmaster2_p & !v8455ab;
assign v3a5d03e = hlock7 & v3a6f6e8 | !hlock7 & v3762ac3;
assign v3745bdc = hmaster2_p & v3a635ea | !hmaster2_p & v3727943;
assign v3a71132 = hbusreq5 & v372abac | !hbusreq5 & v3762dc3;
assign v3746200 = hmaster0_p & v3a6f7dd | !hmaster0_p & v3769d48;
assign v3a59e87 = hbusreq1_p & v3a6f814 | !hbusreq1_p & !v3a58aa5;
assign v373a11f = hbusreq5_p & v376e6ac | !hbusreq5_p & !v37431bb;
assign v3a70f4d = hmaster0_p & v37635ab | !hmaster0_p & v35b71da;
assign v375da36 = hmaster2_p & v373ad95 | !hmaster2_p & !v8455ab;
assign v3762fc4 = hmastlock_p & v3727fe3 | !hmastlock_p & !v8455ab;
assign v372febd = hbusreq0 & v376af98 | !hbusreq0 & v3770f55;
assign v3747dd8 = hmaster2_p & v3a7093c | !hmaster2_p & v377a9e7;
assign v3a6906e = hbusreq5_p & v3a5d96d | !hbusreq5_p & v374819d;
assign v3753ee0 = hbusreq0 & v3a70960 | !hbusreq0 & v3a71473;
assign v37462ed = hmaster2_p & v8455ab | !hmaster2_p & !v3a7053b;
assign v2092f90 = hlock3_p & v3a70e71 | !hlock3_p & v8455b0;
assign v372a288 = hlock7 & v3743cf5 | !hlock7 & v3a70454;
assign v3a5f83e = hgrant6_p & v3a708bd | !hgrant6_p & v377094b;
assign v372e466 = hmaster2_p & v8455e7 | !hmaster2_p & v3a70641;
assign v3755305 = hgrant6_p & v3a6eeef | !hgrant6_p & v372d434;
assign v8455bb = hlock2_p & v8455ab | !hlock2_p & !v8455ab;
assign v372d939 = hmaster2_p & v3a68838 | !hmaster2_p & v375070c;
assign v376051c = hbusreq0 & v3739c81 | !hbusreq0 & v374fa4d;
assign v373f19e = hbusreq1 & v3743b9e | !hbusreq1 & v3a6a195;
assign v3a70cc6 = hgrant5_p & v8455ab | !hgrant5_p & v3a6850e;
assign v3761ae0 = hmaster2_p & v372707d | !hmaster2_p & v372615f;
assign v3759584 = hmaster2_p & v376fbe0 | !hmaster2_p & v3763d20;
assign v3a6f676 = hmaster2_p & v3a635ea | !hmaster2_p & v3750adf;
assign v3a685c7 = hbusreq6_p & v373f0ee | !hbusreq6_p & v3a69946;
assign v3736aaa = hgrant6_p & v3779c33 | !hgrant6_p & v8455ab;
assign v3737aee = hmaster1_p & v3a61a7f | !hmaster1_p & v373a876;
assign v37649ee = hbusreq3_p & v3a6edb1 | !hbusreq3_p & bc7f17;
assign v3a70ab1 = hbusreq5 & v377c67b | !hbusreq5 & v3756a5f;
assign v375f8dd = hgrant6_p & v3737571 | !hgrant6_p & v94e000;
assign v3776751 = hbusreq2_p & v3a6a261 | !hbusreq2_p & v37649ab;
assign v3a59cf3 = hbusreq5 & db32f1 | !hbusreq5 & v8455ab;
assign v372f2ed = hmaster2_p & v35772a5 | !hmaster2_p & !v373bd76;
assign v37285a1 = hbusreq3 & v37794fa | !hbusreq3 & !v8455ab;
assign v376112d = hgrant4_p & v8455ab | !hgrant4_p & v3a6ffcc;
assign v374159f = hbusreq8 & v3a710ff | !hbusreq8 & v3a6abfe;
assign v374a98e = hlock7 & v373f6f7 | !hlock7 & v3a6a8b4;
assign v3737b54 = hmaster0_p & v373e74b | !hmaster0_p & v37291e7;
assign v3a5d48f = hbusreq2_p & v3749a38 | !hbusreq2_p & v374abc9;
assign v37467a3 = hlock0_p & v3a70385 | !hlock0_p & !v3744710;
assign v3751539 = hbusreq8_p & v3a6f121 | !hbusreq8_p & v8455ab;
assign v3764761 = hmaster0_p & v3a5d217 | !hmaster0_p & v373e16b;
assign v37523dd = hmaster0_p & v3a60a24 | !hmaster0_p & v3761719;
assign v374e0ba = hbusreq1_p & bda6d5 | !hbusreq1_p & !v3a58836;
assign v3a708a7 = hmaster2_p & v3746806 | !hmaster2_p & v376d882;
assign v3a7155c = hgrant4_p & v8455b2 | !hgrant4_p & v377f785;
assign v3759ff9 = hbusreq8_p & v37550ac | !hbusreq8_p & !v8455ab;
assign v3735ad2 = hbusreq4 & v376f2a7 | !hbusreq4 & v37496fa;
assign v3a5a45e = hmaster0_p & v37606f0 | !hmaster0_p & v3a62a6d;
assign v372c7b7 = jx0_p & v375b0f9 | !jx0_p & v3726111;
assign v2092b23 = hbusreq2 & v372f3f7 | !hbusreq2 & v3a6a393;
assign v37701af = hmaster2_p & v3a635ea | !hmaster2_p & v37330dc;
assign v3727d18 = hmaster0_p & c0c2de | !hmaster0_p & !v3733cd1;
assign v3a6fcea = hmaster2_p & v377169f | !hmaster2_p & v37716c3;
assign v3a58971 = hmaster2_p & v3729421 | !hmaster2_p & !v8455ab;
assign v375029a = hmaster0_p & v37486de | !hmaster0_p & v37614c1;
assign v38064dd = hlock5_p & v3a71585 | !hlock5_p & v3a2abf5;
assign v3a592be = hbusreq4_p & v3752707 | !hbusreq4_p & v377d8b3;
assign v37752be = hmaster0_p & v37445a8 | !hmaster0_p & v3776cbb;
assign v374a343 = hbusreq6_p & v3a58d7a | !hbusreq6_p & v8455ab;
assign v3a703dd = hburst1 & v3749a12 | !hburst1 & v3753a28;
assign v3746efb = hlock6_p & v374f87c | !hlock6_p & v8455b0;
assign v373aa47 = hbusreq7 & v377b94e | !hbusreq7 & v3751012;
assign v3770af6 = hmaster0_p & v3a6c4e4 | !hmaster0_p & v3769280;
assign v3a683a4 = hbusreq2_p & v3a6c688 | !hbusreq2_p & v8455ab;
assign v3754f54 = hgrant3_p & v35b7299 | !hgrant3_p & !v3733d5a;
assign v3745939 = hbusreq5_p & v3737415 | !hbusreq5_p & dac24d;
assign v375bfa6 = hlock6_p & v3773b23 | !hlock6_p & v8455b0;
assign v3a70467 = hmaster0_p & v8455ab | !hmaster0_p & v3731d76;
assign v377606f = hburst1 & v3a6f776 | !hburst1 & v37618dc;
assign v3a6039a = hgrant4_p & v373b3a8 | !hgrant4_p & v3749c8a;
assign v3764ed7 = hmaster2_p & v375166c | !hmaster2_p & v373ad7b;
assign v3752dc7 = hlock5 & v3a6bbe3 | !hlock5 & v3a709fb;
assign v3a70971 = hmaster0_p & v3a6fab6 | !hmaster0_p & v377312f;
assign v3a5e81d = hgrant3_p & v3723b00 | !hgrant3_p & v3750037;
assign v376f409 = hgrant4_p & v8455ab | !hgrant4_p & v3763d79;
assign v3a6f28b = hbusreq7 & v3806c04 | !hbusreq7 & v37644b7;
assign v372b847 = hbusreq0 & v3740469 | !hbusreq0 & v3773434;
assign v373f051 = hgrant3_p & v3774416 | !hgrant3_p & !v3a6442f;
assign v377226d = hgrant6_p & v3752a0d | !hgrant6_p & v3766c7b;
assign v3a6ff29 = hbusreq4_p & v374a2f3 | !hbusreq4_p & v3731a1f;
assign v3746fdb = hbusreq5 & v375977c | !hbusreq5 & v377bcb3;
assign v3a6f886 = jx0_p & v37465d7 | !jx0_p & v3750f3b;
assign v3a58b13 = hmaster2_p & v3758fa8 | !hmaster2_p & v373bcb6;
assign v375899b = hbusreq3 & v374ec84 | !hbusreq3 & v3a6c5fc;
assign v3762f76 = hbusreq0 & v375c317 | !hbusreq0 & v3a6a6c1;
assign v3748e0c = hlock5 & v3730fbd | !hlock5 & v3a6a6e1;
assign v377a275 = hbusreq1 & v3a7151d | !hbusreq1 & !v8455ab;
assign v3755cb2 = hbusreq2_p & v3a71652 | !hbusreq2_p & !v8455ab;
assign v377576e = hmaster2_p & v3769e7f | !hmaster2_p & v8455ab;
assign v37532cd = hmaster1_p & v3a70675 | !hmaster1_p & v37402ee;
assign v37c00b6 = hbusreq2_p & v375e4a0 | !hbusreq2_p & v3724f7b;
assign v3724c35 = hgrant6_p & v8455ab | !hgrant6_p & v3727849;
assign v376beb4 = hlock6 & v374376b | !hlock6 & v373b11b;
assign v3a70279 = hbusreq6 & v3766a74 | !hbusreq6 & v3a5a8bf;
assign v372dfc3 = hmaster0_p & v3a67d66 | !hmaster0_p & v3758a96;
assign v373ae6a = hmaster0_p & v3a68848 | !hmaster0_p & v373e2e5;
assign v3a7127d = hbusreq5_p & v373946b | !hbusreq5_p & v3a5b615;
assign v376aa99 = hlock0 & v372348c | !hlock0 & v375a7d3;
assign v3806f67 = hbusreq1_p & v37c101a | !hbusreq1_p & !v8455ab;
assign v3a631d0 = hmaster1_p & v3a6ae45 | !hmaster1_p & v3748229;
assign v3738a93 = hmaster0_p & v3742f0b | !hmaster0_p & v3722caa;
assign v373de18 = hmaster2_p & v3a707c4 | !hmaster2_p & !v3a713c9;
assign v372fd0a = hlock4_p & v373aaa8 | !hlock4_p & !v8455ab;
assign v376f549 = hmaster1_p & v8455e7 | !hmaster1_p & v3a69d8f;
assign v3a6e08c = hmaster0_p & v8455ab | !hmaster0_p & v3771e6f;
assign v37361a0 = hbusreq5 & v37665c5 | !hbusreq5 & v37744a3;
assign v374b237 = hmaster3_p & v3a2986b | !hmaster3_p & v3a70a53;
assign v376824b = hmaster0_p & v3a5c3a0 | !hmaster0_p & v376d93b;
assign v2092b2f = stateA1_p & v3757c6f | !stateA1_p & !v3a71085;
assign v375ad79 = hbusreq8 & v3a60f1a | !hbusreq8 & v375538e;
assign v37304a0 = hgrant5_p & v8455ab | !hgrant5_p & v376d7d5;
assign v3a6d9fa = hbusreq6 & v3806ec4 | !hbusreq6 & v3a59391;
assign v3a5e859 = hmaster0_p & v3779d33 | !hmaster0_p & v374e519;
assign v3a5b925 = hbusreq7 & v3a70d7e | !hbusreq7 & v375b56c;
assign v376e00a = hgrant1_p & v8455b6 | !hgrant1_p & v3774b25;
assign v3772a3f = hbusreq4_p & v325b59f | !hbusreq4_p & v3a588a0;
assign v37249ff = hbusreq5_p & v3759bf4 | !hbusreq5_p & v375c9b9;
assign v3760ff4 = hbusreq2_p & v3a635ea | !hbusreq2_p & v377c6b3;
assign v3740171 = locked_p & v8455ab | !locked_p & v39a537f;
assign v37234e0 = hbusreq2_p & v3a5b42a | !hbusreq2_p & !v3773e09;
assign v3737c0d = hgrant4_p & v3a6f312 | !hgrant4_p & v37292df;
assign v3729f64 = hbusreq5_p & v377d077 | !hbusreq5_p & c6053a;
assign v3758ee1 = hmaster0_p & v2acaf2d | !hmaster0_p & v375fe03;
assign v3a7033f = hmaster1_p & v325c94d | !hmaster1_p & v372bc4c;
assign v3a6d621 = hgrant3_p & v372d828 | !hgrant3_p & !v8455ab;
assign v37367f1 = hbusreq6 & v3a67118 | !hbusreq6 & v8455ab;
assign v37653ef = hlock5_p & v3a6d9da | !hlock5_p & v37742a4;
assign v3a71504 = hmaster1_p & v8455ab | !hmaster1_p & v376b4a2;
assign v37581a6 = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v3728e1d;
assign v3a702a0 = hbusreq2_p & v375c705 | !hbusreq2_p & v3754871;
assign v3a6d329 = hmaster0_p & v3807aa1 | !hmaster0_p & v375dc9b;
assign v3776d33 = hgrant3_p & v377499f | !hgrant3_p & !v3a6ca1d;
assign v3a6f3a8 = hlock6_p & v376e914 | !hlock6_p & !v3a658bf;
assign v3758b78 = hmaster2_p & v374ccb7 | !hmaster2_p & v3a709e2;
assign v375d4f9 = hbusreq2_p & v3757598 | !hbusreq2_p & v37747b4;
assign v3730055 = hbusreq5 & v3a6178c | !hbusreq5 & v357742d;
assign v3a70e70 = hbusreq0 & v377a180 | !hbusreq0 & v3779925;
assign bb41ad = hmaster1_p & v3760091 | !hmaster1_p & v3a655e9;
assign v372ab85 = hbusreq1 & v3a70459 | !hbusreq1 & v373b288;
assign v37773c1 = hgrant3_p & v373cdbf | !hgrant3_p & v3726668;
assign v3a6d89d = hgrant5_p & v3a661d0 | !hgrant5_p & v372cace;
assign v375039e = hbusreq1_p & v3747302 | !hbusreq1_p & v360d03f;
assign v377ac7e = hgrant3_p & v8455be | !hgrant3_p & v3778765;
assign v3725b1f = hbusreq8_p & v373923a | !hbusreq8_p & v3a70472;
assign v376c611 = hmaster0_p & v3a6f942 | !hmaster0_p & v3a61e33;
assign v3a56c60 = hlock5 & v3a554f0 | !hlock5 & v373b380;
assign v3754e5e = hburst1 & v3a6ac2a | !hburst1 & v1e37cec;
assign v37775c7 = hgrant5_p & v3773e8d | !hgrant5_p & v37770df;
assign v9c492b = hbusreq2 & v374caab | !hbusreq2 & v8455ab;
assign v3a61b7f = hlock3 & v39eb4de | !hlock3 & v376e568;
assign v377a27f = hmaster1_p & v3a6efe8 | !hmaster1_p & v37266d1;
assign v376b088 = hbusreq6_p & v3763668 | !hbusreq6_p & v377167e;
assign v377d3bf = hbusreq7 & v373c2e1 | !hbusreq7 & v8455ab;
assign v3a6f22e = hbusreq6_p & v37243e6 | !hbusreq6_p & !v37450cb;
assign v3755220 = hmaster0_p & v3729187 | !hmaster0_p & v37276a8;
assign v3a711c0 = hmaster2_p & v3a63ea7 | !hmaster2_p & v373f058;
assign v3a7051c = hgrant3_p & v372ad53 | !hgrant3_p & v3a59833;
assign v3a576bd = hmaster1_p & v8455ab | !hmaster1_p & v3a5fd0a;
assign v373de86 = hlock5_p & v3a6a8ee | !hlock5_p & v8455c3;
assign v3a70aa2 = hbusreq0_p & v377094b | !hbusreq0_p & v8455ab;
assign v3a7050e = hmaster2_p & v3779801 | !hmaster2_p & !v3751510;
assign v377f6ff = hbusreq0_p & v374f0c1 | !hbusreq0_p & v3739e4c;
assign v376b678 = hbusreq7_p & v3738373 | !hbusreq7_p & v3a70c90;
assign v377807f = hmaster1_p & v376d1dd | !hmaster1_p & v3a298b6;
assign v3806599 = hlock5 & v37576e7 | !hlock5 & v37706ae;
assign v3766d5a = hlock0 & v376c76d | !hlock0 & v3a66c6c;
assign v38095b2 = hgrant2_p & v375d38f | !hgrant2_p & !v372e88a;
assign v3729700 = hbusreq2_p & v3767561 | !hbusreq2_p & !v8455ab;
assign v375ad90 = hmaster1_p & v3763175 | !hmaster1_p & v377f298;
assign v377cbc9 = hbusreq6_p & v374f0c1 | !hbusreq6_p & v376e1b7;
assign v3766de9 = hmaster0_p & v3a6af93 | !hmaster0_p & v375c278;
assign v373b76d = hgrant6_p & v373d35f | !hgrant6_p & !v8455ab;
assign v37697d0 = hlock8_p & v3a70e91 | !hlock8_p & v3777f6f;
assign v37408e1 = hbusreq6_p & v3a62a6d | !hbusreq6_p & v3a70b17;
assign v2092ffc = hgrant0_p & v3747302 | !hgrant0_p & v372dadb;
assign v3725578 = hbusreq0 & v373481c | !hbusreq0 & v3752eda;
assign v37299b3 = hgrant0_p & v8455ab | !hgrant0_p & v373905f;
assign v374f707 = hbusreq4_p & v375ff94 | !hbusreq4_p & v37651c2;
assign v377b3b0 = hlock5 & v3730651 | !hlock5 & ae0bd0;
assign v3724b1c = hlock6_p & v8455ab | !hlock6_p & v3a6ab5f;
assign v3a6ff06 = jx1_p & v3745196 | !jx1_p & v3a705c0;
assign v3779f68 = hlock7 & v37503f5 | !hlock7 & v3775903;
assign v37743c6 = hmaster1_p & v879494 | !hmaster1_p & v8455ab;
assign v3749ec1 = hmaster2_p & v3a6ffb6 | !hmaster2_p & !v3a5ef5c;
assign v377df77 = hbusreq8 & v98d1dc | !hbusreq8 & v3741e61;
assign v375ccf3 = hmaster1_p & v9af7ec | !hmaster1_p & v374c679;
assign v37652b1 = hbusreq3 & v3a6fe6a | !hbusreq3 & !v8455ab;
assign v3a6fbd4 = hbusreq6 & v374424e | !hbusreq6 & v8455ab;
assign v37594d4 = hmaster2_p & v8455ab | !hmaster2_p & v3a714cf;
assign v3748d3c = hbusreq7 & v3771633 | !hbusreq7 & v372863f;
assign v3750d06 = hlock0_p & v8455ab | !hlock0_p & v374b962;
assign v374e77f = hlock0_p & v3a6ac2a | !hlock0_p & v8455ab;
assign v3a7141d = hlock7_p & v92a8d7 | !hlock7_p & v3a6caab;
assign v3732899 = hmaster1_p & v375c740 | !hmaster1_p & v8455ab;
assign v3765af5 = hmaster0_p & v3a6f693 | !hmaster0_p & !v8455ab;
assign v3a53c50 = hbusreq6_p & v377e71d | !hbusreq6_p & v8455ab;
assign v3763dd5 = hbusreq4_p & db86c8 | !hbusreq4_p & !v8455ab;
assign v3767ba9 = jx3_p & v1e37b52 | !jx3_p & v3779b96;
assign v3a66747 = hgrant5_p & v3752def | !hgrant5_p & v3776f93;
assign v3a57b5a = hbusreq7 & v3a71008 | !hbusreq7 & v3a592d8;
assign v376157e = hbusreq4 & v375ac23 | !hbusreq4 & v8455ab;
assign v373541f = hbusreq0_p & v37744f5 | !hbusreq0_p & v3a6b4ae;
assign v3749a7c = hmaster1_p & v3a5af94 | !hmaster1_p & v3808531;
assign c29340 = hbusreq6 & v373ec72 | !hbusreq6 & v372cc25;
assign v3726838 = hbusreq6 & v8455cb | !hbusreq6 & !v8455ab;
assign v377b2f3 = hmaster2_p & v3a70172 | !hmaster2_p & v3a70d64;
assign v372d75d = hmaster0_p & v3735324 | !hmaster0_p & v3a6fbaa;
assign v8907fb = hbusreq6_p & v3a70893 | !hbusreq6_p & v373cd16;
assign v3a7089d = hgrant4_p & v8455ab | !hgrant4_p & v375cd5d;
assign v374ee77 = jx3_p & v374a7c3 | !jx3_p & v3a54a24;
assign v37487ca = hlock0_p & v3733e9e | !hlock0_p & v1e38224;
assign v3a6ab5e = hmaster2_p & v375808f | !hmaster2_p & v3a63bb7;
assign v377c490 = hmaster0_p & v39ea76e | !hmaster0_p & v9d7045;
assign v3755ed8 = hlock0 & v38072fd | !hlock0 & v3a636a7;
assign v3a614b1 = hbusreq4_p & v37259cc | !hbusreq4_p & !v8455ab;
assign v3770a5b = hbusreq5 & v3777d63 | !hbusreq5 & v3764a8a;
assign v97f405 = hgrant6_p & v8455c9 | !hgrant6_p & v3a5a853;
assign d2819e = hbusreq3 & v3752bcc | !hbusreq3 & v3a70452;
assign v3a6c922 = hmaster2_p & v375bb51 | !hmaster2_p & v37320ff;
assign v372eb0f = hmaster1_p & v373a2f4 | !hmaster1_p & v3a5744d;
assign v3771e95 = hgrant3_p & v3a5fcbc | !hgrant3_p & v376ab72;
assign v373d40a = hmaster2_p & v3a6126c | !hmaster2_p & v3a57593;
assign v376eca3 = hbusreq3 & v376bc4b | !hbusreq3 & v8455ab;
assign v3a5d7bf = hgrant0_p & v37356d4 | !hgrant0_p & v377a110;
assign v374068b = hbusreq2_p & v37431eb | !hbusreq2_p & v3a6f947;
assign v37599cb = hlock3 & v376a87b | !hlock3 & v3a6430c;
assign v3737a5a = hgrant4_p & v3738006 | !hgrant4_p & v871244;
assign v3a70397 = hgrant2_p & v377fc87 | !hgrant2_p & v3a701d1;
assign v377d60e = hbusreq0 & v3a6fc1d | !hbusreq0 & v376c203;
assign v3777a8a = hmaster0_p & v3a619c0 | !hmaster0_p & !v3a5c945;
assign v372ee41 = hgrant6_p & v3a6fbe4 | !hgrant6_p & v3770dcb;
assign v3a62bc6 = hmaster1_p & v974eb9 | !hmaster1_p & v8455ab;
assign v375295a = hmaster1_p & v377234d | !hmaster1_p & v3759a67;
assign v373c916 = hmaster0_p & v3a541f5 | !hmaster0_p & v8455ab;
assign v3763cf5 = hgrant1_p & v375c7b9 | !hgrant1_p & !v8455e1;
assign v3771be6 = hmaster0_p & v3a6fdd1 | !hmaster0_p & v37462ee;
assign v3a57f42 = hlock0_p & v375444e | !hlock0_p & v8455b0;
assign v3746f46 = hgrant6_p & v8455ca | !hgrant6_p & v3a6eb76;
assign v377a99d = hbusreq0 & v2ff8f8e | !hbusreq0 & v8455ab;
assign v3a59d6b = hbusreq8 & v3725e9a | !hbusreq8 & v3a60276;
assign v376e02e = hbusreq6 & v37495dc | !hbusreq6 & v3773b7b;
assign v3a70c4b = hbusreq5 & v372c3d7 | !hbusreq5 & v376c0c8;
assign v3722b91 = hbusreq5 & v3760644 | !hbusreq5 & v3767e7f;
assign v3736613 = hmaster2_p & v3a7002c | !hmaster2_p & v373891b;
assign v3763a20 = hlock3_p & v3a6a939 | !hlock3_p & !v8455ab;
assign v37497eb = hgrant1_p & v8455ab | !hgrant1_p & !v375003c;
assign v3a6f9bc = hlock6_p & v3a6eb39 | !hlock6_p & v35772a6;
assign v376e580 = hmaster2_p & v377fb09 | !hmaster2_p & v8455ab;
assign v3a69c98 = hgrant4_p & v3a5dd86 | !hgrant4_p & v8455ab;
assign aba148 = hbusreq4_p & v3a6a3ac | !hbusreq4_p & v8455ab;
assign v3a70bfa = hgrant2_p & v376218c | !hgrant2_p & v3809427;
assign v372b1dc = hbusreq3_p & v3a6241d | !hbusreq3_p & v8455ab;
assign v3a61b13 = hbusreq7 & v1e37a35 | !hbusreq7 & v3a684ee;
assign v3757a2b = hlock7 & v3734279 | !hlock7 & v3754c4a;
assign v3760464 = hlock0 & v37651c2 | !hlock0 & v3746ef3;
assign v376b3d0 = hmaster0_p & v3a5ff4b | !hmaster0_p & v3753b80;
assign v374db6a = hbusreq4_p & v376e041 | !hbusreq4_p & v3748d67;
assign v3772b00 = hgrant4_p & v3a53eeb | !hgrant4_p & v3a56aae;
assign v37730cd = hbusreq8 & v3a6f820 | !hbusreq8 & v3777d70;
assign v3a67f5c = jx1_p & v3a6f827 | !jx1_p & v3749762;
assign v3765321 = hbusreq4_p & v3a6f5a1 | !hbusreq4_p & v8455ab;
assign v3a6494a = hgrant0_p & v3740083 | !hgrant0_p & !v3a714f0;
assign v373a9ef = hmaster0_p & v372455c | !hmaster0_p & v3a5d763;
assign v3a6f778 = hbusreq2_p & v3a58218 | !hbusreq2_p & v3770578;
assign v374d451 = hbusreq5_p & v3a5f33d | !hbusreq5_p & fc6f92;
assign v376dcd0 = hlock6_p & v373fe5e | !hlock6_p & !v8455ab;
assign v37321b8 = hbusreq2_p & v3a5fe72 | !hbusreq2_p & v373cb2d;
assign v3a5cf53 = hlock3 & v3747c93 | !hlock3 & v374cc2a;
assign v3746289 = hbusreq6_p & v3772add | !hbusreq6_p & v377957e;
assign v3577392 = hmaster2_p & v3a6fa88 | !hmaster2_p & v3775684;
assign v3a70d67 = hlock3_p & v3a6c063 | !hlock3_p & !v8455ab;
assign v37424b5 = hgrant3_p & v9f7a48 | !hgrant3_p & v3751d87;
assign v3a62d48 = hbusreq4_p & v373b838 | !hbusreq4_p & !v37287bd;
assign aadac1 = hbusreq3 & v372fc81 | !hbusreq3 & !v8455ab;
assign v3729972 = hlock5 & v37542a0 | !hlock5 & v3a5ef9d;
assign v360caba = hgrant5_p & v8455c6 | !hgrant5_p & v3769141;
assign v3a7069e = hlock1_p & v8455e7 | !hlock1_p & !v37547c9;
assign v3a6f41f = hlock8_p & v3a5e874 | !hlock8_p & !v8455ab;
assign v3a67555 = hbusreq5_p & v3a5d522 | !hbusreq5_p & v3777da6;
assign v376ac9b = hlock2_p & v3a6a1b9 | !hlock2_p & !v8455ab;
assign v3741f08 = hlock0 & v374165f | !hlock0 & v372a13a;
assign v3a6ca0b = hmaster0_p & v3a7167d | !hmaster0_p & v3a583b0;
assign v3a61bef = hgrant5_p & v3725626 | !hgrant5_p & v3a6f7f2;
assign v372a4ae = hlock8 & dbf06b | !hlock8 & v3a5be3f;
assign v3a65da2 = hbusreq2 & v3a70923 | !hbusreq2 & v3a641d5;
assign v376f903 = hgrant4_p & v3775537 | !hgrant4_p & v3a6ffd5;
assign v3a69a4c = hbusreq5 & v3763b37 | !hbusreq5 & v3a70448;
assign v3742fc4 = hbusreq7_p & v3a61a37 | !hbusreq7_p & v375bed5;
assign v39ebab4 = hbusreq0 & v3729cfe | !hbusreq0 & v374052a;
assign v3a58e44 = hmaster0_p & v372ae6f | !hmaster0_p & !v37744d9;
assign v3a5abf4 = hlock4_p & v377ea86 | !hlock4_p & !v8455ab;
assign v373ea09 = hlock5 & v3759786 | !hlock5 & v375aff6;
assign v3745ae6 = jx0_p & v376aaf5 | !jx0_p & v3a6360c;
assign v3a711cb = hmaster0_p & v3a635ea | !hmaster0_p & v374aacc;
assign v3748f33 = hbusreq4 & v375d0ed | !hbusreq4 & v3757559;
assign v3742d2a = hmaster1_p & v3a697d2 | !hmaster1_p & v3a6f937;
assign v3753e49 = hgrant6_p & v37418ac | !hgrant6_p & v3728526;
assign v38073fd = hbusreq3 & v373fe5e | !hbusreq3 & !v3753f1a;
assign v3a63af6 = hbusreq1 & v3a568f7 | !hbusreq1 & !v8455ab;
assign v3a66e70 = hgrant3_p & v3a6f2b8 | !hgrant3_p & v8455ab;
assign v3a679e2 = hmaster0_p & v376342f | !hmaster0_p & v3761c61;
assign v375f90e = hmaster0_p & v3735b31 | !hmaster0_p & v3775219;
assign v373291e = hlock0 & v373bd6c | !hlock0 & v376d05f;
assign v3759a27 = hgrant4_p & v8455ab | !hgrant4_p & v372b4a0;
assign v3768495 = hgrant4_p & v376a6f1 | !hgrant4_p & v3a63f0c;
assign v37561e0 = hbusreq8_p & v374e08e | !hbusreq8_p & v3a6f951;
assign v373a973 = hbusreq5_p & v3a71459 | !hbusreq5_p & v3a6fd31;
assign v37509c4 = hbusreq8 & v372c1bb | !hbusreq8 & v373168f;
assign v3a6d951 = hbusreq6 & v376a14f | !hbusreq6 & v8455ab;
assign v3a70955 = hmaster1_p & v3a640e3 | !hmaster1_p & v3745b39;
assign v372d360 = hbusreq8_p & v375f2ab | !hbusreq8_p & !v374b8fe;
assign v37473ca = hbusreq4 & v376a21e | !hbusreq4 & v3768751;
assign v3a6f45d = hmaster1_p & v374e784 | !hmaster1_p & v3773ab1;
assign v3a7001c = hbusreq7_p & v3a5b3dc | !hbusreq7_p & v376e66e;
assign v372f192 = hgrant2_p & v3a5ff76 | !hgrant2_p & v37565ae;
assign v3760d16 = hbusreq4 & v372313c | !hbusreq4 & v37285eb;
assign v3a65241 = hbusreq6 & v3a70200 | !hbusreq6 & !v37621b5;
assign v372546e = hgrant2_p & v376218c | !hgrant2_p & v377437f;
assign v3733d4f = hlock5_p & v376b438 | !hlock5_p & v8455bf;
assign v3723185 = hmaster2_p & v373f058 | !hmaster2_p & v375070c;
assign v3763a29 = hlock7_p & v3809fbb | !hlock7_p & v3a6f00d;
assign v3a71483 = hgrant5_p & v3a700c1 | !hgrant5_p & v372f739;
assign v3a6eee4 = hgrant6_p & v8455ab | !hgrant6_p & v3775a7d;
assign v375ed37 = hbusreq5 & v3a57de9 | !hbusreq5 & v3744aa9;
assign v3755549 = hgrant5_p & v8455ab | !hgrant5_p & b5da28;
assign v3a62812 = hmaster1_p & v37557a0 | !hmaster1_p & v8e42b4;
assign v3a6f1a5 = hgrant6_p & v3a71304 | !hgrant6_p & !v8ed2d8;
assign v9e8d30 = hmaster0_p & v377d107 | !hmaster0_p & v3a7029e;
assign v374b077 = hbusreq0 & v372d8e2 | !hbusreq0 & v377caa3;
assign v373940c = hmaster1_p & v372f2fe | !hmaster1_p & v3743b2c;
assign v377574b = hmaster2_p & v8455ab | !hmaster2_p & v3a68ef7;
assign v3764437 = hmaster0_p & v373a27c | !hmaster0_p & v374b204;
assign v3772add = hbusreq3_p & v37734ba | !hbusreq3_p & !v8455ab;
assign v91a14c = hgrant2_p & v3a5b90b | !hgrant2_p & !v8455ab;
assign v374837b = hmaster1_p & b3a152 | !hmaster1_p & !v3777efb;
assign v37512b3 = hmaster2_p & v37245f8 | !hmaster2_p & v2ff9314;
assign v375c52f = hlock4 & v3a6afef | !hlock4 & v3a710ad;
assign v376e76f = hgrant0_p & v374306c | !hgrant0_p & v3750deb;
assign v373422b = hbusreq0 & v37509a3 | !hbusreq0 & v3a6f5fe;
assign v3747b74 = hmaster1_p & v373a1b4 | !hmaster1_p & v3777763;
assign v373ef01 = hlock4_p & v377b8ee | !hlock4_p & !v8455ab;
assign v3a6d299 = hlock6 & v3753923 | !hlock6 & v38090f6;
assign v376cba1 = hbusreq8 & v3a64bb1 | !hbusreq8 & v374c790;
assign v372e8cc = hgrant6_p & v8455ab | !hgrant6_p & v376780f;
assign v3a71506 = hmaster0_p & v3a6f2f5 | !hmaster0_p & v3762ffa;
assign v374039d = hmaster1_p & a33229 | !hmaster1_p & v376ad8c;
assign v37572b6 = hmaster1_p & v376634c | !hmaster1_p & v3a5cfbb;
assign v3a5faba = hbusreq4 & v377834b | !hbusreq4 & v3a62a6d;
assign v376d45f = locked_p & v3a563ad | !locked_p & v3a70c07;
assign v3747ea2 = hbusreq5 & v3a5e496 | !hbusreq5 & v374851a;
assign v3a6fc75 = hmaster0_p & v8455b0 | !hmaster0_p & v3a59e1c;
assign v35b7771 = hmaster0_p & v377348f | !hmaster0_p & v373ef01;
assign v3771ce2 = busreq_p & v3a715fd | !busreq_p & !v3748529;
assign v3745b15 = hbusreq6_p & v3a6e699 | !hbusreq6_p & v37542af;
assign v3a67d4a = hlock0 & v3a70ad6 | !hlock0 & v3759ee4;
assign v375e577 = hbusreq2 & b3d3ad | !hbusreq2 & v3a70d64;
assign v372a347 = hlock6_p & v37604e9 | !hlock6_p & v35772a6;
assign v37585bd = hmaster1_p & v3a6fed7 | !hmaster1_p & v3a6f3f2;
assign v375e9a7 = hgrant2_p & v3758472 | !hgrant2_p & v3743c44;
assign v3746085 = hbusreq8_p & v37431c0 | !hbusreq8_p & v3732a95;
assign v376fbff = hbusreq5 & v3759b09 | !hbusreq5 & v8455ab;
assign v376fefa = hmaster2_p & v8455ab | !hmaster2_p & v3a70ab0;
assign v3744c95 = hgrant1_p & v376e139 | !hgrant1_p & v8455ab;
assign v3a6fef5 = hbusreq5_p & v3770e0e | !hbusreq5_p & v9a3ffa;
assign v3778967 = hbusreq6_p & v3751af0 | !hbusreq6_p & v377d7db;
assign v37261b2 = hbusreq8 & v1e37368 | !hbusreq8 & v3a70e37;
assign v37370c6 = hmaster2_p & v3a635ea | !hmaster2_p & v3a65762;
assign v375a235 = hgrant3_p & v8455ab | !hgrant3_p & !bdb49d;
assign v376f7a7 = hbusreq2 & v38099e8 | !hbusreq2 & v3a6c5ee;
assign v3744f80 = jx2_p & v3a6e7ae | !jx2_p & v3761aa3;
assign v3a6f4c5 = hbusreq2 & v3a58218 | !hbusreq2 & v8455ab;
assign v3a65546 = hgrant0_p & v372beb8 | !hgrant0_p & v3a5cfdb;
assign v3742aae = hlock6 & v3742290 | !hlock6 & v3a70cc2;
assign v3736012 = hlock5_p & v3a7066b | !hlock5_p & v3754a39;
assign v3725395 = hbusreq2_p & v20d166d | !hbusreq2_p & v3a6fbf7;
assign v3a676aa = hmaster2_p & v377152e | !hmaster2_p & v3756cb8;
assign v377d496 = hmaster1_p & v3778372 | !hmaster1_p & !v3a7124d;
assign v3a66460 = hbusreq1_p & b4fa3c | !hbusreq1_p & v372a201;
assign v3738944 = hmaster0_p & v2889709 | !hmaster0_p & v3761719;
assign v376faea = hmastlock_p & v37444d0 | !hmastlock_p & !v8455ab;
assign v3765a4a = hbusreq8 & v3809e72 | !hbusreq8 & v376a58a;
assign v3764f5c = hbusreq5_p & v3743a49 | !hbusreq5_p & !v8455ab;
assign v3a7113d = hbusreq8_p & v3a70578 | !hbusreq8_p & a80fe2;
assign v3726638 = hbusreq7_p & v377bac7 | !hbusreq7_p & v3a5fcf0;
assign v3a695c2 = hbusreq5 & v37738ae | !hbusreq5 & v8455ab;
assign v3a6eb6e = hbusreq4_p & v374e542 | !hbusreq4_p & v373a755;
assign v372f553 = hbusreq0 & v3726505 | !hbusreq0 & v3a7102b;
assign v3a6b8a0 = hmaster0_p & v3a706d3 | !hmaster0_p & v3a706e3;
assign v374eedb = hgrant4_p & v37541ff | !hgrant4_p & v3740b01;
assign v3a7035a = hgrant6_p & v3752a0d | !hgrant6_p & v377e9aa;
assign v3a6f48a = hmaster0_p & v375a268 | !hmaster0_p & v3756764;
assign v375c003 = hbusreq5_p & v3a5d644 | !hbusreq5_p & v3809388;
assign v3a5c50b = hbusreq0 & v3723dae | !hbusreq0 & v3a6546f;
assign v37715b9 = hbusreq7_p & v3727cec | !hbusreq7_p & v3769310;
assign v3a6bbf0 = hbusreq4 & v3772404 | !hbusreq4 & v1e378b4;
assign v373e2c3 = hbusreq2_p & v3740171 | !hbusreq2_p & v37457fb;
assign v373b295 = hbusreq4_p & v3731549 | !hbusreq4_p & v3751862;
assign v3a5a805 = hbusreq5 & v375345f | !hbusreq5 & v8455ab;
assign v3a6ab14 = hbusreq5 & v37647fc | !hbusreq5 & v3a5e030;
assign v3a70778 = hlock4_p & v374e855 | !hlock4_p & v8455cb;
assign v3744877 = hbusreq6 & v3742905 | !hbusreq6 & v373f0ee;
assign v3741d2d = hlock0_p & v3a66aa4 | !hlock0_p & v3a6fe0d;
assign v374165a = hbusreq4 & v3a6fb27 | !hbusreq4 & v8455ab;
assign v37597c4 = hmaster0_p & v373d0a3 | !hmaster0_p & v374e288;
assign v375a135 = hbusreq1_p & v3a625ee | !hbusreq1_p & !v8455ab;
assign v376d1dd = hlock5 & v3377aee | !hlock5 & v3728493;
assign v375b48b = hmaster0_p & v3a6bddf | !hmaster0_p & v8455e7;
assign v3a57ce9 = hmaster0_p & v37593cb | !hmaster0_p & v3767121;
assign v375be00 = hbusreq7_p & v37240c0 | !hbusreq7_p & v374a7f2;
assign v37419da = hbusreq8_p & v376ce90 | !hbusreq8_p & v373d142;
assign v372bbd2 = hgrant4_p & v375624b | !hgrant4_p & v3778a8b;
assign v3726f2e = hbusreq6_p & v375b2fe | !hbusreq6_p & v376dab5;
assign v3a6f448 = hbusreq5 & v374e4c5 | !hbusreq5 & !v3a6f5d4;
assign v3a705e0 = hmaster2_p & v37270d9 | !hmaster2_p & v37395e6;
assign v3751eb6 = hbusreq5 & v377fc45 | !hbusreq5 & v3a6edb5;
assign v3767a2f = hbusreq8 & v37685fe | !hbusreq8 & v8455ab;
assign v37496b5 = hbusreq6 & v3a70200 | !hbusreq6 & !v374caae;
assign v372a6c2 = hbusreq6 & v3a5c700 | !hbusreq6 & v3a70a88;
assign v37773fa = hgrant3_p & v37645ec | !hgrant3_p & v372dddc;
assign v37541d3 = hbusreq4_p & v377a551 | !hbusreq4_p & v3758700;
assign v377dadb = hmaster3_p & v375a455 | !hmaster3_p & v373f5fc;
assign v375a0b3 = hbusreq6 & v8f64f2 | !hbusreq6 & v3a56e79;
assign v375e624 = hmaster2_p & v372c5e4 | !hmaster2_p & !v8455ab;
assign v3770538 = hmaster0_p & v3724ab6 | !hmaster0_p & v373fdfb;
assign v37316b7 = hgrant3_p & v8455ab | !hgrant3_p & v375cdb1;
assign v3764a2d = hgrant4_p & v37786a6 | !hgrant4_p & v373b0d0;
assign v37332bf = hmaster1_p & v3a58fe2 | !hmaster1_p & v8455b3;
assign v3739fff = hbusreq4 & d44200 | !hbusreq4 & v374e35e;
assign v38097d8 = hlock4_p & v373aecf | !hlock4_p & v373ad95;
assign v373c8ba = hmaster0_p & v372b20b | !hmaster0_p & v23fe28c;
assign v3a7018e = hbusreq4_p & v3752fe6 | !hbusreq4_p & !v37234c3;
assign v372e537 = hmaster1_p & v37272ca | !hmaster1_p & v3726da1;
assign v3760f62 = hlock4_p & v3763fdf | !hlock4_p & v3754a27;
assign v3a6f4d0 = hgrant2_p & v3773048 | !hgrant2_p & v3761b3d;
assign v878208 = hmaster0_p & v3761d4c | !hmaster0_p & v37697ed;
assign v376fbe5 = hbusreq7_p & v3a5b819 | !hbusreq7_p & v3a71279;
assign v3a70464 = hgrant4_p & v37497dd | !hgrant4_p & v37539fc;
assign v3a5a8a4 = hbusreq5_p & v376a755 | !hbusreq5_p & v372ef17;
assign v3a66ca4 = hbusreq8_p & v37458a2 | !hbusreq8_p & v3766853;
assign v3a54b63 = hgrant4_p & v3a702c1 | !hgrant4_p & v375cd4c;
assign v3a6f9cb = hmaster2_p & v377db14 | !hmaster2_p & v3a707ce;
assign v3a70d3e = hmaster2_p & v372b780 | !hmaster2_p & v92e6f3;
assign v372ecab = hburst0 & v2aca977 | !hburst0 & v3a6ac2a;
assign v3746a81 = hmaster2_p & v1e38275 | !hmaster2_p & v3a695fc;
assign v3a5b9d6 = hmaster0_p & v8455ab | !hmaster0_p & v3771b83;
assign v3a62e01 = hgrant6_p & v8455ca | !hgrant6_p & v3a6fdf0;
assign v3a700b2 = hbusreq6 & v3a661fe | !hbusreq6 & v8455ab;
assign v375c62d = hbusreq5_p & v374ac78 | !hbusreq5_p & !v37323c5;
assign v375b342 = hmaster0_p & v374729b | !hmaster0_p & v3a6fcb6;
assign v3a70419 = hbusreq5_p & v37482bb | !hbusreq5_p & v3a56a86;
assign v3a59545 = hbusreq2 & v3806b35 | !hbusreq2 & v8455ab;
assign v3a6199f = hbusreq7 & bca64b | !hbusreq7 & !v8455c6;
assign v375e53a = hbusreq4_p & v8455ab | !hbusreq4_p & v8455c9;
assign v3a6fae5 = stateG10_1_p & v35772a5 | !stateG10_1_p & !v372e8ed;
assign v8c8903 = hlock6_p & v374306c | !hlock6_p & v3a6ffae;
assign v3753994 = hbusreq5 & v37480b3 | !hbusreq5 & v3774bad;
assign v37437cf = hbusreq5 & v3a546a2 | !hbusreq5 & v3a6f5a2;
assign v377cdea = hgrant2_p & v3808ed4 | !hgrant2_p & v37325ad;
assign v3749b84 = hgrant0_p & v3a5d48b | !hgrant0_p & v8455ab;
assign v3a6f64c = jx1_p & v373cc48 | !jx1_p & v372b46a;
assign v374474d = hmaster1_p & v377ceb5 | !hmaster1_p & v8455ab;
assign stateG2 = !v292500d;
assign v37242cb = hmaster2_p & v3757966 | !hmaster2_p & v3a5c4e8;
assign v3748f03 = hlock4 & v3a57658 | !hlock4 & v373303f;
assign v3a66a01 = hgrant4_p & v377d01e | !hgrant4_p & v3750c59;
assign v3a66737 = hbusreq0_p & v8455ab | !hbusreq0_p & v373905f;
assign v3a71394 = hmaster2_p & v3a6fdd1 | !hmaster2_p & v37306c2;
assign v3a6ef42 = hlock4_p & v372fe10 | !hlock4_p & v8455ab;
assign v3737c0a = hbusreq3 & v37401f0 | !hbusreq3 & v8455ab;
assign v373a2b4 = hlock5_p & v8455ab | !hlock5_p & v37308bc;
assign v3729f41 = hmaster2_p & v3a6d569 | !hmaster2_p & v3a6f641;
assign v37370f1 = hbusreq8_p & v3a55aea | !hbusreq8_p & v3776018;
assign v3a66f35 = hbusreq0 & v374a297 | !hbusreq0 & v377085b;
assign v374e5eb = hgrant7_p & v8455ab | !hgrant7_p & v3a70cc6;
assign v37281be = hbusreq8 & v3a704fb | !hbusreq8 & v3774f1e;
assign v376256c = hmaster0_p & v3739082 | !hmaster0_p & v376cd84;
assign v3a70f08 = hmaster2_p & v377b774 | !hmaster2_p & v3a5f0b2;
assign v372f62a = hgrant6_p & v374f511 | !hgrant6_p & v3726098;
assign v3a7150e = hbusreq2 & v374212e | !hbusreq2 & v3a708c2;
assign a72a7c = hgrant5_p & v3727d4c | !hgrant5_p & v3753fc9;
assign v3772c21 = hgrant2_p & v20930ad | !hgrant2_p & v375d4f9;
assign v3766238 = hlock0_p & v373aecf | !hlock0_p & v376430b;
assign v3740489 = hmaster1_p & v377e089 | !hmaster1_p & v377109a;
assign v3762e85 = hmaster2_p & v8455ab | !hmaster2_p & !v380760a;
assign v3a708a2 = hbusreq6 & v8455b0 | !hbusreq6 & v8455ab;
assign v376aa7a = hbusreq3 & v372d880 | !hbusreq3 & v3726006;
assign v374b0d9 = hbusreq8 & v3765433 | !hbusreq8 & v35b71fc;
assign v3743a2c = hgrant1_p & v3a6d684 | !hgrant1_p & v1e38224;
assign v3755a70 = hgrant6_p & v8455ab | !hgrant6_p & v37668cb;
assign v3770ea8 = hmaster0_p & v3a7144d | !hmaster0_p & v3760513;
assign v3a58530 = hlock2 & v377bbbb | !hlock2 & v3778251;
assign v3758dfe = hgrant3_p & v3a70ee7 | !hgrant3_p & v3a6d1a4;
assign v375ecab = hbusreq5_p & v37255f6 | !hbusreq5_p & !v3a58e44;
assign v3808904 = hgrant7_p & v3770362 | !hgrant7_p & v373a79f;
assign v377cf20 = hmaster0_p & v37737aa | !hmaster0_p & v3770ee9;
assign v3758187 = hbusreq0 & v374b9f9 | !hbusreq0 & v3a71660;
assign v376b063 = hlock7_p & v8455ab | !hlock7_p & v374be0c;
assign v9762fd = hbusreq4 & v37615aa | !hbusreq4 & v375b9c1;
assign v372886c = stateG10_1_p & v2aca977 | !stateG10_1_p & v3a6fd79;
assign v373d4a6 = hmaster2_p & v3741240 | !hmaster2_p & v3a66822;
assign v372adc8 = hbusreq6 & v376245d | !hbusreq6 & v8455ab;
assign v3770621 = hmaster2_p & v374c5b2 | !hmaster2_p & v8455bf;
assign v3a6fbe4 = hbusreq6_p & v3748e0b | !hbusreq6_p & v3762498;
assign v3a6fac0 = hgrant4_p & v37697a3 | !hgrant4_p & v377206b;
assign v375c28e = hbusreq7 & v35b86d1 | !hbusreq7 & v373264f;
assign v3a6a580 = hgrant4_p & v8455ab | !hgrant4_p & v3a6ffe7;
assign v37470e2 = hmaster2_p & v8455ab | !hmaster2_p & !v8455c2;
assign v3749106 = hgrant5_p & v3734ab5 | !hgrant5_p & v377584f;
assign v37514c2 = hmaster0_p & v3771ce2 | !hmaster0_p & v23fe295;
assign v377ecd4 = hlock4 & v38072fd | !hlock4 & v37355ce;
assign v37771e3 = hbusreq6 & v375de18 | !hbusreq6 & v8455ab;
assign v3745bbe = hmaster0_p & v8455b2 | !hmaster0_p & v3a7155c;
assign v374774d = hmaster2_p & v3762870 | !hmaster2_p & a4764c;
assign v2acaec4 = hbusreq5_p & v374156a | !hbusreq5_p & v374597c;
assign v3a70301 = hgrant5_p & v3808f5d | !hgrant5_p & v37550bd;
assign v376c235 = hgrant3_p & v3a615f7 | !hgrant3_p & v37299b3;
assign v3760b17 = hgrant6_p & v374bc10 | !hgrant6_p & v372d5bb;
assign v3a6ef8f = hgrant5_p & v8455ab | !hgrant5_p & v3a6926b;
assign v3a71558 = hgrant2_p & v8455ab | !hgrant2_p & !v3736319;
assign v3751983 = hbusreq8_p & v375515c | !hbusreq8_p & v3771182;
assign v2ff9268 = hgrant2_p & v376b5f8 | !hgrant2_p & v373243e;
assign v3772aaf = hgrant5_p & v377af89 | !hgrant5_p & v2acb0e4;
assign v3759e9d = hbusreq1 & v373fe5e | !hbusreq1 & !v376430b;
assign v3a68af5 = hbusreq8_p & v37499a4 | !hbusreq8_p & v35772a6;
assign v39eb569 = hbusreq3_p & v3a6f314 | !hbusreq3_p & v8455ab;
assign v374e019 = hmaster2_p & v3743ff2 | !hmaster2_p & v3a5c562;
assign v3a552c9 = hlock4 & v3a55f2b | !hlock4 & v37413b6;
assign v376ca93 = hbusreq6 & v3a71314 | !hbusreq6 & v8455ab;
assign v37509c7 = hgrant0_p & v37773a9 | !hgrant0_p & v375e309;
assign v3744539 = hbusreq8 & v3a65c81 | !hbusreq8 & v3a67beb;
assign v3809eab = hmaster2_p & v3a633ac | !hmaster2_p & v8455ab;
assign v376af8d = hmaster0_p & v3769c47 | !hmaster0_p & v3770fef;
assign v3a550e2 = hmaster1_p & v373e873 | !hmaster1_p & v3a683c6;
assign v3a5cca9 = jx0_p & v3a653d5 | !jx0_p & v375994d;
assign v8ad83a = hbusreq6_p & v3a5a397 | !hbusreq6_p & v3742eaf;
assign v3a56512 = hmaster2_p & v372c007 | !hmaster2_p & v3a56e63;
assign v3728203 = hbusreq5_p & v3a6d7cd | !hbusreq5_p & v3a6fb1b;
assign v3760aa7 = hbusreq6_p & v3737c86 | !hbusreq6_p & v37474e8;
assign v372bfd0 = hmaster0_p & v28896b4 | !hmaster0_p & v3a6f871;
assign v372570c = hbusreq6_p & v3769010 | !hbusreq6_p & v3722bc2;
assign v377ed8c = hgrant1_p & v8455b6 | !hgrant1_p & !v8455b0;
assign v375fdc9 = hmaster2_p & v3753d94 | !hmaster2_p & v3a70384;
assign v3722f50 = jx0_p & v3740247 | !jx0_p & v376a74a;
assign v3a700b9 = hmaster1_p & v3a70641 | !hmaster1_p & v375d889;
assign d5c12b = jx1_p & v375d85b | !jx1_p & v8455ab;
assign v3a701c7 = hbusreq4 & v38090e9 | !hbusreq4 & v8455ab;
assign v3a71264 = hmaster1_p & v377e056 | !hmaster1_p & v3a70859;
assign v373b9a9 = hbusreq3 & v3a6469c | !hbusreq3 & v1e37c3e;
assign v3739021 = hbusreq3 & v37457fb | !hbusreq3 & v8455ab;
assign v374366a = hmaster1_p & v3747554 | !hmaster1_p & v374e86a;
assign v375a858 = hmaster0_p & v375787b | !hmaster0_p & v373ca5f;
assign v373040e = hbusreq0_p & v8a7f7e | !hbusreq0_p & v3a70bce;
assign v3809968 = hmaster0_p & v372301d | !hmaster0_p & v376a094;
assign v3a69239 = hbusreq7_p & v37374e5 | !hbusreq7_p & !v3766852;
assign v3763364 = hmaster0_p & v3a61a7f | !hmaster0_p & v3a702bd;
assign v3808c89 = hbusreq7_p & v3738b7e | !hbusreq7_p & !v3726ed7;
assign v37624a5 = hlock5_p & v3a60836 | !hlock5_p & !v3775c51;
assign bb4062 = hmaster2_p & v375d263 | !hmaster2_p & v373891b;
assign v377c185 = hgrant0_p & v374c01f | !hgrant0_p & v3a7168a;
assign v376d52a = hmaster1_p & v376501e | !hmaster1_p & v375e06b;
assign v372cd7e = hready_p & v3751a4f | !hready_p & v3793188;
assign v3753055 = hmaster2_p & v372976e | !hmaster2_p & v3772608;
assign v3a68a8b = hmaster0_p & v3770f96 | !hmaster0_p & v377346e;
assign v3a6a5a8 = hgrant5_p & v8455ab | !hgrant5_p & v3a29850;
assign v37702f3 = hmaster0_p & v3a5ade4 | !hmaster0_p & v37654c4;
assign v3753a1d = hbusreq5 & v3728eca | !hbusreq5 & v3a6f9ce;
assign v3a5e0b8 = hmaster0_p & v3a6fb37 | !hmaster0_p & v377fad8;
assign v3747178 = hgrant6_p & v37517d2 | !hgrant6_p & !v3a7030f;
assign v3a59158 = hbusreq4 & v375b64b | !hbusreq4 & v8455ab;
assign v3a63699 = hmaster0_p & v8637a5 | !hmaster0_p & v8455ab;
assign v3728f64 = hbusreq2 & v377ba55 | !hbusreq2 & v3724940;
assign v37318e3 = hmaster0_p & v376b65a | !hmaster0_p & v3733d02;
assign v377e8ca = hgrant6_p & v8455ab | !hgrant6_p & v3770173;
assign v3a7161f = hmaster2_p & v3746c51 | !hmaster2_p & v373cd16;
assign v2925cf2 = hlock5 & v377600d | !hlock5 & v3725b77;
assign v3a6f61a = hbusreq5 & v37599a4 | !hbusreq5 & !v377cc7b;
assign v38069c8 = hlock5_p & v8455ab | !hlock5_p & v374f8da;
assign v3753825 = hmaster2_p & v3753dab | !hmaster2_p & v3753329;
assign v373ac52 = hbusreq2 & v3a6f018 | !hbusreq2 & !v3a5db8a;
assign v3a62f50 = hmaster0_p & v3a62113 | !hmaster0_p & v3a71202;
assign b2ea29 = hmaster2_p & v3a70f8f | !hmaster2_p & v372912f;
assign v377982c = hmaster2_p & v377ca49 | !hmaster2_p & v3764418;
assign v376fc80 = hbusreq5 & v3775f56 | !hbusreq5 & !v3a5fc70;
assign v3a585f1 = hmaster1_p & v3739112 | !hmaster1_p & v3a6f2ce;
assign v377086c = hmaster0_p & v3a65c2c | !hmaster0_p & v373594b;
assign v3778c14 = hbusreq5_p & v377ef71 | !hbusreq5_p & v3a70f27;
assign v377c06f = hmaster3_p & v376b14c | !hmaster3_p & v3743eed;
assign v3a57ad0 = hgrant2_p & v3a5f50e | !hgrant2_p & v377613d;
assign v376d05f = hlock4 & v377d6d3 | !hlock4 & v376b57f;
assign v373ce2b = hmaster0_p & v3a58a34 | !hmaster0_p & v376bae4;
assign v374b27d = hbusreq6_p & v377b24b | !hbusreq6_p & v372be8e;
assign v3763e76 = hbusreq0 & v2092bcb | !hbusreq0 & v374e085;
assign v3749a89 = hlock3_p & v373c151 | !hlock3_p & !v8455ab;
assign v375e217 = hmaster2_p & v8455ab | !hmaster2_p & !v374044c;
assign v3754f0f = hgrant6_p & v377bd79 | !hgrant6_p & v3746e47;
assign v3a56417 = hbusreq1_p & v3a6f1c6 | !hbusreq1_p & !v8455ab;
assign v3a70827 = hbusreq4_p & v373552a | !hbusreq4_p & v3a5dd1a;
assign v3755f4a = hgrant6_p & v377f09a | !hgrant6_p & !v373f224;
assign v3746145 = hlock2 & v3258db3 | !hlock2 & v3a5eafa;
assign v3a53dfc = hlock7_p & v3a6a0c4 | !hlock7_p & !v3739e0e;
assign v3778a8b = hbusreq4_p & v3726d1f | !hbusreq4_p & v3a64aa0;
assign v3773e8d = hmaster1_p & v3a63777 | !hmaster1_p & v374e016;
assign v3723ac4 = hmaster0_p & v3a5a807 | !hmaster0_p & v2ff8e8b;
assign v3a71002 = hmaster0_p & v3743ff2 | !hmaster0_p & v3774492;
assign v39372d9 = hbusreq5 & v3a62d5d | !hbusreq5 & v3740c5f;
assign v374b564 = hlock5 & v376cd09 | !hlock5 & v376c422;
assign v372f74f = hlock6_p & v8455ab | !hlock6_p & v3a601a0;
assign v3a6f900 = jx0_p & v376cc0e | !jx0_p & v373b4c8;
assign v3759b20 = hbusreq5_p & v373efee | !hbusreq5_p & v8455ab;
assign v3777311 = hbusreq3_p & v3778834 | !hbusreq3_p & v8455ab;
assign v3724014 = hmaster1_p & v3731724 | !hmaster1_p & v3735bbb;
assign v374d490 = hbusreq5 & v372f2ae | !hbusreq5 & v3734331;
assign v3736b19 = hmaster0_p & v373a4e4 | !hmaster0_p & v376d7a5;
assign v3a70ee7 = hlock0_p & v3a5891c | !hlock0_p & v3759032;
assign v3773a00 = hmaster0_p & v8455ab | !hmaster0_p & v3747238;
assign v37557c6 = hlock7 & v3a6fd41 | !hlock7 & v3a5f458;
assign v376382f = hgrant5_p & v376934b | !hgrant5_p & v373c334;
assign v3748494 = hlock8 & v3729a07 | !hlock8 & v375f2c7;
assign v3a6abe5 = hbusreq4 & v3a6a939 | !hbusreq4 & v8455ab;
assign v3734279 = hmaster1_p & v377de7f | !hmaster1_p & v8455ab;
assign v37676dc = hmaster2_p & v372433d | !hmaster2_p & v3753ccf;
assign v374e168 = hmaster0_p & v3750f60 | !hmaster0_p & !v373ad3f;
assign v3735e52 = hlock5 & v377de7f | !hlock5 & v3a701b1;
assign v3735468 = hgrant8_p & v374ef8d | !hgrant8_p & v37472b6;
assign v3a70f14 = hbusreq6_p & v3a64252 | !hbusreq6_p & v374ec22;
assign v3a71527 = hbusreq4 & v3a70006 | !hbusreq4 & !v8455ab;
assign v3751d16 = hlock4_p & v3732415 | !hlock4_p & v3a5e7fe;
assign v375fbb7 = hbusreq6 & v37616e0 | !hbusreq6 & v3a6ebcc;
assign v3731a49 = hgrant4_p & v373ff91 | !hgrant4_p & v372f5ec;
assign v372a939 = hgrant6_p & v8455ab | !hgrant6_p & v3774c77;
assign v3a7131c = hbusreq4 & v3a63dbb | !hbusreq4 & v8455ab;
assign v3755af9 = hmaster0_p & v374571a | !hmaster0_p & v375355a;
assign v3a5a28b = hmaster2_p & v376f569 | !hmaster2_p & v3751510;
assign v375afe9 = hgrant4_p & v376a6f1 | !hgrant4_p & v3765576;
assign v3a6184c = hlock5_p & v3753fb7 | !hlock5_p & !v3750e0b;
assign v377c4bf = hlock7_p & v373651a | !hlock7_p & v377c9f3;
assign v376ef7a = hlock6_p & v3773ee6 | !hlock6_p & v8455b3;
assign v2092f41 = hbusreq4 & v3a65da7 | !hbusreq4 & v8455bb;
assign v3a70e37 = hmaster1_p & v374e855 | !hmaster1_p & v3758a7c;
assign v3a60924 = hmaster0_p & v3a7116a | !hmaster0_p & v374476d;
assign v3a71112 = hgrant7_p & v37283ea | !hgrant7_p & v37279df;
assign cd348d = hbusreq2 & v37234f5 | !hbusreq2 & !v8455ab;
assign v35b6167 = decide_p & v3a6f3d6 | !decide_p & v3757047;
assign v37566a2 = hgrant3_p & v3776c43 | !hgrant3_p & v37293b1;
assign v3a70abd = jx1_p & v37291e4 | !jx1_p & v3a700d0;
assign v376c17d = hgrant5_p & v3754086 | !hgrant5_p & v377a4e5;
assign v377664f = hbusreq7 & v3a70194 | !hbusreq7 & v377b735;
assign v3759fd0 = hmaster2_p & v3760513 | !hmaster2_p & v3736cb3;
assign v375b9b0 = hbusreq5_p & v3756d57 | !hbusreq5_p & v8455ab;
assign v3806ce9 = hbusreq4 & v3767f52 | !hbusreq4 & v3a56049;
assign v376bc6a = hbusreq6 & v3a6a939 | !hbusreq6 & v8455ab;
assign v372ef7c = hbusreq1 & v3a6ab5f | !hbusreq1 & !v2acb5a2;
assign v3773633 = hmaster0_p & v3a624e7 | !hmaster0_p & v3769923;
assign v3a6f764 = hbusreq2 & v3a703ad | !hbusreq2 & v8455ab;
assign v3726277 = hgrant1_p & v374306c | !hgrant1_p & v3751fa8;
assign v373c5b5 = hmaster1_p & v373aa91 | !hmaster1_p & v3a6fef5;
assign v3a6b288 = hmaster1_p & v8455ab | !hmaster1_p & v3a5b0a6;
assign v377a36e = hlock6_p & v8455ab | !hlock6_p & v3a70cc0;
assign dc6ab1 = hmaster3_p & v8455ab | !hmaster3_p & a0a219;
assign v37681a3 = hlock5 & v37261ad | !hlock5 & v37785f8;
assign v3a5e91b = hbusreq3 & v373d7fe | !hbusreq3 & v8455ab;
assign v375d34f = hbusreq8_p & v3753f71 | !hbusreq8_p & v375e3a5;
assign v3a6fb85 = hmaster0_p & v8455dd | !hmaster0_p & v8455ab;
assign v375a52a = hbusreq3_p & v373db5d | !hbusreq3_p & v8455ab;
assign v372cdc9 = hgrant2_p & v8455ab | !hgrant2_p & v3a6c390;
assign v3777412 = hbusreq2 & v3a6f7bf | !hbusreq2 & v8455ab;
assign v376f542 = hlock6_p & v2acb5a2 | !hlock6_p & v3a6ac2a;
assign v372a478 = hmaster3_p & v3a6cac4 | !hmaster3_p & v3a709c2;
assign bfa92a = hbusreq8 & v3a7151f | !hbusreq8 & v372cf51;
assign v375c3c5 = hlock7 & v3728990 | !hlock7 & v372af95;
assign v3a63ea7 = hlock2_p & v3763175 | !hlock2_p & !v8455ab;
assign v375478f = hmaster1_p & v8455ab | !hmaster1_p & v377de7f;
assign v3727a2f = hmaster2_p & v374449e | !hmaster2_p & v37615ce;
assign v3756d28 = hmaster2_p & v325c960 | !hmaster2_p & v37422f3;
assign v3778454 = hbusreq4 & v374d28d | !hbusreq4 & v3a6bf41;
assign v3765699 = hgrant6_p & v376d882 | !hgrant6_p & !v3a682a1;
assign v37791a5 = hgrant4_p & v8455ab | !hgrant4_p & v372e3ea;
assign v3758f94 = hgrant6_p & v3726be0 | !hgrant6_p & v3745df8;
assign v3a5a798 = hgrant0_p & v3765b30 | !hgrant0_p & !v3750d06;
assign v3731fb9 = hbusreq5 & v3777362 | !hbusreq5 & v3a656a4;
assign v37448f2 = hbusreq2 & v3771c59 | !hbusreq2 & d1bf3b;
assign v3728990 = hbusreq7 & v377a3af | !hbusreq7 & v3a6b303;
assign v373a2cc = jx1_p & v375d1e1 | !jx1_p & v8455ab;
assign v3a65d33 = hmaster0_p & v37793a6 | !hmaster0_p & v3775100;
assign v3775ca5 = locked_p & v37481c3 | !locked_p & v8455ab;
assign v3771fb7 = hmaster2_p & v377f526 | !hmaster2_p & v3769374;
assign v3a5f7f3 = hlock3 & v3a70910 | !hlock3 & v3733cca;
assign v377d8dd = hbusreq1_p & v372dec8 | !hbusreq1_p & v3732b98;
assign c58ea1 = hgrant3_p & v3a712e6 | !hgrant3_p & !v3a6efd1;
assign v3a70029 = hmaster2_p & v3a6a3e6 | !hmaster2_p & v37514c7;
assign v375881d = hmaster2_p & v3a70ed7 | !hmaster2_p & v37351f5;
assign v3a6ff80 = hlock4_p & v37625a8 | !hlock4_p & v3a5ace5;
assign v37691e2 = hmaster2_p & v3a62ad5 | !hmaster2_p & v3742953;
assign v3a6a0aa = hbusreq4_p & v3724c25 | !hbusreq4_p & v3a66273;
assign v37268cc = hmaster2_p & v37342f2 | !hmaster2_p & v3741906;
assign v377640c = hbusreq0 & v37724db | !hbusreq0 & v3750f49;
assign v3a6802f = hmaster0_p & v3779183 | !hmaster0_p & d1e3dd;
assign v3a59720 = hbusreq1_p & v3a70d65 | !hbusreq1_p & !v3737f5f;
assign v372f4e6 = hlock5 & v372a39a | !hlock5 & v376430d;
assign v374fb02 = hmaster0_p & v3a66110 | !hmaster0_p & v377f505;
assign v372c5bc = hbusreq7 & v3a6ff9a | !hbusreq7 & v3749503;
assign v37280f3 = hmaster2_p & v8455ab | !hmaster2_p & !v374e0f6;
assign v37544fa = hgrant0_p & v8455ab | !hgrant0_p & v3a67370;
assign v3763898 = hgrant2_p & v8455ab | !hgrant2_p & v376c12e;
assign v3a7166a = hmaster1_p & v3a66232 | !hmaster1_p & v3a53ce6;
assign v3a555e5 = hgrant5_p & v3808d74 | !hgrant5_p & v376ce59;
assign v3a6a7a1 = hbusreq1_p & v3a6fc6c | !hbusreq1_p & v37616e1;
assign v3806df2 = hlock7 & v3a54d25 | !hlock7 & v3a70129;
assign v372dadb = hbusreq1_p & v372e8ed | !hbusreq1_p & !v3a6fae5;
assign v373e944 = hmaster0_p & v3a70987 | !hmaster0_p & v377e6fc;
assign v3758cec = hbusreq1_p & v8455e7 | !hbusreq1_p & v8455ab;
assign v3764a6c = hmaster2_p & v3a6ff99 | !hmaster2_p & v3756304;
assign v23fe324 = hgrant4_p & v37665e2 | !hgrant4_p & v372b24d;
assign v3a6f6fa = hgrant3_p & v8455ab | !hgrant3_p & v373abbe;
assign v3757188 = hmaster0_p & v3a70f68 | !hmaster0_p & v3745cc6;
assign v3a5c3ef = hmaster0_p & v3a61a7f | !hmaster0_p & v3a2a0f9;
assign v3a61d77 = hbusreq4_p & v374525d | !hbusreq4_p & v373abde;
assign v3a5e4e5 = hmaster0_p & v3a62965 | !hmaster0_p & v373185b;
assign v3a669e9 = hmaster2_p & v374dc13 | !hmaster2_p & v3733440;
assign v3760233 = hlock7_p & v374361e | !hlock7_p & v3764238;
assign v372c064 = hmaster2_p & v3754b66 | !hmaster2_p & v8455b2;
assign v3a6fc81 = hbusreq8_p & v37784a9 | !hbusreq8_p & v3a6d80d;
assign v3735179 = hgrant2_p & v3a6eb39 | !hgrant2_p & v37483db;
assign v376926f = hbusreq4_p & v3a5841e | !hbusreq4_p & v8455ab;
assign v37375ed = hgrant5_p & v376219d | !hgrant5_p & v3a709b5;
assign v37428ac = hgrant4_p & v3a5c58f | !hgrant4_p & v8455ab;
assign v373facf = hbusreq0 & v37512dc | !hbusreq0 & v375dba4;
assign v3a6f5e7 = jx0_p & v376b56b | !jx0_p & v3764f2d;
assign v37295ce = hlock5_p & v3a70fe6 | !hlock5_p & v3a6eff3;
assign v3808ed2 = locked_p & v3a70521 | !locked_p & v3a6e7b3;
assign v37648af = hbusreq3_p & v8455ab | !hbusreq3_p & v374fb58;
assign v3763c09 = hbusreq4_p & v37721df | !hbusreq4_p & !v8455ab;
assign v376c789 = hbusreq5 & v3750d19 | !hbusreq5 & v3809f0e;
assign v376984f = hbusreq5_p & v3729f7b | !hbusreq5_p & v3769740;
assign v372f91d = hbusreq0 & v3732246 | !hbusreq0 & v3758a10;
assign v3a60a68 = hbusreq6_p & v3a635ea | !hbusreq6_p & v373b288;
assign v3a6fd82 = hgrant3_p & v37c1a6f | !hgrant3_p & v373ee70;
assign v3a59819 = hmaster2_p & v3a70fb2 | !hmaster2_p & v3752e63;
assign v3727ad4 = hgrant4_p & v8455ab | !hgrant4_p & v3a70308;
assign v3a6db06 = hbusreq2_p & v3737ca3 | !hbusreq2_p & v3a5afe8;
assign v377a6ce = hbusreq3 & v375de18 | !hbusreq3 & !v373c755;
assign v373c7db = hbusreq4 & v3729b6a | !hbusreq4 & v3a6403e;
assign v377c3f5 = hlock7_p & v376d007 | !hlock7_p & !v8455ab;
assign v3a71085 = hmastlock_p & v37524c6 | !hmastlock_p & !v8455ab;
assign v377f64b = hmaster0_p & v37737aa | !hmaster0_p & v373eff1;
assign v3730b77 = hbusreq2_p & v377005e | !hbusreq2_p & v3754f54;
assign v3a71439 = hmaster2_p & v3769093 | !hmaster2_p & v3a70a5c;
assign v375b626 = hbusreq4_p & v3777ce4 | !hbusreq4_p & v376871e;
assign v3779491 = hmaster0_p & v3a6f781 | !hmaster0_p & v376c854;
assign v377ce1a = hbusreq4 & v3a6e5f0 | !hbusreq4 & v8455ab;
assign v375c111 = hlock8 & v3746df7 | !hlock8 & v373c7aa;
assign v3741e54 = hgrant4_p & v8455e7 | !hgrant4_p & !v3775269;
assign v3a6b864 = hmaster3_p & v373fe61 | !hmaster3_p & v3745ae6;
assign v3a702c5 = hmaster0_p & v375a500 | !hmaster0_p & v377402f;
assign v3724cce = hmaster1_p & v3735c84 | !hmaster1_p & v3a5d3f6;
assign v3769a16 = hmaster1_p & v3a6efe8 | !hmaster1_p & v374d01c;
assign v337905c = hbusreq5_p & v374851a | !hbusreq5_p & v37790c8;
assign v3749242 = hbusreq5 & v3a6fd12 | !hbusreq5 & v3724060;
assign v3761cd2 = hlock5 & v3a6275e | !hlock5 & v374ad45;
assign v3739246 = hgrant8_p & v8455d2 | !hgrant8_p & v3747c9f;
assign v372cea0 = hmaster2_p & v3a635ea | !hmaster2_p & v3a6e6fa;
assign v377ac8a = hbusreq3 & v3a6f757 | !hbusreq3 & v3a635ea;
assign v37254d2 = hgrant6_p & v8455ab | !hgrant6_p & v372d96e;
assign v3a704f2 = hbusreq6 & v3a6fa2c | !hbusreq6 & v3a6fdef;
assign v377498e = hbusreq4_p & v375aafe | !hbusreq4_p & !v3727976;
assign v3774737 = hmaster2_p & v375a52a | !hmaster2_p & v8455bf;
assign v3770331 = hmaster2_p & v3761b5e | !hmaster2_p & v35772a6;
assign v3742395 = hlock8 & v3807748 | !hlock8 & v3a5bc76;
assign v374d2d5 = hmaster2_p & v3a635ea | !hmaster2_p & v377b330;
assign v37731d8 = hmaster2_p & v8455ab | !hmaster2_p & v37271e7;
assign v3769cd7 = hgrant4_p & v8455ab | !hgrant4_p & v376ee7c;
assign v3761ac9 = hbusreq7_p & v372706f | !hbusreq7_p & v37626ae;
assign v37343bc = hgrant4_p & v3768857 | !hgrant4_p & v3777bf9;
assign v37649ab = hbusreq3_p & v3a6ebbc | !hbusreq3_p & v3732302;
assign v3a6f374 = hbusreq0 & v3a5334f | !hbusreq0 & v1e37cd6;
assign v37435e9 = hbusreq5_p & v3728a45 | !hbusreq5_p & v37313fa;
assign v3743017 = hbusreq5_p & v3777647 | !hbusreq5_p & v3746a67;
assign v3744efc = hmaster0_p & d58c24 | !hmaster0_p & v3a6af83;
assign v372e77b = hmaster1_p & v3757568 | !hmaster1_p & v3723a30;
assign v3742f64 = hbusreq4_p & v3754b66 | !hbusreq4_p & v3728d14;
assign v3768d8f = hbusreq7_p & v3a70428 | !hbusreq7_p & v374b8fe;
assign v3a6ef89 = hbusreq2_p & v3763344 | !hbusreq2_p & v8455ab;
assign v3a6cbfa = hmaster1_p & v39ea76e | !hmaster1_p & v3a5be0b;
assign v374d1dc = hmaster2_p & v372625f | !hmaster2_p & v37297d0;
assign v373bf4f = hbusreq6 & v3778fec | !hbusreq6 & v3762502;
assign v3a5de35 = hgrant6_p & v37395e8 | !hgrant6_p & v373c628;
assign v372b4b4 = hbusreq5 & v372c0d6 | !hbusreq5 & v3a6c0ba;
assign v38092a9 = hmaster1_p & v3a65e9d | !hmaster1_p & c46b05;
assign v374bf93 = hgrant5_p & v373e743 | !hgrant5_p & v3764983;
assign v374182b = hmaster2_p & v3a700e2 | !hmaster2_p & v8455ab;
assign v37667ed = hmaster2_p & v3a69591 | !hmaster2_p & !v37598ab;
assign v377d23d = hbusreq7 & v3a5bfbd | !hbusreq7 & v3749ca6;
assign v3761c61 = hmaster2_p & v3a6ff32 | !hmaster2_p & v8455ab;
assign v3a5e10c = hgrant6_p & v3a6fd6a | !hgrant6_p & v3a60fd6;
assign v375e8d9 = hmaster0_p & v373f9bf | !hmaster0_p & v3a710c3;
assign cc8b5a = hbusreq5 & v3769c6d | !hbusreq5 & v377234d;
assign v3a709db = hbusreq8_p & v3730a22 | !hbusreq8_p & v3734473;
assign v377d45b = hgrant7_p & v3770648 | !hgrant7_p & v374f273;
assign v3a5b6a3 = hbusreq8 & v3a5f51c | !hbusreq8 & v3a70e3c;
assign v3a6f073 = hmaster2_p & v3a6f942 | !hmaster2_p & v376d268;
assign v3a7030f = hgrant2_p & v8455e7 | !hgrant2_p & !v3a63329;
assign v3753d60 = hbusreq3_p & v8455b7 | !hbusreq3_p & v3a61c5a;
assign v3753073 = hlock4 & v3a6ed4c | !hlock4 & v376f0a0;
assign v376cdf6 = hbusreq0 & v3748f33 | !hbusreq0 & !v1e37cd6;
assign v3a54478 = hmaster0_p & v372d727 | !hmaster0_p & v3a70aef;
assign v3a676f1 = hgrant5_p & v375d23b | !hgrant5_p & v3a6f891;
assign v373b203 = hmaster2_p & v372d299 | !hmaster2_p & v37512ca;
assign v37607c6 = jx0_p & v3a6471e | !jx0_p & v3a70816;
assign v377e639 = hgrant6_p & v8455ab | !hgrant6_p & v35b9d5e;
assign v3a6f226 = hbusreq8 & v3737711 | !hbusreq8 & v376e9ed;
assign v3732b81 = hlock3 & v3a70ea0 | !hlock3 & v3760e47;
assign b65b94 = hbusreq0 & v3a70532 | !hbusreq0 & v3728a76;
assign v3768ed2 = hmaster1_p & v3a6fe0d | !hmaster1_p & v3763f30;
assign v3775806 = hgrant5_p & v8455ab | !hgrant5_p & v3731312;
assign v3a6177b = hmaster1_p & v3a661fe | !hmaster1_p & v3774c25;
assign v3a7024f = hbusreq0 & v375491e | !hbusreq0 & v372e3f5;
assign v3a5b89a = hbusreq5 & v3a7017d | !hbusreq5 & v3a6fd98;
assign v3a6ef17 = hbusreq5 & v372b50b | !hbusreq5 & v372a0e3;
assign v3a5815e = busreq_p & v3a70b53 | !busreq_p & v3a5e0cc;
assign v3773d27 = hmaster0_p & v3747130 | !hmaster0_p & v3768495;
assign v3743094 = hmaster0_p & v3755774 | !hmaster0_p & b0e59c;
assign v3a701c2 = hgrant6_p & v374fa4c | !hgrant6_p & v3a64252;
assign v3759ad6 = hmaster2_p & v3732dac | !hmaster2_p & v373a415;
assign v3726379 = hmaster0_p & v3a6eb6a | !hmaster0_p & v3750088;
assign v375c98d = hbusreq0 & v2acaed3 | !hbusreq0 & v3779c2b;
assign v37308b0 = hgrant2_p & v8455ab | !hgrant2_p & !v3a6d621;
assign v3a5be41 = hmaster0_p & v3771d75 | !hmaster0_p & v3a7026a;
assign d62aa6 = hmaster1_p & v8455ab | !hmaster1_p & v372790e;
assign v375538a = hgrant2_p & v3770559 | !hgrant2_p & v374d552;
assign v3a617fa = stateA1_p & v8455ab | !stateA1_p & !v3a65206;
assign v374052a = hbusreq4 & v375179a | !hbusreq4 & v8455ab;
assign v3a62c46 = hmaster0_p & v3778ac5 | !hmaster0_p & v376ef9f;
assign v3a6eb9e = hgrant5_p & v3a6fc07 | !hgrant5_p & v3a70656;
assign v3766a28 = hbusreq6 & v3a6fbd0 | !hbusreq6 & !v3a683e2;
assign v3722fb7 = hmaster1_p & v3764dac | !hmaster1_p & v3a5e030;
assign v376f499 = hlock5 & v37499a0 | !hlock5 & v32574c7;
assign v377f170 = hmaster2_p & v37367a0 | !hmaster2_p & !v3739ab6;
assign v3a6f387 = hmaster0_p & v3746496 | !hmaster0_p & v374f6f9;
assign v3735274 = hmaster0_p & v3a6dc83 | !hmaster0_p & v37466b7;
assign v373ca1a = hlock0 & v376e041 | !hlock0 & v3a6f9c7;
assign v373b2ba = hbusreq5_p & v37781d4 | !hbusreq5_p & !v8455ab;
assign d0e017 = hmaster0_p & v3a6a8c0 | !hmaster0_p & v3730a61;
assign v3a715c3 = hmaster2_p & v375a6a7 | !hmaster2_p & v374f968;
assign v372facf = jx0_p & v3a673fa | !jx0_p & v374aa0f;
assign v3759263 = hmaster0_p & v3a60a6e | !hmaster0_p & v37614c1;
assign v3a70e9a = hbusreq1 & v3749cea | !hbusreq1 & v8455ab;
assign v3738877 = hgrant6_p & v3775b4d | !hgrant6_p & v3734e58;
assign v3a62b5f = hgrant4_p & v8455ab | !hgrant4_p & !v37781b8;
assign v3756205 = hbusreq0 & v377cdbe | !hbusreq0 & v3724667;
assign v3755ad5 = hbusreq4_p & v3758d18 | !hbusreq4_p & v8455ab;
assign v374d042 = hmaster0_p & v3753418 | !hmaster0_p & v3a5c9d7;
assign v23fde61 = hbusreq5 & v374ad5f | !hbusreq5 & v3722e04;
assign v375089b = hbusreq7_p & v3776fec | !hbusreq7_p & v3a5646d;
assign v3a6fcd3 = hlock4_p & v3a70385 | !hlock4_p & !v8455ab;
assign v377d302 = hbusreq5 & v3764306 | !hbusreq5 & v374930c;
assign v37651e0 = hmaster2_p & v3a653e4 | !hmaster2_p & !v37346be;
assign v3771df4 = hbusreq8 & v8455e7 | !hbusreq8 & v377bde3;
assign v37345f3 = hbusreq3_p & v9d7b97 | !hbusreq3_p & v35772a6;
assign v3768737 = hbusreq8 & v37513e6 | !hbusreq8 & v3743a4c;
assign v3a6f523 = hmaster3_p & v3a5d94f | !hmaster3_p & !v373e121;
assign v3726c47 = hmaster1_p & v3a565a1 | !hmaster1_p & v8455ab;
assign v374e34f = hmaster0_p & v1e382c4 | !hmaster0_p & c3f48e;
assign v3a67d59 = hgrant3_p & v3764d17 | !hgrant3_p & !v3a6c0e4;
assign v3a6fa15 = hbusreq2 & v3a5e81d | !hbusreq2 & v8455ab;
assign v3741f5e = hgrant6_p & v377f09a | !hgrant6_p & !v377af34;
assign v37289bb = hmaster1_p & v3a7169d | !hmaster1_p & v372690e;
assign v3768870 = hlock6 & v373f7b7 | !hlock6 & v377b84e;
assign v37435b9 = hlock8 & v376ae9f | !hlock8 & v376f0cd;
assign v37377d2 = hbusreq5_p & v3770a5b | !hbusreq5_p & v376360a;
assign v3768889 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f8cc;
assign v375bb51 = hbusreq4_p & v373cf9c | !hbusreq4_p & v373b288;
assign v377a3da = hgrant4_p & v8455ab | !hgrant4_p & be9654;
assign cc2999 = hmaster0_p & v372ed51 | !hmaster0_p & v377d142;
assign v3a5b563 = hbusreq1_p & v3a635ea | !hbusreq1_p & v3a55271;
assign v3a70225 = hbusreq5_p & v3739120 | !hbusreq5_p & v35772a6;
assign v3a70120 = jx3_p & v375f3bc | !jx3_p & v3763f1d;
assign v3742e40 = hlock5_p & v3a6eb0e | !hlock5_p & !v8455ab;
assign v373d791 = hgrant4_p & v3748797 | !hgrant4_p & v8455ab;
assign v372d9b0 = hbusreq0 & b95629 | !hbusreq0 & v37612d4;
assign v3769af4 = hlock5_p & v8455ab | !hlock5_p & v3a67471;
assign v39ed7e6 = hgrant6_p & v3a6dae2 | !hgrant6_p & v3a70788;
assign v3736026 = hgrant4_p & v376ce77 | !hgrant4_p & v37759e3;
assign v3a61c41 = hlock0_p & v95d97e | !hlock0_p & !v2aca977;
assign v3a6f5fe = hgrant6_p & v8455c9 | !hgrant6_p & v3a70e62;
assign v377af60 = hbusreq5_p & v3a5b20c | !hbusreq5_p & a9ca33;
assign v3a6ec28 = hbusreq7 & v3726e7b | !hbusreq7 & v373e2b7;
assign v375aafe = hbusreq4 & v3809ebc | !hbusreq4 & v3738510;
assign v37546a9 = hbusreq5_p & v3741a07 | !hbusreq5_p & v3731508;
assign v3771f50 = hmaster1_p & v3a6f5bf | !hmaster1_p & v8455ab;
assign v3a5d36a = hgrant4_p & v8455ab | !hgrant4_p & v3a6bf89;
assign v374e28f = hbusreq2_p & v3a70319 | !hbusreq2_p & !v8455ab;
assign v3a675df = hmaster2_p & v375571d | !hmaster2_p & v8455e7;
assign v375297d = hlock0_p & v3a7136f | !hlock0_p & !v8455ab;
assign v372d6fa = hlock8_p & v3769712 | !hlock8_p & !v3749a7c;
assign v3730e71 = hbusreq1 & v376a14f | !hbusreq1 & v8455ab;
assign v3a6fe59 = hmaster0_p & v3732d0f | !hmaster0_p & v8455ab;
assign v374af0d = hlock3_p & v8455ab | !hlock3_p & v375338a;
assign v37330d6 = hgrant8_p & v8455ab | !hgrant8_p & !v8455f7;
assign v3a6fff6 = hbusreq3_p & v37655d6 | !hbusreq3_p & v3a70547;
assign v373f47b = hmaster0_p & v3a57584 | !hmaster0_p & v3763055;
assign v3728a3d = hmaster0_p & v3a6c8c0 | !hmaster0_p & v3a70574;
assign v373bf6a = hbusreq4_p & v377eb2d | !hbusreq4_p & v8455b0;
assign v373bbce = hbusreq7 & v3a70b61 | !hbusreq7 & v8455ab;
assign v377a461 = hbusreq6 & v3a6f68f | !hbusreq6 & v8455ab;
assign v377afb7 = hmaster1_p & v3755002 | !hmaster1_p & v3a70427;
assign v3778bde = hgrant4_p & v8455ab | !hgrant4_p & v3a6f044;
assign v37542b2 = hmaster1_p & v3a5a801 | !hmaster1_p & v3a6c8e4;
assign v3758c35 = hbusreq3_p & c22b44 | !hbusreq3_p & v377bdbe;
assign v372ddde = hmaster2_p & v37784b9 | !hmaster2_p & v3770bd5;
assign v373a1dc = hbusreq5_p & v3a6f6cb | !hbusreq5_p & v8455ab;
assign v377204f = hbusreq0 & v373d8f2 | !hbusreq0 & v3a710d9;
assign v376b21a = hbusreq3_p & v39a537f | !hbusreq3_p & !v39a5381;
assign v3764daf = hbusreq5_p & v3747de2 | !hbusreq5_p & v3a614fe;
assign v3a70d88 = hmaster3_p & v3a56b80 | !hmaster3_p & !v3740f89;
assign v375595c = hbusreq7_p & v3a6fbd3 | !hbusreq7_p & v37287fb;
assign v3a6eeca = hgrant3_p & v3a6505b | !hgrant3_p & v3758c62;
assign v3a7087d = hmaster0_p & v3a63805 | !hmaster0_p & v3a59905;
assign v37431d8 = hmaster0_p & v8455ab | !hmaster0_p & v376ae07;
assign v3a6d364 = hbusreq2_p & v3a6fc63 | !hbusreq2_p & v8455ab;
assign v3a55b91 = hmaster2_p & v37282cf | !hmaster2_p & !v37521ed;
assign v373d8ec = hlock4 & v3770d22 | !hlock4 & v3a5dc35;
assign v373d5df = hmaster0_p & v376df25 | !hmaster0_p & v3774a9c;
assign v3735f25 = hbusreq4 & v3a6143b | !hbusreq4 & !v8455b5;
assign v3a5e394 = jx3_p & v3774618 | !jx3_p & v3a6dada;
assign v3a6ed27 = hbusreq5 & v373240c | !hbusreq5 & v3a71149;
assign v3a66037 = hbusreq4_p & v37373af | !hbusreq4_p & v372c197;
assign v3a6a089 = hmaster2_p & v20d166d | !hmaster2_p & v372a20c;
assign v3a706cb = hmaster2_p & v3a66ada | !hmaster2_p & v372edd9;
assign v3a70175 = hbusreq7_p & v3a5e7e0 | !hbusreq7_p & v3761026;
assign v37655ff = hbusreq5 & v373b732 | !hbusreq5 & v3a61dd0;
assign v3724026 = hbusreq0_p & v3a562a9 | !hbusreq0_p & v8455ab;
assign v3a5f449 = hmaster0_p & v3a56243 | !hmaster0_p & !v37455cd;
assign v377eb2d = hready & v8455ab | !hready & v376c211;
assign v3776670 = hbusreq1_p & v3a5c5ae | !hbusreq1_p & !v39a537f;
assign v375ac16 = hbusreq5 & v3759007 | !hbusreq5 & v3a706f6;
assign v3a55542 = hbusreq5_p & v3a65552 | !hbusreq5_p & v3a71435;
assign v372967b = hgrant5_p & v37650e4 | !hgrant5_p & v3a5e985;
assign v376b03a = jx0_p & v8455c5 | !jx0_p & v8455ab;
assign v3a58b28 = hgrant2_p & v3a6f46a | !hgrant2_p & v373e1a6;
assign v3733e88 = hbusreq3_p & v376ff61 | !hbusreq3_p & v372b5b0;
assign v373b9ab = hmaster0_p & v3a6f6e2 | !hmaster0_p & v372e5fb;
assign v37272ca = hlock5 & v3728793 | !hlock5 & v3a5b310;
assign v3a6c7fe = hbusreq6_p & v373c23e | !hbusreq6_p & v3742140;
assign v372d1d7 = hbusreq4_p & v3759886 | !hbusreq4_p & !v8455ab;
assign v3764334 = hlock5_p & v37314f0 | !hlock5_p & v3a69674;
assign v1e3824a = hbusreq0 & v964c47 | !hbusreq0 & v8455ab;
assign v373b95e = hmaster1_p & v377d077 | !hmaster1_p & v3a6f937;
assign v3a54393 = hgrant6_p & v377938d | !hgrant6_p & v376d240;
assign v8455ab = 1;
assign v3773b2f = hgrant3_p & v8455ab | !hgrant3_p & v37462ca;
assign v3727c3c = hmaster0_p & v3a661fe | !hmaster0_p & v375d832;
assign v377074b = hlock8_p & v3808884 | !hlock8_p & !v372704f;
assign v3731bb5 = hmaster2_p & v375b0d5 | !hmaster2_p & v3a67403;
assign v3a6abcc = hlock0 & v3757009 | !hlock0 & v374586b;
assign v3a6d642 = hlock2_p & v375eb97 | !hlock2_p & v8455e7;
assign v375eeb9 = hmaster0_p & v8455ab | !hmaster0_p & v3a694ec;
assign v37503c9 = hbusreq0 & v37612dd | !hbusreq0 & v377722d;
assign v3748146 = hbusreq4 & v3760f64 | !hbusreq4 & v8455bb;
assign v3a6b1e4 = hbusreq2_p & v377395b | !hbusreq2_p & v8455ab;
assign v1e37cd6 = hbusreq6_p & v8455ab | !hbusreq6_p & v3a5eadd;
assign v3774655 = hbusreq8 & v3732511 | !hbusreq8 & v3a5857c;
assign v3728793 = hbusreq5 & v3a5b310 | !hbusreq5 & v374decf;
assign v3a5755b = hmaster2_p & v2ff8cfd | !hmaster2_p & v37325f4;
assign v375d94c = hmaster0_p & v3744e13 | !hmaster0_p & v3774d9a;
assign v37504f2 = jx0_p & v375038a | !jx0_p & v3a6fe7c;
assign v375c4e6 = hbusreq4 & v3730755 | !hbusreq4 & v8455ab;
assign v374e873 = hbusreq7 & v375194a | !hbusreq7 & v3723025;
assign v3a6c5ed = hbusreq8_p & v373562f | !hbusreq8_p & v3a70fcc;
assign v375156a = hgrant2_p & v8455ba | !hgrant2_p & v3a6f1b2;
assign v3747824 = hmaster2_p & v3752a7a | !hmaster2_p & v374e124;
assign v372349f = hmaster1_p & v373e5c8 | !hmaster1_p & v374d9b7;
assign v377a039 = hbusreq2_p & v3752511 | !hbusreq2_p & v3a6e8fa;
assign v3a6fe0e = hlock4_p & v377169f | !hlock4_p & v3a65da7;
assign v3757dd1 = hbusreq5_p & v3a696a7 | !hbusreq5_p & v377e784;
assign v377b860 = hgrant2_p & v376bb26 | !hgrant2_p & v374abc9;
assign v375da9c = hlock2 & v3a6f4d2 | !hlock2 & v3809b31;
assign v3777da2 = hlock0 & v3a5f9e6 | !hlock0 & v3a7168b;
assign v3a69fbe = hbusreq2_p & v374978c | !hbusreq2_p & !v8455ab;
assign v3a2a911 = hlock5 & v372668c | !hlock5 & v325c90f;
assign v37583ea = hgrant5_p & v3773530 | !hgrant5_p & v374b225;
assign v3a69f36 = hgrant3_p & v8455b5 | !hgrant3_p & v377514f;
assign v377050c = hbusreq5_p & v3733711 | !hbusreq5_p & v373373d;
assign v3737d90 = hmaster2_p & v377308e | !hmaster2_p & v372346b;
assign v3a701af = hbusreq8 & v374891f | !hbusreq8 & !v37316f3;
assign v376b44a = hbusreq8 & v3a5511c | !hbusreq8 & v3a712b5;
assign v377d671 = hmaster1_p & v376f017 | !hmaster1_p & v37542d8;
assign v374a0f0 = hbusreq8 & v373e0b5 | !hbusreq8 & v3749f3b;
assign v376c87d = hgrant6_p & v8455ab | !hgrant6_p & v1e37721;
assign v3a711f8 = hbusreq7_p & v3751210 | !hbusreq7_p & !v3740328;
assign v3a7128b = hmaster2_p & v3770e95 | !hmaster2_p & v3771d4f;
assign v3a6f887 = hlock5 & v3778bef | !hlock5 & v8639e9;
assign v372ab42 = jx1_p & v3a6b864 | !jx1_p & v3728581;
assign v3731304 = hgrant3_p & v3a635ea | !hgrant3_p & v3769510;
assign v3a61375 = hmaster1_p & v3808cf7 | !hmaster1_p & v372fbb1;
assign v3a6617b = hbusreq0 & v8827d7 | !hbusreq0 & v373a18b;
assign v3a704af = hmaster0_p & v3a6dfb2 | !hmaster0_p & !v3736d5e;
assign v3806465 = hbusreq7 & v377cb3d | !hbusreq7 & v3746f9d;
assign v3765f61 = jx0_p & v374474d | !jx0_p & v3745928;
assign v377278b = hmaster2_p & v3a6f963 | !hmaster2_p & !v8455ab;
assign v3a7093d = hmaster0_p & v377234d | !hmaster0_p & v372ee4b;
assign v3a6b462 = hlock5_p & v373a8c0 | !hlock5_p & v372c8d0;
assign v3a6143b = hbusreq1_p & v3a71424 | !hbusreq1_p & v8455ab;
assign v3749a1d = hgrant2_p & v8455ab | !hgrant2_p & !v372ead5;
assign v375818b = hmaster0_p & v8455e7 | !hmaster0_p & v3a6a2f8;
assign v3a715a2 = hbusreq8_p & v3a6c0b7 | !hbusreq8_p & v3778211;
assign v373d4c6 = hbusreq2 & v372e27f | !hbusreq2 & v374dfea;
assign v3739d4a = stateG10_1_p & v3723430 | !stateG10_1_p & v3764834;
assign v1e37c79 = hmaster3_p & v3a710d8 | !hmaster3_p & !v3734a96;
assign v3764141 = hbusreq6_p & v3a635ea | !hbusreq6_p & cb1cc0;
assign v3a6d48a = hmaster2_p & v3769740 | !hmaster2_p & v3a61cd7;
assign v377c28e = hgrant4_p & v376a6f1 | !hgrant4_p & v375887e;
assign v3a6fabe = hbusreq6_p & v37790ef | !hbusreq6_p & v374c4e9;
assign v375fbc6 = hbusreq4_p & v37639b1 | !hbusreq4_p & v8455b0;
assign v374f501 = hgrant4_p & v8455ab | !hgrant4_p & v3a65aca;
assign v3a66f40 = hmaster1_p & v3a70478 | !hmaster1_p & !v3779ac0;
assign v3a714ff = hbusreq2_p & v3726609 | !hbusreq2_p & !v3a68591;
assign v3762802 = hbusreq7_p & v3767a08 | !hbusreq7_p & v373af15;
assign v3a69b77 = hmaster0_p & v3a6e37c | !hmaster0_p & !v377ba8a;
assign v3a6f0f3 = hlock7 & v372a2ff | !hlock7 & v3a700ef;
assign v3a6f21c = hgrant4_p & v3a6ac66 | !hgrant4_p & v8455ab;
assign v3724667 = hlock0 & v38072fd | !hlock0 & v377cdbe;
assign v377cf7f = hbusreq4 & v39a4f09 | !hbusreq4 & v375b233;
assign v3a6e57f = hgrant4_p & v8455ab | !hgrant4_p & !v372ed88;
assign v3774200 = hmaster0_p & v3a576c0 | !hmaster0_p & v8455ab;
assign v3723dae = hgrant6_p & v3a6f2d4 | !hgrant6_p & v3a5fb37;
assign v3734d8a = hbusreq0 & v3a58d67 | !hbusreq0 & v3a64af7;
assign v374da61 = hbusreq4_p & c39398 | !hbusreq4_p & !v8455ab;
assign v37431b5 = hbusreq3 & v3a63abb | !hbusreq3 & v8455ab;
assign v3a55b1d = hbusreq0 & v376fb6b | !hbusreq0 & v375f8dd;
assign v3741f69 = hgrant6_p & v3754fd2 | !hgrant6_p & v37709bb;
assign v37560b4 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3736968;
assign v3765dbc = hmaster2_p & v376bca9 | !hmaster2_p & v37763d1;
assign v3a6953d = hmaster2_p & ae317f | !hmaster2_p & v8455ca;
assign v3a70b4a = hmaster2_p & v3771c85 | !hmaster2_p & v372f853;
assign v3734aae = hbusreq4 & v8455ab | !hbusreq4 & v8455b0;
assign v3a56aee = hmaster3_p & v373d8e4 | !hmaster3_p & !v376b1ee;
assign v372f7ca = hmaster0_p & v377040f | !hmaster0_p & v375881d;
assign v374c720 = hbusreq5_p & v3779cf6 | !hbusreq5_p & v37c36bf;
assign v372948c = hbusreq2_p & v2ff9190 | !hbusreq2_p & v37390c4;
assign v3a6f2c0 = hbusreq6 & v3a644cd | !hbusreq6 & v8455ab;
assign v373f95b = hgrant4_p & v37444b4 | !hgrant4_p & v373ebf9;
assign v372b4ba = stateG10_1_p & v3a6f646 | !stateG10_1_p & v37353c0;
assign v3744b87 = hbusreq5_p & v374c007 | !hbusreq5_p & v372ea5d;
assign v3767d2c = hmaster3_p & v373ca17 | !hmaster3_p & v3a70f05;
assign v373cdb7 = hlock3_p & v3a68426 | !hlock3_p & v8455b7;
assign v3744999 = hbusreq4 & v373fe74 | !hbusreq4 & v23fdaed;
assign v372b3b6 = jx1_p & v3a70fb1 | !jx1_p & v374b364;
assign v3774385 = hmaster0_p & v3a635ea | !hmaster0_p & v37461d9;
assign v375f6ef = hgrant6_p & v3727713 | !hgrant6_p & v3763af8;
assign v37476c5 = hmaster1_p & v3726c61 | !hmaster1_p & v377f6c3;
assign v3a70116 = hmaster2_p & v3755002 | !hmaster2_p & v3a5fdfc;
assign v3737b1a = hmaster1_p & v2678bee | !hmaster1_p & v375ea13;
assign v374549a = hmaster2_p & v3a627a4 | !hmaster2_p & v373015f;
assign v377d2ee = hlock0 & v377b7f9 | !hlock0 & v37513bc;
assign v3a6cedc = hbusreq3_p & v3737c13 | !hbusreq3_p & v8455ab;
assign v3a6fb0c = hgrant4_p & v3a70b5e | !hgrant4_p & v8455ab;
assign v3a652de = hbusreq4_p & v3724c25 | !hbusreq4_p & v377bca1;
assign v3a6ffe1 = hbusreq2_p & v8c34b7 | !hbusreq2_p & !v8455ab;
assign v37235fa = hmaster1_p & v376edbb | !hmaster1_p & v8455ab;
assign v3a5715d = hbusreq4 & v37285ad | !hbusreq4 & v3a5408c;
assign v37384a9 = hmaster0_p & v376f56d | !hmaster0_p & v3a5ed31;
assign v375a0ed = hmaster3_p & v3a712a6 | !hmaster3_p & v372775f;
assign v3753fe6 = hbusreq8_p & v373bd5e | !hbusreq8_p & v37389b1;
assign v375579f = hmaster3_p & v3a6f701 | !hmaster3_p & a5d7b0;
assign v3743e90 = hgrant5_p & v8455ab | !hgrant5_p & v376abd9;
assign v3a710f4 = hmaster2_p & v37294d3 | !hmaster2_p & v3739ab6;
assign v37291e4 = hmaster3_p & v37377f0 | !hmaster3_p & v377457e;
assign v375a754 = hbusreq5_p & v376626a | !hbusreq5_p & v373930f;
assign v3a53e50 = hbusreq0 & v37254d2 | !hbusreq0 & v3762f1a;
assign v3762d3e = hbusreq6_p & v37265f6 | !hbusreq6_p & v37471e0;
assign v3a6b575 = hgrant4_p & v37521f6 | !hgrant4_p & v3a611e6;
assign v3a5ff09 = hbusreq6 & v3a6f612 | !hbusreq6 & v8455ab;
assign v3a70b62 = hbusreq7 & v3a685ee | !hbusreq7 & v3760617;
assign v372e661 = hlock0 & v373eaee | !hlock0 & v373ac12;
assign v3a709a0 = stateG10_1_p & v35772a5 | !stateG10_1_p & !b6b4ea;
assign v3771739 = hmaster0_p & v37398e5 | !hmaster0_p & !v3a62dfa;
assign v3743fe3 = hlock0 & v3a685c7 | !hlock0 & v3764270;
assign v3a6ef26 = hmaster2_p & v3807aa1 | !hmaster2_p & !v375c9f0;
assign stateG10_5 = !v39ed7ea;
assign v3760279 = hgrant3_p & v8455ab | !hgrant3_p & v376897b;
assign v3773e77 = hbusreq4 & v3752933 | !hbusreq4 & v3a641d5;
assign v375d06d = hmaster2_p & v2aca977 | !hmaster2_p & !v3a6ab5f;
assign v3a5f154 = hlock4 & v3a605af | !hlock4 & v374c3d0;
assign v3a6f54b = hbusreq5_p & v39ebb2e | !hbusreq5_p & v37266df;
assign v39a4dd4 = hlock0_p & v375803a | !hlock0_p & v372bcbc;
assign v3739ab2 = hbusreq5 & v3732bb6 | !hbusreq5 & !v377f61c;
assign v3a713e7 = hmaster2_p & v37468e5 | !hmaster2_p & v377e825;
assign v373803a = hbusreq8_p & v3779d06 | !hbusreq8_p & b0ac65;
assign b0e59c = hmaster2_p & v37668e9 | !hmaster2_p & v372edf6;
assign v3a6fccc = hmaster0_p & v3a6fe0d | !hmaster0_p & v373b599;
assign v3a6eb1d = hbusreq4 & v3a667e7 | !hbusreq4 & !v8455ca;
assign v3a7090f = hmaster2_p & v3745828 | !hmaster2_p & v3724fdb;
assign v3a67588 = hbusreq0 & v3770e2d | !hbusreq0 & v3a70f5d;
assign v376749b = hmaster1_p & v372cdde | !hmaster1_p & v3a5a05d;
assign v372e0b7 = jx1_p & v373f13e | !jx1_p & v3a66039;
assign v377ccb7 = hlock8 & v38069c0 | !hlock8 & v376af8e;
assign v3757301 = hmaster0_p & v8455b9 | !hmaster0_p & v373ea7f;
assign v374c4bc = hgrant3_p & v372d02d | !hgrant3_p & v3753fe0;
assign v377326a = hmaster0_p & v376efaa | !hmaster0_p & b8f82c;
assign v376e507 = hlock7 & v3a712f5 | !hlock7 & v3779593;
assign v3744458 = hgrant2_p & v37467f7 | !hgrant2_p & v372fb9d;
assign v376b38c = hmaster0_p & v3758ce2 | !hmaster0_p & v3a669e9;
assign v3a669be = hmaster1_p & v37365f8 | !hmaster1_p & v3a6574d;
assign v3a7061f = hmaster3_p & v3a70013 | !hmaster3_p & v377c47c;
assign v37367da = hlock3_p & v375a18e | !hlock3_p & !v8455ab;
assign v3a6ceb7 = hbusreq2_p & v1e37b65 | !hbusreq2_p & v373ef30;
assign v372f0c7 = hmaster0_p & v8455b0 | !hmaster0_p & v37684c3;
assign v372d435 = hgrant4_p & v37319cd | !hgrant4_p & v3a64722;
assign v3a6eb45 = hgrant1_p & v374f307 | !hgrant1_p & !v8455ab;
assign v3772310 = hbusreq4_p & v3726d1f | !hbusreq4_p & v373f3b5;
assign v3726b10 = hbusreq0 & v3a64374 | !hbusreq0 & v3a71295;
assign v3729c9a = hbusreq7_p & v3734279 | !hbusreq7_p & v3a5f609;
assign v372b813 = hbusreq5_p & v3a70cd6 | !hbusreq5_p & v35b987f;
assign v3a53a43 = hmaster3_p & v376f250 | !hmaster3_p & v3762324;
assign v3768429 = hmaster0_p & v3760750 | !hmaster0_p & v3776f07;
assign v377c271 = hgrant7_p & v3744f1e | !hgrant7_p & v3743d47;
assign v3730cc8 = hgrant0_p & v8455ab | !hgrant0_p & v3a56417;
assign v3771633 = hmaster1_p & v3a635ea | !hmaster1_p & v372f4e6;
assign v3756057 = hlock6 & v3a6fffc | !hlock6 & ae0781;
assign v3778b8c = hbusreq3_p & v37533e3 | !hbusreq3_p & v35772a6;
assign v3a6992f = hmaster2_p & v3a637dd | !hmaster2_p & !v374109e;
assign v3a706a6 = hbusreq4_p & v39a5420 | !hbusreq4_p & v3727486;
assign v3724665 = hmaster1_p & v3a29814 | !hmaster1_p & v3750cfa;
assign v3a624ec = hlock5_p & v3773eee | !hlock5_p & !v374e21d;
assign v377bd63 = hmaster0_p & v377234d | !hmaster0_p & v3a6facb;
assign v3a60cf8 = hmaster1_p & v8455ab | !hmaster1_p & v373beae;
assign v3740681 = hmaster0_p & v3808d56 | !hmaster0_p & v372efee;
assign v3753f77 = hbusreq5 & v374314f | !hbusreq5 & v3a58c07;
assign v3747552 = hgrant2_p & v8455ab | !hgrant2_p & v3a6eac1;
assign v37454cc = hlock0 & v3730695 | !hlock0 & v3759edb;
assign v3a67d83 = hmaster0_p & v3772696 | !hmaster0_p & !v3807765;
assign v3778a89 = hbusreq2 & v1e38224 | !hbusreq2 & v8455ab;
assign v3733384 = hmaster0_p & v3a7058d | !hmaster0_p & v8455ab;
assign v376fdfb = hbusreq7_p & v372e5a8 | !hbusreq7_p & v3a6ef61;
assign v380937f = hbusreq8 & v3739b6a | !hbusreq8 & v3a60276;
assign v372e550 = hmaster1_p & v35b774b | !hmaster1_p & v373f691;
assign v377db89 = hlock5_p & v8455ab | !hlock5_p & v375f888;
assign v3761ad0 = hbusreq3_p & v37674c1 | !hbusreq3_p & v3a5c1a5;
assign v377a4bd = hmaster1_p & v375a268 | !hmaster1_p & v3a6f48a;
assign v3734bf8 = hbusreq4 & v376b21a | !hbusreq4 & !v8455ab;
assign v3779595 = hbusreq5_p & v376f56d | !hbusreq5_p & v3739ab4;
assign v372a00b = hbusreq2_p & v377b774 | !hbusreq2_p & v3724e8e;
assign v373104a = hbusreq0 & v37637ef | !hbusreq0 & v8455ab;
assign v373b92c = hbusreq4 & v3378e07 | !hbusreq4 & v37285eb;
assign v374069b = hmaster1_p & v377bac2 | !hmaster1_p & v3769d79;
assign v3730181 = hlock3_p & v8455ab | !hlock3_p & !v3726ef1;
assign v3730252 = hmaster1_p & v3760276 | !hmaster1_p & v37558f2;
assign v3a7113b = hbusreq5 & v3a6f335 | !hbusreq5 & v8455ab;
assign v3a70e72 = hbusreq5_p & v374478f | !hbusreq5_p & v3a5f648;
assign v3779b5b = hgrant5_p & v3727a6d | !hgrant5_p & v3a656c7;
assign v37586cd = hmaster1_p & v3a71215 | !hmaster1_p & !v377d080;
assign v3758b8b = hlock5 & v3a70af0 | !hlock5 & v3a70a75;
assign v374ba65 = hbusreq2 & v373d78b | !hbusreq2 & v8455ab;
assign v3a5eadd = hbusreq2_p & v8455ab | !hbusreq2_p & v3a6c2b6;
assign v3a297f5 = hmaster1_p & v372ba66 | !hmaster1_p & v372b12d;
assign v9c8578 = hbusreq7_p & v3a70cb3 | !hbusreq7_p & v375d966;
assign v3a665b3 = hmaster2_p & v3a582c5 | !hmaster2_p & v37793a4;
assign v3a6e9b0 = hlock5 & v3772021 | !hlock5 & v374d13d;
assign v3767471 = hbusreq5_p & v3a59c21 | !hbusreq5_p & !v8455ab;
assign v3a60882 = hgrant2_p & v377d4a0 | !hgrant2_p & v3a58a16;
assign v375e120 = hbusreq5 & v373796a | !hbusreq5 & v3a7157d;
assign v3779003 = hbusreq5_p & v374de25 | !hbusreq5_p & !v3724325;
assign d8c443 = hmaster2_p & v373fa89 | !hmaster2_p & v3a705a6;
assign v3735c9d = hgrant6_p & v376bb26 | !hgrant6_p & v377b860;
assign v375d182 = hlock1_p & v3a61237 | !hlock1_p & v3a6ebe7;
assign v3777417 = hgrant3_p & v3739018 | !hgrant3_p & !v37794fa;
assign v374cda5 = hlock1_p & v3a622c0 | !hlock1_p & !v8455b6;
assign v39a4e8f = hgrant3_p & v8455ab | !hgrant3_p & v3a6cedc;
assign v3731d76 = hmaster2_p & v8455ab | !hmaster2_p & v3738dac;
assign v3a6eaf4 = hbusreq2_p & v3a70ee7 | !hbusreq2_p & v3733d6e;
assign v3728ea7 = hgrant6_p & v3a70e75 | !hgrant6_p & v376804b;
assign v375bf12 = hmaster1_p & v3766185 | !hmaster1_p & !v3779a66;
assign v3a5ce55 = hbusreq5_p & v3762806 | !hbusreq5_p & !v8455ab;
assign v372ccea = stateG3_2_p & v8455ab | !stateG3_2_p & v845601;
assign v37702e8 = hbusreq8_p & v3775729 | !hbusreq8_p & v3a58c95;
assign v3739e0e = hbusreq7 & v3734e0b | !hbusreq7 & v3a6f2fd;
assign v37762cd = hmaster2_p & v3a6935c | !hmaster2_p & v37747f8;
assign v3a65e6a = hmaster0_p & v37570f8 | !hmaster0_p & v3725e0d;
assign v3a57584 = hbusreq1_p & v3a6f5df | !hbusreq1_p & v8455ab;
assign v3739dae = hgrant6_p & v3777996 | !hgrant6_p & v37737c9;
assign v37325ed = hbusreq5 & afadd1 | !hbusreq5 & v3a5e030;
assign v376f0a0 = hgrant6_p & v8455ab | !hgrant6_p & v3a6190f;
assign v3a6fbec = hbusreq5 & v3754a8e | !hbusreq5 & v8455ab;
assign v377934a = hlock3_p & v3a6fa6e | !hlock3_p & v8455b7;
assign v3a6f588 = hbusreq3 & v3a6ad8b | !hbusreq3 & v38072fd;
assign v3744501 = hbusreq6_p & v8455e1 | !hbusreq6_p & v375dbd4;
assign v3a70bb3 = hbusreq0_p & v372dadb | !hbusreq0_p & v375fbd7;
assign v377a110 = hbusreq0_p & v3760d83 | !hbusreq0_p & v8455ab;
assign v374e353 = hbusreq4 & v3a6f0e9 | !hbusreq4 & v3730695;
assign v3a6ef64 = hbusreq7_p & v375c99d | !hbusreq7_p & v377acde;
assign v372e4a7 = hmaster0_p & v3a6f541 | !hmaster0_p & v3739b7a;
assign v3a57046 = hgrant4_p & v8455c2 | !hgrant4_p & v373d737;
assign v3732e1b = hbusreq1_p & v3809adf | !hbusreq1_p & !v3a70c07;
assign v3778173 = hgrant2_p & v372abd8 | !hgrant2_p & v3761678;
assign v376d36a = hlock7 & v3a71512 | !hlock7 & v3a6f5aa;
assign v375524f = hbusreq4 & v374db79 | !hbusreq4 & !v3a70dae;
assign v3773bb0 = hgrant6_p & v373ee17 | !hgrant6_p & v3a6f4d0;
assign v380732c = hmaster1_p & v3743287 | !hmaster1_p & v3378f5d;
assign v3750025 = hgrant0_p & v8455ab | !hgrant0_p & v3a6fae2;
assign v3a6d6fe = hlock0_p & v3758cec | !hlock0_p & !v8455ab;
assign v3a702f2 = hmaster0_p & v3a711df | !hmaster0_p & v1e37cf9;
assign v3a6fdf8 = hgrant3_p & v8455e7 | !hgrant3_p & !v3a5f0a7;
assign v3728992 = hmaster1_p & v377b6ce | !hmaster1_p & v3733cfb;
assign v3a70ee9 = hbusreq0 & v3a67cfe | !hbusreq0 & !v8455ab;
assign v377673f = hmaster1_p & v37534c6 | !hmaster1_p & v28896cd;
assign v376648e = hbusreq6 & v372c3df | !hbusreq6 & v38097f6;
assign v376d7c6 = hlock4 & v3a6fbc5 | !hlock4 & v375d10e;
assign v3737ada = hlock3_p & v3772cf2 | !hlock3_p & v3a6ebfd;
assign v37611b7 = hbusreq0_p & v3a635ea | !hbusreq0_p & v3a63621;
assign v3a6fc48 = hlock4_p & v372b231 | !hlock4_p & v8455cb;
assign v374cc7f = hgrant3_p & v372493b | !hgrant3_p & v377d7dd;
assign v3806c9a = hgrant4_p & v3a53eeb | !hgrant4_p & v3750d09;
assign v3a7112d = jx3_p & v3a71156 | !jx3_p & v1e382dc;
assign v3807341 = hlock6 & v38074bc | !hlock6 & v376bfc3;
assign v3a6abfe = hmaster1_p & v3767e7f | !hmaster1_p & v374bd4a;
assign v3a700be = hmaster1_p & v3a635ea | !hmaster1_p & v372610c;
assign v3a712f0 = hbusreq3_p & v3806818 | !hbusreq3_p & !v3a5df97;
assign v3a6cc2a = hmaster1_p & v3a6b931 | !hmaster1_p & v3742a61;
assign v3a70fbf = hmaster2_p & v8455ab | !hmaster2_p & v374f82e;
assign v3a6fd12 = hmaster0_p & v3760452 | !hmaster0_p & v373058e;
assign v375df5a = hbusreq5 & v3808db6 | !hbusreq5 & v3a5514a;
assign v3a69ad9 = hbusreq5_p & v3741197 | !hbusreq5_p & v3735afe;
assign v376b908 = hgrant4_p & v3a5aaed | !hgrant4_p & v3a70674;
assign v3a70454 = hmaster1_p & v3a635ea | !hmaster1_p & v3a6279c;
assign v37297af = hbusreq0 & v3774791 | !hbusreq0 & v3755f9a;
assign v372372d = hbusreq0 & v37706bf | !hbusreq0 & v3745e1f;
assign v374571a = hmaster2_p & adf78a | !hmaster2_p & v372b5f5;
assign v3732df3 = jx0_p & v3724a15 | !jx0_p & v37332ca;
assign v372bffa = hgrant6_p & v3735906 | !hgrant6_p & v3732202;
assign v376f814 = hbusreq5 & v376fe90 | !hbusreq5 & v3a70ae8;
assign v3a6b266 = hbusreq5_p & v3a633c5 | !hbusreq5_p & v1e3737d;
assign v373168f = hmaster1_p & v3760a0b | !hmaster1_p & v8f1dd1;
assign b8f82c = hmaster2_p & v8455ab | !hmaster2_p & v377234d;
assign v375495e = hmaster0_p & v373580d | !hmaster0_p & v3742cd4;
assign v3a62bd5 = hbusreq5 & v377d107 | !hbusreq5 & v3a6ff4e;
assign v3759e3c = hbusreq6_p & v3a6fdb4 | !hbusreq6_p & v372ade8;
assign v3745536 = stateA1_p & v8455ab | !stateA1_p & v8455ff;
assign v3a658bf = locked_p & v3806a74 | !locked_p & v35772a6;
assign v376930a = hbusreq8_p & v375a1fd | !hbusreq8_p & v376ce1a;
assign d2e9f6 = hlock6 & v3757ec4 | !hlock6 & v3a6c63e;
assign v37379a2 = hmaster1_p & v376111d | !hmaster1_p & v372e754;
assign v3754727 = hmaster2_p & v3a5665e | !hmaster2_p & v372912f;
assign v3a71028 = hbusreq4_p & v3a6f505 | !hbusreq4_p & v3a613cc;
assign v377b311 = hmaster2_p & v8455ab | !hmaster2_p & !v8455e7;
assign v3a6c933 = hmaster2_p & v8455e1 | !hmaster2_p & !v1e37370;
assign v8455ce = hbusreq7 & v8455ab | !hbusreq7 & !v8455ab;
assign v3734a99 = busreq_p & v3a635ea | !busreq_p & v37353d9;
assign v3735930 = hmaster0_p & v376d9ad | !hmaster0_p & v3a6f427;
assign v375b24f = hbusreq7 & v374c3bf | !hbusreq7 & v3a71448;
assign v374f528 = hgrant4_p & v8455ab | !hgrant4_p & v3742ec5;
assign v3a7036b = hgrant5_p & v8455ab | !hgrant5_p & v3724a6d;
assign v3a58d68 = hmaster2_p & v373badc | !hmaster2_p & v3763191;
assign v3a6e804 = hlock6 & v37326a5 | !hlock6 & v375d05d;
assign v3759dfb = hmaster2_p & v3a637dc | !hmaster2_p & v3a653e4;
assign v372777c = hgrant3_p & v8455ab | !hgrant3_p & v3806bc8;
assign v3a707b7 = hbusreq6_p & v377b774 | !hbusreq6_p & v3724e8e;
assign v3769cc2 = hlock0_p & v35b9d52 | !hlock0_p & v2aca977;
assign v3762807 = hbusreq4_p & v3a70ee7 | !hbusreq4_p & v3733d6e;
assign v374890e = hgrant4_p & v8455ab | !hgrant4_p & v3734913;
assign v3a71012 = hgrant6_p & v3733e9e | !hgrant6_p & v372ef40;
assign v3a70519 = hbusreq5_p & v3a6eed9 | !hbusreq5_p & v3a707a7;
assign v3751faf = hgrant3_p & v3a6f627 | !hgrant3_p & v375a02d;
assign v372ea02 = hmaster0_p & v3763bb8 | !hmaster0_p & v1e37c38;
assign v3772470 = hmaster1_p & v8455ab | !hmaster1_p & v374a8da;
assign v376d1cb = hmaster2_p & v3a62c12 | !hmaster2_p & v2619b04;
assign v373e760 = hbusreq3_p & v3747302 | !hbusreq3_p & v3762389;
assign v375cfa5 = hlock6 & v373087b | !hlock6 & v373c2ec;
assign v3771971 = hmaster0_p & v37291c0 | !hmaster0_p & v3743c40;
assign v3732e45 = hmaster2_p & v3a60b2e | !hmaster2_p & v372d8f9;
assign v3765a69 = hmaster0_p & v3a6f3ec | !hmaster0_p & v8455ab;
assign v3a700d2 = hmaster3_p & v8455ab | !hmaster3_p & v3a7050d;
assign v3762929 = hgrant4_p & v37350b7 | !hgrant4_p & v3a6783b;
assign v3737f8b = hbusreq5_p & v377de57 | !hbusreq5_p & a15d51;
assign v3a6a42a = jx0_p & b85e8b | !jx0_p & v3a5ca22;
assign v3a62322 = hmaster2_p & v37c0382 | !hmaster2_p & !v8455ab;
assign v376942f = hlock2 & v2092b23 | !hlock2 & v372f3f7;
assign v3a7017b = hmaster1_p & v3733d3f | !hmaster1_p & v3761719;
assign v37536b8 = hmaster1_p & v3a6fd10 | !hmaster1_p & v37298be;
assign v8f2b25 = hmaster3_p & v372c6b3 | !hmaster3_p & v8455ab;
assign v377098c = hmaster0_p & v377989c | !hmaster0_p & v3723023;
assign v377b8b9 = hbusreq3 & v3776ce0 | !hbusreq3 & v377c6b3;
assign v376eaca = hlock2 & v3a590fb | !hlock2 & v29256bb;
assign v3a5770f = hbusreq8 & v3a6fb9e | !hbusreq8 & v373be73;
assign v3732359 = hbusreq0 & v372904d | !hbusreq0 & v8455ab;
assign v373db68 = hbusreq5_p & v3a6f2e5 | !hbusreq5_p & v376140e;
assign v37279df = jx1_p & v3a71545 | !jx1_p & bdbe8b;
assign v372edf8 = hgrant4_p & v37782c9 | !hgrant4_p & v93144b;
assign v3a674c4 = hbusreq7 & v3a707ef | !hbusreq7 & v3a67312;
assign v374b19b = hmaster1_p & v3a635ea | !hmaster1_p & v3a714f1;
assign v3a69e8c = hgrant2_p & v8455ab | !hgrant2_p & v3754260;
assign v3754bd4 = hmaster2_p & v1e382e7 | !hmaster2_p & v39a537f;
assign v3a5c7be = hmaster2_p & v3a6f42e | !hmaster2_p & v373c21c;
assign v37356ec = hmaster0_p & v37356f0 | !hmaster0_p & v3722dfb;
assign v9684f8 = hbusreq4 & v373fe5e | !hbusreq4 & v8455e7;
assign v373198c = hmaster0_p & v37242cb | !hmaster0_p & v3757966;
assign v377c307 = hbusreq5 & v376b290 | !hbusreq5 & v3a2a107;
assign v35b7070 = hlock8_p & v33789d2 | !hlock8_p & v3a5b4a0;
assign v373d593 = hmaster2_p & v3a5a510 | !hmaster2_p & v3733e9e;
assign v3725819 = hbusreq4 & v3a696ed | !hbusreq4 & v8455ab;
assign v3744cfe = hbusreq6_p & v377f2ea | !hbusreq6_p & v3754237;
assign v3a6119e = hmaster2_p & v3735d9c | !hmaster2_p & v3778afd;
assign v3255a07 = hgrant3_p & v3a6432d | !hgrant3_p & v1e3741b;
assign v372a071 = hbusreq4_p & v3a667e7 | !hbusreq4_p & v375331e;
assign v37411c6 = hmaster2_p & v374be59 | !hmaster2_p & v373fb71;
assign v3a71458 = hbusreq6_p & v3733f37 | !hbusreq6_p & v380730d;
assign v3749846 = hmaster2_p & v3736610 | !hmaster2_p & v3a70957;
assign v3a6fc6b = hbusreq7 & v3775303 | !hbusreq7 & v8455ab;
assign v3746ac7 = hgrant0_p & v8455ab | !hgrant0_p & v38097fc;
assign v3772c7a = hlock4_p & v1e38241 | !hlock4_p & v373e827;
assign v3722dd6 = hbusreq7_p & v3809386 | !hbusreq7_p & !v8455ab;
assign v372a2ae = hmaster2_p & v3a5f41b | !hmaster2_p & !v8455ab;
assign v3743f9a = hlock8 & v3731579 | !hlock8 & v375f86d;
assign v373ccb9 = hgrant0_p & v3a6ffb6 | !hgrant0_p & v3a6f6de;
assign v3a6f6b8 = hgrant2_p & v8455ab | !hgrant2_p & v3a70ffb;
assign v37283c8 = hbusreq5 & v376293f | !hbusreq5 & v3a6ff4e;
assign v375a930 = hbusreq0 & v3a5d63f | !hbusreq0 & v3751238;
assign v3726098 = hgrant2_p & v37598dc | !hgrant2_p & v37566a2;
assign v3a709d6 = hbusreq7_p & v373db07 | !hbusreq7_p & !v3a6fb38;
assign v37344c6 = hgrant3_p & v3775aea | !hgrant3_p & v37555cd;
assign v3a71167 = hmaster1_p & v3773c5d | !hmaster1_p & v8455ab;
assign v3757811 = hbusreq0_p & v3a6b2ef | !hbusreq0_p & v376e611;
assign v376959b = jx0_p & v3a6f2bb | !jx0_p & v374b0e3;
assign v37462e3 = hbusreq6 & v3a55cd6 | !hbusreq6 & !v8455b5;
assign v3726006 = hgrant0_p & v3a70a88 | !hgrant0_p & v375d84b;
assign v3a6f317 = hbusreq7 & v3767415 | !hbusreq7 & v3a62236;
assign v37513fa = hgrant4_p & v3a70ac9 | !hgrant4_p & v37592a3;
assign v372e53f = hmaster1_p & v372b29d | !hmaster1_p & v372c762;
assign v374e418 = hgrant0_p & v3a6c860 | !hgrant0_p & v37772bf;
assign v3743e83 = hgrant6_p & v3766b5e | !hgrant6_p & v375b04f;
assign v3733ba7 = hmaster2_p & v377d74c | !hmaster2_p & v3a5b51a;
assign v376d657 = hbusreq8_p & v3746e30 | !hbusreq8_p & v3a67beb;
assign v3a5f439 = hmaster1_p & v3774e33 | !hmaster1_p & v3a706eb;
assign v39ebbae = hlock4_p & v2acb5a2 | !hlock4_p & v8455ab;
assign v372c3a4 = hbusreq6_p & v3a6cc72 | !hbusreq6_p & v8455ab;
assign v3744e11 = hgrant6_p & v377b6ce | !hgrant6_p & v375bd9c;
assign v3a6d175 = hgrant4_p & v377b6ce | !hgrant4_p & v3750b03;
assign v374a23a = hgrant2_p & v8455ab | !hgrant2_p & v3a6f581;
assign v374e8b5 = hmaster2_p & v3777da6 | !hmaster2_p & v3761719;
assign v3a6ffb2 = hbusreq7 & v376cb10 | !hbusreq7 & v3a707e3;
assign v3769c81 = hbusreq2 & v3a603bb | !hbusreq2 & v3a598a0;
assign v377d27f = hlock7_p & v3a70777 | !hlock7_p & v37506fe;
assign v377b5c4 = hgrant2_p & v3a6c580 | !hgrant2_p & v3738766;
assign v3a6ef73 = hbusreq5_p & v3a70000 | !hbusreq5_p & v2092a7a;
assign v3a714d5 = hmaster2_p & v3a62184 | !hmaster2_p & v37484e0;
assign v37416ea = hbusreq6 & v3a6f018 | !hbusreq6 & !v3740f3d;
assign v3a70e03 = hlock3_p & v377b8ee | !hlock3_p & !v8455ab;
assign v3773bf5 = hlock8 & v376ae9f | !hlock8 & v1e37916;
assign v3a6ecdf = hmaster1_p & v3a6fee7 | !hmaster1_p & v376f051;
assign v3779e21 = hbusreq8_p & v8455e7 | !hbusreq8_p & v3a6299c;
assign v3a70d92 = hbusreq7_p & v374445b | !hbusreq7_p & v3a6ef63;
assign v37721cd = hbusreq2_p & v377fb84 | !hbusreq2_p & v3758950;
assign v3749535 = hgrant5_p & v8455c6 | !hgrant5_p & b3b89e;
assign v3751905 = hgrant3_p & v8455ab | !hgrant3_p & !v1e3757b;
assign v3738c75 = hlock4 & v3a70e60 | !hlock4 & v375b9a0;
assign v37489ea = hgrant2_p & v3725230 | !hgrant2_p & v3a6e622;
assign v3729864 = hbusreq2_p & v374d04b | !hbusreq2_p & v3a6f9f6;
assign v3a6f729 = jx0_p & v3a60e6d | !jx0_p & v3728b47;
assign v37299e2 = hgrant3_p & v37c1a6f | !hgrant3_p & v373d34e;
assign v372343e = hbusreq4 & v3a6f520 | !hbusreq4 & !v8455ab;
assign v374254d = hmaster2_p & v3a5ef5c | !hmaster2_p & !v8455ab;
assign v3a6fb2a = hlock2_p & v372abd8 | !hlock2_p & v35772a6;
assign v374f4a0 = stateG10_1_p & v3a7048a | !stateG10_1_p & v3a568ac;
assign v8f1dd1 = hbusreq5_p & v3764e69 | !hbusreq5_p & v3a2976c;
assign v3762cd8 = hbusreq5 & v3a6f9a1 | !hbusreq5 & !v8455ab;
assign v3758e3c = hbusreq3_p & v3774c3f | !hbusreq3_p & v8455ab;
assign v374a50a = hmaster1_p & v374729b | !hmaster1_p & v375b342;
assign v377c97f = hbusreq7_p & v3a7066d | !hbusreq7_p & v3a6dac0;
assign v3764f2d = hbusreq8_p & v37431ac | !hbusreq8_p & v376df68;
assign v3733be1 = hgrant6_p & v3a5cb5f | !hgrant6_p & v3a6802b;
assign v3a67beb = hmaster1_p & v3a5d8a9 | !hmaster1_p & v8455ab;
assign v374afa3 = hmaster0_p & v3771ddb | !hmaster0_p & v3a59a05;
assign v3a685db = hmaster2_p & v375c791 | !hmaster2_p & v375f619;
assign v37575fd = hmaster1_p & v3809f73 | !hmaster1_p & v3a682f9;
assign v374fc20 = hmaster0_p & v375fcbf | !hmaster0_p & v377de50;
assign v3754ba1 = hbusreq5 & v375129f | !hbusreq5 & v37577cd;
assign v37252b7 = hmaster1_p & v374da8a | !hmaster1_p & v3a5efc4;
assign v3a710e3 = hmaster2_p & v37294d3 | !hmaster2_p & v376e854;
assign v37425a5 = hgrant4_p & v3776c04 | !hgrant4_p & v3a60a23;
assign v3a6fc99 = hbusreq5_p & v377ba7d | !hbusreq5_p & !v3a66110;
assign v3a6f360 = hmaster0_p & v376a2d6 | !hmaster0_p & v3a5c94c;
assign v3a647ce = hmaster1_p & v37bfc97 | !hmaster1_p & v8455ab;
assign v3a6f391 = jx0_p & v3741abc | !jx0_p & v3a705cf;
assign v3a5d673 = hbusreq1_p & v3a71456 | !hbusreq1_p & !v3a67d2e;
assign v3a6fd9f = hbusreq5_p & v375a16a | !hbusreq5_p & !v3a70ab1;
assign v372ac3a = hlock2_p & v3770559 | !hlock2_p & v35772a6;
assign v3764461 = hlock7 & v33789d0 | !hlock7 & v3723b33;
assign v3a71417 = hlock2_p & v8455ab | !hlock2_p & v3a5d923;
assign v3a6416b = hmaster2_p & v3a61397 | !hmaster2_p & v8455ab;
assign v3754328 = hmaster1_p & v8455ab | !hmaster1_p & v3775b7e;
assign v376e4a6 = hlock4_p & v3a5be93 | !hlock4_p & v3a702c2;
assign v3723549 = hbusreq6_p & v37709bb | !hbusreq6_p & v374fac6;
assign v3765cec = hmaster2_p & v375bfdf | !hmaster2_p & v377a356;
assign v374b310 = hbusreq2 & v3757d20 | !hbusreq2 & v376bb88;
assign v372dc35 = hbusreq8 & v3a64f1f | !hbusreq8 & v3a6e404;
assign v37302ea = hbusreq3_p & v3a707d1 | !hbusreq3_p & v8455ab;
assign v3728962 = hmaster2_p & v3763c09 | !hmaster2_p & v3a5d5a4;
assign v374ed4b = hgrant1_p & v8455b6 | !hgrant1_p & v8455ab;
assign v3762c8e = jx0_p & v3a59bf7 | !jx0_p & v375a56b;
assign v3777abf = hbusreq0 & v376d6b2 | !hbusreq0 & v376be60;
assign v376a3aa = hmaster0_p & v3a70987 | !hmaster0_p & v373026f;
assign v375586c = hmaster1_p & v377766c | !hmaster1_p & v375f0f8;
assign v372e4de = hgrant6_p & v3728d72 | !hgrant6_p & v3a6ec17;
assign v375fa7a = hmaster2_p & v3a5f8d0 | !hmaster2_p & v8455ab;
assign v3a63f9a = hmaster0_p & v372954c | !hmaster0_p & v8455ab;
assign v373f057 = hgrant5_p & v3a62a6d | !hgrant5_p & v3748eaa;
assign v3a6f626 = jx1_p & v375b61a | !jx1_p & v37384cb;
assign v3738b7e = hlock7_p & v3742dcb | !hlock7_p & !v3726ed7;
assign v3768c2e = hmaster1_p & v3777853 | !hmaster1_p & v37685bf;
assign v3750d6d = hgrant5_p & v8455ab | !hgrant5_p & !v3a6f1eb;
assign v3748d1f = hlock4 & v372dec3 | !hlock4 & v376ba2e;
assign v377e70d = hbusreq0 & v3764ad1 | !hbusreq0 & v8455ab;
assign v374525d = hbusreq0 & v377723a | !hbusreq0 & v928541;
assign v3773536 = hmaster1_p & v8455b5 | !hmaster1_p & v3a6d2d3;
assign v3a67755 = hbusreq7_p & v3745e54 | !hbusreq7_p & v37240c0;
assign v3a67d7b = hlock7 & v374c9d1 | !hlock7 & v3a6062e;
assign v1e37a72 = hlock0 & v3a5378e | !hlock0 & v3a603ad;
assign v3758e7b = hbusreq0 & v3770769 | !hbusreq0 & v8455ab;
assign v3a703d9 = hgrant6_p & v8455ab | !hgrant6_p & v376f7ab;
assign v37750f7 = hbusreq6_p & v3a70425 | !hbusreq6_p & v8455ab;
assign v377d91c = hmaster1_p & v3a6f443 | !hmaster1_p & v3773eee;
assign v3725f48 = hbusreq3_p & v376e06b | !hbusreq3_p & v373b17c;
assign v3a63b69 = hmaster1_p & v8455ab | !hmaster1_p & v37425ab;
assign v337900b = hbusreq4 & v375153e | !hbusreq4 & v3a678d2;
assign v374c0d0 = hbusreq5_p & v372ba66 | !hbusreq5_p & v3730c3c;
assign v3722e90 = hbusreq4 & v3a6af71 | !hbusreq4 & v8455ab;
assign v376ccdf = hgrant4_p & v3a6d627 | !hgrant4_p & v3a6c7ab;
assign v3a71219 = hgrant2_p & v373dbb0 | !hgrant2_p & !v3a713ee;
assign v37370f8 = hbusreq2 & v3a67eec | !hbusreq2 & v37496fa;
assign v3a70c57 = hgrant5_p & v3736b0e | !hgrant5_p & v37611df;
assign v3a70088 = hgrant6_p & v9ed516 | !hgrant6_p & v3770f6e;
assign v374d529 = hbusreq8_p & v37421c0 | !hbusreq8_p & v375c54c;
assign v3777995 = hbusreq7_p & v3746045 | !hbusreq7_p & v3740ad9;
assign v3a6124f = hbusreq2 & v3379037 | !hbusreq2 & v8455ab;
assign v3739eed = hlock5 & v3a6fab1 | !hlock5 & v376a47b;
assign v372a94f = hmaster2_p & v3a70fd5 | !hmaster2_p & v37294d3;
assign v3a64288 = hmaster1_p & v3a6a332 | !hmaster1_p & v3a70ca8;
assign v3770072 = hlock5 & v374d7ec | !hlock5 & v374f712;
assign v37334a3 = hbusreq6_p & v3a555d7 | !hbusreq6_p & v8455ab;
assign v374d339 = hmaster2_p & v3806ff6 | !hmaster2_p & v37313e5;
assign v374ea7e = hbusreq8_p & v372ee8a | !hbusreq8_p & v2092f1b;
assign v374dfd9 = hgrant0_p & v3a57f59 | !hgrant0_p & v3a6ea51;
assign v3753ca0 = hgrant3_p & v8455ab | !hgrant3_p & v372b74c;
assign v374eef1 = hbusreq6_p & v38092b4 | !hbusreq6_p & v3a658bf;
assign v3a53f85 = hbusreq5 & v376c5af | !hbusreq5 & v3745e51;
assign v3779a88 = hbusreq4 & v375c976 | !hbusreq4 & v3a64af7;
assign v376cda5 = hmaster0_p & v373c3e1 | !hmaster0_p & v372cc01;
assign v3753927 = hmaster0_p & v3a6e31f | !hmaster0_p & v37565af;
assign v3754d82 = hmaster2_p & v3a58d22 | !hmaster2_p & v3764978;
assign v375be5b = hgrant1_p & v3766ef9 | !hgrant1_p & v375aa47;
assign v3a6f436 = locked_p & v372cb88 | !locked_p & !v8455ab;
assign v3778362 = hbusreq8 & v377eac3 | !hbusreq8 & !v37366da;
assign v373b2da = hbusreq7 & v3a70fca | !hbusreq7 & v375af91;
assign v3a6f233 = hgrant7_p & v374f048 | !hgrant7_p & v3a56f2e;
assign v3a5d417 = hmaster0_p & v37356f0 | !hmaster0_p & v3a67ab5;
assign v3a70a8a = hgrant0_p & v3a59b87 | !hgrant0_p & v3a6325a;
assign v3a663d6 = hbusreq8 & cda4f0 | !hbusreq8 & v3a63d0f;
assign v373f012 = hmaster0_p & v376e72d | !hmaster0_p & v37754e6;
assign v3763eac = hgrant3_p & v3a64f9b | !hgrant3_p & c0b4d9;
assign v3a6d958 = hbusreq4_p & v3a6dd5a | !hbusreq4_p & v8455ab;
assign v3764448 = hbusreq7 & v32587ac | !hbusreq7 & v377234d;
assign v3a714a2 = hbusreq6_p & v374faa9 | !hbusreq6_p & v37372c9;
assign v376ed91 = hgrant0_p & v35b774b | !hgrant0_p & v3a65934;
assign v376ba47 = locked_p & v3a5e24e | !locked_p & v3a619c0;
assign v2092faa = hlock0_p & v3756bc9 | !hlock0_p & v3727740;
assign v3a6843c = jx0_p & v3a710e0 | !jx0_p & v3772112;
assign v37517d2 = hbusreq6_p & v3a6867e | !hbusreq6_p & v3a6c6cf;
assign v3a6eb69 = hbusreq5_p & v3809964 | !hbusreq5_p & v3a5ba93;
assign v375af36 = hlock4 & v374a4ca | !hlock4 & v3a70791;
assign v37354b5 = hbusreq4 & v37376f9 | !hbusreq4 & v3730d6a;
assign v3725fe1 = hbusreq6_p & v3725152 | !hbusreq6_p & v3735c95;
assign v3740953 = hmaster2_p & v3723fcc | !hmaster2_p & v37786a6;
assign v3777a7f = hburst0 & v3757c6f | !hburst0 & v2092b2f;
assign v3a700b0 = hbusreq2 & v3747e8e | !hbusreq2 & v3a70b92;
assign v373b838 = hbusreq4 & v37457fb | !hbusreq4 & v8455e7;
assign v3a609bb = hbusreq2_p & v3a66d7e | !hbusreq2_p & !v35772a6;
assign v37410b9 = jx0_p & v3751bf3 | !jx0_p & v3733e04;
assign v3a6320d = hbusreq3 & v3a5600a | !hbusreq3 & v8455ab;
assign v3734930 = hlock7_p & v3738f8a | !hlock7_p & v3753e74;
assign v3758e1c = hbusreq4_p & v376574a | !hbusreq4_p & v3a69c57;
assign v372eb90 = hbusreq5 & v375671a | !hbusreq5 & v380760a;
assign v3732569 = hbusreq2_p & v3732e1b | !hbusreq2_p & v3728e09;
assign v375fc83 = hmaster2_p & v3a7142f | !hmaster2_p & v37249cc;
assign v3744fc9 = hlock4_p & v3a607af | !hlock4_p & v8455e7;
assign v3748d6c = hbusreq8 & v37401bb | !hbusreq8 & v3a704ff;
assign v373578f = hgrant8_p & v37451db | !hgrant8_p & v3a57210;
assign v3736db2 = hbusreq4_p & v3a70e3d | !hbusreq4_p & v8455ab;
assign v3768ec3 = jx0_p & v3a6909f | !jx0_p & v3738d86;
assign v3a6f9f7 = hmaster2_p & v373366b | !hmaster2_p & v3a5b978;
assign v3a71454 = hgrant6_p & v3a69487 | !hgrant6_p & v373867c;
assign v3729ee6 = hmaster0_p & v372c064 | !hmaster0_p & v3a7155c;
assign v372351f = hmaster1_p & v3a70a37 | !hmaster1_p & v3a6f3f2;
assign v3a60e5d = hbusreq7 & v374e82c | !hbusreq7 & v375d661;
assign v3774e2b = hbusreq7 & v3735a25 | !hbusreq7 & v3a6fddb;
assign v37492bc = hbusreq0 & v3768622 | !hbusreq0 & v8455ab;
assign v3743726 = hmaster2_p & v3a70374 | !hmaster2_p & v3a70891;
assign v922c1b = hgrant6_p & v375641f | !hgrant6_p & v3745a7b;
assign v3a6b60d = hgrant4_p & v37350b7 | !hgrant4_p & v377c6d0;
assign v3777f05 = hmaster0_p & v372de68 | !hmaster0_p & v3a70c8c;
assign v37380e2 = hmaster2_p & v3a5db8a | !hmaster2_p & !v377b576;
assign v3a70401 = hbusreq4_p & v3a70f20 | !hbusreq4_p & v373ad95;
assign v3a5865e = hmaster2_p & v3757765 | !hmaster2_p & v3a70e9e;
assign v3a645f6 = stateG10_1_p & v39ebac7 | !stateG10_1_p & v3737fe0;
assign v377b94e = hmaster1_p & v376e795 | !hmaster1_p & v376314e;
assign v37647fc = hmaster0_p & v374b0fb | !hmaster0_p & v3a6f134;
assign v37512c0 = hgrant4_p & v8455ab | !hgrant4_p & v37749c3;
assign v377734d = hbusreq8_p & v373f9eb | !hbusreq8_p & v372bb5d;
assign v37354da = hmaster2_p & v3a5f41b | !hmaster2_p & v8455ab;
assign v3a70d7b = hlock5 & v372a1d4 | !hlock5 & v3a63ece;
assign v3a5e02b = hgrant0_p & v3759032 | !hgrant0_p & v373da69;
assign v372efcb = hbusreq5 & v37418bf | !hbusreq5 & !v8455c2;
assign v3a6f4ee = hbusreq5_p & v3a6fe75 | !hbusreq5_p & !v3a5a805;
assign v3a56e03 = hlock5 & v3a69583 | !hlock5 & v3a5b86c;
assign v3a7151b = hmaster0_p & v3763175 | !hmaster0_p & v376a14f;
assign v3a66232 = hlock5 & v3729dea | !hlock5 & v3a60feb;
assign v37331d1 = hbusreq5_p & v8455ab | !hbusreq5_p & v3a70359;
assign v376cc23 = hgrant6_p & v377938d | !hgrant6_p & v3724200;
assign v3a6f639 = hgrant6_p & v377f09a | !hgrant6_p & v374611e;
assign v3a710c8 = hbusreq0 & v2acae4c | !hbusreq0 & v3a58dce;
assign v373c688 = hbusreq5 & v3776ae5 | !hbusreq5 & v374de73;
assign v376c841 = jx0_p & v3a558e5 | !jx0_p & v372ddea;
assign v1e382e7 = hbusreq3_p & v3a619c0 | !hbusreq3_p & v3a66110;
assign v37248e4 = hbusreq6 & v3a582d6 | !hbusreq6 & v3a6f20d;
assign v3a702bb = hbusreq6_p & v3756b78 | !hbusreq6_p & !v8455ca;
assign v372d434 = hgrant2_p & v8455ab | !hgrant2_p & v3742dc6;
assign v374020a = jx3_p & v3a6519c | !jx3_p & v3730e8f;
assign v3a6e29c = hgrant4_p & v8455ab | !hgrant4_p & v37317c4;
assign v376376a = hmaster1_p & v3a62a6d | !hmaster1_p & v3724882;
assign v3a6d4bf = hlock4 & v376b5ad | !hlock4 & v372a939;
assign v3741d11 = hbusreq5 & v3726013 | !hbusreq5 & v37438ca;
assign v3a633ca = hmaster1_p & v8455ab | !hmaster1_p & v3761950;
assign v3a6fa5c = hlock0 & v373a341 | !hlock0 & v3a6f430;
assign v3a6c2ad = hlock2 & v37543ae | !hlock2 & v37486c2;
assign v3a5c2d6 = hmaster1_p & v3a6f7d0 | !hmaster1_p & v37650d7;
assign v3724060 = hmaster0_p & v3a63ae9 | !hmaster0_p & v373058e;
assign v3a70dc1 = jx2_p & v37353be | !jx2_p & v3754ca0;
assign v372c8bc = hbusreq4 & v3777d2e | !hbusreq4 & !v3757f0d;
assign v3a6e857 = hbusreq4_p & v374f654 | !hbusreq4_p & v375a918;
assign v3a596a5 = hmaster1_p & v3760b03 | !hmaster1_p & v374d6ff;
assign v3771203 = hbusreq2_p & v38072fd | !hbusreq2_p & v372eaf0;
assign d3ed45 = hmaster0_p & v3a70fd5 | !hmaster0_p & v372a94f;
assign v3729511 = hgrant6_p & v8455ca | !hgrant6_p & v375156a;
assign v373e2d3 = hlock4 & v3749a6b | !hlock4 & v3754e78;
assign v3724394 = hbusreq4_p & v3a701c7 | !hbusreq4_p & v8455ab;
assign v37386fb = hbusreq4_p & v3a6fce1 | !hbusreq4_p & v3809127;
assign v376981e = hmaster2_p & v3776ada | !hmaster2_p & v3728230;
assign v3a70100 = hmaster0_p & v3744d99 | !hmaster0_p & v3a58d68;
assign v3a70259 = hbusreq5_p & ae5f9e | !hbusreq5_p & !v372e759;
assign v3807183 = hmaster0_p & v3754d82 | !hmaster0_p & v3a539bf;
assign v3772404 = hlock6 & v3a70df4 | !hlock6 & v3a69544;
assign v374d3b8 = hbusreq6 & v3a709d0 | !hbusreq6 & v3a6ebcc;
assign v3748900 = hburst1 & v2aca977 | !hburst1 & v3744577;
assign v377671e = hbusreq6 & v3775bd3 | !hbusreq6 & !v8455b9;
assign v376ad46 = hgrant4_p & v8455ab | !hgrant4_p & !v8455f5;
assign v3724ee0 = hgrant2_p & dbdbc5 | !hgrant2_p & v3a6e8fa;
assign v3a662a2 = hmaster1_p & v3a70fce | !hmaster1_p & v3a707cc;
assign b41a29 = hgrant2_p & v3750269 | !hgrant2_p & v3752c61;
assign v3761f22 = hgrant2_p & v3a5f50e | !hgrant2_p & v372e751;
assign v375b3f0 = hgrant6_p & v375b98c | !hgrant6_p & !v3727dd4;
assign v377c6b3 = hbusreq1_p & v3a635ea | !hbusreq1_p & v3a63621;
assign v3765a2e = hbusreq7 & v377265b | !hbusreq7 & !v3a70aa6;
assign v3a70e46 = hbusreq4_p & v37560ff | !hbusreq4_p & v3744131;
assign v3a70cf4 = hmaster0_p & v3a708c3 | !hmaster0_p & v3a71667;
assign v3a5da31 = hbusreq5_p & v375cd8c | !hbusreq5_p & !v3758a23;
assign v3a67a73 = hmaster0_p & v8455ab | !hmaster0_p & !v373bf74;
assign v376d15d = hbusreq0_p & v375863a | !hbusreq0_p & v8455ab;
assign v380a189 = hmaster0_p & v3a64320 | !hmaster0_p & v3757966;
assign v3a5f8b2 = hgrant7_p & v8455b5 | !hgrant7_p & v372a3dc;
assign v23fe10d = hbusreq2_p & v3777c39 | !hbusreq2_p & v376f938;
assign v37287be = hmaster2_p & v3a5e24e | !hmaster2_p & !v3733d6e;
assign v3a70621 = hbusreq2 & v3755bc2 | !hbusreq2 & v8455ab;
assign v3a68310 = hlock4 & v3a70e97 | !hlock4 & v3a614cb;
assign v3740c92 = hmaster2_p & v374314f | !hmaster2_p & v37737aa;
assign v3731e60 = hgrant2_p & v374068b | !hgrant2_p & v3757182;
assign v3741694 = hbusreq3 & v39a4e5f | !hbusreq3 & v374f35a;
assign v373f6f7 = hbusreq7 & v3a6a8b4 | !hbusreq7 & v373a8a1;
assign v39eb5b0 = hbusreq5 & v3a63ea7 | !hbusreq5 & v8455ab;
assign v3a6fa8e = hgrant4_p & v37432c6 | !hgrant4_p & v3a6f997;
assign v375fbef = hmaster0_p & v3753dab | !hmaster0_p & v3a70666;
assign v37533f6 = hmaster0_p & v3764f48 | !hmaster0_p & v3a5c3d3;
assign v3a6be50 = hmaster0_p & v3742f0b | !hmaster0_p & v37455cd;
assign v3743b63 = hbusreq7 & v37235fa | !hbusreq7 & v3779749;
assign v3753b70 = hmaster1_p & v38094b8 | !hmaster1_p & v374e7fa;
assign v3743327 = hmaster0_p & v3755002 | !hmaster0_p & v3739934;
assign v37793c8 = hgrant6_p & v374c91a | !hgrant6_p & v3769f88;
assign v3a64cfa = hlock4 & v3a711fc | !hlock4 & v3756057;
assign v377bf88 = hgrant4_p & v375058e | !hgrant4_p & v3756516;
assign v372f570 = hgrant6_p & v377f09a | !hgrant6_p & !v3743f5a;
assign v3a699f5 = hgrant3_p & v3a70351 | !hgrant3_p & v3a704c0;
assign v376ce77 = hbusreq0 & v372ec1c | !hbusreq0 & v8455ab;
assign v3a5bbc1 = hgrant5_p & v3a6f36f | !hgrant5_p & v372e99c;
assign v23fdbca = hbusreq3 & v3a5b213 | !hbusreq3 & v8455ab;
assign v3a588ec = hbusreq0 & v3a702a8 | !hbusreq0 & v3748f17;
assign v3755c19 = hmaster0_p & v8455ab | !hmaster0_p & v3a70eba;
assign v3a5fd54 = jx0_p & v372648f | !jx0_p & v375f238;
assign v3a6f9ff = hlock5 & v3744f48 | !hlock5 & v3766160;
assign v373dc55 = hlock5 & v3a5aa5c | !hlock5 & v38073e8;
assign v3a58924 = hlock4_p & v37556fd | !hlock4_p & v8455e7;
assign v3a70890 = hmaster2_p & v37793e4 | !hmaster2_p & v3a6f998;
assign v2092a9a = hlock5_p & v376204f | !hlock5_p & v3a6f387;
assign v377c500 = hmaster0_p & v8455ab | !hmaster0_p & v3a709b9;
assign v3722b6c = hmaster0_p & v374db8d | !hmaster0_p & v3a2a422;
assign v3739b4c = hbusreq4_p & v3730be2 | !hbusreq4_p & v8455ab;
assign v3a57ccf = hmaster2_p & v2ff9314 | !hmaster2_p & v37369b2;
assign v374950c = hbusreq4_p & v3749a32 | !hbusreq4_p & v375f1ee;
assign v3a6f6bd = hbusreq4 & v3a5a158 | !hbusreq4 & v3a62a6d;
assign v372df76 = hmaster0_p & v3754ddd | !hmaster0_p & !v8455ab;
assign v3766c86 = hmaster2_p & v375f2ba | !hmaster2_p & v8455ab;
assign v377a0d8 = hmaster0_p & v3a61a7f | !hmaster0_p & v37467be;
assign v372dd09 = hbusreq2_p & v373d78b | !hbusreq2_p & v3a6fcb9;
assign v3a60620 = hbusreq4 & v3a5fe39 | !hbusreq4 & !v3a640a0;
assign v38072fd = locked_p & v20d166d | !locked_p & v8455ab;
assign v372cdb0 = hmaster0_p & v37386c6 | !hmaster0_p & v3761d47;
assign v3744792 = hbusreq0 & v3a6f2cf | !hbusreq0 & v373dd27;
assign v372b17b = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a6fdef;
assign v3750a9c = hbusreq4_p & v3763056 | !hbusreq4_p & v8455ab;
assign v3a5e591 = hlock3_p & v375ca08 | !hlock3_p & !v2acb5a7;
assign v325b5ea = hburst0 & v37295fe | !hburst0 & v3a6046c;
assign v3775654 = hbusreq4_p & v3767a93 | !hbusreq4_p & v3a7029f;
assign v376539b = hbusreq5 & v292556b | !hbusreq5 & v3a6810b;
assign v37520b7 = hgrant5_p & v373f6b1 | !hgrant5_p & v376a5c1;
assign c6053a = hmaster0_p & v374a65c | !hmaster0_p & v3762ffa;
assign v377a2d1 = jx0_p & v3a61100 | !jx0_p & v3751b6b;
assign v3778cdb = hlock4 & v3740bb4 | !hlock4 & v375df95;
assign v3769424 = hmaster2_p & v3a6f7dd | !hmaster2_p & v375e721;
assign v372ad34 = hmaster2_p & v3755dcd | !hmaster2_p & v37564e4;
assign v3a667e7 = hbusreq6 & v377e181 | !hbusreq6 & v8455ab;
assign v375e133 = hmaster2_p & v8455ab | !hmaster2_p & v373cbf9;
assign v37597f7 = hbusreq8_p & v3a706f0 | !hbusreq8_p & v375be00;
assign v3740aa8 = hmaster3_p & v8455ab | !hmaster3_p & v3a6ef77;
assign v373aa0e = hbusreq5_p & v3a6ac33 | !hbusreq5_p & v3a6fb73;
assign v3a5406b = hbusreq8 & v375586c | !hbusreq8 & v3a6f4ab;
assign v3743690 = locked_p & v3a6ef8c | !locked_p & v373a26e;
assign v372b0cd = stateA1_p & v3a6841c | !stateA1_p & v3739e55;
assign v374c33a = hbusreq6 & v375fec7 | !hbusreq6 & v8455ab;
assign v3733d3f = hmaster0_p & v3a5918c | !hmaster0_p & v3761719;
assign v376a92f = hbusreq5_p & v3745706 | !hbusreq5_p & v38072fe;
assign v3a670e4 = hmaster2_p & v37356f0 | !hmaster2_p & v3753dab;
assign v374db79 = hlock4_p & b0c091 | !hlock4_p & !v8455ab;
assign v3777cb2 = hmaster2_p & v3807aa1 | !hmaster2_p & !v3778cf7;
assign v3774438 = hmaster2_p & v3767b70 | !hmaster2_p & v8455ab;
assign v375b349 = hlock6 & v3754777 | !hlock6 & v3723e1f;
assign v3a6df6c = hmaster1_p & v3a700c8 | !hmaster1_p & v37438ca;
assign v3a6fadd = hlock0_p & v37356ce | !hlock0_p & v3a54f04;
assign v373339b = hgrant4_p & v372f216 | !hgrant4_p & !v375e3d1;
assign v373dfff = hgrant6_p & v3a7124c | !hgrant6_p & v3a5d923;
assign v3739769 = hbusreq8_p & v37362dc | !hbusreq8_p & v3734279;
assign v376d2f4 = hlock4_p & v3a6267f | !hlock4_p & v372ab46;
assign v3758eb3 = hmaster0_p & v3a6f45b | !hmaster0_p & !v376ef9f;
assign v3a6fcd8 = hgrant5_p & v8455ab | !hgrant5_p & v3808eb7;
assign v3756f9b = hmaster0_p & v376c902 | !hmaster0_p & v3a60fa3;
assign v37790fb = hlock4 & v37674a3 | !hlock4 & v373ab15;
assign v372ecd8 = hgrant6_p & v3a65eba | !hgrant6_p & v3741020;
assign v3a5e09d = hbusreq3_p & v374578a | !hbusreq3_p & v3754c2d;
assign v37571c5 = hmaster2_p & v3a60b2e | !hmaster2_p & v372346b;
assign v3a6f556 = hmaster0_p & v375f15c | !hmaster0_p & !v3726991;
assign v375dba4 = hlock0 & v37512f3 | !hlock0 & v37512dc;
assign v377316f = hbusreq5_p & v1e37a8d | !hbusreq5_p & v3a7096d;
assign v3a60205 = hgrant1_p & v3762de1 | !hgrant1_p & !v8455e7;
assign v377cfd9 = hlock0_p & v3809adf | !hlock0_p & v37528b0;
assign v3a5b841 = hlock6 & v3731a3b | !hlock6 & v373d4fc;
assign v3a649c2 = hmaster3_p & v37414be | !hmaster3_p & v3a681f5;
assign v3a6107c = hlock5 & v377de7f | !hlock5 & v3a70854;
assign v3a6ec06 = hbusreq0_p & v372dadb | !hbusreq0_p & v3775bf6;
assign v3774e64 = hbusreq1_p & d0a687 | !hbusreq1_p & !v8455ab;
assign v3a558e5 = hbusreq8_p & v37c025b | !hbusreq8_p & v3a29814;
assign v93c94e = hbusreq5 & v37795d9 | !hbusreq5 & v8455ab;
assign v3a575a5 = hgrant5_p & v3744f6f | !hgrant5_p & v3a713d1;
assign v3a550c2 = hlock5_p & v3a5beb8 | !hlock5_p & !v8455ab;
assign v3a568f7 = locked_p & v3a6885a | !locked_p & v8455ab;
assign v3a64539 = hlock7 & v3a5f6a8 | !hlock7 & v37745e9;
assign v3779403 = hmaster0_p & v37798da | !hmaster0_p & v3a5cf5e;
assign v3724ced = hbusreq5_p & v3a6f3f0 | !hbusreq5_p & v37245a1;
assign v9aea50 = hgrant6_p & v8455ca | !hgrant6_p & v3a6f1ae;
assign v3735a7f = hbusreq7 & v3765998 | !hbusreq7 & v375b801;
assign v3a6ec0e = hbusreq8_p & v377d23c | !hbusreq8_p & v3a667d2;
assign v3a715ae = hbusreq6 & v372c903 | !hbusreq6 & v38072fd;
assign v3a69529 = hlock3_p & v1e37915 | !hlock3_p & !v8455ab;
assign v3a71291 = hmaster2_p & v375649e | !hmaster2_p & v3a5d5a4;
assign v3750aea = hbusreq2 & v3a6c23b | !hbusreq2 & v3a70cdb;
assign v376c02d = hbusreq2 & v373cd16 | !hbusreq2 & v8455ab;
assign v3753903 = hlock0 & v3809ec3 | !hlock0 & v3764a07;
assign v373b91e = hmaster1_p & v377296d | !hmaster1_p & v3744fb6;
assign v377de56 = hmaster1_p & v3778c64 | !hmaster1_p & v3a6073f;
assign v3a59fd0 = hgrant8_p & v8455d2 | !hgrant8_p & v37317b4;
assign v374ba3c = hlock8_p & v3a70713 | !hlock8_p & v39eb56d;
assign v3732c51 = hbusreq4_p & v37796c6 | !hbusreq4_p & v38073b0;
assign v3a6ebe2 = hmaster0_p & v8455ab | !hmaster0_p & !v3a714c7;
assign v3724204 = hlock0_p & v8455ab | !hlock0_p & !v2aca977;
assign v377fad8 = hmaster2_p & v374f3a3 | !hmaster2_p & v3a7082d;
assign v94faa4 = hmaster0_p & adf78a | !hmaster0_p & v3a5f495;
assign v3736684 = hgrant5_p & v375c85c | !hgrant5_p & v3754c99;
assign v3735b3e = hbusreq2_p & v3764d1f | !hbusreq2_p & v8455ab;
assign v3747e8e = hbusreq3_p & v373e521 | !hbusreq3_p & v3743b9e;
assign v37742f1 = hbusreq4 & v3763398 | !hbusreq4 & v8455ab;
assign v3a5db83 = hgrant5_p & v37324e7 | !hgrant5_p & !v8455ab;
assign v373b0e7 = hmaster2_p & v373be25 | !hmaster2_p & v3728e09;
assign v372e868 = hmaster0_p & v8455e7 | !hmaster0_p & v3a6f70a;
assign v3a70c30 = hmaster2_p & v3a70d99 | !hmaster2_p & v3759379;
assign v372b931 = hlock0_p & v3733383 | !hlock0_p & v3753dab;
assign v3a70ed9 = hlock4 & v3761a96 | !hlock4 & v38097ca;
assign v3a6dd65 = hgrant3_p & v376b363 | !hgrant3_p & v374578a;
assign v3a711c3 = hbusreq7_p & d320a7 | !hbusreq7_p & v374ca2e;
assign v3a6fd5a = hgrant4_p & v3a6b7e9 | !hgrant4_p & v375a463;
assign v3a6eed9 = hmaster0_p & v377c7d3 | !hmaster0_p & v37787f5;
assign v3a57f7d = hlock8 & v3a711b4 | !hlock8 & v375be90;
assign v373905f = hbusreq1_p & v3728760 | !hbusreq1_p & v3730ca3;
assign ce378e = hlock2 & v373cf8f | !hlock2 & aa3e48;
assign v3a60a24 = hmaster2_p & v3761719 | !hmaster2_p & v3731b41;
assign v37487b0 = hlock3_p & v3a653e4 | !hlock3_p & !v8455ab;
assign v373d735 = hgrant6_p & v8455ab | !hgrant6_p & v374bdfe;
assign v3727d45 = hmaster0_p & v3a6f6d5 | !hmaster0_p & v372a520;
assign v1e3733c = hmaster0_p & v3753eb2 | !hmaster0_p & v372ba93;
assign v3750e4b = hbusreq8_p & v37523de | !hbusreq8_p & v373e792;
assign bbab81 = hbusreq2_p & v8455b0 | !hbusreq2_p & v3753dab;
assign v3725198 = hbusreq2_p & v3766f7d | !hbusreq2_p & v8455ab;
assign v37306ec = hmaster1_p & v3a6fcc9 | !hmaster1_p & v374e86a;
assign v3a6f9bf = jx0_p & v373a7b4 | !jx0_p & v375c2e6;
assign v375c621 = hmaster2_p & v372689b | !hmaster2_p & v3a69796;
assign v3756343 = hlock8_p & v373d235 | !hlock8_p & v8455ab;
assign v3748a87 = hbusreq4 & v372ae9d | !hbusreq4 & ae317f;
assign v3a5a585 = hbusreq1_p & v375a842 | !hbusreq1_p & v375ac6a;
assign v3a6eb54 = hbusreq5 & c4d63a | !hbusreq5 & v377c174;
assign dc3a01 = jx3_p & v3772f09 | !jx3_p & v3a70500;
assign v3a6332f = hbusreq7 & v3776779 | !hbusreq7 & v3767b5a;
assign v37491af = hmaster1_p & v3a65b0a | !hmaster1_p & v37629b0;
assign v3762a9c = hbusreq3_p & v37431b5 | !hbusreq3_p & v8455ab;
assign v37629b4 = hlock4 & v375ff0d | !hlock4 & v3737e04;
assign v3a71009 = hbusreq8_p & v374c98c | !hbusreq8_p & v3745e12;
assign v374e4c5 = hmaster0_p & v3739517 | !hmaster0_p & v3741bce;
assign v3a65b87 = hmaster2_p & v3a70c39 | !hmaster2_p & v3750a9c;
assign v3763b9e = hbusreq0 & v3a6f2a4 | !hbusreq0 & v3a5ab84;
assign v376f29d = hgrant4_p & v3a653e4 | !hgrant4_p & !v3a71232;
assign v373ee41 = hbusreq6 & v3767578 | !hbusreq6 & v374d4ca;
assign v374bd38 = hbusreq5 & v3a6fd64 | !hbusreq5 & !v373ec1f;
assign v97b684 = hmaster1_p & v372d35f | !hmaster1_p & v373d32e;
assign v3806821 = hbusreq6_p & v374bcb4 | !hbusreq6_p & v376acbb;
assign v3a70308 = hbusreq4_p & v3a6677e | !hbusreq4_p & v8455ab;
assign v374e1f0 = hmaster3_p & v373fe61 | !hmaster3_p & v3768734;
assign v37255a1 = hbusreq5_p & v360d2c6 | !hbusreq5_p & v3a70b19;
assign v377e8be = hlock1_p & v376e914 | !hlock1_p & !v3a658bf;
assign v373dec1 = hlock2 & v38072fd | !hlock2 & v3753b5e;
assign v3749e48 = hlock3 & v3751831 | !hlock3 & v3763d3a;
assign v3a6a76d = hbusreq8 & v3758892 | !hbusreq8 & v3a70242;
assign v37526af = hgrant4_p & v373af21 | !hgrant4_p & v3a62fc4;
assign v3a571fd = hlock4 & v3757091 | !hlock4 & v3753d51;
assign v3732b3c = hmaster0_p & v3766b94 | !hmaster0_p & v377ea20;
assign v373894a = hlock5 & v3a6f621 | !hlock5 & v3755c19;
assign v337947a = hbusreq1 & v373f06b | !hbusreq1 & v8455e7;
assign v3a6df5a = hbusreq3_p & v3a54344 | !hbusreq3_p & v8455ab;
assign v3739faf = hbusreq0_p & v376430b | !hbusreq0_p & v376653d;
assign v3a603fc = hgrant4_p & v3a53eeb | !hgrant4_p & v3a62550;
assign v3a5cf6f = hlock7 & v3a679fd | !hlock7 & v374d612;
assign v3a6f573 = hlock5 & v3a7013a | !hlock5 & v3a5f451;
assign v37524b4 = hbusreq5 & v3746200 | !hbusreq5 & v3773f2b;
assign v3a6f5ea = hlock0_p & v374f87c | !hlock0_p & v3770fb6;
assign v375a4b3 = hbusreq3 & v3a6f586 | !hbusreq3 & !v3a6f3cf;
assign v3730bf9 = hlock6 & v37501ad | !hlock6 & v3a6f49e;
assign v3a711ab = hbusreq5 & v3770367 | !hbusreq5 & v37494ce;
assign v3a6fab5 = hbusreq3_p & v35b9d52 | !hbusreq3_p & v3733ea2;
assign v3a590d1 = hbusreq5_p & v372bc0c | !hbusreq5_p & v375237c;
assign v3a59f74 = hlock3_p & aefb3e | !hlock3_p & v372e59e;
assign v3731f7a = hgrant6_p & v3a705bf | !hgrant6_p & v37610f8;
assign v92e6f3 = hgrant4_p & v377e618 | !hgrant4_p & v3751cc4;
assign v372f56c = hmaster1_p & v3a635ea | !hmaster1_p & v3a5f0a5;
assign v3737143 = hlock8 & v3737808 | !hlock8 & v376a94b;
assign v3727bcb = hlock0 & v1e37bf6 | !hlock0 & v374f7ec;
assign v3a7062b = hgrant2_p & b0f188 | !hgrant2_p & v374fae5;
assign v376530c = hmaster1_p & bc3d4a | !hmaster1_p & v3736358;
assign ac8c4a = hlock7 & v377e31d | !hlock7 & v37499ac;
assign v3771656 = hbusreq2_p & v3a6f918 | !hbusreq2_p & v3744fbb;
assign v373a29c = hgrant2_p & v8c4a86 | !hgrant2_p & v37c0190;
assign v37684cf = hbusreq3 & v375e6b3 | !hbusreq3 & v8455ab;
assign v3769740 = hgrant4_p & v8455c2 | !hgrant4_p & v380919d;
assign v375b445 = hbusreq2 & v3a676d6 | !hbusreq2 & v8455ab;
assign v376c7d1 = hbusreq4_p & v3a62caa | !hbusreq4_p & v3a63621;
assign v37725c4 = hlock5 & v3a70854 | !hlock5 & v3755f9d;
assign v376bc9b = hgrant5_p & v3a6fc07 | !hgrant5_p & v3753900;
assign v3763571 = hlock5 & v3a6ef17 | !hlock5 & v372b50b;
assign v37756ef = hlock5_p & b77306 | !hlock5_p & v8455b7;
assign v3a63d77 = hbusreq5_p & v37709d8 | !hbusreq5_p & v37235b8;
assign v3a56f2d = hmaster1_p & v3a5e24e | !hmaster1_p & v376df3c;
assign v376c51e = hmaster1_p & v8455b0 | !hmaster1_p & v3a70d4d;
assign v3a69e59 = hmaster1_p & v37725c4 | !hmaster1_p & v8455ab;
assign v3754b83 = hgrant6_p & v3a6eeef | !hgrant6_p & v3a5b774;
assign v372dbe1 = hbusreq8 & v373172e | !hbusreq8 & v3729555;
assign v373e712 = hmaster1_p & v3740d05 | !hmaster1_p & v37242b9;
assign v3a6b18b = hlock0 & v3748797 | !hlock0 & v3748560;
assign v3724974 = hbusreq7 & v3a6177b | !hbusreq7 & v3776337;
assign v3752400 = hbusreq2 & v3a67603 | !hbusreq2 & v3a6f949;
assign v3a5fe9e = hgrant4_p & v3a7048e | !hgrant4_p & v3a56f9f;
assign v373b7f5 = hgrant1_p & v37502b7 | !hgrant1_p & v3809adf;
assign v3808f3c = hbusreq7_p & v376d892 | !hbusreq7_p & v3a71239;
assign v38067ba = jx0_p & v374c256 | !jx0_p & v3a71593;
assign v3739f0e = hbusreq0 & v3748f03 | !hbusreq0 & v2aca783;
assign v3776f2c = hbusreq5_p & v37763b2 | !hbusreq5_p & v374a369;
assign v37614c8 = hgrant0_p & v374306c | !hgrant0_p & v374db93;
assign v3757194 = hbusreq8 & v3a626d4 | !hbusreq8 & v3a713f6;
assign v377d821 = hbusreq4_p & v3731f7a | !hbusreq4_p & v3724fe7;
assign v3a6f154 = hbusreq8 & v3756780 | !hbusreq8 & v3774859;
assign v373d41a = hgrant6_p & v374c91a | !hgrant6_p & v3a712d6;
assign v3a592d8 = hgrant5_p & v373ad69 | !hgrant5_p & v37400d8;
assign v3a708d1 = hlock2_p & v3a2a2ee | !hlock2_p & v37c0297;
assign v372bdcf = hmaster0_p & v373c5a6 | !hmaster0_p & v375d77d;
assign v3769ba0 = hmaster1_p & v3a5a807 | !hmaster1_p & v373ce4e;
assign v8fffa6 = hlock0 & v376bade | !hlock0 & v3765219;
assign v3a67b7f = hmaster2_p & v3742995 | !hmaster2_p & v3741e54;
assign v39a5381 = hmastlock_p & v3745b85 | !hmastlock_p & v8455ab;
assign v37393f0 = hgrant1_p & v3577306 | !hgrant1_p & v372fc51;
assign v37543ae = hbusreq2 & v37486c2 | !hbusreq2 & v3a6a82a;
assign v3a6096a = hbusreq5_p & v3a707e0 | !hbusreq5_p & v3a715d9;
assign v3a5744d = hbusreq5_p & v37589e1 | !hbusreq5_p & v3758b05;
assign v3a7060a = hmaster2_p & v3a70f68 | !hmaster2_p & v3a58b20;
assign v376dad7 = hmaster2_p & v377bb3a | !hmaster2_p & adf78a;
assign v376e795 = hlock5 & v377d2bb | !hlock5 & v373c8ba;
assign v3755928 = hgrant6_p & v3a6ffb6 | !hgrant6_p & v377702c;
assign v3750f20 = hmaster0_p & v373959b | !hmaster0_p & v3a702ce;
assign v3762cf7 = hbusreq7_p & v3a5520d | !hbusreq7_p & v33789f3;
assign v23fe37e = hlock5_p & v3a6fd0c | !hlock5_p & v37720f9;
assign v3742f52 = hmaster2_p & v3775dbc | !hmaster2_p & !v3777790;
assign v3a710d1 = jx1_p & v376062b | !jx1_p & v3755898;
assign v372eaf3 = hbusreq6_p & v37535e7 | !hbusreq6_p & v37439b2;
assign v3744452 = hlock0 & v377c6b3 | !hlock0 & v375add0;
assign v37477d2 = hgrant0_p & v8455e1 | !hgrant0_p & !v3a635ff;
assign v3774d9a = hmaster2_p & v376a3fe | !hmaster2_p & v3a563af;
assign v37426ed = hgrant1_p & v373ad95 | !hgrant1_p & v3a637dd;
assign v3729a7a = hmaster2_p & v8455ab | !hmaster2_p & v3a7156d;
assign v3733e56 = hmaster1_p & v3729f64 | !hmaster1_p & v3737421;
assign v3a56898 = hgrant2_p & v373dbb0 | !hgrant2_p & !v3743eda;
assign v37291c0 = hmaster2_p & v37430e7 | !hmaster2_p & v3766ce0;
assign v3763224 = hmaster0_p & v376093b | !hmaster0_p & !v37670ac;
assign v3729ed7 = hbusreq4 & v3a61c49 | !hbusreq4 & v3a63a66;
assign v3a60a6e = hmaster2_p & v3747302 | !hmaster2_p & v3771d4f;
assign v3a5a954 = hmaster1_p & v3746ae3 | !hmaster1_p & !v8455bb;
assign v3a5b955 = hmaster0_p & v3a6604e | !hmaster0_p & v8455ab;
assign v3a6872e = hbusreq6 & v3725556 | !hbusreq6 & v3a6efad;
assign v3a5ba6d = hlock3_p & v375f046 | !hlock3_p & !v8455ab;
assign v3a6499e = hbusreq4 & v37721df | !hbusreq4 & !v8455ab;
assign v3737e21 = hbusreq2 & v37401f0 | !hbusreq2 & v8455ab;
assign v372d538 = hlock5_p & v377703d | !hlock5_p & !v8455ab;
assign v3a7162e = hgrant2_p & v3808ed4 | !hgrant2_p & v3772f4d;
assign v3a60b2e = hbusreq4_p & v3a569b7 | !hbusreq4_p & !v8455ab;
assign v3a71420 = hmaster2_p & v3a6f54d | !hmaster2_p & v3761adc;
assign v3740e5a = hbusreq0 & v3750df3 | !hbusreq0 & v8455ab;
assign v3a64f5e = hbusreq4_p & v3779924 | !hbusreq4_p & !v8455ab;
assign v375d43d = hmaster1_p & v3a70236 | !hmaster1_p & v373443d;
assign v373055b = hlock7 & v37514f1 | !hlock7 & v33790a4;
assign v3a71585 = hmaster0_p & v3a6fe72 | !hmaster0_p & v373e267;
assign v37332ca = hbusreq8_p & v3a71380 | !hbusreq8_p & v3a6ebea;
assign v3763011 = hbusreq6 & v3728e09 | !hbusreq6 & !v8455ab;
assign v3a5a2be = hgrant2_p & v8455ab | !hgrant2_p & v375647e;
assign v377dedb = hmaster2_p & v3a68793 | !hmaster2_p & v3258762;
assign v9ed516 = hbusreq1_p & db0673 | !hbusreq1_p & v8455ab;
assign v375fcab = hmaster1_p & v373a945 | !hmaster1_p & v37709ec;
assign v3a68967 = hbusreq2_p & v3a6f9c3 | !hbusreq2_p & v3a62a96;
assign v37401c2 = hmaster0_p & v375a397 | !hmaster0_p & v373025a;
assign v373e689 = hbusreq2 & v3740171 | !hbusreq2 & v8455ab;
assign v373b4e3 = hmaster2_p & v3765e79 | !hmaster2_p & v3745f9b;
assign v3a707ce = hbusreq0 & v3a697e4 | !hbusreq0 & v3758299;
assign v3746cc1 = hmaster0_p & v375e6a0 | !hmaster0_p & v377904f;
assign v3751cc4 = hbusreq0 & v374b60b | !hbusreq0 & v3a5d93f;
assign v372895b = hbusreq5_p & v37530c7 | !hbusreq5_p & v374f21c;
assign v37233a4 = hgrant1_p & v3a5e7fd | !hgrant1_p & v374e06f;
assign v3a6ad44 = hbusreq4 & v37422b5 | !hbusreq4 & !v8455ab;
assign v376681a = hbusreq4_p & v37759e3 | !hbusreq4_p & v3a626e4;
assign v3a6f7a3 = hmaster1_p & v3770f96 | !hmaster1_p & v3a68a8b;
assign v373114f = hbusreq4_p & v373cbc2 | !hbusreq4_p & v8455ab;
assign bdda12 = hgrant0_p & v3a6c5ee | !hgrant0_p & v377d8dd;
assign v3a6206d = hbusreq6_p & v377aa17 | !hbusreq6_p & !v8455ab;
assign v3a706c8 = hgrant5_p & v3a6f19b | !hgrant5_p & v37252b7;
assign v3a5dbd7 = hmaster0_p & v3738b8a | !hmaster0_p & !v8455ab;
assign v3a6fda1 = hmaster0_p & v376e87e | !hmaster0_p & v377cccb;
assign v373029d = hlock4 & v37327ee | !hlock4 & cfe9c3;
assign v37364cf = hgrant4_p & v374378e | !hgrant4_p & v3756930;
assign v376dacb = hmaster1_p & v380974c | !hmaster1_p & v3a53e45;
assign v3a57c47 = hbusreq5_p & v3729381 | !hbusreq5_p & v37625a7;
assign v3a638e9 = hgrant3_p & v3a69c6f | !hgrant3_p & v3a711c9;
assign v3a6eb33 = hbusreq6_p & v377fb00 | !hbusreq6_p & v3776e85;
assign v3a6a195 = hready & v3743b9e | !hready & v37496fa;
assign v3a623c7 = hbusreq3_p & v2092ffc | !hbusreq3_p & v3772a87;
assign v3a6ebf2 = hbusreq0 & v3757440 | !hbusreq0 & v3739849;
assign v3a70a2e = busreq_p & v372295a | !busreq_p & v8455ab;
assign v3774fa8 = stateG10_1_p & v376d327 | !stateG10_1_p & v376dc21;
assign v3a64e40 = hgrant6_p & v3755e4e | !hgrant6_p & v3a6effa;
assign v3762244 = hbusreq0_p & v375098f | !hbusreq0_p & v3a59720;
assign v360d10b = hbusreq5 & v376f56d | !hbusreq5 & v3a5dbd7;
assign v3a5f984 = hbusreq6_p & v3750dd3 | !hbusreq6_p & v3777009;
assign v3a6fa56 = hmaster3_p & v372b689 | !hmaster3_p & v8455ab;
assign v3770b89 = hgrant1_p & v3733e9e | !hgrant1_p & v1e38224;
assign v37500ae = hlock5_p & v376ccd6 | !hlock5_p & v374ac2e;
assign v3a712d4 = hmaster2_p & v942053 | !hmaster2_p & v3a69946;
assign v375269c = hgrant5_p & v3a578ef | !hgrant5_p & v3806579;
assign v3770559 = hbusreq1_p & v3722e5c | !hbusreq1_p & v35772a6;
assign v374be0c = hbusreq7 & v372fade | !hbusreq7 & !v3a6f944;
assign v9f45ca = hmaster2_p & v372342b | !hmaster2_p & v8455ab;
assign v374a9d4 = hmaster0_p & v3763863 | !hmaster0_p & !v373cde7;
assign v3a5730e = hbusreq7_p & v375320f | !hbusreq7_p & v373867a;
assign v372ac03 = hgrant2_p & v377f812 | !hgrant2_p & v3776415;
assign v377011b = hmaster0_p & v37368ce | !hmaster0_p & v3771ddb;
assign v3a6e96b = hmaster2_p & a747d7 | !hmaster2_p & v376fe6e;
assign v3742feb = hbusreq3 & v3768ecc | !hbusreq3 & v8455ab;
assign v374ec91 = hbusreq6 & v3767561 | !hbusreq6 & v8455bb;
assign v372a39a = hbusreq5 & v376430d | !hbusreq5 & v375d9df;
assign v37356ce = hbusreq1_p & v372692d | !hbusreq1_p & v376f45e;
assign v373d62f = hmaster1_p & v8455ab | !hmaster1_p & v3a6c908;
assign v3a5ddaa = hmaster0_p & v376397d | !hmaster0_p & v3a7114b;
assign v3a5a0e2 = hgrant6_p & v3a70283 | !hgrant6_p & !v37485ec;
assign v3742efa = hmaster0_p & v376a0f6 | !hmaster0_p & v374953c;
assign v3a6fb78 = hgrant0_p & v8455ab | !hgrant0_p & v3a6fbf4;
assign v3a697cc = hgrant4_p & v8455ab | !hgrant4_p & v3747fa9;
assign v3a70f80 = hbusreq3 & v3746063 | !hbusreq3 & v374b3bf;
assign v37795e0 = hbusreq8_p & v37635d6 | !hbusreq8_p & v37434bc;
assign v3729561 = hgrant2_p & v3779cf9 | !hgrant2_p & v3a6fee9;
assign v3724811 = hbusreq5 & v3a71332 | !hbusreq5 & v3a5b514;
assign v3751d33 = hmaster0_p & v374fbb6 | !hmaster0_p & !v3741bce;
assign v3723ee7 = hgrant2_p & v3733e9e | !hgrant2_p & v372949c;
assign v3a5ad4f = hbusreq5_p & v3a70b2f | !hbusreq5_p & v3a60b1b;
assign v375e60f = hbusreq1_p & v376f9a8 | !hbusreq1_p & v376d856;
assign v376f49f = hmaster2_p & v3778ed4 | !hmaster2_p & !v8455ab;
assign v3a7027a = hmaster1_p & v3757966 | !hmaster1_p & v380a189;
assign v3752e82 = hgrant5_p & v3a5cb95 | !hgrant5_p & v374a66c;
assign v3a585d3 = hmaster2_p & d44200 | !hmaster2_p & v3723b00;
assign v3378535 = hmaster1_p & v376e150 | !hmaster1_p & !v3a6f33e;
assign v37579c1 = hbusreq4_p & v3a6f922 | !hbusreq4_p & !v8455ab;
assign v375a697 = hgrant4_p & v3770559 | !hgrant4_p & v374da36;
assign v3a714e6 = hgrant1_p & v377e52e | !hgrant1_p & !v37270d9;
assign v1e37921 = hgrant0_p & v3758b3f | !hgrant0_p & ae6485;
assign v372ded7 = hmaster2_p & v377bf88 | !hmaster2_p & v374bfcf;
assign v37570db = hbusreq4 & v377b67d | !hbusreq4 & v373f0ee;
assign v374df25 = hmaster1_p & v377aaba | !hmaster1_p & v3731eca;
assign v377007d = hmaster0_p & v37355d6 | !hmaster0_p & v374677a;
assign v374da21 = hbusreq8 & v375ca45 | !hbusreq8 & v8455ab;
assign v3a6c8cc = hgrant4_p & v1e37b99 | !hgrant4_p & v3737d95;
assign v373c2e3 = hmaster1_p & v38072dc | !hmaster1_p & v3724798;
assign v372c095 = hlock4_p & v376e9b7 | !hlock4_p & v8455bb;
assign v372a6de = hlock7 & v376eb3c | !hlock7 & v3a70879;
assign v3a62f68 = hmaster3_p & v8455ab | !hmaster3_p & v3a6f391;
assign v3752115 = hmaster0_p & v3a661fe | !hmaster0_p & v3744b55;
assign v3a5beb5 = hbusreq2_p & v3739336 | !hbusreq2_p & v375c1d1;
assign v3a65bb1 = hbusreq7 & v377661b | !hbusreq7 & v3768734;
assign v374dd4c = hmaster2_p & v35772a5 | !hmaster2_p & !v3a635ea;
assign v39a4eaa = hgrant5_p & v8455ab | !hgrant5_p & v377946d;
assign v375ae0a = jx0_p & v37614a9 | !jx0_p & v373d238;
assign v37282f3 = hgrant6_p & v3768633 | !hgrant6_p & v372cdc9;
assign v3742f1b = jx1_p & v3744dda | !jx1_p & v374dae3;
assign v3733c51 = hmaster2_p & v372615f | !hmaster2_p & v3a6039a;
assign v37766fb = hmaster2_p & v3a59d5f | !hmaster2_p & v3768fe7;
assign v3756087 = hbusreq8 & v3749a46 | !hbusreq8 & v373f537;
assign v3a5732f = hbusreq5 & v3a70db3 | !hbusreq5 & v37307a7;
assign v3a64931 = hlock5_p & v3a70c85 | !hlock5_p & v3776abb;
assign b3f461 = hgrant6_p & v377f09a | !hgrant6_p & !v374b894;
assign v373a8be = hlock8_p & v374b7b2 | !hlock8_p & v8455cf;
assign v3a6ae14 = hmaster0_p & v3a635ea | !hmaster0_p & v3741a71;
assign v3724f7b = hgrant3_p & v3a5bb64 | !hgrant3_p & v3759947;
assign v3a6afcd = hmaster1_p & v37570eb | !hmaster1_p & v3778aac;
assign v23fda4e = hbusreq8 & v3747fbf | !hbusreq8 & v372f464;
assign v39a52b7 = hmaster2_p & v3771ce2 | !hmaster2_p & !v8455ab;
assign v3733d71 = hgrant6_p & v8455ab | !hgrant6_p & v3749d58;
assign v3a606d2 = hgrant5_p & v8455ab | !hgrant5_p & v375f777;
assign v3761d84 = hgrant5_p & v37418ab | !hgrant5_p & v375a513;
assign v3a6f3ae = hmaster0_p & v377b0f8 | !hmaster0_p & !v3741bce;
assign v3767b75 = hbusreq0 & v3728a6a | !hbusreq0 & v376938e;
assign v3a6ff58 = hbusreq6_p & bee241 | !hbusreq6_p & ad7e3b;
assign v3766345 = hgrant2_p & v3a70272 | !hgrant2_p & v374b8cb;
assign v3765998 = hmaster1_p & v375a0ad | !hmaster1_p & v3a70cc7;
assign v374732a = hlock3 & v3a6fbed | !hlock3 & v3a590de;
assign v3766105 = hgrant0_p & v37773a9 | !hgrant0_p & v3731e8c;
assign v3769157 = hgrant0_p & v377b6ce | !hgrant0_p & v374790d;
assign v374bd23 = hlock5_p & v375c94e | !hlock5_p & v376f017;
assign v37296a5 = hmaster0_p & v3753dab | !hmaster0_p & v3a5f495;
assign v3765b77 = hbusreq5_p & v3a70134 | !hbusreq5_p & v3737b54;
assign v3750296 = hmaster2_p & v3731210 | !hmaster2_p & v372ec78;
assign v3764a8a = hlock5_p & v377b774 | !hlock5_p & v8455bf;
assign v372d3f1 = hbusreq7 & v3a6ff70 | !hbusreq7 & v35b71fc;
assign v373db51 = hburst1_p & v8455ab | !hburst1_p & !v3a7111f;
assign v3a5de5f = hbusreq7 & v374b19b | !hbusreq7 & v3a71146;
assign v3a712e7 = hlock3_p & v8455ab | !hlock3_p & v373e21a;
assign v372e426 = hlock5_p & v3a5f4e0 | !hlock5_p & v3a7087d;
assign v3753258 = hbusreq0 & v3a69b93 | !hbusreq0 & v3a5bbec;
assign v373e1cc = hbusreq7 & v377073b | !hbusreq7 & !v3a6f234;
assign v375c573 = hbusreq5_p & v8455ab | !hbusreq5_p & v3762651;
assign v3779e72 = hmaster0_p & ca9b68 | !hmaster0_p & !v373aec4;
assign v3a5aaee = hlock4 & v3a701c3 | !hlock4 & v372879a;
assign v376b11a = hbusreq6_p & v3a70641 | !hbusreq6_p & v3733383;
assign v37741f0 = hgrant5_p & v37523f8 | !hgrant5_p & v3722bb0;
assign v3a7088a = hmaster1_p & v376d1b4 | !hmaster1_p & !v373bbb4;
assign v376073d = hbusreq2 & v377efdc | !hbusreq2 & v375c1d1;
assign v373da7d = hmaster2_p & v376d9ad | !hmaster2_p & v8455ab;
assign v3a63fd2 = hmaster0_p & v892398 | !hmaster0_p & v377904f;
assign v3a6e675 = hbusreq5_p & v8455cb | !hbusreq5_p & v3a71133;
assign v3730b15 = hmaster0_p & v3a635ea | !hmaster0_p & v3a64709;
assign v3a6fcc0 = hbusreq2_p & v3750e83 | !hbusreq2_p & v3731666;
assign v3774db3 = hbusreq5_p & v376f56d | !hbusreq5_p & v3a65b4a;
assign v373436a = jx0_p & v375df97 | !jx0_p & v8455ab;
assign v3748c34 = hbusreq3_p & v376f56d | !hbusreq3_p & v372a732;
assign v37275cf = hbusreq2_p & v3a61298 | !hbusreq2_p & v377a345;
assign v374a4d2 = hmaster2_p & v3a70b80 | !hmaster2_p & v3749ff9;
assign v372ce4b = jx0_p & v3a71523 | !jx0_p & v3759b61;
assign v3756018 = hgrant6_p & v3771b2c | !hgrant6_p & v3755c8b;
assign v377e2a4 = hbusreq4 & v374ccb7 | !hbusreq4 & v8455ab;
assign v3808d85 = hbusreq5 & v3a56f0b | !hbusreq5 & v3a61d5b;
assign v372e8d8 = hbusreq0 & v3767f06 | !hbusreq0 & v377205d;
assign v37686c7 = hmaster2_p & v8455ab | !hmaster2_p & !v377b576;
assign v375f97d = hbusreq7_p & v3a5df33 | !hbusreq7_p & v3a539c3;
assign v3a6ef06 = hgrant4_p & v8455ab | !hgrant4_p & v37748f0;
assign v3a70716 = hmaster2_p & v37651c2 | !hmaster2_p & v372348c;
assign v360c1bf = hbusreq4 & cfe9c3 | !hbusreq4 & v37651c2;
assign v375e037 = hmaster0_p & v374bece | !hmaster0_p & v376132a;
assign v375d832 = hmaster2_p & v3a661fe | !hmaster2_p & v3a5be93;
assign v377b61e = hmaster3_p & v3a6f729 | !hmaster3_p & v8455ab;
assign v374640f = hmaster0_p & v3a6605d | !hmaster0_p & v3764d26;
assign v375f302 = hlock6 & v3a704f2 | !hlock6 & v3a6fa2c;
assign v3a71381 = hmaster2_p & v3a6f32f | !hmaster2_p & v3a713c9;
assign v3753638 = hbusreq3 & v377094b | !hbusreq3 & v8455ab;
assign v3a70641 = hready & v8455ab | !hready & v8455e7;
assign v376b0fb = hgrant1_p & v3774f45 | !hgrant1_p & v375f077;
assign v372cdd4 = hbusreq8 & v3a6f600 | !hbusreq8 & v376ae9f;
assign v376b6c8 = hlock4_p & v3a6ac26 | !hlock4_p & v8455ab;
assign v3a6d34c = hmaster1_p & v376d876 | !hmaster1_p & v8455ab;
assign v377459d = hbusreq6_p & v3764d9e | !hbusreq6_p & v376b3bc;
assign v3a6ef4c = hbusreq6_p & v372391f | !hbusreq6_p & !v375c5a8;
assign v20930fa = hbusreq7 & v376d6d9 | !hbusreq7 & v8455ab;
assign v3a6fb73 = hmaster0_p & v3a571fa | !hmaster0_p & v373d43a;
assign v377a27c = hlock5 & v375c4b0 | !hlock5 & v35b9d58;
assign v376f5fb = stateA1_p & v8455ab | !stateA1_p & !v372fc17;
assign v3a57b0d = hbusreq3_p & v2092ffc | !hbusreq3_p & v372842d;
assign v3758ab0 = hgrant4_p & v3762502 | !hgrant4_p & v3725799;
assign v3a6f194 = hlock7 & v360d105 | !hlock7 & v3772b81;
assign v3773838 = hmaster0_p & v3a6eebd | !hmaster0_p & v3a7074e;
assign v3a7158f = hbusreq0 & v3778454 | !hbusreq0 & v3a6e5e8;
assign v3a53d2b = hbusreq8 & v3a70442 | !hbusreq8 & v374757c;
assign v3a6f123 = hgrant5_p & v3a70578 | !hgrant5_p & v3a71055;
assign v377ce00 = hbusreq1 & v3a5600a | !hbusreq1 & v373b3fb;
assign v3808cee = hgrant3_p & v373447d | !hgrant3_p & !v8455ab;
assign v3a703b9 = hlock2 & v3727703 | !hlock2 & v3a6ad59;
assign v376430b = locked_p & v3a5f308 | !locked_p & v8455ab;
assign v37341bc = hbusreq1_p & v37286bb | !hbusreq1_p & v3a70c66;
assign ccdd71 = hbusreq1_p & v377dc15 | !hbusreq1_p & !v377913f;
assign v3a57c0b = hgrant6_p & v377297e | !hgrant6_p & !v8455ab;
assign v374d9b7 = hbusreq5_p & v3a71015 | !hbusreq5_p & v372fe3c;
assign v3732d4b = hburst1 & v3a6ac2a | !hburst1 & v3a5b850;
assign v3a5e846 = hmaster2_p & v3a635ea | !hmaster2_p & v3753258;
assign v375995f = hgrant4_p & v8455ab | !hgrant4_p & v37750c2;
assign v374e1dc = hmaster2_p & v3a70c8c | !hmaster2_p & v3a66387;
assign v376b2a3 = hbusreq5 & v3730e01 | !hbusreq5 & v8455ab;
assign v3728621 = hbusreq6_p & v3a7030f | !hbusreq6_p & v3732759;
assign v375b7bd = hbusreq3_p & v37549e1 | !hbusreq3_p & v8455ab;
assign v377f3ba = hbusreq7_p & v37645c9 | !hbusreq7_p & v3771e26;
assign v3a6f6fe = hbusreq5_p & v3a6015c | !hbusreq5_p & v3a6c8b0;
assign v3a580e3 = hlock8_p & v3737103 | !hlock8_p & v8455ab;
assign v374b5bc = hbusreq7 & v3a626bd | !hbusreq7 & b5a5ab;
assign v373496c = hbusreq7 & v3a66724 | !hbusreq7 & v374dc3c;
assign v375c1fd = hbusreq7_p & v373d6dd | !hbusreq7_p & v3747630;
assign v3a6f8d1 = hgrant6_p & v8455ab | !hgrant6_p & v3a6dfc6;
assign v3771c59 = hbusreq3_p & v373b719 | !hbusreq3_p & !v8455ab;
assign v3a6ef60 = hbusreq8_p & v372d33c | !hbusreq8_p & v3a54519;
assign v3a656c7 = hmaster1_p & v3736d47 | !hmaster1_p & v375f0c9;
assign v3a70a08 = hbusreq2_p & v375c482 | !hbusreq2_p & v8455ab;
assign v37366ed = hlock4 & v209300d | !hlock4 & v3a70317;
assign v38063a0 = hbusreq0 & v3763150 | !hbusreq0 & v3a64af7;
assign v3746ab1 = hbusreq4_p & v37310be | !hbusreq4_p & v3a66f07;
assign v3a70da4 = hmaster2_p & v37651c2 | !hmaster2_p & v374e9c0;
assign v374b3e2 = hlock0 & v3731230 | !hlock0 & v3757c10;
assign v3739ea5 = hmaster2_p & v3a6f48c | !hmaster2_p & !v3775b82;
assign v3a5c860 = hbusreq5_p & v8455ab | !hbusreq5_p & v377efe7;
assign v3a54242 = hbusreq8_p & v3a65b3e | !hbusreq8_p & v3a5d41e;
assign v3757f45 = hgrant6_p & v8455ab | !hgrant6_p & v3770c66;
assign v3a701bf = hmaster1_p & v3749091 | !hmaster1_p & v377c977;
assign v3765d2a = hbusreq2_p & v37693a9 | !hbusreq2_p & v37491b7;
assign v3762475 = hbusreq0 & v3a6267f | !hbusreq0 & v8455ab;
assign v3757fde = hgrant2_p & v8455b9 | !hgrant2_p & v37278c2;
assign v372f747 = hgrant0_p & v3765a98 | !hgrant0_p & v3a68426;
assign v3a7076a = hmaster1_p & v3746c1d | !hmaster1_p & v3a5e7f7;
assign v3a62875 = hbusreq7_p & v37386af | !hbusreq7_p & !v375de73;
assign v37751b2 = hgrant8_p & v8455ab | !hgrant8_p & v3a6b49a;
assign v372ae4c = hgrant2_p & v377182c | !hgrant2_p & v372396a;
assign v374d409 = hgrant5_p & v3a6337a | !hgrant5_p & v377af8e;
assign v3a5b93f = hmaster1_p & v3a574fc | !hmaster1_p & !v3a55d78;
assign v373418b = hmaster2_p & v39a537f | !hmaster2_p & v3a695fc;
assign v3a6af1d = hgrant6_p & v37623b8 | !hgrant6_p & v8455ab;
assign v37578bd = hgrant6_p & v8455ca | !hgrant6_p & v3a5bda1;
assign v375917f = hbusreq3_p & v3734967 | !hbusreq3_p & !v374729b;
assign v3727da5 = jx0_p & v3767091 | !jx0_p & v8455ab;
assign v3766b5e = hbusreq6_p & v376aa5e | !hbusreq6_p & v35772a6;
assign v3769f88 = hgrant2_p & v377182c | !hgrant2_p & v37693cf;
assign v37645c9 = hbusreq8 & v3749283 | !hbusreq8 & v3774bad;
assign v3a68dfd = hgrant4_p & v3a53eeb | !hgrant4_p & v3a71513;
assign v3750178 = hbusreq3_p & v373e877 | !hbusreq3_p & v374f106;
assign v3a66593 = hbusreq0_p & v3a68c1f | !hbusreq0_p & v3a57f59;
assign v3768c01 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v376ab53;
assign v3a6f70c = hgrant6_p & v3727d95 | !hgrant6_p & v3a69b5c;
assign v3736adf = hbusreq7 & v376d3cb | !hbusreq7 & v373653b;
assign v3a5ecb9 = jx0_p & v3a69203 | !jx0_p & v375b84e;
assign v3a5d527 = hmaster0_p & v3765385 | !hmaster0_p & v8455ab;
assign v3a58980 = hmaster1_p & v3727d4c | !hmaster1_p & v373e806;
assign v3a70365 = hbusreq5_p & v38079d5 | !hbusreq5_p & v3774901;
assign v3377adc = hlock7 & v3772a27 | !hlock7 & v39ea259;
assign v3a6c672 = hbusreq3 & v37407b3 | !hbusreq3 & v3a559f0;
assign v37393cc = hlock0_p & v3779324 | !hlock0_p & v3769039;
assign v373a772 = hlock6_p & ca01e4 | !hlock6_p & v8455bb;
assign v96020f = hbusreq0_p & v376d45f | !hbusreq0_p & v3a5bf04;
assign v373adea = hbusreq7 & v325c957 | !hbusreq7 & v373049b;
assign v3a58554 = hgrant2_p & v3a5e221 | !hgrant2_p & v373df3d;
assign v3745a7b = hgrant2_p & v375641f | !hgrant2_p & !v3771026;
assign v3756cb8 = hbusreq4_p & v3a69796 | !hbusreq4_p & v3744cb5;
assign v37431eb = hlock2_p & v3a5a76b | !hlock2_p & v3773aa0;
assign v376047f = hlock0 & v373abde | !hlock0 & v377db1f;
assign v376a97b = hlock4 & v3750fbb | !hlock4 & v3a61cb2;
assign v3738be9 = hbusreq6_p & v376847d | !hbusreq6_p & v3a700f8;
assign v3a5d9bc = hgrant8_p & v8455ab | !hgrant8_p & v3a70f2a;
assign v374877e = hbusreq0 & v3a60258 | !hbusreq0 & v3752ac9;
assign v3746045 = hgrant5_p & v8455ab | !hgrant5_p & v3a5e015;
assign v377a865 = hgrant4_p & v8455ab | !hgrant4_p & v373c61e;
assign v3808e82 = hmaster2_p & v3a5c945 | !hmaster2_p & v3a6d684;
assign v374adfa = hbusreq8_p & v3a68467 | !hbusreq8_p & v373c1e4;
assign v373c01b = hbusreq3_p & v375d689 | !hbusreq3_p & v3a5bb64;
assign v3759c6c = hgrant2_p & v8455ab | !hgrant2_p & ce378e;
assign v3a70a9e = hbusreq5_p & v3738e62 | !hbusreq5_p & !v8455ab;
assign v3a53977 = hgrant5_p & v375c573 | !hgrant5_p & v3a2aed2;
assign v377faff = hgrant5_p & v373875c | !hgrant5_p & v3a6f345;
assign v372bb72 = hmaster2_p & v3a71377 | !hmaster2_p & v3a290f9;
assign v374d383 = hmaster0_p & v376f49f | !hmaster0_p & !v8455ab;
assign v3a682b1 = hlock0_p & v374f307 | !hlock0_p & v377dc0c;
assign v3732d8f = hgrant2_p & v8455ab | !hgrant2_p & v373c924;
assign v374caae = hlock6_p & v3a62072 | !hlock6_p & v8455ab;
assign ad7e3b = hgrant2_p & v3a5eadd | !hgrant2_p & v3a60638;
assign v3a5ec7a = hbusreq0 & v3754c8d | !hbusreq0 & v374518b;
assign v3a656ca = hmaster0_p & v373014d | !hmaster0_p & v3a55392;
assign v3777a07 = hmastlock_p & v373180e | !hmastlock_p & !v8455ab;
assign v3a5fc64 = hgrant7_p & v374d998 | !hgrant7_p & v3763f3f;
assign v9230c3 = hlock1_p & cc809f | !hlock1_p & v8455ab;
assign d3c22f = hgrant2_p & v3730e2a | !hgrant2_p & v3764a1c;
assign v3a5f744 = hmaster2_p & v37430e7 | !hmaster2_p & v3a5d46c;
assign v3740194 = hlock6_p & v37718fb | !hlock6_p & v3a57309;
assign v373b6ee = hlock5 & v37392e0 | !hlock5 & v3773633;
assign v3a69ed4 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f7b2;
assign v3a6ff67 = hbusreq6_p & v376e2ac | !hbusreq6_p & v8455ab;
assign v3a6b19d = hbusreq4_p & v3726a86 | !hbusreq4_p & v8455ab;
assign v375c92f = hmaster0_p & v3a58971 | !hmaster0_p & !v3775f27;
assign v3757e4a = hmaster1_p & v376740f | !hmaster1_p & v8455ab;
assign v372adb5 = hbusreq2_p & v375e2ab | !hbusreq2_p & v8455ab;
assign v380930a = hgrant3_p & v8455ab | !hgrant3_p & v3a5c27f;
assign v3a71632 = hlock6_p & v3a70d57 | !hlock6_p & v3a714e8;
assign v37332fa = hmaster0_p & v3774647 | !hmaster0_p & v3724596;
assign v3725ad3 = hmaster1_p & v37474df | !hmaster1_p & v3a6ffc0;
assign v37763c2 = hgrant6_p & v3a6f71a | !hgrant6_p & v3725564;
assign v375026b = hbusreq4_p & v1e38282 | !hbusreq4_p & v8455ab;
assign v37bfc8c = hgrant6_p & v3723430 | !hgrant6_p & v3a5b7b5;
assign v377d742 = hmaster2_p & v8455ab | !hmaster2_p & v37331ff;
assign v37379bb = hbusreq3_p & v3a70c4d | !hbusreq3_p & v8455ab;
assign v3a5bead = hgrant3_p & v3757568 | !hgrant3_p & v3a6a259;
assign v3a61388 = hbusreq8 & v3a637fd | !hbusreq8 & v3768734;
assign v3a6f76d = hgrant5_p & v8455ab | !hgrant5_p & v3771088;
assign v373ae1e = hgrant4_p & v8455ab | !hgrant4_p & v3a611be;
assign v3a709ee = hgrant4_p & v3751389 | !hgrant4_p & v376a39c;
assign v3a58cc0 = hburst0 & v2aca977 | !hburst0 & v375c7b6;
assign v372cf1f = hmaster2_p & v3724940 | !hmaster2_p & v8455ab;
assign v3a58306 = hlock5 & v3a7085c | !hlock5 & v3a58687;
assign v373552a = hbusreq0 & v377492b | !hbusreq0 & v8455ab;
assign v373d78f = hbusreq5 & v3a61724 | !hbusreq5 & v3a68356;
assign v3808eb7 = hmaster1_p & v374ba57 | !hmaster1_p & v376abd9;
assign v3759b71 = hbusreq0 & v3a5ffac | !hbusreq0 & v380946b;
assign v3758f3c = hbusreq1_p & v3773016 | !hbusreq1_p & v3a71208;
assign v37477d5 = hmaster3_p & v8455ab | !hmaster3_p & v372f744;
assign v3a66c2f = hbusreq6_p & v374bcfb | !hbusreq6_p & v8455ab;
assign v376df68 = hlock8 & v3a615f5 | !hlock8 & v3750857;
assign v376a11d = hmaster2_p & v37784b9 | !hmaster2_p & v3a6595f;
assign v374ab1e = hbusreq6 & v373ac39 | !hbusreq6 & v3732cb4;
assign v3723eef = hgrant6_p & v377d7a4 | !hgrant6_p & v37757e0;
assign v3736b1d = hmaster2_p & v376111d | !hmaster2_p & v3a64ee3;
assign v3a56094 = hgrant3_p & v8455ab | !hgrant3_p & v372b0f9;
assign v374db93 = hbusreq1_p & v3726277 | !hbusreq1_p & v3770d70;
assign v3a6e468 = hlock4_p & v3a6fd47 | !hlock4_p & v3a6f8f9;
assign v8455b6 = hbusreq1 & v8455ab | !hbusreq1 & !v8455ab;
assign v3723ace = hgrant6_p & v374f307 | !hgrant6_p & v3773d82;
assign v3759663 = hbusreq7 & d692cc | !hbusreq7 & v3a56918;
assign ac438c = hgrant3_p & cb9412 | !hgrant3_p & v3732f66;
assign v3a71497 = hmaster2_p & v3750e32 | !hmaster2_p & v3774cde;
assign v373adf1 = hmaster1_p & v3a5b289 | !hmaster1_p & v373cdba;
assign v373fd58 = hmaster1_p & v3a70fa3 | !hmaster1_p & v3a5a6cc;
assign v3a6fa02 = hmaster1_p & v3a6f158 | !hmaster1_p & v23fda78;
assign v3a6fc58 = hbusreq8 & v3734e23 | !hbusreq8 & a0a219;
assign v377c41b = hgrant6_p & v8455ab | !hgrant6_p & v3748d17;
assign v3a6329a = hmaster0_p & v3744d54 | !hmaster0_p & v373dbfe;
assign v3774b56 = hgrant2_p & v3a696ed | !hgrant2_p & v3a6b77d;
assign v3a6d3c9 = hmaster3_p & v8455ab | !hmaster3_p & v3778211;
assign v910050 = hgrant2_p & v8455ab | !hgrant2_p & v3807740;
assign v377e962 = jx3_p & v3a67133 | !jx3_p & v3727171;
assign v3735fc8 = hbusreq7_p & v373a1a4 | !hbusreq7_p & v377a0a1;
assign v3a62a25 = hmaster0_p & v3a56644 | !hmaster0_p & v3745b9c;
assign v3a7042d = hbusreq7_p & v372b172 | !hbusreq7_p & v3771d70;
assign v3a71646 = hgrant3_p & v3733d6e | !hgrant3_p & a21c18;
assign v3a6e868 = hlock2 & v37477dd | !hlock2 & v372da76;
assign a3cddb = hbusreq6 & v373b5d8 | !hbusreq6 & v8455ab;
assign v3751004 = hbusreq0 & v37430c6 | !hbusreq0 & v377a121;
assign v373959b = hmaster2_p & v3a6ab5f | !hmaster2_p & v3a714aa;
assign v3807a47 = hbusreq4_p & v3a6b8aa | !hbusreq4_p & v3751ab7;
assign v3a6f7e1 = hmaster1_p & v3a712e2 | !hmaster1_p & v373ee3e;
assign v3749a38 = hlock2 & v3752400 | !hlock2 & v3725f9b;
assign v3a55c44 = hbusreq7 & v372700b | !hbusreq7 & v37532cd;
assign v3a70c1b = hbusreq6 & v373ac39 | !hbusreq6 & v8455ab;
assign v3a60f1a = hlock7 & v3a572e2 | !hlock7 & v3a567ea;
assign v37322d8 = hbusreq7_p & v3a6eb88 | !hbusreq7_p & v376243f;
assign v3722b5c = hgrant5_p & v374eb3b | !hgrant5_p & v3a6f19d;
assign v90a475 = jx0_p & v3734c0f | !jx0_p & v374f749;
assign v3750a6f = hbusreq5 & v374f8da | !hbusreq5 & v3a5d644;
assign v3775311 = hgrant2_p & v3a6a213 | !hgrant2_p & !v3776d33;
assign v3a7091c = hbusreq2_p & v37693cf | !hbusreq2_p & v375b269;
assign v375887e = hbusreq4_p & v3746259 | !hbusreq4_p & v375f1ee;
assign v376b1a1 = hmaster2_p & v3768e79 | !hmaster2_p & v374e124;
assign v3a6e8b1 = hbusreq5_p & v3a70c87 | !hbusreq5_p & !v8455ab;
assign v377b5dc = hgrant5_p & v3a62fd2 | !hgrant5_p & v3a65e1a;
assign v37305b9 = hbusreq6 & v375aeca | !hbusreq6 & v3765261;
assign v3a6f4de = hbusreq4_p & v373ac67 | !hbusreq4_p & v3749b62;
assign v376f3ae = hlock8 & v3737808 | !hlock8 & v3a6f6cd;
assign v375dfcf = hmaster2_p & v3731724 | !hmaster2_p & v8455ab;
assign v3a64fee = hmaster1_p & v37432cd | !hmaster1_p & v3a60a9f;
assign v3a6f707 = hmaster2_p & v377766c | !hmaster2_p & !v3779801;
assign v3758eae = hbusreq3_p & v3761932 | !hbusreq3_p & v8455ab;
assign v3a6ff4e = hmaster0_p & v3735afb | !hmaster0_p & v3742cd4;
assign v3a5c0e1 = hmaster2_p & v372d299 | !hmaster2_p & v3a70172;
assign v3a70d07 = hmaster0_p & v3762a37 | !hmaster0_p & !v3752281;
assign v3a715cd = hbusreq5_p & v3747389 | !hbusreq5_p & v3a711d1;
assign v3a70cf2 = hmaster0_p & v37566b2 | !hmaster0_p & v372525e;
assign v3733887 = hlock2_p & v3a653e4 | !hlock2_p & !v8455ab;
assign bf5753 = hmaster0_p & v373d27f | !hmaster0_p & v3746d49;
assign v3a71065 = hlock0_p & v3809adf | !hlock0_p & v3730343;
assign v3a6589b = hbusreq4 & v3a6392b | !hbusreq4 & v8455ab;
assign v3730b84 = hbusreq8 & v3771d56 | !hbusreq8 & v8455ab;
assign v3a70041 = hlock5_p & v3a61d9f | !hlock5_p & !v8455ab;
assign v37613a8 = hgrant4_p & v8455ab | !hgrant4_p & !v3a6eebf;
assign v376cd0a = hmaster1_p & v373ad69 | !hmaster1_p & v377432b;
assign v373ad2b = hgrant4_p & v3a70ee7 | !hgrant4_p & v377594d;
assign v372f997 = hmaster2_p & v372ea51 | !hmaster2_p & v3a56ca1;
assign v3a6f7b4 = hlock5 & v3731e0e | !hlock5 & v376ea5c;
assign v3740bce = hmaster0_p & v3a6afdd | !hmaster0_p & v3809d9e;
assign v3a5be8a = hbusreq7_p & v372a7c1 | !hbusreq7_p & !v3768678;
assign v3a6c063 = hbusreq3 & v3a70385 | !hbusreq3 & !v3378ef7;
assign v372f03c = hlock7_p & v3a7078d | !hlock7_p & v3a6f98e;
assign v3a7068a = hlock4 & v3a64b0f | !hlock4 & v372e244;
assign v376f2f8 = hbusreq3_p & v3723430 | !hbusreq3_p & v8455e7;
assign v37325a2 = hbusreq4_p & v37541f4 | !hbusreq4_p & v8455ab;
assign v3a6d70a = hbusreq3_p & v374e20c | !hbusreq3_p & v8455ab;
assign v37578a2 = hgrant2_p & v8455ab | !hgrant2_p & v3779d16;
assign v372402f = hbusreq5 & v375be9f | !hbusreq5 & v8455ab;
assign v374036a = hgrant4_p & v8455ab | !hgrant4_p & v3a70dea;
assign v3a5864f = hbusreq4_p & v3739ea3 | !hbusreq4_p & v3763b0a;
assign v37773c4 = hbusreq1 & v37482f8 | !hbusreq1 & v8455ab;
assign v377d7a8 = hmaster2_p & v374158d | !hmaster2_p & v3759387;
assign v37401bb = hlock7 & v37242fa | !hlock7 & v3a5b925;
assign v374980f = hlock5_p & v3a6ff24 | !hlock5_p & !v37419b2;
assign v23fdd8d = hmaster2_p & v377d107 | !hmaster2_p & v3766a8d;
assign v3726c8d = hgrant6_p & v377e13b | !hgrant6_p & !v1e382a5;
assign v3a708fa = hlock2_p & v373c631 | !hlock2_p & v373f91b;
assign v3731ea5 = hgrant5_p & v374fd12 | !hgrant5_p & v3753a9f;
assign v3a628cf = hbusreq5_p & v3a5d96d | !hbusreq5_p & v2889706;
assign v3a7025d = hbusreq4_p & v37580d5 | !hbusreq4_p & v375c910;
assign v3a6fbf7 = hbusreq3_p & v20d166d | !hbusreq3_p & v3a53f4c;
assign v375b90a = hbusreq6 & v374f351 | !hbusreq6 & v3a5ee6e;
assign v374b429 = hgrant2_p & v3a5cfac | !hgrant2_p & v3739311;
assign v3779cc0 = hbusreq4_p & v37229c2 | !hbusreq4_p & v3a71353;
assign v3a6d5e9 = hbusreq4 & v377f5cb | !hbusreq4 & v3763104;
assign v3758c13 = hmaster0_p & v3a6eb72 | !hmaster0_p & v3770cb8;
assign v3a5a452 = hlock1_p & v3a6f81f | !hlock1_p & v3722dba;
assign v372610c = hlock5 & v376e1d4 | !hlock5 & v3735b0b;
assign v3a7116a = hmaster2_p & v8455ab | !hmaster2_p & v3725e96;
assign v376d060 = hmaster2_p & v3a54350 | !hmaster2_p & v375626c;
assign v37725d6 = hbusreq5 & v376c7f9 | !hbusreq5 & v8455ab;
assign v3751aaa = hgrant2_p & v3a69fbe | !hgrant2_p & !v8455ab;
assign v37311a4 = hbusreq2_p & v3772326 | !hbusreq2_p & v8455ab;
assign v3a56b80 = jx0_p & v377a4bd | !jx0_p & !v37650c4;
assign v373d957 = hbusreq5 & v3a625eb | !hbusreq5 & v373f08d;
assign v375bd9c = hgrant2_p & v377b6ce | !hgrant2_p & v374a9e7;
assign v375098f = hbusreq1_p & v373b7f5 | !hbusreq1_p & !v3a53f1a;
assign v3763e44 = hbusreq4_p & v3767a93 | !hbusreq4_p & v372a3af;
assign v3a7010f = hbusreq2_p & v37658af | !hbusreq2_p & v8455ab;
assign v375c652 = hbusreq8 & v372f49f | !hbusreq8 & v8455ab;
assign v373ba93 = jx0_p & v3767830 | !jx0_p & v377053a;
assign v3a6f5aa = hgrant5_p & v3763b4d | !hgrant5_p & v3735abc;
assign v37c1a73 = hmaster0_p & v3a62322 | !hmaster0_p & v8455b5;
assign v373f3ac = hlock7 & v3a68c87 | !hlock7 & v373149a;
assign v375b15b = hlock7_p & v33789ca | !hlock7_p & v8455ab;
assign v37747f8 = hgrant4_p & v8455ab | !hgrant4_p & v3a6d958;
assign v373e2e5 = hmaster2_p & v3a68848 | !hmaster2_p & v3773262;
assign v372a98e = hbusreq2 & v3a6ab5f | !hbusreq2 & !v3a6ac26;
assign v3a299c1 = stateA1_p & v3762fc4 | !stateA1_p & !v3739e55;
assign v3739c76 = hlock6_p & v374f87c | !hlock6_p & v3724940;
assign v37619dc = hlock0_p & v373905f | !hlock0_p & v3724112;
assign v3a6deec = hmaster3_p & v373553c | !hmaster3_p & v376b1ee;
assign v37461d8 = hmaster3_p & v375259d | !hmaster3_p & v373803a;
assign v3749686 = hgrant6_p & v374a664 | !hgrant6_p & v3a6f5d1;
assign v3a70831 = hgrant5_p & v377d146 | !hgrant5_p & v374072b;
assign v376a47e = hbusreq5 & v3a71427 | !hbusreq5 & v3742950;
assign v373c8ac = hbusreq5_p & v3a5a615 | !hbusreq5_p & v3a61d1f;
assign v3a6f730 = hbusreq5_p & v1e37b76 | !hbusreq5_p & v3a6eb3d;
assign v377beba = hbusreq5 & v3a5637b | !hbusreq5 & v8455ab;
assign v3a7071f = hmaster1_p & v3771e69 | !hmaster1_p & v23fd89c;
assign v3737de9 = hlock7_p & v375e566 | !hlock7_p & v3a5e998;
assign v3a64bc8 = hmaster2_p & v375e682 | !hmaster2_p & bbab81;
assign v3750fa9 = hmaster1_p & v8455ab | !hmaster1_p & v3778bb4;
assign v3733a6c = hburst0_p & v3a7111f | !hburst0_p & v3a6f056;
assign v37652d4 = hmaster2_p & v3a5d079 | !hmaster2_p & v3a71526;
assign v3a62c12 = hgrant4_p & v375e400 | !hgrant4_p & v375c845;
assign v3a6242b = hbusreq8 & v3a6f371 | !hbusreq8 & v8455ab;
assign v3a65dbb = hbusreq8_p & v3a63e51 | !hbusreq8_p & !v8455ab;
assign v38076c9 = hlock5_p & v3a5f449 | !hlock5_p & v3738bf6;
assign bd3fa8 = stateG10_1_p & v8455ab | !stateG10_1_p & v37247e2;
assign v373efee = hbusreq5 & v3a70dca | !hbusreq5 & v8455ab;
assign v3a6869f = hbusreq7 & v3743012 | !hbusreq7 & !v8455c6;
assign v3a6bd0f = hmaster1_p & v3a71585 | !hmaster1_p & !v3738eb0;
assign v3a6f1b2 = hgrant3_p & v8455be | !hgrant3_p & !v3748d3b;
assign v3a701b3 = hgrant3_p & v8455be | !hgrant3_p & !v375ef27;
assign v3a6fce5 = hbusreq6 & v375c2b1 | !hbusreq6 & v8455ab;
assign v3a5ef37 = hbusreq3_p & v3769f95 | !hbusreq3_p & v372c6fb;
assign v3a5ace5 = hlock0_p & v376f9a8 | !hlock0_p & v3a6eb66;
assign v3a6f52a = hmaster1_p & v377c174 | !hmaster1_p & v8455ab;
assign v3759f66 = hlock4 & v373d0d1 | !hlock4 & v3768288;
assign v3a6432d = hbusreq3_p & v3744752 | !hbusreq3_p & v3a70182;
assign v3a5efb2 = hlock6_p & v374f96e | !hlock6_p & v8455b7;
assign v3a5b642 = hlock8 & v3a7165e | !hlock8 & v3a6a084;
assign v376b87b = hbusreq5_p & v373700d | !hbusreq5_p & !v8455ab;
assign v3a7156c = hgrant5_p & v3a67dd8 | !hgrant5_p & v374b199;
assign v3a6b597 = hmaster2_p & v3745a5f | !hmaster2_p & v3744f62;
assign v1e3787a = hbusreq6_p & v37738d4 | !hbusreq6_p & v8455ab;
assign v3a69765 = hbusreq3 & v377b8ee | !hbusreq3 & v8455ab;
assign v380919d = hbusreq0 & v23fdaed | !hbusreq0 & v3a70d32;
assign v375f906 = hmaster0_p & v373b48c | !hmaster0_p & v3a62a6d;
assign d22727 = hgrant3_p & v3a615f7 | !hgrant3_p & v3729823;
assign v374bdcb = jx1_p & v375d41f | !jx1_p & v3a6f8a2;
assign v37316cb = hmaster0_p & v374dd4c | !hmaster0_p & !v3a635ea;
assign v372ebd5 = hmaster0_p & v3a7115e | !hmaster0_p & v3a669e9;
assign v3727b18 = hbusreq4_p & v3751e80 | !hbusreq4_p & v374673a;
assign v3a5d51a = hbusreq8_p & v3740b58 | !hbusreq8_p & v3777186;
assign v376e1c4 = hbusreq6 & v376bb04 | !hbusreq6 & v375f020;
assign v373471a = hmaster1_p & v375f071 | !hmaster1_p & v37617b9;
assign v3758e5f = hlock0_p & v37621ee | !hlock0_p & v3724c95;
assign v375913f = hgrant6_p & v37418ac | !hgrant6_p & v3a6f687;
assign v374ffb8 = hlock7 & v3a6bba4 | !hlock7 & v3a6fdf5;
assign v3a5334f = hbusreq6_p & v3a6f37f | !hbusreq6_p & v37316d9;
assign v3a66d1b = hbusreq0_p & v3a5891c | !hbusreq0_p & v376ef42;
assign v3a5c015 = hbusreq6 & v3778e03 | !hbusreq6 & v3a6a116;
assign v377681e = hmaster0_p & v3724947 | !hmaster0_p & !v373f2a6;
assign v373ecb2 = hmaster2_p & v3a70da3 | !hmaster2_p & v373a415;
assign v3a701fe = hmaster1_p & v3a6f5ae | !hmaster1_p & v8455ab;
assign v3a56187 = hbusreq2_p & v37274be | !hbusreq2_p & cc2c2e;
assign v3a6890e = hgrant4_p & v3a70827 | !hgrant4_p & v374550d;
assign v3a636a7 = hlock4 & v38072fd | !hlock4 & v3a7019a;
assign v372b607 = hmaster0_p & v35b774b | !hmaster0_p & v3a70b87;
assign v37273d7 = hbusreq3_p & v3778937 | !hbusreq3_p & v8455ab;
assign v3a70c8f = hbusreq5_p & v3a70f93 | !hbusreq5_p & !v8455ab;
assign v3763b6c = hmaster2_p & v8455ab | !hmaster2_p & !v377957e;
assign v374ef20 = hmaster0_p & v373703c | !hmaster0_p & v3a62a6d;
assign v374e82c = hmaster1_p & v375870e | !hmaster1_p & v8a7af6;
assign v374b47b = hgrant2_p & v374bf8a | !hgrant2_p & v3a6d74f;
assign v3752c4d = hbusreq0 & v37287bd | !hbusreq0 & !v8455ab;
assign v3734419 = hmaster0_p & v3753093 | !hmaster0_p & v3a6a1af;
assign v3a7031e = hmaster1_p & v376f56d | !hmaster1_p & v3777647;
assign v374e51a = hbusreq0 & v376f56d | !hbusreq0 & !v8455ab;
assign v37628f3 = hlock8 & v3737808 | !hlock8 & v37c0170;
assign v3a71128 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a6fdef;
assign v3a64bb1 = hlock7 & v372f5c5 | !hlock7 & v3a70f63;
assign v373a802 = hbusreq2 & v377c929 | !hbusreq2 & v3a6fefa;
assign v3772596 = hlock3 & v373c3e4 | !hlock3 & v372d880;
assign v374be32 = hbusreq0 & v375bdd4 | !hbusreq0 & !v3a701c2;
assign v374c23c = hbusreq3_p & v37311d6 | !hbusreq3_p & !v374f318;
assign v3762455 = hmaster2_p & v37793a4 | !hmaster2_p & v3728dc7;
assign v3a7028a = hbusreq5 & v3745db5 | !hbusreq5 & v372edf8;
assign v3a6fe7e = hmaster0_p & v377234d | !hmaster0_p & v8af425;
assign v376a3cb = hgrant5_p & v3806bd9 | !hgrant5_p & v3a6377a;
assign v3764ca7 = hmaster1_p & v3a6fe99 | !hmaster1_p & v8455e7;
assign v3a5f2c7 = hgrant6_p & v377ab1f | !hgrant6_p & v3773f4e;
assign v3a6f04a = stateA1_p & v8455ab | !stateA1_p & !v3a6f8a1;
assign v376f9d9 = hbusreq0_p & v374e35e | !hbusreq0_p & !v3a7151d;
assign v3765627 = hbusreq6_p & v3739b80 | !hbusreq6_p & !v8455ab;
assign v3756c25 = hlock2 & v374c9f0 | !hlock2 & v3a67aaa;
assign v373b5c1 = hmaster0_p & v3a5ba8f | !hmaster0_p & !v3764683;
assign v3747a36 = hmaster2_p & v377d1a3 | !hmaster2_p & !v3766ff7;
assign v3771ea2 = hbusreq7_p & v3a6fab3 | !hbusreq7_p & v376a26b;
assign v3744df8 = hgrant4_p & v37369b2 | !hgrant4_p & v377021d;
assign v3a6b68e = hbusreq5_p & v37609e3 | !hbusreq5_p & v3a5bda4;
assign cd5e35 = hmaster1_p & v376665a | !hmaster1_p & v374221c;
assign v373cb13 = jx1_p & v3768522 | !jx1_p & v373fb32;
assign v3a5561b = hgrant3_p & v372f657 | !hgrant3_p & v37655d6;
assign v376e6e2 = hmaster1_p & v3755002 | !hmaster1_p & v3a6f47f;
assign v3757d76 = hmaster0_p & v3777628 | !hmaster0_p & v3a713a7;
assign v373c404 = hmaster1_p & v3767b70 | !hmaster1_p & v3769adb;
assign v37229e0 = hmaster0_p & v3a635ea | !hmaster0_p & d438fc;
assign v3a6fb41 = hbusreq7_p & v373a58c | !hbusreq7_p & !v3767261;
assign v3753317 = hgrant2_p & v3a637dc | !hgrant2_p & v3a70286;
assign v3a70510 = hlock8 & v3a6f91b | !hlock8 & v3a579e2;
assign v3a70d97 = hbusreq5 & v8455ab | !hbusreq5 & v8455b0;
assign v3a66724 = hmaster1_p & v37430c6 | !hmaster1_p & v3727540;
assign v37270d9 = locked_p & v8455ab | !locked_p & !v1e38224;
assign v3a695f1 = hbusreq7 & v375e1de | !hbusreq7 & v3a5af68;
assign v3a6bdca = hbusreq6_p & v3777692 | !hbusreq6_p & v37370b9;
assign v3a70e90 = hbusreq8 & v3a64539 | !hbusreq8 & v3770edc;
assign v37311da = hgrant7_p & v3776479 | !hgrant7_p & v37632c3;
assign v373421c = hbusreq3 & v3a6dc08 | !hbusreq3 & v37406d2;
assign v376c89f = hmaster2_p & v377ba59 | !hmaster2_p & v3a63df4;
assign v375c90c = hbusreq5 & c4dd17 | !hbusreq5 & v3a70515;
assign v377e698 = hgrant6_p & v8455ab | !hgrant6_p & v3754940;
assign v377db8a = hbusreq6_p & v3a6fe6a | !hbusreq6_p & v3a703df;
assign v3a61724 = hmaster0_p & v377c9a1 | !hmaster0_p & v8455ab;
assign v374d037 = hburst0 & v3771ce2 | !hburst0 & v8455e1;
assign v375a55d = hbusreq7_p & v3767d4a | !hbusreq7_p & v375830c;
assign v373e154 = hbusreq4 & v3754b2c | !hbusreq4 & v375cfa5;
assign v372de8f = hmaster1_p & v380777c | !hmaster1_p & v37440e4;
assign v3777216 = hbusreq7 & v3a5fed1 | !hbusreq7 & v3a6c3ae;
assign v3779734 = hbusreq4 & v3743a66 | !hbusreq4 & v3728196;
assign v3729bd1 = hbusreq5_p & v376de00 | !hbusreq5_p & !v8455ab;
assign v376a26b = hgrant5_p & v3a608c4 | !hgrant5_p & v37518ac;
assign v37436bc = hbusreq2_p & v3723430 | !hbusreq2_p & v8455e7;
assign v3a6681e = hbusreq7 & v374d010 | !hbusreq7 & v3762db6;
assign v37730d2 = hmaster0_p & v3a70f68 | !hmaster0_p & v376ee20;
assign v3769ad5 = hmaster2_p & v8455b0 | !hmaster2_p & v373bf45;
assign v373124d = hbusreq5 & v3a6f7b3 | !hbusreq5 & v374c6b8;
assign v1e37397 = hmaster0_p & v3a65671 | !hmaster0_p & v375d2b3;
assign v3a6a02a = hbusreq5 & v3730778 | !hbusreq5 & v3a6ff12;
assign v374ff5a = hgrant6_p & v8455ab | !hgrant6_p & v3738910;
assign v373628a = hmaster3_p & v375a26b | !hmaster3_p & v3a6f058;
assign v3a6f269 = hmaster3_p & v8455ab | !hmaster3_p & v375ae0a;
assign v375c379 = hlock2_p & v3759b11 | !hlock2_p & v3a701a6;
assign v372b9d7 = hmaster0_p & v375e5bb | !hmaster0_p & v3a59905;
assign v3775aef = hbusreq6_p & v3a69b5c | !hbusreq6_p & v3733dd3;
assign v376d172 = hmaster0_p & v373d5ab | !hmaster0_p & v3748b9d;
assign v37699f2 = hlock3 & v337859c | !hlock3 & v37246f1;
assign v375929c = hmaster0_p & v3728d9c | !hmaster0_p & v374486d;
assign v376c248 = hgrant4_p & v8455c2 | !hgrant4_p & v3a54ba7;
assign v3733138 = hlock7_p & v376f14f | !hlock7_p & !v8455ab;
assign v3a6b8a2 = hbusreq3 & v23fe0bb | !hbusreq3 & v3a6c5ee;
assign v373dc73 = hbusreq6 & v8455b0 | !hbusreq6 & v373cc68;
assign v3a65e1a = hmaster1_p & v37327fe | !hmaster1_p & v3a5591a;
assign v3751734 = hbusreq1_p & v39a537f | !hbusreq1_p & !v39a5381;
assign v3a704a3 = hbusreq5_p & v372625f | !hbusreq5_p & v3755000;
assign v37733e3 = hmaster2_p & v37481e4 | !hmaster2_p & v3a700ec;
assign v374b86c = hbusreq7_p & v372dd2a | !hbusreq7_p & v35b91ba;
assign v3a6c6b1 = hbusreq5_p & v3778a97 | !hbusreq5_p & !v8455ab;
assign v9ecbe0 = hmaster2_p & v3a6fd81 | !hmaster2_p & v3766202;
assign v3a67f12 = hmaster1_p & v3a6fe0d | !hmaster1_p & v3a5dec3;
assign v376ae94 = hbusreq7 & v3741ac2 | !hbusreq7 & v3730595;
assign v3737d55 = hlock1_p & v3a655c3 | !hlock1_p & !v8455ab;
assign v374f8da = hmaster0_p & v3776ada | !hmaster0_p & v3729f41;
assign b1f79b = hbusreq8_p & v3a57913 | !hbusreq8_p & v376fe7d;
assign v3a70b7c = hbusreq4_p & v3a64190 | !hbusreq4_p & v3a5b826;
assign v38073b5 = hmaster0_p & v3a6f7dd | !hmaster0_p & v3769424;
assign v3768551 = hmaster0_p & v3747243 | !hmaster0_p & v3a69606;
assign v372a1b5 = hmaster2_p & v3753dab | !hmaster2_p & v3a704e5;
assign v375d4fa = hbusreq3_p & v37741bc | !hbusreq3_p & v37441b5;
assign v376f2f4 = hmaster3_p & v376cc0e | !hmaster3_p & !v3a66988;
assign v3771042 = hbusreq4_p & v377af47 | !hbusreq4_p & v3a5ad12;
assign v375c4ab = hmaster1_p & v3a70987 | !hmaster1_p & v3a700e9;
assign v3a6088f = hmaster1_p & v3a70a78 | !hmaster1_p & v3759b46;
assign v37507f4 = hbusreq4_p & v3a70c5d | !hbusreq4_p & v3a576d3;
assign v3a5de73 = hbusreq6 & v3a6f2bf | !hbusreq6 & v3725564;
assign v374b65e = hlock6_p & v37674c1 | !hlock6_p & v8455ab;
assign v3747c20 = hbusreq5 & v374b42b | !hbusreq5 & v374e78a;
assign v3a713ec = hbusreq4 & v3a70dbe | !hbusreq4 & v374acbe;
assign v3a612a9 = hlock6_p & b0c091 | !hlock6_p & !v8455ab;
assign v3725c6c = hbusreq5 & v3738f30 | !hbusreq5 & v3a700af;
assign v3a56644 = hmaster2_p & v8455ab | !hmaster2_p & v376f2f8;
assign v3a70fd5 = hbusreq0 & v3745f76 | !hbusreq0 & v8455ab;
assign v3a54427 = hmastlock_p & v3a6af99 | !hmastlock_p & v8455ab;
assign v37265d6 = hbusreq2_p & v372bf93 | !hbusreq2_p & v373125c;
assign v3a5b8b9 = hbusreq0 & v375ac20 | !hbusreq0 & v8455ab;
assign v372b219 = hmaster0_p & v3a5a01b | !hmaster0_p & v3a715c5;
assign v37657ef = hbusreq4 & v3757f45 | !hbusreq4 & v3a70ad6;
assign v3a6f495 = hmaster2_p & v37640e9 | !hmaster2_p & v3747d68;
assign v3a70b80 = hgrant4_p & v3a6f35c | !hgrant4_p & v3764870;
assign v1e37e4f = hmaster0_p & v376bf97 | !hmaster0_p & !v3750403;
assign v376bb43 = hmaster0_p & v376a63f | !hmaster0_p & v3a67b7f;
assign v3a70b3f = hmaster1_p & v3a7012a | !hmaster1_p & !v373bbb4;
assign v3755744 = hgrant6_p & v8455c9 | !hgrant6_p & v3746ab6;
assign v376c88f = jx0_p & v3740a1e | !jx0_p & v3749535;
assign v3a6b1ab = hbusreq5_p & v3733711 | !hbusreq5_p & !v3729ddd;
assign v372404f = hmaster2_p & v3762f51 | !hmaster2_p & v3a706f1;
assign v3a6ef2c = hmaster0_p & v3744ef1 | !hmaster0_p & d4d3bb;
assign v3747271 = hbusreq5_p & v373afe9 | !hbusreq5_p & v375aba9;
assign v3745ac6 = hbusreq4_p & v3776022 | !hbusreq4_p & v37247f2;
assign v374897d = hbusreq7_p & v372e0fc | !hbusreq7_p & v377ea1b;
assign v3a5979e = hbusreq1_p & v3769d19 | !hbusreq1_p & !v37497eb;
assign v3729829 = hbusreq2_p & v3a6eb6b | !hbusreq2_p & c0d46a;
assign v3a54b43 = hlock7_p & v377baf9 | !hlock7_p & v376c322;
assign v360c6b6 = hbusreq2 & v3a55ba9 | !hbusreq2 & v3778cdd;
assign v376a966 = hgrant5_p & v8455ab | !hgrant5_p & v3a563ed;
assign v3a6f5e8 = hlock5 & v3a6efb0 | !hlock5 & a50cea;
assign v3a577de = hmaster2_p & v37469c4 | !hmaster2_p & v3a70147;
assign v3a55723 = hbusreq2_p & v3a6a213 | !hbusreq2_p & !v373e8ad;
assign v3723614 = hlock4_p & v3732b75 | !hlock4_p & v3a6f9c3;
assign v3742afe = hmaster0_p & v3766c86 | !hmaster0_p & v374549a;
assign v3a6ead8 = hmaster2_p & v8455e1 | !hmaster2_p & !v377597f;
assign v3a6a64f = hgrant5_p & v374a35d | !hgrant5_p & v3a6973f;
assign v3a71329 = hbusreq5_p & v3a63f9a | !hbusreq5_p & v3a573d2;
assign v3a66d43 = hgrant4_p & v8455ab | !hgrant4_p & !v3a634c9;
assign v3a6fa3c = hbusreq5_p & v37731ec | !hbusreq5_p & v374e401;
assign v3775234 = hbusreq6_p & v3768c3c | !hbusreq6_p & !v374c7f4;
assign v376b734 = hbusreq3 & v37678fc | !hbusreq3 & v8455b3;
assign v374680c = hmaster1_p & v37251f1 | !hmaster1_p & v3735bbc;
assign v3a70ec7 = hmaster2_p & v3a6143b | !hmaster2_p & v3a55cd6;
assign v3a70cef = hbusreq7_p & v373e87e | !hbusreq7_p & !v8455ab;
assign v3722b10 = hmaster1_p & v375c791 | !hmaster1_p & v3a55eda;
assign bae881 = hbusreq4_p & v372874c | !hbusreq4_p & v3777955;
assign v3a700d3 = hlock8_p & v3a70a58 | !hlock8_p & v38078ea;
assign v3730052 = hbusreq4 & v3a2a33d | !hbusreq4 & v3757009;
assign v37705ec = hbusreq5_p & v3770072 | !hbusreq5_p & v3750ba3;
assign d2ccfa = hmaster0_p & v209312a | !hmaster0_p & v377ce47;
assign v377aaa9 = hbusreq7 & v3726c47 | !hbusreq7 & v3734279;
assign v3a67577 = hgrant4_p & v8455ab | !hgrant4_p & v38072f9;
assign v37463de = hbusreq6_p & v3741d99 | !hbusreq6_p & v39ebb20;
assign v373c76c = hmaster1_p & v3772f0f | !hmaster1_p & v37736b3;
assign v375df28 = hmaster1_p & v3724bf3 | !hmaster1_p & v3747271;
assign v3a6fd7e = hmaster2_p & v3723da9 | !hmaster2_p & !v3739ab6;
assign v3a67251 = hbusreq8 & v376625e | !hbusreq8 & v37391e5;
assign v3767a08 = hlock7_p & v374aab3 | !hlock7_p & v373af15;
assign v3a6cccd = hmaster2_p & v375c9f0 | !hmaster2_p & !v3760700;
assign v37605fb = hbusreq4_p & v376ca13 | !hbusreq4_p & v37562a5;
assign v3a6fbd1 = hmaster2_p & v3a59f9b | !hmaster2_p & v3758869;
assign v37381bb = hbusreq6_p & v377edba | !hbusreq6_p & !v3a5c5f4;
assign v3a6677e = hbusreq0 & v373a891 | !hbusreq0 & abddc4;
assign v372fb63 = hmaster1_p & v3758fa8 | !hmaster1_p & v3a70356;
assign v3753592 = hmaster1_p & v3a6d1ea | !hmaster1_p & v37536bf;
assign v373f5ab = hmaster2_p & v3736610 | !hmaster2_p & v2acafcc;
assign v3738844 = hmaster0_p & v3a6f164 | !hmaster0_p & v377376d;
assign v3725042 = hbusreq5_p & v3737dc7 | !hbusreq5_p & !d8fb57;
assign v3764fe1 = hlock8_p & v8455ab | !hlock8_p & !v3757858;
assign v3760ac5 = hbusreq7_p & v376f4b9 | !hbusreq7_p & v8455ab;
assign v377baf9 = hmaster1_p & v375384f | !hmaster1_p & !v3a70516;
assign v2aca977 = hmastlock_p & v373f4d3 | !hmastlock_p & v8455ab;
assign v3a70c54 = hgrant2_p & v3a6fda7 | !hgrant2_p & v35b70e6;
assign v3774055 = hmaster2_p & v376ce4d | !hmaster2_p & v3771102;
assign v373a791 = hmaster0_p & v209312a | !hmaster0_p & v3a6f195;
assign v3740546 = hbusreq4_p & v372e562 | !hbusreq4_p & v3763b0a;
assign v3a6ff8f = hlock4 & v374a115 | !hlock4 & cb1cc0;
assign v3743b2c = hbusreq5 & v3a53b8b | !hbusreq5 & v3726521;
assign v3770bc0 = hmaster2_p & v3757966 | !hmaster2_p & v3a68697;
assign v375eb99 = hmaster2_p & v3a6f9e8 | !hmaster2_p & v37799f4;
assign v3770ee4 = hbusreq8_p & v39748fd | !hbusreq8_p & v3a701b9;
assign v3a6b916 = hbusreq6_p & v372ae9d | !hbusreq6_p & !v8455ab;
assign v1e37869 = hlock3_p & v3732034 | !hlock3_p & v8455ab;
assign v374c9e4 = hlock5 & v3772318 | !hlock5 & v3a56ba2;
assign v373e750 = hmaster0_p & v3746846 | !hmaster0_p & v3809eab;
assign v3a5af82 = hbusreq2_p & v3a5fc3c | !hbusreq2_p & v3757fcc;
assign v372c6fb = hgrant0_p & v8455ab | !hgrant0_p & !v376bbe8;
assign v3a70eeb = hmaster0_p & v3a5b8b9 | !hmaster0_p & v3776c9c;
assign v3a6f456 = hburst0 & v3a6ac2a | !hburst0 & v37353c6;
assign v37381af = hmaster0_p & v3a66aa4 | !hmaster0_p & v377d19f;
assign v375c9a3 = hgrant5_p & v8455c6 | !hgrant5_p & v3724b78;
assign v23fd886 = hgrant3_p & v373e642 | !hgrant3_p & v3753186;
assign v3739c05 = hbusreq0_p & v38097fc | !hbusreq0_p & v8455ab;
assign v3756f8a = hmaster2_p & v374362e | !hmaster2_p & v3a6f7bf;
assign v373d3dd = hgrant2_p & v3750269 | !hgrant2_p & v3a7051c;
assign v3761175 = hbusreq4_p & v3a635ea | !hbusreq4_p & v372348c;
assign v3764af7 = hbusreq2 & v376fd05 | !hbusreq2 & v8455b3;
assign v3751c4c = hbusreq4_p & v8455ab | !hbusreq4_p & v374fb58;
assign v3771b2c = hbusreq6_p & v37645a4 | !hbusreq6_p & v3768d3e;
assign v3733fd0 = hmaster0_p & v37460cd | !hmaster0_p & v3759584;
assign v375d98f = hmaster3_p & v377e73f | !hmaster3_p & v3a70406;
assign v3a6fd4a = hmaster0_p & v8455ab | !hmaster0_p & !v1e37c38;
assign v375a12e = hmaster0_p & v376e7a5 | !hmaster0_p & v3a702ce;
assign v37677d8 = hbusreq2_p & v374d218 | !hbusreq2_p & v3a6fdf7;
assign v375d25d = hbusreq2 & v3748ca3 | !hbusreq2 & v373006f;
assign v91cdff = hbusreq6_p & v373be21 | !hbusreq6_p & v3806f24;
assign v375637c = hmaster0_p & v3735a94 | !hmaster0_p & !v3a5ed4a;
assign v375d05d = hlock2 & v3a5a16b | !hlock2 & v3a5617a;
assign v37685ea = hbusreq6 & v3a6f0fd | !hbusreq6 & v3a70d64;
assign v377489e = hbusreq4_p & v3a635ea | !hbusreq4_p & v377abcb;
assign v372e3e7 = hmaster0_p & v3a700b2 | !hmaster0_p & v3a711db;
assign v3a70925 = hmaster2_p & v8455ab | !hmaster2_p & v375cda2;
assign v3a70b06 = hlock0 & v3a6bf41 | !hlock0 & v3751291;
assign v37308bc = hmaster0_p & v8455e7 | !hmaster0_p & v3a6fb00;
assign v3a6f008 = hmaster2_p & v3743ff2 | !hmaster2_p & v3a712e2;
assign v3764dac = hmaster0_p & v3762158 | !hmaster0_p & v3a667cf;
assign v3723d4b = hlock4 & v3730a93 | !hlock4 & v380879c;
assign v3776756 = hlock5_p & v3759031 | !hlock5_p & v3a6efd9;
assign v3773650 = hbusreq6_p & v376f56d | !hbusreq6_p & v38099c8;
assign v3749381 = hbusreq5 & v3a64483 | !hbusreq5 & v372a6c8;
assign v375d758 = hmaster3_p & v375b344 | !hmaster3_p & v37754ac;
assign v8c34b7 = hbusreq2 & v8455e1 | !hbusreq2 & v8455ab;
assign v3a6f8c9 = hmaster2_p & v3a5e24e | !hmaster2_p & !v3a6fa93;
assign v3a7020e = hbusreq0 & v377a8e0 | !hbusreq0 & v37445e5;
assign v3a5d8e8 = hbusreq8 & v375eeaf | !hbusreq8 & v3a7160a;
assign v3a6da3b = hgrant4_p & v209310e | !hgrant4_p & v375dd29;
assign v374f557 = hbusreq6_p & v3a705de | !hbusreq6_p & !v3725f77;
assign v376195b = hgrant5_p & v3a64c14 | !hgrant5_p & v3761847;
assign v3753526 = hlock4 & v377e85a | !hlock4 & v3754e78;
assign v3746dbf = hmaster0_p & v3a70b4a | !hmaster0_p & v38087ba;
assign v3766c7b = hgrant2_p & v3752a0d | !hgrant2_p & v3a5e686;
assign v3a70e69 = hbusreq0 & v3766b27 | !hbusreq0 & v380954b;
assign v3a5aee5 = hgrant2_p & v3730e2e | !hgrant2_p & v376c235;
assign v376ff42 = hbusreq8_p & v3a5907f | !hbusreq8_p & v3770a83;
assign v37567d3 = hbusreq2 & v373e760 | !hbusreq2 & v3a57959;
assign v3a68977 = hlock8_p & v8455ab | !hlock8_p & v3777070;
assign v3a5fe2f = hgrant4_p & v8455c1 | !hgrant4_p & v3738adf;
assign v3767848 = hgrant4_p & v3759379 | !hgrant4_p & v37246a5;
assign v3a5c640 = hbusreq6_p & v3724543 | !hbusreq6_p & v8455ab;
assign v3756899 = hlock0_p & v38072fd | !hlock0_p & v3737bff;
assign v3a71137 = start_p & v8455ab | !start_p & v3a6b463;
assign v37711e2 = hgrant0_p & v8455ab | !hgrant0_p & v3a70c61;
assign v3a616fb = hbusreq5_p & v3724a65 | !hbusreq5_p & !v3750e0b;
assign v37447b4 = hbusreq5_p & v3749899 | !hbusreq5_p & v3763043;
assign v3776081 = hmaster1_p & v3a6256a | !hmaster1_p & v374610d;
assign v3a67f97 = hlock4 & v37664e7 | !hlock4 & v37266cb;
assign v373193a = hlock2 & v374b256 | !hlock2 & v3a66e70;
assign v37695e0 = hmaster1_p & v3a62a25 | !hmaster1_p & v376dce5;
assign v374fa1e = hlock8 & v3737808 | !hlock8 & v3755901;
assign v372dc20 = hlock8_p & v3a6205a | !hlock8_p & v3744539;
assign v3727a6c = hlock1_p & v3a61310 | !hlock1_p & v374d260;
assign v3754202 = hbusreq2 & v374ccb7 | !hbusreq2 & v8455ab;
assign v37726bf = hmaster1_p & v3a70f68 | !hmaster1_p & v37485e2;
assign v3749969 = hmaster2_p & v3a70374 | !hmaster2_p & v373511d;
assign v375889d = hbusreq8_p & v3a6b896 | !hbusreq8_p & v3726a09;
assign v3a5dde7 = hbusreq0 & v3a711e7 | !hbusreq0 & db9e30;
assign v3731e5c = hbusreq7_p & v3a6f7ae | !hbusreq7_p & v3767fa4;
assign v3a70099 = hmaster0_p & v374089d | !hmaster0_p & !v377e51b;
assign v3a70b55 = hgrant2_p & v3758fa7 | !hgrant2_p & v3a7028d;
assign v3a6f4cb = hmaster2_p & v33789b9 | !hmaster2_p & v3a68d2e;
assign v3764552 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a60a68;
assign v372dee5 = hmastlock_p & v3750fea | !hmastlock_p & !v8455ab;
assign v375c263 = hgrant6_p & v3a605b5 | !hgrant6_p & a61f6b;
assign v3a6af4d = hbusreq7_p & v372f96d | !hbusreq7_p & v3765ed6;
assign v3746d52 = hmaster2_p & v3a71026 | !hmaster2_p & v372d2dc;
assign v373d10a = hmaster1_p & v8455ab | !hmaster1_p & !v374d383;
assign v3728389 = hbusreq7_p & v372cd8b | !hbusreq7_p & dc33c0;
assign v3a63a46 = hlock4 & v3a5d882 | !hlock4 & v3741afa;
assign v3a6fdca = hmaster1_p & v37656be | !hmaster1_p & v3a299f8;
assign v37537ef = hgrant2_p & v3a5c700 | !hgrant2_p & v3a7047e;
assign v3723e2f = hmaster0_p & v374743d | !hmaster0_p & v372e9ef;
assign v3774664 = hbusreq8 & v3a62dae | !hbusreq8 & v3723025;
assign v3729a2a = hgrant4_p & v37510a5 | !hgrant4_p & v3768c5d;
assign v3a54aa0 = hgrant4_p & v3734967 | !hgrant4_p & v37612f7;
assign v3a6ef6e = hgrant3_p & v8455ab | !hgrant3_p & v3a55d2f;
assign v3725770 = hmaster2_p & v3766a8d | !hmaster2_p & !v8455ab;
assign v3773bbc = hbusreq4 & v3767f33 | !hbusreq4 & v8455e7;
assign v373db5d = hlock3_p & v8455ab | !hlock3_p & v39a5265;
assign v372ef16 = hlock6_p & v373b3fb | !hlock6_p & v8455b0;
assign v377fb00 = hbusreq6 & v3a5e0f7 | !hbusreq6 & v3776e85;
assign v3a67862 = hmaster0_p & v374e52d | !hmaster0_p & v3a5fd4a;
assign v3725a0b = hbusreq5_p & v374e78a | !hbusreq5_p & v3a61d1f;
assign v375ae8d = hbusreq7_p & v3748a5d | !hbusreq7_p & v3a5df82;
assign v3a70e71 = hbusreq3 & v3a5600a | !hbusreq3 & v3a299d4;
assign v376906d = hbusreq0_p & v3a66e91 | !hbusreq0_p & v38072fd;
assign v3a6e065 = hmaster2_p & v3a60787 | !hmaster2_p & v372493b;
assign v3735b0b = hmaster0_p & v3a635ea | !hmaster0_p & v3a70c75;
assign v374f8a1 = jx0_p & v3a70089 | !jx0_p & v3a6cb5b;
assign v3a6f96b = hmaster1_p & v373aaed | !hmaster1_p & v3734081;
assign v1e3751e = hbusreq5 & v3a6ae14 | !hbusreq5 & v3730b15;
assign v96c77f = hbusreq7_p & v3a70892 | !hbusreq7_p & v374af1f;
assign v3728343 = hbusreq5 & v376ac56 | !hbusreq5 & v372e3e7;
assign v3729597 = hbusreq5 & v3a689e5 | !hbusreq5 & v3764dac;
assign v373ccbc = hmaster0_p & v8455ab | !hmaster0_p & !v375789b;
assign v3a61b63 = hlock0_p & d44200 | !hlock0_p & v3a7008b;
assign v374fad8 = hmaster0_p & v3a5a28b | !hmaster0_p & v375f664;
assign v3a70822 = hgrant6_p & v377f09a | !hgrant6_p & v3a6186a;
assign v3a64ebb = hmaster0_p & be145a | !hmaster0_p & v374549a;
assign v3a6fb8b = hlock8 & v3a70d6d | !hlock8 & v3723db5;
assign v3736d3a = hgrant5_p & v3765e47 | !hgrant5_p & v3754a0d;
assign v372a13a = hlock4 & v374145b | !hlock4 & v3a70bb7;
assign v372c676 = hmaster0_p & v3a70e6a | !hmaster0_p & v3746a7e;
assign v3a6062e = hgrant5_p & v3742005 | !hgrant5_p & v3723220;
assign v3a53e5b = hbusreq4 & v3a58429 | !hbusreq4 & v3736679;
assign aca44a = hbusreq4 & v3733471 | !hbusreq4 & v8455ab;
assign v3735a71 = hbusreq4 & v373cc51 | !hbusreq4 & v8455ab;
assign v3a57baa = hmaster0_p & v375789e | !hmaster0_p & v3758d6c;
assign v3725d18 = hlock5_p & v3750d8e | !hlock5_p & v37472b9;
assign v3a6d7cd = hbusreq5 & v3a6fd3f | !hbusreq5 & v37676cd;
assign v372e40f = hlock5_p & v3a702f2 | !hlock5_p & !v2092ac3;
assign v376803b = hbusreq6 & v3735f9b | !hbusreq6 & v8455ab;
assign a5d7b0 = jx0_p & v372bee9 | !jx0_p & v8455ab;
assign v3a6ffe0 = stateG2_p & v8455ab | !stateG2_p & v3a5cf0b;
assign v3a70970 = hgrant2_p & v3759032 | !hgrant2_p & v3a2981b;
assign v37431a0 = hgrant5_p & v375cda1 | !hgrant5_p & v374620b;
assign v3779b31 = hbusreq5 & v37496fc | !hbusreq5 & aac06c;
assign v37701cf = hlock2 & v377542e | !hlock2 & v373413c;
assign v3a6b572 = hbusreq0 & v374f126 | !hbusreq0 & v373f125;
assign v3760b46 = hbusreq5 & v377521b | !hbusreq5 & v3a58c07;
assign v3a5a484 = hlock5_p & v37463d4 | !hlock5_p & v3a701f2;
assign v3a6fe8a = hgrant6_p & v8455ab | !hgrant6_p & v37535f2;
assign v376934b = hmaster1_p & v372a465 | !hmaster1_p & v3a6ffec;
assign v376871e = hgrant6_p & v8455ab | !hgrant6_p & !v3a6eff7;
assign v3a70240 = hbusreq6_p & v375cfd7 | !hbusreq6_p & v3a5cd88;
assign v372bd5e = hmaster0_p & v373c583 | !hmaster0_p & v3732c95;
assign v376fd4e = hgrant4_p & v8455ab | !hgrant4_p & v375d924;
assign v3a6376d = hmaster1_p & v3a704ca | !hmaster1_p & v3a70bee;
assign v37269a2 = hbusreq0_p & v372391f | !hbusreq0_p & !v375c5a8;
assign v372dcc0 = hmaster0_p & v37469c4 | !hmaster0_p & v373e8df;
assign v3a6fdd1 = hbusreq0 & v380974c | !hbusreq0 & !v8455ab;
assign v376ee62 = hbusreq5_p & v3a5f946 | !hbusreq5_p & v3a708d7;
assign v377d789 = hmaster0_p & v3a6e7b3 | !hmaster0_p & v3779c7e;
assign v3a299d7 = hbusreq6 & v37796c6 | !hbusreq6 & v8455ab;
assign v375d9df = hmaster0_p & v3a635ea | !hmaster0_p & v3a5e62b;
assign v375b93d = hgrant3_p & v8455ab | !hgrant3_p & v37278c8;
assign v360d2ce = hmaster2_p & v3a661fe | !hmaster2_p & v374d057;
assign v375abf4 = hmaster2_p & v3748ca3 | !hmaster2_p & v373f503;
assign v3724f1d = hmaster0_p & v372455c | !hmaster0_p & v37273b0;
assign v2aca783 = hlock0 & v3a5e2e1 | !hlock0 & v3748f03;
assign v3a6d590 = hbusreq4_p & v3a5f239 | !hbusreq4_p & v8455ab;
assign v3a6d686 = hbusreq5 & v3736113 | !hbusreq5 & v3a5e030;
assign v3776c87 = hlock5_p & v375841a | !hlock5_p & v3a6fe59;
assign v372ead6 = hbusreq4 & v37667b3 | !hbusreq4 & v37512f3;
assign v3751338 = hbusreq0 & v37297b2 | !hbusreq0 & v376022e;
assign v373d0d3 = hmaster2_p & v374f5e0 | !hmaster2_p & v38092e6;
assign v3769a62 = hbusreq7_p & v3764de1 | !hbusreq7_p & !v3a6fb3e;
assign v3771609 = hbusreq0 & v373fe74 | !hbusreq0 & a0d21b;
assign v3742e30 = hbusreq4 & v3a6f018 | !hbusreq4 & !v3a6fcba;
assign v372fb9d = hgrant3_p & v37777a2 | !hgrant3_p & v3754c2d;
assign v3731123 = hbusreq5_p & v3756031 | !hbusreq5_p & v3a5de32;
assign v3a70239 = hgrant7_p & v3762ec5 | !hgrant7_p & v377a65c;
assign v373f0a3 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v3738d63;
assign v3745bdf = hmaster2_p & v3747302 | !hmaster2_p & v3a65762;
assign v3a7039a = hbusreq4_p & v377a7e9 | !hbusreq4_p & v3a6c2a9;
assign v3a65019 = hlock5 & v377cda9 | !hlock5 & c81b97;
assign v3a5657a = hmaster3_p & v8455ab | !hmaster3_p & v3a5d474;
assign v3a706d5 = hmaster2_p & a96343 | !hmaster2_p & v3a6fac0;
assign v3a558dc = hmaster1_p & v8455ab | !hmaster1_p & v3772ab6;
assign v3731afc = hbusreq3 & d435c2 | !hbusreq3 & v372842d;
assign v3737200 = hmaster1_p & v376fbfd | !hmaster1_p & v374b074;
assign v3a6fff9 = hgrant2_p & v374d542 | !hgrant2_p & v3753ff9;
assign v374dc3c = hmaster1_p & v3754a54 | !hmaster1_p & v3a64d8f;
assign v3a5db7b = jx0_p & v374b9bb | !jx0_p & v37569b8;
assign v3753f71 = hgrant5_p & v8455c6 | !hgrant5_p & v373a438;
assign v37541f4 = hbusreq4 & v3745529 | !hbusreq4 & v8455ab;
assign beab35 = hbusreq5_p & v372630c | !hbusreq5_p & v372549f;
assign v3a70ab7 = hbusreq1_p & v3a70c73 | !hbusreq1_p & !v3a55b6c;
assign v3a5c11a = hmaster2_p & v8455ab | !hmaster2_p & v3a55773;
assign v377a577 = hmaster2_p & v3748451 | !hmaster2_p & v37318d7;
assign v3a5d1fb = hgrant3_p & v376ea4a | !hgrant3_p & v373632b;
assign v377c7d3 = hmaster2_p & v8455ab | !hmaster2_p & v3a70cee;
assign v3a6b41e = hbusreq4 & v3723e64 | !hbusreq4 & v8455ab;
assign v3a6f986 = hbusreq3 & v3a6a939 | !hbusreq3 & v8455ab;
assign v3a60ba3 = hgrant2_p & v3771203 | !hgrant2_p & v8455ab;
assign v373a972 = hgrant6_p & v3a70d99 | !hgrant6_p & v3776db6;
assign v376dd3d = hbusreq6_p & v3a6146a | !hbusreq6_p & v8455b0;
assign v3a715df = hlock5_p & v3726ea3 | !hlock5_p & v3a5605f;
assign v3a6dfdb = hmaster2_p & v375e657 | !hmaster2_p & v37598ab;
assign v3a5d644 = hmaster0_p & v8455ab | !hmaster0_p & v3729f41;
assign v3a5c41b = hbusreq5_p & v3a67dd5 | !hbusreq5_p & v3a55a75;
assign v373d97a = hmaster1_p & v3a61714 | !hmaster1_p & v3731349;
assign v376d07b = hmaster2_p & v376b81b | !hmaster2_p & v3727b0e;
assign v373b8c6 = hmaster1_p & v8455ab | !hmaster1_p & v3255a34;
assign v3771e60 = hgrant3_p & v8455ab | !hgrant3_p & v377437a;
assign v374efad = hlock7 & v3a70b52 | !hlock7 & v3756d6e;
assign v37374d6 = hlock5_p & v3a5ada9 | !hlock5_p & !v3773acc;
assign v3724e7d = hmaster2_p & v3a70d99 | !hmaster2_p & !v37234c3;
assign v3763b9b = hbusreq4_p & v3734967 | !hbusreq4_p & !v374729b;
assign v373cdea = hlock0 & v3a70a7f | !hlock0 & v23fe27f;
assign v3724fe8 = hgrant6_p & v3744cfe | !hgrant6_p & v3a6bdca;
assign v3a6efdd = hbusreq3 & v3a66aa4 | !hbusreq3 & v35b774b;
assign v3a70f78 = hbusreq6 & v3a6ff85 | !hbusreq6 & v3a70d77;
assign v3a5690f = jx1_p & v3a2a128 | !jx1_p & v372fd11;
assign v3725091 = hlock6_p & v377c7c0 | !hlock6_p & v373014d;
assign v373c441 = hgrant6_p & v3754fd2 | !hgrant6_p & v3730bf5;
assign b1fcb7 = hmaster1_p & a65142 | !hmaster1_p & be54b2;
assign v375bcf2 = hgrant6_p & v3741acc | !hgrant6_p & v375ed9f;
assign v376ce59 = hmaster1_p & v37678eb | !hmaster1_p & v372ee5a;
assign v3744990 = hbusreq7_p & v3a6f938 | !hbusreq7_p & !v3a6eb09;
assign v3a5ec2d = hbusreq2 & v3726df4 | !hbusreq2 & !v8455ab;
assign v3a7006d = hmaster0_p & v3a672a8 | !hmaster0_p & v3746a7e;
assign v37233e4 = hmaster2_p & v376f56d | !hmaster2_p & v8455ab;
assign v3766cfb = hmaster0_p & v377b66a | !hmaster0_p & v376ff64;
assign v377d4ab = hbusreq2_p & v3a6f807 | !hbusreq2_p & v372949c;
assign v3766d04 = hgrant3_p & v8455ab | !hgrant3_p & v3735580;
assign v3a6f98c = hbusreq2_p & v372e61a | !hbusreq2_p & v3a70b6e;
assign v1e37eb7 = hgrant5_p & v375dc25 | !hgrant5_p & !v3724aa4;
assign v37607a7 = hgrant4_p & v3a6eb95 | !hgrant4_p & v3a702e7;
assign v8dc5a6 = hbusreq7_p & v38068c1 | !hbusreq7_p & !v3a6aaa4;
assign v3a60836 = hmaster0_p & v3a57f59 | !hmaster0_p & v3760e51;
assign v375f030 = hburst0 & v3757c6f | !hburst0 & v3723118;
assign v3a558be = jx1_p & v3746138 | !jx1_p & v8455ab;
assign v3a70ad6 = hgrant6_p & v8455ab | !hgrant6_p & v372781d;
assign v3723ef8 = hbusreq5_p & v3732736 | !hbusreq5_p & v37523c6;
assign v3774ae5 = hbusreq5 & v376c1d6 | !hbusreq5 & v373db50;
assign v3a5473a = hmaster2_p & v374158d | !hmaster2_p & v1e37519;
assign v3762385 = hlock6 & v3a62fa7 | !hlock6 & v3a710e4;
assign v3731688 = hgrant0_p & v8455ab | !hgrant0_p & !v3a6efaa;
assign v376f175 = hbusreq6_p & v3a56e79 | !hbusreq6_p & v8455bf;
assign v3764b6e = hmaster2_p & v3a6fbf1 | !hmaster2_p & v374fe0f;
assign v373e114 = hbusreq0 & v3736679 | !hbusreq0 & v8455ab;
assign v3a66983 = hgrant3_p & v3a5e485 | !hgrant3_p & !v374910b;
assign v3a6f45a = hbusreq4_p & v39ebab4 | !hbusreq4_p & v372d967;
assign v3a59833 = hbusreq3_p & v8455ab | !hbusreq3_p & v37299b3;
assign v3a71312 = jx0_p & v373a3a7 | !jx0_p & !v3a70bdf;
assign v3761466 = hbusreq4 & v37255a7 | !hbusreq4 & v374e9c0;
assign v3758fa8 = hgrant4_p & v8455ab | !hgrant4_p & v377349f;
assign v3772935 = hgrant4_p & v375b7bd | !hgrant4_p & v377ce7d;
assign v3745d0a = hgrant5_p & v372d70c | !hgrant5_p & v3741872;
assign v3a70e84 = hbusreq3 & v376d327 | !hbusreq3 & v3a635ea;
assign a36719 = hbusreq7 & v373d26a | !hbusreq7 & v8455ab;
assign v373562f = hgrant5_p & v3a58980 | !hgrant5_p & v37548b3;
assign v3756e63 = hbusreq7_p & v377e871 | !hbusreq7_p & v373f1aa;
assign v3a70b73 = stateG10_1_p & v8455ab | !stateG10_1_p & v3756971;
assign v3757996 = hbusreq5_p & v377e904 | !hbusreq5_p & v373561e;
assign v377e033 = hlock6_p & v37681fa | !hlock6_p & v3a6f48b;
assign v3a701d7 = hbusreq2_p & v377e9a4 | !hbusreq2_p & v35772a6;
assign v373dff6 = hmaster1_p & v3a6f2d2 | !hmaster1_p & ca11a2;
assign v3754b03 = hgrant4_p & v8455c1 | !hgrant4_p & v3745ce4;
assign v3763eb0 = hbusreq8_p & v3761ac9 | !hbusreq8_p & v8455ab;
assign b4f354 = hbusreq7_p & v374c6c5 | !hbusreq7_p & !v3a70981;
assign v3a61853 = hlock3_p & v8455ab | !hlock3_p & !v2aca977;
assign v3a70398 = hbusreq5 & v3a70033 | !hbusreq5 & v3a5a1ef;
assign v3a6950d = hmaster2_p & v372e821 | !hmaster2_p & v8455ab;
assign c5ed52 = hmaster1_p & v3a669c6 | !hmaster1_p & v3a5f946;
assign v3a674ac = hlock3_p & v8455e7 | !hlock3_p & !v8455ab;
assign v3756f10 = hbusreq4_p & v3767e76 | !hbusreq4_p & v3808f6f;
assign v372b009 = hgrant5_p & v37467e9 | !hgrant5_p & v375b597;
assign v376dad0 = hlock8_p & v3a6eb8f | !hlock8_p & !v3766852;
assign cb09e1 = hlock5 & v37551c4 | !hlock5 & v3768904;
assign v3a5c196 = hlock5 & v3724028 | !hlock5 & v374ad17;
assign v377ce1c = hlock5_p & v3a704cb | !hlock5_p & v2092ac3;
assign v377cc25 = hgrant3_p & v376c72f | !hgrant3_p & !v37346be;
assign v3a6fb77 = hmaster0_p & v377b429 | !hmaster0_p & v37482c3;
assign v3731dc6 = stateG10_1_p & v8455ab | !stateG10_1_p & v2619ad0;
assign v3a6f613 = hbusreq2 & v372b7b7 | !hbusreq2 & v3a635ea;
assign v372539e = hlock4 & v372a04c | !hlock4 & v3a5548b;
assign v3a59da9 = hburst0_p & v8455ab | !hburst0_p & v3a69555;
assign v3a56c6d = hbusreq4 & v3a67967 | !hbusreq4 & v8455ab;
assign v3a6fc78 = hgrant4_p & v37354f8 | !hgrant4_p & v8455ab;
assign v3744c08 = hbusreq5 & v374f3ad | !hbusreq5 & v3a635ea;
assign v374c22d = hbusreq8_p & v3746676 | !hbusreq8_p & v8455ab;
assign v3734caf = hmaster0_p & v37617ed | !hmaster0_p & !v373bf1d;
assign v3742a62 = hbusreq6_p & v3a6fc6a | !hbusreq6_p & v376dab5;
assign v372781d = hgrant2_p & v8455ab | !hgrant2_p & v3a6a4d4;
assign v3766573 = hmaster2_p & v37526af | !hmaster2_p & v8455ab;
assign v3744593 = hmaster0_p & v3725901 | !hmaster0_p & v3a6a1af;
assign v372f4fe = hlock5 & v3724811 | !hlock5 & v3a71332;
assign v3737846 = hgrant5_p & v374fd12 | !hgrant5_p & v3730828;
assign v374aa46 = hmaster2_p & v374ad7d | !hmaster2_p & v373186a;
assign v3a70beb = hbusreq4 & v3a66606 | !hbusreq4 & v8455ab;
assign v37452e7 = hlock5_p & v375706b | !hlock5_p & v3754981;
assign v2ff9353 = hgrant8_p & v3742f7f | !hgrant8_p & v3a57646;
assign v360d029 = hmaster1_p & v3a6f96e | !hmaster1_p & !v374b36f;
assign v372313c = hgrant6_p & v8455ab | !hgrant6_p & v3a65f32;
assign v3a66dcf = hbusreq3_p & v37447bf | !hbusreq3_p & v3a6f483;
assign v3741f3c = hbusreq6_p & v3724887 | !hbusreq6_p & v375f0ba;
assign v3985138 = hgrant6_p & v8455ab | !hgrant6_p & v8455c9;
assign cea55f = hgrant4_p & v377eaf2 | !hgrant4_p & v8455ab;
assign cb9412 = hbusreq3_p & v372ba4d | !hbusreq3_p & v37480a7;
assign v3577338 = hlock6 & v3a66b88 | !hlock6 & v3778fda;
assign v3a70df6 = hmaster1_p & v37710c7 | !hmaster1_p & v35b779c;
assign v3a59548 = hbusreq0 & v3a627b3 | !hbusreq0 & v3a5a93a;
assign v3a6f1c8 = hmaster1_p & v3a700af | !hmaster1_p & v8f1dd1;
assign v3809439 = hbusreq5_p & be54b2 | !hbusreq5_p & v3a5ddc1;
assign v3a6f7b8 = hmaster1_p & v3a5c945 | !hmaster1_p & v37297c0;
assign v38099ce = hgrant3_p & v8455ab | !hgrant3_p & v3a7143f;
assign v39eb4e4 = hmaster0_p & v3a5d2f0 | !hmaster0_p & v375d4aa;
assign v3729f05 = hbusreq6 & v37574d2 | !hbusreq6 & v3a635ea;
assign b52e7d = hbusreq5_p & v3725058 | !hbusreq5_p & v376bf83;
assign v377142b = hbusreq5 & v3a705d1 | !hbusreq5 & v3764e69;
assign v37591da = hbusreq6_p & v372781d | !hbusreq6_p & v3a6fddd;
assign v3a55cc4 = hmaster2_p & v373ac1c | !hmaster2_p & v3767aae;
assign v375647e = hbusreq2_p & v3746e4e | !hbusreq2_p & v3757fcc;
assign v373485b = hmaster2_p & v3733d6e | !hmaster2_p & v3a6f312;
assign v3762100 = hbusreq5_p & v8455bf | !hbusreq5_p & v3742cd4;
assign v3a7007b = hbusreq2_p & v3732c24 | !hbusreq2_p & !v37448f2;
assign v3a700da = hgrant1_p & v3a61fc9 | !hgrant1_p & !v8455ab;
assign v372b20b = hmaster2_p & v376489b | !hmaster2_p & v373ae83;
assign v3a6d574 = hmaster2_p & v3a672c9 | !hmaster2_p & !v3a6b0c7;
assign v3750eaa = hbusreq2 & v3a7156d | !hbusreq2 & v8455ab;
assign v373a782 = hbusreq8_p & v3757066 | !hbusreq8_p & v3a66d2e;
assign v377fc4b = hbusreq6_p & v8455bb | !hbusreq6_p & v37338d8;
assign v372b418 = hmaster0_p & v372a49a | !hmaster0_p & v1e37c38;
assign v3a6f418 = hbusreq2 & v3a5cf53 | !hbusreq2 & v3a7162d;
assign v3a6f08a = hlock4 & v376d29a | !hlock4 & v3a5cd72;
assign v3754682 = hlock4 & v376c80f | !hlock4 & v39eb4cb;
assign v2092fa9 = hmaster3_p & v373fe61 | !hmaster3_p & v373c8a4;
assign v3a6dae0 = hbusreq8 & v375f938 | !hbusreq8 & v2acb0d7;
assign v3728d5a = hbusreq4 & v3a70cc3 | !hbusreq4 & v8455ab;
assign v372535d = hmaster0_p & v373a1b4 | !hmaster0_p & v373fa04;
assign v373b87c = hbusreq6_p & v3a71071 | !hbusreq6_p & v8455ab;
assign v3a6a973 = hgrant4_p & v8455ab | !hgrant4_p & v3a5d156;
assign v3736e7d = hbusreq6_p & v374a9a0 | !hbusreq6_p & v8455ab;
assign v372363e = hbusreq8_p & v3771162 | !hbusreq8_p & v3a70d99;
assign v3a538b9 = hgrant6_p & v3a61a7f | !hgrant6_p & v3a60faf;
assign v372f039 = hbusreq8_p & v372af35 | !hbusreq8_p & v8455ab;
assign v3729785 = hlock4 & v37577b6 | !hlock4 & v3a654c1;
assign v377a12e = hbusreq8_p & v3a6f569 | !hbusreq8_p & v37741f0;
assign v3742af4 = hbusreq4_p & v3a55641 | !hbusreq4_p & v3a67a85;
assign v3747edc = hmaster2_p & v3736d47 | !hmaster2_p & v372af77;
assign v374a0c4 = hmaster1_p & v3a6dc83 | !hmaster1_p & v3735274;
assign v3a70ce7 = hmaster2_p & v3a6ef01 | !hmaster2_p & v3741be8;
assign v3772616 = hbusreq8_p & v3747079 | !hbusreq8_p & v377987e;
assign v3736515 = hbusreq7 & v3a66c94 | !hbusreq7 & v3774f1e;
assign v3a5aff3 = hbusreq7 & v3a6c2d2 | !hbusreq7 & v8455b3;
assign v3807bf7 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v375d559;
assign v373afa4 = hmaster1_p & v3779060 | !hmaster1_p & v3a58640;
assign v373d032 = hbusreq4 & v376a715 | !hbusreq4 & v3a71454;
assign v3749ed5 = hmaster1_p & v3775dfb | !hmaster1_p & !v3734d9a;
assign v3756012 = hbusreq5 & v987445 | !hbusreq5 & v373de86;
assign v3744dd2 = hbusreq3_p & v37487f5 | !hbusreq3_p & !v8455ab;
assign v3a5df82 = hlock8 & v3a702e0 | !hlock8 & v3a5d99f;
assign v376013c = hmaster3_p & v376c841 | !hmaster3_p & v3753f85;
assign v3737bfb = hmaster0_p & v3a619c0 | !hmaster0_p & v3a57867;
assign v3a71263 = hbusreq3 & v3a660f2 | !hbusreq3 & v8455ab;
assign v23fe0be = hbusreq2_p & v3a6b423 | !hbusreq2_p & v8455ab;
assign v37298b2 = hmaster3_p & v8455ab | !hmaster3_p & v376d657;
assign v3731b72 = hbusreq2 & v372eaaf | !hbusreq2 & v377395f;
assign v3a6fd45 = hmaster2_p & v37795d3 | !hmaster2_p & v37745c3;
assign v3a69676 = hmaster2_p & v3a70374 | !hmaster2_p & v374b526;
assign v3764eff = hgrant5_p & v8a0a3d | !hgrant5_p & v37293e9;
assign v3733412 = hlock0_p & v3a6fdb4 | !hlock0_p & v3761224;
assign v3a71150 = hbusreq8_p & v376fc23 | !hbusreq8_p & v96c77f;
assign v372d8fa = hlock3_p & v3a62973 | !hlock3_p & !v3a704a8;
assign v3a65911 = hlock5_p & v374774a | !hlock5_p & v3a540f8;
assign v3752536 = hbusreq4 & v37583be | !hbusreq4 & !v8455ab;
assign v37269f6 = hbusreq4 & v373340d | !hbusreq4 & v3730695;
assign v374851a = hmaster0_p & v376f0f6 | !hmaster0_p & v3a6f81b;
assign v374fe65 = jx0_p & v3759ec7 | !jx0_p & v3773f70;
assign v3a5d438 = hbusreq5 & v3a63c3b | !hbusreq5 & v372f04d;
assign v372d905 = hbusreq0 & v8455e7 | !hbusreq0 & v8455ab;
assign v3a6f261 = hbusreq8_p & v3808d68 | !hbusreq8_p & v3740b8c;
assign v3809427 = hgrant3_p & v3a70710 | !hgrant3_p & v374bee4;
assign v3a6f896 = hbusreq6_p & v3a6fb7a | !hbusreq6_p & v37443ab;
assign v3731f9a = hmaster2_p & v3a70374 | !hmaster2_p & v3a70384;
assign v375b8cf = hmaster0_p & v3a6dcf5 | !hmaster0_p & v3764d26;
assign v3a6a73d = hgrant5_p & v3728876 | !hgrant5_p & v3741fe8;
assign v376d1b3 = hmaster2_p & v3a6f018 | !hmaster2_p & v377b576;
assign v372d0ad = hbusreq2_p & v37406d2 | !hbusreq2_p & v376648d;
assign v3a710b3 = hmaster1_p & a747d7 | !hmaster1_p & v3752798;
assign v3779d16 = hbusreq2_p & v3a6f975 | !hbusreq2_p & v8455ab;
assign v372dc2b = hgrant5_p & v373557e | !hgrant5_p & v3a6f6ca;
assign v3a7148c = hbusreq6_p & v3a6f87f | !hbusreq6_p & v374569b;
assign v37765e1 = hgrant3_p & v3747302 | !hgrant3_p & v2092ffc;
assign v374fa94 = hlock0_p & v3a67dd0 | !hlock0_p & v3775341;
assign v3778ac5 = hmaster2_p & v37482f8 | !hmaster2_p & v3a5f83e;
assign v3a6f3c6 = hbusreq6_p & v376e041 | !hbusreq6_p & v3748d67;
assign v3776c82 = hmaster0_p & v3a619a2 | !hmaster0_p & v3a5c3d3;
assign v3767cc0 = hmaster1_p & v3a6ef4e | !hmaster1_p & v8455ab;
assign v3748966 = hbusreq5 & v37631a9 | !hbusreq5 & v373bac6;
assign ade6f1 = hbusreq8_p & v372eec6 | !hbusreq8_p & v3a5902d;
assign v37311d6 = hgrant0_p & v3738c99 | !hgrant0_p & v8455ab;
assign v3a7004f = hmaster2_p & v3a6e5f0 | !hmaster2_p & v3a6f6a4;
assign v372775f = hbusreq8_p & v3a6f766 | !hbusreq8_p & v8455ab;
assign v376b5ad = hbusreq4 & v372a939 | !hbusreq4 & v3731230;
assign v37496fc = hmaster0_p & v8455ab | !hmaster0_p & v377b981;
assign v3760bb4 = stateG10_1_p & v3735ed0 | !stateG10_1_p & v3766035;
assign v3762cc4 = hlock3 & v3a6f588 | !hlock3 & v3a6ad8b;
assign v3a707e9 = hbusreq4 & v3a70893 | !hbusreq4 & v8455ab;
assign v3775393 = hbusreq5 & v376f182 | !hbusreq5 & v3a70d99;
assign v3760582 = stateG10_1_p & v39ebac7 | !stateG10_1_p & v3a70593;
assign d2728f = hbusreq4 & v38073b0 | !hbusreq4 & v8455ab;
assign v373d199 = hmaster0_p & v377700a | !hmaster0_p & v3a5a807;
assign v377c3a1 = hgrant3_p & v3a5a7c6 | !hgrant3_p & v3a6fe6a;
assign v3757727 = hgrant6_p & v3a5b5d3 | !hgrant6_p & !v3a6c835;
assign v3a64c14 = hmaster1_p & v372a0e3 | !hmaster1_p & v377e915;
assign v373db50 = hlock5_p & v3a6810b | !hlock5_p & !v3732510;
assign v37330ca = hbusreq5_p & v375c90c | !hbusreq5_p & v375aacf;
assign v3a6f52e = hgrant6_p & v3a6b873 | !hgrant6_p & v3777386;
assign v3757556 = hmaster0_p & v3a713f0 | !hmaster0_p & v3753a65;
assign v3733711 = hbusreq5 & v37742ca | !hbusreq5 & v8455ab;
assign v3a694b4 = hmaster0_p & v3a6f443 | !hmaster0_p & v37780fd;
assign v3a5ffbf = hbusreq6 & v3734af2 | !hbusreq6 & v8455ab;
assign v8455cd = hbusreq7_p & v8455ab | !hbusreq7_p & !v8455ab;
assign v3a5c00e = hlock6_p & v8455ab | !hlock6_p & v3761f22;
assign v3776413 = jx1_p & v8455ab | !jx1_p & v3741890;
assign v3a6fbc6 = jx0_p & v3a558ce | !jx0_p & v9c9282;
assign v3a5de59 = hlock7 & v3a6b57d | !hlock7 & v2092ee9;
assign v3a6edb1 = hgrant0_p & v3759b2f | !hgrant0_p & v8a7f7e;
assign v3a604bc = hbusreq0 & v373cd41 | !hbusreq0 & v3775252;
assign v3a70e52 = hbusreq1_p & v3a6eb45 | !hbusreq1_p & !v3a6eb81;
assign v3725bf4 = hbusreq6 & v3a673d6 | !hbusreq6 & v8455ab;
assign v3a5e1b7 = hlock7 & v373efdf | !hlock7 & v374457b;
assign v3a6b92c = hlock0 & v3a612a4 | !hlock0 & v3723d4b;
assign v3a6ba88 = hgrant5_p & v373f53e | !hgrant5_p & !v8455ab;
assign v372ebaa = hbusreq0_p & v3748797 | !hbusreq0_p & v3736e1d;
assign v3762453 = hgrant1_p & v3a5b5d3 | !hgrant1_p & v35772a6;
assign v3a704d0 = hlock2 & aebd68 | !hlock2 & v3751dc9;
assign v3a6f145 = hgrant6_p & v377f09a | !hgrant6_p & v374dafa;
assign v3740dc8 = hbusreq8_p & v3750ac3 | !hbusreq8_p & v3776eef;
assign v372d8e2 = hbusreq4 & v3a5b121 | !hbusreq4 & v377caa3;
assign v3a6f9a7 = hmaster0_p & v3757568 | !hmaster0_p & v374cd43;
assign v3a6bada = hlock6 & v373c377 | !hlock6 & v910050;
assign v375cc06 = hbusreq4 & v372d95c | !hbusreq4 & v3753dd4;
assign v37429cc = hmaster2_p & v3a6fe1a | !hmaster2_p & v8455b5;
assign v375dd60 = hlock2_p & v3770d6d | !hlock2_p & v37c02a0;
assign v377866b = hbusreq8_p & v3742dcb | !hbusreq8_p & v3747465;
assign v373d0af = hgrant3_p & v8455ab | !hgrant3_p & v3a70f64;
assign v376e5fe = hgrant6_p & v8455ab | !hgrant6_p & v37690ea;
assign v3a62fc4 = hbusreq4_p & v37704dc | !hbusreq4_p & v3757f01;
assign v3a70d7d = hbusreq7_p & v3730d77 | !hbusreq7_p & v375ed19;
assign v372e8ae = hgrant5_p & v374cd6b | !hgrant5_p & v3731476;
assign v3a6c43c = hmaster1_p & v373ad69 | !hmaster1_p & v37447b4;
assign v3730ad2 = hbusreq0 & v3a713ae | !hbusreq0 & v372eec5;
assign v3a63d0f = hmaster1_p & v8455ab | !hmaster1_p & v3777d6c;
assign v3a6fe27 = hmaster2_p & v374e51a | !hmaster2_p & !v8455ab;
assign v37770f5 = hmaster2_p & v376158d | !hmaster2_p & v8455ab;
assign v3a6a78c = hbusreq6 & v372f231 | !hbusreq6 & v8455ab;
assign v3a714f2 = hbusreq6_p & v376a4dd | !hbusreq6_p & v3a6b4a6;
assign v372459b = hbusreq8_p & v377a87d | !hbusreq8_p & v377601b;
assign v376495e = hlock0_p & v8455e7 | !hlock0_p & v3727eb2;
assign v373ae84 = hmaster1_p & v3756c2e | !hmaster1_p & v3a5fe51;
assign v3a5b109 = hlock5 & v3a63b7a | !hlock5 & v37229e0;
assign v37400fe = hmaster1_p & v38087c5 | !hmaster1_p & v3751e07;
assign v3739d49 = jx0_p & v377065f | !jx0_p & v374bd13;
assign v375d507 = hmaster2_p & v3758c65 | !hmaster2_p & v3a6f244;
assign ce4abb = hgrant4_p & v8455c1 | !hgrant4_p & v374e7e6;
assign v37549eb = hbusreq4 & v373d78b | !hbusreq4 & v8455ab;
assign v373bca5 = hlock8_p & v3756c19 | !hlock8_p & v3760ba7;
assign v3a64643 = hbusreq3_p & v3a55a19 | !hbusreq3_p & !v3a672c9;
assign v3731803 = hbusreq0 & v39ed7e6 | !hbusreq0 & v8455ab;
assign v375f159 = hmaster0_p & v3726e1f | !hmaster0_p & v3728fda;
assign v3772904 = hbusreq5_p & v3a5bf28 | !hbusreq5_p & v373ff04;
assign v377f264 = hbusreq5_p & v377e9b0 | !hbusreq5_p & v3a66856;
assign v3740f3d = hburst1 & v3757c6f | !hburst1 & v3a70b94;
assign v374195f = hbusreq4_p & v377445c | !hbusreq4_p & !v3777790;
assign b96080 = hlock0 & v3a6a934 | !hlock0 & v3747c90;
assign v3769c2e = hgrant2_p & v3771137 | !hgrant2_p & v374e6ec;
assign v373a496 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f8d1;
assign v372d2dc = hgrant4_p & v37747db | !hgrant4_p & v3736ea1;
assign v3760b03 = hbusreq5_p & v377dacb | !hbusreq5_p & v3a6f887;
assign v3772326 = hbusreq2 & v3a63abb | !hbusreq2 & v8455ab;
assign v3a61516 = hmaster0_p & v3a6f04d | !hmaster0_p & v8455ab;
assign v376d215 = hbusreq5_p & v375e30b | !hbusreq5_p & v3a66e6f;
assign v1e37405 = hmaster0_p & v3a70771 | !hmaster0_p & v3777536;
assign v373b8e2 = hbusreq0 & v3760854 | !hbusreq0 & v372c706;
assign v37575e7 = hbusreq2 & v39a5265 | !hbusreq2 & !v376f665;
assign v3a6f15c = hmaster2_p & v3730e7d | !hmaster2_p & v3a6f806;
assign v8cf677 = hmaster2_p & v3a701a1 | !hmaster2_p & v375ed6f;
assign v37463d4 = hmaster0_p & v376111d | !hmaster0_p & v376e562;
assign v373e87e = hlock7_p & v3730f5d | !hlock7_p & !v8455ab;
assign v37315fd = jx0_p & v8455ab | !jx0_p & v3724b94;
assign v3a708ce = hmaster2_p & v3a56531 | !hmaster2_p & v3766ff7;
assign v3a5d6b7 = hbusreq7_p & v37341ff | !hbusreq7_p & !v3751929;
assign v3a62c7d = hbusreq6_p & v372c713 | !hbusreq6_p & v377d714;
assign v3a6fb51 = hgrant6_p & v372ec1c | !hgrant6_p & v3726d2a;
assign v3a6900c = hbusreq0_p & v8455ab | !hbusreq0_p & v8455b0;
assign v372ab6c = hmaster0_p & v3742725 | !hmaster0_p & v37662e7;
assign d52046 = hgrant5_p & v3755082 | !hgrant5_p & v3a70276;
assign v377c3ad = hlock0 & v373bd6c | !hlock0 & v3a70c55;
assign v1e37a8d = hbusreq5 & v3726ee7 | !hbusreq5 & v8455ab;
assign v360d016 = hgrant1_p & v8455ab | !hgrant1_p & !v3761785;
assign v374f82e = hgrant4_p & v8455ab | !hgrant4_p & v3758d7e;
assign v88e7d1 = hbusreq5 & v3778619 | !hbusreq5 & v3a711e6;
assign v377d06b = hmaster0_p & v3a6f833 | !hmaster0_p & v374953c;
assign v373e4db = hlock4 & v375e815 | !hlock4 & v37413d8;
assign v3735760 = hbusreq5 & v373809d | !hbusreq5 & v376784b;
assign v3a6d434 = hlock8 & v3a5d55b | !hlock8 & v3a70cac;
assign v1e37ab9 = hlock3_p & v3a622d0 | !hlock3_p & v37658b1;
assign v377814b = hbusreq2 & v3a70cea | !hbusreq2 & v8455ab;
assign v3779b96 = hgrant7_p & v3a6f2d5 | !hgrant7_p & v3756bd2;
assign v372ec6d = hgrant4_p & v376428f | !hgrant4_p & dac328;
assign v3762924 = hbusreq4_p & v373ec24 | !hbusreq4_p & !v3a56cdb;
assign v3742275 = hmaster0_p & v3a66c66 | !hmaster0_p & v374eaf4;
assign v3762870 = hgrant4_p & v3759b2f | !hgrant4_p & v3a6a442;
assign v3738a87 = hmaster0_p & v3a70ca8 | !hmaster0_p & v8455e7;
assign v3a5b87f = hmaster2_p & v3a635ea | !hmaster2_p & v373cf9c;
assign v3a6ffc1 = hlock5 & v3a6d792 | !hlock5 & v3a70c33;
assign v3731f07 = hgrant8_p & v8455ab | !hgrant8_p & v377815d;
assign v3a705d1 = hmaster0_p & v374faf5 | !hmaster0_p & v3a7026a;
assign v380952f = hmaster2_p & v3a70f5e | !hmaster2_p & !v374ab8d;
assign v375070a = hbusreq8 & a5c257 | !hbusreq8 & v376d66c;
assign a8c5c5 = hbusreq4_p & v325c960 | !hbusreq4_p & v3752446;
assign v23fe27f = hlock4 & v3777daa | !hlock4 & cff2df;
assign v373c331 = hgrant0_p & c51df8 | !hgrant0_p & v3a6f562;
assign v3a57bb0 = hbusreq6 & v3775750 | !hbusreq6 & v35b774b;
assign v3738ed8 = hmaster2_p & v373a822 | !hmaster2_p & v37788a6;
assign v3a6145f = hgrant3_p & v3739018 | !hgrant3_p & !v3771bed;
assign v3a70abc = hlock6_p & v3a6f880 | !hlock6_p & v8455ab;
assign v3a60fa7 = hgrant5_p & v3728992 | !hgrant5_p & v3378996;
assign v377ed25 = hmaster0_p & v3a5b6ac | !hmaster0_p & v374549a;
assign v3761a8f = hmaster0_p & v372b6d0 | !hmaster0_p & v376a6f1;
assign v3a6f9e8 = hgrant4_p & v8455ab | !hgrant4_p & v3725dce;
assign v37473a3 = hgrant6_p & v375f653 | !hgrant6_p & v3776f7f;
assign v3a59ce1 = hbusreq5_p & v3727bc1 | !hbusreq5_p & v3a2a107;
assign v35b7153 = hbusreq5 & v3a60f21 | !hbusreq5 & v3a2a107;
assign v3728bc3 = hmaster1_p & v3779183 | !hmaster1_p & v375705a;
assign v3764d9e = hgrant2_p & v3757c37 | !hgrant2_p & v3745a47;
assign v2092baa = hbusreq6_p & v373f492 | !hbusreq6_p & v372f16b;
assign v373313b = hbusreq6_p & v3a5bd48 | !hbusreq6_p & v3a6bc78;
assign v374b5a8 = hbusreq4_p & v3a6fd81 | !hbusreq4_p & v3a702c2;
assign v3a70cfa = hmaster1_p & v3a6eecb | !hmaster1_p & v37420de;
assign v375964f = hbusreq2_p & v37291d1 | !hbusreq2_p & v372e27f;
assign v374999b = hbusreq4 & v3723ace | !hbusreq4 & v3722e7a;
assign v3a6bef4 = hmaster2_p & v8455ab | !hmaster2_p & v3a6a580;
assign v375f486 = hbusreq4_p & v3722b92 | !hbusreq4_p & !v8455ab;
assign v3a69444 = hgrant4_p & v3a592be | !hgrant4_p & v3763d52;
assign v377affd = hgrant3_p & v3a6c2b6 | !hgrant3_p & !v3767904;
assign v380a0c2 = hbusreq6_p & v37583be | !hbusreq6_p & v3a5be20;
assign v3751a86 = hlock0 & v375da10 | !hlock0 & v3729785;
assign v3755c0e = hlock5_p & v3a6b5ba | !hlock5_p & !v3a6ff71;
assign v372b8eb = hbusreq4_p & v374853c | !hbusreq4_p & v3748d67;
assign v3779e45 = hbusreq2_p & v3748d3e | !hbusreq2_p & !v8455ab;
assign v377b6fc = hbusreq6 & v380663a | !hbusreq6 & !v3727e59;
assign v3757765 = hbusreq0 & v376f56d | !hbusreq0 & v8455ab;
assign v3a709d3 = hlock5_p & v3748990 | !hlock5_p & !v376faf6;
assign v3a6fc5e = hgrant4_p & v8455c2 | !hgrant4_p & v377b4cc;
assign v3732bff = hmaster2_p & v3a635ea | !hmaster2_p & v3a6f71a;
assign v3a710ad = hlock6 & v3759536 | !hlock6 & v3a7116e;
assign v37477dd = hbusreq2 & v3744cea | !hbusreq2 & v3a6fdef;
assign v375b5ce = hmaster2_p & v23fe0be | !hmaster2_p & v3736ded;
assign v3a5d989 = hbusreq5_p & v3761719 | !hbusreq5_p & v3731b41;
assign v3774bc0 = hgrant5_p & v3a5ff7c | !hgrant5_p & v372d378;
assign v3769041 = hbusreq3_p & v37482be | !hbusreq3_p & v3a640c5;
assign v374bb74 = jx0_p & v3756723 | !jx0_p & v8455ab;
assign v3a701a2 = hgrant4_p & v3766e55 | !hgrant4_p & v372e25b;
assign v3a540f8 = hmaster0_p & v3a6a56e | !hmaster0_p & v37390c9;
assign v3a71121 = hbusreq2_p & v3734967 | !hbusreq2_p & !v374729b;
assign v3735293 = hgrant6_p & v376a040 | !hgrant6_p & !v375135a;
assign v3761351 = hgrant5_p & v3757f6d | !hgrant5_p & v3770bca;
assign v37555fd = hlock5_p & v3a70c8e | !hlock5_p & !v8455ab;
assign v3a6f717 = hgrant2_p & v8455b5 | !hgrant2_p & v3a69f36;
assign v3a6613e = hgrant3_p & dab321 | !hgrant3_p & !v375bc6e;
assign v374abb5 = hmaster1_p & v37245f8 | !hmaster1_p & v3723ee4;
assign v3753c8c = hmaster1_p & v372580e | !hmaster1_p & v374c69c;
assign v3a58e93 = hmaster2_p & v3a70e2e | !hmaster2_p & v3735b3e;
assign v3a5c904 = hgrant0_p & v3722eaf | !hgrant0_p & !v3a664b8;
assign v375e91e = hbusreq7_p & v3727699 | !hbusreq7_p & v376ca61;
assign v3a6841c = hmastlock_p & v376b164 | !hmastlock_p & v8455ab;
assign v3722b42 = hbusreq3 & v3a617b4 | !hbusreq3 & v3773ee6;
assign v3806ff0 = hbusreq2 & v374fd4a | !hbusreq2 & v3a5b2fd;
assign v3a667d2 = hbusreq7_p & v3746a45 | !hbusreq7_p & v3a6d8a9;
assign ab11fe = hbusreq5 & v3258dd9 | !hbusreq5 & v3771c85;
assign v3a70c0b = hbusreq2_p & v3733887 | !hbusreq2_p & v373ad95;
assign v374140e = hgrant8_p & v372d86d | !hgrant8_p & v3770dbf;
assign v377b2d0 = hgrant6_p & v8455ab | !hgrant6_p & v376cd14;
assign v37764c0 = hgrant4_p & v8455ab | !hgrant4_p & v3777abf;
assign v2ff9287 = hbusreq3_p & v3752ec0 | !hbusreq3_p & v8455e9;
assign v3747926 = hmaster0_p & v3a6b100 | !hmaster0_p & v37429c2;
assign v377bf0d = hbusreq0_p & v3a6f316 | !hbusreq0_p & v3738f04;
assign v3a5b45b = hmaster0_p & v37312e3 | !hmaster0_p & v3a70f68;
assign v3745714 = hmaster2_p & v1e38224 | !hmaster2_p & !v37521ed;
assign v3734c60 = hbusreq1_p & v38071c1 | !hbusreq1_p & !v3748d8c;
assign v3a70d78 = hbusreq7 & v3a6f55d | !hbusreq7 & v3733173;
assign v377ad76 = hbusreq0 & v3a56cca | !hbusreq0 & v375a635;
assign v3a55fc1 = jx1_p & v3a7049d | !jx1_p & v375745a;
assign v3723749 = hmaster1_p & v3a700d9 | !hmaster1_p & v3736ea9;
assign v3765109 = hmaster2_p & v3723af9 | !hmaster2_p & v3a6ac60;
assign v374b10b = hgrant4_p & v8455e1 | !hgrant4_p & !v377762d;
assign v3a71025 = hbusreq0 & v3775831 | !hbusreq0 & v3a70417;
assign v3748ff3 = hmaster0_p & v3749649 | !hmaster0_p & v2092ec6;
assign v3733da4 = hbusreq0 & v373d8ec | !hbusreq0 & v3774e32;
assign v3a68728 = hbusreq0 & v3749e96 | !hbusreq0 & v376beed;
assign v3746aa9 = hlock7 & v3a615c7 | !hlock7 & v3a5bed2;
assign v373fdae = hmaster2_p & v374bfd2 | !hmaster2_p & v37745c3;
assign v3806fa6 = hgrant3_p & v3a6f627 | !hgrant3_p & v37258c9;
assign v376beee = stateA1_p & v376a35c | !stateA1_p & !v8455e1;
assign v3a70799 = hgrant3_p & v3a5e1a5 | !hgrant3_p & v377af98;
assign v373f17f = hbusreq4_p & v37fca8d | !hbusreq4_p & v3a704ea;
assign v3a6ff07 = hmaster1_p & v3a5aaca | !hmaster1_p & v209300b;
assign v3773250 = hbusreq2 & v39a5265 | !hbusreq2 & !v2aca977;
assign v3a603f3 = hbusreq5_p & v3a700ea | !hbusreq5_p & v3a7055a;
assign v373471f = hbusreq4 & v2925d19 | !hbusreq4 & v3749bf0;
assign v373dcb6 = hgrant1_p & v375cd0c | !hgrant1_p & v8455ab;
assign v377c44f = hgrant4_p & v3a6b873 | !hgrant4_p & v3a6f52e;
assign v3766e8b = hlock2 & v3a6a4cf | !hlock2 & v373d0af;
assign v3a5ec6b = hgrant5_p & v372bbab | !hgrant5_p & v3a5dc2a;
assign v3748446 = hmaster0_p & v8455b0 | !hmaster0_p & v3a70641;
assign v3745e51 = hmaster0_p & v3808e85 | !hmaster0_p & v376981e;
assign v375c99d = hbusreq8 & v377929d | !hbusreq8 & v376b504;
assign v3a6f89d = hbusreq6 & v3a6fe0d | !hbusreq6 & !v8455b5;
assign v3757575 = hlock4_p & v3756fba | !hlock4_p & v3a5b213;
assign v360cffa = hlock8_p & v373ec92 | !hlock8_p & v8455b7;
assign v372a9a5 = hbusreq5 & v3740d05 | !hbusreq5 & v3a71530;
assign v377d95a = hmaster2_p & v373b87c | !hmaster2_p & v3756cee;
assign v3a6ff39 = hlock5_p & v375bb26 | !hlock5_p & v3738f35;
assign v3a70e9b = hgrant6_p & v3761fb5 | !hgrant6_p & v3a59df2;
assign v377e328 = hmaster0_p & v3a64421 | !hmaster0_p & v3a70f66;
assign v3a714f8 = hbusreq8 & v3a67c6d | !hbusreq8 & v8455ab;
assign v3a6fa22 = hmaster2_p & v2ff9314 | !hmaster2_p & v3759379;
assign v377aa17 = hbusreq6 & v3a70200 | !hbusreq6 & !cfe6df;
assign v3a67c34 = hbusreq7 & v3a6f20c | !hbusreq7 & v3a71082;
assign v3a6f2c9 = hmaster2_p & v8455ab | !hmaster2_p & v3733b37;
assign hmaster1 = !v190eb62;
assign v3a640e3 = hlock5 & v37287d2 | !hlock5 & v373666f;
assign v3753278 = hbusreq8 & v3a708a6 | !hbusreq8 & v3774452;
assign v3735f7a = hgrant2_p & v8455b9 | !hgrant2_p & v3809f5f;
assign v376ef46 = hgrant6_p & v8455ab | !hgrant6_p & v372d7ed;
assign v905dc4 = hbusreq8_p & v3743dff | !hbusreq8_p & v3a5f853;
assign v3729a1c = hbusreq6_p & v3734c20 | !hbusreq6_p & v3a641d5;
assign v3a6f072 = hbusreq5_p & v37c01ec | !hbusreq5_p & v374c9ab;
assign v3728685 = hgrant4_p & v3759886 | !hgrant4_p & !v8455ab;
assign v38071c7 = hbusreq7_p & v3a712d2 | !hbusreq7_p & v3a664ed;
assign v3a66ada = hgrant4_p & v3a6d48c | !hgrant4_p & v3774a12;
assign v3a6eb7e = hmaster2_p & v3a6fcb0 | !hmaster2_p & v377988b;
assign v3a6eb4b = hmaster1_p & v3728a3d | !hmaster1_p & v3a6f937;
assign v376bb64 = hgrant0_p & v8455ab | !hgrant0_p & v3755e29;
assign v37559ea = hbusreq6 & v374956a | !hbusreq6 & v3a635ea;
assign v3a6ded8 = hbusreq7 & v3748efb | !hbusreq7 & a18d54;
assign d648e4 = hbusreq0 & v377873a | !hbusreq0 & v376c490;
assign v3728963 = hbusreq0 & v3a6f477 | !hbusreq0 & v3a714cc;
assign v3a6a82d = hbusreq7_p & v3778e98 | !hbusreq7_p & v3a61375;
assign v3772e3f = hmaster1_p & v8455ab | !hmaster1_p & !v3778b83;
assign v3776d62 = hgrant5_p & v3a58604 | !hgrant5_p & v373c074;
assign v3a70453 = hmaster2_p & v3a6e57f | !hmaster2_p & v3728d9c;
assign v3768c08 = hmaster0_p & v3a66d94 | !hmaster0_p & v372e213;
assign v3a6c0fb = hbusreq6_p & v376eb1f | !hbusreq6_p & v8455ab;
assign v3766438 = hbusreq0_p & v2ff9190 | !hbusreq0_p & v3a6da9c;
assign v375973d = hgrant5_p & v3736ae6 | !hgrant5_p & v3726d4a;
assign v37296f0 = hgrant0_p & v3a69e18 | !hgrant0_p & v375803a;
assign v3a5a73d = hbusreq6_p & v372904d | !hbusreq6_p & v373650c;
assign v375a938 = hlock4_p & v373aed4 | !hlock4_p & v8455bf;
assign v3a6d9da = hmaster0_p & v373cedd | !hmaster0_p & !v3a658cf;
assign v3a6fb69 = hbusreq5 & v3a69fde | !hbusreq5 & v375d417;
assign v376de00 = hbusreq5 & v37555fd | !hbusreq5 & v372c6ce;
assign v3a710f6 = hgrant6_p & v377f09a | !hgrant6_p & !v3a6fb7c;
assign v3a647cd = hbusreq8_p & v3a6f569 | !hbusreq8_p & b5394c;
assign c8bdc6 = jx1_p & v373627b | !jx1_p & v3a6efc3;
assign v37572f7 = hlock6 & v375d4d9 | !hlock6 & v37526d6;
assign v3736eff = hmaster2_p & v3a635ea | !hmaster2_p & v3a63621;
assign v3a63033 = hmaster2_p & v375e75d | !hmaster2_p & v3a66822;
assign v3a70524 = hbusreq3_p & v37777d2 | !hbusreq3_p & v8455ab;
assign v3758c72 = hmaster2_p & v3a6ebed | !hmaster2_p & v377eb45;
assign v3772a87 = hlock3 & v3769616 | !hlock3 & v372d880;
assign b0b0c6 = hbusreq7_p & v3a693ca | !hbusreq7_p & v374d41e;
assign v373b4e6 = hbusreq4 & v3759970 | !hbusreq4 & v373f647;
assign v3722a0a = hgrant2_p & v372f09a | !hgrant2_p & v3a654c4;
assign v3255a0f = hbusreq7_p & v375f848 | !hbusreq7_p & v373c7af;
assign v3a711e8 = hgrant4_p & v376a6f1 | !hgrant4_p & v3726810;
assign v3728b2f = hbusreq3_p & v37401f0 | !hbusreq3_p & v374ea45;
assign v37434bc = hbusreq7_p & v3a6ef27 | !hbusreq7_p & v372dd94;
assign v372760c = hbusreq7_p & v376ad33 | !hbusreq7_p & v376ce17;
assign v3a6fc2b = hmaster2_p & v3a6dfb2 | !hmaster2_p & !v372935c;
assign v3a6360c = hlock8 & v3a61388 | !hlock8 & v3a637fd;
assign v3a714c3 = hlock0_p & v8455ab | !hlock0_p & v376915a;
assign v3a6ffea = hbusreq4_p & v3a6f92f | !hbusreq4_p & !v377adf5;
assign v372ce45 = hlock0 & v3a70c74 | !hlock0 & v3a70ed9;
assign v3a66773 = hbusreq6 & v3a7025f | !hbusreq6 & v375b9c1;
assign v3a70968 = hgrant7_p & v3a649c2 | !hgrant7_p & v376f2f4;
assign v3a6fe74 = hbusreq4_p & v3731803 | !hbusreq4_p & v37785be;
assign v360d147 = hlock4_p & v375ec98 | !hlock4_p & v375c845;
assign v3757e15 = hmaster1_p & v372d891 | !hmaster1_p & v3735bbc;
assign v3a55aa3 = hmaster0_p & v8455e7 | !hmaster0_p & v37788d5;
assign v3750559 = hbusreq8 & v3753404 | !hbusreq8 & v3737808;
assign v377f76a = hbusreq3_p & v3a71528 | !hbusreq3_p & !v3a71065;
assign v37358ab = hbusreq4_p & v8455c2 | !hbusreq4_p & !v8455ab;
assign v372e885 = hmaster0_p & v372ef36 | !hmaster0_p & v37341d3;
assign v3a6fa57 = hlock8_p & v3767a2f | !hlock8_p & v3746a45;
assign v3743434 = hbusreq0 & v372ab46 | !hbusreq0 & !v8455ab;
assign v3779810 = hmaster1_p & v8455ab | !hmaster1_p & v374dabe;
assign v372cd61 = hmaster0_p & v3a6f7ee | !hmaster0_p & v3a70bf3;
assign v3725eb6 = hbusreq8_p & v37585c9 | !hbusreq8_p & b0ac65;
assign v3764e95 = hgrant2_p & v372abd8 | !hgrant2_p & v374fb93;
assign v3a70593 = hgrant1_p & v376d45f | !hgrant1_p & v3a70c07;
assign v1e37721 = hlock6 & v376ee03 | !hlock6 & v3a644e6;
assign v3a70119 = hbusreq5 & v3a71375 | !hbusreq5 & v3770aee;
assign v3742b54 = hbusreq0 & v3a710cb | !hbusreq0 & !v37298b9;
assign v377c546 = hgrant3_p & v3a6ffb6 | !hgrant3_p & d39337;
assign v3a587f6 = hbusreq0 & v3733412 | !hbusreq0 & v372cc25;
assign v1e3786e = hgrant4_p & v8455ab | !hgrant4_p & v947c98;
assign v375b0f9 = hbusreq7_p & v8455cf | !hbusreq7_p & !v8455ab;
assign v3777888 = hbusreq5 & v3774385 | !hbusreq5 & v3a70582;
assign v373a09f = hmaster0_p & v3a635ea | !hmaster0_p & v3a57f6c;
assign v3a6fb1b = hbusreq5 & v37553b9 | !hbusreq5 & v8455bb;
assign v3a656dd = hmaster1_p & v3a6e5f0 | !hmaster1_p & v37576b1;
assign v373d9b3 = hmaster2_p & v373eaf6 | !hmaster2_p & v372c257;
assign v37283fe = hgrant4_p & v8455ab | !hgrant4_p & v372fb48;
assign v3764378 = hbusreq7 & v3774b71 | !hbusreq7 & v3a5fb90;
assign v380719b = hgrant6_p & v3a6f3a1 | !hgrant6_p & v3a6fe94;
assign v376eb2b = hgrant1_p & v3a6e591 | !hgrant1_p & v3a6f252;
assign v3a70dd9 = hmaster2_p & v3a704cc | !hmaster2_p & v3750a9c;
assign v3a5b7ad = hlock5 & v3744c08 | !hlock5 & v376aae5;
assign v8f9a63 = hmaster1_p & v3a63ea7 | !hmaster1_p & v372e332;
assign v3760646 = hbusreq5_p & v377de7f | !hbusreq5_p & v3764caa;
assign v3a70b2c = hbusreq6 & v3765e46 | !hbusreq6 & v8455ab;
assign v2678c40 = hbusreq1_p & v3758c64 | !hbusreq1_p & !v376db07;
assign v37243fe = hmaster2_p & v3a5ee73 | !hmaster2_p & v3774c1b;
assign v3a60f9b = hbusreq5 & bf6c15 | !hbusreq5 & v8455ab;
assign v3a62122 = hgrant3_p & v3a6c2b6 | !hgrant3_p & !v37440ff;
assign v3808865 = hmaster0_p & v37430fb | !hmaster0_p & v3750edc;
assign v372d02d = hbusreq3_p & v3726f6c | !hbusreq3_p & !v3a6ff7d;
assign v373bafb = jx1_p & v3a5cd0e | !jx1_p & v3740aa8;
assign v3752ef1 = hgrant1_p & v372fc81 | !hgrant1_p & v8455ab;
assign adaeff = hmaster3_p & v3a69203 | !hmaster3_p & v375b84e;
assign v37723c6 = hbusreq7 & v38098b0 | !hbusreq7 & v3a666a9;
assign v37619b8 = hgrant0_p & v3726806 | !hgrant0_p & v23fe285;
assign v372721d = hgrant5_p & v8455c6 | !hgrant5_p & v37289f0;
assign v3765e6a = hgrant6_p & v3a6984f | !hgrant6_p & v3727ff7;
assign v3a61d83 = hlock4_p & v376a14f | !hlock4_p & v8455e7;
assign v376daf6 = hbusreq2_p & v37765e1 | !hbusreq2_p & v380917f;
assign v3a70b5d = hlock2 & v3759ffd | !hlock2 & v375767e;
assign v3765f8e = hmaster1_p & v3727fa7 | !hmaster1_p & v3a61ff9;
assign v3a70057 = hgrant2_p & v376b5f8 | !hgrant2_p & v3762934;
assign v3a57741 = hmaster2_p & v373096c | !hmaster2_p & v3742e6b;
assign v37666d7 = hbusreq7_p & v3745e54 | !hbusreq7_p & v374a7f2;
assign v3a6f518 = hbusreq7 & v3a6fd9c | !hbusreq7 & v3a6f435;
assign v3772bb3 = hmaster0_p & v3a661fe | !hmaster0_p & v377a615;
assign v3752edc = hmaster1_p & v374a1f5 | !hmaster1_p & v3739589;
assign v3a6ff99 = hbusreq0 & v375cb14 | !hbusreq0 & v3807a2e;
assign v372d33c = hbusreq7_p & v3a67a02 | !hbusreq7_p & v3a698d8;
assign v372fe64 = hbusreq8_p & v3a57796 | !hbusreq8_p & !v8455ab;
assign v37391b4 = hgrant2_p & v377db21 | !hgrant2_p & v3806b87;
assign v374d162 = hmaster1_p & v377d76b | !hmaster1_p & v3a5a8a4;
assign v373d8c3 = hbusreq5 & v3a71002 | !hbusreq5 & v3767a21;
assign v3a714fc = hbusreq4 & v373935b | !hbusreq4 & v376e513;
assign v3733ae1 = hbusreq0 & v3a6f326 | !hbusreq0 & v3a67e53;
assign v37319c5 = hlock5 & v3757537 | !hlock5 & v3a53ed2;
assign v372ca24 = hlock5_p & v376b2ab | !hlock5_p & v3a7045d;
assign v3a605af = hbusreq4 & v374c3d0 | !hbusreq4 & v373031f;
assign v3731b28 = hbusreq5 & v377aed1 | !hbusreq5 & v375e512;
assign v3743df6 = hbusreq8 & v3a6d2e2 | !hbusreq8 & v372d827;
assign v37512a0 = hbusreq2_p & v374125a | !hbusreq2_p & v3a6eeca;
assign v3a5fa82 = hmaster0_p & v3a60c4f | !hmaster0_p & v37429c2;
assign v3a60a75 = hbusreq0 & v372807c | !hbusreq0 & v3745366;
assign v3a69f9e = hbusreq6_p & v3a70cf0 | !hbusreq6_p & v375e00a;
assign v377ccba = hbusreq4_p & v3a7094d | !hbusreq4_p & v3a66750;
assign v374fd32 = hbusreq5 & v3a69b77 | !hbusreq5 & v37358ab;
assign v3a6b6d2 = hbusreq2 & v3a619c0 | !hbusreq2 & !v8455ab;
assign v376b03d = hmaster0_p & v3577306 | !hmaster0_p & v380886b;
assign v377e871 = hgrant5_p & v8455ab | !hgrant5_p & !v37536b8;
assign v3733234 = hgrant2_p & v377b6ce | !hgrant2_p & v374262d;
assign v3a71308 = hgrant4_p & v372298c | !hgrant4_p & v3809112;
assign v3a6b51f = hbusreq0 & v3a66c6c | !hbusreq0 & v3766d5a;
assign v3757b0f = hmaster1_p & v37519a8 | !hmaster1_p & v375d78f;
assign v3729988 = hbusreq5_p & v37280a3 | !hbusreq5_p & v37719a0;
assign v37753b4 = hmaster0_p & v3a70630 | !hmaster0_p & v3809d9e;
assign v20930c9 = hmaster2_p & v3a637dd | !hmaster2_p & !v37346be;
assign hgrant8 = v3a28da6;
assign v3736104 = hmaster2_p & v3759032 | !hmaster2_p & v37432c6;
assign v373df0d = hbusreq2_p & v3750b04 | !hbusreq2_p & v35772a6;
assign v3777d95 = hbusreq6 & v1e38224 | !hbusreq6 & v8455ab;
assign v3725cc8 = hlock4 & v37233d2 | !hlock4 & v3a6db1a;
assign v3a60bee = hmaster0_p & v8455ab | !hmaster0_p & v3738321;
assign v374cf68 = jx0_p & v3778e46 | !jx0_p & v3a70a21;
assign v374871a = hlock5 & v3a656be | !hlock5 & v3a5a5a7;
assign v373a327 = hmaster0_p & v3761947 | !hmaster0_p & v8455ab;
assign v376a04d = hmaster0_p & v3748fde | !hmaster0_p & v3768495;
assign v3778998 = hmaster0_p & v3a67d66 | !hmaster0_p & v3776f42;
assign v3a70a81 = hbusreq0 & v3a6b62d | !hbusreq0 & v3a70d32;
assign v3a6eb0e = hmaster0_p & v3755002 | !hmaster0_p & v23fd858;
assign v3732511 = hmaster1_p & v3725198 | !hmaster1_p & v3762969;
assign v3a5b89b = hbusreq6_p & v372493b | !hbusreq6_p & !v3a6febd;
assign v3775f27 = hmaster2_p & v373c4c2 | !hmaster2_p & v37302f1;
assign v37390ce = hbusreq0 & v377831d | !hbusreq0 & v8455ab;
assign v372baaf = hbusreq4 & v373f42f | !hbusreq4 & v8455ab;
assign v3768e31 = hbusreq8_p & v375c724 | !hbusreq8_p & v373df91;
assign v3729c71 = hgrant7_p & v37530cf | !hgrant7_p & v3a5858c;
assign v3779477 = hmaster0_p & v376589f | !hmaster0_p & v3757ffa;
assign v37664e7 = hbusreq4 & v37266cb | !hbusreq4 & v3725799;
assign v3774bad = hbusreq4_p & v8455c3 | !hbusreq4_p & !v8455ab;
assign v3a6a8c5 = hgrant0_p & v8455ab | !hgrant0_p & v8455eb;
assign v375c8c4 = hmaster2_p & v8455ab | !hmaster2_p & v374f87c;
assign v3a6f929 = hlock5_p & v3a619c0 | !hlock5_p & !v8455ab;
assign v380755c = hmaster1_p & v372e443 | !hmaster1_p & v3a6eb7a;
assign v3769f95 = hlock3_p & v3767885 | !hlock3_p & v37488ed;
assign v3750775 = hbusreq2 & v3a69bf4 | !hbusreq2 & v8455bf;
assign v377f3ae = hbusreq5 & v373b16f | !hbusreq5 & v8455ab;
assign v374bda9 = hgrant6_p & v8455ab | !hgrant6_p & v3a6f457;
assign v37548e9 = hbusreq5 & v3a5c4c6 | !hbusreq5 & v37494c3;
assign v376efdb = hgrant2_p & v8455ab | !hgrant2_p & v3a70f01;
assign v374b923 = hbusreq6_p & v3744640 | !hbusreq6_p & v8455ab;
assign abddc4 = hbusreq4 & v373f954 | !hbusreq4 & v8455ab;
assign v3a6f505 = hbusreq0 & v3a70f67 | !hbusreq0 & v376c5f5;
assign v3725152 = hbusreq6 & v3a660f2 | !hbusreq6 & v8455ab;
assign v37513d1 = hgrant1_p & v373c4e4 | !hgrant1_p & v3740171;
assign v376b4ad = hbusreq6_p & v376a015 | !hbusreq6_p & v8455ab;
assign v3764c0d = hmaster0_p & v377027e | !hmaster0_p & !v3777f6e;
assign v3a5bc04 = hbusreq0 & v3a70966 | !hbusreq0 & v3a68822;
assign v3a6faf0 = hlock7 & v372a0cb | !hlock7 & v3a70f38;
assign v375a7fc = hbusreq0_p & v3723ac5 | !hbusreq0_p & v8455ab;
assign v3808cbf = hmaster1_p & v3748e5a | !hmaster1_p & v372ee5a;
assign v376b036 = hmaster0_p & v3a70029 | !hmaster0_p & v3a6fd53;
assign v3775b3a = hbusreq5 & v3a6f76a | !hbusreq5 & v8455ab;
assign v374e109 = hmaster0_p & v8455ab | !hmaster0_p & v3741dea;
assign v373aed4 = hbusreq3_p & v376d955 | !hbusreq3_p & v8455ab;
assign v375bc70 = hmaster0_p & v37782c9 | !hmaster0_p & v3757888;
assign v3a6fc94 = hmaster1_p & v3a6b27d | !hmaster1_p & v374e7fa;
assign v3a709ae = hbusreq5 & v3a6faff | !hbusreq5 & v375cbcb;
assign v3a70e86 = hbusreq3_p & v3a6a8d2 | !hbusreq3_p & v8455b0;
assign v37514f7 = hbusreq5_p & v373e12b | !hbusreq5_p & !v37682ce;
assign v37317da = hbusreq5_p & v3726eea | !hbusreq5_p & c7ae7d;
assign v3731164 = hmaster2_p & v375dcd5 | !hmaster2_p & v3a5bb42;
assign v3a70170 = hbusreq7_p & v3a638f4 | !hbusreq7_p & v3a5aa93;
assign v3809879 = hgrant6_p & v375d861 | !hgrant6_p & v373f028;
assign v3727de3 = hmaster3_p & v3724579 | !hmaster3_p & v377435f;
assign v373d071 = hmaster1_p & v377accc | !hmaster1_p & v3738666;
assign v3a6756b = jx1_p & v8455ab | !jx1_p & v9a641e;
assign v3a6f227 = hbusreq7_p & v3a63cf5 | !hbusreq7_p & c8ca6f;
assign v377455b = jx1_p & v375e29c | !jx1_p & v374fa2a;
assign v377d146 = hmaster1_p & v3a547ff | !hmaster1_p & v374925f;
assign v373feaa = hbusreq4_p & v375f169 | !hbusreq4_p & !v3749bba;
assign v3767420 = hgrant2_p & v3722e5c | !hgrant2_p & v3738d68;
assign v3a620ef = hgrant4_p & v8455ab | !hgrant4_p & v3a70255;
assign v3760a6e = hbusreq7 & v3768ed2 | !hbusreq7 & !v8455b5;
assign v3758a23 = hbusreq5 & v8455ab | !hbusreq5 & v3a59a2b;
assign v377682d = hlock0_p & v373aecf | !hlock0_p & !v3724026;
assign v3806f08 = hlock0 & v3a641d5 | !hlock0 & v3769e70;
assign v948ef2 = hmaster2_p & v3a62bae | !hmaster2_p & v37449fc;
assign v2acb068 = hbusreq5 & v373dd5a | !hbusreq5 & v372c85e;
assign v3a7126e = hmaster0_p & v37712aa | !hmaster0_p & v3a6567f;
assign v3730019 = hmaster1_p & v3734f6d | !hmaster1_p & v3a69949;
assign v3749d86 = hmaster2_p & v3a59c65 | !hmaster2_p & v377f2a9;
assign v373664d = hbusreq5_p & v3765463 | !hbusreq5_p & v3738a59;
assign v375be90 = hlock7 & v375554d | !hlock7 & v3739621;
assign v375be11 = hmaster1_p & v374c34d | !hmaster1_p & b736f4;
assign v372cfd5 = hlock4 & v376c30a | !hlock4 & v3a703bb;
assign v373e3d5 = hbusreq6 & v372d7a4 | !hbusreq6 & v372e83f;
assign v39eb519 = hbusreq5_p & v376de5c | !hbusreq5_p & v3a7088b;
assign v3a5bab6 = hlock6_p & v376a8d5 | !hlock6_p & !v8455ab;
assign v3726bb8 = hlock0_p & v375323b | !hlock0_p & v8455ab;
assign v3731dfd = hbusreq4_p & v376ce77 | !hbusreq4_p & v3a5fc34;
assign v37277c3 = hbusreq3_p & v37289ee | !hbusreq3_p & v3770f51;
assign v374bbc7 = hbusreq4_p & v3a5cebb | !hbusreq4_p & v377c6cf;
assign v3a70746 = hmaster1_p & v3725a2e | !hmaster1_p & v3a70144;
assign v37512ca = hbusreq4_p & v374f35a | !hbusreq4_p & v3a68d2e;
assign v376d66c = hmaster1_p & v3a6c4e4 | !hmaster1_p & v3a700ea;
assign v3a5a397 = hbusreq6 & v3a7162e | !hbusreq6 & v376005f;
assign v3749408 = hbusreq3_p & v3757388 | !hbusreq3_p & v8455ab;
assign v374d479 = hbusreq3_p & v8455b7 | !hbusreq3_p & v3732302;
assign v374a66c = hmaster1_p & v3770b73 | !hmaster1_p & v377af60;
assign v3756a09 = hbusreq0_p & v37376c8 | !hbusreq0_p & v377c3fb;
assign v3a70236 = hbusreq5_p & v3763f8e | !hbusreq5_p & v374c9ab;
assign v3a2a128 = hmaster3_p & v8455ab | !hmaster3_p & !v372dc34;
assign v3a6fe96 = hgrant4_p & v374ad16 | !hgrant4_p & v375b64b;
assign v37470eb = hbusreq1 & v39a5381 | !hbusreq1 & v8455ab;
assign v3743c44 = hgrant3_p & v35b7299 | !hgrant3_p & v3766105;
assign v3754922 = hgrant6_p & v37517d2 | !hgrant6_p & !v3a702f7;
assign v3a70e54 = hbusreq8 & v3a5d6f3 | !hbusreq8 & v3773ccd;
assign v37639c6 = hlock2 & v376e833 | !hlock2 & v3735809;
assign v3a5cb20 = hlock7_p & v8455ab | !hlock7_p & v3772f3c;
assign v37644ee = hlock7 & v3766232 | !hlock7 & v374b972;
assign v373cbc2 = hbusreq4 & v3779860 | !hbusreq4 & v8455ab;
assign v3a70b2a = hmaster3_p & v37478dd | !hmaster3_p & !v3759d9c;
assign v372797f = hbusreq6 & v3a6f2d7 | !hbusreq6 & v376ef7a;
assign v3a70986 = hbusreq6_p & v372ea14 | !hbusreq6_p & v37571f1;
assign v37447f7 = hmaster2_p & v375d3cd | !hmaster2_p & v3a700d8;
assign v373e891 = hlock5 & v3765f5c | !hlock5 & v3a7040e;
assign v377b690 = hgrant1_p & v3a55e7d | !hgrant1_p & !v8455ab;
assign v37698a1 = hmaster2_p & v3734062 | !hmaster2_p & v374f178;
assign v37658f9 = hgrant4_p & v8455ab | !hgrant4_p & v3a70a5e;
assign v374f077 = hmaster0_p & v3758672 | !hmaster0_p & v373185b;
assign v374510a = hbusreq8_p & v3a580e3 | !hbusreq8_p & v8455ab;
assign v3a630db = hlock4_p & v372abd8 | !hlock4_p & v35772a6;
assign v3a70976 = hgrant3_p & v372919a | !hgrant3_p & v373d139;
assign v3a54120 = hlock8_p & v375eea5 | !hlock8_p & v3a5a2e5;
assign v3a7115c = hlock5 & v3a60826 | !hlock5 & v377efa7;
assign v3725e4b = hmaster2_p & v375121b | !hmaster2_p & !v3a6f59d;
assign v3577421 = hbusreq4_p & v3726d1f | !hbusreq4_p & v376c76d;
assign v3a6ffe7 = hgrant6_p & v8455ab | !hgrant6_p & v3746cdc;
assign v37774d3 = hmaster2_p & v376fe6e | !hmaster2_p & v37425a5;
assign v374ff02 = hbusreq7_p & v3a6d5a8 | !hbusreq7_p & !v377a9b2;
assign v3727dd4 = hbusreq6_p & v3a6ef23 | !hbusreq6_p & v377bb21;
assign v37243d7 = hbusreq3_p & v3759b2f | !hbusreq3_p & !v373be25;
assign v3a6738e = hbusreq7_p & v376bd2f | !hbusreq7_p & v37446e0;
assign v3a6bdd7 = hgrant1_p & v3a70e9a | !hgrant1_p & v8455ab;
assign v377d999 = hbusreq8 & v372aff0 | !hbusreq8 & v37395d4;
assign v3754422 = hlock6 & v3734f70 | !hlock6 & v3a6f77e;
assign v3738b4c = hmaster2_p & v37738fc | !hmaster2_p & v3a6773a;
assign v3723923 = hmaster0_p & v377d1dc | !hmaster0_p & v3745589;
assign v3735d9c = hgrant4_p & v3a6f35c | !hgrant4_p & v3a5f26f;
assign v3a65a33 = hgrant3_p & v8455ab | !hgrant3_p & v37435f6;
assign v3a712b2 = hgrant6_p & v3a5b5d3 | !hgrant6_p & v376fafe;
assign v373e827 = hgrant6_p & v3a71685 | !hgrant6_p & !v8455ab;
assign v3737dad = hbusreq0 & v373f8b1 | !hbusreq0 & v3a6f322;
assign v374407c = hmaster1_p & v8455ab | !hmaster1_p & !v3767471;
assign v37435f1 = hbusreq8 & v3a6869d | !hbusreq8 & v3a70f23;
assign v3a584d6 = hbusreq5_p & v3a635ea | !hbusreq5_p & v377af11;
assign v372bdd9 = hbusreq4 & v377349f | !hbusreq4 & v37684a8;
assign v3a658c0 = hlock6_p & v8455ab | !hlock6_p & !v374e77f;
assign v3a712c4 = hgrant4_p & v8455ab | !hgrant4_p & v3a713c8;
assign v375b5eb = hbusreq5_p & v3739ab2 | !hbusreq5_p & !v3a5c998;
assign v376075c = hmaster0_p & v3a6dfb2 | !hmaster0_p & v3a6fc2b;
assign v376dad4 = hmaster0_p & v3a61480 | !hmaster0_p & v3753a65;
assign v3a70f8c = hbusreq5 & v3a6ef2c | !hbusreq5 & v376cd02;
assign v3a70d21 = hbusreq5 & v3769d4c | !hbusreq5 & v39a4e1f;
assign v37530d1 = hgrant5_p & v8455c9 | !hgrant5_p & v2ff8d08;
assign v373149a = hmaster1_p & v8455ab | !hmaster1_p & v3778f19;
assign v372de68 = hgrant4_p & v3a6f585 | !hgrant4_p & v3774075;
assign v3a6a493 = hgrant6_p & v8455ab | !hgrant6_p & v3775d76;
assign v3a5d34b = hbusreq0_p & v3737462 | !hbusreq0_p & v35772a6;
assign v375ceff = hmaster2_p & v372424e | !hmaster2_p & v38092e6;
assign v3a5b86c = hmaster0_p & v3a635ea | !hmaster0_p & v3755738;
assign v3a6eefb = hmaster2_p & v3a5d4d0 | !hmaster2_p & v96dd76;
assign v3a6a187 = stateA1_p & v8455e1 | !stateA1_p & !v3749e1c;
assign v3774e8c = hgrant0_p & v8455ab | !hgrant0_p & v376d15d;
assign v3734ab5 = hmaster1_p & v376c2e6 | !hmaster1_p & v3a70217;
assign v375306b = hlock6_p & v3a68426 | !hlock6_p & v8455b7;
assign v372a64f = hbusreq7_p & v375b84e | !hbusreq7_p & v3a69203;
assign v3770717 = hbusreq5 & v3a66ade | !hbusreq5 & v3778c64;
assign v3a6fbf4 = hbusreq1_p & v3a6fc6c | !hbusreq1_p & v3752dbb;
assign v374b225 = hmaster1_p & v3a56230 | !hmaster1_p & v3770eeb;
assign v374c164 = hmaster2_p & v3752d2c | !hmaster2_p & v377b94f;
assign v3a70ede = hmaster2_p & v37672af | !hmaster2_p & v3a5d36a;
assign v37441a3 = hbusreq7 & v3a65755 | !hbusreq7 & v372fdd0;
assign v37640de = hmaster2_p & v372e0b0 | !hmaster2_p & v3a67869;
assign v376711c = hgrant2_p & v8455ab | !hgrant2_p & bf3e2b;
assign v3724581 = hready & v8455ab | !hready & v373d9e5;
assign v37596fd = hgrant1_p & v3a6f10f | !hgrant1_p & v8455ab;
assign v37521f6 = hbusreq4_p & v3729ed7 | !hbusreq4_p & cbd026;
assign v374dd8f = hmaster2_p & v375d3cd | !hmaster2_p & v3a705a8;
assign v3a71193 = hgrant5_p & v3a6f5ff | !hgrant5_p & v37476c5;
assign v3740aa7 = hmaster2_p & v8455c3 | !hmaster2_p & v3a6f0f9;
assign v3a6f322 = hgrant6_p & v3727cd0 | !hgrant6_p & v377e2f7;
assign v376832f = hmaster0_p & v3a61410 | !hmaster0_p & v3a6e8d9;
assign v3751925 = hmaster2_p & v374ad7d | !hmaster2_p & v3724a4b;
assign v3a6c6ad = hmaster2_p & v3a5a807 | !hmaster2_p & v376b4ad;
assign v3735134 = hbusreq6 & v373d551 | !hbusreq6 & v374aca8;
assign v37287f6 = hmaster2_p & v376ce77 | !hmaster2_p & v373c21c;
assign v374eab3 = hmaster2_p & v37590a2 | !hmaster2_p & v37697a3;
assign v3a70ca8 = hbusreq2_p & v8455e7 | !hbusreq2_p & v8455ab;
assign v375789b = hmaster2_p & v39a4dac | !hmaster2_p & !v8455ab;
assign v37702c5 = hbusreq5_p & v37337f1 | !hbusreq5_p & !v372e6d3;
assign v373385b = hmaster0_p & v23fe361 | !hmaster0_p & v377f5db;
assign v37357d9 = hmaster0_p & v373a222 | !hmaster0_p & !v3a61c70;
assign v3a5aa42 = hmaster3_p & v8455ab | !hmaster3_p & v372dbb0;
assign v377cc7b = hlock5_p & b6a7cc | !hlock5_p & v8455ab;
assign v3a63ff3 = hgrant3_p & v372d02d | !hgrant3_p & v375c806;
assign v3a661d0 = hmaster1_p & v3a299cd | !hmaster1_p & v3a64879;
assign v3a70d5d = hmaster0_p & v372fa3a | !hmaster0_p & v372efcd;
assign v375f84b = hmaster2_p & v3743ff2 | !hmaster2_p & v9bf1d8;
assign v3a7153c = hbusreq4_p & v3a668a4 | !hbusreq4_p & v8455ab;
assign v377981a = hgrant5_p & v3756d6e | !hgrant5_p & v372a704;
assign v3a5cc77 = hmaster2_p & v3752536 | !hmaster2_p & !v3a70fec;
assign v3a6a295 = hbusreq0 & v37621eb | !hbusreq0 & v3742a27;
assign v37596c8 = hbusreq3_p & v37729ac | !hbusreq3_p & v8455ab;
assign v3769310 = hmaster1_p & v377050c | !hmaster1_p & v3a6f54b;
assign v376ab39 = hmaster0_p & v377e31b | !hmaster0_p & v3738ed8;
assign v3739078 = hbusreq0 & v3a62f06 | !hbusreq0 & v38072fd;
assign v37737d2 = hmaster1_p & v3a6f443 | !hmaster1_p & v3a6d140;
assign v3777d79 = hbusreq3_p & v377934a | !hbusreq3_p & v3732302;
assign v3767e7f = hmaster0_p & v37564d1 | !hmaster0_p & v3a59649;
assign v3778e03 = hgrant2_p & v3751a33 | !hgrant2_p & v3761cbb;
assign v3738dac = hbusreq4_p & v3a603a1 | !hbusreq4_p & v3778528;
assign v37741bd = hmaster0_p & v8455ab | !hmaster0_p & v3a625a1;
assign v3a59b42 = jx0_p & v377dac2 | !jx0_p & v374d529;
assign v37300d3 = hmaster1_p & v8455ab | !hmaster1_p & v373d5f0;
assign v377b4f2 = hgrant3_p & v8455ab | !hgrant3_p & v3a61b7f;
assign v3a62e77 = hmaster1_p & v3726c61 | !hmaster1_p & v373e941;
assign v3a70b8a = hgrant6_p & v377938d | !hgrant6_p & v3a70d57;
assign v3a5aef6 = hmaster1_p & v3754892 | !hmaster1_p & v23fe052;
assign v373b46b = hgrant6_p & v375d861 | !hgrant6_p & v37407f5;
assign v374f178 = hgrant4_p & v3760bdd | !hgrant4_p & v375ecff;
assign v3a70a5c = hbusreq4_p & v37748b7 | !hbusreq4_p & v8455ab;
assign v37262ad = hlock5_p & v3a70641 | !hlock5_p & v3748446;
assign v3778023 = hbusreq8 & v374373a | !hbusreq8 & v3744c88;
assign v3747fda = hmaster2_p & v3740d3b | !hmaster2_p & v3725827;
assign v3a6fa06 = hgrant2_p & v8455ab | !hgrant2_p & v3a6de73;
assign v3734a4f = hlock5 & v373124d | !hlock5 & v3a6f7b3;
assign v373a33d = hbusreq4 & v37740d0 | !hbusreq4 & v3a62a6d;
assign v372479c = hbusreq2_p & v372493b | !hbusreq2_p & !v3a6febd;
assign v3a56ca1 = hgrant4_p & v3771697 | !hgrant4_p & v3a66381;
assign v3766c60 = hgrant4_p & v3a6fea9 | !hgrant4_p & v3a6b14a;
assign v3a59cde = hbusreq7_p & v376147a | !hbusreq7_p & !v8455ab;
assign v3a6f90f = hmaster2_p & v3a708a2 | !hmaster2_p & v8455ab;
assign v3730778 = hmaster0_p & v3a7113c | !hmaster0_p & v3753055;
assign v3a56b05 = hgrant4_p & v8455ab | !hgrant4_p & v37605fb;
assign v373568c = hgrant3_p & v37647e7 | !hgrant3_p & v3a6f9f8;
assign a97cd0 = hmaster2_p & v3763030 | !hmaster2_p & v8455ab;
assign v3748e9d = hbusreq0 & c3d672 | !hbusreq0 & v37362d7;
assign v3a6f78a = hlock0 & v376c76d | !hlock0 & v3765021;
assign v209300d = hbusreq4 & v377a1d3 | !hbusreq4 & v374f35a;
assign v375b92a = hlock4_p & v3a5be93 | !hlock4_p & v3a6fd81;
assign v375d30b = hgrant3_p & v3a6c2b6 | !hgrant3_p & !v2ff8f1e;
assign v3a6cf7f = hmaster2_p & v37632f8 | !hmaster2_p & v3734067;
assign v3764af3 = hgrant2_p & v8455ab | !hgrant2_p & v3a70a55;
assign v37599b8 = jx0_p & v3728d75 | !jx0_p & v37708bb;
assign v3a6f537 = hbusreq5 & v3a71133 | !hbusreq5 & v3a5f12b;
assign v3759837 = hbusreq4 & v373a4e4 | !hbusreq4 & v3a70d99;
assign beb1cf = hbusreq6_p & v3a70937 | !hbusreq6_p & !v374e28f;
assign v37479b4 = hgrant0_p & v8455ab | !hgrant0_p & v2619ad3;
assign v3806a7a = hbusreq8 & v373e8e3 | !hbusreq8 & v374a39f;
assign v377c261 = hmaster0_p & v377d742 | !hmaster0_p & v3a5c3ba;
assign v3748251 = hbusreq8_p & v37539c8 | !hbusreq8_p & v377f501;
assign v374f351 = hgrant2_p & v375b7b5 | !hgrant2_p & v8455ab;
assign v374df1b = hbusreq6 & v3729f32 | !hbusreq6 & v8455ab;
assign v373c768 = hgrant6_p & v3755785 | !hgrant6_p & v3a5c2df;
assign v37492d2 = hmaster1_p & v3a64361 | !hmaster1_p & v375a51f;
assign v3a61f46 = hmaster0_p & v3736ded | !hmaster0_p & v3a57e6d;
assign v3a71393 = hlock6 & v3a643d7 | !hlock6 & v3a714b3;
assign v37314cb = hlock4_p & v37565c7 | !hlock4_p & v3a6cdd4;
assign v37367a0 = hbusreq0 & v374cab9 | !hbusreq0 & !v8455ab;
assign v3773e09 = hbusreq2 & v372ee9a | !hbusreq2 & v3a6be44;
assign v377ed71 = stateG10_1_p & v35772a5 | !stateG10_1_p & !v3774d04;
assign v372a399 = hbusreq0_p & v3a5e9d3 | !hbusreq0_p & v3743b9e;
assign v3a714ed = hbusreq7 & v3a5e245 | !hbusreq7 & !v8455b9;
assign v3769f7f = hbusreq5_p & v3a63f66 | !hbusreq5_p & v8455ab;
assign v3a60826 = hbusreq5 & v377efa7 | !hbusreq5 & v374f345;
assign v1e382f1 = hbusreq8 & v37383b1 | !hbusreq8 & v3735049;
assign v37572c1 = hgrant4_p & v8455ab | !hgrant4_p & v3754a4d;
assign v3747398 = hgrant1_p & v3728ea6 | !hgrant1_p & v8455ab;
assign v3a5a09c = hbusreq3_p & v3733c39 | !hbusreq3_p & v3754e7b;
assign v3a629a9 = hmaster3_p & v3a65760 | !hmaster3_p & v3a628ef;
assign v374592e = start_p & v8455ab | !start_p & v3a5a496;
assign v374641d = hbusreq4 & v3a70e5b | !hbusreq4 & v373031f;
assign v372b906 = hbusreq4 & v3753d51 | !hbusreq4 & v3a70bb7;
assign v377348f = hmaster2_p & v3a70c39 | !hmaster2_p & v37386cb;
assign v1e37a30 = hbusreq7_p & v3a62f05 | !hbusreq7_p & v375be2d;
assign v3761b23 = hlock5 & v3a58bae | !hlock5 & v376c5d3;
assign v377bb57 = hmaster2_p & v3a70326 | !hmaster2_p & v3a5fdd3;
assign v3a66464 = hburst0 & v8455ab | !hburst0 & !v3745b85;
assign v3a64045 = hbusreq6_p & v376c6ed | !hbusreq6_p & v3776b9a;
assign v3742a4b = hbusreq5 & v373e93e | !hbusreq5 & v3752321;
assign b5f474 = hlock4 & v3a6f139 | !hlock4 & v376cf3f;
assign v3746c8d = hburst1_p & v845605 | !hburst1_p & v8455ab;
assign v3a6d8a9 = hbusreq8 & v372d561 | !hbusreq8 & v8455ab;
assign v377894b = hgrant2_p & v375975b | !hgrant2_p & v3a71098;
assign v3a59bbd = hmaster2_p & v3a6e985 | !hmaster2_p & v3751081;
assign v3748ca5 = hbusreq3_p & v3749ea2 | !hbusreq3_p & v8455ab;
assign v3a6087b = hmaster0_p & v374749d | !hmaster0_p & v3774bdf;
assign v372e27b = hbusreq4_p & v8455c3 | !hbusreq4_p & !v3a6a036;
assign v3a5bc5f = hmaster0_p & v3723211 | !hmaster0_p & v3a5a226;
assign v376a915 = hmaster0_p & v377766c | !hmaster0_p & v37334fc;
assign v37286a2 = hgrant2_p & v8455b5 | !hgrant2_p & v3a5ccfd;
assign v375e50c = hbusreq5_p & v3a6eb22 | !hbusreq5_p & v3a6fbda;
assign v374fb8d = hbusreq4_p & v3a61ce7 | !hbusreq4_p & v8455cb;
assign v3731511 = hbusreq4_p & v373330f | !hbusreq4_p & v377aa06;
assign v3a69091 = jx0_p & v37466a5 | !jx0_p & v374da33;
assign v3729708 = hmaster0_p & v3a661fe | !hmaster0_p & v3a6fcd2;
assign v3747389 = hbusreq5 & v3a6f93b | !hbusreq5 & v8455ab;
assign v3741793 = hlock7 & v3a6f83b | !hlock7 & v373c4a7;
assign v3761f2b = hbusreq7_p & v3777d51 | !hbusreq7_p & v3731ea5;
assign v3749c27 = hlock0_p & v3778ed4 | !hlock0_p & v8455e7;
assign v37248c1 = hbusreq4 & v375f423 | !hbusreq4 & v8455ab;
assign v3772cc3 = hmaster1_p & v8455b5 | !hmaster1_p & v3a707b1;
assign v380925f = hmaster0_p & v37386c6 | !hmaster0_p & v3732c86;
assign v3a6ff9b = hbusreq2 & v37348ee | !hbusreq2 & v3a69487;
assign v3756305 = hbusreq5 & v375138c | !hbusreq5 & v3722a6f;
assign v3a6f4b2 = hlock6_p & v3722e5c | !hlock6_p & v35772a6;
assign v372a9c7 = hgrant4_p & v374f4a3 | !hgrant4_p & v2ff91fe;
assign v3809282 = hbusreq3 & v37270d9 | !hbusreq3 & v8455e7;
assign v3772c4d = jx0_p & v3a70605 | !jx0_p & v3a70c31;
assign v375c44b = hlock4_p & v377a965 | !hlock4_p & v374b18c;
assign v374db33 = hbusreq8 & v3a6fbfd | !hbusreq8 & !v3a70157;
assign v3a71254 = hgrant5_p & v8455ab | !hgrant5_p & v3a6ef01;
assign v375b483 = hlock5_p & v8455e7 | !hlock5_p & !v3a6fd3d;
assign v3765a79 = hmaster2_p & v8455ab | !hmaster2_p & v3732dc6;
assign v3a5e020 = hbusreq2 & v3751e09 | !hbusreq2 & v8455ab;
assign v377955b = hbusreq0 & v375ef36 | !hbusreq0 & v8455ab;
assign v3a6600a = hbusreq2 & v377e089 | !hbusreq2 & !v8455bd;
assign v3a5a6f4 = hbusreq2_p & v3778fb2 | !hbusreq2_p & v3a70d05;
assign v2aca789 = hgrant3_p & v376ace9 | !hgrant3_p & v3a6eab0;
assign v3a672de = hlock5_p & v374d383 | !hlock5_p & v3a672e6;
assign v3a62f60 = hlock4_p & v37716c3 | !hlock4_p & v3a7084e;
assign v3732da0 = hready_p & v374efeb | !hready_p & v3a6fceb;
assign v3a572ea = hmaster0_p & v3a5a807 | !hmaster0_p & v374c02e;
assign v3754c02 = hmaster0_p & v3734bd2 | !hmaster0_p & v375b0e4;
assign v375f883 = jx1_p & v3a607c3 | !jx1_p & v377c6b0;
assign v37471a7 = hmaster2_p & v374502e | !hmaster2_p & v3a6ab5f;
assign v3a65d93 = hmaster2_p & v3736f61 | !hmaster2_p & v376856b;
assign v3807bfa = hmaster1_p & v3a5762d | !hmaster1_p & v376abdf;
assign v376a907 = hmaster2_p & v3a702c2 | !hmaster2_p & v3a5f40e;
assign v3749eb2 = hbusreq0 & v3a6c39b | !hbusreq0 & v8455ab;
assign v37758de = hbusreq7 & v3776066 | !hbusreq7 & v375075b;
assign v3a70866 = hmaster0_p & v375bd8c | !hmaster0_p & v372e05a;
assign v375d95f = hmaster1_p & v37325c5 | !hmaster1_p & v374e21e;
assign v3764a58 = hbusreq8_p & v375a4c4 | !hbusreq8_p & v3722dd6;
assign v3a6cf88 = hgrant5_p & v3a70220 | !hgrant5_p & v3730094;
assign v3a707e5 = hbusreq7 & v37342cd | !hbusreq7 & !v8455ab;
assign v37654c4 = hmaster2_p & v3725c63 | !hmaster2_p & v3758166;
assign v3a64aa0 = hbusreq0 & v3727c62 | !hbusreq0 & v374d33d;
assign v3a70d9b = hgrant5_p & v377d91c | !hgrant5_p & v373fdf0;
assign v3a57867 = hmaster2_p & v3a619c0 | !hmaster2_p & !v3a5bf04;
assign v3723d55 = hbusreq3_p & v3760073 | !hbusreq3_p & v8455ab;
assign v3a6255b = hlock0_p & v8455ab | !hlock0_p & v8455b5;
assign v3a7062e = hgrant6_p & v3741acc | !hgrant6_p & v3774a7e;
assign v3a6f647 = hbusreq0 & v377293c | !hbusreq0 & v3a7159c;
assign v3a6f12a = hbusreq0 & v3a5a967 | !hbusreq0 & v3a7012d;
assign v3774cee = hbusreq6 & v37510b1 | !hbusreq6 & !v8455ab;
assign v3a7102a = jx1_p & v3a709de | !jx1_p & v3761930;
assign v3a70ed8 = hbusreq8_p & v3a713a9 | !hbusreq8_p & v3740e9c;
assign v376aad2 = hgrant6_p & v3a6f17e | !hgrant6_p & v3a5c350;
assign v373bdac = hburst1 & v8455ab | !hburst1 & v3758079;
assign v373593a = hbusreq0_p & v376d327 | !hbusreq0_p & v3a63621;
assign v377a1ee = hbusreq5_p & v3731724 | !hbusreq5_p & v1e3786e;
assign v3766472 = hmaster1_p & v37494c3 | !hmaster1_p & v3735d84;
assign v3a6a0b0 = hbusreq2 & v8455b0 | !hbusreq2 & v37406d2;
assign v3779c2b = hlock0 & v3a6efad | !hlock0 & v2acaed3;
assign v375f9ec = hbusreq0 & v373e09b | !hbusreq0 & v373c768;
assign v3734291 = hbusreq3 & v374f87c | !hbusreq3 & v8455ab;
assign v3a57912 = hmaster2_p & v3a70f7f | !hmaster2_p & v3764568;
assign v2925c67 = hbusreq3 & v3a7037c | !hbusreq3 & v8455ab;
assign v3730fcd = hlock4_p & v3a6910c | !hlock4_p & v3731e7b;
assign v3a5af41 = hbusreq7_p & v375075b | !hbusreq7_p & v3a6fe04;
assign v360d1ca = hgrant1_p & v3777705 | !hgrant1_p & v8455ab;
assign v372588c = hmaster1_p & v373a1d0 | !hmaster1_p & v37418db;
assign v38068ec = hmaster2_p & v3a6e31f | !hmaster2_p & v3a6d684;
assign v3a6eb6a = hmaster2_p & v3a5fc34 | !hmaster2_p & v373c21c;
assign v375e29b = hmaster1_p & v3750f77 | !hmaster1_p & v8455ab;
assign v3747db9 = hmaster3_p & v372c49f | !hmaster3_p & v377a2d1;
assign v3a6eb86 = hgrant0_p & v37773a9 | !hgrant0_p & v3777fc5;
assign v372c571 = hgrant4_p & v8455ab | !hgrant4_p & v372cfbf;
assign v373cca3 = hready & v37563eb | !hready & !v8455ab;
assign v3a6f3fb = hbusreq0 & v37463e5 | !hbusreq0 & v3a5cf78;
assign v375d161 = hgrant3_p & v372d02d | !hgrant3_p & v3a6eb01;
assign v3a705c5 = hbusreq2_p & v375b445 | !hbusreq2_p & v8455ab;
assign v375f071 = hbusreq5_p & v3a71116 | !hbusreq5_p & !v8455ab;
assign v373cf42 = hlock0_p & v376ef42 | !hlock0_p & v3a70c07;
assign v37315ae = hgrant8_p & v377fc58 | !hgrant8_p & v3a71112;
assign v376f693 = start_p & v845605 | !start_p & v865472;
assign v3756045 = hmaster0_p & v3a6aef7 | !hmaster0_p & v372c46e;
assign v376799e = hbusreq2_p & v3a6eb6b | !hbusreq2_p & v372f532;
assign v3768b46 = hbusreq4_p & v8455bf | !hbusreq4_p & v3a55bd0;
assign v37702a1 = hbusreq5 & v372e40f | !hbusreq5 & !v377ce1c;
assign v3737ca2 = hbusreq8_p & v3736b0e | !hbusreq8_p & v35b774b;
assign v3a290f9 = hgrant4_p & v3a62508 | !hgrant4_p & v3a715b2;
assign v3a7130f = hbusreq5 & v375b483 | !hbusreq5 & v8455c7;
assign v375ac20 = hlock0_p & v372feb2 | !hlock0_p & !v8455ab;
assign v3a5857c = hmaster1_p & v3736ded | !hmaster1_p & v3a61f46;
assign v3776e45 = hlock7 & v3a6f31e | !hlock7 & v3739493;
assign v37317ba = hbusreq3 & v377989c | !hbusreq3 & v8455ab;
assign v377b07a = hmaster2_p & v3760f87 | !hmaster2_p & v8455ab;
assign v3a5f1d4 = hbusreq4_p & v3747302 | !hbusreq4_p & v3743b9e;
assign v37585c9 = hgrant5_p & v8455ab | !hgrant5_p & v3756c22;
assign v3770c4c = hgrant6_p & v373c81c | !hgrant6_p & v3a59dc4;
assign v3a6a2b5 = hbusreq6_p & v372864a | !hbusreq6_p & v3776e85;
assign v3743cf5 = hbusreq7 & v3a70454 | !hbusreq7 & v374d617;
assign v3a6fa97 = hmaster2_p & v8455ab | !hmaster2_p & !v3742cd4;
assign v3a6fbc2 = hlock8_p & v372dbe1 | !hlock8_p & !v8455ab;
assign v3a5846c = hgrant2_p & v8455ab | !hgrant2_p & v3a66c5c;
assign v373a85c = hmaster2_p & v3a6f8af | !hmaster2_p & v8455ab;
assign v3a70479 = hmaster2_p & v3a62a6d | !hmaster2_p & v3a5cfac;
assign v3a5ce1e = hgrant2_p & v377cbad | !hgrant2_p & v37798aa;
assign v3a6ebd3 = hgrant2_p & v3748792 | !hgrant2_p & v3a70f37;
assign v3a6cb5b = hmaster1_p & v8455ab | !hmaster1_p & v372b7a5;
assign v376bf8d = hlock0_p & v3770993 | !hlock0_p & v3a6f4b6;
assign v3a66e6f = hmaster0_p & v3a53a2d | !hmaster0_p & v3a700db;
assign v37790df = hgrant2_p & v3a6305e | !hgrant2_p & v3742655;
assign v3734913 = hgrant6_p & v8455ab | !hgrant6_p & v376efdb;
assign v3a70bf9 = hbusreq8 & v374cd15 | !hbusreq8 & v376cef0;
assign v3a700ce = hmaster2_p & v3739b80 | !hmaster2_p & !v374a2cc;
assign v3a705f4 = hlock6_p & v8455ab | !hlock6_p & v3a5e363;
assign v3a6fd22 = hbusreq5 & v3a695a8 | !hbusreq5 & v3a692da;
assign v377a083 = hmaster2_p & v3a6e13d | !hmaster2_p & v3732b75;
assign v374da93 = hlock5_p & v3771fec | !hlock5_p & !v377c500;
assign v3a5d704 = hbusreq8_p & v39ebb5d | !hbusreq8_p & v377bf2b;
assign v3a71248 = hmaster2_p & v37390c5 | !hmaster2_p & v3754aa3;
assign v3748e0b = hbusreq6 & v3725091 | !hbusreq6 & v3a56e79;
assign v1e37d82 = hmaster2_p & v8455ab | !hmaster2_p & !v3772add;
assign v37665c5 = hgrant4_p & v8455ab | !hgrant4_p & v3a6ebb8;
assign v3a700f8 = hbusreq6 & v37521ed | !hbusreq6 & !v8455ab;
assign v37502b7 = locked_p & v3a5bd24 | !locked_p & v3809adf;
assign v37719a0 = hlock5 & v3777d37 | !hlock5 & v372cb8c;
assign v3a5c9df = hbusreq5_p & v3a6fb2f | !hbusreq5_p & v3738666;
assign v3a6fee9 = hgrant3_p & v3779cf9 | !hgrant3_p & v3a5a09c;
assign v37348c9 = jx1_p & v3758a11 | !jx1_p & v8455ab;
assign v37751cb = hmaster1_p & v3a70987 | !hmaster1_p & v376a3aa;
assign v3726777 = hbusreq3 & v3807c0c | !hbusreq3 & v375cf36;
assign v3a71030 = hgrant5_p & v372b0b0 | !hgrant5_p & v372d59d;
assign v3725d48 = hbusreq5_p & v3a6b29f | !hbusreq5_p & v3747e73;
assign v37233a7 = hlock4 & v3736b57 | !hlock4 & v3750f8f;
assign v37615ce = hgrant4_p & v373f17f | !hgrant4_p & v3774653;
assign v3a6f557 = hbusreq2_p & v37510ae | !hbusreq2_p & v37563fe;
assign v375e6fc = hgrant5_p & v376bd96 | !hgrant5_p & v373ce36;
assign v3a70d69 = hlock5_p & v373c15d | !hlock5_p & v37251f1;
assign v3756f77 = hmaster2_p & v377d74c | !hmaster2_p & v3a55419;
assign v377caa3 = hlock3_p & v3379037 | !hlock3_p & !v8455ab;
assign v37793b9 = hmaster2_p & v3770bcd | !hmaster2_p & v377c28e;
assign v3a70562 = hbusreq4 & v374922a | !hbusreq4 & !v8455ab;
assign v3a58dfb = hmaster3_p & v3771232 | !hmaster3_p & v3a6f232;
assign v37720e5 = hbusreq3 & v3a57309 | !hbusreq3 & v8455ab;
assign v376660c = hbusreq6 & v3a70d79 | !hbusreq6 & v8455ab;
assign v372981a = hmaster1_p & v1e37bde | !hmaster1_p & v376fcd6;
assign v3745706 = hbusreq5 & v3729fa4 | !hbusreq5 & v3a55bd3;
assign v37627a8 = hmaster1_p & v3a6fdb3 | !hmaster1_p & v3a6f5c6;
assign v373ae0a = hbusreq0 & v372edf9 | !hbusreq0 & v3a69d13;
assign v37610ce = hmaster1_p & v375ede6 | !hmaster1_p & v3a683c6;
assign v376d883 = hbusreq5_p & v372998e | !hbusreq5_p & v377249b;
assign v3748262 = hmaster2_p & v3a70374 | !hmaster2_p & v3a70e28;
assign v3773a45 = hgrant2_p & v3758472 | !hgrant2_p & v3a70568;
assign v373c4d4 = hbusreq0 & v3a702de | !hbusreq0 & v3a588ef;
assign v37409cd = hmaster2_p & v37289f0 | !hmaster2_p & v3769740;
assign v3a6a880 = hbusreq6 & v3764f27 | !hbusreq6 & v8455ab;
assign v373f06c = hlock5_p & v3a6f749 | !hlock5_p & v37511c6;
assign v3a68463 = hbusreq2 & v3a598a0 | !hbusreq2 & v376e041;
assign v3a6f352 = hmaster0_p & v3735891 | !hmaster0_p & v374c5c5;
assign v37378ca = hbusreq3_p & v3777870 | !hbusreq3_p & v8455ab;
assign v375d886 = hlock5 & v3a71687 | !hlock5 & v3724c63;
assign v3a6f09c = hbusreq6 & v374362e | !hbusreq6 & v3a676d6;
assign v3a67dc7 = hlock3_p & v2925c39 | !hlock3_p & !v8455ab;
assign v3768c25 = hmaster2_p & v3735272 | !hmaster2_p & v3a5b576;
assign v38097f6 = hlock6_p & v3a6f213 | !hlock6_p & !v3a6fe1a;
assign v373146d = hgrant6_p & v3a5cb5f | !hgrant6_p & v3737bc8;
assign v3a7129b = hgrant6_p & v372bfa1 | !hgrant6_p & v3a5b3d8;
assign v2acaf41 = hlock6_p & v3806db7 | !hlock6_p & v8455b0;
assign v3732558 = hlock5_p & v3770827 | !hlock5_p & !v8455ab;
assign v3a5841e = hbusreq4 & v37457fb | !hbusreq4 & v8455ab;
assign v2acaeaa = hmaster1_p & v373fa3d | !hmaster1_p & v3772409;
assign v372f85e = hgrant0_p & v8455e7 | !hgrant0_p & v3766e3a;
assign v23fe052 = hbusreq5_p & v3767744 | !hbusreq5_p & v3749cf4;
assign v3754379 = hmaster0_p & v3a635ea | !hmaster0_p & v3a6fcfd;
assign v373197c = hmaster2_p & v3a5be74 | !hmaster2_p & v3750d27;
assign v3749bef = hgrant2_p & v3767304 | !hgrant2_p & v3a6f5f6;
assign v3777610 = hlock5 & v3a63f9a | !hlock5 & v3734fba;
assign v377f526 = hbusreq0 & v3746063 | !hbusreq0 & v8455ab;
assign v3a69123 = hmaster2_p & v3777bde | !hmaster2_p & v374892a;
assign v372945c = hmaster0_p & v3742582 | !hmaster0_p & v3a706cb;
assign v3378b6c = hmaster1_p & v3758fa8 | !hmaster1_p & v3a7031c;
assign v3744824 = hlock7 & v372f3a4 | !hlock7 & v3a6b0eb;
assign v37751c3 = jx0_p & v377c97f | !jx0_p & v3a706e6;
assign v37645a4 = hbusreq6 & v3a55173 | !hbusreq6 & v8455ab;
assign v3768774 = hbusreq5_p & v3a6eede | !hbusreq5_p & !v3745b66;
assign v3a62e1e = hlock2 & v373a802 | !hlock2 & v3a6440f;
assign v376c9a5 = jx0_p & v376596c | !jx0_p & v372d764;
assign v3a5bf04 = locked_p & v3a563ad | !locked_p & v1e38224;
assign v23fdea8 = jx1_p & v3734c59 | !jx1_p & v375d758;
assign v372883e = hmaster2_p & v3a70374 | !hmaster2_p & v3a71134;
assign v372e30d = hlock2 & v3748797 | !hlock2 & v2092f5e;
assign v373040b = hmaster2_p & v3a6f213 | !hmaster2_p & v8455ab;
assign v3729022 = hbusreq6_p & v376f56d | !hbusreq6_p & v374c6b1;
assign v372a0a1 = hbusreq5_p & v372f1e9 | !hbusreq5_p & v3756dd6;
assign v375548b = hbusreq5_p & v8dfd63 | !hbusreq5_p & v37541b4;
assign v377a2e1 = hmaster0_p & v3738253 | !hmaster0_p & v376a941;
assign v373120c = hbusreq6 & v373abb7 | !hbusreq6 & v3a702a7;
assign v3a65b00 = hbusreq7_p & v3768f71 | !hbusreq7_p & !v3736d1d;
assign v3752da9 = hbusreq8 & v3a57b5a | !hbusreq8 & v3a592d8;
assign v37381eb = hgrant2_p & v375d12e | !hgrant2_p & v3a5a1ba;
assign v374243d = hbusreq0 & v3a6f4af | !hbusreq0 & v372e873;
assign v3a5fa25 = hbusreq2 & v372c3df | !hbusreq2 & !v3a69515;
assign v373052f = hmaster1_p & v37640e9 | !hmaster1_p & v3743018;
assign v3776c43 = hbusreq3_p & v3a682cb | !hbusreq3_p & v3a658bf;
assign v3a6fc11 = hgrant2_p & v90829e | !hgrant2_p & v3a6613e;
assign v3a715f7 = hmaster2_p & v376a31b | !hmaster2_p & v376da22;
assign v377b946 = hbusreq6_p & v37496fa | !hbusreq6_p & v3743b9e;
assign v3a54bc5 = hbusreq3 & v3745f76 | !hbusreq3 & !v8455ab;
assign v3a70f3f = jx1_p & v866387 | !jx1_p & v8455ab;
assign v3756de3 = hbusreq4 & v376e17e | !hbusreq4 & v3724be1;
assign v374d648 = hgrant6_p & v372825b | !hgrant6_p & b1ca9b;
assign v3777c0c = hmaster0_p & v3a70d99 | !hmaster0_p & v3728cdc;
assign v3751100 = hlock4_p & v3a70cdb | !hlock4_p & v3755791;
assign v37389b1 = hbusreq7_p & v3a710ae | !hbusreq7_p & v3752f43;
assign v3a555ae = hmaster0_p & v3a6fe8d | !hmaster0_p & v8455ab;
assign v3a70cf1 = hbusreq5_p & v372b164 | !hbusreq5_p & v374a11d;
assign v3a6efb0 = hbusreq5 & a50cea | !hbusreq5 & v374e016;
assign v373b744 = hgrant1_p & v376bf04 | !hgrant1_p & !v37270d9;
assign v3a63dde = hbusreq8_p & v3a5567a | !hbusreq8_p & v3756b7b;
assign v3a6f9f6 = hbusreq2 & v8455b0 | !hbusreq2 & v3a63805;
assign v3a53962 = hgrant7_p & v3a70a85 | !hgrant7_p & v373d119;
assign v3a598a9 = hbusreq6_p & v3773e34 | !hbusreq6_p & v3750c0d;
assign v373a4b2 = hmaster1_p & v377cc6d | !hmaster1_p & v375e62f;
assign v3777517 = hbusreq5 & v3a6bf3c | !hbusreq5 & v373790d;
assign v375aa07 = hmaster1_p & v372455c | !hmaster1_p & v376f9a1;
assign v3724a10 = hgrant5_p & v8455b5 | !hgrant5_p & v3a709da;
assign v3a6f42a = hbusreq4_p & v377d9aa | !hbusreq4_p & !v8455ab;
assign v3746404 = hlock0_p & v3a70cdb | !hlock0_p & v3755791;
assign v3727849 = hbusreq6_p & v3731599 | !hbusreq6_p & v8455ab;
assign v37719b4 = hlock0_p & v3747c3e | !hlock0_p & v8455ab;
assign v3a567ec = hbusreq0 & v37438ab | !hbusreq0 & v3757921;
assign v3a5373e = hbusreq5_p & v37731ce | !hbusreq5_p & v374bfd2;
assign v3a7151e = hlock4 & v3751090 | !hlock4 & v1e37b3f;
assign v3a708c8 = hmaster0_p & v37469c4 | !hmaster0_p & v2ff8c74;
assign v3764811 = hbusreq5_p & v1e3737d | !hbusreq5_p & v3a5fc48;
assign v376441d = hgrant3_p & v8455ab | !hgrant3_p & v3a70418;
assign v3776e8b = hbusreq6_p & v3742b24 | !hbusreq6_p & v376dab5;
assign v3779627 = hmaster2_p & v3736ded | !hmaster2_p & v37716c3;
assign v3a7102f = hmaster0_p & v3a61a7f | !hmaster0_p & v37777d5;
assign v3a6f063 = hbusreq8_p & v3808f3c | !hbusreq8_p & ac6831;
assign v3758fae = jx1_p & v374b237 | !jx1_p & !v375811b;
assign v373a02b = hmaster2_p & v37520c4 | !hmaster2_p & v3756ecd;
assign v376663a = hlock0 & v3745f9b | !hlock0 & v37522ff;
assign v372b1e3 = hlock0 & v3a5b6de | !hlock0 & v3735051;
assign v373e09b = hgrant6_p & v3755785 | !hgrant6_p & v23fe098;
assign v3747d69 = jx0_p & v3a66988 | !jx0_p & v3a7162b;
assign v374430e = hmaster2_p & v3a67d66 | !hmaster2_p & v3770415;
assign v375355c = hlock5_p & v3a70348 | !hlock5_p & v372d92b;
assign v3a5a801 = hbusreq5_p & v8455ab | !hbusreq5_p & v3a7079f;
assign v377f2ea = hbusreq6 & v37740d0 | !hbusreq6 & v3a62a6d;
assign v3a6f71a = hbusreq2_p & v375da10 | !hbusreq2_p & v376bb26;
assign v3a616aa = hbusreq8 & v3a711c8 | !hbusreq8 & v3a6f95b;
assign v377816f = hmaster0_p & v3a5f744 | !hmaster0_p & v3a6a998;
assign v3a59d47 = hbusreq6_p & v3a62a8c | !hbusreq6_p & v3a70d42;
assign v374b64d = jx2_p & v37662f4 | !jx2_p & v3a61c5e;
assign v3a70aa3 = hmaster1_p & v2619aa7 | !hmaster1_p & v377e904;
assign v3778352 = hbusreq4 & v3a6fb2b | !hbusreq4 & v8455bf;
assign v3a5bf5f = hgrant4_p & v374f95d | !hgrant4_p & v3a6827b;
assign v3a70c9b = hgrant6_p & v3773044 | !hgrant6_p & v3a5ce1e;
assign v3760ba8 = hbusreq6_p & v95d97e | !hbusreq6_p & v373a391;
assign v3749a6b = hbusreq4 & v3754e78 | !hbusreq4 & v377b946;
assign v37528b9 = hbusreq3 & v3747994 | !hbusreq3 & v8455ab;
assign v3743040 = hlock6_p & aab2b0 | !hlock6_p & v8455e7;
assign v3a57508 = hbusreq5 & v375029a | !hbusreq5 & v372620f;
assign v3a70ab0 = hbusreq0 & v3777071 | !hbusreq0 & v3748797;
assign v3776be1 = hgrant2_p & v3a6f46a | !hgrant2_p & v3a5d717;
assign v3776685 = hbusreq2_p & v373e524 | !hbusreq2_p & v8455ab;
assign v374e531 = hbusreq6_p & v3a69f17 | !hbusreq6_p & !v35772a6;
assign v3a71448 = hgrant5_p & v373b91e | !hgrant5_p & v375dc43;
assign v3729798 = hbusreq5_p & v3a70f93 | !hbusreq5_p & v1e3737d;
assign v3a5e244 = hbusreq0 & v3a6f08a | !hbusreq0 & v3a712d1;
assign v3743eda = hgrant3_p & v8455e7 | !hgrant3_p & !v3738b0c;
assign v3a70c4c = hlock5_p & v37739ed | !hlock5_p & !v8455ab;
assign v37789a0 = hlock2 & v3a64e29 | !hlock2 & v3a67284;
assign v380946b = hlock0 & v1e378b4 | !hlock0 & v38078e5;
assign v374f307 = hready & v8455e7 | !hready & !v8455ab;
assign v3727a4d = hmaster2_p & v3764276 | !hmaster2_p & v3a653e4;
assign v3a6c9ab = hbusreq6_p & v3a6fb2b | !hbusreq6_p & v3749149;
assign v375c009 = hmaster1_p & v3a6546b | !hmaster1_p & v37542d8;
assign v3736e12 = hbusreq5 & v37450aa | !hbusreq5 & v3a709d3;
assign v3a65c2c = hmaster2_p & v3723eef | !hmaster2_p & v3754c5e;
assign v37321c2 = hlock4 & v3733716 | !hlock4 & v3a5b885;
assign v377ca3b = hgrant2_p & v3a5eadd | !hgrant2_p & v376f277;
assign v375d3bc = hbusreq4 & v3a58218 | !hbusreq4 & v8455ab;
assign v3770fef = hmaster2_p & v3759007 | !hmaster2_p & v37590d1;
assign v373ce74 = hgrant6_p & v37648af | !hgrant6_p & v3763299;
assign v373e642 = hbusreq3_p & v3a5a824 | !hbusreq3_p & v3a706b1;
assign v3739a9f = jx0_p & v376827d | !jx0_p & v376321e;
assign v375feb1 = hgrant3_p & v8455ab | !hgrant3_p & v3a6a8c5;
assign v3809af2 = hbusreq5_p & v8455ab | !hbusreq5_p & v3750c0c;
assign v3749580 = hbusreq5 & v3a6f106 | !hbusreq5 & v8455ab;
assign v3771a11 = hbusreq4_p & v3a5a807 | !hbusreq4_p & v3728c23;
assign v3a70964 = hbusreq0_p & v3735e39 | !hbusreq0_p & !v3a6d684;
assign v3a590de = hlock0_p & v3a635ea | !hlock0_p & !v3a65a24;
assign v3a71546 = hbusreq8 & v376cd19 | !hbusreq8 & v37431a0;
assign v3740bba = jx1_p & v37351a7 | !jx1_p & v8455ab;
assign v3a6fffc = hbusreq6 & ae0781 | !hbusreq6 & v3a708c2;
assign v37738d4 = hbusreq6 & v376dbdf | !hbusreq6 & v8455ab;
assign v373f996 = hbusreq5 & v372a77a | !hbusreq5 & v8455ab;
assign v3744d18 = hgrant2_p & v372493b | !hgrant2_p & v3759181;
assign v377529a = hmaster2_p & v8455ab | !hmaster2_p & v3a6cc65;
assign v374486d = hmaster2_p & v376e3fb | !hmaster2_p & v3728d9c;
assign v37602b1 = hmaster3_p & v377a916 | !hmaster3_p & v3754956;
assign v372dd2a = hlock7_p & v3a71124 | !hlock7_p & v374e5ab;
assign v3751364 = hbusreq3_p & v3a6fa9f | !hbusreq3_p & v3771c3a;
assign v377e784 = hgrant4_p & v3a637dc | !hgrant4_p & v3a66037;
assign v37331ff = hgrant4_p & v3a647df | !hgrant4_p & v372f91d;
assign a0d21b = hgrant6_p & v8455ca | !hgrant6_p & v3a5e0f7;
assign v3740690 = stateA1_p & v8455e1 | !stateA1_p & v3a293c5;
assign v3a70421 = hlock5_p & v3a640d1 | !hlock5_p & v3732871;
assign v373a9ee = hlock0 & v3a6fdef | !hlock0 & v37266c2;
assign v373049b = hmaster1_p & v373927b | !hmaster1_p & v3a566c1;
assign v373aaed = hmaster0_p & v3a6119e | !hmaster0_p & v3764015;
assign v3775750 = hbusreq2_p & v373997b | !hbusreq2_p & v37738fc;
assign v3761bb6 = hgrant2_p & v3779e45 | !hgrant2_p & v3730fd2;
assign v377a35c = hlock4_p & v373e209 | !hlock4_p & v377af44;
assign v3740451 = hbusreq7 & v3756afd | !hbusreq7 & v37332bf;
assign v37628f6 = hmaster1_p & v3a6ffb6 | !hmaster1_p & v3a5a806;
assign a7adce = hbusreq0 & v377ad57 | !hbusreq0 & v8455ab;
assign cdcddf = hmaster1_p & v8455ab | !hmaster1_p & v375a563;
assign v373eadd = hmaster0_p & v3a6a56e | !hmaster0_p & v8455ab;
assign v3a6efc4 = hmastlock_p & v3a648f2 | !hmastlock_p & v8455ab;
assign v3a6f40f = hmaster0_p & v3a6e5f0 | !hmaster0_p & v3a6dd80;
assign v360ba91 = decide_p & v3748851 | !decide_p & v3a5d9bc;
assign v3768695 = hmaster0_p & v8455ab | !hmaster0_p & v374636c;
assign v372d1ae = hlock5 & v3769cc4 | !hlock5 & v3a7017d;
assign v3745e54 = hgrant5_p & v8455ab | !hgrant5_p & v3758fa8;
assign v1e3780f = hgrant0_p & v3a64c10 | !hgrant0_p & !v3757082;
assign v374a096 = hlock6 & v372fe1b | !hlock6 & v3a5a8c3;
assign v3a64df4 = hlock5_p & v37596de | !hlock5_p & v2acb006;
assign v37693a3 = hbusreq5 & v3755aca | !hbusreq5 & v374e784;
assign v37390c4 = hbusreq3_p & v2ff9190 | !hbusreq3_p & v37508b2;
assign v373eb03 = hlock8 & v23fda4e | !hlock8 & v3747fbf;
assign v3a6958b = hbusreq3 & v3a64ee3 | !hbusreq3 & !v3a70131;
assign v37305e6 = hgrant5_p & v37530e8 | !hgrant5_p & v3731a95;
assign v372f2ae = hmaster0_p & v3a585d3 | !hmaster0_p & d26e1e;
assign v376de5c = hmaster0_p & v3728179 | !hmaster0_p & v3741357;
assign v3a551a4 = hbusreq1_p & v375356f | !hbusreq1_p & v8455ab;
assign v3750faa = hmaster2_p & v372ae9d | !hmaster2_p & !v3764978;
assign v3809505 = hlock5_p & v374e855 | !hlock5_p & v8455cb;
assign v375ab04 = hmaster3_p & v3a634b9 | !hmaster3_p & v3a66988;
assign v3726e81 = hlock6 & v3776125 | !hlock6 & v372310a;
assign v3a709cd = hlock8_p & v3727699 | !hlock8_p & !v3a6d5a8;
assign v377eb9d = hready & v8455ab | !hready & !v375e373;
assign v3756e87 = hmaster1_p & v3a6fa7a | !hmaster1_p & v3a6294e;
assign v37562fd = stateA1_p & v8455e1 | !stateA1_p & !v377c2e6;
assign v3766e4a = hgrant2_p & v38072fd | !hgrant2_p & v8455ab;
assign v31c329f = hready_p & v37346c5 | !hready_p & v8455df;
assign v376a943 = hbusreq4 & v3765739 | !hbusreq4 & v8455ab;
assign v3a70878 = hmaster1_p & v3749580 | !hmaster1_p & v3a2abf4;
assign v3a6c636 = hgrant2_p & v8455ab | !hgrant2_p & v3a53dff;
assign v3741ac2 = hmaster1_p & v377bb3a | !hmaster1_p & v374d645;
assign v3a6f7dd = hgrant4_p & v3775dbc | !hgrant4_p & v3a62070;
assign v3762d6e = hbusreq4_p & v3a6b3d4 | !hbusreq4_p & v3765f60;
assign v3739d9b = jx0_p & v3a70afd | !jx0_p & v9381f3;
assign v3a70380 = hlock5_p & v3a6ff8d | !hlock5_p & v8455e7;
assign v3a695c1 = hmaster1_p & v374729b | !hmaster1_p & v3a64b57;
assign v3735a25 = hgrant5_p & v3a5e684 | !hgrant5_p & v3a6fc61;
assign v374de7f = hburst0 & v376c211 | !hburst0 & v39ebb49;
assign v3a6bb65 = hbusreq5_p & v3a62b09 | !hbusreq5_p & v37654e7;
assign v373d4ff = hbusreq2_p & v3747302 | !hbusreq2_p & v3a6c5ee;
assign v3a706d1 = hbusreq1_p & v3a705e1 | !hbusreq1_p & v8455ab;
assign v3a57aad = hlock6_p & v376430b | !hlock6_p & v8455ab;
assign v3a56194 = hmaster3_p & v3722a42 | !hmaster3_p & v3a71125;
assign v3742cce = hbusreq7_p & v372f357 | !hbusreq7_p & v3764210;
assign v37798da = hmaster2_p & v3774bad | !hmaster2_p & a34d2b;
assign v2889705 = hbusreq2_p & v3a6c688 | !hbusreq2_p & v373125c;
assign v3a6f2bf = hgrant2_p & v3a6f718 | !hgrant2_p & v3a5d48f;
assign v375970d = hbusreq5 & v376256c | !hbusreq5 & v375e512;
assign v37506d8 = hgrant2_p & v3758472 | !hgrant2_p & v3767a5b;
assign v3a6f801 = hgrant6_p & v377097a | !hgrant6_p & v3a53c9d;
assign v3a6eaff = hgrant4_p & v8455ab | !hgrant4_p & v373bd6c;
assign v3736a37 = hbusreq1 & v3a6ab5f | !hbusreq1 & !v3748900;
assign v3a6931f = hmaster2_p & v373d825 | !hmaster2_p & v8455e7;
assign v37268b6 = hbusreq7_p & v3809e77 | !hbusreq7_p & v3a54e0c;
assign v3730a3d = hbusreq4_p & v3a70bc6 | !hbusreq4_p & v8455ab;
assign v373d687 = hbusreq8 & v3734a93 | !hbusreq8 & v3a6818c;
assign v3809f61 = hlock5_p & v37315af | !hlock5_p & v3a6fce0;
assign v3a5cae1 = hlock8_p & v3741920 | !hlock8_p & !v8455ab;
assign v375d7b6 = hgrant0_p & v3a70233 | !hgrant0_p & v376a8cf;
assign v3765406 = hgrant5_p & v8455ab | !hgrant5_p & v373127a;
assign v375921f = hmaster2_p & v8455ab | !hmaster2_p & !v373f503;
assign v3a70d59 = hlock8_p & v3740da1 | !hlock8_p & v8455ab;
assign v372c3e9 = hgrant7_p & v8455ab | !hgrant7_p & v3a6f49b;
assign v3735ea8 = hgrant6_p & v35b774b | !hgrant6_p & v374e9ac;
assign v375efe8 = hbusreq8_p & v372cf41 | !hbusreq8_p & !v8455ab;
assign v376c590 = hbusreq5_p & v3a6eec4 | !hbusreq5_p & v373e750;
assign v377e7f8 = jx1_p & v374cad6 | !jx1_p & v3744aca;
assign v3a594f1 = hgrant6_p & v374a664 | !hgrant6_p & v37506d8;
assign v374deab = hbusreq5 & v3729e17 | !hbusreq5 & v374949d;
assign v3a6fe15 = hbusreq8_p & v3769db7 | !hbusreq8_p & v3a6fb42;
assign v37388ce = hbusreq3_p & v375c939 | !hbusreq3_p & !v377b3a8;
assign v3a5e998 = hbusreq7 & v8455b0 | !hbusreq7 & v8455ab;
assign v3a59b8a = hbusreq0 & v3757adc | !hbusreq0 & v8455ab;
assign v3806542 = hmaster1_p & v37524b4 | !hmaster1_p & v3727ee9;
assign v3a62f75 = hmaster2_p & v3a5e2a3 | !hmaster2_p & v8455ab;
assign v3739fb8 = hbusreq5_p & v3a5fabd | !hbusreq5_p & v374e079;
assign v3737ce6 = hgrant3_p & v8455ab | !hgrant3_p & v372da87;
assign v3772962 = hmaster2_p & v3a712e2 | !hmaster2_p & v37711c3;
assign v3a63043 = hburst1 & v3745509 | !hburst1 & v374c862;
assign v3a709da = hmaster1_p & v3774a95 | !hmaster1_p & v373499c;
assign v372f3e0 = hbusreq4_p & v373330a | !hbusreq4_p & v3a6c515;
assign v3761224 = hbusreq1_p & v37c011c | !hbusreq1_p & !v8455ab;
assign v37c038c = hbusreq6_p & v3a7145f | !hbusreq6_p & v3a6b688;
assign v3749b62 = hbusreq4 & v37290af | !hbusreq4 & v8455ab;
assign v3a6fc53 = hgrant1_p & v3735593 | !hgrant1_p & v3743690;
assign v373c07d = hgrant4_p & v375413c | !hgrant4_p & v88c50b;
assign v3779c7e = hmaster2_p & v3a6e7b3 | !hmaster2_p & !v8455ab;
assign v3751f34 = hbusreq4_p & v3a709e2 | !hbusreq4_p & v37388ce;
assign v376605a = hbusreq0_p & v372b351 | !hbusreq0_p & v8455b6;
assign v3765d9e = hmaster1_p & v372f309 | !hmaster1_p & v3a6f3fa;
assign v39a5359 = hgrant5_p & v377e319 | !hgrant5_p & v3779852;
assign v3a5610f = hbusreq3_p & v3a56e5e | !hbusreq3_p & v38072fd;
assign v373f27d = hbusreq5_p & v3a61f83 | !hbusreq5_p & !v376b012;
assign v374c88a = hbusreq0 & v37476f7 | !hbusreq0 & v376a1a3;
assign v3741357 = hmaster2_p & v33781df | !hmaster2_p & v374220d;
assign v376a31b = hgrant4_p & v3779060 | !hgrant4_p & v377c7ce;
assign v37634d8 = hgrant4_p & v8455ab | !hgrant4_p & v376ebe6;
assign v3770366 = hmaster0_p & v374184c | !hmaster0_p & v3a669e9;
assign v377b3df = hmaster0_p & v3a6d499 | !hmaster0_p & v3a70716;
assign v37309ae = hmaster1_p & v35b7168 | !hmaster1_p & v3a656b2;
assign v37580b6 = jx3_p & v3742f1b | !jx3_p & v360cd91;
assign v3758c62 = hgrant0_p & v8455ab | !hgrant0_p & v37703c6;
assign v3a6f522 = hbusreq0_p & v377606f | !hbusreq0_p & v8455b5;
assign v3a7128e = hmaster2_p & v8455ab | !hmaster2_p & v3a6422d;
assign v377ef47 = hbusreq2_p & v3748ca5 | !hbusreq2_p & v376ba33;
assign v3a70931 = jx0_p & v2ff8e61 | !jx0_p & v3774d13;
assign v3a6ceb0 = hbusreq5_p & v3742649 | !hbusreq5_p & v375c740;
assign v3a70d94 = hbusreq0 & v3a63d63 | !hbusreq0 & v3777e69;
assign v373dd4a = hlock0 & v3a70244 | !hlock0 & d5ffe1;
assign v3752798 = hmaster0_p & a747d7 | !hmaster0_p & v3a6e96b;
assign v37425ad = hgrant6_p & v37658d7 | !hgrant6_p & v3a70986;
assign v3a6f160 = hlock4 & v373a5a6 | !hlock4 & v372bf7f;
assign v3a70a2b = hmaster2_p & v3736ded | !hmaster2_p & v8455ab;
assign v3a70ebc = hmaster0_p & v375fa16 | !hmaster0_p & !v37243fe;
assign v377b7f9 = hlock4 & v3775c0b | !hlock4 & v377f73c;
assign v3a63f06 = hgrant6_p & v8455ab | !hgrant6_p & v3759d52;
assign v3758174 = hmaster2_p & v3a578e2 | !hmaster2_p & v3a685e1;
assign v3a70795 = hlock8 & v3774664 | !hlock8 & v3a62dae;
assign v3a5f0a7 = hbusreq3_p & v3751161 | !hbusreq3_p & v8455ab;
assign v377492b = hbusreq4 & v376d1e2 | !hbusreq4 & v3a69487;
assign v3735ac3 = hmaster2_p & b0c091 | !hmaster2_p & v8455e7;
assign v3a68399 = hbusreq5 & v3a697d2 | !hbusreq5 & v373d68a;
assign v3a63938 = hbusreq0 & v372cb28 | !hbusreq0 & !v8455ab;
assign v3a71006 = hbusreq2_p & v3a68016 | !hbusreq2_p & v373e98b;
assign v376d972 = hlock8 & v376366a | !hlock8 & v3a6022f;
assign v3a5e5f3 = hbusreq4 & v3729004 | !hbusreq4 & v8455ab;
assign v3777996 = hbusreq6_p & v3a7125f | !hbusreq6_p & v37387ed;
assign v3775684 = hgrant4_p & v37386fb | !hgrant4_p & v2092aaa;
assign v376e0cb = hbusreq8_p & v373293c | !hbusreq8_p & v1e3737f;
assign v3760e51 = hmaster2_p & v3a57f59 | !hmaster2_p & v3759032;
assign v373d2e3 = hmaster0_p & v3a711ec | !hmaster0_p & v8455ab;
assign v372b1b5 = hmaster2_p & v3770415 | !hmaster2_p & v376a96b;
assign v37402cd = hbusreq4_p & v38072fd | !hbusreq4_p & v372cb99;
assign v3a55fe8 = hlock7 & v376d0b5 | !hlock7 & v3766f51;
assign v37361e7 = hbusreq6_p & v3731c79 | !hbusreq6_p & !v8455ab;
assign v37418dc = hmaster2_p & v374bb76 | !hmaster2_p & v37320ff;
assign v3723e1f = hlock2 & v3a6f613 | !hlock2 & v372b7b7;
assign v3727e66 = hgrant4_p & v3a63a7a | !hgrant4_p & v3758850;
assign hmaster0 = !v28e9804;
assign v377757b = hbusreq6 & v37366d0 | !hbusreq6 & v8455ab;
assign v3a670fb = hmaster0_p & v3a6d1aa | !hmaster0_p & v373a3c8;
assign v372c921 = hbusreq7_p & v377e568 | !hbusreq7_p & v372f765;
assign v373eeec = hbusreq7 & v87762a | !hbusreq7 & v377b774;
assign a4764c = hgrant4_p & v375641f | !hgrant4_p & v922c1b;
assign v375dc25 = hmaster1_p & v3a61532 | !hmaster1_p & v3a573c2;
assign v3a70214 = hbusreq6 & v376111d | !hbusreq6 & v8455ab;
assign v380714f = hmaster2_p & v8455ab | !hmaster2_p & !v375aaca;
assign v3a55349 = hgrant2_p & v8455ab | !hgrant2_p & v3742d37;
assign v3722e5e = hbusreq4 & v3a5fd6a | !hbusreq4 & v3737028;
assign v37531fd = hbusreq5 & v37730ff | !hbusreq5 & v37371df;
assign v37613d3 = hbusreq6_p & v374c33a | !hbusreq6_p & v373a2f2;
assign v3747006 = hmaster0_p & v3762557 | !hmaster0_p & v376730a;
assign v3a68aa8 = hbusreq3_p & v3a6e47f | !hbusreq3_p & v3a6c355;
assign v3a715d9 = hmaster0_p & v375607f | !hmaster0_p & v37696c4;
assign v373a333 = hbusreq6_p & v3a635ea | !hbusreq6_p & v377aeba;
assign v37518fb = hbusreq6 & v3773d82 | !hbusreq6 & v8455b0;
assign v3a6fca7 = jx3_p & v375e34d | !jx3_p & v372c3e9;
assign v3762847 = hlock5_p & v375dda4 | !hlock5_p & v8455ab;
assign v3a54a76 = hgrant3_p & v376ace9 | !hgrant3_p & v373b197;
assign v375e4d9 = jx0_p & v3a70175 | !jx0_p & v3766846;
assign v37411c1 = hmaster1_p & v37640dc | !hmaster1_p & v372e1bb;
assign v37742a4 = hmaster0_p & v37539cd | !hmaster0_p & !v3a658cf;
assign v375178f = hbusreq6 & v376bf0a | !hbusreq6 & v8455ab;
assign v3748451 = hgrant4_p & v375bde1 | !hgrant4_p & v3741c76;
assign v3743fea = hgrant5_p & v373ae84 | !hgrant5_p & v3754eca;
assign c75852 = hbusreq3 & v3a70a8a | !hbusreq3 & v8455ab;
assign v3a70221 = hbusreq5_p & v3a62542 | !hbusreq5_p & v377accc;
assign cf8423 = hlock5 & v3754ce8 | !hlock5 & v38097c0;
assign v3a55ec0 = hbusreq7_p & v3a5a4ce | !hbusreq7_p & v8455ab;
assign v3a71302 = hgrant2_p & v374d542 | !hgrant2_p & v3a6eab3;
assign v3a62c28 = hmaster1_p & v3771ce8 | !hmaster1_p & v3736358;
assign v3723d1a = hgrant5_p & v8455ab | !hgrant5_p & v376a847;
assign v3a5c3d3 = hmaster2_p & v373133d | !hmaster2_p & v375b7bd;
assign v372e1bb = hbusreq5_p & v373d957 | !hbusreq5_p & v3a6ea2b;
assign af345a = hbusreq8_p & v376a3cb | !hbusreq8_p & v3a65b64;
assign v377d367 = hbusreq4_p & v3724731 | !hbusreq4_p & v3735c9d;
assign v3a71288 = hmaster2_p & v3a5b289 | !hmaster2_p & v3767561;
assign v3a709df = hbusreq2_p & v3a6a831 | !hbusreq2_p & v3725092;
assign v3754fc8 = hbusreq0 & v375c423 | !hbusreq0 & v8455ab;
assign v380761d = hgrant6_p & v3742c16 | !hgrant6_p & v2aca977;
assign v377a43e = hgrant3_p & v360d0db | !hgrant3_p & v3729115;
assign v3a6f733 = hmaster1_p & v3a5c3a0 | !hmaster1_p & v3a707e0;
assign v3732688 = hbusreq5 & v374558a | !hbusreq5 & v8455ab;
assign v3a702b0 = hbusreq4 & v3a6f5fb | !hbusreq4 & v8455ab;
assign v3a6cfa7 = hburst0 & v373bf7c | !hburst0 & v372dd8e;
assign v3744adf = hbusreq6 & v374401a | !hbusreq6 & v376bade;
assign v3a5a158 = hbusreq3_p & v37591b4 | !hbusreq3_p & v8455ab;
assign v375214d = hmaster2_p & v8455e1 | !hmaster2_p & !v8455ab;
assign v375e7cc = hbusreq2_p & v377af0a | !hbusreq2_p & !v377408e;
assign v3a71146 = hmaster1_p & v3a635ea | !hmaster1_p & v3a5e783;
assign v3748eff = hmaster1_p & v3a65aa5 | !hmaster1_p & v3747fd2;
assign v3763e6c = hmaster3_p & v3a5a814 | !hmaster3_p & v3734a96;
assign v374fac7 = hmaster2_p & v3747302 | !hmaster2_p & v3a57959;
assign v3a6741a = hgrant3_p & v376f768 | !hgrant3_p & ca602f;
assign v3734b97 = hbusreq4_p & v3a60787 | !hbusreq4_p & !v377cfd9;
assign v376c028 = hlock5 & v372494a | !hlock5 & v3763f13;
assign v3a63d7a = hbusreq2 & v374e35e | !hbusreq2 & v8455ab;
assign v3728fe7 = hbusreq4 & v3a5f642 | !hbusreq4 & v8455ab;
assign v3a6f31d = hmaster1_p & v37249c7 | !hmaster1_p & !v377167d;
assign v3a6fe6a = hburst1 & v3757c6f | !hburst1 & v3777a7f;
assign v3a6dcbf = hbusreq7 & v3a5bc27 | !hbusreq7 & v3758435;
assign v3a6ff23 = hbusreq4_p & v374e28d | !hbusreq4_p & v8455ab;
assign v3762116 = hgrant5_p & v3a6d3b6 | !hgrant5_p & v37306ec;
assign v374ace7 = hgrant0_p & v3a714f5 | !hgrant0_p & v374059d;
assign v3730d64 = hbusreq5 & v3a7130b | !hbusreq5 & v3a58c07;
assign v3a6f8ce = jx0_p & v375c358 | !jx0_p & v3a63dde;
assign v3a61fc9 = hlock1_p & v3750d37 | !hlock1_p & !v8455ab;
assign v3727420 = hbusreq0 & v3778cdb | !hbusreq0 & v3747193;
assign v3a57836 = hbusreq3_p & v37581c0 | !hbusreq3_p & v8455b0;
assign v374500f = hgrant2_p & v375975b | !hgrant2_p & v373913a;
assign v3742dce = hbusreq0 & v376a348 | !hbusreq0 & v374b30b;
assign v3a5cdf4 = hbusreq5_p & v3a57db6 | !hbusreq5_p & v375a64f;
assign v375de72 = hbusreq8_p & v3a6fdce | !hbusreq8_p & v3726f76;
assign v377af64 = hbusreq0_p & v3a5b563 | !hbusreq0_p & v372998c;
assign v3a708e7 = hmaster2_p & v3775f1f | !hmaster2_p & v3754d3a;
assign v375b56c = hmaster1_p & v3a635ea | !hmaster1_p & v3809964;
assign v37660d2 = hbusreq3_p & v3a635ea | !hbusreq3_p & v3a70eb6;
assign v37327c3 = hbusreq5 & v3761b24 | !hbusreq5 & v373d964;
assign v377d2a0 = hgrant4_p & v3751d73 | !hgrant4_p & v3a64e40;
assign v37571c0 = hgrant4_p & v372b77b | !hgrant4_p & v3a6aaaa;
assign v374586a = hbusreq4_p & v373d7f9 | !hbusreq4_p & v374877e;
assign bdb49d = hbusreq3_p & v3752ec0 | !hbusreq3_p & v3724d93;
assign v3733998 = hbusreq8 & v3740cd2 | !hbusreq8 & v3a5bb57;
assign v3739c6f = hbusreq5_p & v3a6f9d3 | !hbusreq5_p & v3a708c9;
assign v3a6d558 = hbusreq4 & v3747b3c | !hbusreq4 & v3a5f9e6;
assign v37408a3 = hbusreq3 & v37416b5 | !hbusreq3 & v37496fa;
assign v376e844 = hbusreq4_p & v372b2ab | !hbusreq4_p & v3739e25;
assign v37765fb = hgrant2_p & v3a5872b | !hgrant2_p & v3751f67;
assign v3a700ec = hbusreq2_p & v3a6c40f | !hbusreq2_p & !v3a68591;
assign v375c0cd = hgrant2_p & v8455ab | !hgrant2_p & v376fb18;
assign v3741bce = hmaster2_p & v3a7015f | !hmaster2_p & v8455ab;
assign v37532ac = hgrant6_p & v3a2a8f2 | !hgrant6_p & d78807;
assign v3a6f96f = hbusreq2 & v3a5600a | !hbusreq2 & v375444e;
assign v372ed88 = hgrant6_p & v37361e7 | !hgrant6_p & !v8455ab;
assign v375c317 = hbusreq4 & v373933b | !hbusreq4 & v8455ab;
assign v372fa9d = hbusreq5 & v3a70ca5 | !hbusreq5 & v377a2f3;
assign v1e37bab = hbusreq3 & v3754ec1 | !hbusreq3 & !v3a6fe1a;
assign v3a625ac = hmaster0_p & v8455ab | !hmaster0_p & v373a0ea;
assign v373796a = hmaster0_p & v37430c6 | !hmaster0_p & v3a6fe4d;
assign v3747167 = hbusreq6 & v37282cf | !hbusreq6 & v37674c1;
assign v376e1fd = hmaster0_p & v3a64421 | !hmaster0_p & v3a6c6ce;
assign v3744ae4 = hbusreq4 & v3a5408c | !hbusreq4 & v3762502;
assign v3761af1 = hgrant0_p & v8455ab | !hgrant0_p & v3a6b18a;
assign v3a55377 = hmaster2_p & v376bca9 | !hmaster2_p & v373b02e;
assign v3752616 = hbusreq5_p & v3a635ea | !hbusreq5_p & v37c36bf;
assign v3770f97 = hmaster1_p & v375a1a7 | !hmaster1_p & v373e27e;
assign v3a70a05 = hgrant2_p & v3a5f50e | !hgrant2_p & v35b70e6;
assign v374cf82 = hbusreq5 & v372bfd0 | !hbusreq5 & v374514e;
assign v3754eb4 = hmaster1_p & v37281ca | !hmaster1_p & v3a6a73a;
assign v373bc2f = hmaster0_p & v3770ff4 | !hmaster0_p & v3a70ede;
assign v372b721 = hlock7 & a0a219 | !hlock7 & v377ebf3;
assign v3742146 = hmaster1_p & v3a5e24e | !hmaster1_p & v376e074;
assign v37278f5 = hbusreq5 & v3a70ff7 | !hbusreq5 & v8455ab;
assign v37530c7 = hbusreq5 & v3724b74 | !hbusreq5 & v3a59de6;
assign v37761e4 = stateG10_1_p & v35772a6 | !stateG10_1_p & !v377217f;
assign v374bae0 = hbusreq0_p & v35772a5 | !hbusreq0_p & !v3806507;
assign v372c1b0 = hbusreq4 & v3728ea7 | !hbusreq4 & v3759361;
assign v3746f18 = jx0_p & v3759d9c | !jx0_p & v3a6f223;
assign v376ad8c = hbusreq5_p & v37661dc | !hbusreq5_p & !v375e167;
assign v3766452 = hgrant1_p & v3759032 | !hgrant1_p & !v39a537f;
assign v3a66492 = hlock0_p & v377eaf2 | !hlock0_p & v3a6946d;
assign v3a6f880 = hgrant2_p & v3771656 | !hgrant2_p & v3a6f918;
assign v3763055 = hmaster2_p & v3a57584 | !hmaster2_p & v3a6f32f;
assign v9ca2d6 = hlock5 & v3a6d686 | !hlock5 & v3736113;
assign v3a6b6f3 = hbusreq1_p & v2aca977 | !hbusreq1_p & v372b819;
assign v23fde92 = hbusreq2 & v376d1e2 | !hbusreq2 & v3a69487;
assign v375b84e = hgrant5_p & v8455ab | !hgrant5_p & v377ba29;
assign v3a6fcc9 = hmaster0_p & v3a70d3e | !hmaster0_p & v3722ae9;
assign a9e394 = hmaster2_p & v3735afb | !hmaster2_p & v8455b3;
assign v3a70c72 = hbusreq0 & v3a6d840 | !hbusreq0 & v372f76c;
assign v3809390 = hmaster0_p & v8455ab | !hmaster0_p & v374d847;
assign v3a697b9 = hbusreq5_p & v3735324 | !hbusreq5_p & v373b11a;
assign v3a5902f = hmaster2_p & v3a716a0 | !hmaster2_p & v3730a3d;
assign v3a6616c = hbusreq4_p & v3a714fc | !hbusreq4_p & v8455b0;
assign v3a5d186 = hmaster1_p & v3a70377 | !hmaster1_p & v3728d9c;
assign v3743f5a = hbusreq6_p & v37586c0 | !hbusreq6_p & v8455ab;
assign v372433d = hbusreq4_p & v8455b7 | !hbusreq4_p & v37759b6;
assign v374aa73 = stateA1_p & v20d166d | !stateA1_p & v374ceec;
assign v376c569 = hbusreq2 & v3749435 | !hbusreq2 & v8455ab;
assign v3a6fcb2 = hmaster0_p & v8455e7 | !hmaster0_p & v373e13a;
assign v3a703a7 = hmaster0_p & v8455e7 | !hmaster0_p & v372e466;
assign v3726b63 = hbusreq8_p & v3a7104f | !hbusreq8_p & v3a711c3;
assign v3766eef = hbusreq2_p & v8455ab | !hbusreq2_p & v37758ce;
assign v3a64b0f = hbusreq4 & v372e244 | !hbusreq4 & v374d0e3;
assign v3a6fd5d = hmaster1_p & v3a6dfb2 | !hmaster1_p & v376075c;
assign v37307d7 = hbusreq0 & v3a6ef2e | !hbusreq0 & v1e37cd6;
assign v3a6f616 = hgrant6_p & v376a040 | !hgrant6_p & !v3725786;
assign v3a5ae2f = hbusreq1_p & v3a70334 | !hbusreq1_p & v3a6ec94;
assign v3a6da08 = hmaster1_p & v3a58ddb | !hmaster1_p & v3a6f790;
assign v325c974 = hmaster1_p & v3753a34 | !hmaster1_p & v375b389;
assign v377b292 = hbusreq3 & v3a70321 | !hbusreq3 & v375cf36;
assign v3a6ac2c = hmaster1_p & v373f7ef | !hmaster1_p & !v3a6a33a;
assign v3774df5 = hbusreq5 & v375f368 | !hbusreq5 & !v3a60301;
assign v3a70666 = hmaster2_p & v8907fb | !hmaster2_p & v373b5d8;
assign v3727e25 = hmaster1_p & v37660f0 | !hmaster1_p & v8455ab;
assign v37483c5 = hgrant6_p & v3a5a63c | !hgrant6_p & v376e4da;
assign v375067d = hmaster0_p & v3a6dc08 | !hmaster0_p & v3a5f495;
assign v3762cb2 = hmaster2_p & v8455ab | !hmaster2_p & !v3a6419e;
assign v373fe1f = hmaster2_p & v3a66aa4 | !hmaster2_p & v373997b;
assign v3a53cf5 = hbusreq4 & v3a697f1 | !hbusreq4 & !v3731c4b;
assign a6859a = hbusreq6_p & v3770dcb | !hbusreq6_p & v374f630;
assign v380693e = hbusreq1 & v3743b9e | !hbusreq1 & v37496fa;
assign v374731f = hmaster1_p & v377007d | !hmaster1_p & v375918d;
assign v372456f = hgrant1_p & v3730e71 | !hgrant1_p & v373df21;
assign v373cdef = hmaster3_p & v372c30a | !hmaster3_p & v3725eb6;
assign v37582e0 = hlock7 & v3a5de5f | !hlock7 & v374b19b;
assign v377f108 = start_p & v845605 | !start_p & v8455ab;
assign v374523d = hmaster2_p & v3757b9b | !hmaster2_p & v3a6ef89;
assign v9450a2 = hbusreq6 & v374a134 | !hbusreq6 & v8455ab;
assign v3765463 = hbusreq5 & v3a5dad5 | !hbusreq5 & v373de86;
assign v3726df4 = hbusreq1_p & v35b9d52 | !hbusreq1_p & v2acb0c1;
assign v3a5cf22 = hgrant2_p & v374068b | !hgrant2_p & v3766d0d;
assign v3774d15 = hgrant6_p & v373ba4a | !hgrant6_p & v3731a29;
assign v3a68e39 = hgrant3_p & v3775aea | !hgrant3_p & v373687f;
assign v374e74c = hmaster1_p & v3a63ea7 | !hmaster1_p & v3a54264;
assign v37759e3 = hbusreq0 & v3a6fb51 | !hbusreq0 & v8455ab;
assign v3730617 = jx0_p & v374fd1f | !jx0_p & v8455ab;
assign v377408e = hbusreq2 & v374cab9 | !hbusreq2 & v37674c1;
assign v377dae3 = hgrant6_p & v3a62a6d | !hgrant6_p & v3a711dd;
assign v3779f43 = hbusreq0 & v3764bd6 | !hbusreq0 & v37285eb;
assign v3a712ae = hbusreq8_p & v2acaeaa | !hbusreq8_p & v3745b51;
assign v3a6be05 = hbusreq5 & v3a6f740 | !hbusreq5 & v373f06c;
assign v372d10e = hgrant6_p & v8455ab | !hgrant6_p & v2ff8e00;
assign v37243e6 = hbusreq6 & v3a705ad | !hbusreq6 & v964c47;
assign v8455b9 = hbusreq2_p & v8455ab | !hbusreq2_p & !v8455ab;
assign v3806c04 = hgrant5_p & v8455ab | !hgrant5_p & v374069b;
assign v3a6ff32 = hbusreq6_p & v37728a5 | !hbusreq6_p & v3a70d99;
assign v377dbd7 = hmaster2_p & v3779183 | !hmaster2_p & v375f2ba;
assign v3766e3a = hbusreq1_p & v377c2ba | !hbusreq1_p & !v3752648;
assign v372d827 = hgrant5_p & v3769559 | !hgrant5_p & v3809e3c;
assign v35b779e = hmaster0_p & v8455ab | !hmaster0_p & v377d945;
assign v373484e = hgrant6_p & v3735525 | !hgrant6_p & v3739da7;
assign v3a69671 = hbusreq3 & v37274c2 | !hbusreq3 & !v8455b5;
assign v3756c22 = hmaster1_p & v375a4d0 | !hmaster1_p & v3770b26;
assign v372f260 = hmaster2_p & v3a71162 | !hmaster2_p & v372a85f;
assign v377115d = hmaster0_p & v3a6f62b | !hmaster0_p & v374e855;
assign v3a70c8c = hgrant4_p & v3a6f585 | !hgrant4_p & v3a6e0f4;
assign v3725994 = hbusreq3 & v3753dab | !hbusreq3 & v8455ab;
assign v376888c = hgrant4_p & v372abd8 | !hgrant4_p & v37765d0;
assign v3a7044e = hbusreq8 & v3746ed6 | !hbusreq8 & v376b3d4;
assign v37507dd = hlock4 & v1e379ef | !hlock4 & v377a5a9;
assign v3750e94 = hbusreq4 & v3a6f018 | !hbusreq4 & !v3a5db8a;
assign v3757c10 = hlock4 & v372cfd2 | !hlock4 & v3769e3a;
assign v3a7142e = hmaster1_p & v3757568 | !hmaster1_p & v3a5d431;
assign v37410bd = hmaster0_p & v3a70b71 | !hmaster0_p & v3a70574;
assign v3744cf7 = hmaster1_p & v37245f8 | !hmaster1_p & v3a700c6;
assign v3a5fbad = hgrant6_p & v374cb44 | !hgrant6_p & !v3764114;
assign v376d82f = hbusreq2_p & v375a235 | !hbusreq2_p & v375d30b;
assign v37562f2 = hgrant3_p & v37761ae | !hgrant3_p & !v3a5c904;
assign v377629f = hlock6 & v375d4d9 | !hlock6 & v374d8bb;
assign v37484df = hbusreq2_p & v374cab9 | !hbusreq2_p & c61447;
assign v3a6eec9 = hbusreq0 & v2678c95 | !hbusreq0 & v3767258;
assign v3767b77 = hgrant5_p & v3a7150f | !hgrant5_p & v374e4bd;
assign v3749e96 = hgrant6_p & v8455ab | !hgrant6_p & v376ed1f;
assign v377704c = hgrant6_p & v3a635ea | !hgrant6_p & v3750f72;
assign v3737554 = busreq_p & v373deb5 | !busreq_p & v3748422;
assign v3a6947c = hmaster1_p & v37744a3 | !hmaster1_p & v3a59de6;
assign v3728b05 = hgrant0_p & v37301f5 | !hgrant0_p & v376ef3f;
assign v376f0c3 = hgrant7_p & v8455ab | !hgrant7_p & v372bb4b;
assign v3a70f53 = hgrant4_p & v377c931 | !hgrant4_p & v3753030;
assign v3764f6a = hgrant5_p & v37378d4 | !hgrant5_p & v3806542;
assign v3a6b27e = hmaster2_p & v377e784 | !hmaster2_p & v3a637dd;
assign v3754ec1 = hbusreq1_p & v3a540f3 | !hbusreq1_p & v8455ab;
assign v3773043 = hbusreq2 & v3a5eafa | !hbusreq2 & v375cf36;
assign v3a62079 = hmaster2_p & v3a70987 | !hmaster2_p & v3739d88;
assign v377fb84 = hbusreq2 & v3747994 | !hbusreq2 & v8455ab;
assign v39a53eb = hmaster0_p & v37356f0 | !hmaster0_p & v3a670e4;
assign v3a62f06 = hlock4 & v38072fd | !hlock4 & v375ff0d;
assign v3762ca2 = hbusreq5_p & v3a5c3eb | !hbusreq5_p & v377b3df;
assign v374d0f9 = hlock6 & v3758f1b | !hlock6 & v3756c25;
assign v3765f13 = hlock4 & v3733690 | !hlock4 & v377c214;
assign v3763311 = hbusreq7 & v376e822 | !hbusreq7 & v3a63368;
assign v3768751 = hgrant6_p & v3a6f3c6 | !hgrant6_p & v37533ea;
assign v3a70b43 = hlock7_p & v3752781 | !hlock7_p & v37572b6;
assign v37379fc = hbusreq6_p & v375306b | !hbusreq6_p & v8455b7;
assign v3a70cd0 = jx0_p & v373bb89 | !jx0_p & v374de47;
assign v3a70e60 = hbusreq4 & v375b9a0 | !hbusreq4 & v3a64af7;
assign v376f7ab = hgrant2_p & v8455ab | !hgrant2_p & v3752b4b;
assign v3773b23 = hready & v3726dfa | !hready & !v375e373;
assign v374221c = hbusreq5_p & v37384a9 | !hbusreq5_p & v3a70b4b;
assign v3a5c5e5 = hmaster2_p & v3757966 | !hmaster2_p & v3776196;
assign v372834c = hgrant3_p & v372ad53 | !hgrant3_p & v373dfcc;
assign v3a6fe5d = hgrant3_p & v3a56aeb | !hgrant3_p & v3772dc6;
assign v3a709fc = hmaster0_p & v3a71133 | !hmaster0_p & !v3807765;
assign v3a6ac60 = hgrant2_p & v37646c7 | !hgrant2_p & v3748ca5;
assign v3a6c4c3 = hbusreq5 & v3758bc2 | !hbusreq5 & v1e37405;
assign v3a71601 = hgrant4_p & v3a6ef50 | !hgrant4_p & !v3809d87;
assign v3736913 = hbusreq2 & v3806db7 | !hbusreq2 & v374f87c;
assign v377e1e8 = hbusreq2_p & v3765901 | !hbusreq2_p & v3a709aa;
assign v3775a7d = hgrant2_p & v8455ab | !hgrant2_p & v377d7e1;
assign v37c028d = hbusreq8 & v3a68057 | !hbusreq8 & v3a6194e;
assign v373ef10 = hbusreq5_p & v3a6eb22 | !hbusreq5_p & v3744898;
assign v3a6feb4 = hmaster0_p & v3745ece | !hmaster0_p & v3745b9c;
assign v3737d95 = hgrant6_p & v3a70a41 | !hgrant6_p & v3a6f5d1;
assign v375cf7d = hbusreq6 & v3738d0b | !hbusreq6 & v3a70f74;
assign v3a67983 = hready & v8455ab | !hready & !v373dceb;
assign v1e37b76 = hmaster0_p & v3a6fd72 | !hmaster0_p & v3735272;
assign v3749975 = hbusreq7 & v372a636 | !hbusreq7 & v374dc1b;
assign v375eefe = hmaster0_p & v374bf36 | !hmaster0_p & v377f34a;
assign v3a6e031 = hlock5_p & v3725198 | !hlock5_p & v3a5b289;
assign v3729031 = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3738d63;
assign v3a708b6 = hmaster1_p & v3748451 | !hmaster1_p & v3a68c7d;
assign v3a709ef = hbusreq0_p & v3747302 | !hbusreq0_p & v3743b9e;
assign v3728cfe = hgrant3_p & v3a5978c | !hgrant3_p & v8455ab;
assign v3a6842c = hmaster2_p & v8455e7 | !hmaster2_p & v3723430;
assign v3a5d3fc = hbusreq5 & v3753bfb | !hbusreq5 & v3a6f462;
assign v37386cb = hlock4_p & v3a6fa39 | !hlock4_p & !v8455ab;
assign v3a70daf = hmaster1_p & v8455ab | !hmaster1_p & !v3a6fac3;
assign v377a522 = hmaster1_p & v3779060 | !hmaster1_p & v3a5cb4c;
assign v3a70145 = hlock5_p & v3734967 | !hlock5_p & !v3768de8;
assign v39ebacc = hbusreq5 & v377f64b | !hbusreq5 & v8455ab;
assign v3a6f598 = hlock3_p & v375b902 | !hlock3_p & !v3a6ac26;
assign v376ec1d = hbusreq7_p & v3a69c7b | !hbusreq7_p & v8455ab;
assign v3726d4a = hmaster1_p & v375c381 | !hmaster1_p & v376d215;
assign v39a5420 = hbusreq4 & v373a972 | !hbusreq4 & v3a6faef;
assign v3a5e8a1 = hmaster2_p & v3757568 | !hmaster2_p & !v3732dc6;
assign v3a6f213 = hbusreq1_p & v375ff95 | !hbusreq1_p & v8455ab;
assign v3a6f10f = hbusreq1 & v3a6ffca | !hbusreq1 & v8455ab;
assign v374445b = hgrant5_p & v8455ab | !hgrant5_p & v3a6a093;
assign v3a71561 = hmaster2_p & v8455ab | !hmaster2_p & !v373f2d8;
assign v376e04c = hbusreq2_p & v3778fec | !hbusreq2_p & v3a5bb64;
assign v3a6e552 = hgrant5_p & v373c5ea | !hgrant5_p & v3a70d23;
assign v377c147 = hbusreq6_p & v3a70ed6 | !hbusreq6_p & v37642f9;
assign v3903ee6 = hready_p & v3a70400 | !hready_p & b15d44;
assign v3a58967 = hmaster0_p & v3a709ed | !hmaster0_p & v376d07b;
assign v372dc8e = hmaster0_p & v8455ab | !hmaster0_p & v3a58519;
assign v376819e = hbusreq0 & v372e88f | !hbusreq0 & v3724859;
assign v3a64fe0 = hbusreq3 & v3733ea2 | !hbusreq3 & !v8455ab;
assign v375a261 = hbusreq4 & v372ea4b | !hbusreq4 & v3a70a88;
assign v3a71688 = hgrant0_p & v37773a9 | !hgrant0_p & v3a60bc8;
assign v376eef5 = hmaster1_p & v3a70db1 | !hmaster1_p & v3a60e4c;
assign v3756d57 = hbusreq5 & v3a6396b | !hbusreq5 & v8455ab;
assign v3a6f56a = hmaster2_p & v3a5a807 | !hmaster2_p & !v374f547;
assign v372b3cf = stateA1_p & v373f4d3 | !stateA1_p & v3a6ffe0;
assign v3a6ab55 = hmaster0_p & v3748451 | !hmaster0_p & v372a246;
assign v37741ca = hbusreq0 & v3774d15 | !hbusreq0 & v3a70190;
assign v3a71332 = hmaster0_p & v3734534 | !hmaster0_p & v8d4314;
assign v372ec78 = hbusreq0 & v3a6f5fb | !hbusreq0 & v8455ab;
assign v3a634fa = hlock7_p & v3a6f2be | !hlock7_p & !v3768d7e;
assign v3775653 = hbusreq2_p & v376f56d | !hbusreq2_p & v3a54c8d;
assign v376f8ba = hmaster2_p & v3a703c3 | !hmaster2_p & !v3739ddf;
assign v3a714b0 = hmaster1_p & v3727d4c | !hmaster1_p & v374c000;
assign v37571a9 = hbusreq3_p & v372f391 | !hbusreq3_p & v8455b0;
assign v37366d5 = hmaster0_p & v3763c39 | !hmaster0_p & v8455ab;
assign v3a555a9 = hbusreq7 & v3a6f474 | !hbusreq7 & v377386a;
assign v373c9b1 = hbusreq2 & v3a6f4ac | !hbusreq2 & v374acbe;
assign v37493ce = start_p & v8455d5 | !start_p & v3a712be;
assign v3a53c21 = hbusreq6_p & v374bec6 | !hbusreq6_p & v3750c47;
assign v3a70736 = hmaster0_p & v3807aa1 | !hmaster0_p & v374cdc4;
assign v3a299ba = hbusreq8 & v375ef7b | !hbusreq8 & v375e8d2;
assign v3a643d6 = hbusreq7 & v375580b | !hbusreq7 & cb85ef;
assign v3a70ec3 = hbusreq3_p & v377094b | !hbusreq3_p & v3a71422;
assign v3a6f2d1 = hbusreq0 & v3729030 | !hbusreq0 & v3727ed2;
assign v3a5a039 = hmaster2_p & v3763a86 | !hmaster2_p & v377bbd9;
assign v3a7160a = hmaster1_p & v3a5b8b9 | !hmaster1_p & v3778aa0;
assign v3751de0 = hlock5_p & v3743613 | !hlock5_p & v3a6f86b;
assign v3a70771 = hmaster2_p & v377b946 | !hmaster2_p & v3a6f3c6;
assign v376a054 = jx0_p & v3a5c484 | !jx0_p & v374beb6;
assign v3a5e1e8 = hmaster2_p & v377adf5 | !hmaster2_p & v374c7f4;
assign v3a7088f = hbusreq4 & d44200 | !hbusreq4 & v8455ab;
assign v3770bcd = hgrant4_p & v376a6f1 | !hgrant4_p & v374950c;
assign v3742f7f = hmaster3_p & v3750382 | !hmaster3_p & v8455ab;
assign v3724872 = hmaster1_p & v3a70e2f | !hmaster1_p & v3a5ce55;
assign v39a53e9 = hmaster0_p & v3759519 | !hmaster0_p & v373d67c;
assign v3a60ce2 = decide_p & v3a70b11 | !decide_p & v3a69c73;
assign v3a6439a = hbusreq4 & v377dae3 | !hbusreq4 & v3750c52;
assign v3a70d2c = hbusreq2 & v3a696ed | !hbusreq2 & v8455ab;
assign v3a70854 = hbusreq5 & v3755f9d | !hbusreq5 & v377de7f;
assign v3a56ba2 = hmaster0_p & v3771076 | !hmaster0_p & v3768070;
assign v3a5c4b0 = hgrant5_p & v8455c6 | !hgrant5_p & v3732e48;
assign v3753a34 = hlock5 & v374cef4 | !hlock5 & v1e37397;
assign v3a5d8e0 = hmaster1_p & v3752fcb | !hmaster1_p & v3a70cc7;
assign v3733440 = hgrant4_p & v3a7129f | !hgrant4_p & v376c26e;
assign v3a6c066 = hbusreq6 & v3a58218 | !hbusreq6 & v8455ab;
assign v3a6f08d = hbusreq5 & v3763f30 | !hbusreq5 & !v8455b5;
assign v3770ff9 = hmaster0_p & v3a5fc34 | !hmaster0_p & v3746b73;
assign v372b9c5 = hmaster0_p & v3a70f68 | !hmaster0_p & v37565b0;
assign v3775b2f = hbusreq7 & v3a705ee | !hbusreq7 & v3a62bc6;
assign v3a6f66d = hbusreq7_p & v3767fd7 | !hbusreq7_p & v3a70b50;
assign v373f72a = hbusreq1_p & v3a70415 | !hbusreq1_p & v8455ab;
assign v90fd44 = hready & v3758615 | !hready & v3a713e1;
assign v3a626d4 = hbusreq7 & v3a635b9 | !hbusreq7 & a6c8aa;
assign v3a6c725 = hbusreq0_p & v3a5f8d0 | !hbusreq0_p & v3775303;
assign v3744fb6 = hbusreq5_p & v3736e12 | !hbusreq5_p & v37257e9;
assign v37677a3 = hlock6_p & v3806db7 | !hlock6_p & v3a54c77;
assign v3a6a332 = hmaster0_p & v3a70ca8 | !hmaster0_p & v3733b4b;
assign v2ff8ce3 = hmaster2_p & v373114f | !hmaster2_p & v3752dd0;
assign v3a6f997 = hgrant6_p & v37432c6 | !hgrant6_p & v37474f3;
assign v3a6eaf8 = hmaster0_p & v3a635ea | !hmaster0_p & v374b080;
assign v37286d3 = hbusreq4_p & v3a71415 | !hbusreq4_p & v37676d0;
assign v37673f7 = hbusreq1 & v37718fb | !hbusreq1 & v8455ab;
assign v1e3741b = hgrant0_p & v37773a9 | !hgrant0_p & v380853c;
assign v3778921 = hbusreq0 & v3a53329 | !hbusreq0 & v3743c22;
assign v38074c2 = hbusreq6_p & v374c7f4 | !hbusreq6_p & !v3766bc8;
assign v3a5beb6 = hbusreq6 & v35b7808 | !hbusreq6 & v37425c0;
assign v3a7037a = hmaster0_p & v3a704e9 | !hmaster0_p & v8455ab;
assign v3a6bce9 = hgrant5_p & v375133a | !hgrant5_p & v37239a5;
assign v3a64e29 = hbusreq2 & v3a67284 | !hbusreq2 & b755d3;
assign v374868d = hbusreq2 & v3a70eb6 | !hbusreq2 & v372b7b7;
assign v37434f6 = hbusreq6 & v374362e | !hbusreq6 & v3757024;
assign v3766101 = hmaster0_p & v3a6eb72 | !hmaster0_p & v3a5f992;
assign v374f2fb = hgrant5_p & v373e76c | !hgrant5_p & !v8455ab;
assign v3767e47 = hmaster0_p & v8455bd | !hmaster0_p & v3a6f6c5;
assign ac043d = hbusreq5_p & v3a697d2 | !hbusreq5_p & v376ee43;
assign v3740c8e = hbusreq4 & v37436bc | !hbusreq4 & v8455ab;
assign v3778bef = hbusreq5 & v8639e9 | !hbusreq5 & v377dacb;
assign v3779ea0 = hlock0_p & v3770559 | !hlock0_p & v35772a6;
assign v3728a77 = hbusreq4_p & v37643b5 | !hbusreq4_p & v8455ab;
assign v375003c = locked_p & v3a70278 | !locked_p & !v8455ab;
assign v3776c6e = hlock7 & a0a219 | !hlock7 & v3a5874e;
assign v376166b = hmaster2_p & v3a70374 | !hmaster2_p & v375b880;
assign v3723988 = hmaster2_p & v374f658 | !hmaster2_p & v374f5e0;
assign v376e9b7 = hbusreq2_p & v372cfec | !hbusreq2_p & v8455ab;
assign v377abe1 = hbusreq5 & v374314f | !hbusreq5 & v377edd6;
assign v3a6e5f4 = hbusreq2_p & v3742d37 | !hbusreq2_p & v372f532;
assign v3a67aa1 = hmaster1_p & v3a67d66 | !hmaster1_p & v3a6f426;
assign v37357ce = hlock5_p & v37502f1 | !hlock5_p & !v376bb7a;
assign v3751e8d = hbusreq3 & v37482f8 | !hbusreq3 & !v3a703df;
assign v37717f4 = hbusreq1_p & v373df14 | !hbusreq1_p & v374f4a0;
assign v3a6f408 = hgrant2_p & v3a70645 | !hgrant2_p & v3742655;
assign v3a5e783 = hmaster0_p & v3a635ea | !hmaster0_p & v3a6fb57;
assign v3a5b70a = hlock4 & v37667f7 | !hlock4 & v3723fce;
assign v3742a78 = hbusreq2_p & v376de4e | !hbusreq2_p & v39eb569;
assign v3a6c050 = hmaster2_p & v8455ab | !hmaster2_p & v3a56b05;
assign v372e544 = hmaster0_p & v3729178 | !hmaster0_p & !v3764585;
assign v3a58b8f = hbusreq0 & v3754421 | !hbusreq0 & v377e24d;
assign v3a5c33d = hbusreq4_p & v3767b75 | !hbusreq4_p & v8455b3;
assign v3a706e2 = hbusreq6_p & v37272ed | !hbusreq6_p & !v3767cb7;
assign v3a635f8 = hbusreq0 & v3742723 | !hbusreq0 & v3a6d1fa;
assign v3723747 = hbusreq2 & v3754ec1 | !hbusreq2 & !v3a6fe1a;
assign v377e406 = hbusreq5_p & v37267f3 | !hbusreq5_p & v3742275;
assign v3746b73 = hmaster2_p & v3a5fc34 | !hmaster2_p & v373e114;
assign v3a5958e = hmaster0_p & v3808ed2 | !hmaster0_p & v3742322;
assign v3a6f087 = hmaster1_p & v3745754 | !hmaster1_p & v3a60b37;
assign v37450b8 = hbusreq3_p & v374f35a | !hbusreq3_p & v3a68d2e;
assign v35b774b = hbusreq1_p & v37547c9 | !hbusreq1_p & v8455ab;
assign v3a6ef6d = hgrant6_p & v3743eae | !hgrant6_p & v37384ee;
assign v373dcad = hlock3_p & v94ce87 | !hlock3_p & v3a6958b;
assign v3a2abf5 = hmaster0_p & v3763863 | !hmaster0_p & v373e267;
assign v373e046 = hbusreq2 & v3a5600a | !hbusreq2 & v37757e0;
assign decide = !v3806640;
assign v374ae7a = hmaster0_p & a26fed | !hmaster0_p & v3762ffa;
assign v374faa2 = hlock0 & v376e041 | !hlock0 & v3a71425;
assign v3a6ff24 = hmaster0_p & v375abf4 | !hmaster0_p & v3732c95;
assign v377661b = hgrant5_p & v37742d2 | !hgrant5_p & v3a6ff89;
assign v8ac028 = hmaster3_p & v376fe00 | !hmaster3_p & v3a6b72a;
assign v37271f9 = locked_p & v23fd98d | !locked_p & !v8455ab;
assign v3a71631 = hbusreq0 & v3760f4e | !hbusreq0 & !v8455ab;
assign v373df5c = hgrant7_p & v376636b | !hgrant7_p & v3743038;
assign v3748e5a = hmaster0_p & v360c5d9 | !hmaster0_p & v377402f;
assign v3a714c9 = hbusreq1_p & v372a7c9 | !hbusreq1_p & v376cf85;
assign v37367e3 = hmaster2_p & v372d905 | !hmaster2_p & v8455ab;
assign v3774f4e = hbusreq4 & v37556ec | !hbusreq4 & v375e12d;
assign v3752577 = hgrant6_p & v3777996 | !hgrant6_p & v374b47b;
assign v3a7011c = hbusreq0_p & v39a537f | !hbusreq0_p & !v1e38224;
assign v3734862 = hbusreq8 & v3a71315 | !hbusreq8 & !v8455ab;
assign v3a61cb2 = hbusreq6_p & v375cfa5 | !hbusreq6_p & v3725717;
assign v375ef1e = hbusreq2_p & v3765013 | !hbusreq2_p & v8455ab;
assign v3a71493 = hgrant5_p & v3a70dfd | !hgrant5_p & v3752bbd;
assign v3a65856 = hbusreq0 & v374cd7e | !hbusreq0 & v3740de5;
assign v3a6f508 = jx0_p & v3a711f7 | !jx0_p & !v3773847;
assign v3a6fdc9 = hbusreq2_p & v3a6143b | !hbusreq2_p & !v39a4ca8;
assign v37400bc = hgrant3_p & v3754227 | !hgrant3_p & v375f30d;
assign v377b1db = hlock2_p & v3729b33 | !hlock2_p & v8455ab;
assign v3a67f5b = hbusreq5_p & v375b046 | !hbusreq5_p & v376cfae;
assign v374f2d2 = hlock5 & v3a70119 | !hlock5 & v3a71375;
assign v23fde7f = hbusreq8_p & v3a7101a | !hbusreq8_p & v3a6a03c;
assign v372fd11 = hmaster3_p & v3734b6e | !hmaster3_p & !v3a6fb4e;
assign v3770367 = hmaster0_p & v374ae00 | !hmaster0_p & v3757ffa;
assign v377a6dc = hlock0 & v377bfc0 | !hlock0 & v3734e69;
assign v3a5bd58 = hgrant4_p & v3a6d809 | !hgrant4_p & v3748e9d;
assign v3730dc1 = hbusreq7_p & v3734862 | !hbusreq7_p & v8455ab;
assign v376b087 = hbusreq2_p & v3736785 | !hbusreq2_p & v37672ac;
assign v37360df = hmaster1_p & v377a1ef | !hmaster1_p & v3769d79;
assign v3a60008 = hlock2 & v374cd48 | !hlock2 & v377825c;
assign v3774878 = hmaster2_p & v3a714b1 | !hmaster2_p & v8455ab;
assign v372d5ba = hgrant5_p & v375afbf | !hgrant5_p & v3a6fdca;
assign v1e38262 = hbusreq5_p & v3741438 | !hbusreq5_p & !v8455ab;
assign v3742521 = hbusreq6_p & v374faa9 | !hbusreq6_p & v3a6fba1;
assign v372ddea = hbusreq8_p & v3a5aef8 | !hbusreq8_p & v377234d;
assign v374925f = hbusreq5_p & v37374d6 | !hbusreq5_p & !v3a7115d;
assign v376c0c8 = hmaster0_p & v375cddb | !hmaster0_p & v377291b;
assign v377c620 = hmaster1_p & v374bdea | !hmaster1_p & v3a706eb;
assign v375069a = hbusreq4_p & v3806ce9 | !hbusreq4_p & v2092abe;
assign v3a6be6d = hgrant2_p & v8455b9 | !hgrant2_p & v2889705;
assign v375e512 = hmaster0_p & v373a9fb | !hmaster0_p & v3a5992f;
assign v3769a71 = hbusreq5_p & v3a70642 | !hbusreq5_p & v3a62bd5;
assign v3757cd6 = hbusreq0 & v3a6e50e | !hbusreq0 & v3a6ffbd;
assign v37296ca = hmaster3_p & v37410b9 | !hmaster3_p & !v376b1ee;
assign v3762c4c = hgrant5_p & v8455c6 | !hgrant5_p & v375242f;
assign v2619b26 = locked_p & v8455ab | !locked_p & v3735ed0;
assign v3a70a01 = hmaster0_p & v3a67577 | !hmaster0_p & v375e6ff;
assign v3a60c86 = hbusreq4_p & v3a5a72a | !hbusreq4_p & v37331df;
assign v377b732 = hmaster1_p & v374a9e4 | !hmaster1_p & v3752ebb;
assign v373d268 = hbusreq7 & v35b70c9 | !hbusreq7 & v3750fa9;
assign v374373a = hmaster1_p & v3a70a9e | !hmaster1_p & !v373a265;
assign v3a70b37 = hbusreq4 & v3729421 | !hbusreq4 & v8455bd;
assign v372c0d6 = hmaster0_p & v377bb3a | !hmaster0_p & v374ad7d;
assign v377ebf3 = hbusreq7 & v374b4c5 | !hbusreq7 & a0a219;
assign v3735cb3 = hbusreq4_p & v3778355 | !hbusreq4_p & v1e378da;
assign v3751f67 = hgrant3_p & v35b7299 | !hgrant3_p & v3756943;
assign v3a6f149 = hlock0_p & v372e169 | !hlock0_p & v373df9c;
assign v3775e82 = hbusreq4 & v377d785 | !hbusreq4 & v8455ab;
assign v3a603ad = hlock4 & v376f87a | !hlock4 & v3730c26;
assign v3a6f10e = hbusreq6_p & v374875d | !hbusreq6_p & v376dab5;
assign v3808eed = hgrant4_p & v375c170 | !hgrant4_p & v3a6eba9;
assign v3a6a41e = hlock3_p & v3a70a6f | !hlock3_p & v375ea58;
assign v3a6e40b = hbusreq5 & v373a27c | !hbusreq5 & v8455e7;
assign v37745a0 = hgrant4_p & v3733e9e | !hgrant4_p & v37711c5;
assign v39a535f = hbusreq3_p & v2acb5a2 | !hbusreq3_p & !v8455ab;
assign v3770bf5 = hlock6 & v3a6f659 | !hlock6 & v3a6f914;
assign v3751d6f = hmaster2_p & v37430c6 | !hmaster2_p & v3a68838;
assign v3a66110 = busreq_p & v39a537f | !busreq_p & !v1e38224;
assign v3733e62 = hbusreq4_p & v373d7f9 | !hbusreq4_p & v3a70315;
assign v3758869 = hbusreq0 & v373bda7 | !hbusreq0 & v377f104;
assign v375cade = hgrant3_p & v376f0c1 | !hgrant3_p & v3777baa;
assign v377057c = hlock4_p & v3a6eb39 | !hlock4_p & v35772a6;
assign v3766448 = hlock1_p & v3778ed4 | !hlock1_p & v8455e7;
assign v3759b63 = hbusreq4_p & v373ccde | !hbusreq4_p & v372348c;
assign v374cd7e = hlock4 & v373d753 | !hlock4 & v376b1be;
assign v3726efd = hbusreq7_p & v373bfd3 | !hbusreq7_p & v3807bfa;
assign v373e80b = start_p & v845605 | !start_p & v372ccea;
assign v37458a2 = hmaster1_p & v376bd2c | !hmaster1_p & v374016f;
assign v374c120 = hmaster0_p & v8455e7 | !hmaster0_p & v3756954;
assign v372d49e = jx0_p & v3a6af4d | !jx0_p & v3a70ebb;
assign v3a71686 = hbusreq6_p & v3a703d3 | !hbusreq6_p & v39eb4a7;
assign v3a709f2 = hbusreq0 & v23fdf30 | !hbusreq0 & v3736d43;
assign v3a70e4b = hgrant4_p & v8455ab | !hgrant4_p & v37562a5;
assign v373d9e4 = hmaster0_p & v3765c35 | !hmaster0_p & v3a5cf5e;
assign v37276f2 = hbusreq0 & v376a9de | !hbusreq0 & v37662e2;
assign v377bd81 = hbusreq5_p & v377de7f | !hbusreq5_p & v3734ca9;
assign v3a5cb57 = hbusreq6_p & v3a5f8d0 | !hbusreq6_p & v3775303;
assign v37758d3 = hbusreq8 & v375d102 | !hbusreq8 & v8455ab;
assign v374915c = jx0_p & v3747e71 | !jx0_p & v3a6338d;
assign v374c88d = hmaster2_p & v8455ab | !hmaster2_p & v292555a;
assign v337897a = hgrant2_p & v8c4a86 | !hgrant2_p & v3760279;
assign v377657c = hbusreq6 & v3a69062 | !hbusreq6 & v3a70e8d;
assign v3a56dff = jx0_p & v9259bc | !jx0_p & v372509d;
assign v3732736 = hbusreq5 & v3378f4e | !hbusreq5 & v3739b5c;
assign v3378b65 = jx0_p & v3a5e2af | !jx0_p & v3a6f973;
assign v3a5b687 = hmaster1_p & v3a5fabd | !hmaster1_p & v37612c1;
assign v3735f79 = hmaster2_p & v3a6fe52 | !hmaster2_p & v3a6ffd0;
assign v37706ae = hmaster0_p & v3a635ea | !hmaster0_p & v3a594fe;
assign v376fbce = hbusreq8 & v3763046 | !hbusreq8 & v3a6fd20;
assign v3776cda = hbusreq8_p & v3a64e13 | !hbusreq8_p & v3a6fdec;
assign v3a70ad2 = hbusreq2 & v3776aa8 | !hbusreq2 & v8455ab;
assign v3750c0c = hbusreq5 & v376a6f1 | !hbusreq5 & v3742be5;
assign v374d4d3 = hmaster2_p & v373b9d6 | !hmaster2_p & v3a6f8d0;
assign v3a675f7 = hbusreq0 & v3759f66 | !hbusreq0 & v3728213;
assign v3724200 = hgrant2_p & v377182c | !hgrant2_p & v375b9c3;
assign v3742be5 = hmaster0_p & v375248f | !hmaster0_p & v376a6f1;
assign v3726344 = hbusreq0 & v3a6d4bf | !hbusreq0 & v37502ca;
assign v372b8a5 = hmaster0_p & v3730829 | !hmaster0_p & !v37670ac;
assign v3a70853 = hgrant4_p & v37245f8 | !hgrant4_p & v3a64225;
assign v3759b7c = hbusreq3 & v37481f3 | !hbusreq3 & v37735ec;
assign v3768421 = hmaster2_p & v37737aa | !hmaster2_p & v3758133;
assign v377ea6c = hmaster0_p & v39ea76e | !hmaster0_p & v3a533d8;
assign v3777692 = hgrant2_p & v37234e0 | !hgrant2_p & !v375e1a2;
assign v39ebb63 = hbusreq5_p & v37551b0 | !hbusreq5_p & v3729b52;
assign v2ff9314 = hbusreq2_p & v3764efe | !hbusreq2_p & v8455ab;
assign v377217f = hgrant1_p & v377b6ce | !hgrant1_p & !v35772a6;
assign v3724621 = hlock4_p & v3733c46 | !hlock4_p & v3778993;
assign v3a6ec83 = hmaster1_p & v3778372 | !hmaster1_p & v3762145;
assign v3a60a9f = hmaster0_p & v37432cd | !hmaster0_p & v3a624d1;
assign v3735f67 = hbusreq5_p & v3758fa8 | !hbusreq5_p & v3a6eb3d;
assign v3761a32 = hlock5_p & v3a5f9d5 | !hlock5_p & v3a704ca;
assign v3a69a04 = hbusreq6 & v3756e01 | !hbusreq6 & v3744724;
assign v3759421 = hlock7_p & v3808f2f | !hlock7_p & v37770ab;
assign v3778c9a = hmaster3_p & v3732cdc | !hmaster3_p & v377afaa;
assign v37710a1 = hmaster2_p & v373a341 | !hmaster2_p & v3a6efad;
assign v3a7096f = hmaster2_p & v376285a | !hmaster2_p & !v3730749;
assign b3ccfa = hbusreq7_p & v373250a | !hbusreq7_p & !v8455ab;
assign v3a6fa53 = hmaster0_p & v3730e7d | !hmaster0_p & v3a70585;
assign v3737423 = hgrant6_p & v375034b | !hgrant6_p & v3a64252;
assign v373b7c8 = hgrant0_p & v3749529 | !hgrant0_p & v3770e2b;
assign v37494c3 = hmaster0_p & v376c25c | !hmaster0_p & v3777536;
assign v375b01e = hlock5 & v1e379cc | !hlock5 & v3770366;
assign v3772347 = hmaster2_p & v3a5d079 | !hmaster2_p & v3a70891;
assign v3740f9c = hmaster2_p & v375c9f0 | !hmaster2_p & !v3a70fec;
assign v3723227 = hbusreq5 & v373375c | !hbusreq5 & v3760bda;
assign v372dcf7 = hmaster2_p & c5fc63 | !hmaster2_p & v3758df6;
assign v3a710b2 = hbusreq0_p & v37787ec | !hbusreq0_p & v3778528;
assign v3a7071b = hbusreq0 & v3779316 | !hbusreq0 & v376fa94;
assign v3740b8b = hbusreq4 & v373dd77 | !hbusreq4 & v8455ab;
assign v377d2e7 = hbusreq3_p & v37708f1 | !hbusreq3_p & v372cc25;
assign v3a5d841 = hgrant6_p & v3a5cd51 | !hgrant6_p & v3766f2e;
assign v3a6d9ca = hmaster0_p & v373c3e1 | !hmaster0_p & v1e37d8e;
assign v37722cc = hbusreq1 & v3a706c0 | !hbusreq1 & v3a635ea;
assign d1bf3b = hbusreq3_p & v3a71391 | !hbusreq3_p & !v8455ab;
assign v3a61dd0 = hlock5_p & v3a71245 | !hlock5_p & !v8455ab;
assign v2092b90 = hlock8_p & v3a7110f | !hlock8_p & v3762121;
assign v3a56bf0 = hbusreq6_p & v3a6a78c | !hbusreq6_p & v373a2f2;
assign v3a6065f = hbusreq6_p & v3a5988f | !hbusreq6_p & v3731e60;
assign v3750e23 = hmaster2_p & v373997b | !hmaster2_p & v8455ab;
assign v3755793 = hbusreq4_p & v377b4c9 | !hbusreq4_p & v374145d;
assign v3744c9d = hbusreq2_p & v372324a | !hbusreq2_p & v8455ab;
assign v373b9d6 = hbusreq4_p & v3a635ea | !hbusreq4_p & v374aece;
assign v1e3771d = hbusreq0 & v8cb684 | !hbusreq0 & v374999b;
assign v23fe28c = hmaster2_p & v37796ce | !hmaster2_p & v3725717;
assign v3a5d97a = hmaster1_p & v37731ce | !hmaster1_p & acbf77;
assign v3a6c9c2 = hmaster2_p & v3758fa8 | !hmaster2_p & v3a6fd72;
assign v3a712bf = hgrant4_p & v3770719 | !hgrant4_p & v3a5d08e;
assign v3a710f7 = hmaster2_p & v3a54aa0 | !hmaster2_p & v3a6f995;
assign v3763175 = hready & v3727345 | !hready & !v8455ab;
assign v375e99f = hbusreq4_p & v3a551f9 | !hbusreq4_p & v377eb00;
assign v376d0b5 = hbusreq7 & v3766f51 | !hbusreq7 & v3a6f1e8;
assign v372e669 = hbusreq0 & v372e468 | !hbusreq0 & v3a6ec03;
assign v3770ae6 = hlock3 & v3a56e5e | !hlock3 & v3a66e91;
assign v377db14 = hbusreq0 & v3a68954 | !hbusreq0 & v3754176;
assign v376791c = hgrant6_p & v3a65eba | !hgrant6_p & v3a5faaa;
assign v3a6abf7 = hgrant4_p & v375058e | !hgrant4_p & v376725e;
assign v375e85e = hbusreq8_p & v3a6f88a | !hbusreq8_p & v37c37ed;
assign v37323a1 = hbusreq0 & v377fc15 | !hbusreq0 & v3759fb4;
assign v3a662c7 = hbusreq6 & v3743879 | !hbusreq6 & v376ef7a;
assign v372e5d3 = hgrant1_p & v3a6ffae | !hgrant1_p & v372dab1;
assign v376ea99 = hbusreq4_p & v3a585fd | !hbusreq4_p & v3756524;
assign v3a693ca = hlock8_p & v374da21 | !hlock8_p & v37343bd;
assign v3a6f7b5 = hmaster0_p & v3a6ffd3 | !hmaster0_p & ab15ca;
assign v3a6767a = hlock1_p & v3a63e82 | !hlock1_p & !v35772a6;
assign bb49f9 = hmaster0_p & v37388d6 | !hmaster0_p & v3747bfe;
assign v375b980 = hbusreq6 & v372e9f3 | !hbusreq6 & v375da82;
assign v372abc8 = hbusreq6 & v375a4fa | !hbusreq6 & !v8455ab;
assign v3749cea = locked_p & v376402f | !locked_p & v39a5381;
assign v37320bf = hgrant4_p & v3769f61 | !hgrant4_p & v377a942;
assign v3a7005e = hbusreq4 & v3739635 | !hbusreq4 & v37285eb;
assign v3a6cc67 = hlock4 & v3a700e5 | !hlock4 & v377d10c;
assign v3740349 = hbusreq3 & v373a841 | !hbusreq3 & v8455ab;
assign v372f96d = hlock7_p & v3a5770f | !hlock7_p & v3765ed6;
assign v3758d18 = hbusreq0 & v3a6e5e1 | !hbusreq0 & v377871a;
assign v376e2bb = hmaster2_p & v376c4f9 | !hmaster2_p & v8455ab;
assign v3733de8 = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v3739b80;
assign v3752222 = hbusreq6_p & v3a5b286 | !hbusreq6_p & v377a511;
assign v3a7106c = hgrant4_p & v8455ab | !hgrant4_p & v3a6fc96;
assign v374f243 = hbusreq7_p & v373432d | !hbusreq7_p & v3759b93;
assign v3779233 = hbusreq5 & bfe049 | !hbusreq5 & !v3745bbe;
assign v3726609 = hbusreq2 & v37482f8 | !hbusreq2 & !v3a6fe6a;
assign v373ca9e = hbusreq5_p & v3a59de6 | !hbusreq5_p & v3a61f85;
assign v3758c5c = hmaster0_p & v3a5e24e | !hmaster0_p & v3735ec7;
assign v3a2981e = hgrant2_p & v8455ba | !hgrant2_p & v375865a;
assign v372f87c = hlock6 & v3733103 | !hlock6 & v37440a8;
assign v1e37a69 = hbusreq3_p & v37390ba | !hbusreq3_p & v8455ab;
assign v377444f = hbusreq8 & v3a5b979 | !hbusreq8 & v8455b3;
assign v3a65369 = hgrant4_p & v3a67e67 | !hgrant4_p & v373f94e;
assign v376ba89 = hlock4 & v360c1bf | !hlock4 & cfe9c3;
assign v375fb00 = hmaster0_p & v3738686 | !hmaster0_p & v937864;
assign v3a70dfe = hbusreq0 & v3a66e41 | !hbusreq0 & v373e4c0;
assign dc5778 = hmaster1_p & v3752f9b | !hmaster1_p & v2acb110;
assign v3752986 = hmaster3_p & v3767e6a | !hmaster3_p & v3a6ff9c;
assign v374cd43 = hmaster2_p & v3757568 | !hmaster2_p & !v8455ab;
assign v23fd858 = hmaster2_p & v3755002 | !hmaster2_p & v8455b0;
assign v374d6de = hbusreq5_p & v3a6feb8 | !hbusreq5_p & v3a6ffae;
assign v3a71380 = hgrant5_p & v373a4a8 | !hgrant5_p & v373a999;
assign v3a70e3c = hmaster1_p & v3a5b8b9 | !hmaster1_p & v3a613f2;
assign v3a56396 = stateG10_1_p & v37270d9 | !stateG10_1_p & !v373b744;
assign v376db6d = hmaster1_p & v3a638fb | !hmaster1_p & v3779a3c;
assign v372f3fc = hgrant5_p & v3a71576 | !hgrant5_p & v377258d;
assign v374cd18 = hbusreq4_p & v3807a32 | !hbusreq4_p & !v372d60f;
assign d66718 = hbusreq8_p & v3a70d7d | !hbusreq8_p & v3a6eed1;
assign v3a6393d = hbusreq7_p & v8455b7 | !hbusreq7_p & v23fe156;
assign v3758b05 = hmaster0_p & v3a6f04e | !hmaster0_p & v3a658cf;
assign v3766f14 = hbusreq4_p & v3769945 | !hbusreq4_p & v3a6ebf2;
assign v374bc3e = hgrant2_p & v8ef654 | !hgrant2_p & v8455ab;
assign v37637ef = hbusreq4 & v3749435 | !hbusreq4 & v8455ab;
assign v3a6de73 = hgrant3_p & v8455ab | !hgrant3_p & v37533c3;
assign v3a5ef59 = hlock0_p & v374ab5b | !hlock0_p & v3a6fb64;
assign v377195f = hbusreq5_p & v3a71118 | !hbusreq5_p & !v8455ab;
assign v3a65bad = hbusreq4 & v3737ea9 | !hbusreq4 & v8455ab;
assign v376be4c = hbusreq3 & v3a6ca99 | !hbusreq3 & v3a6fdef;
assign v3726a2c = hgrant3_p & v8455be | !hgrant3_p & v3a6f41c;
assign v3a71279 = hgrant5_p & v3764fad | !hgrant5_p & v3725e33;
assign v3a7062c = hbusreq6_p & v376a7b5 | !hbusreq6_p & v8455ab;
assign v3808e85 = hmaster2_p & v376081b | !hmaster2_p & v3a7160f;
assign v374b383 = hgrant0_p & v375a288 | !hgrant0_p & !bbbe50;
assign v3807008 = hbusreq7 & v3744daa | !hbusreq7 & v3a701ad;
assign v376ba53 = hlock2_p & v3a5788f | !hlock2_p & v8455ab;
assign v3a6eebf = hgrant6_p & v3a709a3 | !hgrant6_p & !v8455ab;
assign v374e58f = hmaster1_p & v3a58218 | !hmaster1_p & v3a706be;
assign v3738666 = hmaster0_p & v377accc | !hmaster0_p & v3a672c8;
assign v377a393 = hlock2_p & v372b726 | !hlock2_p & v3a5ab9d;
assign v2aca76c = hmaster3_p & v3733cf4 | !hmaster3_p & v3733955;
assign v3730b5e = hbusreq2_p & v372673b | !hbusreq2_p & v372f532;
assign v377cc6d = hbusreq5_p & v3a61b45 | !hbusreq5_p & v8455ab;
assign v376d3a6 = hlock8 & v376f5ed | !hlock8 & v375c735;
assign d3a479 = hlock5_p & v375abc2 | !hlock5_p & v375f888;
assign v3748229 = hbusreq5_p & v3735050 | !hbusreq5_p & v3a6d9ca;
assign v376cffc = hmaster2_p & v374b8fa | !hmaster2_p & v3a68dfd;
assign v3759aec = hlock5_p & v3761db0 | !hlock5_p & v375cbcb;
assign v37533b4 = stateG10_1_p & v35772a5 | !stateG10_1_p & !v3a63621;
assign v3776974 = jx1_p & v3735d9e | !jx1_p & b4ede7;
assign v375518f = hgrant4_p & v3754b58 | !hgrant4_p & v3743e83;
assign v3a70c95 = hbusreq0 & v3757c10 | !hbusreq0 & v374b3e2;
assign v376b012 = hmaster0_p & v374254d | !hmaster0_p & !v3a6af83;
assign v3a6dc60 = hmaster2_p & v8455ab | !hmaster2_p & v3742122;
assign v37684e6 = hmaster1_p & v3a5a24b | !hmaster1_p & v372873a;
assign v3724744 = stateA1_p & v8455ab | !stateA1_p & !v3727e15;
assign v3741218 = hlock0 & v3a635ea | !hlock0 & v37420e2;
assign v377ee74 = hmaster2_p & v3a6ffca | !hmaster2_p & v3a6a939;
assign v3a5f974 = hbusreq4 & v3733b37 | !hbusreq4 & v8455ab;
assign v209324e = hgrant2_p & v376ddfb | !hgrant2_p & v3a6feaa;
assign v3739743 = hbusreq2 & v3757ae7 | !hbusreq2 & v374a637;
assign v376495c = hlock7_p & v3745e29 | !hlock7_p & v375101b;
assign v3764f27 = hlock6_p & v8455ab | !hlock6_p & v373e21a;
assign v3a70fd9 = hbusreq8 & v37325e0 | !hbusreq8 & v8455ab;
assign v3a5e63b = hbusreq4_p & c7d127 | !hbusreq4_p & v37621e9;
assign v3749ba6 = hbusreq5_p & v3a65088 | !hbusreq5_p & v35772a6;
assign v374b918 = hgrant3_p & v8455be | !hgrant3_p & v3a707f1;
assign v373dd36 = hmaster2_p & v376285a | !hmaster2_p & !v8455ab;
assign v3775ee8 = hgrant0_p & v8455ab | !hgrant0_p & v374b4d6;
assign v3a6a895 = hlock2_p & v376a08d | !hlock2_p & !v8455ab;
assign v373a79f = hmaster3_p & v3a71493 | !hmaster3_p & !v3a62e20;
assign v3739f1f = hbusreq2 & v3a7154e | !hbusreq2 & v3753b7d;
assign v3772e82 = hmaster0_p & v3a5af94 | !hmaster0_p & !v3a6e31f;
assign v3744a67 = hbusreq8 & v3755783 | !hbusreq8 & v373b8c6;
assign v3a6b381 = hbusreq1 & v3a685cd | !hbusreq1 & v377eaf2;
assign v3a71474 = hbusreq4_p & v3756930 | !hbusreq4_p & v37369f2;
assign v3a679ae = hbusreq6_p & v3a6fb7a | !hbusreq6_p & v8455bb;
assign v374e21d = hmaster0_p & v3a58cfc | !hmaster0_p & !v376eaf2;
assign v3a5b8e4 = hlock6 & v3774209 | !hlock6 & v3a6cf19;
assign v3a58378 = hmaster0_p & v3735796 | !hmaster0_p & v37662e7;
assign v380922b = hbusreq4 & v373f8d4 | !hbusreq4 & v3a6df9a;
assign v3772f32 = hmaster0_p & v3806ff5 | !hmaster0_p & v3770cb8;
assign v375c956 = hgrant1_p & v372373f | !hgrant1_p & v373df21;
assign v3a627cc = hbusreq2_p & v37662dc | !hbusreq2_p & v37521ed;
assign v3a6f3d5 = hbusreq2_p & v376e040 | !hbusreq2_p & v3a6ef5f;
assign v3a5e784 = hmaster2_p & v3a6dc08 | !hmaster2_p & v37386cb;
assign v3a70ce4 = hbusreq5 & v23fdead | !hbusreq5 & v8455ab;
assign v3a6dc57 = hmaster2_p & v3a6ffca | !hmaster2_p & v8455ab;
assign c0c2de = hmaster2_p & v375bfdf | !hmaster2_p & v374b5c5;
assign v1e38291 = hmaster1_p & v3a57584 | !hmaster1_p & v373f47b;
assign aed6c7 = hmaster0_p & ce4d7a | !hmaster0_p & v3775f27;
assign v3769d5c = hgrant2_p & v375d12e | !hgrant2_p & v3751faf;
assign v3a60bc8 = hbusreq1_p & v3749c22 | !hbusreq1_p & v3751ca5;
assign v37459dd = hbusreq3 & v3767437 | !hbusreq3 & v8455b3;
assign v3a64225 = hgrant6_p & v37245f8 | !hgrant6_p & v373c983;
assign v37683c2 = hgrant4_p & v3a53eeb | !hgrant4_p & v376067f;
assign v37483dd = hbusreq6_p & v3a5a510 | !hbusreq6_p & !v1e382e7;
assign v3a5e647 = hmaster2_p & v3a635ea | !hmaster2_p & v3a57384;
assign v374b36e = hgrant2_p & v37432c6 | !hgrant2_p & !v376454b;
assign v3a6eb53 = hmaster1_p & v3766799 | !hmaster1_p & v376a40c;
assign v9af5fc = hmaster2_p & v3a70d99 | !hmaster2_p & v37728a5;
assign v3779c38 = hmaster2_p & v8455b0 | !hmaster2_p & v3754c5e;
assign v3a56804 = jx3_p & v3751fde | !jx3_p & v3a70b5c;
assign v3a5fed1 = hmaster1_p & v372fe58 | !hmaster1_p & v3749139;
assign c76b50 = hbusreq8_p & v3a6fbc9 | !hbusreq8_p & !v3a6ebc6;
assign v3a5946d = hgrant8_p & v8455ab | !hgrant8_p & v374e5eb;
assign v372f532 = hgrant3_p & v3a6c2b6 | !hgrant3_p & !v375fabf;
assign v3a6f8cc = hgrant6_p & v8455ab | !hgrant6_p & !v3809399;
assign v3742aff = hlock6_p & v1e38275 | !hlock6_p & v39a537f;
assign v3a70c11 = hgrant0_p & v8455ab | !hgrant0_p & v3a71287;
assign v3a638fe = hlock2 & v3770855 | !hlock2 & v86d3dc;
assign v3a57d9f = hbusreq0 & v372f6ab | !hbusreq0 & v3a6d69b;
assign v375682e = hmaster1_p & v3745c84 | !hmaster1_p & v375d78f;
assign v374546c = hmaster0_p & v3743ff2 | !hmaster0_p & v374e019;
assign v969d5b = hmaster1_p & v3a6f2ba | !hmaster1_p & v3777efb;
assign v3a6b161 = hbusreq8_p & v37605a5 | !hbusreq8_p & v377435f;
assign aa421e = hmaster2_p & v1e377ba | !hmaster2_p & v3a7119c;
assign v3725a56 = hbusreq6 & v39a537f | !hbusreq6 & !v8455ab;
assign v374e3c2 = hgrant3_p & v3752a0d | !hgrant3_p & v373c668;
assign v3a7039e = hlock6_p & v372b24d | !hlock6_p & v3740f3d;
assign v3a710d8 = hbusreq8_p & v37c028b | !hbusreq8_p & v3763c20;
assign v3738ce7 = hbusreq3_p & v3a5e02b | !hbusreq3_p & v37498be;
assign v374cba0 = hgrant3_p & v3a71145 | !hgrant3_p & v3762fc2;
assign v3a5c5b5 = hbusreq6 & v3a6f9c3 | !hbusreq6 & v8455bf;
assign v3808f5d = hmaster1_p & v8455ab | !hmaster1_p & v3758d1e;
assign v373cbc5 = hbusreq5_p & v3744887 | !hbusreq5_p & v8455ab;
assign v3a6effa = hgrant2_p & v38095ed | !hgrant2_p & v377911e;
assign v3756810 = hmaster0_p & v37592d0 | !hmaster0_p & v3a5cf5e;
assign v3753418 = hbusreq0 & v37453d8 | !hbusreq0 & v8455ab;
assign v374f1a1 = hbusreq1_p & v372b0ac | !hbusreq1_p & !v3749ece;
assign v376fc1c = hbusreq4_p & v3a6ef3f | !hbusreq4_p & v37477aa;
assign v1e3828a = hgrant4_p & v3a62184 | !hgrant4_p & v3a59ff7;
assign v3a5966b = hgrant6_p & v3739334 | !hgrant6_p & v8455ab;
assign v3753af9 = hbusreq8_p & v3a6eac2 | !hbusreq8_p & !v3a695c1;
assign v373fe7b = hbusreq6 & v376d081 | !hbusreq6 & v372c500;
assign v3a58da1 = hlock6_p & v3741cda | !hlock6_p & v37506d8;
assign v37577cd = hmaster0_p & v3a7160d | !hmaster0_p & v3a5992f;
assign v3a70796 = hbusreq5 & v372e263 | !hbusreq5 & v374c679;
assign v376363f = hmaster2_p & v374db8d | !hmaster2_p & v8455c3;
assign v376a6bc = hbusreq6_p & b2271d | !hbusreq6_p & v8455ab;
assign cd0aed = hlock5 & v3747452 | !hlock5 & v373c005;
assign v374d63f = hgrant6_p & v1e378b4 | !hgrant6_p & v3a6ebcc;
assign v3a5c733 = hmaster1_p & v3a5a807 | !hmaster1_p & v3a6b6a3;
assign v372b652 = hmaster0_p & v38087ee | !hmaster0_p & !v372ee6a;
assign v3a69957 = hmaster3_p & v3a69203 | !hmaster3_p & v3a71031;
assign v375754a = hmaster2_p & v377766c | !hmaster2_p & v376f569;
assign v3739748 = hbusreq5 & v3a58378 | !hbusreq5 & v3742ca7;
assign v375bbe9 = locked_p & v374c9c7 | !locked_p & v3a66110;
assign v3a7105c = hgrant6_p & v3755e4e | !hgrant6_p & v372ad52;
assign v3a63de8 = hlock0_p & v8455ab | !hlock0_p & v8455b1;
assign v3a6dada = hgrant7_p & v8455ab | !hgrant7_p & v3a678f9;
assign v3a55d4c = hmaster0_p & v373f75b | !hmaster0_p & !v372cdd5;
assign v372e790 = hbusreq0 & v377150c | !hbusreq0 & v3a6ff10;
assign v375da17 = hgrant3_p & v375a268 | !hgrant3_p & v23fdbdc;
assign v3a5a0b3 = hbusreq1 & v374362e | !hbusreq1 & !v3a568f7;
assign v3749a98 = jx3_p & v376f0c3 | !jx3_p & v3a577ed;
assign v3761785 = locked_p & v3a6e7b3 | !locked_p & !v8455ab;
assign v374c679 = hmaster0_p & v9af7ec | !hmaster0_p & v3a6fdbc;
assign v37787d1 = hmaster2_p & v37430c6 | !hmaster2_p & v8455b0;
assign v3764c8a = hgrant6_p & v3a53fa4 | !hgrant6_p & v3772c21;
assign v375b02a = hlock4_p & v377c7c0 | !hlock4_p & v373014d;
assign v37371be = hmaster1_p & v3772374 | !hmaster1_p & v3a6fe83;
assign v3a6783b = hbusreq4_p & v3764702 | !hbusreq4_p & v3a66f07;
assign v3a5e665 = hmaster2_p & v3a713df | !hmaster2_p & v3766202;
assign v374f3a9 = hbusreq7 & v377cb05 | !hbusreq7 & v3a6ffdd;
assign v37400ab = hmaster0_p & v374b887 | !hmaster0_p & v3a6fd0a;
assign v374a41b = hmaster0_p & v376d0bc | !hmaster0_p & v3754d88;
assign v1e3780d = hmaster1_p & v8455b0 | !hmaster1_p & v23fda7e;
assign v374fde8 = hlock5_p & v360d2c6 | !hlock5_p & !v8455ab;
assign v377de4d = hlock7_p & c8ca6f | !hlock7_p & !v37738b2;
assign v9ec00e = hgrant6_p & v3a6eb39 | !hgrant6_p & v3735179;
assign v372a674 = hmaster2_p & v8455ab | !hmaster2_p & v3a709e5;
assign v377e018 = hmaster0_p & v37287e1 | !hmaster0_p & v3a5ac38;
assign v374f0af = hbusreq5 & v3a70706 | !hbusreq5 & !v8455ab;
assign v3a5ace8 = hmaster2_p & v3a6ffb6 | !hmaster2_p & v35b774b;
assign v3a58732 = hbusreq4 & v3a619c0 | !hbusreq4 & !v8455ab;
assign v3a5fabd = hgrant4_p & v3751389 | !hgrant4_p & v3768e70;
assign v3a6b6ef = hgrant4_p & v3739896 | !hgrant4_p & v375b878;
assign v3a6b405 = hbusreq2_p & v3732949 | !hbusreq2_p & !v8455ab;
assign c118e3 = hmaster2_p & v374306c | !hmaster2_p & v3a5b5d3;
assign v373e163 = hmaster0_p & v1e382e7 | !hmaster0_p & !v3a5a510;
assign v3770d93 = hgrant6_p & v209323b | !hgrant6_p & v37463de;
assign v3a7047e = hlock2 & d9a7db | !hlock2 & v3771e95;
assign v3809d53 = hgrant5_p & v8455c6 | !hgrant5_p & v3a6fef2;
assign v372d8bd = jx1_p & v374b237 | !jx1_p & !v3a56194;
assign v3755a2f = hgrant2_p & v3a710f9 | !hgrant2_p & !v8455ab;
assign v377b233 = hlock8_p & v373afa4 | !hlock8_p & !v37519dd;
assign v3a70530 = hbusreq6_p & v8455ab | !hbusreq6_p & v3a6a939;
assign v3a65dce = hmaster1_p & v8455e7 | !hmaster1_p & v3730d6e;
assign v376f942 = hbusreq5_p & v374b8fa | !hbusreq5_p & v375ee68;
assign v3a70832 = hgrant2_p & v376dcdc | !hgrant2_p & v3a29842;
assign v374b879 = hmaster0_p & v377adf5 | !hmaster0_p & v37234d1;
assign v2ff9371 = hmaster0_p & v3a6fcea | !hmaster0_p & v373d67c;
assign v374a39f = hmaster1_p & v3a29814 | !hmaster1_p & v375c7cd;
assign v3a70b52 = hbusreq7 & v3756d6e | !hbusreq7 & v3a6f6e0;
assign v3778f83 = hbusreq0_p & v372c3d4 | !hbusreq0_p & !v3a5ef5c;
assign v3762f5b = hmaster1_p & v3a704a3 | !hmaster1_p & v3a5eb8f;
assign v375370a = hlock4 & v3a70fc9 | !hlock4 & v3a6fe44;
assign v376dc2e = hgrant1_p & v8455ab | !hgrant1_p & v3a635ea;
assign v37699a0 = hbusreq2_p & v3763e88 | !hbusreq2_p & !v8455ab;
assign v3a709bf = hlock0_p & v373da69 | !hlock0_p & v37c014e;
assign v3a657d3 = hlock8_p & v375c648 | !hlock8_p & v3a7064e;
assign v37519dd = hmaster1_p & v3a6dfb2 | !hmaster1_p & v37270ad;
assign v374e085 = hlock0 & v3a6f044 | !hlock0 & v2092bcb;
assign v3755e29 = hlock0_p & v372ac5c | !hlock0_p & v3773ba2;
assign v377aa4d = hbusreq8 & v3a7117d | !hbusreq8 & v375c8db;
assign v3a71678 = hgrant4_p & v3a62a6d | !hgrant4_p & v377dae3;
assign v906a66 = hmaster0_p & v3a5e9a8 | !hmaster0_p & v37399d0;
assign v3a6fd37 = hgrant6_p & v376f2f8 | !hgrant6_p & v37705de;
assign v3756b7b = hbusreq7_p & v3a6f414 | !hbusreq7_p & v3a6f8b7;
assign v23fdbfc = hbusreq8_p & v3726fff | !hbusreq8_p & v3a6e152;
assign v37360c8 = hlock5_p & v3a712d8 | !hlock5_p & !v3a61e9f;
assign v377e9a5 = hmaster0_p & v3a6d499 | !hmaster0_p & v3774bdf;
assign v3a6ebe6 = hbusreq6_p & v37432c6 | !hbusreq6_p & !v37521ed;
assign v39e9ca4 = decide_p & v37304a2 | !decide_p & v376a27b;
assign v377184d = hgrant2_p & v377b6ce | !hgrant2_p & !v3a5c2f4;
assign v3775d76 = hlock6 & v3729e5f | !hlock6 & v375f317;
assign v3a6fa17 = hlock5_p & v372b219 | !hlock5_p & v3a714a3;
assign v3a6d2ed = hlock5 & v3727830 | !hlock5 & v376c6fb;
assign v3769cac = hmaster0_p & v3750746 | !hmaster0_p & v3a710c4;
assign v37764d7 = hbusreq1 & v372b24d | !hbusreq1 & !v8455ab;
assign v3a58022 = hmaster0_p & v3725589 | !hmaster0_p & v3758395;
assign v37510b9 = hmaster0_p & v373f11a | !hmaster0_p & v8455e7;
assign v3764bca = hgrant2_p & v8455ab | !hgrant2_p & !v3a7041e;
assign v375caa0 = hbusreq5 & v3a6f2dc | !hbusreq5 & v35ba1cf;
assign v3a70aa4 = hgrant3_p & v8455be | !hgrant3_p & !v3a704d9;
assign v373782c = jx1_p & v3742472 | !jx1_p & v1e37c79;
assign v3765322 = jx0_p & v374e2a0 | !jx0_p & !v3725b1f;
assign v3750d44 = hgrant6_p & v8455ca | !hgrant6_p & v3a6eb33;
assign v2092ec6 = hmaster2_p & v3a63eaf | !hmaster2_p & v373ee17;
assign v3739509 = hbusreq2 & v3a5600a | !hbusreq2 & v3773b23;
assign v3a6dcf3 = hbusreq5_p & v374e5fa | !hbusreq5_p & v3a656a4;
assign v375b659 = hbusreq5_p & v3a58ddb | !hbusreq5_p & v377a865;
assign v3a644e6 = hgrant2_p & v8455ab | !hgrant2_p & v37789a0;
assign v3a71360 = hmaster1_p & v8455ab | !hmaster1_p & v3a703f7;
assign v3770957 = hmaster2_p & v377de7b | !hmaster2_p & v3776685;
assign v3a68dab = hmaster0_p & v3764e37 | !hmaster0_p & !v3741922;
assign v3a66f81 = hgrant0_p & v3a635ea | !hgrant0_p & v376b269;
assign v3757182 = hbusreq2_p & v376278c | !hbusreq2_p & v376c747;
assign v377541e = jx0_p & v3734ed6 | !jx0_p & v8455ab;
assign v37674fb = hbusreq8_p & v3a6f123 | !hbusreq8_p & v3a712b7;
assign v376af20 = hmaster2_p & v374f307 | !hmaster2_p & !v3a7151d;
assign v3a6fcb9 = hbusreq0_p & v3733383 | !hbusreq0_p & v8455ab;
assign v3764684 = hmaster2_p & v3a635ea | !hmaster2_p & v3a687a7;
assign v3763f48 = hbusreq2 & v3730e7d | !hbusreq2 & v3a62a6d;
assign v3a70113 = hbusreq6 & v37489ea | !hbusreq6 & v8455ab;
assign v3744898 = hbusreq5 & v3a701a1 | !hbusreq5 & v3764ee3;
assign v3a6f4f8 = hbusreq4_p & v3a70893 | !hbusreq4_p & v373cd16;
assign v3a6178e = hbusreq7 & v372b59f | !hbusreq7 & v377e3fe;
assign v373ead8 = hbusreq0_p & v3a635ea | !hbusreq0_p & v373b288;
assign v373e55b = hlock5_p & v377a887 | !hlock5_p & !v8455ab;
assign v3a53d44 = hmaster1_p & v3a6f617 | !hmaster1_p & v37579f1;
assign v3a6efc7 = hmaster2_p & v37356b4 | !hmaster2_p & v376d1bb;
assign v3a6a87d = hbusreq7_p & v3778ae9 | !hbusreq7_p & v3a5445e;
assign v3a605e2 = hbusreq6_p & v3749bef | !hbusreq6_p & v373376b;
assign v376a84d = hbusreq5_p & cc8b5a | !hbusreq5_p & v3a7110e;
assign v2092eb6 = hmaster1_p & v374f0c1 | !hmaster1_p & v37680de;
assign v375e34d = hgrant7_p & v8455ab | !hgrant7_p & v37629d2;
assign v3a6f5d1 = hgrant2_p & v3758472 | !hgrant2_p & v3751f67;
assign v3a62ad0 = hmaster2_p & v37665bf | !hmaster2_p & v373a841;
assign v3a5dd1a = hbusreq0 & v3731596 | !hbusreq0 & v8455ab;
assign v3a7108a = hbusreq2 & v375de18 | !hbusreq2 & !v373c755;
assign v3a6becc = hbusreq7_p & v3a6f7b6 | !hbusreq7_p & v372fff7;
assign cd3c6e = hbusreq2_p & v37430c2 | !hbusreq2_p & v3778cdd;
assign v37486de = hmaster2_p & v3a7024f | !hmaster2_p & v3771d4f;
assign v375f504 = hgrant6_p & v377f21b | !hgrant6_p & v3a6f408;
assign v372edf9 = hgrant6_p & v8455ca | !hgrant6_p & v377c7cf;
assign v3722de8 = hmaster2_p & v374f307 | !hmaster2_p & v3a7156d;
assign v37403ea = hgrant2_p & v3a5f50e | !hgrant2_p & v3a6f77a;
assign v37249fe = hmaster1_p & v3742649 | !hmaster1_p & v8455ab;
assign v3744fbb = hbusreq3_p & v3745291 | !hbusreq3_p & !v8455ab;
assign v3755066 = hmaster1_p & v374306c | !hmaster1_p & v3a70c85;
assign v377abb1 = hbusreq2 & v3775c0a | !hbusreq2 & v3a6f6fa;
assign v3731bcf = hlock0_p & v3a69515 | !hlock0_p & v3727638;
assign v3734a96 = hbusreq7_p & v3a69da8 | !hbusreq7_p & v372eb0f;
assign v373c72a = hgrant5_p & v8455ab | !hgrant5_p & v3a5d186;
assign v3751159 = hbusreq5_p & v3757ee7 | !hbusreq5_p & v8455ab;
assign v3742441 = jx3_p & v3a64c32 | !jx3_p & v958697;
assign v3754717 = hbusreq5 & v3725371 | !hbusreq5 & !v8455c2;
assign v3a5c188 = hmaster0_p & v3a71189 | !hmaster0_p & !v3746ea0;
assign v37504fd = hmaster2_p & v3a69727 | !hmaster2_p & v3728d9c;
assign v3722a46 = hmaster0_p & v376e5ab | !hmaster0_p & v373dbfe;
assign v3774cf5 = hbusreq8_p & v3a71076 | !hbusreq8_p & v37523f8;
assign d7e38d = hlock5_p & v3a715d1 | !hlock5_p & !v3a6f5cd;
assign v3723b5b = hbusreq0 & v3754a42 | !hbusreq0 & v3a53873;
assign v3a5d90d = hbusreq8_p & v3a69ce6 | !hbusreq8_p & v380880f;
assign v3a6f06a = hmaster1_p & v3a5e24e | !hmaster1_p & v3a53f38;
assign v375ad94 = hbusreq4 & v3a5b7b9 | !hbusreq4 & v372e83f;
assign v37618ad = hbusreq6 & v3723495 | !hbusreq6 & v372dd89;
assign v3a6fc35 = hlock5_p & v3a6fa7a | !hlock5_p & v3a6f632;
assign v376cf3f = hgrant6_p & v8455ab | !hgrant6_p & v3807ac3;
assign v372eae4 = hbusreq2 & v3a55b2d | !hbusreq2 & v376bade;
assign v375899a = hmaster2_p & v37718cc | !hmaster2_p & v3728d9c;
assign v3727f3b = hmaster2_p & v3806db0 | !hmaster2_p & v3727ad4;
assign v3a6f751 = hbusreq4 & cff2df | !hbusreq4 & v376beb4;
assign v3748f40 = hbusreq8 & v3a64f1f | !hbusreq8 & v3740922;
assign v3736ef2 = hbusreq5_p & v3a70642 | !hbusreq5_p & v37536b2;
assign v373a47e = hbusreq6_p & v3751734 | !hbusreq6_p & v3746265;
assign v3a6146c = hbusreq8 & v377f35c | !hbusreq8 & !v8455ab;
assign v3a7091d = hmastlock_p & v376282b | !hmastlock_p & !v8455ab;
assign v3779801 = hbusreq0 & v3a6f3cf | !hbusreq0 & !v8455ab;
assign v9a2413 = hlock0 & v3a635ea | !hlock0 & v3a68310;
assign v376ccd6 = hmaster0_p & afa913 | !hmaster0_p & v375d3fd;
assign v3779e29 = hmaster1_p & v375db64 | !hmaster1_p & v3a59c1d;
assign v3a6480b = hbusreq6 & v3754c86 | !hbusreq6 & v8455ab;
assign v376e5de = hbusreq5 & v3758c41 | !hbusreq5 & v3a6c7e8;
assign v3a6f5a4 = hmaster1_p & v8455ab | !hmaster1_p & v3764869;
assign v377c07a = hbusreq6 & v37547ad | !hbusreq6 & v3a5641a;
assign v3737d3f = hlock4 & v3749d3f | !hlock4 & v374852b;
assign v3a64474 = hlock3 & v38072fd | !hlock3 & v376a87b;
assign v3776d32 = hgrant5_p & v37300d7 | !hgrant5_p & v917443;
assign v37477b7 = hbusreq7 & v373852b | !hbusreq7 & v373ba25;
assign v375fc73 = hbusreq7 & v3a70727 | !hbusreq7 & v3749503;
assign v373026f = hmaster2_p & v3a70987 | !hmaster2_p & v3746d2a;
assign v3a714cd = hmaster0_p & v372bfcc | !hmaster0_p & v3a6c803;
assign v3729480 = stateA1_p & v8455e1 | !stateA1_p & !v3a54427;
assign v3806bd9 = hmaster1_p & v376fe0c | !hmaster1_p & v3765960;
assign v3a60b1b = hbusreq5 & v3a5ce0f | !hbusreq5 & v8455ab;
assign v376f516 = hgrant5_p & v8455ab | !hgrant5_p & v3a6adf2;
assign v374e124 = hgrant4_p & v3a7133d | !hgrant4_p & v37696a2;
assign v3727eb8 = hbusreq2 & v374c5b2 | !hbusreq2 & v3730122;
assign v3809d9e = hmaster2_p & v373daa8 | !hmaster2_p & v3731991;
assign v3a5c1e7 = hbusreq7 & v375f938 | !hbusreq7 & v8455c3;
assign v373e4a7 = hmaster1_p & v3806f0b | !hmaster1_p & v37477cb;
assign v374cb44 = hbusreq6_p & v372a347 | !hbusreq6_p & v35772a6;
assign v3a70b39 = hgrant6_p & v377f09a | !hgrant6_p & v37403ea;
assign v374e4ec = hmaster2_p & v374e0f6 | !hmaster2_p & v3a6f23a;
assign v3a70356 = hmaster0_p & v3758fa8 | !hmaster0_p & v3a576a4;
assign v3748179 = hmaster2_p & v372ccbe | !hmaster2_p & v37284d5;
assign v37504a9 = hlock6 & ce69d1 | !hlock6 & v376e02e;
assign v372dcac = hmaster0_p & v3768c97 | !hmaster0_p & v3a6ef7f;
assign v3a63ae9 = hmaster2_p & v3a6f4ba | !hmaster2_p & v376e35e;
assign v3a6f9bb = hmaster3_p & v8455ab | !hmaster3_p & v23fdaf1;
assign v37746ea = hgrant6_p & v3776d97 | !hgrant6_p & v3a6f6b6;
assign v373ab2b = hbusreq8 & v3740a1e | !hbusreq8 & v3777d70;
assign v377c4b7 = hbusreq0 & v3809879 | !hbusreq0 & v373b46b;
assign v3a569e1 = hbusreq2_p & v3a66983 | !hbusreq2_p & v376454b;
assign v3759611 = hbusreq5_p & v8455ab | !hbusreq5_p & v3a5b875;
assign v37628cd = hmaster2_p & v2092ba8 | !hmaster2_p & v3a6932d;
assign v37680de = hmaster0_p & v374f0c1 | !hmaster0_p & v3a6f64a;
assign v3752e42 = hmaster2_p & v3a56cdb | !hmaster2_p & !v3732569;
assign v377df60 = hbusreq2_p & v37273be | !hbusreq2_p & v376fa76;
assign v3737928 = hmaster0_p & v3a70af6 | !hmaster0_p & !v377f34a;
assign v375237c = hmaster0_p & v3a5ddc1 | !hmaster0_p & v9c0027;
assign v37333bb = hlock4 & v372eb1a | !hlock4 & v3727580;
assign v376fdd6 = hbusreq6 & v376dcd0 | !hbusreq6 & v373daac;
assign v372b6a1 = hbusreq7_p & v3744a67 | !hbusreq7_p & v375de66;
assign v377695e = hbusreq5_p & v8455ab | !hbusreq5_p & c9c058;
assign v377476b = hbusreq6 & v375859f | !hbusreq6 & v3766e4a;
assign v3a57660 = hbusreq6 & v372ff9e | !hbusreq6 & v8455ab;
assign v39ebb20 = hbusreq6 & v3736f3b | !hbusreq6 & v3770f6e;
assign v3740ad9 = hgrant5_p & v8455ab | !hgrant5_p & v3a5d989;
assign v37422af = jx0_p & v374c885 | !jx0_p & d60033;
assign v3a70d65 = hgrant1_p & v3735e39 | !hgrant1_p & v39a537f;
assign v3a6ff2c = hbusreq0 & d5ffe1 | !hbusreq0 & v376a0fc;
assign v375cebd = hbusreq7_p & v1e3778c | !hbusreq7_p & v8c9ea7;
assign v3727cd0 = hbusreq6_p & v3a6fbe6 | !hbusreq6_p & v3766d1b;
assign v3a566eb = hgrant4_p & v3a6ffea | !hgrant4_p & v3a70c9b;
assign v3739768 = hbusreq7_p & v3a70195 | !hbusreq7_p & v3a6c43c;
assign v3808874 = hbusreq0 & v372a886 | !hbusreq0 & v8455ab;
assign v1e37b65 = hbusreq2 & v377834b | !hbusreq2 & v3a62a6d;
assign v374c95a = hbusreq0 & v3a69dc1 | !hbusreq0 & v3755820;
assign v3a6dbbf = hlock8 & ac4b49 | !hlock8 & v37517f7;
assign v3a6c73d = hmaster3_p & v374915c | !hmaster3_p & v3a6f886;
assign v3a6628b = hmaster2_p & v3747302 | !hmaster2_p & v377d58d;
assign v3753e8e = hgrant5_p & v3759758 | !hgrant5_p & !v8455ab;
assign v3750c50 = hbusreq4_p & v20d166d | !hbusreq4_p & v3776386;
assign v372a966 = hmaster2_p & v373186a | !hmaster2_p & v8455ab;
assign v3a5e7f7 = hbusreq5_p & v3744593 | !hbusreq5_p & v376ba56;
assign v3a538bd = hbusreq0 & v2aca778 | !hbusreq0 & v375c944;
assign v375df77 = hbusreq3_p & v374f0e7 | !hbusreq3_p & v8455b3;
assign v3a66a6e = hbusreq6 & v3a5952d | !hbusreq6 & v3a707c4;
assign v3a6ff87 = hlock4_p & v3739dae | !hlock4_p & v377c34f;
assign v3766607 = hmaster1_p & v374193d | !hmaster1_p & v3a6b78f;
assign v3753a9f = hmaster1_p & v3a6ad46 | !hmaster1_p & v372ffd3;
assign v376269a = hbusreq4_p & v3a5fa81 | !hbusreq4_p & v375cc11;
assign v3a6dca6 = hmaster1_p & v377b9fd | !hmaster1_p & v8455ab;
assign v374b549 = hmaster0_p & v373b18b | !hmaster0_p & v3a70574;
assign v3a701e4 = hbusreq2_p & v3745f76 | !hbusreq2_p & v3a67c13;
assign v377c7cf = hgrant2_p & v8455ba | !hgrant2_p & v3a29706;
assign v3743a4c = hmaster1_p & v3a635ea | !hmaster1_p & v3a69923;
assign v3a70063 = hbusreq8 & v3758e73 | !hbusreq8 & v3765e47;
assign v37273b0 = hmaster2_p & v372455c | !hmaster2_p & !v3a55033;
assign v3a57672 = hmaster2_p & v3757966 | !hmaster2_p & v3775688;
assign v3776996 = hlock3_p & v37507be | !hlock3_p & v2aca977;
assign v3a6dd1a = hmaster0_p & v373ff04 | !hmaster0_p & v3a5d8bb;
assign v3a6fb29 = hlock4_p & v37556fd | !hlock4_p & v3a70530;
assign v374e4c9 = stateG10_1_p & v8455ab | !stateG10_1_p & !v3a6db4b;
assign v376f345 = hgrant2_p & v3758472 | !hgrant2_p & !v3a6d364;
assign v373d449 = hgrant5_p & v8455c6 | !hgrant5_p & v380755c;
assign v3756e01 = hlock6_p & v3a5600a | !hlock6_p & v8455b0;
assign v376e029 = hbusreq5 & d3ed45 | !hbusreq5 & !v3745bbe;
assign v37734d2 = hlock7 & v37441a3 | !hlock7 & v3a65755;
assign v3a5f3f0 = hmaster1_p & v3a6f433 | !hmaster1_p & v8455ab;
assign v3729793 = hmaster2_p & v8455ab | !hmaster2_p & v39eb590;
assign v376de99 = hbusreq0 & v3767437 | !hbusreq0 & v8455ab;
assign v3a6fdde = hbusreq4_p & v3757aa1 | !hbusreq4_p & v377b576;
assign v3a69973 = hmaster1_p & v8455ab | !hmaster1_p & v37381c2;
assign v375f71d = hbusreq2_p & v37765e1 | !hbusreq2_p & v3a6a393;
assign v3a5f0a5 = hlock5 & v3a6913c | !hlock5 & v3a62250;
assign v3760927 = hmaster0_p & v3a5a04c | !hmaster0_p & v3742b6a;
assign v375fe15 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3749f9d;
assign v3a6708c = hbusreq0 & v372cbfc | !hbusreq0 & v8455ab;
assign v3a67bbd = hbusreq5 & v3a674fd | !hbusreq5 & v8455ab;
assign bc3d4a = hbusreq5_p & v3a70ed4 | !hbusreq5_p & v3a695c2;
assign v3776db0 = hmaster0_p & v3a63166 | !hmaster0_p & v377d95a;
assign v3a7089b = hmaster2_p & v377989c | !hmaster2_p & v37665bf;
assign v3766b6e = hlock5 & v377de7f | !hlock5 & v37786f3;
assign v377224f = hmaster2_p & v3a619c0 | !hmaster2_p & v39a537f;
assign v3766727 = hbusreq4 & v3a71540 | !hbusreq4 & v3a6bf41;
assign v376f938 = hgrant3_p & v375917f | !hgrant3_p & v3809f1c;
assign v375c0c4 = hlock4 & v373d0d1 | !hlock4 & v377e29a;
assign v375add8 = hgrant2_p & v8455ab | !hgrant2_p & v3724b93;
assign v375f0c9 = hlock5 & v375eaea | !hlock5 & v3806575;
assign v372d75a = hbusreq5 & v37591e8 | !hbusreq5 & v3a585b7;
assign v1e37349 = hbusreq5_p & v3a6ffdc | !hbusreq5_p & v37783ba;
assign v37297e8 = hmaster2_p & v3779680 | !hmaster2_p & v3a60b2e;
assign v377ece3 = hlock8 & v375c7a3 | !hlock8 & v3a6fbf6;
assign v3768ecc = hlock0_p & v3740171 | !hlock0_p & v3726464;
assign v376ac10 = hbusreq7 & v3727e25 | !hbusreq7 & v3734279;
assign v3a671de = hbusreq4_p & v3a68d70 | !hbusreq4_p & v3a6fa3f;
assign v37283a8 = hlock3_p & v3735e39 | !hlock3_p & v376d856;
assign v372be59 = hlock6_p & v37569ec | !hlock6_p & v37506d8;
assign v377012f = hbusreq8_p & v3771303 | !hbusreq8_p & v374637b;
assign v3722e04 = hlock5_p & v3a7110d | !hlock5_p & v3a70448;
assign v3a70275 = hlock0 & v377b946 | !hlock0 & v373e2d3;
assign v373bbe6 = hmaster1_p & v3757dc4 | !hmaster1_p & v3a5d3f6;
assign v3733c46 = hbusreq3_p & v3a70641 | !hbusreq3_p & v3733383;
assign v376a3f5 = hbusreq5_p & v37365fa | !hbusreq5_p & !v372b91e;
assign v3742b79 = hbusreq5_p & v3a5bf4c | !hbusreq5_p & v3744081;
assign v3a71105 = hbusreq5 & v3768888 | !hbusreq5 & v3a6dfa3;
assign v3725b9b = hmaster2_p & v3a6f018 | !hmaster2_p & v3757aa1;
assign v3763868 = hgrant6_p & v2acaf72 | !hgrant6_p & !v375f326;
assign v3a70ff2 = hbusreq7_p & v376da21 | !hbusreq7_p & v37550ac;
assign v3767985 = hmaster2_p & v8455ab | !hmaster2_p & !v377b4c9;
assign v3737e2c = hmaster2_p & v3747302 | !hmaster2_p & v3735525;
assign v3a5e4f4 = hgrant6_p & v3739884 | !hgrant6_p & v3a70057;
assign v375a6be = hmaster0_p & v373cd03 | !hmaster0_p & v3733d02;
assign v3a69a39 = hbusreq4 & v372952e | !hbusreq4 & v3a708c2;
assign v376a96b = hbusreq2_p & v3729991 | !hbusreq2_p & v8455bf;
assign v37786bb = hbusreq6 & v3a5e748 | !hbusreq6 & !v8455ab;
assign v2ff8be4 = hgrant3_p & v8455ab | !hgrant3_p & v373ca0e;
assign v3a706f4 = hbusreq5_p & v3a5d3fc | !hbusreq5_p & !v37291f4;
assign v37785be = hbusreq0 & v3723048 | !hbusreq0 & v8455ab;
assign v3a6b924 = hgrant4_p & v376d2b7 | !hgrant4_p & v377d377;
assign v3a6aaed = hlock5_p & v3a65ee0 | !hlock5_p & v8455ab;
assign v377da1e = hmaster0_p & v376a31b | !hmaster0_p & v3a715f7;
assign v372bd23 = hbusreq4 & v3a5cb57 | !hbusreq4 & v8455ab;
assign v37242b9 = hbusreq5_p & v38093c2 | !hbusreq5_p & v3a70100;
assign v3806624 = jx0_p & v3729844 | !jx0_p & v3a66998;
assign v373d203 = hmaster3_p & v374307e | !hmaster3_p & v3745473;
assign v3a6e721 = hgrant5_p & v37683bf | !hgrant5_p & v376592b;
assign v3a6f0a5 = hbusreq4 & v3762312 | !hbusreq4 & v3a5aacb;
assign v3775636 = hlock0 & v3755a05 | !hlock0 & v375c52f;
assign v3740212 = hmaster2_p & v8455ab | !hmaster2_p & v374821f;
assign v2ff8cae = hgrant4_p & v373ade9 | !hgrant4_p & v3768a37;
assign v376abdf = hbusreq5_p & v3a5e2c8 | !hbusreq5_p & v3a6a199;
assign v3a6f97f = hbusreq8_p & v373d449 | !hbusreq8_p & v3a554c5;
assign v3a6fe41 = hlock5_p & v8455ab | !hlock5_p & v37549cd;
assign v372cbdf = hmaster1_p & v3764a2c | !hmaster1_p & v3759c8c;
assign v3a61acf = hbusreq4_p & v3a672cb | !hbusreq4_p & v3761866;
assign v3a70bf3 = hmaster2_p & v3a6f130 | !hmaster2_p & v377e002;
assign v3a6fd3f = hlock5_p & v3a70922 | !hlock5_p & v37267f3;
assign v373cf4e = hbusreq1 & v8455ab | !hbusreq1 & !v373ad95;
assign v374b025 = hmaster0_p & v3a6e5f0 | !hmaster0_p & v3767e7e;
assign v372bc46 = hbusreq5_p & v3769d07 | !hbusreq5_p & !v373e6eb;
assign v3a708ee = hmaster0_p & v9d35e2 | !hmaster0_p & v377fad8;
assign v3745239 = hlock5_p & v3a71674 | !hlock5_p & v3724325;
assign v376fe88 = hbusreq6_p & v3747f5d | !hbusreq6_p & v377baeb;
assign v377a50f = hlock0 & v3754682 | !hlock0 & v3735051;
assign v373b671 = hbusreq0 & v376410a | !hbusreq0 & c7355c;
assign v374ce46 = hbusreq8_p & v376e113 | !hbusreq8_p & v3723686;
assign v374a9eb = hbusreq5_p & v3757c7d | !hbusreq5_p & !v372ab80;
assign v3734967 = hlock0_p & v3a68c1f | !hlock0_p & v3a66593;
assign v376aa98 = hbusreq4_p & v3a71617 | !hbusreq4_p & v3a63559;
assign v3724f4f = hbusreq5_p & v376fa43 | !hbusreq5_p & v376ce06;
assign v3a6f11c = hmaster0_p & v37517f4 | !hmaster0_p & d8c443;
assign v1e379cc = hbusreq5 & v3770366 | !hbusreq5 & v373c1ff;
assign v3a6f2f2 = stateG10_1_p & v8455ab | !stateG10_1_p & v377051a;
assign v3739732 = hgrant2_p & v377a9e7 | !hgrant2_p & v3772c57;
assign v376a941 = hmaster2_p & v3738253 | !hmaster2_p & v3766484;
assign v3730e98 = hbusreq1_p & v37749f0 | !hbusreq1_p & v8455ab;
assign v3a70d7a = hgrant2_p & v3a6ae68 | !hgrant2_p & v380761c;
assign v373cd8a = hbusreq5 & v3729cfa | !hbusreq5 & v37b64f8;
assign v3751aab = hbusreq8 & v3a70482 | !hbusreq8 & v3774bc0;
assign v37260fc = hmaster1_p & v8455e7 | !hmaster1_p & bc8871;
assign v376f4b9 = hlock8_p & v3a5cb20 | !hlock8_p & v376b063;
assign v376f1c0 = hbusreq4_p & b4ac83 | !hbusreq4_p & v373cf96;
assign v3a6f6e7 = hgrant3_p & v373ea3f | !hgrant3_p & v3a5e3bb;
assign v3a6faaa = hmaster1_p & v23fe361 | !hmaster1_p & v373385b;
assign v37626a4 = hgrant2_p & v373a568 | !hgrant2_p & v377c160;
assign v3771c5f = hmaster0_p & v37455ff | !hmaster0_p & v3735485;
assign v3777666 = hgrant6_p & v3750c38 | !hgrant6_p & v376005f;
assign v3774791 = hgrant6_p & v3747a53 | !hgrant6_p & v3734778;
assign v3767e76 = hbusreq0 & v376b4e1 | !hbusreq0 & !v8455ab;
assign v3752a7e = hgrant1_p & v8455ab | !hgrant1_p & !v372361c;
assign v37642e6 = hmaster0_p & v37434b2 | !hmaster0_p & !v3a6bc9a;
assign v3777631 = hbusreq8 & v375f5c1 | !hbusreq8 & v376e66e;
assign v377b27b = hbusreq2 & v37599cb | !hbusreq2 & v38072fd;
assign v3747816 = hmaster2_p & v3a6f443 | !hmaster2_p & !v3735e39;
assign v37552cb = hmaster0_p & v3a5af94 | !hmaster0_p & v3747737;
assign v375199d = hgrant4_p & v372b1e6 | !hgrant4_p & v3a70114;
assign v3741b5a = hgrant8_p & v3a7102a | !hgrant8_p & v3a5b6c8;
assign v3a592bc = hgrant5_p & v8455ab | !hgrant5_p & !v37763d1;
assign v37611c3 = hbusreq6 & v375aa2d | !hbusreq6 & v8455ab;
assign v373c21c = hbusreq0 & v372919a | !hbusreq0 & v8455ab;
assign a0715f = hlock5_p & v375345f | !hlock5_p & v8455ab;
assign v3779fd9 = hbusreq0 & v3755199 | !hbusreq0 & v3a581e4;
assign v3745f8d = hbusreq6_p & v376e040 | !hbusreq6_p & v3a6f3d5;
assign v375ff94 = hbusreq0 & v1e37339 | !hbusreq0 & v374518c;
assign v372dc5c = hbusreq2 & v3a6f70d | !hbusreq2 & v3a635ea;
assign v3761b3d = hbusreq2_p & v3a6cf5d | !hbusreq2_p & v374ad1e;
assign v377730a = hlock5_p & v375b97a | !hlock5_p & v373285d;
assign v3763dd4 = hmaster0_p & v3725bdc | !hmaster0_p & v3a70f44;
assign v37591b4 = hbusreq3 & v3a6f7bf | !hbusreq3 & v8455ab;
assign v377a887 = hmaster0_p & v3a619c0 | !hmaster0_p & v3a6f9ab;
assign v372d851 = hgrant2_p & v3774dbe | !hgrant2_p & v377ef47;
assign v374a510 = hgrant5_p & v377e493 | !hgrant5_p & v3a682f7;
assign v37738b2 = hmaster1_p & v3a66110 | !hmaster1_p & v376bc8c;
assign v23fdead = hlock5_p & v3a71509 | !hlock5_p & v37637d4;
assign v376ff61 = hbusreq3 & v373e5fb | !hbusreq3 & v372b5b0;
assign v3730fc4 = hmaster2_p & v3a58218 | !hmaster2_p & v37406d2;
assign v373fa33 = hgrant5_p & v8455c6 | !hgrant5_p & v3a61cd7;
assign v3a7021a = hbusreq7_p & v37610ce | !hbusreq7_p & v3a550e2;
assign v3a70cc7 = hbusreq5_p & v375f3ac | !hbusreq5_p & v373547f;
assign v3a5b42a = hbusreq2 & v3a6f806 | !hbusreq2 & v37453d7;
assign v3a6ee22 = hburst1 & v2aca977 | !hburst1 & v3a58cc0;
assign v374102a = hlock2_p & v37318da | !hlock2_p & v3763e88;
assign v3760681 = hmaster0_p & v3a70abe | !hmaster0_p & v3a70641;
assign v377aa5d = hmaster2_p & v373366b | !hmaster2_p & b66167;
assign v37592d0 = hmaster2_p & v37326a0 | !hmaster2_p & a34d2b;
assign v37601d6 = hbusreq6 & v374f754 | !hbusreq6 & v8455ab;
assign v3745e63 = hmaster3_p & v3a704e6 | !hmaster3_p & v375df4f;
assign v3a6fe5b = hbusreq0_p & v372dadb | !hbusreq0_p & v3a5a585;
assign v3747d30 = hmaster2_p & v373d219 | !hmaster2_p & v377baf4;
assign v3a6fe91 = hmaster0_p & v3764203 | !hmaster0_p & v3a71498;
assign v3772f3c = hbusreq8 & v3a6f356 | !hbusreq8 & v377e905;
assign v375ad9f = hmaster2_p & v39a5265 | !hmaster2_p & v3a70cc0;
assign v372bb0f = hmaster0_p & v372def3 | !hmaster0_p & !v3a56b7c;
assign v37299dc = hmaster0_p & v8455ab | !hmaster0_p & v3742efb;
assign v3738a94 = hmaster3_p & v3776c6b | !hmaster3_p & v37240c8;
assign v375ed60 = hmaster1_p & v3a71194 | !hmaster1_p & !v377167d;
assign v3a6f20d = hlock2 & v3a68463 | !hlock2 & v3a598a0;
assign v376455c = hgrant6_p & v8455ab | !hgrant6_p & v3752c99;
assign v3758e68 = hgrant2_p & v8455ab | !hgrant2_p & v373c99b;
assign v3a6632a = hlock0 & v3749d78 | !hlock0 & v374ba61;
assign v3777071 = hlock4 & v3a6f2ad | !hlock4 & v3a6e804;
assign v3a6ff8d = hmaster0_p & v376d9ad | !hmaster0_p & v37293f2;
assign v37606e5 = hlock4_p & v3739c30 | !hlock4_p & !v372c9ac;
assign v3a70286 = hbusreq2_p & d27546 | !hbusreq2_p & v376640b;
assign v3769215 = hmaster0_p & v3a58bb0 | !hmaster0_p & v37508b9;
assign v3777a7e = hbusreq2 & v3a6f5fb | !hbusreq2 & v8455ab;
assign v3a6968b = hbusreq2_p & v3744794 | !hbusreq2_p & v8455ab;
assign v376626a = hmaster0_p & v37334c5 | !hmaster0_p & v3742851;
assign v3a659d0 = hmaster2_p & v3a70b80 | !hmaster2_p & v37462e7;
assign v3723a00 = hgrant4_p & v3a7106e | !hgrant4_p & v372f2b7;
assign v3768636 = hbusreq8 & v3a570cd | !hbusreq8 & v376ec0d;
assign v3a5bc0a = hbusreq8 & v3a7031e | !hbusreq8 & v373e1cc;
assign v3a66ac0 = hgrant6_p & v372ffaa | !hgrant6_p & v375bc38;
assign v3a70011 = hlock1_p & v3735e39 | !hlock1_p & v376d856;
assign v3a7083e = hbusreq3 & v23fd7d9 | !hbusreq3 & v8455ab;
assign v3739ca8 = hbusreq2_p & v372c8d1 | !hbusreq2_p & !v8455ab;
assign v3740893 = hmaster2_p & v3a635ea | !hmaster2_p & v373ae83;
assign v372e562 = hbusreq0 & v376352a | !hbusreq0 & abddc4;
assign v3a6c908 = hbusreq5_p & v37c00f6 | !hbusreq5_p & v3a7122f;
assign v3741608 = hmaster1_p & v8455ab | !hmaster1_p & v35b7805;
assign v375a563 = hmaster0_p & v8455ab | !hmaster0_p & v3774882;
assign v374cc40 = hmaster2_p & v35772a6 | !hmaster2_p & !v3a56c66;
assign v3a714bd = hlock2_p & v3a68426 | !hlock2_p & v8455b7;
assign v377ec50 = hbusreq4 & v3a6ebfb | !hbusreq4 & v3a6bf41;
assign v3a70cec = hgrant4_p & v8455ab | !hgrant4_p & v3736aaa;
assign v375ebc3 = hbusreq5 & v376ffb4 | !hbusreq5 & v8455ab;
assign v3a66381 = hbusreq0 & v3a58e7f | !hbusreq0 & v3747178;
assign v376dea1 = hmaster0_p & v3728d9c | !hmaster0_p & v372f38e;
assign v3a5a258 = hbusreq6_p & v374b697 | !hbusreq6_p & v375c7d3;
assign v3745a5f = hbusreq4 & v39a537f | !hbusreq4 & v8455ab;
assign v3a702e7 = hbusreq4_p & v28896e3 | !hbusreq4_p & v3a705a9;
assign v3749f86 = hmaster2_p & v3a54aa0 | !hmaster2_p & v23fdd06;
assign v375314d = hgrant6_p & v37c039c | !hgrant6_p & v3a53c21;
assign v3a6fdb0 = hlock6 & v37391a1 | !hlock6 & v3a58530;
assign v3734534 = hmaster2_p & v3733da4 | !hmaster2_p & v3759f09;
assign v3745f4a = hlock3 & v3809b44 | !hlock3 & v3a6c672;
assign v3a711ac = hlock4_p & v374d99a | !hlock4_p & v3a5f20d;
assign v37765a3 = hlock0 & v3a70a7f | !hlock0 & v3738e63;
assign v37463ef = hmaster1_p & v3757261 | !hmaster1_p & v3a6fafb;
assign v23fe152 = hbusreq7 & v377f37e | !hbusreq7 & v376fff8;
assign v3777191 = hmastlock_p & v3a6cd1b | !hmastlock_p & !v8455ab;
assign v376f71a = hmaster1_p & v3723134 | !hmaster1_p & v3a70e0e;
assign v3763590 = jx0_p & v3a681f5 | !jx0_p & v8dc5a6;
assign v3762552 = hmaster0_p & v8455ab | !hmaster0_p & v375100c;
assign v375b239 = hbusreq7_p & v8455ab | !hbusreq7_p & v373c921;
assign v3764331 = hgrant5_p & v3724872 | !hgrant5_p & !v8455ab;
assign v3a58b20 = hgrant4_p & v8455ab | !hgrant4_p & v3a7167e;
assign v3a29a44 = hmaster0_p & v3a70051 | !hmaster0_p & v3758c58;
assign v3a5688f = hgrant2_p & v8455ab | !hgrant2_p & v3730b6d;
assign v3736cc7 = hbusreq3 & v3776b61 | !hbusreq3 & bdda12;
assign v37419fa = hmaster1_p & v3a6b1ab | !hmaster1_p & v3a63d05;
assign v3742e25 = hbusreq8 & v374bec2 | !hbusreq8 & v373d62f;
assign v3747586 = hmaster2_p & a568f8 | !hmaster2_p & !v372e0b0;
assign v3737186 = jx2_p & v3a6b478 | !jx2_p & v3736518;
assign v377baf4 = hgrant4_p & v8455ab | !hgrant4_p & v3809d8b;
assign v3777ca9 = hgrant0_p & v3a5a80c | !hgrant0_p & v3a65934;
assign v3a704a8 = hbusreq3 & v3732d4b | !hbusreq3 & !v8455ab;
assign v37576e7 = hbusreq5 & v37706ae | !hbusreq5 & v3a5e783;
assign v3730627 = hbusreq1_p & v37419a9 | !hbusreq1_p & v8455ab;
assign v3a6ffbe = stateG10_1_p & v8455ab | !stateG10_1_p & v3770548;
assign a36a2a = hlock3 & v377f149 | !hlock3 & v3a6c0b3;
assign v376b40c = hmaster0_p & v37640e9 | !hmaster0_p & v3761178;
assign v3742cd5 = hmaster0_p & v3a57672 | !hmaster0_p & v3757966;
assign v3a5ee85 = hbusreq5 & v374cfd9 | !hbusreq5 & v373d2e3;
assign v3776d72 = hmaster1_p & v3a647b8 | !hmaster1_p & v373a1dc;
assign v372fc77 = hbusreq2_p & v374e753 | !hbusreq2_p & v3a6fca5;
assign c6fb51 = hbusreq5_p & v3a7130f | !hbusreq5_p & !v8455ab;
assign v372d733 = hmaster1_p & v3a676c6 | !hmaster1_p & v37270dc;
assign v3730057 = hmaster0_p & v3a70bf6 | !hmaster0_p & v3a708e7;
assign v373ea19 = hmaster2_p & v38087c5 | !hmaster2_p & v8455ab;
assign v374e436 = hbusreq4 & v373de13 | !hbusreq4 & v3a71267;
assign v372ca99 = hmaster0_p & v3a5cc77 | !hmaster0_p & v3a70d93;
assign v3a70cea = hgrant3_p & v3a68aa8 | !hgrant3_p & v3a59351;
assign v37600c0 = hgrant4_p & v373828a | !hgrant4_p & !v374679f;
assign v39eb30a = hbusreq8_p & v3a6f634 | !hbusreq8_p & v37279dc;
assign v373ab4a = hbusreq2 & v3a6fa39 | !hbusreq2 & v8455ab;
assign v3a6f35c = hbusreq4_p & v377a606 | !hbusreq4_p & !v3a5dde0;
assign v3735abc = hmaster1_p & v37793e4 | !hmaster1_p & v3a70d7b;
assign v3a70938 = hmaster1_p & v37325c5 | !hmaster1_p & v3a6efb9;
assign v3a6ee78 = hbusreq6_p & v3748797 | !hbusreq6_p & v3a71131;
assign v3a5c25e = hlock4 & v3768723 | !hlock4 & v374d0f9;
assign v3732c0a = hmaster0_p & v3a6eef5 | !hmaster0_p & v3758ff0;
assign v3762f6e = hmaster0_p & v3776767 | !hmaster0_p & v8455ab;
assign v3764c9c = hlock0 & v3a6efad | !hlock0 & v3749008;
assign v3a70c04 = hbusreq5 & v3a67f13 | !hbusreq5 & v373a327;
assign v373bfdd = hlock7 & v3a6ffe2 | !hlock7 & v3768c76;
assign v372d8f9 = hbusreq4_p & v3771394 | !hbusreq4_p & !v8455ab;
assign v3745c20 = hbusreq8_p & v3a7008a | !hbusreq8_p & v1e37c44;
assign v3a5b12c = hbusreq2_p & v37431eb | !hbusreq2_p & v3773aa0;
assign v3a5db8a = hburst1 & v3757c6f | !hburst1 & v375f030;
assign v3a6ea51 = hbusreq1_p & v3a64566 | !hbusreq1_p & !v3a55b6c;
assign v3760e1b = hlock7 & v3a6f7c6 | !hlock7 & v3731f7f;
assign v372fb60 = hgrant6_p & v375b01a | !hgrant6_p & v376655b;
assign v23fe098 = hbusreq6_p & v3a5d90a | !hbusreq6_p & v3724ee0;
assign v372a683 = hmaster2_p & v3a635ea | !hmaster2_p & v3a567ec;
assign v3a65587 = hmaster1_p & v8455ab | !hmaster1_p & v2ff87d2;
assign v3767a42 = hgrant7_p & v37744e3 | !hgrant7_p & v373a79f;
assign v3748b43 = hmaster2_p & v3724394 | !hmaster2_p & v3a6b2c9;
assign v374270c = hmaster1_p & v3770b04 | !hmaster1_p & v3a70519;
assign v3734b80 = hbusreq6 & v3a66aa4 | !hbusreq6 & v35b774b;
assign v37404c5 = hmaster0_p & v376f5d9 | !hmaster0_p & v37654c4;
assign v3a6aabc = hbusreq4_p & v377349f | !hbusreq4_p & v37684a8;
assign v3a698c3 = hgrant2_p & v8455ba | !hgrant2_p & v37257c8;
assign v3752511 = hgrant3_p & v3a5f9f2 | !hgrant3_p & v3775a84;
assign dc571e = hbusreq7 & v375e0cc | !hbusreq7 & v8455ab;
assign v3a62396 = hbusreq1_p & v3a70672 | !hbusreq1_p & !v8455ab;
assign v3a5a3c7 = hbusreq2_p & v3a6f43e | !hbusreq2_p & v372935c;
assign v3a70481 = hbusreq4 & v3a70cb1 | !hbusreq4 & v3a6c5ee;
assign v3a6e7b3 = busreq_p & v376faea | !busreq_p & !v3a6841c;
assign v374b3b5 = hlock5_p & v3a6f336 | !hlock5_p & v376a863;
assign v3a669dc = hmaster1_p & v3733d3f | !hmaster1_p & v3a57c47;
assign v3776923 = hbusreq5_p & v3a70e45 | !hbusreq5_p & v3a60a9b;
assign v3736d58 = hmaster2_p & v3766d07 | !hmaster2_p & v372912f;
assign v37522a0 = hmaster0_p & v8455ab | !hmaster0_p & v3a6fa4d;
assign v37754f6 = hmaster0_p & v3a6f7dd | !hmaster0_p & v3757735;
assign v3732c72 = hbusreq2_p & v3a70635 | !hbusreq2_p & v8455b7;
assign v375b044 = hlock2 & v3a55bf6 | !hlock2 & v3a66051;
assign v38071bb = hmaster2_p & v3731857 | !hmaster2_p & !v3756f10;
assign v37523f4 = hbusreq2_p & v3a60618 | !hbusreq2_p & v37521af;
assign v374b228 = hmaster3_p & v3a6f5e7 | !hmaster3_p & v3748472;
assign v374a9db = hmaster1_p & v3a6f781 | !hmaster1_p & v3a58fa7;
assign v3a5e7a5 = hlock2_p & v3734af6 | !hlock2_p & v372c4c6;
assign v3a65552 = hbusreq5 & v3a6dc83 | !hbusreq5 & v377234d;
assign v3a5395c = hmaster0_p & v3737e2c | !hmaster0_p & v3a7074e;
assign v3750edc = hgrant4_p & v8455c2 | !hgrant4_p & v3732968;
assign v377028b = hgrant2_p & v8455ab | !hgrant2_p & v373193a;
assign v3748797 = locked_p & v2ff9190 | !locked_p & v8455ab;
assign v377bd5c = hbusreq4_p & v374612b | !hbusreq4_p & v8455ab;
assign v3743407 = hbusreq7_p & v3a634fa | !hbusreq7_p & !v3768d7e;
assign v3a644ac = hmaster3_p & v377cbb6 | !hmaster3_p & v3734a96;
assign v3771bed = hgrant0_p & v377682d | !hgrant0_p & !v3752e8e;
assign v3a707e7 = hmaster1_p & v3a663ef | !hmaster1_p & v375a754;
assign v3a71569 = hbusreq4 & cc4895 | !hbusreq4 & v375c70c;
assign v3726c5b = hlock6_p & v3725198 | !hlock6_p & v3a5b289;
assign v376a236 = hmaster1_p & v375af0b | !hmaster1_p & v3727f9c;
assign v373aeb3 = hbusreq4_p & v3a6fff0 | !hbusreq4_p & v3743393;
assign b038e6 = hbusreq4_p & v3727ee4 | !hbusreq4_p & v8455ab;
assign v3a698e1 = hbusreq7_p & v3a69ec5 | !hbusreq7_p & !v3a70333;
assign v3779b03 = hburst0 & v8455ab | !hburst0 & !v3a67851;
assign v3763498 = stateG10_1_p & v3a6f646 | !stateG10_1_p & v3a5db66;
assign v377824e = hbusreq2_p & v3764c4c | !hbusreq2_p & v3759512;
assign v374fd1f = hbusreq8_p & v3745e0d | !hbusreq8_p & v3a69239;
assign v377317d = hgrant4_p & v3a57b88 | !hgrant4_p & v377c4b7;
assign v374b887 = hgrant4_p & v8455c1 | !hgrant4_p & v37368e1;
assign v375ce98 = hbusreq4_p & v3722e5c | !hbusreq4_p & v35772a6;
assign v372362a = hmaster2_p & v376c2b7 | !hmaster2_p & !v3a632d8;
assign v3a6a051 = hlock6 & v3a714d2 | !hlock6 & v3723495;
assign v372ff6d = hmaster2_p & v380881d | !hmaster2_p & v3a5a8ce;
assign v3a5e2af = hbusreq8_p & v372e1bc | !hbusreq8_p & !v3768d8f;
assign v3a6fae3 = hmaster2_p & v8455e7 | !hmaster2_p & !v3a568f7;
assign v3733350 = stateG10_1_p & v35772a6 | !stateG10_1_p & !v373ae2e;
assign v377e27e = hmaster2_p & v3a70374 | !hmaster2_p & v377bbd9;
assign v37621d5 = hmaster0_p & v3a5a807 | !hmaster0_p & v3a66d14;
assign v376b0e6 = hgrant1_p & v3a57445 | !hgrant1_p & !v8455ab;
assign v3a63f43 = hgrant5_p & v373b71f | !hgrant5_p & v375ed43;
assign v37577a4 = hmaster2_p & v3763dd5 | !hmaster2_p & !v8455ab;
assign v3a5dad5 = hlock5_p & v3769093 | !hlock5_p & v374db8d;
assign v37435e1 = hmaster1_p & v3760690 | !hmaster1_p & v373ca9e;
assign v3722e4c = hbusreq2 & v3a6741a | !hbusreq2 & v3a6f949;
assign v375567c = hmaster1_p & v373d9e4 | !hmaster1_p & v3a62ad8;
assign v3a6e305 = hbusreq2_p & v3a6eb52 | !hbusreq2_p & !v3a68591;
assign v375842f = hmaster2_p & v3a635ea | !hmaster2_p & v373f0ee;
assign v3a70b3a = hbusreq3_p & v3749e48 | !hbusreq3_p & v3759947;
assign v3778ae9 = hmaster1_p & v377b24b | !hmaster1_p & v377cf4f;
assign v374597c = hmaster0_p & v3741249 | !hmaster0_p & v37358ab;
assign v3a7074d = hgrant4_p & v3776e5b | !hgrant4_p & v3a5417e;
assign v3a70f41 = hmaster2_p & v3777b00 | !hmaster2_p & v37745c3;
assign v372c00a = hbusreq7 & v3779b5b | !hbusreq7 & v375bfc4;
assign v3762b32 = hlock5 & v3723227 | !hlock5 & v373375c;
assign v377e319 = hmaster1_p & v3a7046c | !hmaster1_p & v3a706f4;
assign v3a6ae45 = hbusreq5_p & v3a70fd5 | !hbusreq5_p & v373c3e1;
assign v3732f19 = hmaster0_p & v373f9df | !hmaster0_p & v3a6f633;
assign v375f6f6 = hgrant1_p & v3750d37 | !hgrant1_p & !v8455ab;
assign v375fc0a = hgrant4_p & v3734292 | !hgrant4_p & v373df89;
assign v3a6bbe5 = hmaster2_p & v3755002 | !hmaster2_p & v8455ab;
assign a3d29c = hmaster2_p & v372d8e8 | !hmaster2_p & !v8455ab;
assign v372494a = hbusreq5 & v3763f13 | !hbusreq5 & v3806636;
assign v3762f2d = hbusreq8 & v3745e0e | !hbusreq8 & !v3768048;
assign v374ad96 = hbusreq6 & v3a6f018 | !hbusreq6 & !v3a5db8a;
assign v3a29856 = hbusreq7_p & v3732eaa | !hbusreq7_p & !v3a61b13;
assign v3a709cb = hgrant5_p & v35b774b | !hgrant5_p & v3a569dd;
assign v375aba9 = hlock5 & v3a57508 | !hlock5 & v375cf04;
assign v37506d6 = hbusreq4 & v376d488 | !hbusreq4 & v3741022;
assign v3761bd6 = hbusreq5_p & v3749381 | !hbusreq5_p & v3a6eec8;
assign v3a55640 = hgrant6_p & v376ea4a | !hgrant6_p & v37770d2;
assign v3809e25 = hgrant5_p & v8455ab | !hgrant5_p & v374caa8;
assign v3a6ff36 = hbusreq5_p & v375b046 | !hbusreq5_p & v3753d03;
assign v3a658b0 = hbusreq2_p & v3764994 | !hbusreq2_p & v374b4a4;
assign v3747fbc = hmaster2_p & d1bf3b | !hmaster2_p & v377957e;
assign v3728ae9 = hmaster1_p & v3a70c51 | !hmaster1_p & v3750113;
assign v373c1d7 = hbusreq2 & v3732b75 | !hbusreq2 & v377b774;
assign v8455bf = hlock3_p & v8455ab | !hlock3_p & !v8455ab;
assign v374249f = hbusreq6 & v374362e | !hbusreq6 & v8455ab;
assign v3759c49 = hbusreq6_p & v3a6f9c3 | !hbusreq6_p & v3a68967;
assign v3770c59 = hmaster2_p & v3a6908b | !hmaster2_p & v375ab02;
assign v3806a1c = hmaster1_p & v377854f | !hmaster1_p & v3736ded;
assign v3a6f043 = hbusreq4 & v37447e1 | !hbusreq4 & v377193a;
assign v3758357 = hbusreq8 & v3806df2 | !hbusreq8 & v3737808;
assign v374c801 = hbusreq6_p & v37610f8 | !hbusreq6_p & v3808eaa;
assign v375d84b = hlock0_p & v375fbd7 | !hlock0_p & v375bebd;
assign v37617ad = hbusreq4_p & v38072fd | !hbusreq4_p & v3a710dd;
assign v3a70094 = hgrant6_p & v374f557 | !hgrant6_p & !v3a61fcc;
assign v3a70209 = hbusreq6 & v3a71524 | !hbusreq6 & v8455ab;
assign v3756516 = hbusreq4_p & v377349f | !hbusreq4_p & v3a5bb4f;
assign v3737517 = hmaster1_p & v377d76b | !hmaster1_p & v372b813;
assign v3a672cb = hbusreq4 & v3763191 | !hbusreq4 & v35b774b;
assign v3728ced = hmaster0_p & v3a708e3 | !hmaster0_p & v3a553db;
assign v37736b4 = hbusreq5_p & v3a675dc | !hbusreq5_p & v374c9ab;
assign v3a680f4 = hbusreq6 & v3a55673 | !hbusreq6 & v3577376;
assign v3a705e8 = hlock0 & v38073c9 | !hlock0 & v3752002;
assign v37287d2 = hbusreq5 & v373666f | !hbusreq5 & v3a6542a;
assign v3a59d00 = jx1_p & v3a6f407 | !jx1_p & v3a6fa18;
assign v3767fa4 = hmaster1_p & v3a29a44 | !hmaster1_p & v3a70f10;
assign v37701a5 = jx0_p & v3a57dbb | !jx0_p & v377734d;
assign v3765370 = hbusreq0 & v3763186 | !hbusreq0 & v373f9ad;
assign v37521af = hbusreq2 & v380974c | !hbusreq2 & v8455b3;
assign v3761d5a = hbusreq6_p & v37474c2 | !hbusreq6_p & v3761eb6;
assign v3761b90 = hbusreq3_p & v3750d37 | !hbusreq3_p & !v3732dc6;
assign v376305d = hmaster2_p & v372d299 | !hmaster2_p & v3a69946;
assign v3a5f5ec = hlock7_p & v375bdd6 | !hlock7_p & v375b3b7;
assign v3764678 = hmaster1_p & v374e033 | !hmaster1_p & v3a59314;
assign v3a715e1 = hbusreq2_p & v3a5fc3c | !hbusreq2_p & v8455ab;
assign v3a71519 = stateA1_p & v3743bc5 | !stateA1_p & v3a70e3a;
assign v3730bd8 = hmaster2_p & v3a6a3e6 | !hmaster2_p & v374355e;
assign v3a70503 = hbusreq5_p & v373cd8a | !hbusreq5_p & !v3771e6d;
assign v3762bdf = hbusreq8 & v372cae4 | !hbusreq8 & v3a5f626;
assign v377bac7 = hlock8_p & v3a69da8 | !hlock8_p & !v3a69ec5;
assign v3a6fc9f = hmaster2_p & v39a5265 | !hmaster2_p & !v8455ab;
assign v3a5a591 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3770bf5;
assign v377ec9b = busreq_p & v3a703cf | !busreq_p & v3a6a187;
assign v3a633a7 = hbusreq6 & v377028b | !hbusreq6 & v377728d;
assign v2acb0b1 = hbusreq7_p & v3a704b3 | !hbusreq7_p & v374df3c;
assign v3751c77 = hbusreq4 & v374663d | !hbusreq4 & v3731230;
assign v373ddca = hbusreq2_p & v374074d | !hbusreq2_p & !v8455ab;
assign v374998d = hbusreq0 & v37264c9 | !hbusreq0 & v377e9d7;
assign v3742698 = hmaster2_p & v3a7151d | !hmaster2_p & !v3a7156d;
assign v3746d57 = hbusreq5_p & v377a13b | !hbusreq5_p & v3a57108;
assign v377ce96 = hgrant5_p & v3a6ff28 | !hgrant5_p & v3a6a8aa;
assign v373d239 = hgrant5_p & v3a579d1 | !hgrant5_p & v372d733;
assign v37444b2 = hgrant6_p & v373a013 | !hgrant6_p & v39eb532;
assign v3a6f0b8 = hbusreq6 & v3a676a9 | !hbusreq6 & v373fc8a;
assign v3a6f79f = hmaster0_p & v3743ff2 | !hmaster0_p & v3a66e30;
assign v3a56323 = hbusreq5_p & v37555b4 | !hbusreq5_p & v372de6f;
assign v377586c = hbusreq4 & v3a5e817 | !hbusreq4 & v37c0382;
assign v377cb2b = hbusreq6_p & v374f78c | !hbusreq6_p & v3a57836;
assign v376c1f7 = hbusreq4_p & v3740b8b | !hbusreq4_p & !v8455c2;
assign v373f2a6 = hmaster2_p & v3739ca5 | !hmaster2_p & v3a7007b;
assign v3772183 = hmaster0_p & v3a6a0a6 | !hmaster0_p & v377972c;
assign v376769e = hbusreq7 & v3763b4d | !hbusreq7 & v3723d79;
assign v3a6f81b = hmaster2_p & v3a67cff | !hmaster2_p & v375da82;
assign v3a712b9 = hbusreq8 & v3a56bb5 | !hbusreq8 & v8455ab;
assign v37776eb = hgrant5_p & ca32a1 | !hgrant5_p & v3a70a2c;
assign v3a5be70 = hmaster2_p & v3726c61 | !hmaster2_p & v37745a0;
assign v3a70025 = hbusreq6_p & v373325f | !hbusreq6_p & !v8455ab;
assign v3734de2 = hgrant5_p & v3774fee | !hgrant5_p & v375005c;
assign cc9e54 = hmaster3_p & v3778f32 | !hmaster3_p & v3778fae;
assign v337948a = hbusreq3_p & v372493b | !hbusreq3_p & !v3a6febd;
assign v372ab0f = hmaster0_p & v37565c3 | !hmaster0_p & v3774a9c;
assign v37328bf = hready & v3724994 | !hready & !v8455ab;
assign v3749caa = hbusreq2 & v3a6ab5f | !hbusreq2 & !v3a6ec7a;
assign v3a6c2df = hgrant6_p & a0503f | !hgrant6_p & v3a65b5d;
assign v3a5f711 = hmaster0_p & v37428b3 | !hmaster0_p & v375f014;
assign v3a70247 = hmaster1_p & v23fd9e7 | !hmaster1_p & v37289f0;
assign v373502a = hlock3 & v376be2c | !hlock3 & v3a66b2b;
assign v3741438 = hbusreq5 & v372571e | !hbusreq5 & v8455c7;
assign v3a706fe = hgrant4_p & v3743b9e | !hgrant4_p & v3a6bb84;
assign v3a61d67 = hbusreq5_p & v3756f41 | !hbusreq5_p & v3a5b3e6;
assign v3754a54 = hbusreq5 & v376b67d | !hbusreq5 & v3743d30;
assign v3a59bb4 = hbusreq2_p & v3a70e02 | !hbusreq2_p & v3a713c7;
assign v377e586 = hbusreq2 & v37718fb | !hbusreq2 & v8455ab;
assign v3a69dbd = hbusreq5 & v3a6d874 | !hbusreq5 & v3a6c5e5;
assign v3a602a4 = hbusreq4_p & v3775a4a | !hbusreq4_p & v375e64c;
assign v3a61302 = hbusreq5 & v3a62819 | !hbusreq5 & v3a70582;
assign v372e58c = hmaster2_p & v3752147 | !hmaster2_p & v3764cea;
assign v3736107 = hbusreq8 & v3756e87 | !hbusreq8 & v3752f15;
assign cceefd = hbusreq5_p & v3a6f66a | !hbusreq5_p & v372f93c;
assign v375a94a = hbusreq4_p & v374b077 | !hbusreq4_p & v374c95a;
assign v37648f2 = hlock0 & v373d10f | !hlock0 & v325b5df;
assign v3732cb4 = hgrant2_p & v8455e7 | !hgrant2_p & v1e3755f;
assign v375c771 = hgrant3_p & v377dd3b | !hgrant3_p & !v3a6f8dc;
assign v3765aa0 = hbusreq7 & v35b70ed | !hbusreq7 & v3a6a8ee;
assign v3a70319 = hbusreq2 & v3a7151d | !hbusreq2 & !v8455ab;
assign v374a67d = hlock4 & v3a552f7 | !hlock4 & v3a59dab;
assign v3725932 = hmaster2_p & v3730627 | !hmaster2_p & v8455ab;
assign v3724887 = hgrant2_p & v3a6fcc0 | !hgrant2_p & v3757598;
assign v375c32d = hbusreq8_p & v375ad7d | !hbusreq8_p & v8455ab;
assign v374e455 = hbusreq7_p & v3759fda | !hbusreq7_p & !v8455ab;
assign v3773e5f = hbusreq4_p & v376ddc6 | !hbusreq4_p & v37685bb;
assign v372b8d7 = hlock0 & v3760ff4 | !hlock0 & v3a70322;
assign v3741c3d = hmaster1_p & v3757966 | !hmaster1_p & v3742cd5;
assign v3728ca9 = hgrant0_p & v3a5b71a | !hgrant0_p & !v37381f0;
assign v3723fcc = hbusreq0 & v372c5da | !hbusreq0 & v372ff9a;
assign v375ea85 = hgrant4_p & v8455b0 | !hgrant4_p & v375b828;
assign v3a620d3 = hgrant6_p & v8455ab | !hgrant6_p & v376711c;
assign v374668d = hbusreq1 & v3a57309 | !hbusreq1 & v8455ab;
assign v3a6f2e5 = hbusreq5 & v376a94e | !hbusreq5 & v3749a06;
assign d7669b = hmaster0_p & v372aec7 | !hmaster0_p & v3774e4f;
assign v372754b = hmaster2_p & v3a62a6d | !hmaster2_p & !v37392ad;
assign v3754d21 = hgrant4_p & v8455ab | !hgrant4_p & v3a70c2e;
assign v3a5f413 = hgrant4_p & v3747c3e | !hgrant4_p & v8455ab;
assign v3a6eec8 = hbusreq5 & v372bdcf | !hbusreq5 & v3a6f1ea;
assign v3a6eb2d = hbusreq6_p & v373e933 | !hbusreq6_p & v8455b7;
assign v377038e = hmaster2_p & v372b231 | !hmaster2_p & v37229c2;
assign v3a5f76b = hmaster2_p & v3737478 | !hmaster2_p & v376a1dd;
assign v3724f9c = hbusreq3_p & v3a6cef4 | !hbusreq3_p & cf1ae7;
assign v37755ff = hmaster2_p & v3725f77 | !hmaster2_p & !v373e8ad;
assign v3a5cb0e = hbusreq5 & v37680a7 | !hbusreq5 & v3a63f9a;
assign v374d9b3 = hbusreq6 & v372fd12 | !hbusreq6 & v377bfc0;
assign v3a70990 = hbusreq5 & v376d9ad | !hbusreq5 & v373755a;
assign v3741d7c = hmaster1_p & v3756996 | !hmaster1_p & v3755508;
assign v3768e14 = hmaster1_p & v374fba1 | !hmaster1_p & v3740466;
assign v3a7045b = hlock6_p & v373621d | !hlock6_p & v37765fb;
assign v37381f0 = hlock0_p & v377c3fb | !hlock0_p & v374047d;
assign v3779227 = hlock2_p & v3779fb2 | !hlock2_p & v377613d;
assign v372cd8b = hgrant5_p & v3a6f290 | !hgrant5_p & v3a7164f;
assign v3770700 = hmaster0_p & v372ed51 | !hmaster0_p & v3a62d82;
assign v3760bda = hmaster0_p & v3a635ea | !hmaster0_p & v3a67c3b;
assign v3a67131 = jx3_p & v3769d3d | !jx3_p & v8455ab;
assign v3a6ad8b = hlock0_p & v3a66e91 | !hlock0_p & v376906d;
assign v3750978 = hbusreq3 & v39a5381 | !hbusreq3 & !v8455ab;
assign v37556ce = jx1_p & v3a6ecee | !jx1_p & v3a5d8f6;
assign v3a6776f = hbusreq5_p & v3770690 | !hbusreq5_p & v3779233;
assign a0503f = hbusreq6_p & v3a708a2 | !hbusreq6_p & v8455ab;
assign v3a7168b = hbusreq4 & v3577354 | !hbusreq4 & v3a5f9e6;
assign v37357d0 = hmaster0_p & v3a6f4d6 | !hmaster0_p & v8455ab;
assign v375babe = hmaster2_p & v37590d1 | !hmaster2_p & v3a54b46;
assign v374a3b2 = hgrant6_p & v8455ab | !hgrant6_p & v37531af;
assign v3772a57 = hmaster1_p & v376a4ec | !hmaster1_p & v37558f2;
assign v3a66538 = hgrant3_p & d284a6 | !hgrant3_p & v8455ab;
assign v3a70a3a = hmaster0_p & v376da3f | !hmaster0_p & !v3a610a4;
assign v375415d = hmaster0_p & v3a6ff25 | !hmaster0_p & v3732d3e;
assign v3a59d80 = hmaster1_p & v3a6906e | !hmaster1_p & v3774cc2;
assign v3a6912a = hgrant4_p & v3761e19 | !hgrant4_p & !d648e4;
assign v3a5618d = hbusreq0 & v3a6ffda | !hbusreq0 & v3a70d32;
assign v373f90a = hbusreq5 & v376a6f1 | !hbusreq5 & v3a6eb02;
assign v37792cf = hlock6 & v3a67b86 | !hlock6 & v3a69488;
assign v3758524 = hmaster2_p & v376b11e | !hmaster2_p & v23fd83f;
assign v375e8c1 = hmaster1_p & v375cab5 | !hmaster1_p & v3a70e72;
assign v3a706d2 = hlock0 & v3731230 | !hlock0 & v3753073;
assign v3752a0d = hlock0_p & v35b774b | !hlock0_p & v3753189;
assign v3a6fdea = hmaster2_p & v373aeb3 | !hmaster2_p & v3755417;
assign v3a5f07a = hgrant6_p & v3771b2c | !hgrant6_p & v372cfdf;
assign v3a636fe = hgrant6_p & v8455ca | !hgrant6_p & v373c423;
assign v37251b9 = hlock3 & v3a70dd0 | !hlock3 & a9f66a;
assign v375be25 = jx0_p & v3727b7f | !jx0_p & v3779c40;
assign v3742a61 = hbusreq5 & v23fdbe3 | !hbusreq5 & v3a67095;
assign v373d40c = hgrant5_p & v3769323 | !hgrant5_p & v3a6257d;
assign v374fa0a = hgrant0_p & v8455e7 | !hgrant0_p & !v372475a;
assign v3a5ea7b = hgrant0_p & v3779ea0 | !hgrant0_p & !v3a6b083;
assign v374f485 = hgrant3_p & v360d1cb | !hgrant3_p & v37296f0;
assign v3a6f834 = hbusreq8_p & v3740a8a | !hbusreq8_p & v3755066;
assign v9ae4c2 = hmaster0_p & v3a5687e | !hmaster0_p & v37328f1;
assign v37545a0 = hmaster2_p & v377bb3a | !hmaster2_p & v3724a4b;
assign v37395e6 = hbusreq3_p & v3740171 | !hbusreq3_p & v37270d9;
assign v3a70d44 = hlock0 & v376c76d | !hlock0 & v3a70336;
assign v3766ef7 = jx1_p & v3a6fe76 | !jx1_p & v3766f8a;
assign v3750f2a = hlock0_p & v3a708ec | !hlock0_p & c858c6;
assign v372e967 = hlock5 & v3a701b1 | !hlock5 & v2ff918d;
assign v3a54344 = hlock3_p & v3727ec9 | !hlock3_p & v37598c6;
assign v3a708ed = hmaster3_p & v373087c | !hmaster3_p & v377a0be;
assign v3a66e63 = hbusreq8 & v373d268 | !hbusreq8 & v3750fa9;
assign v3808f45 = hgrant6_p & v3770c9d | !hgrant6_p & v372d630;
assign v377762d = hgrant6_p & v375c7b9 | !hgrant6_p & v3a6b23f;
assign v375c70c = hgrant6_p & v374acbe | !hgrant6_p & v3767429;
assign v3a68825 = hbusreq7 & v377ef0b | !hbusreq7 & v373dafe;
assign v374f34b = hgrant7_p & v3768ba9 | !hgrant7_p & v376f2f4;
assign v39eb520 = hmaster0_p & v3762929 | !hmaster0_p & v3723e15;
assign v3a2986f = hbusreq5_p & v3a63f9a | !hbusreq5_p & v3777610;
assign v3a6f995 = hgrant4_p & v3a60787 | !hgrant4_p & v377a551;
assign c61447 = hbusreq3_p & v374cab9 | !hbusreq3_p & v376b509;
assign bbeeaf = hbusreq4_p & v8455bb | !hbusreq4_p & v3a65da7;
assign v37298f1 = hlock0 & v377bfc0 | !hlock0 & v3a5aaee;
assign v3a708f9 = hmaster1_p & v3746c51 | !hmaster1_p & v37269bf;
assign v3806a74 = stateA1_p & v8455ab | !stateA1_p & v373e80b;
assign v372fa17 = hmaster0_p & v8455e1 | !hmaster0_p & v3a6c933;
assign v3a7084f = hlock8 & v380937f | !hlock8 & v3739b6a;
assign v3a6ffe2 = hbusreq7 & v3a6fc94 | !hbusreq7 & v3a60859;
assign v375eac3 = hmaster0_p & v3746c51 | !hmaster0_p & v3a7161f;
assign v3a71273 = hmaster0_p & v3a709ee | !hmaster0_p & v37323a2;
assign v37796ce = hbusreq0 & v3a70765 | !hbusreq0 & v3770f54;
assign v3a7080b = hlock0 & v373484e | !hlock0 & v3a70405;
assign v374e401 = hbusreq5 & v37296f5 | !hbusreq5 & v8455bb;
assign v3733e1f = hlock5 & v3a70613 | !hlock5 & v3a6fb7f;
assign v375f9f1 = hlock5 & v3a70feb | !hlock5 & v3a58527;
assign v37583f0 = hmaster0_p & v3a6f550 | !hmaster0_p & v373185b;
assign v372dccf = hbusreq0_p & v373f06b | !hbusreq0_p & v8455ab;
assign v377849a = hmaster2_p & v3a6f42a | !hmaster2_p & !v376d86c;
assign v377b66a = hmaster2_p & v3a635ea | !hmaster2_p & v3779cf9;
assign v3743b98 = hbusreq4 & v3762072 | !hbusreq4 & v3a6ec0a;
assign v374284d = hbusreq0 & v37629b4 | !hbusreq0 & v38072fd;
assign v3a69949 = hbusreq5_p & v374943a | !hbusreq5_p & !v37552cb;
assign v377aed3 = hmaster3_p & v8455ab | !hmaster3_p & v37488d2;
assign v3a70a31 = hmaster0_p & v3a5e24e | !hmaster0_p & v3378a2d;
assign v373fede = hbusreq8_p & v375d20f | !hbusreq8_p & v37266d9;
assign v3762d5f = hlock2_p & v373712d | !hlock2_p & v8455b0;
assign v374bddc = hmaster2_p & v373ad2b | !hmaster2_p & v3737c0d;
assign v374172f = hbusreq2 & v373502a | !hbusreq2 & v373f0ee;
assign v3736bcd = hlock4 & v375c3a2 | !hlock4 & v3a6f709;
assign v372af30 = hbusreq2 & v3755002 | !hbusreq2 & v8455ab;
assign v3757ca4 = hmaster0_p & v3735d6f | !hmaster0_p & !v3a5a807;
assign v3a6a075 = hbusreq2_p & v3a63805 | !hbusreq2_p & v8455b0;
assign v375e30f = hmaster0_p & v377ef09 | !hmaster0_p & v373ec8f;
assign v37689aa = hmaster3_p & v3a5aa64 | !hmaster3_p & v3a6c5ed;
assign v3756e20 = hmaster2_p & v373195f | !hmaster2_p & a39369;
assign v37663b5 = hbusreq6_p & v3a715e3 | !hbusreq6_p & v8455ab;
assign v372efbe = hgrant3_p & v8455e7 | !hgrant3_p & v372f85e;
assign v376f8bf = hbusreq0 & v3a62082 | !hbusreq0 & v37480fe;
assign v373f06b = locked_p & v8455ab | !locked_p & v3745f76;
assign v3724e2a = hbusreq4 & v374dffc | !hbusreq4 & v373abde;
assign v3a6f6e1 = hbusreq7_p & v375c9a3 | !hbusreq7_p & v37335a5;
assign v373af21 = hbusreq4_p & v3740e5a | !hbusreq4_p & v372eeda;
assign v37722e5 = hbusreq6_p & v3a662c7 | !hbusreq6_p & v377c671;
assign v3a715f8 = hgrant5_p & v8455ab | !hgrant5_p & v3a6d926;
assign v3759c5d = hgrant3_p & v3728b2f | !hgrant3_p & v37401f0;
assign v376f661 = hbusreq2_p & v37c0190 | !hbusreq2_p & v3779e66;
assign v37501f3 = hgrant6_p & v8455ab | !hgrant6_p & v3a5846c;
assign v3733e30 = hmaster0_p & v3775d26 | !hmaster0_p & !v372cdd5;
assign v37685fe = hmaster1_p & v3726ea3 | !hmaster1_p & v3774399;
assign v3761769 = hmaster2_p & v3a5f6d5 | !hmaster2_p & v375518f;
assign v3a6ffcf = hbusreq3 & v3a6772f | !hbusreq3 & v3a68523;
assign v373ec98 = hbusreq4_p & v3758187 | !hbusreq4_p & v3a55584;
assign v3a7005f = hbusreq0 & v3a702e1 | !hbusreq0 & v3a70088;
assign v37742c5 = hbusreq7_p & v373aa76 | !hbusreq7_p & !v3a6c9c7;
assign v3a705ea = hmaster1_p & v3a6f6c0 | !hmaster1_p & v3777da6;
assign v3a6fd91 = hgrant6_p & v374233c | !hgrant6_p & v3779cb7;
assign v3730e4c = jx0_p & v374c885 | !jx0_p & v377b209;
assign v376ace9 = hbusreq3_p & v3a70a6f | !hbusreq3_p & v3764dc2;
assign v2092f20 = hgrant0_p & v376866e | !hgrant0_p & !v373b0e5;
assign v3756263 = hmaster0_p & v3a715fc | !hmaster0_p & v3a6ef7f;
assign v37656ec = hburst1 & v8455ab | !hburst1 & v3a6f909;
assign v37538e4 = hgrant3_p & v360d1cb | !hgrant3_p & v3730cda;
assign v39a4db0 = hgrant3_p & v38070c1 | !hgrant3_p & v3a66476;
assign v3736968 = hbusreq4_p & v377a9cb | !hbusreq4_p & v37721e3;
assign v376fe00 = hgrant5_p & v8455ab | !hgrant5_p & v3a706de;
assign v3771e23 = hmaster2_p & v3a708c6 | !hmaster2_p & v3a60a32;
assign v37325b9 = hbusreq7 & v376910a | !hbusreq7 & v3761351;
assign v3a6eb7d = hbusreq5_p & v3a6fd66 | !hbusreq5_p & v374fe63;
assign v3a70b11 = hready_p & v3749293 | !hready_p & v373c553;
assign v3725bba = hbusreq5 & v3766160 | !hbusreq5 & v9ae4c2;
assign v377327b = hlock2_p & v1e37dd9 | !hlock2_p & v377c7b2;
assign v372874e = hmaster1_p & v376c3fd | !hmaster1_p & v374fc17;
assign v37551b0 = hmaster0_p & v3724394 | !hmaster0_p & v3a714b4;
assign v373bbb4 = hbusreq5_p & v37316ec | !hbusreq5_p & !v8455ab;
assign v3a63bb7 = hbusreq0 & v3753dab | !hbusreq0 & v8455ab;
assign v39eb56d = hbusreq8 & v3a62027 | !hbusreq8 & v8455ab;
assign v3a6724f = hgrant5_p & v3a60cf8 | !hgrant5_p & v3a551e2;
assign v3742d37 = hgrant3_p & v8455ab | !hgrant3_p & !v8455e9;
assign v3a62a14 = hmaster1_p & v3778484 | !hmaster1_p & v37242b9;
assign v2093005 = jx1_p & v3a70dad | !jx1_p & v8455ab;
assign v3a60bc1 = hmaster1_p & v3a62542 | !hmaster1_p & v3a5c066;
assign v374ccb3 = hgrant4_p & v1e37b99 | !hgrant4_p & !v3a7119f;
assign v37366d0 = hlock0_p & v3a70641 | !hlock0_p & v3766c8c;
assign v37327c5 = hmaster2_p & v8455ca | !hmaster2_p & ae317f;
assign v372e36d = hmaster0_p & v376142c | !hmaster0_p & v37509a9;
assign v3740f65 = hmaster0_p & v3a706a1 | !hmaster0_p & v37660f2;
assign a5c619 = hbusreq8 & v376b7ff | !hbusreq8 & v3762100;
assign v37724db = hlock4 & v372fecf | !hlock4 & v3741338;
assign v3a70de5 = hbusreq7 & v374a79e | !hbusreq7 & v372863f;
assign v3a71658 = hmaster0_p & v3a6e130 | !hmaster0_p & v374e519;
assign v37746d7 = hbusreq1_p & v3a700da | !hbusreq1_p & !v8455ab;
assign v3a6f5fb = hbusreq3_p & v373d78b | !hbusreq3_p & v3a6fcb9;
assign v3739062 = hbusreq2_p & v374fd8d | !hbusreq2_p & v373125c;
assign v374f0c1 = busreq_p & v3732a41 | !busreq_p & !v37687ce;
assign v3a6f38c = hbusreq6 & v3a6a075 | !hbusreq6 & v8455ab;
assign v3a55491 = hmaster1_p & v3a6f86a | !hmaster1_p & v374975c;
assign v375c791 = hgrant4_p & v3a61a7f | !hgrant4_p & v3a538b9;
assign v23fda7e = hmaster0_p & v8455b0 | !hmaster0_p & v3a710b4;
assign v375f169 = hbusreq4 & v375139d | !hbusreq4 & !v37706b3;
assign v372c500 = hgrant2_p & v3a70b92 | !hgrant2_p & v37730bf;
assign v3a70cdd = hgrant6_p & v377f09a | !hgrant6_p & v3730646;
assign v3a67284 = hgrant3_p & v8455ab | !hgrant3_p & v372aa99;
assign v377f865 = hlock4_p & v3a607af | !hlock4_p & v373aaa8;
assign v937864 = hmaster2_p & v3a6ef50 | !hmaster2_p & v209310e;
assign v3a6f2a2 = hbusreq0_p & v375e309 | !hbusreq0_p & v8455b5;
assign v3a70b6e = hgrant3_p & v8455be | !hgrant3_p & v3a66dcf;
assign v37551ec = hbusreq0 & v37717a4 | !hbusreq0 & v8455ab;
assign v3770651 = hgrant3_p & v8455ab | !hgrant3_p & v375ed5a;
assign v3758c06 = hgrant6_p & v8455ab | !hgrant6_p & v3747276;
assign v3728b1d = hbusreq8_p & v375e737 | !hbusreq8_p & d70cde;
assign v3768ac9 = jx0_p & v37370a1 | !jx0_p & v3726efd;
assign v3258760 = hmaster1_p & v376c0a0 | !hmaster1_p & v376c590;
assign v3735eb8 = hbusreq2 & v37652a5 | !hbusreq2 & v39ea7a8;
assign v3a70334 = hgrant1_p & v3a6f4d3 | !hgrant1_p & v3a6f436;
assign v3a58ea7 = hlock4_p & v37315da | !hlock4_p & v3a708a2;
assign v3a7013d = hbusreq7 & v374f6a4 | !hbusreq7 & v8455bb;
assign v3a53fb5 = hbusreq5_p & v35b7771 | !hbusreq5_p & v373f4a9;
assign v377609f = hmaster2_p & v37245f8 | !hmaster2_p & v3a6fdd6;
assign v37302c5 = hlock6 & v373a493 | !hlock6 & cf45c3;
assign v3730e75 = hmaster2_p & v3a57584 | !hmaster2_p & !v3a7101b;
assign v37572eb = hmaster3_p & v3a712b5 | !hmaster3_p & v360d01e;
assign v3a6f91e = hbusreq4_p & v3a58d22 | !hbusreq4_p & !v3a70025;
assign v3a5491d = hmaster2_p & v3775a29 | !hmaster2_p & v3728d9c;
assign v3a6feb9 = hgrant3_p & v8455e7 | !hgrant3_p & !v1e37a69;
assign v3a65b4a = hbusreq4_p & v376f56d | !hbusreq4_p & v3773650;
assign v3a5614c = hbusreq1_p & v3a6d749 | !hbusreq1_p & !v8455ab;
assign v3a6f333 = hlock1 & v37722cc | !hlock1 & v372ab85;
assign v3731974 = hmaster1_p & v3a6373e | !hmaster1_p & v376d896;
assign v3750b9e = hgrant2_p & v2092ac0 | !hgrant2_p & v376f661;
assign v37345aa = hmaster2_p & v2ff8bbc | !hmaster2_p & v3a6eb7b;
assign v3a6ac17 = hmaster2_p & v9ed516 | !hmaster2_p & v8455ab;
assign v372a023 = stateA1_p & v3a6ac94 | !stateA1_p & v3a71137;
assign v3a70704 = hlock4 & v377f171 | !hlock4 & a9c905;
assign v3737103 = hmaster1_p & v8455ab | !hmaster1_p & v3737a06;
assign v3a67f31 = hbusreq4 & v372ca2a | !hbusreq4 & v8455ab;
assign v377244a = hbusreq7_p & v3759421 | !hbusreq7_p & v37770ab;
assign v3a55a58 = hbusreq5_p & v3a55d4c | !hbusreq5_p & v375a804;
assign v3a56197 = hmaster1_p & v375c94e | !hmaster1_p & v3773dc6;
assign v3769759 = hgrant8_p & v8455ab | !hgrant8_p & !v377b074;
assign v374f7f8 = hmaster3_p & v372ad5a | !hmaster3_p & !v3a70657;
assign v3a57be6 = hmaster1_p & v377c7c0 | !hmaster1_p & v3768064;
assign v377918a = hmaster2_p & v3a5b8b9 | !hmaster2_p & v380881d;
assign v374d970 = hbusreq0 & v3a70966 | !hbusreq0 & v377e512;
assign abd043 = hmaster0_p & v3744af9 | !hmaster0_p & v3a6cf7f;
assign v3a6fef1 = hbusreq4_p & v3a5e55e | !hbusreq4_p & v3a5fc8d;
assign v3a615c8 = hgrant6_p & v3a70b9e | !hgrant6_p & v3757ec8;
assign ae6485 = hbusreq1_p & v373dcb0 | !hbusreq1_p & v373d8c0;
assign v377a62e = hmaster0_p & v3730f7e | !hmaster0_p & !v377624b;
assign v3771b2a = hbusreq8_p & v3a70fad | !hbusreq8_p & v376d9ed;
assign v3a70cdb = hbusreq1_p & v3a67a06 | !hbusreq1_p & v8455ab;
assign v3733027 = hbusreq4_p & v374c53a | !hbusreq4_p & v3778567;
assign v3a5b6c8 = hgrant7_p & v3a6eaf7 | !hgrant7_p & v374bdcb;
assign v3a670fe = hbusreq2 & a36a2a | !hbusreq2 & v3a7162d;
assign v377bbbd = hlock4 & v3a70c10 | !hlock4 & v3a62c49;
assign v3a6ad00 = hbusreq0 & v3a7022e | !hbusreq0 & v3a71092;
assign v3774c11 = hgrant1_p & v3a53877 | !hgrant1_p & v8455e7;
assign v372c944 = hbusreq6 & v376c4c5 | !hbusreq6 & v373f492;
assign v37588cf = hmaster0_p & v3773f26 | !hmaster0_p & v37445ff;
assign v377e692 = hmaster2_p & v372b881 | !hmaster2_p & v3722bca;
assign v3a6f9ca = hbusreq3 & v3a6fcb9 | !hbusreq3 & v8455ab;
assign v373bf3c = hbusreq4 & v1e3795b | !hbusreq4 & v8455ab;
assign v3a66545 = hbusreq4_p & v3a620d3 | !hbusreq4_p & v3a6bf89;
assign v374d836 = hlock1 & v375bd8a | !hlock1 & v377836a;
assign v373913a = hbusreq2_p & v3753ca0 | !hbusreq2_p & v3a6d37f;
assign v3a6ff28 = hmaster1_p & v3736ef2 | !hmaster1_p & v373afd5;
assign v375874f = hmaster0_p & v376d9ad | !hmaster0_p & v373da7d;
assign v3a70a75 = hmaster0_p & v3a635ea | !hmaster0_p & v3769e50;
assign v375634b = hmaster1_p & v3773697 | !hmaster1_p & v3759501;
assign v3a6fb53 = jx0_p & v3a682e5 | !jx0_p & v375377b;
assign v3a59de6 = hmaster0_p & v372fd00 | !hmaster0_p & v3768c25;
assign v37255f6 = hmaster0_p & v3a6b597 | !hmaster0_p & v37744d9;
assign v3775f25 = hmaster2_p & v374cfee | !hmaster2_p & v3a55395;
assign v3758225 = hgrant1_p & v3a5e9d3 | !hgrant1_p & v3a5ce2d;
assign v373300a = hbusreq5_p & v3742649 | !hbusreq5_p & v372ebc8;
assign v3758950 = hbusreq2 & v37796c6 | !hbusreq2 & v8455ab;
assign v372a0e3 = hmaster0_p & v377e298 | !hmaster0_p & v3a6adff;
assign v3a7125d = hlock8 & v3a574d7 | !hlock8 & v373db82;
assign v3744aed = hgrant6_p & v376a040 | !hgrant6_p & !v3744dc6;
assign v3a61e95 = hbusreq5_p & v372b164 | !hbusreq5_p & !v8455ab;
assign v3747b29 = hmaster2_p & v2092faa | !hmaster2_p & v3a6a213;
assign v3a69488 = hgrant2_p & v37682c0 | !hgrant2_p & v3739f22;
assign v377e19d = hgrant4_p & v373c21c | !hgrant4_p & v375c1df;
assign v3a6fcdf = hmaster1_p & v3726ddb | !hmaster1_p & v8455c6;
assign v3741f22 = hbusreq6_p & v377b2b6 | !hbusreq6_p & v375ced9;
assign v37560f7 = hlock6_p & v3a653e4 | !hlock6_p & !v8455ab;
assign v3734fc3 = hmaster0_p & v375d4de | !hmaster0_p & v3a5ae95;
assign v3a6867e = hbusreq6 & v376e25b | !hbusreq6 & v3a70d99;
assign v37501ad = hbusreq6 & v3a6f49e | !hbusreq6 & v373b687;
assign v3a704ea = hbusreq4 & v377af09 | !hbusreq4 & v3727084;
assign v3a7160d = hmaster2_p & v3a70374 | !hmaster2_p & v375c903;
assign v3772117 = hgrant3_p & v8455ab | !hgrant3_p & v3723d55;
assign v3758c65 = hgrant4_p & v3a6f32d | !hgrant4_p & !v37739c6;
assign v3773712 = hmaster1_p & v376d883 | !hmaster1_p & !v3a55d78;
assign v3746d31 = hlock5_p & v3a6f92f | !hlock5_p & !v3a6572c;
assign v3a6bf05 = hlock5_p & v376583c | !hlock5_p & v3a6faff;
assign v375d7d2 = hlock7 & v3a6673e | !hlock7 & v3a704f5;
assign v376bfc3 = hgrant2_p & v3a702f8 | !hgrant2_p & v8455ab;
assign v376c1de = hbusreq4_p & v372ff70 | !hbusreq4_p & v8455ab;
assign v3745196 = hmaster3_p & v3a5fd54 | !hmaster3_p & v3769c51;
assign v3a5b01a = hmaster1_p & v3a6fd4f | !hmaster1_p & v3772e4f;
assign v35b70e6 = hgrant3_p & v377dd3b | !hgrant3_p & v37598c6;
assign v374b3f8 = hgrant4_p & v3a5b1ec | !hgrant4_p & v3778a8b;
assign v292554f = hmaster0_p & v3756a6a | !hmaster0_p & v375d2b3;
assign v3727165 = hbusreq1_p & v37368df | !hbusreq1_p & v376cf85;
assign v373d381 = hmaster0_p & v3a637dc | !hmaster0_p & v3a709d9;
assign v372c9ac = hgrant3_p & v3760bf8 | !hgrant3_p & v1e379fe;
assign v3a6f62f = hbusreq5_p & v372416d | !hbusreq5_p & !v374e34d;
assign v380a20c = hmaster3_p & v3a6ff68 | !hmaster3_p & v3a5e0dd;
assign v373790d = hmaster0_p & v8455ab | !hmaster0_p & v3a6a19b;
assign v372c4c6 = hbusreq2 & v8455ab | !hbusreq2 & !v373ad95;
assign v3a7045d = hmaster0_p & v372e250 | !hmaster0_p & v3737721;
assign v3a5d94a = hbusreq4 & v37674c1 | !hbusreq4 & !v8455ab;
assign v377f6af = hbusreq7 & v3a64aa2 | !hbusreq7 & a18d54;
assign v3a6ba54 = hbusreq7 & v376f319 | !hbusreq7 & !v8455ab;
assign v372b164 = hbusreq5 & v376f56d | !hbusreq5 & v374a11d;
assign v3775642 = hbusreq2_p & v375e2d3 | !hbusreq2_p & v3766709;
assign v373bde3 = hlock4 & v3a6bbf0 | !hlock4 & v3772404;
assign v3746e94 = hmaster0_p & v374c78e | !hmaster0_p & v3a6c03d;
assign v375facf = hmaster1_p & v3a6e7ce | !hmaster1_p & !v373b7dd;
assign v3a70bde = hgrant6_p & v8455ab | !hgrant6_p & v375000b;
assign v3a6d930 = hmaster0_p & v3a7002c | !hmaster0_p & v3736613;
assign v373fc36 = hmaster2_p & v3a55ee6 | !hmaster2_p & v3743434;
assign v373f159 = hbusreq4_p & v377a9e7 | !hbusreq4_p & !v3747623;
assign v373cc0f = hgrant4_p & v8455ab | !hgrant4_p & v37293ea;
assign v3765aee = hmaster2_p & v3a6d590 | !hmaster2_p & v375f61e;
assign v3749cf7 = hbusreq4 & v377caa3 | !hbusreq4 & v8455bf;
assign v37535f2 = hgrant2_p & v8455ab | !hgrant2_p & v3a62d36;
assign v3a70a53 = jx0_p & v3773536 | !jx0_p & v8455ab;
assign v3744cf1 = hgrant5_p & v375d43d | !hgrant5_p & v3a5e035;
assign v8455b0 = hready & v8455ab | !hready & !v8455ab;
assign v3a56d04 = hmaster0_p & v3a5b46d | !hmaster0_p & !v8455e7;
assign v31c369c = hgrant6_p & v8455ab | !hgrant6_p & v3a7126c;
assign v375e767 = hbusreq5 & v3a7086d | !hbusreq5 & v375329c;
assign v3757dd4 = hbusreq7 & v37464f3 | !hbusreq7 & v3a6c15c;
assign v373ab7e = hbusreq5_p & v374f0af | !hbusreq5_p & !v8455ab;
assign v375fea8 = jx0_p & v3a6982f | !jx0_p & v3a6a156;
assign v372df2a = hbusreq6 & v37583be | !hbusreq6 & v376b4e1;
assign v373f940 = hmaster0_p & v375d92e | !hmaster0_p & v376730a;
assign v3a55dc3 = hbusreq0 & v3744999 | !hbusreq0 & v3a711b2;
assign v372f441 = hmaster0_p & v376cbbe | !hmaster0_p & !v375fb03;
assign v3a709d9 = hmaster2_p & v3a637dc | !hmaster2_p & v3a637dd;
assign v374a795 = jx0_p & v373f5b1 | !jx0_p & v3807d51;
assign v3734e70 = hlock7 & v3743b63 | !hlock7 & v3731f35;
assign v373df82 = hmaster2_p & v3767561 | !hmaster2_p & v3a5e7fe;
assign v3757e71 = hbusreq7_p & v3a70cb4 | !hbusreq7_p & v3752a6c;
assign v3a67fee = hmaster1_p & v8455ab | !hmaster1_p & v3a7049e;
assign v3a5dd98 = hbusreq8_p & v3a705d3 | !hbusreq8_p & v3a7075c;
assign v374c1a0 = hmaster0_p & v3a582c5 | !hmaster0_p & v3755670;
assign v373f125 = hgrant6_p & v8455ab | !hgrant6_p & v3779337;
assign v374518b = hgrant6_p & v8455ab | !hgrant6_p & v3749caf;
assign v3738510 = hbusreq3_p & v3731eb8 | !hbusreq3_p & v8455ab;
assign v372b9e9 = hmaster2_p & v35772a2 | !hmaster2_p & v3a67967;
assign v374502e = hburst1 & v3771ce2 | !hburst1 & v374d037;
assign v3763da5 = hmaster2_p & v3a635ea | !hmaster2_p & v3a706fe;
assign v3776d4b = hbusreq7_p & a0a219 | !hbusreq7_p & v373121b;
assign v375cce7 = hmaster3_p & v374a36a | !hmaster3_p & v37750e0;
assign v372dddc = hbusreq3_p & v377af98 | !hbusreq3_p & v375f30d;
assign v3a6f8d9 = hbusreq5_p & v38094b8 | !hbusreq5_p & v373e873;
assign v375c4a1 = hgrant0_p & v376102a | !hgrant0_p & v377ae9c;
assign v3a6ef55 = hmaster3_p & v3a70c18 | !hmaster3_p & v3a7058c;
assign v372977b = jx0_p & v3a69a00 | !jx0_p & v39ea2e3;
assign v376d566 = hgrant6_p & v8455ca | !hgrant6_p & v3a711c1;
assign v3730cb5 = hlock7_p & v3728ac4 | !hlock7_p & !v8455ab;
assign v3777d70 = hgrant5_p & v8455c6 | !hgrant5_p & v3769740;
assign v374c582 = hmaster2_p & v8455ab | !hmaster2_p & v372eff2;
assign v3a70cd7 = hbusreq7 & v3a70f92 | !hbusreq7 & v3779d96;
assign v373b16e = hmaster2_p & v376a14f | !hmaster2_p & v3806db7;
assign v3750e8a = hbusreq7_p & v372dc2b | !hbusreq7_p & v3a6a64f;
assign v3a58219 = hbusreq8 & v372b721 | !hbusreq8 & a0a219;
assign v37362ff = hmaster2_p & v3755002 | !hmaster2_p & v3723eef;
assign v373e38a = hgrant4_p & v3a65d01 | !hgrant4_p & v374e768;
assign v372b0f9 = hbusreq3_p & v37714e6 | !hbusreq3_p & v3a70cdf;
assign v373dafe = hgrant5_p & v8455ab | !hgrant5_p & v3a6cdcd;
assign v3763c82 = hgrant3_p & v3734967 | !hgrant3_p & aef136;
assign v3759dda = hbusreq1_p & v3742034 | !hbusreq1_p & v8455ab;
assign v3747210 = hmaster1_p & v377c15d | !hmaster1_p & v372ce29;
assign v375265e = hbusreq4 & v3a6b94f | !hbusreq4 & v8455ab;
assign v377f7e1 = hbusreq6_p & v3a6f898 | !hbusreq6_p & v3a6fe71;
assign v3745069 = hbusreq6 & v372b1ed | !hbusreq6 & v3754940;
assign v374f44c = hmaster0_p & v37758d0 | !hmaster0_p & v8455ab;
assign v3a5b514 = hmaster0_p & v374093f | !hmaster0_p & d54152;
assign v3744c10 = hgrant4_p & v373f159 | !hgrant4_p & v37266c6;
assign v37429a1 = hgrant4_p & v8455ab | !hgrant4_p & v3a5741c;
assign v373427f = hgrant4_p & v3a708c2 | !hgrant4_p & v37519ea;
assign v374a8e2 = hmaster0_p & v374aabf | !hmaster0_p & v8455ab;
assign v374b759 = hmaster2_p & v3a70464 | !hmaster2_p & v377a356;
assign v375eb97 = hbusreq2 & v3a607af | !hbusreq2 & v8455ab;
assign v372dd4b = hbusreq5_p & v3a56794 | !hbusreq5_p & v3762b32;
assign v3a6eba3 = hbusreq0 & v3730043 | !hbusreq0 & v3808cf1;
assign v373af66 = hmaster2_p & v3a6f4c3 | !hmaster2_p & v3747787;
assign v3a6fa0d = hbusreq2_p & v374f29f | !hbusreq2_p & v3735354;
assign v373ba2e = hlock5 & v3a6fb69 | !hlock5 & v37675e9;
assign v3a68f98 = hlock6 & v372d4de | !hlock6 & v3a6f20d;
assign v375de2d = hbusreq6_p & v2889716 | !hbusreq6_p & v3735f7a;
assign v3a658be = hlock2_p & v3a6f96f | !hlock2_p & v8455b0;
assign v3726826 = hbusreq5_p & v37570f8 | !hbusreq5_p & v377437d;
assign v3a6cd87 = hbusreq5_p & v37706ef | !hbusreq5_p & v8455ab;
assign v2092a7a = hbusreq5 & v1e37cd7 | !hbusreq5 & v3766ff3;
assign v375791b = hbusreq0 & v374e19c | !hbusreq0 & v37404b3;
assign v37782a8 = hmaster1_p & v3a556ab | !hmaster1_p & v8455ab;
assign v37710f3 = hmaster1_p & aed6c7 | !hmaster1_p & v37350b2;
assign v3777178 = hgrant6_p & v8455ab | !hgrant6_p & v3a706a2;
assign v375c4c7 = hmaster1_p & v3a29520 | !hmaster1_p & v3a69a1b;
assign v3a5df97 = hbusreq3 & v3a5e817 | !hbusreq3 & v37c0382;
assign v377f037 = jx0_p & v374b589 | !jx0_p & v3762e7a;
assign v38088b6 = hbusreq5 & v3736d0d | !hbusreq5 & v3a58c07;
assign v373d076 = hmaster2_p & v374f707 | !hmaster2_p & v3759b63;
assign v3a6fba6 = hgrant6_p & v3a710f1 | !hgrant6_p & v3a714a2;
assign v374d7fc = hbusreq8 & v37234d5 | !hbusreq8 & !v8455ab;
assign v375fb93 = hmaster2_p & v8455b5 | !hmaster2_p & !v8455ab;
assign v3779e66 = hgrant3_p & v8455bd | !hgrant3_p & v373d932;
assign v3772083 = hbusreq5 & v374c78e | !hbusreq5 & v372ba66;
assign v376969b = hlock0_p & v3a676d6 | !hlock0_p & !v375d453;
assign v37721b2 = hgrant3_p & v360d1cb | !hgrant3_p & v3737ac6;
assign v3a6b94f = hbusreq6_p & v3a63805 | !hbusreq6_p & v8455b0;
assign v3a6a1e8 = hbusreq5 & v3a70d69 | !hbusreq5 & v3733d4f;
assign v37451b6 = hmaster1_p & v3a6f11c | !hmaster1_p & v375548b;
assign v3a68b7b = hmaster2_p & v373ad68 | !hmaster2_p & v375199d;
assign v374394c = hgrant4_p & v376d882 | !hgrant4_p & v3765699;
assign v3776ff3 = hbusreq7_p & v3a6f3be | !hbusreq7_p & v3757311;
assign v3a6a2d7 = hmaster0_p & v380956b | !hmaster0_p & !v8455e7;
assign v375338a = hbusreq3 & v3768931 | !hbusreq3 & v8455ab;
assign v375a4ba = hmaster0_p & v3a70925 | !hmaster0_p & v3a6b8cc;
assign v372664e = hgrant5_p & v377a4bd | !hgrant5_p & v3a683f9;
assign v374f754 = hlock6_p & v37665bf | !hlock6_p & v3a6a939;
assign v375ed5c = hmaster0_p & v3a65b4a | !hmaster0_p & v9e52e0;
assign v3740d9e = hbusreq7_p & v3a5b4d6 | !hbusreq7_p & v374d258;
assign v375a99b = hbusreq2 & v3a5b539 | !hbusreq2 & v8455ab;
assign v3778f6c = hgrant6_p & v376ea51 | !hgrant6_p & v377bf2d;
assign v3a5c6e9 = hgrant6_p & v8455ab | !hgrant6_p & !v3a6fa6f;
assign v3776ce3 = hbusreq8_p & v37312f4 | !hbusreq8_p & v3761f74;
assign v990999 = hbusreq8 & v3a5f51c | !hbusreq8 & v3a67fe2;
assign v3a70a48 = hbusreq3 & v374ccb7 | !hbusreq3 & v8455ab;
assign v3a5b4a0 = hbusreq8 & v3a6376d | !hbusreq8 & v8455ab;
assign v3a71593 = hbusreq8_p & v376ae9f | !hbusreq8_p & v37435b9;
assign v3753e00 = hlock6_p & v3a6267f | !hlock6_p & v372ab46;
assign v3756bb9 = hgrant3_p & v3a55d41 | !hgrant3_p & v3a58520;
assign v3a6567f = hmaster2_p & v3a70083 | !hmaster2_p & v373427f;
assign v374ec8b = hbusreq6 & v3a5bab6 | !hbusreq6 & v373472c;
assign v3a6f8df = busreq_p & v377d219 | !busreq_p & !v3a71519;
assign v87f2ea = jx1_p & v377e710 | !jx1_p & v372c959;
assign v375bbe2 = hbusreq7_p & v376f516 | !hbusreq7_p & v373db92;
assign v3728d75 = hbusreq8_p & v376b678 | !hbusreq8_p & v374b024;
assign v3741325 = hlock2 & v3741cd7 | !hlock2 & v3a6c2d4;
assign v37525e0 = hlock8_p & v8455ab | !hlock8_p & !v35b70fa;
assign a34d2b = hbusreq4_p & v374df64 | !hbusreq4_p & v8455bf;
assign v39a53f3 = hbusreq6_p & v2ff9190 | !hbusreq6_p & v372948c;
assign v3a6e943 = hbusreq8_p & v3a62541 | !hbusreq8_p & v3a61b9d;
assign v37247b3 = hbusreq5 & v3776756 | !hbusreq5 & v8455ab;
assign v3761f4e = hbusreq8 & v3a5d03e | !hbusreq8 & v376a06d;
assign v3779097 = hbusreq7 & v3727c74 | !hbusreq7 & v3767b5a;
assign v373a696 = hbusreq0_p & v3746fce | !hbusreq0_p & v3a707c4;
assign v3a62524 = hbusreq2_p & v3a714bd | !hbusreq2_p & v8455b7;
assign v377c2bc = hbusreq7 & v377f5ca | !hbusreq7 & v3a71146;
assign v3a704b3 = hgrant5_p & v373191d | !hgrant5_p & v374fc95;
assign v3a70d2b = hmaster1_p & v374dcbd | !hmaster1_p & v3763716;
assign v3a6c515 = hbusreq4 & v3775bd3 | !hbusreq4 & !v8455b9;
assign v3769374 = hbusreq0 & v376e040 | !hbusreq0 & v8455ab;
assign v3a6ef7d = hmaster1_p & v375d640 | !hmaster1_p & v3728d9c;
assign v37560c7 = hbusreq3 & v374a266 | !hbusreq3 & v3a70a88;
assign afdeb4 = hgrant4_p & v376a6f1 | !hgrant4_p & v372ec4e;
assign v3779d86 = hbusreq2_p & v3730b23 | !hbusreq2_p & v8455b0;
assign v39a537f = stateA1_p & v8455ab | !stateA1_p & !v39a5381;
assign v3a6910c = hbusreq2_p & v3a70641 | !hbusreq2_p & v3733383;
assign v3729430 = hbusreq6_p & v3755cb2 | !hbusreq6_p & v3a6ffe1;
assign v377a985 = hmaster2_p & v37466d4 | !hmaster2_p & v3a71314;
assign a0a219 = hmaster1_p & v3a63f9a | !hmaster1_p & v8455ab;
assign v372ab8d = hbusreq4_p & v3732359 | !hbusreq4_p & v373a331;
assign v37266cb = hgrant6_p & v3a5408c | !hgrant6_p & v3742b24;
assign v3726654 = hlock8 & v375521a | !hlock8 & v3744824;
assign v2ff8cfd = hgrant4_p & v377b6ce | !hgrant4_p & v3a5f3e3;
assign v375ce35 = hgrant6_p & v8455ab | !hgrant6_p & v37244a0;
assign v3a6f670 = hmaster1_p & v377234d | !hmaster1_p & v3a70ff4;
assign v3a702ce = hmaster2_p & v374a6a5 | !hmaster2_p & v3a66c20;
assign v3a6c1f1 = hbusreq5 & v3a5be41 | !hbusreq5 & v3a2976c;
assign v3a6f144 = hbusreq8 & v376587d | !hbusreq8 & v38074aa;
assign v3a56122 = hgrant4_p & v8455ab | !hgrant4_p & v374f9ce;
assign v3754e5a = hbusreq3_p & v3a5c945 | !hbusreq3_p & !v3a619c0;
assign v3752e46 = hbusreq2 & v375d51e | !hbusreq2 & v375b93d;
assign v375413c = hbusreq4_p & v3a70272 | !hbusreq4_p & !v3a5b68a;
assign v376cdc4 = hmaster1_p & v3735324 | !hmaster1_p & v372d75d;
assign v3a71608 = hmaster0_p & v3a66aa4 | !hmaster0_p & v3739514;
assign v374f35a = hbusreq1_p & v3a635ea | !hbusreq1_p & !v3a6d9c6;
assign v3740bf5 = hmaster0_p & v3747b81 | !hmaster0_p & v376d1cb;
assign v372f11d = hbusreq5_p & v3a68787 | !hbusreq5_p & v3766ff3;
assign v3a70e98 = hbusreq4_p & v3a5fefa | !hbusreq4_p & v3a641d5;
assign v3759a08 = hbusreq5_p & v3a70fed | !hbusreq5_p & v3742a57;
assign v3a5794d = hgrant6_p & v3a5c90c | !hgrant6_p & v3a70e6f;
assign v3a5e684 = hmaster1_p & v3755082 | !hmaster1_p & v377695e;
assign v3a70b57 = hmaster1_p & v377d1dc | !hmaster1_p & v3a6fc91;
assign v3761c4e = hbusreq3 & v373a27c | !hbusreq3 & v8455ab;
assign v374875f = hbusreq5_p & v373e845 | !hbusreq5_p & v3a6f448;
assign v3762f14 = hmaster3_p & v8455ab | !hmaster3_p & v374b88a;
assign v373653b = hmaster1_p & v373ab7e | !hmaster1_p & v373bbb4;
assign v376a7b2 = hbusreq4_p & v3737dad | !hbusreq4_p & v3772541;
assign v3a703bf = hbusreq4_p & v37692c1 | !hbusreq4_p & v373b7c5;
assign v3a5c3d6 = hbusreq5_p & v376f56d | !hbusreq5_p & baec07;
assign v3a70e65 = hlock2_p & v3731aeb | !hlock2_p & v377613d;
assign v375a918 = hbusreq4 & v3a704e5 | !hbusreq4 & v8455ab;
assign v37728a4 = stateG10_1_p & v3743690 | !stateG10_1_p & v3a6fc53;
assign v376f7d1 = hgrant5_p & v3761ff9 | !hgrant5_p & v3a6d84a;
assign v3765a1d = hmaster0_p & v377e089 | !hmaster0_p & v3774ccf;
assign v377d8b3 = hbusreq4 & v3a71416 | !hbusreq4 & !v8455b9;
assign v37798aa = hbusreq2_p & v3765901 | !hbusreq2_p & v37705d1;
assign v375ddaf = hgrant5_p & v377dc72 | !hgrant5_p & v37540e2;
assign v3a67c30 = hlock5 & v3a656be | !hlock5 & v3767797;
assign b7dcc5 = hlock5_p & v375cab5 | !hlock5_p & v3727fa7;
assign v1e37d3f = hgrant1_p & v376ef42 | !hgrant1_p & v3a70c07;
assign v37667f9 = hbusreq3_p & v1e3780f | !hbusreq3_p & v377dfe2;
assign v3a71090 = hmaster1_p & v23fd9e1 | !hmaster1_p & v3a6dcf3;
assign v373b90b = hlock8_p & v3a71386 | !hlock8_p & !v3a70b4f;
assign v374de47 = hbusreq8_p & v374ab76 | !hbusreq8_p & !v8455ab;
assign v3a6f423 = hmaster0_p & v3a5ffdd | !hmaster0_p & v372840a;
assign v3727486 = hgrant6_p & v2ff9314 | !hgrant6_p & v3a6fc54;
assign v3a60c59 = hgrant8_p & v377f7dd | !hgrant8_p & v373b6e4;
assign v3758d6c = hmaster2_p & v3a68e71 | !hmaster2_p & v37740d0;
assign v3747b2b = hmaster2_p & v373aed4 | !hmaster2_p & v8455ab;
assign v374e19c = hgrant6_p & v3a53fa4 | !hgrant6_p & v3a6f72a;
assign v3767938 = hmaster1_p & v374743d | !hmaster1_p & v3733228;
assign v23fe376 = hbusreq3_p & v3727ce4 | !hbusreq3_p & v3727d1e;
assign v3a6442f = hgrant0_p & v3a6f110 | !hgrant0_p & !v3a6f562;
assign v3808e0d = hlock0_p & v3775b81 | !hlock0_p & v8455ab;
assign v376a898 = hgrant3_p & v8455ab | !hgrant3_p & v3729d1b;
assign v3a70362 = hgrant6_p & v8455ab | !hgrant6_p & bee241;
assign v3a6ac9e = hbusreq8 & v3a6faf0 | !hbusreq8 & v3730f6f;
assign v3a665ca = hmaster1_p & v37269b2 | !hmaster1_p & !v3a69fcf;
assign v374dfe3 = hgrant5_p & v3733e56 | !hgrant5_p & v375a8d5;
assign v3a67a48 = hmaster0_p & v3733a17 | !hmaster0_p & v3726983;
assign v3757569 = hmaster2_p & v8455e7 | !hmaster2_p & v377395f;
assign v3735113 = hlock8 & v3727a12 | !hlock8 & v375c10c;
assign v37706ef = hbusreq5 & v373a2b4 | !hbusreq5 & v8455ab;
assign v375870e = hmaster0_p & v374cb62 | !hmaster0_p & v37270b9;
assign v3a7125c = hmaster0_p & v3a5f030 | !hmaster0_p & !v3736dc2;
assign v37786a4 = hgrant2_p & v374bf8a | !hgrant2_p & v23fd886;
assign v37555cd = hbusreq3_p & v3773871 | !hbusreq3_p & v3a5b9ea;
assign v3747133 = hbusreq8_p & v3750d6d | !hbusreq8_p & v3768e15;
assign v3733b37 = hbusreq3_p & v3740171 | !hbusreq3_p & v37457fb;
assign v3a70017 = hmaster1_p & v3765af5 | !hmaster1_p & !v8455ab;
assign v3761cd3 = hbusreq2 & v3a66aa4 | !hbusreq2 & v35b774b;
assign v377260b = hmaster3_p & v3a58d2e | !hmaster3_p & v8455ab;
assign v3a6d10a = hgrant2_p & v8455ab | !hgrant2_p & cd3c6e;
assign v373b380 = hmaster0_p & v3766d29 | !hmaster0_p & v3733d02;
assign v375671a = hmaster0_p & v3779680 | !hmaster0_p & v3a70f45;
assign v3a6f9f9 = hgrant4_p & v8455ab | !hgrant4_p & v373ec8e;
assign v374eb9e = hmaster2_p & v3a6fcb0 | !hmaster2_p & v372ab8d;
assign v3a53cfe = hbusreq6 & v380974c | !hbusreq6 & v8455b3;
assign v376cb9d = hmaster3_p & v3a69203 | !hmaster3_p & v3a5e755;
assign v3751849 = hlock8_p & v37737d2 | !hlock8_p & !v3a582bc;
assign v3a65130 = hbusreq7_p & v377b267 | !hbusreq7_p & v372acd3;
assign v23fe0c9 = hmaster2_p & v372ee98 | !hmaster2_p & v3a6fcc3;
assign v3750c59 = hgrant6_p & v374f511 | !hgrant6_p & v3739f84;
assign v3a6fd72 = hgrant4_p & v8455ab | !hgrant4_p & v37684a8;
assign v374c937 = hbusreq3_p & v95d97e | !hbusreq3_p & v373a391;
assign v375fdf5 = hbusreq0 & v3a70512 | !hbusreq0 & v20930c2;
assign v3a2a422 = hmaster2_p & v374db8d | !hmaster2_p & v377d7dc;
assign v377f15c = hbusreq6_p & v3a6fc11 | !hbusreq6_p & v372a4c3;
assign v3a71267 = hbusreq6_p & v3747302 | !hbusreq6_p & v377bfc0;
assign v3744151 = hmaster0_p & v2aca977 | !hmaster0_p & v3a70afe;
assign v3750d19 = hmaster0_p & v325c93e | !hmaster0_p & !v377211f;
assign v3773c10 = hbusreq7 & v372cbdf | !hbusreq7 & !v360d177;
assign v3a5c562 = hgrant4_p & v37416c6 | !hgrant4_p & v374eaeb;
assign v3a71478 = hgrant5_p & v3a60cf8 | !hgrant5_p & v374270c;
assign v3763562 = hbusreq7_p & v3a560d9 | !hbusreq7_p & v3757194;
assign v3a6fab3 = hgrant5_p & v3a58589 | !hgrant5_p & v3a710b3;
assign v3a5dfe8 = hgrant4_p & v8455ab | !hgrant4_p & !v3747c10;
assign cbd026 = hbusreq4 & v3a5f984 | !hbusreq4 & v3727084;
assign v37287d8 = hbusreq4_p & v3a67f31 | !hbusreq4_p & v8455ab;
assign v37401f0 = hbusreq1_p & v3762815 | !hbusreq1_p & v8455b0;
assign b12fe4 = hgrant6_p & v8455ab | !hgrant6_p & v374b8e2;
assign v3a62184 = hbusreq6_p & v377097a | !hbusreq6_p & v3a62a6d;
assign v3778c64 = hmaster0_p & v3a708c3 | !hmaster0_p & v3a66ade;
assign v3a5a806 = hmaster0_p & v3a6ffb6 | !hmaster0_p & v3749ec1;
assign v3726054 = hbusreq4 & v3a70f3d | !hbusreq4 & v3731230;
assign v3a5f51c = hmaster1_p & v3a5b8b9 | !hmaster1_p & v3a56e53;
assign v37565a6 = hmaster0_p & v372673d | !hmaster0_p & v376739f;
assign v3a5b5c4 = hbusreq6 & v377a36e | !hbusreq6 & v8455ab;
assign v3a70059 = hbusreq4_p & v3778cf7 | !hbusreq4_p & !v8455ab;
assign v3757a88 = hbusreq0 & v3724204 | !hbusreq0 & v8455ab;
assign v3a67ecb = hbusreq0 & v372fecf | !hbusreq0 & v3776516;
assign v3777955 = hgrant6_p & v8455ab | !hgrant6_p & !v373d53f;
assign v3760453 = hgrant4_p & v8455ab | !hgrant4_p & v374ff5a;
assign v37572af = hmaster0_p & v3a6628b | !hmaster0_p & v3a7090f;
assign v38064e4 = hbusreq6_p & v375b68b | !hbusreq6_p & v3a55482;
assign v3764d40 = hbusreq5_p & v376e7e4 | !hbusreq5_p & !v8455ab;
assign v3a64f4f = hbusreq2 & b0c091 | !hbusreq2 & !v3768ac7;
assign v3a6aa15 = hbusreq8 & v374680c | !hbusreq8 & v8455bf;
assign v374fe63 = hbusreq5 & v3740352 | !hbusreq5 & v8455ab;
assign v3a576d0 = hlock4_p & v3753f1a | !hlock4_p & v8455ab;
assign v377c9cb = hmaster2_p & v376926f | !hmaster2_p & v3739b4c;
assign v37254c0 = hbusreq3 & v3806507 | !hbusreq3 & v3a635ea;
assign v3808cf7 = hmaster0_p & v373485b | !hmaster0_p & v37665e1;
assign b33e26 = hgrant1_p & v3a5e24e | !hgrant1_p & v3733b65;
assign v372587b = hmaster0_p & v3762759 | !hmaster0_p & v3762ffa;
assign v3a5f3e3 = hgrant6_p & v377b6ce | !hgrant6_p & v3a6c835;
assign v372b8da = hbusreq5 & v3a6fa17 | !hbusreq5 & v8455ab;
assign v372e684 = hmaster1_p & v3a609da | !hmaster1_p & v374e855;
assign v3a5f50e = hbusreq2_p & v3738dca | !hbusreq2_p & !v8455ab;
assign v3736319 = hgrant3_p & v375ea58 | !hgrant3_p & !v8455ab;
assign v373e32c = hmaster2_p & v3a6dc08 | !hmaster2_p & v3a704e5;
assign v8455dd = hmaster2_p & v8455ab | !hmaster2_p & !v8455ab;
assign v3a70b92 = hbusreq3_p & v37496fa | !hbusreq3_p & v3743b9e;
assign v3725b69 = hmaster2_p & v3a70b17 | !hmaster2_p & v8455ab;
assign v3744cb5 = hbusreq0 & v374bcac | !hbusreq0 & v3733b0c;
assign v3a6f916 = hmaster1_p & v3729792 | !hmaster1_p & !v3a70e0e;
assign v376b744 = hbusreq7_p & v3735055 | !hbusreq7_p & v3748126;
assign v3736260 = hbusreq5 & v3a63556 | !hbusreq5 & v8455ab;
assign v376c25c = hmaster2_p & v3a60a68 | !hmaster2_p & v3a6f3c6;
assign v3743338 = hgrant2_p & v374ca41 | !hgrant2_p & v3a665ab;
assign v357731b = hbusreq0 & v37318e2 | !hbusreq0 & v374b6ac;
assign v375fcfb = hlock3_p & v3740349 | !hlock3_p & v8455e7;
assign v3757bac = hbusreq5_p & v3769740 | !hbusreq5_p & v3a57046;
assign v3a5fbd6 = hgrant4_p & v3a68c72 | !hgrant4_p & v372449f;
assign v373bce7 = stateA1_p & v35772a5 | !stateA1_p & !v8455ab;
assign v3a7069a = hbusreq5 & v3a6fc75 | !hbusreq5 & v3a7142a;
assign v3769ca2 = hmaster0_p & v3a6c1d3 | !hmaster0_p & !v3a6e4cd;
assign v372c9eb = hbusreq5_p & v3a5fb9e | !hbusreq5_p & v3738f35;
assign v3a63eff = hlock6 & v37559ea | !hlock6 & v3a6f914;
assign v37606c7 = stateG10_1_p & v39a537f | !stateG10_1_p & !v3766452;
assign v3a6fc8f = hlock4_p & v3735e39 | !hlock4_p & v376d856;
assign v372dfbe = hbusreq0_p & v3a6ff8a | !hbusreq0_p & v3a635ea;
assign v3a701a9 = hgrant2_p & v3774b89 | !hgrant2_p & !v373ae22;
assign v3759ec7 = hbusreq8_p & v2092abd | !hbusreq8_p & v374f094;
assign v845601 = stateG3_0_p & v8455ab | !stateG3_0_p & !v8455ab;
assign v3a6f9d9 = hbusreq4_p & v3725d7b | !hbusreq4_p & v2925d2c;
assign v3776415 = hbusreq2_p & v3746888 | !hbusreq2_p & v37240e8;
assign v37772d5 = hbusreq4 & v8455b0 | !hbusreq4 & v37406d2;
assign v3a6f47f = hmaster0_p & v3755002 | !hmaster0_p & v3a6bbe5;
assign v37261b3 = hbusreq3_p & v8455e7 | !hbusreq3_p & v8455ab;
assign v3a6e69d = hmaster1_p & v373eadd | !hmaster1_p & v8455ab;
assign v3a6ffe9 = hbusreq7 & v3730b1c | !hbusreq7 & v3a67b58;
assign v3a6fc0b = hgrant2_p & v3a635ea | !hgrant2_p & v3731304;
assign v3a70428 = hmaster1_p & v3a619c0 | !hmaster1_p & v3737bfb;
assign v372d95c = hgrant6_p & v3730bf9 | !hgrant6_p & v3a707a0;
assign v377ba8e = hmaster0_p & v373c897 | !hmaster0_p & v373b30b;
assign v372f3f7 = hgrant3_p & v3a5fcbc | !hgrant3_p & v377b4fb;
assign v3a6f09b = hmaster2_p & v2925c39 | !hmaster2_p & v3a62396;
assign v3739d45 = hbusreq6_p & v3a6cb19 | !hbusreq6_p & v8455b0;
assign v373e113 = hgrant2_p & v8455ab | !hgrant2_p & v3a6968b;
assign v3a5641a = hlock6_p & v23fe0be | !hlock6_p & !v3a70e4f;
assign v3755a83 = hgrant4_p & v8455ab | !hgrant4_p & v37525c7;
assign v376151e = hmaster2_p & v3734827 | !hmaster2_p & v377a657;
assign c17897 = hbusreq3 & v39a4ca8 | !hbusreq3 & v8455b5;
assign v376ad04 = hbusreq7 & v3774b66 | !hbusreq7 & v3774eed;
assign v37283f8 = hbusreq4_p & v3729b2e | !hbusreq4_p & !v3749bba;
assign v3726c99 = hmaster3_p & v37718d5 | !hmaster3_p & v376241e;
assign v377182c = hbusreq2_p & v1e37932 | !hbusreq2_p & v3a5d5d3;
assign v3a6672b = hbusreq3_p & v8455b0 | !hbusreq3_p & v3753dab;
assign v3a714c5 = hbusreq5 & v373fe48 | !hbusreq5 & v3729435;
assign v3748422 = stateA1_p & v3773a3d | !stateA1_p & v3a6efc4;
assign v3a5ed31 = hmaster2_p & v376f56d | !hmaster2_p & !v8455ab;
assign v377ac6f = busreq_p & v376f5fb | !busreq_p & v8455ab;
assign v372baa1 = hmaster2_p & v3727976 | !hmaster2_p & !v8455ab;
assign v3774a12 = hbusreq4_p & v3761cdb | !hbusreq4_p & v37686f3;
assign v3a6e9b1 = hlock1_p & v3a711b7 | !hlock1_p & v37547c9;
assign v3a66d94 = hgrant4_p & v3a631b4 | !hgrant4_p & v373fad7;
assign v3a6f447 = hgrant6_p & v377f7e1 | !hgrant6_p & v373ffa0;
assign v3727f69 = hbusreq7_p & v3a6f9e9 | !hbusreq7_p & v3a7044e;
assign b72b90 = hgrant2_p & v3a5eadd | !hgrant2_p & v376799e;
assign v376c335 = hmaster0_p & v37728dc | !hmaster0_p & v372e05a;
assign v3a700a6 = hmaster0_p & v3577306 | !hmaster0_p & v377d206;
assign v3a6233b = hbusreq4 & v376a14f | !hbusreq4 & v8455ab;
assign v3a70686 = hmaster1_p & v373d79e | !hmaster1_p & v372bef3;
assign v23fdd06 = hgrant4_p & v3733d6e | !hgrant4_p & v3758700;
assign v3a6462c = hmaster0_p & v37330b1 | !hmaster0_p & v3a6fc2d;
assign v3764c7c = hmaster0_p & v3a635ea | !hmaster0_p & v3a60ab2;
assign v375afc7 = hlock4 & v3a6210a | !hlock4 & v37697ba;
assign v3750b0d = hgrant6_p & v8455ab | !hgrant6_p & v3757651;
assign v375bab8 = hmaster0_p & v376654b | !hmaster0_p & v8455ab;
assign v3770b6e = hbusreq3_p & v8455bf | !hbusreq3_p & v8455b3;
assign v3a69c57 = hgrant6_p & v3725717 | !hgrant6_p & v3a629a6;
assign v375c1df = hbusreq0 & v3a6c6d6 | !hbusreq0 & v8455ab;
assign v3a5b9ea = hgrant0_p & v8455b3 | !hgrant0_p & v3a6c6aa;
assign v37586d1 = hlock7 & v3a62b35 | !hlock7 & v373402f;
assign v3a70b74 = hbusreq6_p & v377eb2d | !hbusreq6_p & v8455b0;
assign v3a6efea = hbusreq2_p & v374f35a | !hbusreq2_p & v3a68d2e;
assign v3a59409 = hbusreq3_p & v3751734 | !hbusreq3_p & v3726845;
assign v37523b5 = hbusreq7_p & v377c3f5 | !hbusreq7_p & !v8455ab;
assign v3756bd1 = hmaster3_p & v3a6ebd4 | !hmaster3_p & v1e37938;
assign v373bd77 = hlock2 & v3806a6f | !hlock2 & v3747e8e;
assign v37314f2 = hlock2_p & v373c631 | !hlock2_p & v8455e7;
assign v3a5e827 = hmaster2_p & v3a635ea | !hmaster2_p & v3a5d079;
assign v3a6a208 = hbusreq7 & v3737d23 | !hbusreq7 & v3723e62;
assign v376d79d = hbusreq2 & v3a705ac | !hbusreq2 & v8455ab;
assign v374d3b0 = hbusreq7 & v3735da7 | !hbusreq7 & !v38069e7;
assign v3769d48 = hgrant4_p & v3775dbc | !hgrant4_p & v3a70fe8;
assign v3722eee = hmaster0_p & v372455c | !hmaster0_p & v374249a;
assign v3756beb = hbusreq5 & v375588a | !hbusreq5 & v3764a8a;
assign v375068c = hlock3_p & v3750d37 | !hlock3_p & !v8455ab;
assign v3a6fec9 = hbusreq4_p & v373e0d3 | !hbusreq4_p & v8455ab;
assign v3728fda = hmaster2_p & v377a99d | !hmaster2_p & v37c02a9;
assign v3a6770f = hbusreq6 & v3a58b4c | !hbusreq6 & v373db8f;
assign v3778cf7 = hbusreq4 & v376b4e1 | !hbusreq4 & !v8455ab;
assign v3a607af = hlock0_p & v8455ab | !hlock0_p & v3765436;
assign v377eaf2 = locked_p & v3726dfa | !locked_p & v8455ab;
assign v3a70674 = hbusreq4_p & v3765758 | !hbusreq4_p & v375895e;
assign v372c1fc = hmaster2_p & v3a7137a | !hmaster2_p & v372f100;
assign v3a7104f = hbusreq7_p & v377e67a | !hbusreq7_p & v372a4ae;
assign v374248e = hmaster1_p & v3a70296 | !hmaster1_p & v3a65388;
assign v3a6f4b5 = hmaster1_p & v37281a4 | !hmaster1_p & v3a6ffdc;
assign v37662ac = hmaster0_p & v3728d9c | !hmaster0_p & v3723485;
assign v3a7001d = hgrant6_p & v3a6ee78 | !hgrant6_p & v8455ab;
assign v37759b6 = hbusreq6_p & v8455b7 | !hbusreq6_p & v3756b48;
assign v376cf96 = hbusreq5_p & v375199a | !hbusreq5_p & v3a7105f;
assign v3a70722 = hgrant6_p & v8455ca | !hgrant6_p & v3737d48;
assign v37682bc = hbusreq8 & v3769bb0 | !hbusreq8 & v3768734;
assign v3a70969 = hbusreq4_p & v3a6ef3f | !hbusreq4_p & v372a61c;
assign v377cb41 = hbusreq5_p & v3a62ccf | !hbusreq5_p & !v3a70a3a;
assign v3744daa = hmaster1_p & v3a63039 | !hmaster1_p & v3769ec3;
assign v3742bc1 = hmaster2_p & v3a5fa22 | !hmaster2_p & v375a6d3;
assign v372ad6d = hbusreq4_p & v3747042 | !hbusreq4_p & v3a5a01b;
assign v377bb3a = hlock3_p & v3755002 | !hlock3_p & !v8455ab;
assign v3a69ae7 = hbusreq6_p & v3731749 | !hbusreq6_p & !v3733862;
assign v3a70aeb = hbusreq4_p & v3a6762b | !hbusreq4_p & v372ebbf;
assign v3a61445 = hlock6_p & v3a56eb1 | !hlock6_p & !v3768202;
assign v37597a4 = hbusreq6 & v3a65da7 | !hbusreq6 & v8455bb;
assign v374774a = hmaster0_p & v37765cf | !hmaster0_p & v37390c9;
assign v3a6fcb5 = hmaster1_p & v374c190 | !hmaster1_p & v372e1bb;
assign v373c005 = hmaster0_p & v3762158 | !hmaster0_p & v3731164;
assign v37554c0 = hgrant2_p & v3743425 | !hgrant2_p & v3739f22;
assign v377205d = hlock0 & v3a635ea | !hlock0 & v3767f06;
assign v3764dc2 = hbusreq3 & v3763175 | !hbusreq3 & v8455ab;
assign v23fe209 = hbusreq7 & v375fae9 | !hbusreq7 & v3737808;
assign v3a5ca7b = stateA1_p & v8455ab | !stateA1_p & !v3742b0e;
assign v3772f4d = hbusreq2 & v3749b46 | !hbusreq2 & v376441d;
assign v3a5b4c1 = hgrant2_p & v3758472 | !hgrant2_p & v376efda;
assign v377803a = hbusreq6 & v376b83d | !hbusreq6 & v373c965;
assign v375d12e = hbusreq2_p & v3778425 | !hbusreq2_p & v37500ac;
assign v3751e07 = hmaster0_p & v38087c5 | !hmaster0_p & v372a1b6;
assign v3a70193 = hbusreq6_p & v3a593cb | !hbusreq6_p & v377e05a;
assign v3a5a75c = hgrant5_p & v374e3fa | !hgrant5_p & v37627a8;
assign v3a6c7c6 = hgrant3_p & v3754877 | !hgrant3_p & v3a69043;
assign v377702c = hgrant2_p & v3a6ffb6 | !hgrant2_p & v374d2dd;
assign v3a64abe = hmaster0_p & v3745589 | !hmaster0_p & v372efcd;
assign v3807f45 = hbusreq3_p & v37618e0 | !hbusreq3_p & v8455b0;
assign v38099c1 = hlock0_p & v373be25 | !hlock0_p & v3a5cfd9;
assign v37515a6 = hbusreq4_p & v2ff9291 | !hbusreq4_p & v372874c;
assign v376f0ab = hmaster2_p & v3a69444 | !hmaster2_p & v3778afd;
assign v373389a = hbusreq3_p & v374d184 | !hbusreq3_p & v8455ab;
assign v375d4d4 = hbusreq4_p & v374f543 | !hbusreq4_p & v8455ab;
assign v3730a61 = hmaster2_p & v3a6a8c0 | !hmaster2_p & be54b2;
assign v3752b6a = hbusreq6_p & v3a6e9b8 | !hbusreq6_p & v3749a1d;
assign v374cf79 = hbusreq6 & v3a6006a | !hbusreq6 & v3a70fd2;
assign v3742b84 = hlock6 & v3a6fa7e | !hlock6 & v3740839;
assign v373becf = hmaster1_p & v3747929 | !hmaster1_p & v3a65260;
assign v3741286 = hbusreq8_p & v37715b9 | !hbusreq8_p & ce7a16;
assign v3770f54 = hlock0 & v3a71267 | !hlock0 & v3a70765;
assign v3a5bed2 = hmaster1_p & v375c0e8 | !hmaster1_p & v3a6f6fe;
assign v3a6f5eb = hmaster0_p & v3750218 | !hmaster0_p & v3a70d93;
assign v376cd14 = hbusreq6_p & v3763a84 | !hbusreq6_p & v8455ab;
assign v3808e5b = hbusreq5 & v376086c | !hbusreq5 & v8455ab;
assign v3741edb = hbusreq8_p & v988a3b | !hbusreq8_p & v3772773;
assign v3a6efd2 = hlock6 & v374b20c | !hlock6 & v377228d;
assign v37274a2 = hgrant7_p & v8455ab | !hgrant7_p & v3749412;
assign v374053e = hbusreq1_p & v3730de9 | !hbusreq1_p & v374f033;
assign v37684ed = hlock1_p & v3a70e06 | !hlock1_p & !v374f593;
assign v3a6eebb = hmaster2_p & v3a67458 | !hmaster2_p & v3a6e548;
assign v39a4dbb = hbusreq2_p & v37502b7 | !hbusreq2_p & v3735e39;
assign v3728df3 = stateG10_1_p & v3809adf | !stateG10_1_p & !v37234e7;
assign v3a6a3e6 = hbusreq0 & v3a58429 | !hbusreq0 & v8455ab;
assign v3739e55 = hmastlock_p & v3759020 | !hmastlock_p & v8455ab;
assign v3807686 = hgrant4_p & v1e37b99 | !hgrant4_p & !v372d744;
assign v3767419 = hmaster2_p & v8455e7 | !hmaster2_p & v372eaaf;
assign v377b6b2 = hmaster2_p & v375a95b | !hmaster2_p & v3735272;
assign v3a70b5f = hbusreq0_p & v3a635ea | !hbusreq0_p & v3809093;
assign v3754fd2 = hbusreq6_p & v3a6ae2d | !hbusreq6_p & !v8455ca;
assign v3a6cc72 = hbusreq6 & v3a63abb | !hbusreq6 & v8455ab;
assign v372685c = hlock5 & v3a6f81c | !hlock5 & v376f51c;
assign v3a6d18a = hlock0_p & v3725410 | !hlock0_p & v3770187;
assign v3a70557 = hgrant4_p & v3a5a510 | !hgrant4_p & v374c052;
assign v3736db8 = hgrant6_p & v3a57fff | !hgrant6_p & v377c003;
assign v37576d1 = hgrant2_p & dbdbc5 | !hgrant2_p & v372eecf;
assign v374aece = hbusreq0 & v3a710eb | !hbusreq0 & v3757407;
assign v373703c = hmaster2_p & v37453d7 | !hmaster2_p & v3a62a6d;
assign v377b779 = hgrant2_p & v374d542 | !hgrant2_p & v3a6e516;
assign v374bc02 = hmaster2_p & v37482f8 | !hmaster2_p & v377df2e;
assign v3a57f18 = hbusreq8_p & v37260af | !hbusreq8_p & v375d17d;
assign v37518c9 = hmaster1_p & v3a6f4ee | !hmaster1_p & v374f1e9;
assign v372ef9b = hburst0 & v372b0cd | !hburst0 & b09623;
assign v3744265 = hbusreq1_p & v3a64566 | !hbusreq1_p & !v3a53cc3;
assign v3737a30 = hgrant3_p & v8455be | !hgrant3_p & !v373d434;
assign v3a70629 = hgrant6_p & v3a71411 | !hgrant6_p & v3728f87;
assign v3738bdf = hmaster1_p & v3a5fae2 | !hmaster1_p & v374610d;
assign v37539c8 = hbusreq7_p & v37734cb | !hbusreq7_p & v8455c7;
assign v3724926 = hmaster0_p & v8455b3 | !hmaster0_p & v37364af;
assign v3a64eb3 = hbusreq7_p & v377baf9 | !hbusreq7_p & !v3a6d7a0;
assign v3a634fd = hmaster0_p & v372d939 | !hmaster0_p & v37270b9;
assign v372e083 = hmaster2_p & v8455b0 | !hmaster2_p & v3a6fa39;
assign v3a629a6 = hgrant2_p & v3765e79 | !hgrant2_p & v3a5e6f6;
assign v377fc89 = hmaster1_p & v8455ab | !hmaster1_p & v372e4e1;
assign v3a71101 = hgrant5_p & v37378d4 | !hgrant5_p & v375783b;
assign v37326a5 = hbusreq6 & v375d05d | !hbusreq6 & v3748797;
assign v3747b55 = hmaster1_p & v3a6e5f0 | !hmaster1_p & v376c25b;
assign v376891a = hlock5 & v3738750 | !hlock5 & v3739ec6;
assign v3a57b60 = hbusreq6_p & v3759044 | !hbusreq6_p & v372c37f;
assign v3a6f767 = hbusreq6_p & v3737c86 | !hbusreq6_p & v376a4dd;
assign v377ddae = hlock3_p & v3767d4e | !hlock3_p & !v8455ab;
assign v37611fb = hbusreq5_p & v3a6fc67 | !hbusreq5_p & v37258b4;
assign v377ea1b = hbusreq8 & v3a6f437 | !hbusreq8 & v3809142;
assign a8fc27 = hgrant2_p & v3a70403 | !hgrant2_p & v3a689eb;
assign v37638fe = hmaster0_p & v3a6f359 | !hmaster0_p & v377904f;
assign v374fdc9 = hmaster0_p & v3a5e24e | !hmaster0_p & v372542e;
assign v3744d2b = hmaster0_p & v3a6fa9a | !hmaster0_p & v3a583b0;
assign v3776852 = hlock0 & v38072fd | !hlock0 & v377ecd4;
assign v3a61480 = hmaster2_p & v37270d9 | !hmaster2_p & v3767f33;
assign v373fa07 = hlock3_p & v3759f8b | !hlock3_p & v8455b0;
assign v3a70efe = hmaster0_p & v37c36cb | !hmaster0_p & !v8455b3;
assign v38070c7 = hmaster0_p & v373a4e4 | !hmaster0_p & v37452a4;
assign v3a63004 = hmaster0_p & v376a14f | !hmaster0_p & v373b16e;
assign v3a6f3c2 = hbusreq8 & v3a61820 | !hbusreq8 & v376ae9f;
assign v3a6396b = hmaster0_p & v37737aa | !hmaster0_p & v3a70d3f;
assign v3771715 = hgrant4_p & v8455c1 | !hgrant4_p & v3729b4c;
assign v373ee81 = hmaster0_p & v3a701a1 | !hmaster0_p & v8cf677;
assign v37584fe = hgrant0_p & v3a65596 | !hgrant0_p & v8455ab;
assign v3a6f659 = hbusreq6 & v884deb | !hbusreq6 & v3a635ea;
assign v3777c4e = hmaster1_p & v3a29814 | !hmaster1_p & v3a5afd7;
assign v374a9cd = hbusreq8_p & v3a62c37 | !hbusreq8_p & v89df94;
assign v3760740 = hlock0_p & v3a5f8d0 | !hlock0_p & v3a6c725;
assign v3a7078a = hbusreq3_p & v3a68bf8 | !hbusreq3_p & v377c31a;
assign v3745e0d = hbusreq7_p & v3a6ef38 | !hbusreq7_p & v376dad0;
assign v373e031 = hlock6 & v376d8c1 | !hlock6 & v3a57f8b;
assign v3a6a81f = hbusreq8_p & v372ae4f | !hbusreq8_p & v374c6aa;
assign v3a5a24d = hmaster0_p & v3730ffe | !hmaster0_p & v8455ab;
assign v3729c45 = hbusreq4_p & v3747302 | !hbusreq4_p & v3757cd6;
assign v377e087 = hlock2 & v3728346 | !hlock2 & v3a66538;
assign v3a708af = hgrant0_p & v8455ab | !hgrant0_p & v3776c09;
assign v3779e95 = hgrant4_p & v8455c1 | !hgrant4_p & v3a6f45a;
assign v3777312 = hmaster1_p & v8455b3 | !hmaster1_p & v3a7054c;
assign v373fe48 = hmaster0_p & v375afe9 | !hmaster0_p & v3745d9c;
assign v3753bfb = hmaster0_p & v376801c | !hmaster0_p & v372b7a3;
assign v372e95b = hbusreq4_p & v3a702c2 | !hbusreq4_p & v8455b0;
assign v373a494 = jx0_p & v8455ab | !jx0_p & v375dc63;
assign v3a70ca5 = hlock5_p & v37532ee | !hlock5_p & v3758466;
assign v372a20d = hmaster0_p & v3a65b4a | !hmaster0_p & v3a6402e;
assign v3a62b13 = hmaster0_p & v3769e49 | !hmaster0_p & v37585d8;
assign v3a55352 = hgrant8_p & v372f320 | !hgrant8_p & v373e8de;
assign v372f464 = hmaster1_p & v3757ad8 | !hmaster1_p & v38065f1;
assign v3a6af99 = stateG2_p & v8455ab | !stateG2_p & !v865472;
assign v3a608b9 = hlock4_p & v3a6ab5f | !hlock4_p & !v8455ab;
assign v3741ea8 = hgrant5_p & v8455ab | !hgrant5_p & v3a6e884;
assign v373b59f = hmaster2_p & v325c960 | !hmaster2_p & v3763668;
assign v2925ce0 = hmaster2_p & v3a6ebcd | !hmaster2_p & v372526a;
assign v3a6ffc5 = hbusreq8_p & v372c921 | !hbusreq8_p & v8455ab;
assign v38075aa = hbusreq6_p & v37323a5 | !hbusreq6_p & v8455ab;
assign v3a6f7c5 = hmaster2_p & v3766bc8 | !hmaster2_p & !v3732569;
assign v3764a7d = hmaster2_p & v3a6f65c | !hmaster2_p & v3a71025;
assign v3a69f17 = hlock6_p & v3a63e82 | !hlock6_p & !v35772a6;
assign v373efc2 = hbusreq3_p & v375e657 | !hbusreq3_p & !v3a69591;
assign v3771733 = hbusreq6 & v373a27c | !hbusreq6 & v8455e7;
assign v2aca784 = hbusreq1_p & v37513d1 | !hbusreq1_p & v1e3731f;
assign v37559d6 = hbusreq8_p & v375654b | !hbusreq8_p & v3773040;
assign v372d772 = hbusreq4 & v374eb89 | !hbusreq4 & v3379037;
assign v3a6f5e6 = hgrant5_p & v3755ad0 | !hgrant5_p & v3730895;
assign v3747cfc = hmaster3_p & v374f8b5 | !hmaster3_p & v3730766;
assign v3a59eb3 = hgrant6_p & v8455ab | !hgrant6_p & v373e32a;
assign v3725d5a = hbusreq7 & v3a69c64 | !hbusreq7 & v8455b3;
assign v37299ef = hbusreq8 & v23fe21d | !hbusreq8 & !v8455ab;
assign v3725380 = hlock5 & v3a7152f | !hlock5 & v376d72e;
assign v372946e = hlock0 & v374acbe | !hlock0 & v374b37d;
assign v37538af = hmaster2_p & v3a70a5c | !hmaster2_p & d5f283;
assign v3a652b6 = hmaster0_p & v372e250 | !hmaster0_p & v374e758;
assign v3a70574 = hmaster2_p & v8455ab | !hmaster2_p & v38074ac;
assign v1e37e82 = hlock4_p & v372a4c1 | !hlock4_p & v8455ab;
assign v3a6f1ad = hbusreq4_p & v3a6ac26 | !hbusreq4_p & v3a6ac2a;
assign v375bc08 = hgrant2_p & v8455ba | !hgrant2_p & v3769d3e;
assign v3746dc9 = hbusreq4_p & v37617de | !hbusreq4_p & v3a70952;
assign v3777f86 = hbusreq4_p & v3a6f29a | !hbusreq4_p & v37492bc;
assign v3a63e9d = hbusreq5 & v374a7de | !hbusreq5 & v3a2a107;
assign v377854f = hmaster0_p & v3736ded | !hmaster0_p & v3a70a2b;
assign v3a7093c = hbusreq4_p & v3768c3c | !hbusreq4_p & v3a70326;
assign v38079dc = hbusreq4 & v3a5966b | !hbusreq4 & v3a5741c;
assign v3a6ddea = hmaster2_p & v39a4c67 | !hmaster2_p & v372a85f;
assign v3743d47 = jx1_p & v37352fa | !jx1_p & v3a700e8;
assign d3482c = hmaster1_p & v377ea20 | !hmaster1_p & v3732b3c;
assign v3a6f414 = hgrant5_p & v3a6ff2e | !hgrant5_p & v3a54b2b;
assign v373a629 = hgrant4_p & v372493b | !hgrant4_p & v3752e24;
assign v37369b2 = hbusreq2_p & v3750eaa | !hbusreq2_p & v8455ab;
assign v375cd8b = hbusreq5 & v3755045 | !hbusreq5 & v3759f77;
assign v374074a = hmaster2_p & v3a67de3 | !hmaster2_p & v3767b70;
assign v3a6f533 = hmaster2_p & v8455b3 | !hmaster2_p & !v3768202;
assign v3a55e75 = hbusreq7 & v373e57b | !hbusreq7 & v8455ab;
assign v3750abf = hbusreq7_p & v372cdec | !hbusreq7_p & v3a5cf28;
assign v35b73a5 = hlock5 & v360bedd | !hlock5 & v3731d8f;
assign v37388d6 = hmaster2_p & v8455b0 | !hmaster2_p & v374ebb0;
assign v37235bd = hgrant6_p & v3a6f43e | !hgrant6_p & v37609a6;
assign v3a6c23b = hbusreq1_p & v374c6df | !hbusreq1_p & v8455ab;
assign v373c8c5 = hmaster2_p & v3a6f781 | !hmaster2_p & v37646e1;
assign v375f0ba = hgrant2_p & v377d4a0 | !hgrant2_p & v37747b4;
assign v372bf93 = hlock2_p & v3a57c48 | !hlock2_p & v35b70e6;
assign v3778b83 = hbusreq5_p & v3768172 | !hbusreq5_p & !v8455ab;
assign v372b795 = hbusreq6_p & v37485ec | !hbusreq6_p & c6598e;
assign v374067b = hmaster1_p & v8455ab | !hmaster1_p & v373894a;
assign v37708e7 = hgrant2_p & v3a646f5 | !hgrant2_p & v38099ce;
assign v3a71084 = stateA1_p & v8455ab | !stateA1_p & v3a6a939;
assign v374882c = hbusreq5 & v3a5d678 | !hbusreq5 & v3a635ea;
assign v3a6d69b = hlock0_p & v3a7153a | !hlock0_p & v3a63805;
assign v3730895 = hmaster1_p & v3a5bf5f | !hmaster1_p & v3741c4b;
assign v37422f3 = hgrant6_p & v376b088 | !hgrant6_p & v3763668;
assign v3747bfe = hmaster2_p & v377adf0 | !hmaster2_p & v3a7094d;
assign v3a611d8 = hbusreq8 & b9d061 | !hbusreq8 & v377386a;
assign v3a65dad = hmaster1_p & v3a55a58 | !hmaster1_p & !v3a6f446;
assign v3743dff = hlock8_p & v3724908 | !hlock8_p & v374ddef;
assign v372f231 = hlock6_p & v8455ab | !hlock6_p & v3779582;
assign v374e207 = hbusreq7_p & v3761953 | !hbusreq7_p & !v3736adf;
assign v3a6827b = hbusreq0 & v375a234 | !hbusreq0 & v3732515;
assign v3724947 = hmaster2_p & v3771c59 | !hmaster2_p & v377957e;
assign v373f2d2 = hmaster1_p & v8455ab | !hmaster1_p & v3a6e9b0;
assign v375ed9f = hgrant2_p & v3751931 | !hgrant2_p & v3a699f5;
assign v376f9be = hmaster0_p & v3723a2d | !hmaster0_p & v374523d;
assign v3a6ba77 = hbusreq6_p & v374faa9 | !hbusreq6_p & v37775eb;
assign v373a303 = hbusreq0 & v3a6784d | !hbusreq0 & v8455ab;
assign v377da26 = hlock6 & v3a680f4 | !hlock6 & v3a55673;
assign v3774a8f = hgrant0_p & v3749529 | !hgrant0_p & v3752e8e;
assign v3749831 = hbusreq0 & v3779734 | !hbusreq0 & v3a70ef4;
assign v3762bf1 = hlock0_p & v37775c4 | !hlock0_p & v3a6fe80;
assign v3a6f069 = hmaster1_p & v3769f7f | !hmaster1_p & v3a6fb1d;
assign v3770a3b = hlock5_p & v3735f51 | !hlock5_p & v3775931;
assign v374c154 = hbusreq8_p & v3a62f05 | !hbusreq8_p & v1e37a30;
assign v3a659eb = hmaster2_p & v376285a | !hmaster2_p & v3a6f018;
assign v3a6d84a = hmaster1_p & v3a70e4c | !hmaster1_p & v3731725;
assign v37730b9 = hmaster2_p & v1e3787a | !hmaster2_p & v3739ddf;
assign v37632c6 = hbusreq7_p & v3a713b4 | !hbusreq7_p & v3a6ec83;
assign v3a70f1d = hmaster0_p & v372bb72 | !hmaster0_p & v3766573;
assign v375641f = hbusreq3_p & v3759b2f | !hbusreq3_p & v3a6f43e;
assign v3a6fbed = hbusreq3 & v3a590de | !hbusreq3 & v375b9c1;
assign v3757dad = hbusreq3 & v8455ab | !hbusreq3 & v8455b0;
assign v37320bb = hbusreq2_p & v37400f8 | !hbusreq2_p & v3a6ffae;
assign v39ea7a8 = hlock0_p & v95d97e | !hlock0_p & !v3a6ac26;
assign v3728fd0 = hmaster2_p & v3a57584 | !hmaster2_p & !v3a5952d;
assign v3a658f7 = hmaster2_p & v3a5b7c2 | !hmaster2_p & !v3766ff7;
assign v3757637 = hbusreq6_p & v3747ec5 | !hbusreq6_p & v37311de;
assign v3a5fe1d = hgrant1_p & v3a66110 | !hgrant1_p & v375bbe9;
assign v3a6257d = hmaster1_p & v3a5637b | !hmaster1_p & v3a6f3f2;
assign v3a61202 = hbusreq5 & v37251f1 | !hbusreq5 & v8455bf;
assign b9f474 = hbusreq0_p & v3723430 | !hbusreq0_p & v8455e7;
assign v372594c = hgrant6_p & v8455c9 | !hgrant6_p & v3741e68;
assign v3751af0 = hbusreq6 & v373d78b | !hbusreq6 & v8455ab;
assign v3746d4a = hlock4 & v3a6f0a5 | !hlock4 & v3778dd7;
assign v374d778 = hmaster0_p & v3778d7f | !hmaster0_p & v376b540;
assign v37775ff = hmaster0_p & v376c6ba | !hmaster0_p & v3a57106;
assign v37601df = jx0_p & v8455ab | !jx0_p & v3a6ec10;
assign v3807afa = hbusreq4_p & v372e96f | !hbusreq4_p & v3a6f6b9;
assign v372505f = hmaster0_p & v3734374 | !hmaster0_p & v8455e7;
assign v3a7138c = hlock5 & v3a57c0d | !hlock5 & v372c85f;
assign v3768a79 = hbusreq2_p & v3a6dd65 | !hbusreq2_p & v372fb9d;
assign v377a657 = hgrant4_p & v1e37b99 | !hgrant4_p & v3a65e1e;
assign v3a6f612 = hlock6_p & v372fba5 | !hlock6_p & v3724940;
assign v3a644d3 = hgrant7_p & v8455b9 | !hgrant7_p & v3a6706d;
assign v3a71048 = hbusreq7 & v37305c2 | !hbusreq7 & v3759284;
assign v375d80d = hgrant1_p & v37547c9 | !hgrant1_p & !v8455ab;
assign v373318b = hmaster2_p & v3753dab | !hmaster2_p & v372b5f5;
assign v3a67ec4 = hlock2 & v37477dd | !hlock2 & v3744cea;
assign v3a6fb17 = hbusreq7 & v3726eb4 | !hbusreq7 & v8455ab;
assign v3a70081 = hmaster1_p & v375db64 | !hmaster1_p & v3739e31;
assign v3a577fe = hbusreq4_p & v377c700 | !hbusreq4_p & v8455ab;
assign v377d8f9 = stateG2_p & v8455ab | !stateG2_p & !v3751c12;
assign v3769a63 = jx0_p & v3809d53 | !jx0_p & v3a5c4b0;
assign v37654a9 = hbusreq7 & v3a70abb | !hbusreq7 & v372ab70;
assign v377815d = hgrant7_p & v8455ab | !hgrant7_p & v39372da;
assign v3378a0a = hgrant1_p & v3775b81 | !hgrant1_p & v8455ab;
assign v2ff8f33 = hlock5 & v37523ef | !hlock5 & v372cdb0;
assign v3757e56 = hbusreq7_p & v3a651c8 | !hbusreq7_p & v3a6e29d;
assign v375c062 = hbusreq5 & v372aa71 | !hbusreq5 & v3a70347;
assign v3a6c860 = hlock0_p & v3a706d1 | !hlock0_p & v3770187;
assign v3a707a4 = hmaster0_p & v23fdf1b | !hmaster0_p & v37420bb;
assign v377314f = hburst0 & v3a6ab5f | !hburst0 & v8455e1;
assign v3a713ea = hmaster1_p & v376d1dd | !hmaster1_p & v3747271;
assign v374bcb5 = hmaster0_p & v3a7149d | !hmaster0_p & v37767fa;
assign v3a6850e = hgrant4_p & v8455ab | !hgrant4_p & v377c31d;
assign v3746e79 = hbusreq1_p & v3a6f84d | !hbusreq1_p & v372981e;
assign v3a6fbbd = hlock5_p & v3a6ff31 | !hlock5_p & !v376c7cc;
assign v39eb565 = hmaster2_p & v3a53c18 | !hmaster2_p & v3a6fc5e;
assign v3a6f15a = jx0_p & v3a7014f | !jx0_p & v377f253;
assign v372ee9a = hbusreq3_p & v3a70fa2 | !hbusreq3_p & !v8455ab;
assign v3a704b1 = hlock3_p & v3722b42 | !hlock3_p & v37459dd;
assign v3763548 = hmaster2_p & v3a635ea | !hmaster2_p & v372d299;
assign v3a598a0 = hbusreq3_p & v3747302 | !hbusreq3_p & v3a62fa3;
assign v3a65607 = hmaster0_p & v3a6f97b | !hmaster0_p & v3a6f35b;
assign v3a6464f = hgrant6_p & v8455ca | !hgrant6_p & v3a702ec;
assign v3a71170 = hbusreq4_p & v3a6e81e | !hbusreq4_p & v3a71012;
assign v3747a68 = hlock5_p & v3770c1a | !hlock5_p & v3a6512d;
assign v3a70ecb = hgrant4_p & v3745ac6 | !hgrant4_p & v3a55b1d;
assign v374b0eb = hbusreq7_p & v373c8db | !hbusreq7_p & v8455ab;
assign v3a707f2 = hgrant4_p & v3758bbd | !hgrant4_p & v8455ab;
assign v373a072 = hlock5_p & v3a713cd | !hlock5_p & v8455ab;
assign v3779988 = hmaster2_p & v3759a7f | !hmaster2_p & v374f968;
assign v374e05d = hmaster1_p & v3a7125c | !hmaster1_p & !v3a616fb;
assign v3a713e3 = hgrant3_p & v8455be | !hgrant3_p & !v374f609;
assign v3731aaf = hmaster0_p & v3806ff5 | !hmaster0_p & v373026e;
assign v3725671 = hlock4 & v372a39d | !hlock4 & v374178a;
assign v3749a32 = hbusreq0 & v37684a8 | !hbusreq0 & v377c31d;
assign v3a70474 = hlock5 & v3769069 | !hlock5 & v376ed63;
assign v372af67 = hbusreq2 & v37566b2 | !hbusreq2 & !v8455ab;
assign v3752c73 = hbusreq4_p & v3a5618d | !hbusreq4_p & v375a5b6;
assign v3a6c81d = hmaster1_p & v372f6d3 | !hmaster1_p & v3a6fb0e;
assign v3a55081 = hbusreq5_p & v374f8f6 | !hbusreq5_p & !v3a7113b;
assign v3a5b52c = hbusreq5 & v3a2a0f4 | !hbusreq5 & v3a70484;
assign v3a6ff3e = hmaster0_p & v377989c | !hmaster0_p & v3a7089b;
assign v3766bc8 = hbusreq2_p & v3a70c07 | !hbusreq2_p & v1e38224;
assign v3750b02 = hmaster2_p & v3753d94 | !hmaster2_p & v3a6f3e7;
assign b318d6 = hgrant4_p & v375582f | !hgrant4_p & v3762245;
assign v3a6cc28 = hgrant5_p & v8455ab | !hgrant5_p & v3a70005;
assign v372f2ce = hmaster2_p & v1e3787a | !hmaster2_p & v37466cb;
assign v3378c57 = hlock4_p & v372c6cb | !hlock4_p & v373ddca;
assign v37305c2 = hmaster1_p & v3a635ea | !hmaster1_p & v3745eb8;
assign v3725ceb = hmaster0_p & v3734967 | !hmaster0_p & v377613b;
assign v8e4f94 = hbusreq4_p & v3756de3 | !hbusreq4_p & v8455cb;
assign v3a704f0 = hbusreq5 & v3771c5f | !hbusreq5 & v1e379c4;
assign v372bb25 = hgrant5_p & v3a70769 | !hgrant5_p & v3a5b687;
assign v3769cd6 = hgrant2_p & v375d38f | !hgrant2_p & !v3761fc1;
assign v3985142 = hgrant5_p & v3728876 | !hgrant5_p & v373052f;
assign v373e121 = jx0_p & v377a993 | !jx0_p & v1e37e1f;
assign v37666b4 = hready_p & v376a25e | !hready_p & v372c046;
assign v377825c = hbusreq3_p & v377c103 | !hbusreq3_p & v3778528;
assign v3756ea2 = hbusreq5 & v3a54ebe | !hbusreq5 & v9e8d30;
assign a38ed7 = hbusreq1_p & v3a5c5ae | !hbusreq1_p & !v3809adf;
assign v3a6fc38 = hmaster0_p & v3727a2f | !hmaster0_p & v377376d;
assign v3775790 = hgrant5_p & v3768c01 | !hgrant5_p & v3765f0a;
assign v37c0190 = hgrant3_p & v8455ab | !hgrant3_p & v3769041;
assign v3a70d93 = hmaster2_p & v3759119 | !hmaster2_p & !v3a5dbd1;
assign v372a1d4 = hbusreq5 & v3a63ece | !hbusreq5 & v3763db6;
assign c48c9d = hmaster0_p & v37370c6 | !hmaster0_p & v3a6fb52;
assign v374c8ec = hbusreq0 & v3a714e1 | !hbusreq0 & v3a6cb4e;
assign v3731e16 = hmaster0_p & v3a70c8c | !hmaster0_p & v374e1dc;
assign v377167d = hbusreq5_p & v3a70ebc | !hbusreq5_p & !v3748544;
assign v372667b = hlock7_p & v3a56bb5 | !hlock7_p & !v8455ab;
assign v37280de = hbusreq2_p & v3a5ba97 | !hbusreq2_p & v8455ab;
assign v372295a = stateA1_p & v8455ab | !stateA1_p & v3a58588;
assign v3a64e01 = hbusreq5_p & v3a5949f | !hbusreq5_p & v3a58c07;
assign v37709ec = hbusreq5_p & v373cd8a | !hbusreq5_p & !v3a6355c;
assign v3747e71 = hbusreq8_p & v3a5d1c9 | !hbusreq8_p & v376bc98;
assign v3749283 = hmaster1_p & v3a67862 | !hmaster1_p & v3a6b78f;
assign v374fe39 = hbusreq0 & v3a7145a | !hbusreq0 & v377ca8e;
assign v3746fd4 = hgrant6_p & v1e37cd6 | !hgrant6_p & v3742dae;
assign v3a59505 = hbusreq4_p & v3759b2f | !hbusreq4_p & !v373be25;
assign v3735d84 = hbusreq5_p & v3755731 | !hbusreq5_p & v3a57cc8;
assign v3808d56 = hmaster2_p & v3736afd | !hmaster2_p & v3a6a374;
assign v3756737 = hmaster0_p & v372cec6 | !hmaster0_p & v373026e;
assign v377bb0e = hmaster2_p & v376e717 | !hmaster2_p & v3a70096;
assign v380705b = hmaster1_p & v376f499 | !hmaster1_p & v3a65019;
assign v3a6ef4d = hlock4 & v38072fd | !hlock4 & v3763186;
assign v37293c3 = hmaster0_p & v3747bc9 | !hmaster0_p & !v8455ab;
assign v373c3ac = hmaster1_p & v3774db3 | !hmaster1_p & v376769a;
assign v37667c6 = hmaster2_p & v376dbdf | !hmaster2_p & v376f2f8;
assign v374d86e = hlock5 & v3778c7f | !hlock5 & v9204d4;
assign v377e9cd = hgrant4_p & v8455ab | !hgrant4_p & v3a6b20a;
assign v374dc53 = hlock6 & v3a71064 | !hlock6 & v39a4e43;
assign v37580d5 = hbusreq4 & v3775750 | !hbusreq4 & v35b774b;
assign v373d238 = hbusreq7_p & a0a219 | !hbusreq7_p & v37514dd;
assign v377a0da = hmaster2_p & v3746641 | !hmaster2_p & v3a71308;
assign v374e079 = hgrant4_p & v3751389 | !hgrant4_p & v372b02f;
assign v3750088 = hmaster2_p & v3731dfd | !hmaster2_p & v8455ab;
assign v3a70e91 = hbusreq8 & v3a7076a | !hbusreq8 & v37285cd;
assign v37723ce = hbusreq5 & v37329ec | !hbusreq5 & v3771994;
assign v3a6f6cd = hbusreq8 & v3741793 | !hbusreq8 & v3737808;
assign v3726072 = hbusreq8 & v3a64f96 | !hbusreq8 & v3746f9d;
assign v3738da4 = hmaster1_p & v3742b79 | !hmaster1_p & v2ff9229;
assign v3a701e9 = hgrant6_p & v37483dd | !hgrant6_p & v3762525;
assign v376eed8 = hlock5 & v3770def | !hlock5 & v3763076;
assign v375485b = hbusreq5_p & v3a63f9a | !hbusreq5_p & v3751dcc;
assign v376f665 = hburst1 & v2aca977 | !hburst1 & v372ecab;
assign v37675d5 = hlock0 & v3a6bf41 | !hlock0 & v3a66306;
assign v3a29760 = hlock8_p & v8455ab | !hlock8_p & v3a70311;
assign v374922a = hbusreq6_p & v375a4fa | !hbusreq6_p & v37510b1;
assign v372dec8 = hgrant1_p & v37496fa | !hgrant1_p & v3a635ea;
assign v37263d2 = hlock8 & bd1306 | !hlock8 & v375f28d;
assign v3a5591a = hbusreq5_p & v3736411 | !hbusreq5_p & v374c73c;
assign v37540df = hgrant6_p & v372fb1b | !hgrant6_p & !v3a66584;
assign v37263b9 = hbusreq4 & v3a5e10c | !hbusreq4 & v374d63f;
assign v3a53c18 = hgrant4_p & v8455c2 | !hgrant4_p & v3a6f9f5;
assign v37269bf = hmaster0_p & v3746c51 | !hmaster0_p & v3a70db0;
assign v3748266 = hbusreq5_p & v3a63512 | !hbusreq5_p & v3a6f335;
assign v377aa81 = hbusreq4_p & v376dc91 | !hbusreq4_p & v372a954;
assign v3a70f19 = hgrant3_p & v3a5c945 | !hgrant3_p & v376e41a;
assign v3778546 = hbusreq0 & v3758915 | !hbusreq0 & v372f1b9;
assign v3a5665e = hbusreq4_p & v3a6d625 | !hbusreq4_p & v3a667a7;
assign v372c502 = hlock2_p & v3778425 | !hlock2_p & v3748d3e;
assign v3a70a1f = hmaster1_p & v37384a6 | !hmaster1_p & v375b12b;
assign c2c2bc = hgrant6_p & v3a6fe48 | !hgrant6_p & v3771667;
assign v373261f = hlock6_p & v372adb5 | !hlock6_p & !v8455ab;
assign v3759044 = hbusreq6 & v3733b37 | !hbusreq6 & v8455e7;
assign v373b0d0 = hbusreq0 & v3739e7a | !hbusreq0 & v1e37558;
assign v3757ec8 = hbusreq2_p & v3a563ba | !hbusreq2_p & !v8455ab;
assign v33790a4 = hgrant5_p & v3a6c527 | !hgrant5_p & v37725b5;
assign v3723903 = hlock6 & v3a54f85 | !hlock6 & v3766b81;
assign v380735e = hmaster1_p & v372a465 | !hmaster1_p & v3773ab1;
assign v375706b = hmaster0_p & v3a680bd | !hmaster0_p & v375a086;
assign v3763e92 = hbusreq8_p & v3a6eeb7 | !hbusreq8_p & v3a7021a;
assign v3a70bb8 = hbusreq6 & v3a5a158 | !hbusreq6 & v3a62a6d;
assign v3a6fa4b = hready_p & v8455e7 | !hready_p & v3a58cb2;
assign v37742ca = hlock5_p & v8455ab | !hlock5_p & !v3a641c0;
assign v3a6f0b2 = hbusreq2_p & v374610e | !hbusreq2_p & v8455ab;
assign v3738a2a = hbusreq7_p & v3763813 | !hbusreq7_p & v3a6d88e;
assign v37646a9 = hmaster2_p & v3a635ea | !hmaster2_p & v37697a3;
assign v3769e49 = hmaster2_p & v3736026 | !hmaster2_p & v377e19d;
assign v3725827 = hgrant4_p & v375da10 | !hgrant4_p & v3a5aacb;
assign v3756b78 = hbusreq6 & v35772c9 | !hbusreq6 & v8455ab;
assign v372706d = stateG10_1_p & v2aca977 | !stateG10_1_p & v3a6ee22;
assign v3a5b979 = hmaster1_p & v377f45d | !hmaster1_p & v3759c8c;
assign v3745cc6 = hmaster2_p & v3a70f68 | !hmaster2_p & v377f734;
assign v37688d1 = hmaster2_p & v372b881 | !hmaster2_p & v3a53e66;
assign v3a6a156 = hbusreq8_p & v375c9a3 | !hbusreq8_p & v3a6f6e1;
assign v3a6fd34 = hgrant6_p & v374cb44 | !hgrant6_p & v3737c6c;
assign v3760e7b = hbusreq1_p & v3735826 | !hbusreq1_p & v3a58fef;
assign v37c0296 = hlock5_p & v3a6eb3e | !hlock5_p & v9a3ffa;
assign v376e17e = hlock4_p & v3763295 | !hlock4_p & v8455cb;
assign v375db7f = hlock6_p & v373006f | !hlock6_p & !v8455ab;
assign v376054c = hbusreq7 & v3774f39 | !hbusreq7 & v3768082;
assign v37788ca = hlock0_p & v37682c6 | !hlock0_p & v380989b;
assign v3a705cc = hmaster0_p & v37368c8 | !hmaster0_p & v8455e7;
assign v3766acb = hmaster0_p & v3a635ea | !hmaster0_p & v3a668da;
assign v3a5b4be = hgrant6_p & v3729127 | !hgrant6_p & v3a70409;
assign v374fda4 = hgrant2_p & v374a6fc | !hgrant2_p & v3a6c243;
assign v3a6f998 = hgrant4_p & v3a567ec | !hgrant4_p & v3a61a76;
assign v3a6fa3a = hmaster2_p & v3a70147 | !hmaster2_p & v3809a6a;
assign v376323b = hmaster1_p & v373ad69 | !hmaster1_p & v3738a63;
assign v3734778 = hbusreq6_p & v372cdc9 | !hbusreq6_p & v3a6fc60;
assign v377463a = hbusreq4_p & v2ff9291 | !hbusreq4_p & v3777955;
assign v373a542 = hbusreq6 & v37290af | !hbusreq6 & v8455ab;
assign v3a64868 = hgrant5_p & v3a626da | !hgrant5_p & v3741d7c;
assign v37542a0 = hbusreq5 & v3a5ef9d | !hbusreq5 & v375e512;
assign v3a6f8f6 = hbusreq6_p & v373c965 | !hbusreq6_p & v8455bb;
assign v375c334 = hbusreq6_p & v3a6f8f5 | !hbusreq6_p & v374df14;
assign v3a68e10 = hmaster1_p & v3a6b17e | !hmaster1_p & v375d1d4;
assign v3727823 = hlock8 & v3761f4e | !hlock8 & v3a5d03e;
assign v37352dc = hmaster1_p & v3730e7d | !hmaster1_p & v3a6fa53;
assign v37247cf = hmaster2_p & v374eab4 | !hmaster2_p & v376b4ad;
assign v3732f66 = hbusreq3_p & v3a708af | !hbusreq3_p & v37556cb;
assign v3a71015 = hbusreq5 & v38070c7 | !hbusreq5 & v3a70d99;
assign v3a6b100 = hmaster2_p & v9bf1d8 | !hmaster2_p & v3727e66;
assign v3a6e8d2 = hbusreq4_p & v37704dc | !hbusreq4_p & v377ceea;
assign v8fa780 = hbusreq8 & v372f649 | !hbusreq8 & v8455ab;
assign v3a6134b = hgrant6_p & v8455ab | !hgrant6_p & v3a70a87;
assign v3a70578 = hmaster1_p & v3a635ea | !hmaster1_p & v373a09f;
assign v3759203 = hgrant8_p & a4e409 | !hgrant8_p & v3750553;
assign v3a61820 = hlock7 & v372ce1e | !hlock7 & v377c0c3;
assign v375372b = hmaster1_p & v37597f4 | !hmaster1_p & v3757a04;
assign v3a7048e = hbusreq4_p & v372e096 | !hbusreq4_p & !v3774f3b;
assign v377d080 = hbusreq5_p & v376a8be | !hbusreq5_p & v3a6be50;
assign v372fc07 = hbusreq4 & v3a6fdb0 | !hbusreq4 & v3748797;
assign v37692dc = hlock5 & v373301a | !hlock5 & a19873;
assign v37798bd = hbusreq7_p & v3809d8e | !hbusreq7_p & v3722968;
assign v3777870 = hbusreq3 & v3a57cb4 | !hbusreq3 & v8455ab;
assign v3722f88 = hgrant0_p & v8455ab | !hgrant0_p & !v37746d7;
assign v3a545c8 = hlock7_p & v3778674 | !hlock7_p & !v3257354;
assign v3a711f1 = hgrant1_p & v3a693bf | !hgrant1_p & !v8455ab;
assign v374b15d = hbusreq0 & v37778e2 | !hbusreq0 & v3a6ff1a;
assign v3736d47 = hgrant4_p & v3a635ea | !hgrant4_p & v23fe0c2;
assign v373d993 = hmaster2_p & v3a635ea | !hmaster2_p & v3a54eae;
assign v3755e64 = hmaster0_p & v373b03b | !hmaster0_p & v372ee6a;
assign v3a70652 = hmaster1_p & v3a6ffae | !hmaster1_p & v3776abb;
assign v3a6f5c6 = hbusreq5_p & v8dfd63 | !hbusreq5_p & v37627a2;
assign v373db92 = hbusreq8 & v3736257 | !hbusreq8 & v3748c3f;
assign v372c53a = hmaster2_p & v3a635ea | !hmaster2_p & v377db14;
assign v3763ca1 = hmaster1_p & v372b1dc | !hmaster1_p & v373d029;
assign v3753f17 = hbusreq2_p & v376ea4a | !hbusreq2_p & !v3728e09;
assign v37538ca = hlock5_p & v37558c7 | !hlock5_p & v375456e;
assign v373929f = hbusreq2 & v3766df9 | !hbusreq2 & v8455ab;
assign v376c784 = hmaster1_p & v375637c | !hmaster1_p & !v37605ab;
assign v3a5bdd2 = hgrant4_p & v377a617 | !hgrant4_p & v3756cf0;
assign v373afe9 = hlock5 & v3758c3d | !hlock5 & v3759263;
assign v380971d = hlock5_p & v374d94e | !hlock5_p & v3755af9;
assign v372e741 = hbusreq5_p & v377ee7c | !hbusreq5_p & v3743fc1;
assign v3740fe0 = hbusreq2 & v376bb88 | !hbusreq2 & v3a70a7f;
assign v3762a26 = hmaster0_p & v3775dbc | !hmaster0_p & v373a6ba;
assign v3753b90 = hgrant3_p & v8455ab | !hgrant3_p & v374bc77;
assign db903b = hbusreq6 & v3a5ef89 | !hbusreq6 & v3a641d5;
assign v3a69fe0 = hmaster1_p & v3a6b27d | !hmaster1_p & v37300e3;
assign v3729513 = hgrant0_p & v3741d2d | !hgrant0_p & !v3773a9d;
assign v373086c = hbusreq2 & v8455b0 | !hbusreq2 & v373cc68;
assign v3a6acbb = hgrant0_p & v3a60787 | !hgrant0_p & v37393cc;
assign v3a56d3a = hbusreq8 & v375790e | !hbusreq8 & !v37281a4;
assign v374d43f = hmaster2_p & v372e711 | !hmaster2_p & v374db6a;
assign v3749bf0 = hgrant6_p & v37496fa | !hgrant6_p & v3377b1b;
assign v3752fe9 = hlock3_p & v380713a | !hlock3_p & !v8455ab;
assign v374ed80 = hmaster3_p & v3762c8e | !hmaster3_p & v3770a1c;
assign v3a70905 = hlock6 & v376f584 | !hlock6 & v3a65827;
assign v373aa23 = hlock0_p & v3a635ea | !hlock0_p & v372e474;
assign v3758559 = hbusreq7 & v3a555e5 | !hbusreq7 & v3a6fb8a;
assign v3774a9c = hmaster2_p & v375ce98 | !hmaster2_p & v372abd8;
assign v372f309 = hbusreq0 & v372dccf | !hbusreq0 & v8455ab;
assign v37539ef = hgrant4_p & v209310e | !hgrant4_p & v3740db1;
assign v3a70f2e = hbusreq7 & v3a5a5c4 | !hbusreq7 & v3a71535;
assign v3a6e846 = hmaster2_p & v374d4e6 | !hmaster2_p & v3767848;
assign v3753837 = hgrant4_p & v3a6ff30 | !hgrant4_p & v37600da;
assign v3a61535 = hbusreq0 & v375ba37 | !hbusreq0 & v3a64225;
assign v3729004 = hbusreq6_p & v373f058 | !hbusreq6_p & v3753dab;
assign v375d5e1 = hlock7 & v23fdf14 | !hlock7 & v3a6f750;
assign v35b7b3b = hmaster0_p & v3a65c2a | !hmaster0_p & v37270b9;
assign v373f1d4 = hmaster1_p & v3a6ffca | !hmaster1_p & v377a337;
assign v374bc27 = hlock6 & v3754ec0 | !hlock6 & v3768ef1;
assign v375b65b = hbusreq3_p & v3737c13 | !hbusreq3_p & v3a5cd20;
assign v37355e3 = hlock7 & v375ac88 | !hlock7 & v1e373d9;
assign v3a70ea5 = hbusreq5 & v372c676 | !hbusreq5 & v3746bce;
assign v374763e = hlock7_p & v377664f | !hlock7_p & v3737897;
assign v3a6fd5c = hbusreq6 & v37482f8 | !hbusreq6 & !v3a705f0;
assign v3744f37 = jx0_p & v3806db2 | !jx0_p & v376a74a;
assign v3728608 = hbusreq1 & v37282cf | !hbusreq1 & !v8455ab;
assign v3758663 = hbusreq8_p & v3a704b3 | !hbusreq8_p & v3768036;
assign v3741a9b = hgrant3_p & v3754076 | !hgrant3_p & !v37390ed;
assign v372b61a = hbusreq7 & dc5778 | !hbusreq7 & v376a7da;
assign v373c38b = hmaster1_p & v3a564d9 | !hmaster1_p & v373adb9;
assign v373ad16 = hlock0 & v3a6f3c6 | !hlock0 & v3a63299;
assign v3a70899 = hmaster2_p & v3a6fffd | !hmaster2_p & v8455ab;
assign v375a41b = hbusreq6 & v3a60008 | !hbusreq6 & v374a637;
assign v375a202 = hmaster2_p & v8455ab | !hmaster2_p & v37658f9;
assign v8b1055 = hmaster0_p & v3767b70 | !hmaster0_p & v3774438;
assign v376ddfb = hbusreq2_p & v3777a7e | !hbusreq2_p & v373a188;
assign v3a5e874 = hbusreq8 & v8455e7 | !hbusreq8 & v3a5bb57;
assign v3757f09 = hmaster2_p & v8455ab | !hmaster2_p & v375604f;
assign v372b231 = hbusreq6_p & v37293ee | !hbusreq6_p & v8455ab;
assign v374affb = hgrant6_p & v372493b | !hgrant6_p & v3722f3b;
assign v3a6b768 = hmaster0_p & v3a6efc1 | !hmaster0_p & v8455ab;
assign v377cd7f = hgrant5_p & v8455ab | !hgrant5_p & v3a70baf;
assign v377a470 = hlock5_p & v374d042 | !hlock5_p & v3258dd9;
assign v3a5da57 = hgrant2_p & v3a632f4 | !hgrant2_p & v3743698;
assign v3a6fa6f = hbusreq6_p & v37395bc | !hbusreq6_p & v3737acd;
assign v3775942 = hmaster0_p & v37447df | !hmaster0_p & !v372f1d4;
assign v3773b18 = hmaster2_p & v35b774b | !hmaster2_p & v3a6f213;
assign v374f4a3 = hbusreq4_p & v3778492 | !hbusreq4_p & v3725931;
assign v3724aa0 = hmaster0_p & v377a7f8 | !hmaster0_p & !v3761c61;
assign v37264a2 = hbusreq5_p & v3a5ee85 | !hbusreq5_p & v373d2e3;
assign v372f173 = hmaster2_p & v3a6efe8 | !hmaster2_p & v374c5b2;
assign v373bda7 = hlock0 & v3a630dc | !hlock0 & v375c4ac;
assign v37274e6 = hlock8 & v375e093 | !hlock8 & v3a70a16;
assign v3a63d22 = hmaster2_p & v3a67d8d | !hmaster2_p & v375107e;
assign v3762651 = hbusreq5 & v376a6f1 | !hbusreq5 & v377e345;
assign v373aa96 = hmaster2_p & v3777da6 | !hmaster2_p & v3a6ef01;
assign v37788d7 = hgrant7_p & v3a66039 | !hgrant7_p & v3a570a0;
assign v3764a07 = hbusreq4 & v376e5fe | !hbusreq4 & v3809ec3;
assign v37303aa = jx0_p & v372d24d | !jx0_p & v377504f;
assign v374a3c5 = hbusreq6 & v2acaf41 | !hbusreq6 & v3a714b2;
assign v23fde69 = hlock5_p & v372a02b | !hlock5_p & !v8455ab;
assign v375b143 = hbusreq6_p & v3a5a2be | !hbusreq6_p & v37461e1;
assign v3a5cc4c = hgrant3_p & v37434d6 | !hgrant3_p & v3a5d356;
assign v376cd8f = hbusreq8 & v3762712 | !hbusreq8 & v3a6f0c6;
assign v3766669 = hmaster2_p & v37480b7 | !hmaster2_p & !v3a66910;
assign v374f0f1 = hmaster1_p & v3a6f443 | !hmaster1_p & v3a6b285;
assign v3a6fa5e = hgrant3_p & v3759842 | !hgrant3_p & v3730cc8;
assign v376cc1b = hbusreq6 & v37474b8 | !hbusreq6 & v3a70d64;
assign v3763105 = hlock7 & v376739e | !hlock7 & v3734a80;
assign v3772828 = hgrant6_p & v3a6f3d9 | !hgrant6_p & v37719c6;
assign v374fb40 = hlock6 & v374de48 | !hlock6 & v3a713f4;
assign v3a700d8 = hgrant4_p & v8455ab | !hgrant4_p & v3739f29;
assign v3774492 = hmaster2_p & v372edf8 | !hmaster2_p & v9bf1d8;
assign v3779a66 = hbusreq5_p & v38076c9 | !hbusreq5_p & !v3a6b6f2;
assign v373ab15 = hgrant6_p & v374fafa | !hgrant6_p & v3776e8b;
assign v3a6f475 = hmaster2_p & v373891b | !hmaster2_p & v8455ab;
assign v3751c54 = hmaster1_p & v3768995 | !hmaster1_p & v375a4f8;
assign v3a715d6 = hmaster0_p & v3750cae | !hmaster0_p & !v3778277;
assign v3731d67 = hmaster2_p & v3a70130 | !hmaster2_p & v3769c7f;
assign v377437a = hgrant0_p & v3748797 | !hgrant0_p & v8455ab;
assign v3a5bf99 = hgrant2_p & v8455ba | !hgrant2_p & v3a61d5f;
assign v376a246 = hlock4_p & v3755608 | !hlock4_p & v8455ab;
assign v2092bdc = hbusreq4_p & v377506b | !hbusreq4_p & v3727084;
assign v3a7088b = hmaster0_p & v377a352 | !hmaster0_p & v3741357;
assign v3a57e6d = hmaster2_p & v3736ded | !hmaster2_p & v23fe0be;
assign v3773530 = hmaster1_p & v3777bfc | !hmaster1_p & v37415c3;
assign v3777988 = hgrant5_p & v8455ab | !hgrant5_p & v3a6da08;
assign v373ca5f = hmaster2_p & v3a71601 | !hmaster2_p & v37539ef;
assign v3740140 = hbusreq3 & v374362e | !hbusreq3 & v3a676d6;
assign d9a7db = hbusreq2 & v3771e95 | !hbusreq2 & v3a6a393;
assign v374c6df = hlock1_p & v3739d51 | !hlock1_p & v3a60c77;
assign v376a7e8 = hbusreq2_p & v3a6f989 | !hbusreq2_p & v3a2981b;
assign v3726458 = hmaster2_p & v3772e0c | !hmaster2_p & v3770027;
assign v3745ce4 = hbusreq4_p & v3a6677e | !hbusreq4_p & v377aa06;
assign v37637d6 = hgrant3_p & v376f0c1 | !hgrant3_p & v373adae;
assign v3a5f281 = hmaster2_p & v374314f | !hmaster2_p & v373366b;
assign v3755082 = hbusreq5_p & v8455ab | !hbusreq5_p & v375ecf8;
assign v3378a34 = hbusreq2 & v372f76a | !hbusreq2 & v3a67aaa;
assign v377f812 = hbusreq2_p & v3a71528 | !hbusreq2_p & !v3a5b68a;
assign v3a57b70 = hlock6 & v3378594 | !hlock6 & v37440a8;
assign v3a6a25c = hbusreq8_p & v375fb71 | !hbusreq8_p & v3756526;
assign v3733b02 = hmaster1_p & v9c1340 | !hmaster1_p & v3757272;
assign v374bb56 = hbusreq3 & v373fe5e | !hbusreq3 & !v376430b;
assign v3a6afdd = hmaster2_p & v3a6f806 | !hmaster2_p & v3a5a158;
assign v39af33c = jx2_p & v372bc78 | !jx2_p & !v3a61a1d;
assign v3a70a4c = hbusreq2 & v377881b | !hbusreq2 & v3a70c74;
assign v37690f3 = hbusreq0 & v3a63331 | !hbusreq0 & v3741bb2;
assign v3a70737 = hbusreq3_p & v377eb2d | !hbusreq3_p & v8455b0;
assign v373dc1c = hlock0_p & v373fe5e | !hlock0_p & !v8455ab;
assign v376e72d = hbusreq6_p & v373cb54 | !hbusreq6_p & v8455ab;
assign v377a9cb = hgrant6_p & v8455ab | !hgrant6_p & v37574b0;
assign v375d77d = hmaster2_p & v37513fa | !hmaster2_p & v3a706e4;
assign v3727f14 = hbusreq4_p & v3a5a573 | !hbusreq4_p & v8455ab;
assign v3a6d407 = hmaster2_p & v3a6d71b | !hmaster2_p & v3758df6;
assign v3731088 = hbusreq5_p & v377e328 | !hbusreq5_p & v373f6cf;
assign v375626c = hgrant4_p & v374e849 | !hgrant4_p & v372fe8b;
assign v375c0d6 = hmaster2_p & v3a70374 | !hmaster2_p & v3a55419;
assign v3767dc8 = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v372f071;
assign v3a70a95 = hgrant2_p & v3a70dc4 | !hgrant2_p & v3a701d3;
assign v3767f33 = hbusreq1_p & v3740171 | !hbusreq1_p & v37270d9;
assign v3756ba5 = hmaster1_p & v3a6b27d | !hmaster1_p & v3728435;
assign v374139a = jx0_p & v8455ab | !jx0_p & v374c2e1;
assign v3731415 = hmaster2_p & v8455ab | !hmaster2_p & v376e16e;
assign v376aae5 = hbusreq5 & v374f3ad | !hbusreq5 & v3a70dcb;
assign v374c91a = hbusreq6_p & v3745452 | !hbusreq6_p & v8455b0;
assign v39a4d8a = hmaster2_p & v3752fe6 | !hmaster2_p & v3729f14;
assign v2093252 = hbusreq5_p & v37682ce | !hbusreq5_p & v8455ab;
assign v373b837 = hmaster1_p & v375a510 | !hmaster1_p & v372af06;
assign v3a703a4 = hbusreq3_p & v372b765 | !hbusreq3_p & !v3a640c5;
assign v3723ddc = hmaster1_p & v372d905 | !hmaster1_p & v372fb3c;
assign v3754903 = hgrant2_p & v8455ab | !hgrant2_p & v373b4ad;
assign v92391b = hbusreq8 & v3a6eee7 | !hbusreq8 & v375da55;
assign v377fabb = hbusreq4_p & v375d00a | !hbusreq4_p & v3763b0a;
assign v37547f7 = hlock7_p & v3a673d9 | !hlock7_p & v8455ab;
assign v375501e = hbusreq4_p & v3745539 | !hbusreq4_p & v373769f;
assign v375bb10 = hmaster2_p & v3745a5f | !hmaster2_p & v3777a00;
assign v3753c2a = hgrant4_p & v377d354 | !hgrant4_p & v8455ab;
assign v3727d7e = hmaster2_p & v3a6f43e | !hmaster2_p & v376ea4a;
assign v3a6fd98 = hmaster0_p & v374fe9d | !hmaster0_p & v373185b;
assign v37513bc = hlock4 & v37759b5 | !hlock4 & v372cb44;
assign v3a713d1 = hmaster1_p & v3739fb8 | !hmaster1_p & v3731684;
assign v376025c = hmaster1_p & v375121b | !hmaster1_p & v37418bf;
assign v37551eb = hmaster1_p & v376086c | !hmaster1_p & v3a53fb5;
assign v375de66 = hbusreq8 & v3755783 | !hbusreq8 & v3753f35;
assign v3751db0 = hbusreq1_p & v20d166d | !hbusreq1_p & v8455ab;
assign v3a7143f = hbusreq3_p & v3760073 | !hbusreq3_p & v3a640c5;
assign v373f6d5 = hbusreq4 & v3a5dc82 | !hbusreq4 & v3760ff4;
assign v377d9b2 = hgrant5_p & v373ad69 | !hgrant5_p & v3735f67;
assign v37510d7 = hbusreq8_p & v3740742 | !hbusreq8_p & v23fd9af;
assign v3a70dbb = hlock5 & v3739748 | !hlock5 & v3a58378;
assign v3737fca = hmaster0_p & v372eb5c | !hmaster0_p & v37390c9;
assign v3754bb9 = jx0_p & v3a68af5 | !jx0_p & v3773daf;
assign v372af46 = hbusreq2 & v37395e6 | !hbusreq2 & v8455e7;
assign v3a63dcc = hlock2 & v375fbe8 | !hlock2 & v380930a;
assign v3733168 = hmaster0_p & v376c208 | !hmaster0_p & !v8455ab;
assign v3a6254e = hlock1_p & v375bc4b | !hlock1_p & v8455ab;
assign v3769c72 = hbusreq7_p & v3a6f270 | !hbusreq7_p & v377981b;
assign v37446d8 = hbusreq5 & v375f87a | !hbusreq5 & v377de07;
assign v375527f = hbusreq5_p & v3a70990 | !hbusreq5_p & v3731d06;
assign v3727bc1 = hbusreq5 & v3a70572 | !hbusreq5 & v3a2a107;
assign v3740bb4 = hbusreq4 & v375df95 | !hbusreq4 & v37285eb;
assign v373e553 = hmaster0_p & v375db57 | !hmaster0_p & v372a520;
assign locked = v3a6757a;
assign v3a5d3af = hlock6_p & v3777311 | !hlock6_p & adf78a;
assign v3749942 = hmaster1_p & v1e38283 | !hmaster1_p & v373aee6;
assign v3763d77 = hlock6 & v3a68ed1 | !hlock6 & v372b89e;
assign v3728a53 = hmaster1_p & v373b6ee | !hmaster1_p & v3778c14;
assign v3a66a3b = hlock4_p & v376dd3d | !hlock4_p & v37573f4;
assign v376fc09 = hbusreq5 & v3806def | !hbusreq5 & v37bfc97;
assign v375b880 = hgrant4_p & v374d0e3 | !hgrant4_p & v375aea6;
assign v3773a84 = hbusreq4 & v37406d2 | !hbusreq4 & v8455ab;
assign v3a6fd66 = hbusreq5 & v377c0d5 | !hbusreq5 & v8455ab;
assign v377f4bb = stateA1_p & v376faea | !stateA1_p & v372dee5;
assign v3736a92 = hgrant0_p & v37773a9 | !hgrant0_p & v3a6b2ef;
assign v376726e = hgrant7_p & v8455ab | !hgrant7_p & !b69f28;
assign v3a70937 = hbusreq6 & v3a6fdd6 | !hbusreq6 & v373ea71;
assign v3a709b5 = hmaster1_p & v37533c8 | !hmaster1_p & v372f9b4;
assign v375a4c4 = hbusreq7_p & v3a70176 | !hbusreq7_p & v373178d;
assign v373d26a = hmaster1_p & v3a6ff25 | !hmaster1_p & v375415d;
assign v3a704bf = hbusreq5_p & v3734c40 | !hbusreq5_p & v377ba8e;
assign v3a5621f = hlock0 & v3748797 | !hlock0 & v377c023;
assign v37731ce = hgrant4_p & v3770032 | !hgrant4_p & v3a5ad1d;
assign v37434c6 = hmaster2_p & v37430e7 | !hmaster2_p & v8455b3;
assign v3a70f01 = hgrant3_p & v3a70737 | !hgrant3_p & v8455ab;
assign v3748829 = hmaster0_p & v8455ab | !hmaster0_p & v3a53a8a;
assign v3809388 = hmaster0_p & v3a70c3e | !hmaster0_p & v3a6fd0a;
assign v3a6f110 = hlock0_p & v3a568f7 | !hlock0_p & v3723cc2;
assign v372de49 = hmaster3_p & v3733392 | !hmaster3_p & v3768ac9;
assign v2092b5f = hmaster1_p & v37349e4 | !hmaster1_p & v8455ab;
assign v374005b = hbusreq3_p & v3750025 | !hbusreq3_p & v3a70888;
assign v3a70069 = hready_p & ce3eb4 | !hready_p & !v373281b;
assign v3a71094 = hgrant5_p & v8455c6 | !hgrant5_p & v3a53d44;
assign v37740d0 = hbusreq2_p & v377834b | !hbusreq2_p & v3a6f8de;
assign v3a64c6b = hgrant5_p & v3a58980 | !hgrant5_p & v3a70686;
assign v3577416 = hgrant3_p & v3a5e24e | !hgrant3_p & v3768ab0;
assign v3a66c49 = hlock8_p & v377f2bb | !hlock8_p & v2092eb6;
assign v37414b0 = hbusreq6_p & v3a6480b | !hbusreq6_p & v3a70b2c;
assign v376674a = hbusreq2_p & v3749380 | !hbusreq2_p & v3a71646;
assign v3a65bb5 = hbusreq0_p & cf3b5d | !hbusreq0_p & v372998c;
assign v3734aa5 = hmaster1_p & v3a58218 | !hmaster1_p & v3772140;
assign v375e527 = hbusreq0 & v375d134 | !hbusreq0 & v3a6d81d;
assign v3a633bf = hmaster0_p & v3724da7 | !hmaster0_p & v3770db3;
assign v3a6605d = hmaster2_p & v3a71678 | !hmaster2_p & v3a711f9;
assign v3730e54 = hgrant6_p & v8455ab | !hgrant6_p & v3a6ef75;
assign v3a6fb2f = hmaster0_p & v3a62542 | !hmaster0_p & v377c8d1;
assign v3739938 = hmaster0_p & v3762455 | !hmaster0_p & !v3a6f6cf;
assign v3729ca6 = hbusreq5_p & v3a70ce4 | !hbusreq5_p & v8455ab;
assign v37463bc = hbusreq2 & v3a6ab5f | !hbusreq2 & !v3748900;
assign v374e35e = hready & v373a0bf | !hready & v8455ab;
assign v3a70178 = hgrant2_p & v8455ab | !hgrant2_p & v376e677;
assign v3729852 = hbusreq6_p & v39a5381 | !hbusreq6_p & v372d2ad;
assign v3a6fea3 = hbusreq3_p & v3775ee8 | !hbusreq3_p & v3a6a8c5;
assign v3774372 = hlock8 & v3754445 | !hlock8 & v376b4d4;
assign v3a626e4 = hbusreq0 & v3a71454 | !hbusreq0 & v8455ab;
assign v3741fea = jx1_p & v3763afe | !jx1_p & v8455ab;
assign v3745d9c = hmaster2_p & v375afe9 | !hmaster2_p & v3a6866f;
assign v3769f0f = hgrant2_p & v37699a0 | !hgrant2_p & v373f23c;
assign v376a755 = hmaster0_p & v3a70209 | !hmaster0_p & v377fb81;
assign v374cfd9 = hlock5_p & v3774200 | !hlock5_p & v374893c;
assign v373dd27 = hgrant6_p & v3a70240 | !hgrant6_p & v375de2d;
assign v3731210 = hbusreq0 & v3a6fcb9 | !hbusreq0 & v8455ab;
assign v3762ec5 = jx1_p & v37555cb | !jx1_p & v3a675b2;
assign v3a70605 = hbusreq8_p & v3766664 | !hbusreq8_p & !v3a6f9b6;
assign v3723dc3 = hmaster2_p & v8455b7 | !hmaster2_p & v3a6a261;
assign v3a5f6da = hlock5 & v37261ad | !hlock5 & v3a65e55;
assign v3a6f326 = hlock0 & v3a67f97 | !hlock0 & v3a704e7;
assign v1e37c44 = hbusreq7_p & v3a69063 | !hbusreq7_p & v3767919;
assign v372e47b = hmaster1_p & v3764276 | !hmaster1_p & v3742a8b;
assign v3772e4f = hlock5 & v3725ba5 | !hlock5 & v373497f;
assign v3378992 = hlock5_p & v374cceb | !hlock5_p & !d1375e;
assign v3a6816a = hgrant0_p & v8455e7 | !hgrant0_p & v3a6f40c;
assign v372c029 = hgrant4_p & v3725230 | !hgrant4_p & v375cbe3;
assign v376eb33 = hmaster2_p & v37745c3 | !hmaster2_p & v372d2dc;
assign v3765008 = hlock5 & v3751e62 | !hlock5 & v3768e0e;
assign v3754c4a = hbusreq7 & v3771f50 | !hbusreq7 & v3734279;
assign v376fe30 = hgrant0_p & v37773a9 | !hgrant0_p & v2aca784;
assign v3752ade = hmaster2_p & v3a6fe18 | !hmaster2_p & v8455ab;
assign v376c5de = hmaster0_p & v3a5a39f | !hmaster0_p & !v37590f4;
assign v37283bb = hbusreq6_p & v3747302 | !hbusreq6_p & v3a70b92;
assign v37563eb = busreq_p & v8455ab | !busreq_p & v373b003;
assign v375fecf = hlock8 & v3737808 | !hlock8 & v3750559;
assign v3727699 = hmaster1_p & v376f979 | !hmaster1_p & v377d080;
assign v37711cd = hbusreq8_p & v375b84e | !hbusreq8_p & v3a69203;
assign v3740be8 = hbusreq8 & v376fb07 | !hbusreq8 & v3734279;
assign v3a68fc9 = hbusreq6_p & v3748609 | !hbusreq6_p & !v3732569;
assign v372462b = hgrant2_p & v3a5b6de | !hgrant2_p & v37366b5;
assign v3a63c12 = hbusreq5 & v3a6eb19 | !hbusreq5 & v8455ab;
assign v3a71689 = hbusreq2 & v3a67e64 | !hbusreq2 & !v3746fce;
assign v3725d79 = hmaster2_p & v3a66110 | !hmaster2_p & v376d856;
assign v3a6f35f = hlock0 & v3a64af7 | !hlock0 & v3a7026f;
assign v3a6eb40 = hmaster1_p & v3723ec6 | !hmaster1_p & v3a6ec0b;
assign v373f8a7 = hbusreq0 & v3723dae | !hbusreq0 & v3a5a057;
assign v377b086 = hbusreq2_p & v8455ab | !hbusreq2_p & v3809a76;
assign v3a5ca44 = hbusreq0 & v377135e | !hbusreq0 & v3730e54;
assign v3756d07 = hbusreq2 & v3a6b6f3 | !hbusreq2 & !v8455ab;
assign v373a90e = hlock4 & v3a70525 | !hlock4 & v373b50e;
assign v372641e = hgrant5_p & v3a54ac1 | !hgrant5_p & v377a681;
assign v3753001 = hbusreq0 & v3724048 | !hbusreq0 & v3a61344;
assign v3a70c96 = hbusreq2 & v375e551 | !hbusreq2 & v8455ab;
assign v374a233 = hgrant4_p & v3a53eeb | !hgrant4_p & v3a70b39;
assign v375f74e = hbusreq4 & v3a7084e | !hbusreq4 & v8455bb;
assign v3731859 = hbusreq6_p & v3a7039b | !hbusreq6_p & v8455e7;
assign v3a63d3c = hgrant6_p & v376ea4a | !hgrant6_p & v3a5aa9d;
assign v3a64c73 = jx2_p & v377e7f8 | !jx2_p & !v3806828;
assign v3753940 = hgrant6_p & v377f09a | !hgrant6_p & v374d7dd;
assign v373a756 = hmaster2_p & v375c675 | !hmaster2_p & v374693f;
assign v3730bf5 = hgrant2_p & v376004c | !hgrant2_p & v3a70799;
assign v3a6f791 = hmaster1_p & v3a6f6bf | !hmaster1_p & v37249ff;
assign v3a704fb = hlock7 & v3736515 | !hlock7 & v373c228;
assign v3776f42 = hmaster2_p & v3a67d66 | !hmaster2_p & v8455bb;
assign v373f410 = hgrant4_p & v377015c | !hgrant4_p & v37276f2;
assign v3757d75 = hmaster2_p & v3a6fc74 | !hmaster2_p & ce4abb;
assign v376ebc7 = jx1_p & v3a674d5 | !jx1_p & v3767d2c;
assign v3577487 = hgrant5_p & v3a715e9 | !hgrant5_p & v3a6ec88;
assign v3a5b614 = hgrant3_p & v38072fd | !hgrant3_p & v8455ab;
assign v3a6f4f3 = hmaster0_p & v3a6d1a5 | !hmaster0_p & v372700a;
assign v374e1fd = hlock5_p & v3a6f942 | !hlock5_p & v372580e;
assign v376739e = hbusreq7 & v3734a80 | !hbusreq7 & v373abcf;
assign v3a6fa50 = hbusreq6 & v3a696ed | !hbusreq6 & v8455ab;
assign v3777ee7 = hmaster2_p & v374e079 | !hmaster2_p & v35772a6;
assign v8d3fe3 = hmaster1_p & v373e91a | !hmaster1_p & v3a571de;
assign v35d37b1 = jx2_p & v372bc78 | !jx2_p & !v3737672;
assign v3723025 = hmaster1_p & v374c6b8 | !hmaster1_p & v3a713da;
assign v3776ca9 = hmaster2_p & v3744bfc | !hmaster2_p & !v8455ab;
assign v375ae91 = hbusreq0 & v3a6ef4d | !hbusreq0 & v3a6f44e;
assign v377f5db = hmaster2_p & v23fe361 | !hmaster2_p & v8455ab;
assign v3a70715 = hbusreq2 & v3a61cbf | !hbusreq2 & v3a708c2;
assign v373754d = hbusreq7_p & v3a71591 | !hbusreq7_p & v3722e49;
assign v3a61a3d = hbusreq2 & v8455e7 | !hbusreq2 & v8455ab;
assign v3a61c51 = hmaster2_p & v373a27c | !hmaster2_p & v37457fb;
assign v3763327 = hbusreq4_p & v3a7084c | !hbusreq4_p & v8455b0;
assign v37346dc = hlock4 & v3a57658 | !hlock4 & v3747bea;
assign v3769f84 = hbusreq6_p & v375084d | !hbusreq6_p & v3a6fddd;
assign v3a5604a = hbusreq5 & v373ee81 | !hbusreq5 & v3764ee3;
assign v3779746 = hlock6 & v377550d | !hlock6 & v3a6ff2d;
assign v3a70a64 = hmaster3_p & v8455ab | !hmaster3_p & v374828c;
assign v37548c4 = hmaster2_p & v3a6a8ee | !hmaster2_p & d5f283;
assign v3a70907 = hmaster3_p & v3a6b2ea | !hmaster3_p & v3a6fb41;
assign v3a701c3 = hbusreq4 & v372879a | !hbusreq4 & v377bfc0;
assign v3a6e09b = hmaster2_p & v37282cf | !hmaster2_p & !v3728e09;
assign v3768fba = hbusreq5 & v3728419 | !hbusreq5 & v8455ab;
assign v3756200 = hmaster1_p & v3a57ee9 | !hmaster1_p & v3773ab1;
assign v372d8f7 = hbusreq4 & v373f836 | !hbusreq4 & v3727084;
assign v374424e = hlock6_p & v376ddc6 | !hlock6_p & v373f503;
assign v375a293 = hbusreq3_p & v38072fd | !hbusreq3_p & v375e22b;
assign v3a5585e = hbusreq4 & v38072f9 | !hbusreq4 & v8455ab;
assign v3727b41 = hbusreq6_p & v3a7037c | !hbusreq6_p & v3746f84;
assign v377d8c8 = hmaster2_p & v372f309 | !hmaster2_p & v377bf71;
assign v372bea3 = hmaster2_p & v3778cf7 | !hmaster2_p & !v3760700;
assign v37332c8 = hbusreq6_p & v3a64112 | !hbusreq6_p & v3806f24;
assign v374abcc = hmaster0_p & v377766c | !hmaster0_p & v3a6f707;
assign v3736f2a = hbusreq6_p & v374a192 | !hbusreq6_p & v3a70fdf;
assign v3a6f298 = jx0_p & v8e3f65 | !jx0_p & v3723809;
assign v377ba5a = hgrant3_p & v8455ab | !hgrant3_p & v3a68523;
assign v377a65c = jx1_p & v37573d2 | !jx1_p & v3a675b2;
assign v37461e1 = hgrant2_p & v8455ab | !hgrant2_p & v3724392;
assign v3749ddf = hbusreq6 & v3a54853 | !hbusreq6 & !v3a70abc;
assign v3a668e4 = hmaster0_p & v3a5f08f | !hmaster0_p & v3a6a8ee;
assign v37650e3 = hgrant2_p & v3a5adfd | !hgrant2_p & a7f6c5;
assign v3a709fb = hmaster0_p & v3a5a223 | !hmaster0_p & v373d076;
assign v37657be = hlock5 & v3763478 | !hlock5 & v372c97c;
assign v373beae = hbusreq5_p & v3742649 | !hbusreq5_p & v3a60d50;
assign v377478a = hmaster1_p & v3a58cfc | !hmaster1_p & v3a706c5;
assign v3774a4b = hbusreq8 & v37515a1 | !hbusreq8 & v380735e;
assign v377bb93 = hmaster2_p & v8455ab | !hmaster2_p & !v3a7092a;
assign v37375f3 = hgrant2_p & v3a66671 | !hgrant2_p & v3807ac6;
assign v3a6f681 = hlock7_p & v37790bd | !hlock7_p & !v8455ab;
assign v372afcc = hbusreq5 & v3754379 | !hbusreq5 & v37759a7;
assign v377a916 = jx0_p & v3739731 | !jx0_p & v37738e9;
assign v376069d = hbusreq8_p & v374478a | !hbusreq8_p & v3a6f7fe;
assign v3a70bbe = hbusreq5_p & v372490a | !hbusreq5_p & !v3a6fc41;
assign v23fdb05 = decide_p & v374cca4 | !decide_p & v375a94d;
assign v374e8a2 = hbusreq5 & v376b40c | !hbusreq5 & v3807729;
assign v376c211 = stateA1_p & v8455ab | !stateA1_p & !v3a7147e;
assign v374c048 = hmaster3_p & v8ce84c | !hmaster3_p & v3750e8a;
assign v3a654af = hbusreq6 & v376b7db | !hbusreq6 & v375b2fe;
assign v3a5fc70 = hmaster0_p & v3749c2f | !hmaster0_p & !v374b1a4;
assign v3728a9f = hgrant4_p & v8455b9 | !hgrant4_p & v377882e;
assign v3a6cdd4 = hgrant6_p & v375f653 | !hgrant6_p & v374fac6;
assign c10173 = hmaster2_p & v377eaf2 | !hmaster2_p & v8455ab;
assign v3a6f2de = hmaster2_p & v3a5fc34 | !hmaster2_p & v8455ab;
assign v373df13 = hbusreq0 & v1e3799d | !hbusreq0 & v3749e13;
assign v3744380 = hlock6_p & v3770415 | !hlock6_p & v8455bb;
assign v3a66c22 = hbusreq8 & v374e3ab | !hbusreq8 & v39a4e7e;
assign v376b307 = hbusreq2_p & v3a5d5d3 | !hbusreq2_p & v8455ab;
assign v375b2af = hmaster0_p & v3728646 | !hmaster0_p & v3760951;
assign v3a65752 = hmaster2_p & c0990a | !hmaster2_p & v374916a;
assign v3779df7 = hmaster2_p & v372745b | !hmaster2_p & v3a6f93a;
assign v3a71064 = hbusreq6 & v39a4e43 | !hbusreq6 & v3a5ee6e;
assign v3a68084 = hbusreq4_p & v377caa3 | !hbusreq4_p & v3755820;
assign v3730aaf = hbusreq4 & v3760f62 | !hbusreq4 & v372cc25;
assign v3772f37 = hmaster3_p & v3a712b5 | !hmaster3_p & v375fc79;
assign v3767a93 = hbusreq0 & v3767d1b | !hbusreq0 & v373e814;
assign v3725ba8 = hlock0_p & v3a5980d | !hlock0_p & v8455b7;
assign v372a902 = hbusreq6_p & v375d9a7 | !hbusreq6_p & v8455ab;
assign v3a65ce5 = hbusreq7_p & v3756a8f | !hbusreq7_p & !v374a37e;
assign v3a53986 = hmaster2_p & v373b11a | !hmaster2_p & v8455ab;
assign v3752dbb = stateG10_1_p & v8455ab | !stateG10_1_p & v3a6fc6c;
assign v3a7000a = hmaster2_p & v3756eaf | !hmaster2_p & v3a66750;
assign v374d218 = hgrant3_p & v375c1d1 | !hgrant3_p & v3a640c5;
assign v3a29d87 = hmaster2_p & v8455ab | !hmaster2_p & !v3a71350;
assign v3a71343 = hbusreq5_p & v374b912 | !hbusreq5_p & v377e056;
assign v373178d = hlock8_p & v8455ab | !hlock8_p & v3a63f6d;
assign v372af57 = hlock4 & v372952d | !hlock4 & v3774acc;
assign v3a70208 = hgrant0_p & v3a637dc | !hgrant0_p & v3a66140;
assign v376be82 = hgrant8_p & v3776413 | !hgrant8_p & v3739fc8;
assign v3a6fdab = hgrant5_p & v3758924 | !hgrant5_p & v373b95e;
assign v37612d0 = hbusreq8 & v8455b0 | !hbusreq8 & v3735da3;
assign v3a6d0ae = hbusreq8_p & v3772dcb | !hbusreq8_p & v3768734;
assign v3734292 = hbusreq4_p & v373bfab | !hbusreq4_p & v375fd8d;
assign v376af2d = hgrant6_p & v377f09a | !hgrant6_p & !v3a694bb;
assign v3a6f90e = hmaster2_p & v375d616 | !hmaster2_p & v3776685;
assign v372f759 = hlock4 & v3760d16 | !hlock4 & v372313c;
assign v3734c0f = hbusreq7_p & v373285a | !hbusreq7_p & v3774058;
assign v374f535 = jx3_p & v3751fde | !jx3_p & v373e2bc;
assign v377da14 = hmaster2_p & v373a4e4 | !hmaster2_p & v376b88d;
assign v376d88f = hmaster1_p & v37782c9 | !hmaster1_p & v372b551;
assign v37645eb = hmaster2_p & dc5fea | !hmaster2_p & v37769cc;
assign v3728cdc = hmaster2_p & v3a70d99 | !hmaster2_p & v8455ab;
assign v3a66a6c = hgrant2_p & v3a70dc4 | !hgrant2_p & v3769de7;
assign v3a6f74f = hlock7_p & v3a63cf5 | !hlock7_p & !v3a69df3;
assign v3a6d30c = hbusreq6_p & v375f462 | !hbusreq6_p & v3747cf5;
assign v3a7090b = hmaster1_p & v376501e | !hmaster1_p & v3a64eac;
assign v374648f = hbusreq4 & v3a5d469 | !hbusreq4 & v3a69487;
assign v37466c1 = hbusreq6_p & v37395bc | !hbusreq6_p & v3a635c3;
assign v374cceb = hmaster0_p & v3a5a510 | !hmaster0_p & v374b13e;
assign v3a6e1ed = hmaster0_p & v37701a0 | !hmaster0_p & v3a553db;
assign v37671b7 = hbusreq4 & v3a70188 | !hbusreq4 & v376bade;
assign v3a656f0 = hbusreq8_p & v373b90b | !hbusreq8_p & !v37590d5;
assign v3a70307 = hlock8 & v374ace9 | !hlock8 & v3746aa9;
assign v38067ea = hbusreq5 & be54b2 | !hbusreq5 & v3769740;
assign v3a61ce7 = hbusreq4 & v3a6fc48 | !hbusreq4 & v3a6bdaa;
assign v37266b1 = hbusreq2 & v377989c | !hbusreq2 & v8455ab;
assign v3a6aefd = hgrant6_p & v374eef1 | !hgrant6_p & v3764218;
assign v373fbb4 = hlock2_p & v8455ab | !hlock2_p & !v3a6b714;
assign v3759ffd = hbusreq2 & v375767e | !hbusreq2 & v373c480;
assign v374314f = hgrant4_p & v374f307 | !hgrant4_p & v3723ace;
assign v3a70500 = hgrant7_p & v372af6d | !hgrant7_p & v3a70064;
assign v376ae41 = hlock4 & v3a6f4fd | !hlock4 & v3a5ab85;
assign v3a6fa45 = hmaster2_p & v373f95b | !hmaster2_p & v3775684;
assign v3a64374 = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a6e4de;
assign v3a71675 = hbusreq8 & v375095e | !hbusreq8 & v373e1cc;
assign v3734331 = hmaster0_p & v373ec38 | !hmaster0_p & d26e1e;
assign v3a587bc = hgrant3_p & v8455ab | !hgrant3_p & v376fc36;
assign v23fdbc1 = hmaster2_p & v374f307 | !hmaster2_p & v8455ab;
assign v375e6b3 = hgrant0_p & v376969b | !hgrant0_p & v3755a10;
assign v37617d4 = hbusreq3_p & v3a70159 | !hbusreq3_p & v3743e56;
assign v3747ac9 = hbusreq0 & v373e4db | !hbusreq0 & v3a63873;
assign v3746ef3 = hlock4 & v37327ee | !hlock4 & v37772db;
assign v3743f2c = hbusreq8 & b44720 | !hbusreq8 & v374148a;
assign v3779797 = hmaster0_p & v374ab22 | !hmaster0_p & v3736fb6;
assign v2092f2c = hlock8 & v373f2fe | !hlock8 & v3731370;
assign v3a6c5e5 = hmaster0_p & v8455ca | !hmaster0_p & !v3a70386;
assign v374a70f = hbusreq2 & v375cade | !hbusreq2 & v8455ab;
assign ad3125 = hgrant6_p & v3a682b1 | !hgrant6_p & v3735bdc;
assign ac1a2c = hbusreq0 & v377db1f | !hbusreq0 & v376047f;
assign v3a58aa5 = stateG10_1_p & v39ebac7 | !stateG10_1_p & v1e38224;
assign v3a572b4 = hgrant6_p & v8455ab | !hgrant6_p & v23fdc46;
assign v373dd8a = hbusreq1 & v3a6a195 | !hbusreq1 & v37496fa;
assign v37785a8 = hbusreq6 & v373c01a | !hbusreq6 & v8455ab;
assign v3755b5e = hbusreq3_p & v372ba4d | !hbusreq3_p & v3a71630;
assign v3a6edb5 = hmaster0_p & v37722a0 | !hmaster0_p & v3a6adff;
assign v3735dae = hbusreq6_p & v3a635ea | !hbusreq6_p & v376bade;
assign v3a5cfb0 = hbusreq5_p & v374801c | !hbusreq5_p & v373ee81;
assign v3779f1e = hmaster1_p & v372a0e3 | !hmaster1_p & v372c23b;
assign v375f1ee = hbusreq0 & v3a6a1df | !hbusreq0 & c7355c;
assign v3a53d12 = hbusreq6_p & v376f2a7 | !hbusreq6_p & v3743b9e;
assign v377b735 = hmaster1_p & v8455ab | !hmaster1_p & !v37793cd;
assign v37669d0 = hlock8 & v376cba1 | !hlock8 & v3a64bb1;
assign v3a565eb = hbusreq2 & v3a6c243 | !hbusreq2 & v8455ab;
assign v3a70f4f = hgrant5_p & v325c974 | !hgrant5_p & v3a669be;
assign v3739d2c = hlock5 & v3734c47 | !hlock5 & v374f077;
assign v3a6d03c = hlock4 & v373e6cf | !hlock4 & v372ea4b;
assign v3a64fb4 = hmaster2_p & v3a5b8b9 | !hmaster2_p & v3a64f7e;
assign v3a56e63 = hbusreq2_p & v39a537f | !hbusreq2_p & !v1e38224;
assign v3776135 = hmaster0_p & v8455b0 | !hmaster0_p & v3775303;
assign v3768931 = hbusreq1_p & v376ebdd | !hbusreq1_p & !v8455ab;
assign v3745428 = hmaster1_p & v3a6f7cd | !hmaster1_p & !v3a5733c;
assign v3737280 = hbusreq6 & v8455b0 | !hbusreq6 & v37406d2;
assign v372eb5b = hmaster1_p & v3750735 | !hmaster1_p & v3a6a68c;
assign v37606b8 = hbusreq4_p & v3a63b57 | !hbusreq4_p & v3772c7d;
assign v3a6aa9f = hbusreq0 & v3a64ad2 | !hbusreq0 & v3761d06;
assign v376992a = hlock6 & v373698b | !hlock6 & v3a6f03f;
assign v3731d80 = stateG2_p & v8455ab | !stateG2_p & !v845605;
assign v3a62bce = hbusreq2 & v3768ecc | !hbusreq2 & v8455ab;
assign v3751acf = hbusreq0 & v375a4fa | !hbusreq0 & v8455ab;
assign stateG10_7 = !v397d860;
assign v372beb6 = hgrant5_p & v372bcf2 | !hgrant5_p & v3a6eab2;
assign v376b14c = hbusreq8_p & v3778b73 | !hbusreq8_p & v375b0f9;
assign v372f012 = hlock2_p & v37575e7 | !hlock2_p & !v8455ab;
assign v3757343 = hmaster2_p & v8455ab | !hmaster2_p & !v3748caf;
assign v376130f = hmaster1_p & v8455e1 | !hmaster1_p & v3752fbe;
assign v3a6f469 = hbusreq5_p & v3a6a1e8 | !hbusreq5_p & v3a61202;
assign v3762333 = hbusreq6 & v3773d82 | !hbusreq6 & v8455ab;
assign v3749ae8 = hbusreq7 & v3743798 | !hbusreq7 & v375c8db;
assign v3a6fbd9 = hlock6_p & v3a6c23b | !hlock6_p & v3a63805;
assign v3a57330 = locked_p & v374f0c1 | !locked_p & v3a6ffae;
assign v3768454 = hbusreq6 & v3a612a9 | !hbusreq6 & v372c35a;
assign v3749c8a = hgrant6_p & v3a56d01 | !hgrant6_p & v3808881;
assign v3774add = hbusreq6_p & v373a4f7 | !hbusreq6_p & v8455ab;
assign v2acaf12 = hgrant5_p & v3a70615 | !hgrant5_p & v3a616cb;
assign v3774b12 = hmaster0_p & v8455ab | !hmaster0_p & !v3723211;
assign v377e288 = hbusreq2 & v3a701e7 | !hbusreq2 & v8455ab;
assign v375ced9 = hbusreq6 & v3a6672b | !hbusreq6 & v8455ab;
assign v376640b = hgrant3_p & v3a637dc | !hgrant3_p & v3a6e236;
assign v37602c4 = hmaster1_p & v3778e3f | !hmaster1_p & v3a70cc7;
assign v376a6ae = hgrant5_p & v372c0de | !hgrant5_p & !v372580c;
assign v3a6624e = hbusreq5 & v3775606 | !hbusreq5 & v3764dac;
assign v3766484 = hgrant4_p & v3744b1b | !hgrant4_p & v37323a1;
assign v3771536 = hlock4_p & v373b3fb | !hlock4_p & v8455b0;
assign v3769ad7 = hbusreq0 & v3a63abb | !hbusreq0 & !v37439ad;
assign v3a707cd = hbusreq3_p & v3a5891c | !hbusreq3_p & v376ef42;
assign v3a64ded = hgrant4_p & v377d01e | !hgrant4_p & v372f62a;
assign v3a6157d = hbusreq0 & v3744501 | !hbusreq0 & v8455ab;
assign v3735b3d = hbusreq8 & v3774e2b | !hbusreq8 & v3a6fddb;
assign v3a6f646 = locked_p & v8455ab | !locked_p & v373c3bd;
assign v3a6dfb2 = hbusreq1_p & v3807bf8 | !hbusreq1_p & v3a66110;
assign v3765ce2 = hlock3 & v3731afc | !hlock3 & v3a6fbfc;
assign v3749bba = hbusreq4 & v3765627 | !hbusreq4 & v377a376;
assign v375a842 = hgrant1_p & v3a71452 | !hgrant1_p & v3806507;
assign v37240a4 = hmaster2_p & v3a6ab5f | !hmaster2_p & v373dfff;
assign v374a7ab = hgrant6_p & v3768633 | !hgrant6_p & v3a66ef6;
assign v376978a = jx0_p & v3a6be15 | !jx0_p & v3a6c2b2;
assign v3a579a3 = hbusreq6_p & v374fcd2 | !hbusreq6_p & !v8455ab;
assign v37275f8 = hmaster3_p & v8455ab | !hmaster3_p & v37258d0;
assign v3769b75 = hmaster0_p & v3a6dfb2 | !hmaster0_p & !v37500e0;
assign v3a5d474 = jx0_p & v375b776 | !jx0_p & v3a67fee;
assign v1e37cc1 = hmaster2_p & v3763209 | !hmaster2_p & v373d4ff;
assign v3a6fa63 = hmaster1_p & v374502e | !hmaster1_p & v373e41c;
assign v3a57445 = hlock1_p & v8455e7 | !hlock1_p & !v8455ab;
assign v372c49f = jx0_p & c587b2 | !jx0_p & v3a57e01;
assign v3a70f0c = hlock5 & v3a6c4c3 | !hlock5 & v3758bc2;
assign v376a619 = hbusreq5 & v37752be | !hbusreq5 & v8455ab;
assign v376747e = hmaster0_p & v3a635ea | !hmaster0_p & v377086b;
assign v3779183 = hgrant4_p & v3807f45 | !hgrant4_p & v3a5c80e;
assign v373221a = hmaster2_p & v377d9aa | !hmaster2_p & !v3744f62;
assign v88b8eb = hmaster1_p & v3724bf3 | !hmaster1_p & v3a298b6;
assign v3a66bfa = hmaster1_p & v3a635ea | !hmaster1_p & v377451f;
assign v3723cc2 = hbusreq0_p & v373c755 | !hbusreq0_p & v37674c1;
assign v37567f5 = hmaster0_p & v3a700b2 | !hmaster0_p & v3744b55;
assign v377e825 = hgrant4_p & v8455ab | !hgrant4_p & v3737909;
assign v3a5872a = hbusreq3_p & v3734a79 | !hbusreq3_p & v3a59d40;
assign v373c628 = hgrant2_p & v8455ab | !hgrant2_p & v37767d8;
assign v3731e55 = hmaster1_p & v3771076 | !hmaster1_p & v374c9e4;
assign v376d0d8 = hbusreq7 & v3a6376d | !hbusreq7 & v8455ab;
assign v3747d37 = hgrant4_p & v3750d06 | !hgrant4_p & v376b99f;
assign v373ac08 = hmaster2_p & v3747302 | !hmaster2_p & v3756304;
assign v377e56f = hbusreq6 & v376dcd0 | !hbusreq6 & !v3a69248;
assign v3748299 = hlock7 & v3a66274 | !hlock7 & v3a6f791;
assign v3a6f816 = hbusreq8_p & v3740e8d | !hbusreq8_p & v3a6ef64;
assign v3a611cf = hbusreq5_p & v37485df | !hbusreq5_p & v8455ab;
assign v377dac2 = hbusreq8_p & v376f516 | !hbusreq8_p & v375bbe2;
assign v3752ec0 = hgrant0_p & v37773a9 | !hgrant0_p & !v8455ab;
assign v375a4a0 = hbusreq5_p & v3771204 | !hbusreq5_p & v8455ab;
assign v37738e9 = hbusreq8_p & v3728876 | !hbusreq8_p & v3731780;
assign v3a63597 = hgrant3_p & v3754227 | !hgrant3_p & !v8455ab;
assign v3728419 = hmaster0_p & v37667c6 | !hmaster0_p & v3745b9c;
assign v3a6fdee = hmaster0_p & v3a6a312 | !hmaster0_p & v3a296d8;
assign v3808dca = hgrant6_p & v3a6f18f | !hgrant6_p & v3767e15;
assign v3745cea = hbusreq6_p & v3731a3b | !hbusreq6_p & v391331d;
assign beb41d = hmaster0_p & v372c221 | !hmaster0_p & v3a6f901;
assign v3a5a3be = hbusreq3 & v3a6f757 | !hbusreq3 & v377857d;
assign v373498b = hlock6_p & v373e10c | !hlock6_p & v3762949;
assign v3a5c75c = hbusreq5_p & v374193d | !hbusreq5_p & v3a61cb0;
assign v373a9c4 = hbusreq5 & v3a61a75 | !hbusreq5 & v3a66170;
assign v3744af9 = hmaster2_p & v372935c | !hmaster2_p & !v3a6b0c7;
assign v3746ce0 = hmaster2_p & v37283f8 | !hmaster2_p & v3779eea;
assign v377624b = hmaster2_p & v3758a4b | !hmaster2_p & v376c99e;
assign v3756cee = hbusreq2_p & v373913e | !hbusreq2_p & v8455ab;
assign v3760854 = hgrant6_p & v377f09a | !hgrant6_p & v3779582;
assign v3776c9a = hgrant0_p & v3a5b71a | !hgrant0_p & !v3750f2a;
assign v377e51b = hmaster2_p & v3a6f3a3 | !hmaster2_p & v3a70212;
assign v3775eee = hgrant4_p & v37606b8 | !hgrant4_p & v3761cdb;
assign v3767e71 = hmaster2_p & v3a5f1d4 | !hmaster2_p & v374bd09;
assign v37255a2 = hmaster1_p & v3a6fe0d | !hmaster1_p & v3a6e127;
assign v3754b2c = hlock6 & v375b980 | !hlock6 & v372e9f3;
assign v3258dd9 = hmaster0_p & v374ab22 | !hmaster0_p & v3a70267;
assign v3a557b1 = hbusreq2 & v373997b | !hbusreq2 & v35b774b;
assign v3a5e9a8 = hmaster2_p & v20d166d | !hmaster2_p & v37484de;
assign v3a70db0 = hmaster2_p & v3746c51 | !hmaster2_p & v3777311;
assign v3a5fd2f = jx0_p & v375ca80 | !jx0_p & v377ce91;
assign v3763f20 = hmaster2_p & v3723fcc | !hmaster2_p & v3a6f4c7;
assign v3a6f875 = hmaster0_p & v373dad7 | !hmaster0_p & !v3a705ec;
assign v3a6ff62 = jx1_p & v372b313 | !jx1_p & v37275f8;
assign v3a57ebf = hmaster0_p & v375c791 | !hmaster0_p & v375a4ea;
assign v3a6a7cb = hlock5_p & v89b450 | !hlock5_p & v3a6f423;
assign v37728dc = hmaster2_p & v375ac50 | !hmaster2_p & v38090ee;
assign v3747358 = hbusreq4_p & v3a71077 | !hbusreq4_p & !v3a60340;
assign v377597f = hgrant4_p & v376462a | !hgrant4_p & v3740df7;
assign v3a6cb16 = hbusreq6_p & v3734967 | !hbusreq6_p & !v374729b;
assign v3771913 = hgrant6_p & v8455ab | !hgrant6_p & v3a661b5;
assign v3a687be = hbusreq2_p & v377a393 | !hbusreq2_p & v8455ab;
assign v3731142 = hgrant4_p & v377b6ce | !hgrant4_p & v3759a00;
assign v374891f = hmaster1_p & v37386f5 | !hmaster1_p & v37440af;
assign v3760c3c = hbusreq2_p & v3750ebc | !hbusreq2_p & !v8455ab;
assign b69f28 = jx1_p & cc9e54 | !jx1_p & v373d203;
assign v3735153 = hgrant4_p & v372b77b | !hgrant4_p & v3a6b572;
assign v374f2d1 = hgrant7_p & v8455ce | !hgrant7_p & v3735e18;
assign v3778595 = hmaster1_p & v3a574bf | !hmaster1_p & v3a5da31;
assign v3754488 = hlock5_p & v3a7037a | !hlock5_p & v8455ab;
assign v3a69063 = hlock7_p & v3a65096 | !hlock7_p & v372e479;
assign v373f9eb = hgrant5_p & v373edb9 | !hgrant5_p & v377de56;
assign v373a0f8 = hlock7 & v377034f | !hlock7 & v375caa2;
assign v373f392 = hmastlock_p & v37386f2 | !hmastlock_p & v8455ab;
assign v376f37e = hbusreq7 & v3a5bbaa | !hbusreq7 & v373b837;
assign v3a7119c = hgrant4_p & v8455c1 | !hgrant4_p & v37703a5;
assign v373b887 = hbusreq5_p & v377d1dc | !hbusreq5_p & v373b02e;
assign v3727986 = hbusreq4_p & v376a39c | !hbusreq4_p & v37290a1;
assign v3a70dc0 = hgrant0_p & v8455ab | !hgrant0_p & v377217c;
assign v3738e72 = hbusreq4 & v372c3df | !hbusreq4 & !v373c8d0;
assign v3776859 = hgrant5_p & v3a70de3 | !hgrant5_p & v375a33d;
assign v372a02b = hmaster0_p & v37261b3 | !hmaster0_p & v8455e7;
assign v3724f5d = hbusreq4 & v3a6910c | !hbusreq4 & v8455ab;
assign v3a6fd87 = hmaster1_p & v98bccb | !hmaster1_p & b9675e;
assign v3a557d2 = hmaster1_p & v374dbf7 | !hmaster1_p & v3a5d3f6;
assign v376e316 = hgrant3_p & v3735809 | !hgrant3_p & v37389db;
assign v23fdab8 = locked_p & v376beee | !locked_p & v8455ab;
assign v35b7033 = hbusreq7 & v373edf3 | !hbusreq7 & v373abcf;
assign v3a7165d = hbusreq0 & v37578b4 | !hbusreq0 & v375c674;
assign v377c214 = hgrant6_p & v8455ab | !hgrant6_p & v3a70414;
assign v3a6355c = hbusreq5 & v3a6f07f | !hbusreq5 & v3723add;
assign v3a6fe04 = hgrant5_p & v3739dfa | !hgrant5_p & v3762dd5;
assign v375cd8c = hbusreq5 & v373755a | !hbusreq5 & v38076cf;
assign v372d42d = hmaster2_p & v3750b71 | !hmaster2_p & v374f329;
assign v373dfb4 = hbusreq0 & v37620eb | !hbusreq0 & v3748797;
assign v3756723 = hbusreq7_p & v3748da1 | !hbusreq7_p & v3761916;
assign v3a704ef = hmaster1_p & v37302a2 | !hmaster1_p & v35b6c3a;
assign v3738d68 = hgrant3_p & v3722e5c | !hgrant3_p & v9d7b97;
assign v3731a95 = hmaster1_p & v3766986 | !hmaster1_p & v3a71656;
assign v373ebac = hmaster0_p & v375d337 | !hmaster0_p & v3767e66;
assign v1e37938 = jx0_p & v373bce1 | !jx0_p & v376fdfb;
assign v3a70020 = hbusreq3 & v3741216 | !hbusreq3 & v8455ab;
assign v3a6fc64 = hbusreq3 & v37481f3 | !hbusreq3 & v3749b84;
assign v3763a84 = hbusreq6 & v3732cb4 | !hbusreq6 & v8455ab;
assign v377b330 = hbusreq0 & v3753f0d | !hbusreq0 & v3809a58;
assign v374bf8a = hbusreq2_p & v374df0b | !hbusreq2_p & v373e654;
assign v377a121 = hbusreq2_p & v373b5f5 | !hbusreq2_p & v8455ab;
assign v3740e49 = hbusreq3 & v3a67927 | !hbusreq3 & v38079ff;
assign v3731724 = hgrant4_p & v8455ab | !hgrant4_p & v3755167;
assign v3763e30 = hbusreq5 & v3a66aa6 | !hbusreq5 & v3a6e7ed;
assign v3a7107f = hmaster0_p & v3728c14 | !hmaster0_p & v373026e;
assign v37c0158 = hlock0 & v3a641d5 | !hlock0 & v3a5899d;
assign v3741b28 = hbusreq6_p & v3734b35 | !hbusreq6_p & v3a554a6;
assign v373e5a7 = hbusreq0 & v3a6fee1 | !hbusreq0 & v373d9d3;
assign v3a533d3 = hbusreq6 & v3a6f8f5 | !hbusreq6 & v8455bf;
assign v377a002 = hgrant4_p & v3764552 | !hgrant4_p & v3a61e9a;
assign v375041a = hbusreq8_p & v3a709d6 | !hbusreq8_p & v8455ab;
assign v37272ed = hbusreq6 & v3a6f586 | !hbusreq6 & !v3a6f3cf;
assign v375b4d8 = hbusreq4 & v374e542 | !hbusreq4 & !v8455ca;
assign b20520 = hmaster2_p & v3a70fd5 | !hmaster2_p & !v3723da9;
assign v3735ff7 = hmaster2_p & v3740f5d | !hmaster2_p & v3777c59;
assign v3a6cacb = hgrant0_p & v8455ab | !hgrant0_p & !v3a655cb;
assign v38099c8 = hbusreq2_p & v376f56d | !hbusreq2_p & !v8455ab;
assign v373325f = hbusreq6 & v3a58353 | !hbusreq6 & !v8455ab;
assign v37bfff7 = decide_p & v376b962 | !decide_p & v3a70d4a;
assign v3a634db = hbusreq4 & v3a70468 | !hbusreq4 & v376e4a6;
assign v3757a61 = hbusreq8_p & v3a70578 | !hbusreq8_p & v3a71032;
assign v3a53f1a = stateG10_1_p & v39ebac7 | !stateG10_1_p & v374089e;
assign v3768adf = hmaster3_p & v8455ab | !hmaster3_p & v375b752;
assign v376f178 = hbusreq0_p & v2aca784 | !hbusreq0_p & v8455ab;
assign v372adb6 = hmaster2_p & v3a701a1 | !hmaster2_p & v3744835;
assign v37422d8 = hbusreq1 & v37457fb | !hbusreq1 & v8455e7;
assign v3a6419e = hbusreq2_p & v3748f87 | !hbusreq2_p & !v8455ab;
assign v37269b2 = hbusreq5_p & v3764f06 | !hbusreq5_p & v3772c9f;
assign v3a636d2 = hbusreq7_p & v3a592bc | !hbusreq7_p & v3a65ea7;
assign v3a70424 = jx0_p & v3778a55 | !jx0_p & v8455ab;
assign v3749e33 = hgrant0_p & v3a71387 | !hgrant0_p & v8455ab;
assign v3756ebb = hgrant3_p & v3a55d41 | !hgrant3_p & v3a6eb86;
assign v373859f = hmaster0_p & v3a58287 | !hmaster0_p & v3808e2e;
assign v376ea13 = hmaster0_p & v3752e42 | !hmaster0_p & !v376ff85;
assign v372df82 = hgrant4_p & v375c7b9 | !hgrant4_p & !v3379070;
assign v374c4c0 = jx1_p & v3a6f8c5 | !jx1_p & v3a67a78;
assign v375dab1 = hlock0_p & v3a68c1f | !hlock0_p & !v3807bf8;
assign v373ad3f = hmaster2_p & v3a70a32 | !hmaster2_p & v3a6eb3f;
assign v374ef66 = hbusreq3_p & v3a6dc32 | !hbusreq3_p & v3739417;
assign v37640e9 = hgrant4_p & v37245f8 | !hgrant4_p & v375ba37;
assign v377d497 = hmaster1_p & v3a70592 | !hmaster1_p & v37420de;
assign v3a71175 = hlock5 & v3729597 | !hlock5 & v3a689e5;
assign v373f52e = hbusreq4 & v3a713cc | !hbusreq4 & v3a71554;
assign v3748d3e = hbusreq2 & v3778993 | !hbusreq2 & v8455ab;
assign v3a6e2d0 = hbusreq4_p & v3727c1d | !hbusreq4_p & !v3a573cc;
assign v3a5a868 = hmaster2_p & v372ee9a | !hmaster2_p & !v37564e4;
assign v373472c = hlock6_p & v3a57309 | !hlock6_p & !v8455ab;
assign v3a62ed6 = hgrant0_p & v3a65596 | !hgrant0_p & v3a70c61;
assign v37553b9 = hmaster0_p & v373df82 | !hmaster0_p & v374eaf4;
assign v3773940 = hlock8_p & v373bb3a | !hlock8_p & v3a6aa15;
assign v3a64a9a = hmaster2_p & v3a6f442 | !hmaster2_p & v3a55419;
assign v3724f05 = hmaster1_p & v3a635ea | !hmaster1_p & v3a5ba93;
assign v377c3ea = hgrant2_p & v8455e7 | !hgrant2_p & !v3a70974;
assign v377f24b = hlock5_p & v3765af5 | !hlock5_p & !v8455ab;
assign v377fc45 = hmaster0_p & v3725673 | !hmaster0_p & v3764a7d;
assign v373d9e0 = hgrant4_p & v3733da4 | !hgrant4_p & v373506a;
assign v3a70ac4 = hmaster0_p & v8455ab | !hmaster0_p & !v37590fb;
assign v376f30a = hlock0_p & v376a8cf | !hlock0_p & v3771b20;
assign v374757c = hmaster1_p & v377234d | !hmaster1_p & v3a6fdb6;
assign v37677b4 = hmaster0_p & v37730b9 | !hmaster0_p & v3a713a7;
assign v375e657 = hbusreq1_p & a5679d | !hbusreq1_p & v8455ab;
assign v374e0e9 = hmaster2_p & v3a6908b | !hmaster2_p & v375fc0a;
assign v376a129 = hmaster3_p & v375e23b | !hmaster3_p & v8455ab;
assign v37679b0 = hgrant5_p & v373f909 | !hgrant5_p & v3752759;
assign v3755d64 = hbusreq2 & v376b21a | !hbusreq2 & v8455ab;
assign v3726f38 = hbusreq0 & v3748347 | !hbusreq0 & v377389f;
assign v3a6fac5 = hlock3_p & v2092eac | !hlock3_p & v37720e5;
assign v3761bb7 = hlock0 & v3748797 | !hlock0 & v3a6f9e5;
assign v373e6bc = hlock5_p & v3a56cfd | !hlock5_p & v3a6fabf;
assign v3732586 = hbusreq7_p & v3762363 | !hbusreq7_p & v3809e25;
assign v1e3780e = hmaster2_p & v3753dab | !hmaster2_p & v3a6fa39;
assign v2ff8f8e = hbusreq6_p & v3a70f78 | !hbusreq6_p & v3737280;
assign v372456c = hgrant6_p & d2e9f6 | !hgrant6_p & v37368b3;
assign v3763db6 = hmaster0_p & v37793e4 | !hmaster0_p & v3774deb;
assign v374686d = hgrant4_p & v373b687 | !hgrant4_p & v3753dd4;
assign v3a70055 = hgrant2_p & v8455ab | !hgrant2_p & v376b5bc;
assign v3a605bd = hgrant3_p & v8455be | !hgrant3_p & !v372d6e5;
assign v37551f2 = hgrant1_p & v3748797 | !hgrant1_p & v8455ab;
assign v37528b0 = hbusreq0_p & v3809adf | !hbusreq0_p & v39a537f;
assign v3a70956 = hbusreq7 & v3a54e47 | !hbusreq7 & v8455ab;
assign v375a804 = hmaster0_p & v3a6ce52 | !hmaster0_p & !v377ba8a;
assign v3a5cbd8 = hbusreq6_p & v8455ab | !hbusreq6_p & v374e26d;
assign v3735302 = hbusreq5 & v3a57e27 | !hbusreq5 & !v372b971;
assign v3752556 = hlock0 & v3a5e2e1 | !hlock0 & v37346dc;
assign v375783c = hlock2_p & v3750aea | !hlock2_p & v375361a;
assign v3778cdd = hgrant3_p & v8455ab | !hgrant3_p & v372b5b0;
assign a81487 = hmastlock_p & v3744037 | !hmastlock_p & v8455ab;
assign v3a6fde0 = hmaster2_p & v8455ab | !hmaster2_p & v3748797;
assign v3a6da6b = hbusreq4_p & v3726d1f | !hbusreq4_p & v38073c9;
assign v3729f14 = hbusreq2_p & v373d99d | !hbusreq2_p & v8455ab;
assign v37576ec = hmaster3_p & v372d780 | !hmaster3_p & !v3759d9c;
assign v375859f = hgrant2_p & v2619ada | !hgrant2_p & v8455ab;
assign v3764818 = hmaster0_p & v3a652c7 | !hmaster0_p & !v377fbbf;
assign v375581b = hgrant6_p & v3a6c97d | !hgrant6_p & v3757e4b;
assign v3a66ff2 = hgrant0_p & v37301f5 | !hgrant0_p & v37772bf;
assign v375dda4 = hmaster0_p & v3730288 | !hmaster0_p & v8455ab;
assign b95629 = hlock4 & v3a5dd62 | !hlock4 & v3a59264;
assign v3a5740f = hmaster1_p & v94faa4 | !hmaster1_p & v372dfba;
assign v3a60feb = hmaster0_p & v3755136 | !hmaster0_p & v37268cc;
assign v377d126 = stateA1_p & v37295fe | !stateA1_p & !a81487;
assign v377bb6d = hgrant4_p & v3a6eb39 | !hgrant4_p & v9ec00e;
assign v374a189 = hbusreq7 & v3a710ea | !hbusreq7 & v3a69b91;
assign v37351bc = hbusreq1 & v374362e | !hbusreq1 & v8455ab;
assign v3734f09 = hgrant3_p & v377f342 | !hgrant3_p & !v37293b1;
assign v376a556 = hmaster1_p & v37524b4 | !hmaster1_p & v3a6274c;
assign v372ade8 = hbusreq1_p & v377d408 | !hbusreq1_p & !v8455ab;
assign v3a5a52f = jx0_p & v3a656f0 | !jx0_p & v3775120;
assign v2093059 = hbusreq3 & v8455ab | !hbusreq3 & !v373ad95;
assign c8d28b = hbusreq0 & v3a6f328 | !hbusreq0 & v3731389;
assign v375e039 = hmaster0_p & v3a619c0 | !hmaster0_p & !c60fa0;
assign v3a62c37 = hlock8_p & v3a70618 | !hlock8_p & v3a57f64;
assign v375ff74 = hlock6_p & v3753f1a | !hlock6_p & v376430b;
assign v372fbf4 = hlock3_p & v3a7031d | !hlock3_p & v377a6ce;
assign v37603b3 = hbusreq6 & v37356f0 | !hbusreq6 & v8455ab;
assign v3a5cb5f = hbusreq6_p & v377757b | !hbusreq6_p & v3a70408;
assign v3746202 = hbusreq0 & v3a63884 | !hbusreq0 & v376d86d;
assign v3a6fc70 = hmaster0_p & v3a5c6d0 | !hmaster0_p & v3a70941;
assign v37680af = hgrant6_p & v3735d71 | !hgrant6_p & v377b2ce;
assign v3a6c02f = hbusreq6 & v3a583ee | !hbusreq6 & v3767429;
assign v37705f3 = hmaster2_p & v3a5fc34 | !hmaster2_p & v374693f;
assign v31c3694 = hbusreq2_p & v3779060 | !hbusreq2_p & !v3a6dfb2;
assign v3a68e41 = jx3_p & v3751fde | !jx3_p & v3a585f5;
assign v3759586 = hmaster2_p & v3767e7e | !hmaster2_p & v3a5690e;
assign v3a6f9be = hbusreq8_p & v3a70e7a | !hbusreq8_p & v374ab4c;
assign v377bb62 = hgrant3_p & v35b774b | !hgrant3_p & v3776fe2;
assign v3a6d3b6 = hmaster1_p & v8db8b7 | !hmaster1_p & v374f1e9;
assign v377273d = hbusreq5 & v3a70866 | !hbusreq5 & v376c335;
assign v3a6fffd = hbusreq4_p & v3741cfb | !hbusreq4_p & v3748797;
assign v377389f = hgrant6_p & v377e1d0 | !hgrant6_p & v3775fae;
assign v3a6ec1b = hgrant7_p & v3a59c0b | !hgrant7_p & v3a6f6dd;
assign v3a5cf84 = jx0_p & v3a5d704 | !jx0_p & v37702e8;
assign v37383bb = hmaster3_p & v37288c3 | !hmaster3_p & v376da8d;
assign v377ddc1 = hbusreq4_p & v3727c1d | !hbusreq4_p & !v3a706af;
assign v3a5f83c = hbusreq4 & v3763d77 | !hbusreq4 & v376e90a;
assign v377e36c = hbusreq5 & v375fe02 | !hbusreq5 & aeff0f;
assign v3729421 = hbusreq3_p & v3750978 | !hbusreq3_p & !v8455ab;
assign v3a65a24 = hbusreq0_p & v35772a5 | !hbusreq0_p & !v3776ce0;
assign v3a71130 = hbusreq0_p & v3a5cfdb | !hbusreq0_p & v3774e64;
assign v8455c6 = hbusreq5 & v8455ab | !hbusreq5 & !v8455ab;
assign v3748f81 = hmaster2_p & v3a7112c | !hmaster2_p & v3742cd4;
assign v377fa89 = hbusreq2_p & v374d13c | !hbusreq2_p & v3a713e3;
assign v8dfd63 = hmaster0_p & v39a5380 | !hmaster0_p & v377b6b2;
assign v3a70eb6 = hlock3 & v37254c0 | !hlock3 & v3806507;
assign v3777d2e = hlock4_p & d99853 | !hlock4_p & !v8455ab;
assign v3758bcd = hlock8 & v376956a | !hlock8 & v3a5d8d3;
assign v3a6962d = hbusreq2 & v3a6f7bf | !hbusreq2 & v8455e7;
assign v3776865 = hmaster2_p & v3747302 | !hmaster2_p & v37786a6;
assign v3753328 = hmaster0_p & v8455ab | !hmaster0_p & !v372e3b4;
assign v3a67927 = hgrant0_p & v1e3791d | !hgrant0_p & v3a66460;
assign v3a68f22 = hmaster3_p & v3a7113d | !hmaster3_p & v3723025;
assign v37686af = hbusreq1 & v37270d9 | !hbusreq1 & v8455ab;
assign v3a6fd19 = hmaster0_p & v372bea3 | !hmaster0_p & !v373197c;
assign v3722be8 = hgrant1_p & v8455ab | !hgrant1_p & v8455b0;
assign v3a7127f = hgrant6_p & v377db8a | !hgrant6_p & v3a6fe6a;
assign v3a70e79 = hbusreq0 & v374fc57 | !hbusreq0 & v3a57750;
assign v377d15d = hbusreq7 & v3a5ab7b | !hbusreq7 & v3743a4c;
assign v39e9c98 = hmaster2_p & v3a635ea | !hmaster2_p & v376489b;
assign v373eba7 = hmaster2_p & adf78a | !hmaster2_p & v8455ab;
assign v3732b1e = hbusreq4 & v3a711ac | !hbusreq4 & v8455ab;
assign v3a55b16 = hmaster1_p & v3723211 | !hmaster1_p & v3a5520a;
assign v3769f23 = hbusreq5_p & v374871a | !hbusreq5_p & v374457a;
assign v3a6fc43 = hlock4_p & v126f91f | !hlock4_p & v3760f64;
assign v3741cda = hgrant2_p & v372d1a4 | !hgrant2_p & v3751196;
assign v2ff87a0 = hbusreq5_p & v3728fa6 | !hbusreq5_p & v3a54677;
assign v3a5b5ef = hgrant4_p & v8455ab | !hgrant4_p & v375bb15;
assign v377c94b = hbusreq4_p & v374df45 | !hbusreq4_p & v375fcb7;
assign v3722dd5 = hbusreq7_p & v8455ab | !hbusreq7_p & v373ad69;
assign v3a70c69 = hbusreq5 & v3742303 | !hbusreq5 & v3760bda;
assign v3a70700 = hmaster1_p & v8455c6 | !hmaster1_p & v374bc97;
assign v8455bd = hbusreq3_p & v8455ab | !hbusreq3_p & !v8455ab;
assign v375a637 = hbusreq4_p & v3a58b8f | !hbusreq4_p & v3757a57;
assign v37528b8 = hmaster3_p & v8455ab | !hmaster3_p & v3739769;
assign v374c28d = hmaster1_p & v2acaec4 | !hmaster1_p & v3735a87;
assign v376eb1d = hgrant4_p & v3a6f059 | !hgrant4_p & v8455ab;
assign v3763030 = hgrant4_p & v376ab5d | !hgrant4_p & v3a595b8;
assign v3a5f97f = hmaster0_p & v37651e0 | !hmaster0_p & !v937864;
assign v377c186 = hgrant1_p & v3a7069e | !hgrant1_p & !v3752a45;
assign v3747c3d = hbusreq0 & v3a65b53 | !hbusreq0 & v373e814;
assign v3a703df = hburst1 & v3757c6f | !hburst1 & v3775da7;
assign v372a4c4 = hbusreq2_p & v377636a | !hbusreq2_p & v3a58a16;
assign v37601a1 = hbusreq0 & v374afa4 | !hbusreq0 & !v376ce15;
assign v3a603cf = hbusreq6_p & v3a714e9 | !hbusreq6_p & v3a705ce;
assign c0b985 = hbusreq4_p & v3739594 | !hbusreq4_p & v8455ab;
assign v3749469 = hlock5 & v3763d53 | !hlock5 & v3a6826a;
assign v377c57a = hbusreq2_p & v376ac9b | !hbusreq2_p & !v8455ab;
assign v374ca2d = stateG2_p & v3a5a496 | !stateG2_p & !v372c42d;
assign v372f2fe = hbusreq5 & v373e6d2 | !hbusreq5 & v374f658;
assign v37360b3 = hgrant3_p & v3739018 | !hgrant3_p & v373b7c8;
assign v375a1fd = hmaster1_p & v8455ab | !hmaster1_p & v3726e48;
assign v37657e4 = hmaster2_p & v3a6be44 | !hmaster2_p & v8455bd;
assign v3a713f2 = hmaster2_p & v377b774 | !hmaster2_p & v8455ab;
assign v37682a8 = hbusreq1_p & v372865e | !hbusreq1_p & v372eb43;
assign v372a3cb = hlock6_p & v377de7b | !hlock6_p & v375d616;
assign v3759d08 = hbusreq4_p & v3754b79 | !hbusreq4_p & v3a70210;
assign v3a59b87 = hlock0_p & v376dbdf | !hlock0_p & v3a6e592;
assign v376374e = hbusreq7 & v374067b | !hbusreq7 & v376ae9f;
assign v373a7b4 = hbusreq8_p & v3a54120 | !hbusreq8_p & v3a5a2e5;
assign v3757231 = hlock7_p & v3a67c34 | !hlock7_p & v3a60e78;
assign v3741627 = hmaster0_p & v3a70902 | !hmaster0_p & v37549e2;
assign v3759e04 = hbusreq7 & v3a639a1 | !hbusreq7 & v372d5ba;
assign v3762fcb = hgrant2_p & v3722f85 | !hgrant2_p & v8455ab;
assign v375534a = hbusreq6 & v37642a0 | !hbusreq6 & v374a637;
assign v376a3f7 = hmaster0_p & v3768589 | !hmaster0_p & v374b24a;
assign v375de18 = locked_p & v3a6f958 | !locked_p & v39a537f;
assign v376b97b = hgrant1_p & cc9d04 | !hgrant1_p & v35772a6;
assign v3744161 = hgrant3_p & v37650dd | !hgrant3_p & !v3737ac8;
assign v3a61f82 = hgrant3_p & v8455ab | !hgrant3_p & v37773a2;
assign v374e650 = hbusreq7 & v3a70301 | !hbusreq7 & v3a60276;
assign v374b9e6 = hmaster0_p & v3a6f09b | !hmaster0_p & v377fbbf;
assign v3a6ff8a = hlock1 & v3762434 | !hlock1 & v3770f7a;
assign v3a6ebf1 = hlock0_p & v2acb5a2 | !hlock0_p & v8455ab;
assign v3a6efcd = hmaster2_p & v8455ab | !hmaster2_p & v8455bf;
assign v3739cda = hgrant6_p & v8455ab | !hgrant6_p & v3738762;
assign v35b9d58 = hmaster0_p & v375e9b2 | !hmaster0_p & v3747d30;
assign v372ad5a = jx0_p & v3a6202c | !jx0_p & v37348f8;
assign v372f7d4 = hbusreq3 & v377ba55 | !hbusreq3 & v8455ab;
assign v3770827 = hmaster0_p & v3a619c0 | !hmaster0_p & v372cb9d;
assign v37655d3 = hbusreq3_p & v3a668ec | !hbusreq3_p & v8455b0;
assign v9ae45c = hmaster2_p & v3a6dc08 | !hmaster2_p & v372b5f5;
assign v3a5caf4 = hmaster1_p & v1e38262 | !hmaster1_p & v377104a;
assign v3722f10 = hgrant6_p & v375d877 | !hgrant6_p & v3a58554;
assign v3739589 = hmaster0_p & v374a1f5 | !hmaster0_p & v372ba40;
assign v3736847 = hbusreq2_p & v376f9a8 | !hbusreq2_p & v376d856;
assign v3777b18 = hmaster1_p & v37302a2 | !hmaster1_p & v374bb64;
assign v3775b7e = hbusreq5_p & v3742649 | !hbusreq5_p & v3a61516;
assign v37581d2 = hgrant5_p & v3733c82 | !hgrant5_p & v376d57d;
assign v3a6f442 = hgrant4_p & v3727943 | !hgrant4_p & v3774b98;
assign v373eaf6 = hgrant4_p & v376faab | !hgrant4_p & v8455ab;
assign v3a68e5d = hlock4_p & v375c718 | !hlock4_p & v3a6fac6;
assign v376a8d5 = hready & v375eb9c | !hready & v37295fe;
assign v380749d = hgrant3_p & v8455ab | !hgrant3_p & v3758eae;
assign v374cbe2 = hmaster0_p & v8455ab | !hmaster0_p & v3a6f8ae;
assign cf4a8f = hbusreq0_p & v372dadb | !hbusreq0_p & v3a706c7;
assign v3a7051e = hlock7 & v39eaae4 | !hlock7 & v3774e7b;
assign v3778f46 = hmaster0_p & v373b30b | !hmaster0_p & v3768a78;
assign v3756996 = hmaster0_p & v3742c87 | !hmaster0_p & v23fd8c6;
assign v1e37ae9 = hbusreq7_p & v3726bdb | !hbusreq7_p & v3a63f43;
assign v377dfbd = hgrant5_p & v372a264 | !hgrant5_p & v374e684;
assign v3763f13 = hmaster0_p & v3a635ea | !hmaster0_p & v3a62245;
assign v37380be = hbusreq5 & v374e179 | !hbusreq5 & v374e784;
assign v37342ef = hmaster2_p & v8455b3 | !hmaster2_p & v374b3cf;
assign v377b253 = hmaster0_p & v3a6a089 | !hmaster0_p & v377d95a;
assign v3764fd5 = hmaster3_p & v37377f0 | !hmaster3_p & v3736cd2;
assign v374b256 = hbusreq2 & v3a66e70 | !hbusreq2 & v3a5f5bb;
assign v3806db0 = hgrant4_p & v8455ab | !hgrant4_p & v3732701;
assign v376d488 = hlock4_p & v3a54c77 | !hlock4_p & !v8455ab;
assign v37599a4 = hlock5_p & v377a104 | !hlock5_p & !v8455ab;
assign v3a6f9b9 = hgrant2_p & v8455ab | !hgrant2_p & v3725582;
assign v3a712ca = hmaster2_p & v3a635ea | !hmaster2_p & v37512ca;
assign v375fcfa = hbusreq5 & v3772464 | !hbusreq5 & v8455ab;
assign v37488d2 = jx0_p & v3763474 | !jx0_p & v3a6f645;
assign v3a56c66 = hbusreq1_p & v3a6767a | !hbusreq1_p & !v35772a6;
assign v3a63b90 = hgrant3_p & v3a55d41 | !hgrant3_p & v374a044;
assign v3a65b2b = hmaster0_p & v3779be2 | !hmaster0_p & v3a5ed4a;
assign v37416e1 = hbusreq0_p & v374ccb7 | !hbusreq0_p & v8455ab;
assign v3776b20 = hmaster2_p & v8455c2 | !hmaster2_p & v8455b2;
assign v3735ad0 = hbusreq7 & v37671d3 | !hbusreq7 & v3807969;
assign v3a71509 = hmaster0_p & v3a70641 | !hmaster0_p & v3a677ce;
assign v3a70408 = hbusreq6 & v377b8ee | !hbusreq6 & v8455ab;
assign v3a6eb8c = hmaster1_p & v376964a | !hmaster1_p & v37787dd;
assign v373414c = stateA1_p & v8455ab | !stateA1_p & !v3a6f682;
assign v37522bc = hbusreq3_p & v3a635ea | !hbusreq3_p & v3759f61;
assign v3a6f351 = stateG10_1_p & v3744a2f | !stateG10_1_p & v3a57e21;
assign v37437c1 = hmaster0_p & v374aae0 | !hmaster0_p & v376d07b;
assign v377d219 = stateA1_p & v8455ab | !stateA1_p & !v373fecd;
assign v3a54b84 = hmaster1_p & v3776f2c | !hmaster1_p & v3a2a41f;
assign v3762ba2 = hmaster2_p & v3a67577 | !hmaster2_p & !v8455ab;
assign v3749907 = hbusreq3_p & v3a5f8d0 | !hbusreq3_p & v3775303;
assign v3768062 = hbusreq1_p & v3a71452 | !hbusreq1_p & v3743b9e;
assign v3a709eb = hbusreq7_p & v3a704c4 | !hbusreq7_p & v3773076;
assign v3739334 = hbusreq6_p & v3748797 | !hbusreq6_p & v3a63dbf;
assign v3a6f117 = hbusreq5 & v376293f | !hbusreq5 & v3742cd4;
assign v37599eb = hmaster2_p & v374743d | !hmaster2_p & v372615f;
assign v3738c0a = hgrant4_p & v37479ef | !hgrant4_p & v3738ad8;
assign v377da10 = hlock5_p & v8455ab | !hlock5_p & v3735675;
assign v3a602d7 = hbusreq6_p & v3779544 | !hbusreq6_p & !v8455ab;
assign v373d091 = hbusreq5_p & v3775b3a | !hbusreq5_p & v8455ab;
assign v3a58546 = jx2_p & v372a0e6 | !jx2_p & v377b32c;
assign v3a716a0 = hbusreq4_p & v3a7088f | !hbusreq4_p & v8455ab;
assign v3734cb7 = hbusreq6_p & v377c07a | !hbusreq6_p & v3a67fd9;
assign v37562a5 = hgrant6_p & v8455ab | !hgrant6_p & v3a6fddd;
assign v374bdea = hmaster0_p & v3a71611 | !hmaster0_p & v374fe44;
assign v37596df = hbusreq5 & v377d6fc | !hbusreq5 & v373b9ab;
assign v376b71f = hbusreq8_p & v3a71193 | !hbusreq8_p & v372647c;
assign v377a6fe = hmaster0_p & v375808f | !hmaster0_p & v3a6ab5e;
assign v375f046 = hbusreq3 & v39a5265 | !hbusreq3 & !v2aca977;
assign v37402f0 = hbusreq3_p & v375d7b6 | !hbusreq3_p & v375825a;
assign v3738ea9 = hmaster0_p & v37391ac | !hmaster0_p & v374dad0;
assign v374ef62 = hmaster1_p & v37782c9 | !hmaster1_p & v3753cf6;
assign v373651a = hbusreq7 & v375c4ab | !hbusreq7 & v3a5a807;
assign v3724733 = hmaster0_p & v3a6f75d | !hmaster0_p & v8455ab;
assign v372a22f = hlock5_p & v3747a5b | !hlock5_p & v3a67c50;
assign v3a6f8de = hbusreq3_p & v3739021 | !hbusreq3_p & v8455ab;
assign v3769f01 = hmaster2_p & v374f319 | !hmaster2_p & v8455ab;
assign v3772d6e = hbusreq4_p & v3734aae | !hbusreq4_p & v8455b0;
assign v3769edd = hmaster0_p & v9af7ec | !hmaster0_p & v3777ac3;
assign v39eaae9 = hlock7 & v376769e | !hlock7 & v3763b4d;
assign v3779647 = hlock0_p & v3750d37 | !hlock0_p & !v8455ab;
assign v3773069 = hbusreq0_p & v3771728 | !hbusreq0_p & v3a6918e;
assign v375d40b = hlock2_p & v3770d6d | !hlock2_p & adf78a;
assign v37323c5 = hbusreq5 & v375c92f | !hbusreq5 & v374f9cc;
assign v3a5f26f = hbusreq0 & v374b5da | !hbusreq0 & v3763868;
assign v375cf36 = hlock0_p & v3a635ea | !hlock0_p & v37611b7;
assign v3769c51 = jx0_p & v3a67c9e | !jx0_p & v3a70287;
assign v377d077 = hmaster0_p & v3739ec9 | !hmaster0_p & v3a70574;
assign v3a6dded = hmaster2_p & v374d4e6 | !hmaster2_p & v3a7142f;
assign v372661f = hbusreq5_p & v3a6ff4b | !hbusreq5_p & !v3a7122f;
assign v3730038 = hmaster1_p & v374a9d0 | !hmaster1_p & v38067b3;
assign v3a5b774 = hgrant2_p & v8455ab | !hgrant2_p & v376071e;
assign v372b726 = hbusreq2 & v3806db7 | !hbusreq2 & v8455ab;
assign v3730e2a = hbusreq3_p & v35b774b | !hbusreq3_p & v9ed516;
assign v3765740 = hgrant4_p & v3756304 | !hgrant4_p & v3a710f3;
assign v376c85c = hmaster2_p & v3767e7e | !hmaster2_p & v3a6fc66;
assign v374e620 = hbusreq7_p & v3a6f2f8 | !hbusreq7_p & v3a704d2;
assign v377472b = hgrant4_p & v3a6b7e9 | !hgrant4_p & v37755d5;
assign v37360c0 = hbusreq5 & v377e869 | !hbusreq5 & !v3742b88;
assign v3a7154d = hmaster3_p & v2acafdd | !hmaster3_p & v376b1ee;
assign v3735a7c = hgrant6_p & v3758166 | !hgrant6_p & !v372a7ae;
assign v3730c86 = hbusreq5_p & v373e1fb | !hbusreq5_p & v37541c6;
assign v3a6b20a = hgrant6_p & v8455ab | !hgrant6_p & v37658f5;
assign v3a6f44a = hbusreq7 & v3747f46 | !hbusreq7 & !v373518a;
assign v372e754 = hmaster0_p & v376111d | !hmaster0_p & v376afb1;
assign ae5f9e = hmaster0_p & v372f2ce | !hmaster0_p & v374c164;
assign v375e516 = hbusreq7_p & v3a57fa1 | !hbusreq7_p & v3730f34;
assign v35b9d5e = hbusreq6_p & v373f883 | !hbusreq6_p & v373a2f2;
assign v3731720 = hmaster0_p & v3a5c0e1 | !hmaster0_p & v3774e4f;
assign v3749899 = hmaster0_p & v8455ab | !hmaster0_p & v375a5a1;
assign v39eb413 = hmaster0_p & v3a6eef7 | !hmaster0_p & v3a69606;
assign v3a6f376 = hbusreq7_p & v3737846 | !hbusreq7_p & v3731ea5;
assign v3726810 = hbusreq4_p & v3a71247 | !hbusreq4_p & v3765396;
assign v3a6ffae = busreq_p & v35772a6 | !busreq_p & v3577306;
assign v376d8c1 = hbusreq6 & v3a57f8b | !hbusreq6 & v3a58102;
assign v3777e0e = hlock0 & v3a620d3 | !hlock0 & v37513bc;
assign v3a6a68c = hbusreq5_p & v2acb110 | !hbusreq5_p & v3a6fb77;
assign v377868e = hlock6 & v3a5c015 | !hlock6 & v3778e03;
assign v3737ac6 = hgrant0_p & v8455ab | !hgrant0_p & v3a6d0ef;
assign v3773acc = hmaster0_p & v1e382e7 | !hmaster0_p & !v373d593;
assign v3733ee4 = hmaster1_p & v3a633bf | !hmaster1_p & v373a973;
assign v37474d6 = hmaster0_p & v3a712a2 | !hmaster0_p & !v3a583b0;
assign v3772a27 = hbusreq7 & v39ea259 | !hbusreq7 & v376775d;
assign v37288db = hgrant2_p & v377fc87 | !hgrant2_p & v3737e8c;
assign v3738de9 = hlock0_p & v37397c3 | !hlock0_p & v3a70295;
assign v3758abd = hmaster0_p & beaea1 | !hmaster0_p & v3a7090f;
assign v23fe21d = hbusreq7 & v372b034 | !hbusreq7 & v3a6f52a;
assign v376efda = hgrant3_p & v35b7299 | !hgrant3_p & v377e5fd;
assign v3a6165e = hbusreq8 & v1e37acb | !hbusreq8 & v373c404;
assign v3739bb2 = hbusreq2 & v3a64ee3 | !hbusreq2 & !v3a70131;
assign v3a71125 = jx0_p & v3761da5 | !jx0_p & v8455ab;
assign v3a6e105 = hbusreq6 & v37686f6 | !hbusreq6 & v376711c;
assign v3a5cf3c = hbusreq5_p & v3a6f5cd | !hbusreq5_p & !v3809892;
assign v375e439 = hbusreq7 & v3761d84 | !hbusreq7 & v376e66e;
assign v374057a = stateA1_p & v8455ab | !stateA1_p & v376147f;
assign v98068b = hmaster0_p & v37608ba | !hmaster0_p & v8455ab;
assign v3a67e13 = hmaster0_p & v3728d9c | !hmaster0_p & v3a70375;
assign v3733ac0 = hbusreq8_p & v3a6efb1 | !hbusreq8_p & v373f0c7;
assign v377d595 = hmaster0_p & v3775e03 | !hmaster0_p & v373ac71;
assign v3a708ff = hgrant8_p & v8455ab | !hgrant8_p & !v3775379;
assign v3a6963f = hlock2_p & v3764af7 | !hlock2_p & !v374e459;
assign v372367c = hgrant6_p & v3a68fc9 | !hgrant6_p & v373d338;
assign v3a708f8 = hbusreq7_p & v375dd84 | !hbusreq7_p & v3a70831;
assign v3769325 = hmaster0_p & v3a66d3e | !hmaster0_p & v8455ab;
assign v3a5b1ec = hbusreq4_p & v3a635ea | !hbusreq4_p & v374523b;
assign v3a712a7 = hmaster1_p & v3768a1c | !hmaster1_p & v3a54b77;
assign v3a709d2 = hlock0 & v3a67cff | !hlock0 & v373a90e;
assign v375323b = hbusreq1_p & v373ead4 | !hbusreq1_p & v3760bb4;
assign v373cc95 = hbusreq6_p & v375e657 | !hbusreq6_p & !v3a69591;
assign v3809b53 = hbusreq7_p & v3a6c0b7 | !hbusreq7_p & v3a700d3;
assign v372d2ad = hbusreq2_p & v39a5381 | !hbusreq2_p & v9181c9;
assign v3a66ba8 = hbusreq8 & v373e712 | !hbusreq8 & v372e550;
assign v3a70a4d = hbusreq4 & v3a70d04 | !hbusreq4 & v3a539bb;
assign v9f9402 = hbusreq6 & v3744380 | !hbusreq6 & v373a772;
assign v3a6a036 = hbusreq4 & v8455ab | !hbusreq4 & !v8455c3;
assign a21c18 = hgrant0_p & v3733d6e | !hgrant0_p & v375da3a;
assign v374b6ac = hlock0 & v3762502 | !hlock0 & v3a57ac7;
assign v3a6fab9 = hlock4 & v3a70a4f | !hlock4 & v374ffb7;
assign v3a702c2 = hlock6_p & v8455b0 | !hlock6_p & !v8455ab;
assign v3a6eecb = hmaster0_p & v375d1a1 | !hmaster0_p & v3a708a7;
assign v37656b8 = hbusreq0 & v380719b | !hbusreq0 & v377222a;
assign v3a67447 = hmaster2_p & v373cd16 | !hmaster2_p & v377961f;
assign v2acb0d7 = hmaster1_p & v8455c3 | !hmaster1_p & v373f349;
assign v3a64987 = hmaster2_p & v8455ab | !hmaster2_p & v3760353;
assign v377f118 = hgrant2_p & v3779b95 | !hgrant2_p & !v8455ab;
assign v3a5a985 = hbusreq3 & v373b0a4 | !hbusreq3 & v3a6fdef;
assign v3762d09 = hmaster2_p & v3a635ea | !hmaster2_p & v3754df4;
assign v99b721 = hmaster1_p & v3751dd2 | !hmaster1_p & v3a6e844;
assign v3a6f6c7 = hmaster0_p & v3779183 | !hmaster0_p & v3a60358;
assign v3a6ef1f = hgrant3_p & v3a69487 | !hgrant3_p & v3736fdd;
assign v3a6fa39 = hbusreq1_p & v8455b0 | !hbusreq1_p & v3753dab;
assign v3775630 = hgrant7_p & v3a6eb5b | !hgrant7_p & v3a6f69c;
assign v3743165 = hbusreq5 & v3a707ec | !hbusreq5 & v37404d0;
assign v3766a98 = hlock2 & v37524a6 | !hlock2 & v3a6440f;
assign v37777bf = hlock0_p & v372dadb | !hlock0_p & bc9e23;
assign v3a5f33d = hlock5 & v975066 | !hlock5 & v372d643;
assign v377d042 = hlock0 & v375da82 | !hlock0 & v3778a76;
assign v3a7112a = hbusreq4_p & v37647ce | !hbusreq4_p & v374eaeb;
assign v3a61e59 = hbusreq6_p & v3a6f39b | !hbusreq6_p & !v3727976;
assign v3a70f33 = hmaster0_p & v3a57584 | !hmaster0_p & v3728fd0;
assign v3a6fb44 = hbusreq7_p & v372f3fc | !hbusreq7_p & v8455ab;
assign v374bc77 = hgrant0_p & v37719b4 | !hgrant0_p & v8455ab;
assign v3a6eafc = stateG10_1_p & v3778ed4 | !stateG10_1_p & !v3a6e66e;
assign v37233e7 = hbusreq6 & v375da9c | !hbusreq6 & v37450b8;
assign v3759279 = hmaster2_p & v2acafcc | !hmaster2_p & v374aa71;
assign v3a70550 = hbusreq5_p & v3a6f73c | !hbusreq5_p & v8455ab;
assign v3763f30 = hmaster0_p & v3a6fe0d | !hmaster0_p & v3a6f692;
assign v3758bbf = hmaster1_p & v373ad69 | !hmaster1_p & v376e77e;
assign v3774b16 = hmaster0_p & v3a6b60d | !hmaster0_p & v3761c72;
assign v3730829 = hmaster2_p & v376b4e1 | !hmaster2_p & !v37388ce;
assign v3737dc7 = hbusreq5 & v3a62c46 | !hbusreq5 & !v3766216;
assign v8637a5 = hmaster2_p & v377e9bb | !hmaster2_p & v8455ab;
assign v3a7006e = hmaster1_p & v3733d60 | !hmaster1_p & v38064e3;
assign v3741afa = hgrant6_p & v8455ab | !hgrant6_p & v374a3f3;
assign v37500d0 = jx1_p & v3a70207 | !jx1_p & v37477d5;
assign v3757ce3 = hmaster2_p & v3762870 | !hmaster2_p & v373698e;
assign v37665bf = locked_p & v8455ab | !locked_p & v3a6a939;
assign v3a5d8d3 = hlock7 & v3a68916 | !hlock7 & v3728455;
assign v376b856 = hmaster2_p & v3a6e5f0 | !hmaster2_p & v8455b0;
assign v372549f = hmaster0_p & v376e0cd | !hmaster0_p & v3a57e58;
assign v37333a4 = hmaster2_p & v3a6ff25 | !hmaster2_p & v3732dac;
assign v374e4bd = hmaster1_p & v3a5fe3c | !hmaster1_p & v374f979;
assign v3751860 = start_p & v3730a0f | !start_p & v3a70ce3;
assign v86d306 = hbusreq6_p & v3743ada | !hbusreq6_p & v373619d;
assign v37307d4 = hbusreq4_p & v3a706f1 | !hbusreq4_p & v374b9ee;
assign v375d689 = hlock3 & v3a5cd50 | !hlock3 & v3a59d9d;
assign v372952e = hlock6 & v3a68f4f | !hlock6 & v3a710a2;
assign v3a71579 = hmaster2_p & v8455ab | !hmaster2_p & c7d478;
assign v37706b3 = hlock4_p & v372adaa | !hlock4_p & v372f071;
assign v8bc1c0 = hmaster2_p & v377b24b | !hmaster2_p & v35772a6;
assign v3a5a5ec = hlock3_p & v3734291 | !hlock3_p & v372f7d4;
assign v3a5de18 = hgrant6_p & v3761fb5 | !hgrant6_p & v376993b;
assign v3a6bdaa = hlock4_p & v37767e6 | !hlock4_p & v8455cb;
assign v3754981 = hmaster0_p & v372658a | !hmaster0_p & v375a086;
assign v377de7f = hmaster0_p & v3a70133 | !hmaster0_p & v8455ab;
assign v373b077 = hmaster1_p & v37693fe | !hmaster1_p & v3a5ad4f;
assign v3a60d5e = hmaster2_p & v1e37370 | !hmaster2_p & v3727db5;
assign v373c612 = hgrant4_p & v8455ab | !hgrant4_p & d5959b;
assign v3a7031b = hmaster2_p & v37613a8 | !hmaster2_p & v3a6fad2;
assign v3a69c6f = hbusreq3_p & v3a6f940 | !hbusreq3_p & v37281d0;
assign v375a677 = hgrant6_p & v8455ab | !hgrant6_p & v372f16b;
assign v376aa54 = hmaster0_p & v3a664b5 | !hmaster0_p & v375b0e4;
assign v3739885 = hmaster3_p & v374a20f | !hmaster3_p & v3a6ae54;
assign v377e090 = hbusreq2 & v3a6fdb4 | !hbusreq2 & v372cc25;
assign v376bb7a = hmaster0_p & v372fb58 | !hmaster0_p & !v3771c85;
assign v3a68d3f = hgrant3_p & v8455be | !hgrant3_p & !v3779ac2;
assign v37751d9 = hlock4_p & bbab81 | !hlock4_p & !v8455ab;
assign v377efa7 = hmaster0_p & v375c0d6 | !hmaster0_p & v3a6fec4;
assign v3743113 = hmaster2_p & v372d8e8 | !hmaster2_p & !v3750e32;
assign v373461a = hmaster1_p & v375f852 | !hmaster1_p & v3a7080c;
assign v3a6ffb6 = hbusreq1_p & v3751a0b | !hbusreq1_p & v8455b0;
assign v374e463 = jx0_p & v3758b25 | !jx0_p & v3735a77;
assign v374cb02 = hbusreq7 & v3a69057 | !hbusreq7 & v3728464;
assign v3752535 = hbusreq7_p & v3774314 | !hbusreq7_p & !v374b5bc;
assign v3a5a16a = hbusreq0 & v3a6c007 | !hbusreq0 & v3a5f9e6;
assign v3734df5 = hlock5 & v3a6049f | !hlock5 & v35b779e;
assign v374be59 = hbusreq4_p & v3750e94 | !hbusreq4_p & !v8455ab;
assign v3a59dc4 = hgrant2_p & v375e7cc | !hgrant2_p & v3a6fbb4;
assign v374f526 = hbusreq5_p & v3755aae | !hbusreq5_p & v3a5b9cd;
assign v372fa02 = hbusreq2_p & v3733da3 | !hbusreq2_p & v3763eac;
assign v1e37d3a = hmaster2_p & v373e114 | !hmaster2_p & v3a5fc34;
assign v377f7dd = hbusreq8_p & v8455ab | !hbusreq8_p & v3722dd5;
assign v3a70601 = hbusreq5_p & v96f7ab | !hbusreq5_p & v3727d18;
assign v3a6ecb7 = hgrant5_p & v3770c2a | !hgrant5_p & v3a70015;
assign v3a70a22 = hbusreq8_p & v1e3778c | !hbusreq8_p & v375cebd;
assign v374776e = hbusreq0 & v3749e5a | !hbusreq0 & v372b4c0;
assign v3a59c65 = hgrant4_p & v3a53eeb | !hgrant4_p & v372ed34;
assign v3766da7 = hmaster2_p & v373ea71 | !hmaster2_p & v3759379;
assign v3758f02 = hmaster0_p & v3a70462 | !hmaster0_p & v3a707f5;
assign v1e37a9d = hlock8 & v37667eb | !hlock8 & v3760e1b;
assign v3a680cb = hgrant5_p & v8455ab | !hgrant5_p & v3a6d31d;
assign v37503ec = hbusreq6 & v37738fc | !hbusreq6 & v35b774b;
assign v375ce8d = hmaster0_p & v3765cec | !hmaster0_p & v3766d24;
assign v3742dfb = hmaster0_p & v3744104 | !hmaster0_p & v3758174;
assign v377ec28 = hbusreq6 & v374f307 | !hbusreq6 & v8455ab;
assign v3a56d78 = hgrant6_p & v8455e7 | !hgrant6_p & v3a70a05;
assign v3a70e2f = hbusreq5_p & a85c8e | !hbusreq5_p & !v8455ab;
assign v377d7dd = hgrant0_p & v376ea4a | !hgrant0_p & !v373aa77;
assign v37275a7 = hgrant1_p & v372373f | !hgrant1_p & v37328bf;
assign v37c1a6f = hbusreq3_p & v375c0cb | !hbusreq3_p & v3a69765;
assign v3725bdd = hgrant5_p & v3776cad | !hgrant5_p & v2acaeeb;
assign v3a61cd7 = hgrant4_p & v8455c2 | !hgrant4_p & v3779fd9;
assign v3725360 = hbusreq6 & v373a568 | !hbusreq6 & v3735525;
assign v377e73f = jx0_p & v3a712b5 | !jx0_p & v3748282;
assign v3a5ef6e = hbusreq6 & v37745b8 | !hbusreq6 & v377bfc0;
assign v373b16f = hlock5_p & v8455ab | !hlock5_p & v8455e7;
assign v3a70f6d = hbusreq8_p & v3764e3f | !hbusreq8_p & v3a60276;
assign v374e47e = hmaster2_p & v3776ada | !hmaster2_p & v3a596c4;
assign v3a70107 = hmaster1_p & v374314f | !hmaster1_p & v3778eed;
assign v374c4e1 = hbusreq1 & v375de18 | !hbusreq1 & !v373c755;
assign v377e0b8 = hgrant4_p & v23fde7c | !hgrant4_p & v3778da6;
assign v3a703f7 = hbusreq5_p & v377de7f | !hbusreq5_p & v377b838;
assign v37558d3 = hbusreq5 & v3a6f47a | !hbusreq5 & v3a635ea;
assign v374aa1b = hmaster0_p & v376eb33 | !hmaster0_p & !v3764585;
assign v37448a7 = hmaster1_p & v3a70b35 | !hmaster1_p & v3724df8;
assign v3a633c5 = hbusreq5 & v3729eb0 | !hbusreq5 & v8455ab;
assign v3a6eb2a = hbusreq2 & v39a537f | !hbusreq2 & v8455ab;
assign v3a64235 = stateA1_p & v8455ab | !stateA1_p & !v3a69ad1;
assign v3a6f338 = hbusreq6 & v35b779f | !hbusreq6 & v3765261;
assign v376bc32 = hmaster0_p & v375049a | !hmaster0_p & v376132a;
assign v3a66210 = hbusreq5_p & v37775ff | !hbusreq5_p & v377b706;
assign v3754076 = hbusreq3_p & v376a20e | !hbusreq3_p & v3757663;
assign v3748347 = hgrant6_p & v377e1d0 | !hgrant6_p & v3769f2f;
assign v2acb0e4 = hmaster1_p & v3753e6f | !hmaster1_p & v8e42b4;
assign v376a863 = hmaster0_p & v8455e7 | !hmaster0_p & v3767419;
assign v3775ec8 = hbusreq7_p & v3771622 | !hbusreq7_p & v3a6dbbf;
assign v3753cc4 = hlock0_p & v3757082 | !hlock0_p & v3a6ff43;
assign v374cd37 = hmaster1_p & v8455ab | !hmaster1_p & v376575a;
assign v3a711c9 = hgrant0_p & v3a714c6 | !hgrant0_p & v8455ab;
assign v3a70fa8 = hmaster0_p & v2619aa5 | !hmaster0_p & v3a65752;
assign v3744751 = hbusreq7 & v3741608 | !hbusreq7 & cb0c12;
assign v3762452 = hmaster1_p & v372455c | !hmaster1_p & v373a9ef;
assign v375a28a = hlock3 & v3a583f5 | !hlock3 & v37735ec;
assign v372f3b1 = hmaster2_p & v8455b0 | !hmaster2_p & v377ef4a;
assign v373e57b = hmaster1_p & v3a5d2c5 | !hmaster1_p & beab35;
assign v3734c40 = hmaster0_p & v3a70ce7 | !hmaster0_p & v3a6ef01;
assign v37573d2 = hmaster3_p & v3a709db | !hmaster3_p & v373ce66;
assign v3762037 = hlock0 & v3a635ea | !hlock0 & v374b274;
assign v377a91a = hlock5 & v360d195 | !hlock5 & v37522a0;
assign v3742b88 = hmaster0_p & v3727141 | !hmaster0_p & !v374b68a;
assign v3736ea9 = hbusreq5 & v373e55b | !hbusreq5 & v8455ab;
assign v37255d6 = hgrant8_p & v8455ab | !hgrant8_p & !v3760198;
assign v375c740 = hmaster0_p & v373b1ae | !hmaster0_p & v8455ab;
assign v3a5b903 = hbusreq4_p & v3a5d40d | !hbusreq4_p & v8455ab;
assign v37507be = hbusreq3 & v35b9d52 | !hbusreq3 & !v8455ab;
assign v3a70d19 = hmaster1_p & v3758dcb | !hmaster1_p & v3a6096a;
assign v373a7f7 = hlock7_p & v3a60026 | !hlock7_p & v3a712a5;
assign v376964c = hmaster3_p & v3746085 | !hmaster3_p & v3a66988;
assign v3774fee = hmaster1_p & v373a2f4 | !hmaster1_p & !v3755096;
assign v2678ca9 = decide_p & v3732da0 | !decide_p & v374efeb;
assign v375aa6b = hlock0 & v37771ca | !hlock0 & v3a6b51b;
assign v37469db = hgrant1_p & v3735e39 | !hgrant1_p & v3809adf;
assign v1e3735b = hgrant4_p & v377dee0 | !hgrant4_p & v372372d;
assign v3a7124d = hmaster0_p & v3a712f6 | !hmaster0_p & !v3774a9c;
assign v37718de = hgrant6_p & v3a65eba | !hgrant6_p & v3a56898;
assign v3735ecd = hgrant4_p & v3a2ad1b | !hgrant4_p & v373fd72;
assign v3a6b3d4 = hgrant6_p & v8455ab | !hgrant6_p & v37535bd;
assign v3a7118a = hbusreq6 & v3a703d0 | !hbusreq6 & v3a6f61f;
assign v3739082 = hmaster2_p & v373d9e0 | !hmaster2_p & v375f9e9;
assign v37434ce = hgrant6_p & v37285ad | !hgrant6_p & v3a6fc6a;
assign v3754403 = hgrant4_p & v8455ab | !hgrant4_p & v3a70e70;
assign v375240c = hmaster0_p & v377a121 | !hmaster0_p & v375d8a6;
assign v3746c51 = hbusreq3_p & v3a6a41e | !hbusreq3_p & v8455ab;
assign v375ddb7 = hbusreq2 & v3a5fcbc | !hbusreq2 & v3a70a88;
assign v375da9d = hbusreq0 & v377a9cb | !hbusreq0 & v3a7044a;
assign v3764683 = hmaster2_p & v3a624da | !hmaster2_p & v37604e9;
assign v374a3b7 = hbusreq5 & v373144a | !hbusreq5 & v3a6f45c;
assign v3a55ec8 = jx3_p & v1e37c79 | !jx3_p & v373782c;
assign v9d70f0 = hmaster1_p & v3749469 | !hmaster1_p & v3747271;
assign v372f4ce = hmaster1_p & v3a67b62 | !hmaster1_p & !v375c0f1;
assign v3768953 = hmaster2_p & v3a5979b | !hmaster2_p & v3a70fec;
assign v3a6934e = hmaster0_p & v37712aa | !hmaster0_p & v3a70caa;
assign v372f202 = hmaster0_p & v3777da5 | !hmaster0_p & v3a611bd;
assign v3a6267a = hgrant5_p & v377209b | !hgrant5_p & v3a55861;
assign b4389d = hmaster1_p & v3726339 | !hmaster1_p & v372e749;
assign v3a5574a = hbusreq2_p & v3760343 | !hbusreq2_p & v3724f7b;
assign v3a6e0f2 = hgrant2_p & v8455ba | !hgrant2_p & v3a6b4d7;
assign v3a6f54c = hmaster2_p & v3762e13 | !hmaster2_p & v3a6935c;
assign v3a533d8 = hmaster2_p & v39ea76e | !hmaster2_p & v3a6d684;
assign v377ab1f = hbusreq6_p & v3779060 | !hbusreq6_p & !v3a6dfb2;
assign v3a7167e = hgrant6_p & v8455ab | !hgrant6_p & !v3751aaa;
assign v3a701d1 = hbusreq2_p & v3747346 | !hbusreq2_p & v3773856;
assign v375e3a1 = jx1_p & v375ab04 | !jx1_p & v373628a;
assign v37446b1 = hbusreq7 & v37472ea | !hbusreq7 & v8455ab;
assign v3759efd = hmaster0_p & v3741c91 | !hmaster0_p & v3a708e7;
assign v3a6f31c = hgrant6_p & v372abd8 | !hgrant6_p & v3778173;
assign v3778b8d = hlock2 & v37370f8 | !hlock2 & v373e521;
assign v373b288 = locked_p & v3a635ea | !locked_p & !v35772a5;
assign v3726570 = hgrant1_p & v3a5c945 | !hgrant1_p & !v372c11d;
assign v3a558f6 = hgrant3_p & v8455ab | !hgrant3_p & v3725cbf;
assign v3774eec = hmaster1_p & v3762eeb | !hmaster1_p & v37698c3;
assign v3a6fbe6 = hbusreq6 & v377834b | !hbusreq6 & v3a62a6d;
assign v3809e41 = hgrant7_p & v8455ab | !hgrant7_p & !v3a70306;
assign v3a6b643 = hbusreq5 & v1e377f7 | !hbusreq5 & v3a700af;
assign v376aba9 = hbusreq4 & v3a5dd17 | !hbusreq4 & v3a704b0;
assign v3731780 = hmaster1_p & v37245f8 | !hmaster1_p & v3767ef0;
assign v3a715ac = hgrant4_p & v3a6fc83 | !hgrant4_p & v3a6fef1;
assign v376636b = jx1_p & v3a6f269 | !jx1_p & dc6ab1;
assign v1e37b3f = hgrant6_p & v373f03e | !hgrant6_p & v8455ab;
assign v3a713f6 = hbusreq7 & v374845f | !hbusreq7 & ce8abd;
assign v377a42f = hbusreq0_p & v3723b00 | !hbusreq0_p & v8455ab;
assign v3a70303 = hbusreq2_p & v374513e | !hbusreq2_p & !v37392ad;
assign v3769ce7 = hlock7 & v3a6f7d5 | !hlock7 & v375d997;
assign v374558a = hmaster0_p & v375808f | !hmaster0_p & v37743e0;
assign v3760799 = hmaster2_p & v372424e | !hmaster2_p & v3a5e070;
assign v374f654 = hbusreq4 & v377928c | !hbusreq4 & v8455ab;
assign v3a6f9df = hbusreq6 & v3a58429 | !hbusreq6 & v3736679;
assign v3775072 = hlock5 & v3a63e9d | !hlock5 & v374a7de;
assign v3730ae6 = hmaster1_p & c63c1f | !hmaster1_p & v3a6a68c;
assign v3a6a4b9 = hbusreq5 & v3a69539 | !hbusreq5 & v376bc32;
assign v37297e4 = hgrant6_p & v3730e2a | !hgrant6_p & v3257329;
assign v374e39c = hmaster2_p & v3a6d3c5 | !hmaster2_p & v37283fe;
assign v3775999 = hgrant6_p & v375da82 | !hgrant6_p & v23fd967;
assign v373c00f = hbusreq5 & v3a701a1 | !hbusreq5 & v3760513;
assign v373340f = hmaster1_p & v3776b22 | !hmaster1_p & v3770ecc;
assign v88d9b8 = hmaster2_p & v37550d4 | !hmaster2_p & v3729864;
assign v3a5e0c9 = hgrant8_p & v375023c | !hgrant8_p & v3a7038d;
assign v3a57214 = hbusreq6 & v3a70f43 | !hbusreq6 & v3a58102;
assign v372eec6 = hbusreq7_p & v3a70d29 | !hbusreq7_p & v3a6ebe8;
assign v373b983 = hbusreq2 & v374f87c | !hbusreq2 & v8455ab;
assign v377adf7 = hmaster0_p & v3a7112c | !hmaster0_p & v3748f81;
assign v3735b5a = hbusreq5_p & v37691ab | !hbusreq5_p & v3a6f11b;
assign v3749b2e = hmaster3_p & v375b777 | !hmaster3_p & v375889d;
assign v37695f7 = hbusreq5_p & v3776c82 | !hbusreq5_p & !v372abb9;
assign v3a702aa = hbusreq0_p & v39a537f | !hbusreq0_p & !v39a5381;
assign v372b60b = hmaster0_p & v3a70f08 | !hmaster0_p & v377a083;
assign v3a6eb36 = hmaster0_p & v23fe061 | !hmaster0_p & v3a692f6;
assign v377a88e = hbusreq4_p & v3730aaf | !hbusreq4_p & v372cc25;
assign v377583c = hgrant5_p & v3738a70 | !hgrant5_p & v3258760;
assign v374a36a = jx0_p & v373de83 | !jx0_p & v372cc3d;
assign v3a70a3d = hmaster3_p & v3a68183 | !hmaster3_p & v37256c0;
assign v3a6fed2 = hgrant3_p & v8455ab | !hgrant3_p & v3a6f9a0;
assign v3768a3c = hmaster2_p & v8455ab | !hmaster2_p & v3a6f8af;
assign v3a70df9 = hmastlock_p & v23fda2f | !hmastlock_p & v8455ab;
assign v376b4e5 = hbusreq4_p & v3a6c68c | !hbusreq4_p & v8455ab;
assign v9bd777 = hbusreq5_p & v3724e4b | !hbusreq5_p & v374c837;
assign v3a58cd4 = hlock4 & v377ec50 | !hlock4 & v3a6ebfb;
assign v3a596c4 = hgrant4_p & v8455ab | !hgrant4_p & v377b0f7;
assign v380956b = hmaster2_p & v3753f1a | !hmaster2_p & !v8455e7;
assign v3a53ce6 = hlock5 & v37347b2 | !hlock5 & v372afe7;
assign v3a67095 = hmaster0_p & v3a5b8a2 | !hmaster0_p & v3742f25;
assign v372476f = hmaster0_p & v375ceff | !hmaster0_p & v3a7062d;
assign v3730553 = hmaster2_p & v8455b3 | !hmaster2_p & v3760f4e;
assign v33790c9 = hbusreq8_p & v3a5406b | !hbusreq8_p & v3748e82;
assign v3a6adff = hmaster2_p & v37283bb | !hmaster2_p & v373b687;
assign v38090ee = hgrant4_p & v3a602c3 | !hgrant4_p & v374700b;
assign v3a540a1 = hbusreq5 & v3a673d3 | !hbusreq5 & v3a6fa44;
assign v3772e0c = hgrant4_p & v8455e7 | !hgrant4_p & !v3a6fc7d;
assign v3a6a36d = hmaster2_p & v3757568 | !hmaster2_p & v3750d37;
assign v3775729 = hgrant5_p & v8455ab | !hgrant5_p & v3a70aa3;
assign v37506fe = hbusreq7 & v37551eb | !hbusreq7 & v3768082;
assign v3a5445e = hmaster1_p & v373523c | !hmaster1_p & v3a5b98b;
assign v377d7a0 = hbusreq5 & v3751de0 | !hbusreq5 & v37538ca;
assign v37565a5 = hlock2 & v37567d3 | !hlock2 & v373e760;
assign v372ea51 = hgrant4_p & v376428f | !hgrant4_p & v3734f7b;
assign v39ea2e3 = hbusreq7_p & v3a69118 | !hbusreq7_p & v3764c6c;
assign v37629cf = hbusreq4 & v3a6fdd6 | !hbusreq4 & v373ea71;
assign v373b414 = hlock0_p & v3722e5c | !hlock0_p & v35772a6;
assign v374d7c1 = hbusreq6 & v3a6224d | !hbusreq6 & v3a70a7f;
assign v8a7af6 = hbusreq5_p & v377d7a0 | !hbusreq5_p & v3a68ee5;
assign v374f834 = hgrant5_p & v373a982 | !hgrant5_p & v3a68e10;
assign v374d547 = hgrant5_p & v8455ab | !hgrant5_p & !v3a585f1;
assign v37485c0 = hlock6_p & v28896da | !hlock6_p & v3750dd3;
assign v3748b83 = hmaster2_p & v3807aa1 | !hmaster2_p & v3a5979b;
assign v380958f = hbusreq7_p & v374731f | !hbusreq7_p & !v37678f8;
assign v3a6f901 = hmaster2_p & d1e3dd | !hmaster2_p & v375f2ba;
assign v3762153 = hmaster0_p & v375b0cd | !hmaster0_p & v8455b5;
assign v3a5f08f = hmaster2_p & v37325a2 | !hmaster2_p & v3a6a8ee;
assign v3748b9d = hmaster2_p & v3757863 | !hmaster2_p & v3774f35;
assign v3776615 = hbusreq3 & v3a7066e | !hbusreq3 & v37447bf;
assign v377b4cc = hbusreq0 & v374fb51 | !hbusreq0 & v3734d12;
assign v37739a8 = hgrant5_p & v3745e5e | !hgrant5_p & v3a6f6eb;
assign v372ea4b = hlock6 & v3a70995 | !hlock6 & v377aa23;
assign v3750e89 = hmaster0_p & v376cfc1 | !hmaster0_p & v3a69123;
assign v376f4b2 = hbusreq4_p & v3a5cc1a | !hbusreq4_p & !v3a7107a;
assign b00c46 = hmaster2_p & v8455ab | !hmaster2_p & !v3746289;
assign v3728b31 = hmaster0_p & v374729b | !hmaster0_p & !v3a54f8a;
assign v373e34e = hmaster0_p & v372c221 | !hmaster0_p & v3a60358;
assign v376d2dc = hbusreq4 & v3762a2a | !hbusreq4 & v373abde;
assign v375945f = hmaster2_p & v3a712e2 | !hmaster2_p & v3727e66;
assign v3a667b8 = hbusreq4 & v374ad16 | !hbusreq4 & v8455ab;
assign v3a6d4b7 = hbusreq4_p & v37652eb | !hbusreq4_p & v3736e8e;
assign v3779d91 = hbusreq7_p & v3734279 | !hbusreq7_p & v376ec4f;
assign v3a5c040 = hbusreq8 & v3a5b960 | !hbusreq8 & v3761351;
assign v375e309 = hbusreq1_p & v37345f5 | !hbusreq1_p & v3a5e8f6;
assign v3a703c3 = hbusreq6_p & v374c9cf | !hbusreq6_p & !v8455ab;
assign v3747c3e = locked_p & v3a58cd5 | !locked_p & v8455ab;
assign v3767304 = hbusreq2_p & v37274be | !hbusreq2_p & v3731be6;
assign v3732715 = hbusreq3 & v3a6abaa | !hbusreq3 & v3763d3a;
assign v3a550cd = hmaster2_p & v3731a49 | !hmaster2_p & v37745c3;
assign v3728903 = hmaster0_p & v3a6de4f | !hmaster0_p & v3a59649;
assign v3a6fa88 = hgrant4_p & v374672f | !hgrant4_p & v373ebf9;
assign v3a5e985 = hmaster1_p & v374bfa2 | !hmaster1_p & v3a6fe5f;
assign v3a6f38b = hmaster1_p & v3748e09 | !hmaster1_p & v3a6f6fe;
assign v374ab8d = hbusreq4_p & v3765c6d | !hbusreq4_p & v8455ab;
assign v3a6f0f2 = hlock0 & v37285eb | !hlock0 & v3a71566;
assign v3a7121f = hbusreq5_p & v3a707e0 | !hbusreq5_p & v37780e2;
assign v3732ecb = hmaster2_p & v3740f3d | !hmaster2_p & !v3757aa1;
assign v3753ee5 = hlock8_p & v375e2de | !hlock8_p & v3a63ef6;
assign v375d3fd = hmaster2_p & v3a7010e | !hmaster2_p & v3762475;
assign v3752caa = hbusreq5_p & v3735bbb | !hbusreq5_p & v3806fe2;
assign v373fc52 = hmaster3_p & v3a69203 | !hmaster3_p & v3a5ecb9;
assign v3a6fc4a = hbusreq5_p & v373cae5 | !hbusreq5_p & !v3a6f6a8;
assign v3760343 = hlock2 & v3765c85 | !hlock2 & v3a6e3bb;
assign v3751d73 = hbusreq4_p & v3a630db | !hbusreq4_p & v35772a6;
assign v3a5d822 = hlock0_p & v374362e | !hlock0_p & v3a66673;
assign v37403fe = hmaster2_p & v3a5600a | !hmaster2_p & v374ebb0;
assign v3a6f2ad = hbusreq4 & v3a6e804 | !hbusreq4 & v3748797;
assign v372a0b0 = hbusreq2_p & v376d79d | !hbusreq2_p & v8455ab;
assign v377af5d = hmaster1_p & v3a582c5 | !hmaster1_p & v374c1a0;
assign dcb1a9 = hmaster2_p & v3776ada | !hmaster2_p & v373222d;
assign v3a65df3 = hbusreq5_p & v3753f77 | !hbusreq5_p & v3a58c07;
assign v3731dfe = hmaster2_p & v3a635ea | !hmaster2_p & v377c6ce;
assign v3a70388 = hmaster2_p & v373d791 | !hmaster2_p & v373e1d0;
assign v3736ebd = hbusreq3_p & v37652b1 | !hbusreq3_p & !v8455ab;
assign v3806388 = hbusreq3_p & v2092ffc | !hbusreq3_p & v3772596;
assign v9fc6a0 = hbusreq5 & v377730a | !hbusreq5 & v3770f76;
assign v3a70c85 = hmaster0_p & v374306c | !hmaster0_p & v375b5d3;
assign v3776b18 = hlock2_p & v3750d37 | !hlock2_p & !v8455ab;
assign v373edbe = hbusreq2_p & v3a6efe8 | !hbusreq2_p & v3a5e80e;
assign v3a71345 = stateG10_1_p & v3a635ea | !stateG10_1_p & v372dec8;
assign v37418ac = hbusreq6_p & v3745452 | !hbusreq6_p & v374760a;
assign v3a70dba = hgrant5_p & v37575fd | !hgrant5_p & v380776b;
assign v37283ea = jx1_p & v3765443 | !jx1_p & v3728723;
assign v37784a0 = hmaster0_p & v3a71186 | !hmaster0_p & v3741b5e;
assign v37400f8 = hlock2_p & v374306c | !hlock2_p & v3a6ffae;
assign v3a66c66 = hmaster2_p & v3a65da7 | !hmaster2_p & v3a5e7fe;
assign v3a6f2b8 = hbusreq3_p & v3748797 | !hbusreq3_p & v372f8d3;
assign v375dbeb = hlock0_p & a9f66a | !hlock0_p & v37416f0;
assign v376c7f9 = hmaster0_p & v3777226 | !hmaster0_p & v2092ec6;
assign v3a611e6 = hbusreq4_p & v3778281 | !hbusreq4_p & v37297af;
assign v894fb9 = hgrant5_p & v8455ab | !hgrant5_p & v3753592;
assign v3a70e2d = hmaster1_p & v377d1dc | !hmaster1_p & v3a64abe;
assign v372449f = hbusreq0 & v374b18c | !hbusreq0 & v3a5f20d;
assign v377f730 = hlock3_p & v3724e61 | !hlock3_p & !v8455ab;
assign v3a6f944 = hmaster1_p & v2aca977 | !hmaster1_p & v3a70f51;
assign v3723df5 = hmaster3_p & v3a5ee7e | !hmaster3_p & v3763ca5;
assign v372e61a = hbusreq2 & v373e9a9 | !hbusreq2 & v37749bf;
assign v3a702ee = hbusreq4_p & v37725ea | !hbusreq4_p & !v8455ab;
assign v3a708cf = hlock4 & v3a69a39 | !hlock4 & v372952e;
assign v3771162 = hmaster1_p & v3a70d99 | !hmaster1_p & v3a55c2f;
assign v3a6eac1 = hgrant3_p & v8455ab | !hgrant3_p & v373fff3;
assign v376ee43 = hmaster0_p & v37451b8 | !hmaster0_p & v3762ffa;
assign v3a7140d = hmaster3_p & v8455ab | !hmaster3_p & !v3a71327;
assign v373d89b = hbusreq7 & v3a54769 | !hbusreq7 & v3759284;
assign v3724a6e = hlock0_p & v3a709ea | !hlock0_p & v375ecc7;
assign v376702c = hbusreq7_p & v3757231 | !hbusreq7_p & !v3739368;
assign v373b748 = hbusreq4 & v3a70e5a | !hbusreq4 & v2092abe;
assign v8455b3 = hlock0_p & v8455ab | !hlock0_p & !v8455ab;
assign v3a706c1 = hmaster0_p & v377a477 | !hmaster0_p & !v3758ff0;
assign v3a6ff0c = hlock6_p & v3a70641 | !hlock6_p & v8455ab;
assign v372a77a = hlock5_p & v376e79d | !hlock5_p & v3a7121a;
assign v3a6a07b = hbusreq4 & v37454a8 | !hbusreq4 & v8455ab;
assign v37440a8 = hgrant2_p & v377aa23 | !hgrant2_p & v3a6ec6d;
assign start = v288971d;
assign v3728729 = hbusreq5 & v3a64df4 | !hbusreq5 & v8455ab;
assign v374d313 = hmaster2_p & v3742122 | !hmaster2_p & v8455ab;
assign v3767ee9 = hmaster0_p & v376aa57 | !hmaster0_p & v372a96f;
assign v377a434 = hbusreq4_p & v3a6f9c3 | !hbusreq4_p & v3759c49;
assign v3a6ebaf = hbusreq6 & v37363fd | !hbusreq6 & !v3a6feca;
assign v3a6337a = hbusreq5_p & v3809505 | !hbusreq5_p & v3a71133;
assign v3769c19 = jx0_p & v375e85e | !jx0_p & v3736d87;
assign v377457e = hbusreq8_p & v374d1b8 | !hbusreq8_p & v3a70e73;
assign v3a6faeb = hbusreq4_p & v3723296 | !hbusreq4_p & !v3a658bf;
assign v3a59f5a = hgrant5_p & v8455b5 | !hgrant5_p & v3774a95;
assign v3a5ad13 = hbusreq1_p & v3745b36 | !hbusreq1_p & v3772db0;
assign v3a70131 = hburst1 & v8455ab | !hburst1 & v3734c05;
assign v3735f56 = hlock0_p & v3a57f59 | !hlock0_p & !v3a66110;
assign v3a6982f = hbusreq8_p & v3769dcb | !hbusreq8_p & v3769fe3;
assign v376a7fc = hlock3 & v3a6ad19 | !hlock3 & v376129a;
assign db32f1 = hlock5_p & v8455ab | !hlock5_p & v373f042;
assign v3a5919f = hbusreq6_p & v373374d | !hbusreq6_p & v373dbc5;
assign v377e852 = hgrant5_p & v8455ab | !hgrant5_p & v37411ca;
assign v373e8ad = hbusreq3_p & v377cfd9 | !hbusreq3_p & !v372ee7e;
assign v3727477 = jx0_p & v373f408 | !jx0_p & v3747ced;
assign v374949f = hmaster0_p & v3a6f90e | !hmaster0_p & v3a296d8;
assign v377422b = hbusreq0 & v37772d5 | !hbusreq0 & v8455ab;
assign v3a5912f = hmaster0_p & v1e3780e | !hmaster0_p & v3a71609;
assign v3740e7d = hgrant2_p & v8455ab | !hgrant2_p & v37280de;
assign v375055f = hbusreq7 & v3737298 | !hbusreq7 & v377a2b2;
assign v3a53356 = hlock2 & v376cc8d | !hlock2 & v3728cfe;
assign v3a5dbc7 = hgrant2_p & ae0781 | !hgrant2_p & v3a638fe;
assign v3759d5a = hbusreq2_p & v37705d1 | !hbusreq2_p & v3a709aa;
assign v3758850 = hbusreq0 & v3a69bbd | !hbusreq0 & v8455ab;
assign v37590fb = hmaster2_p & v3a6823d | !hmaster2_p & !v8455ab;
assign v374e210 = hmaster0_p & v3a63ea7 | !hmaster0_p & v3a5ce54;
assign v3754e8c = hbusreq5_p & v3766cfc | !hbusreq5_p & !v377ce5a;
assign v3a5b1a3 = hbusreq4 & v373935b | !hbusreq4 & v3a58ea7;
assign v37308ae = hmaster1_p & v3a5e24e | !hmaster1_p & v1e37d71;
assign v3a69427 = hlock8_p & v3a56a0d | !hlock8_p & !v3774369;
assign v374a516 = jx0_p & v377012f | !jx0_p & v3a65c47;
assign v3767c44 = hbusreq0_p & v3a70e52 | !hbusreq0_p & v8455ab;
assign v3809e72 = hgrant5_p & v373f6b1 | !hgrant5_p & v374801f;
assign v376b28c = hmaster1_p & v3a6fa7a | !hmaster1_p & v3a5c93e;
assign v3a6a2ab = hmaster0_p & v375b282 | !hmaster0_p & !v373ca5f;
assign v3a7022c = hmaster2_p & v377b330 | !hmaster2_p & v3a6f4c7;
assign v37377f0 = hbusreq8_p & v8455ab | !hbusreq8_p & v375b239;
assign v3a70133 = hmaster2_p & v3748797 | !hmaster2_p & v8455ab;
assign v3a61d9f = hmaster0_p & v3a5a807 | !hmaster0_p & v8455e7;
assign v3735708 = hgrant6_p & v3a5a63c | !hgrant6_p & v3724577;
assign v3a62ccf = hmaster0_p & v3742d95 | !hmaster0_p & v3a610a4;
assign v372bdc2 = hbusreq5_p & v3a6eb22 | !hbusreq5_p & v373c00f;
assign v3758c32 = hbusreq0 & v375dcf5 | !hbusreq0 & v37375e4;
assign v374237b = hmaster1_p & v37357d9 | !hmaster1_p & !v3a5744d;
assign v3730e74 = hbusreq4_p & v375ce35 | !hbusreq4_p & v374baac;
assign v3750700 = hgrant5_p & v3a69409 | !hgrant5_p & v3a6f087;
assign v37258e7 = hbusreq5_p & v3a6a7cb | !hbusreq5_p & v3a6f423;
assign v37644ce = hmaster2_p & v8455ab | !hmaster2_p & v3734916;
assign v372d891 = hbusreq5 & v3730bae | !hbusreq5 & v377984a;
assign v3752c29 = hbusreq2 & v3766e5d | !hbusreq2 & v3757955;
assign v3726aa5 = hbusreq1 & v37482f8 | !hbusreq1 & !v372b24d;
assign v3a6fcc5 = hbusreq0_p & v3731e8c | !hbusreq0_p & v8455b5;
assign v3758bc2 = hmaster0_p & v3734585 | !hmaster0_p & v3a6fb52;
assign v3772ee4 = hgrant4_p & v377c94b | !hgrant4_p & v3774d12;
assign v3728179 = hmaster2_p & v3744ada | !hmaster2_p & v37273d2;
assign v3767631 = hmaster2_p & v3a579a3 | !hmaster2_p & !v8455ab;
assign v3763c9c = hmaster2_p & v3a6b94f | !hmaster2_p & v3a6a075;
assign v3759cc1 = hmaster0_p & v8455ab | !hmaster0_p & v3762cb2;
assign v3a70183 = hbusreq4_p & v3a5c65e | !hbusreq4_p & v3a6bb84;
assign v3754caa = hmaster2_p & v3736d47 | !hmaster2_p & v377ba59;
assign v376b031 = hmaster2_p & v373227a | !hmaster2_p & b318d6;
assign v377ca40 = hmaster2_p & v3a6dc08 | !hmaster2_p & v3a6fa39;
assign v3767e38 = hbusreq8_p & v3726980 | !hbusreq8_p & v3a63d5f;
assign v3a7049a = hbusreq4_p & v373a33d | !hbusreq4_p & v373c8cb;
assign v3a5d373 = hgrant2_p & v37516cc | !hgrant2_p & !v376674a;
assign v3809d49 = hbusreq4 & v374f307 | !hbusreq4 & v8455ab;
assign v3a5948d = hgrant6_p & v37379fc | !hgrant6_p & v3741f39;
assign v3755096 = hbusreq5_p & v3a6d9da | !hbusreq5_p & !v3736471;
assign v372e618 = hbusreq4 & v3778390 | !hbusreq4 & v375f9df;
assign v374ab5b = hbusreq1_p & v375cd0c | !hbusreq1_p & !v8455ab;
assign v3a5905e = jx1_p & v3a70eee | !jx1_p & v3a5ac5c;
assign v376ee7c = hgrant6_p & v8455ab | !hgrant6_p & v3747c0b;
assign v3768d56 = hbusreq8 & v3a70434 | !hbusreq8 & v373abcf;
assign v3746cdd = jx1_p & v8455ab | !jx1_p & v3a70681;
assign v37627bd = hbusreq6 & v3a65afa | !hbusreq6 & v8455ab;
assign v3a6ef96 = hbusreq7_p & v3a7067d | !hbusreq7_p & v3a680cb;
assign v374a0ae = hmaster2_p & v3762e13 | !hmaster2_p & v377e419;
assign v3768a7b = hlock8_p & v3757f96 | !hlock8_p & v37546c9;
assign v3765978 = hmaster1_p & v376581d | !hmaster1_p & v8455e7;
assign v38072bc = jx0_p & d66718 | !jx0_p & v37332b8;
assign v372d741 = hbusreq2_p & v37765e1 | !hbusreq2_p & v3a6fefa;
assign v3752333 = hmaster2_p & v375e657 | !hmaster2_p & v8455ab;
assign v372c42d = hburst0_p & v845605 | !hburst0_p & v3746c8d;
assign v3a6f100 = hmaster1_p & a374cd | !hmaster1_p & v3a70fb7;
assign v375e73a = jx0_p & v8455ab | !jx0_p & v3a69dd2;
assign v3a70b10 = hbusreq7 & v3731f35 | !hbusreq7 & v3779749;
assign v3a64566 = hgrant1_p & v3a57f59 | !hgrant1_p & !v3a70ecf;
assign v3a71470 = hbusreq5 & v373a9ac | !hbusreq5 & v8455ab;
assign v33789d2 = hbusreq8 & v3749942 | !hbusreq8 & v8455ab;
assign v3a6f618 = hgrant6_p & v374530a | !hgrant6_p & !v372f1a0;
assign v3a715e8 = jx0_p & v3a6f7fa | !jx0_p & v37561e0;
assign v3a6f4df = hmaster2_p & v8455ab | !hmaster2_p & v3750c27;
assign v374178a = hbusreq4 & v373eecc | !hbusreq4 & v3a614cb;
assign v3779f51 = hmaster2_p & v372e95b | !hmaster2_p & v8455b0;
assign v3a64f2d = hgrant6_p & v37414b0 | !hgrant6_p & v3a6006c;
assign v3762fd0 = hlock8_p & v37376dd | !hlock8_p & v376dc03;
assign v376b5a4 = hmaster2_p & v8455ab | !hmaster2_p & v3774cde;
assign v3a5fc8d = hbusreq0 & v3a67b28 | !hbusreq0 & v3a70c63;
assign v37781b7 = hmaster2_p & v3750e32 | !hmaster2_p & v3744a0c;
assign v3743287 = hmaster0_p & v374d6bd | !hmaster0_p & v372b2ef;
assign v3a70cb1 = hlock6 & v3a6f0be | !hlock6 & v37314b5;
assign v3758dcb = hbusreq5_p & v3a5c3a0 | !hbusreq5_p & v375607f;
assign v3a60301 = hmaster0_p & v3771931 | !hmaster0_p & !v3755914;
assign v3a5a8ce = hbusreq0 & v3a6f993 | !hbusreq0 & v8455ab;
assign v3a6e872 = hmaster2_p & v3a6bf22 | !hmaster2_p & v3a6efeb;
assign v3a7147c = hmaster2_p & v375c5a8 | !hmaster2_p & v376ea4a;
assign v3a6f71d = stateA1_p & v37481c3 | !stateA1_p & !v8455ab;
assign v3a70f64 = hbusreq3_p & v3722f58 | !hbusreq3_p & v3a6c5fc;
assign v376761d = hmaster2_p & v376ccdf | !hmaster2_p & v374d52a;
assign v37277c2 = hbusreq0_p & v375039e | !hbusreq0_p & v376bb26;
assign v3731beb = hbusreq5 & v3744b3d | !hbusreq5 & v372476f;
assign v377cebd = hmaster0_p & v377d745 | !hmaster0_p & v374d339;
assign v3a5d6f9 = hbusreq7_p & v3730fb9 | !hbusreq7_p & v37258d0;
assign v373064e = hlock0_p & v8455ab | !hlock0_p & v39a5265;
assign a22759 = hlock0_p & v372dadb | !hlock0_p & v3a70bb3;
assign v376b6d8 = hmaster0_p & v3774647 | !hmaster0_p & v3a6765d;
assign v3a644ab = hgrant2_p & v3a67403 | !hgrant2_p & v3774cd5;
assign v3a71295 = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a64968;
assign v3766309 = hmaster0_p & baec07 | !hmaster0_p & v3774730;
assign v372e865 = hgrant5_p & v373a267 | !hgrant5_p & v37519e5;
assign v3a6ef5c = hgrant4_p & v374f304 | !hgrant4_p & !v377970b;
assign v3745bc4 = hgrant4_p & v8455ab | !hgrant4_p & v377dab6;
assign v374fad5 = hmaster0_p & v3a66110 | !hmaster0_p & !v372ced7;
assign v373a68a = hlock0 & v377c6b3 | !hlock0 & v3a711de;
assign v3a696ee = hmaster1_p & v3a6ffb6 | !hmaster1_p & v3770a8c;
assign v373bbd0 = hmaster0_p & v377bb57 | !hmaster0_p & v37654c4;
assign v37383da = hmaster0_p & v3748262 | !hmaster0_p & v3a6e318;
assign v2aca987 = hbusreq8 & v3779014 | !hbusreq8 & v375075b;
assign stateG10_1 = !v2678ca9;
assign v3a6ebfd = hbusreq3 & v376f148 | !hbusreq3 & v8455ab;
assign v376cef0 = hmaster1_p & v3a6f5d4 | !hmaster1_p & v8455b9;
assign v3730b23 = hlock2_p & v3739509 | !hlock2_p & v8455b0;
assign v3a5858c = hmaster3_p & v3777988 | !hmaster3_p & v3a5e7be;
assign v374ae00 = hmaster2_p & v8455b0 | !hmaster2_p & v3750a9c;
assign v3a6ac20 = hmaster0_p & v372911f | !hmaster0_p & v377cccb;
assign v3a5c5ca = hbusreq3_p & v3761224 | !hbusreq3_p & v3a6557d;
assign v3a57f59 = locked_p & v8455ab | !locked_p & !v3a66110;
assign v3a64e75 = hgrant5_p & v3a642ab | !hgrant5_p & v3746825;
assign v37621c1 = hmaster1_p & v3a6ffb6 | !hmaster1_p & v377c8fd;
assign v37355c9 = hmaster0_p & v375b429 | !hmaster0_p & v37574c0;
assign v3a67fe2 = hmaster1_p & v3a5b8b9 | !hmaster1_p & v3775610;
assign v377a993 = hbusreq7_p & v3a54b43 | !hbusreq7_p & !v377ed4b;
assign v3756b39 = hbusreq6 & v3760707 | !hbusreq6 & v373c965;
assign v3769948 = hbusreq5_p & v37409c7 | !hbusreq5_p & v3a619b8;
assign v375968a = hbusreq2_p & v8455ab | !hbusreq2_p & v377568c;
assign v3741f67 = hmaster2_p & v3a635ea | !hmaster2_p & v3733da4;
assign v3770f51 = hgrant0_p & v8455ab | !hgrant0_p & v373e8b5;
assign v374cb62 = hmaster2_p & v8455b0 | !hmaster2_p & v375070c;
assign v3a57ee9 = hmaster0_p & v376445f | !hmaster0_p & v377291b;
assign v373db82 = hbusreq8 & v3a6f9b4 | !hbusreq8 & v3741572;
assign v3a7166b = jx0_p & v8455c5 | !jx0_p & !v8455c1;
assign v3a54dfa = hlock4 & v37671b7 | !hlock4 & v3a70188;
assign v3758ff8 = hbusreq5 & v3a6dc91 | !hbusreq5 & v3764dac;
assign v3a5ba8f = hmaster2_p & v376e914 | !hmaster2_p & !v3a6eb39;
assign v37345f5 = hgrant1_p & v3a55e7d | !hgrant1_p & v8455e7;
assign v37706e9 = hmaster2_p & v372d203 | !hmaster2_p & v8455ab;
assign v3a682a1 = hgrant2_p & v3a653e4 | !hgrant2_p & !v3766eef;
assign v372b798 = hmaster0_p & v3772007 | !hmaster0_p & !v3a6e4cd;
assign v3a6f972 = hbusreq0_p & v3a68426 | !hbusreq0_p & v373c627;
assign v3a66920 = hbusreq7 & v377e431 | !hbusreq7 & v374d409;
assign v3a67b28 = hgrant6_p & v373cc5c | !hgrant6_p & v3757637;
assign v3a7131f = hbusreq8 & v37690fe | !hbusreq8 & v3806a1c;
assign v372ab06 = hmaster0_p & v3a6f4cb | !hmaster0_p & v372e58c;
assign v3a6d0ec = hbusreq0 & v3a6d32c | !hbusreq0 & v3a712b1;
assign v3a6a539 = stateA1_p & v2ff9190 | !stateA1_p & v3a70ad0;
assign v3807748 = hbusreq8 & v3a5bc76 | !hbusreq8 & v3a7071f;
assign v37362d7 = hgrant6_p & v3724c77 | !hgrant6_p & v3737511;
assign v373aaa8 = hlock0_p & v8455ab | !hlock0_p & v37700ee;
assign v3a715c4 = hbusreq8_p & v3a7167c | !hbusreq8_p & v3a703a0;
assign v3a71292 = jx0_p & v3729beb | !jx0_p & v37795e0;
assign v373c30e = hbusreq7_p & v3763086 | !hbusreq7_p & v3a578c3;
assign v3729189 = hmaster0_p & v372b32f | !hmaster0_p & v3761bee;
assign v3728d84 = hbusreq6_p & v3734b80 | !hbusreq6_p & v3a6f89d;
assign v3743f3b = hmaster0_p & v376e72d | !hmaster0_p & v3756a04;
assign v3a5ef76 = hmaster2_p & v3a6d1ce | !hmaster2_p & v3759daf;
assign v372c3d4 = hbusreq1_p & v37724ca | !hbusreq1_p & v8455ab;
assign v3766185 = hbusreq5_p & v38064dd | !hbusreq5_p & v374a9d4;
assign v3741343 = hmaster2_p & v375d800 | !hmaster2_p & v3a70e98;
assign v3a6fc08 = hbusreq8_p & v23fd869 | !hbusreq8_p & v3a62875;
assign v3255b53 = hlock5 & v3743165 | !hlock5 & v3744a91;
assign v3729ae9 = hbusreq4 & v3a6eddd | !hbusreq4 & v38078ed;
assign v375b3b7 = hbusreq8 & v3a68789 | !hbusreq8 & v39a53a1;
assign v376f0fb = hbusreq0 & v3a6261b | !hbusreq0 & v37695b1;
assign v376107b = hlock4_p & v3778ed4 | !hlock4_p & v8455e7;
assign v3763ff7 = hbusreq6_p & v3758166 | !hbusreq6_p & !v3a56e63;
assign v3a68916 = hbusreq7 & v3728455 | !hbusreq7 & v3745d1e;
assign v3730695 = hbusreq6_p & v3a7162d | !hbusreq6_p & v3778528;
assign v37476bd = hbusreq0 & v3a64b90 | !hbusreq0 & v37591f3;
assign v372cd50 = hmaster3_p & v3a709f0 | !hmaster3_p & !v3a58a0d;
assign v3770d22 = hbusreq4 & v3a5dc35 | !hbusreq4 & v37496fa;
assign v3728202 = hmaster2_p & v8455b5 | !hmaster2_p & v3a6fe1a;
assign v37293ee = hbusreq6 & v3724b1c | !hbusreq6 & v8455ab;
assign a7394c = hmaster2_p & v376bca9 | !hmaster2_p & v377d1dc;
assign v3a6fb4a = hmaster1_p & v3725198 | !hmaster1_p & a7b390;
assign v375cec2 = hmaster2_p & v376ce77 | !hmaster2_p & v37541ff;
assign v372cfad = hlock6_p & v372a5c8 | !hlock6_p & v3a6f5d1;
assign v3737f5a = hmaster1_p & v373664d | !hmaster1_p & v373cf66;
assign v2acb094 = hbusreq7 & v376e3a3 | !hbusreq7 & v372c83a;
assign v373a6bf = hmaster1_p & v375db64 | !hmaster1_p & b46885;
assign v372c8d1 = hbusreq2 & v35772c9 | !hbusreq2 & v8455ab;
assign v377e08c = hbusreq3 & v3a6fd79 | !hbusreq3 & !v8455ab;
assign v2ff9291 = hgrant6_p & v8455ab | !hgrant6_p & !v3a6f87f;
assign v3769a00 = hmaster0_p & v373359b | !hmaster0_p & !v3745b9c;
assign v376c8a4 = hbusreq7_p & v376bd2f | !hbusreq7_p & v3a5a75c;
assign v3a5f8a2 = hbusreq0 & v3a70261 | !hbusreq0 & v3a55d3b;
assign v3776084 = hbusreq7 & v3730df7 | !hbusreq7 & v8455ab;
assign v3a55290 = hgrant5_p & v8455ab | !hgrant5_p & v3762dc3;
assign v372a39d = hbusreq4 & v376d9aa | !hbusreq4 & v3a635ea;
assign v37486d7 = hmaster3_p & v8455ab | !hmaster3_p & v375b3b9;
assign v377eb7a = hgrant2_p & v31c3694 | !hgrant2_p & v3a6079f;
assign v376db8a = hgrant0_p & v8455ab | !hgrant0_p & !v3a70fc0;
assign v372538b = hbusreq3 & v3730cc8 | !hbusreq3 & v8455ab;
assign v3a700ef = hmaster1_p & v3a584d6 | !hmaster1_p & v37702dc;
assign v3a6efc0 = hbusreq5 & v375977c | !hbusreq5 & v377bc8e;
assign v3a55454 = hmaster2_p & v375fba5 | !hmaster2_p & !v8455ab;
assign v3807a80 = hbusreq4_p & v3774c1b | !hbusreq4_p & !v38099c1;
assign v3775219 = hmaster2_p & v3734f04 | !hmaster2_p & v8455ab;
assign v374074d = hlock2_p & v3749caa | !hlock2_p & !v8455ab;
assign v376c4fe = hbusreq3_p & v3a70cc5 | !hbusreq3_p & v3776fe2;
assign v3a6ebb1 = hgrant0_p & v35b774b | !hgrant0_p & v373eedf;
assign v375f077 = locked_p & v3a6ef8c | !locked_p & v3a619c0;
assign v3a70b0d = hbusreq1_p & v372f576 | !hbusreq1_p & !v8455ab;
assign v3768be2 = hbusreq6 & v3771c59 | !hbusreq6 & d1bf3b;
assign v374e016 = hmaster0_p & v3a63777 | !hmaster0_p & v3a6f529;
assign v375a6e6 = hlock2 & v37434f4 | !hlock2 & v3a5ad94;
assign v374fafa = hbusreq6_p & v3a595ba | !hbusreq6_p & v3a5bb64;
assign v372589e = hbusreq7_p & v37bfc8a | !hbusreq7_p & v3a59900;
assign v3761071 = hmaster0_p & v37400aa | !hmaster0_p & v3757966;
assign v3760e46 = hbusreq6 & v3a7062b | !hbusreq6 & v37452c7;
assign v3a6f662 = hbusreq5_p & v376a3f7 | !hbusreq5_p & v374de73;
assign v376dc6f = hmaster0_p & v3a6f9e4 | !hmaster0_p & v3a713e7;
assign v3a70caa = hmaster2_p & v3740c75 | !hmaster2_p & v3742f0a;
assign v37548be = hlock8_p & v3a68c63 | !hlock8_p & v374d12f;
assign v374ff44 = hbusreq2 & v377caa3 | !hbusreq2 & v8455bf;
assign v3742035 = hmaster2_p & v375ed6f | !hmaster2_p & v3a6eb2f;
assign v373443d = hbusreq5_p & v3765d5e | !hbusreq5_p & v3732c6a;
assign v375f27b = hbusreq5_p & v37281a4 | !hbusreq5_p & v8455ab;
assign v3a5de8f = hbusreq0 & v376dba6 | !hbusreq0 & v37539bc;
assign v3806ed4 = hmaster1_p & v3736d47 | !hmaster1_p & v3a5aad8;
assign v3738fe2 = hbusreq0 & v3a7024b | !hbusreq0 & v37609d6;
assign v375e2bc = hgrant4_p & v8455ab | !hgrant4_p & v3a6ad38;
assign v3a5bd24 = stateA1_p & v8455e1 | !stateA1_p & !v373c3bd;
assign v376ca02 = hbusreq5_p & v374cacb | !hbusreq5_p & !v3a70dab;
assign v372c1cf = hlock6_p & v3724204 | !hlock6_p & v8455b3;
assign v377a5df = hgrant6_p & v37379fc | !hgrant6_p & v3743ada;
assign v376435f = hbusreq4 & v373628e | !hbusreq4 & v3a60a68;
assign v377086b = hmaster2_p & v3a635ea | !hmaster2_p & v376b11e;
assign v3a6f232 = jx0_p & v3765734 | !jx0_p & v3757e56;
assign v8df61b = hbusreq2_p & v3a67629 | !hbusreq2_p & !v3728eeb;
assign v3a71307 = hmaster0_p & v3a582c5 | !hmaster0_p & v3a665b3;
assign v3a53904 = hmaster0_p & a8fef2 | !hmaster0_p & v94e9e0;
assign v373862e = hmaster0_p & v3a6f8ec | !hmaster0_p & v3753a65;
assign v3726cd4 = hmaster0_p & b00c46 | !hmaster0_p & v8455ab;
assign v3a6f411 = hbusreq7_p & v3a6ecd1 | !hbusreq7_p & v3725d5a;
assign cd3a92 = hbusreq2_p & v3760279 | !hbusreq2_p & v376278c;
assign v3a5787a = hbusreq4_p & v3a6fdcc | !hbusreq4_p & v373b671;
assign v3731d89 = hgrant6_p & v3730e2a | !hgrant6_p & d3c22f;
assign v377dab6 = hbusreq4_p & v3a7158f | !hbusreq4_p & v3a6bf41;
assign v375e177 = hbusreq5 & v374314f | !hbusreq5 & v8455b0;
assign v375d152 = hmaster0_p & v377ad9b | !hmaster0_p & v3737721;
assign v3768858 = hbusreq5 & v376e0b6 | !hbusreq5 & v3a5e030;
assign v37664ab = hbusreq3_p & v3a70dc0 | !hbusreq3_p & v37595c8;
assign v376acee = hbusreq0 & v377f4e5 | !hbusreq0 & v377c31d;
assign v373257d = hlock5_p & v3753dbd | !hlock5_p & v3754981;
assign v3764381 = hgrant6_p & v37379fc | !hgrant6_p & v3754543;
assign v3769f5f = hgrant6_p & v3a706b7 | !hgrant6_p & !v8455ab;
assign v23fdad1 = hmaster2_p & v37710c7 | !hmaster2_p & v3a5c85c;
assign v3723cff = hlock0_p & v3768ac7 | !hlock0_p & v8455ab;
assign v377d76b = hbusreq5_p & v3a70209 | !hbusreq5_p & v375fbf2;
assign v37bfc4d = hgrant6_p & v8455ab | !hgrant6_p & !v91a14c;
assign v32587ac = hmaster1_p & v3a6dc83 | !hmaster1_p & v3a6f5cb;
assign v3a55ab6 = hmaster1_p & v3a635ea | !hmaster1_p & v35b73a5;
assign v373b666 = hgrant2_p & v3a6db06 | !hgrant2_p & v372526e;
assign v37426ea = hmaster1_p & v377a18b | !hmaster1_p & v37300e3;
assign v3742c16 = hbusreq6_p & v2aca977 | !hbusreq6_p & v376f665;
assign v3a70ece = hgrant2_p & v374203a | !hgrant2_p & !v3768a79;
assign v3a6f3a1 = hbusreq6_p & v3a67729 | !hbusreq6_p & v37637d5;
assign v37549e2 = hmaster2_p & v375e53a | !hmaster2_p & v3a5bfe6;
assign v3733a17 = hmaster2_p & v3a5600a | !hmaster2_p & v376ddc6;
assign v88c50b = hgrant6_p & v9cc76d | !hgrant6_p & v3735a4f;
assign v3a687a7 = hbusreq0 & v3a71425 | !hbusreq0 & v374faa2;
assign v37285ad = hlock6 & v373bf4f | !hlock6 & v3778fec;
assign v376fac8 = hlock2_p & v8615d7 | !hlock2_p & v3a7108a;
assign v3a6521e = hgrant8_p & v8455ab | !hgrant8_p & v8455d1;
assign v3a584f1 = hbusreq4_p & v373ccc7 | !hbusreq4_p & v3a6f4f1;
assign v3a5617a = hlock3 & v374cb4a | !hlock3 & v3a6f149;
assign b4f302 = hbusreq2 & v377ea86 | !hbusreq2 & !v39a535f;
assign v3a6eeb7 = hbusreq7_p & v3a70795 | !hbusreq7_p & v373945c;
assign v3a66f0d = hgrant6_p & v3778967 | !hgrant6_p & v373fb30;
assign v3a6fd3d = hmaster0_p & v8455ab | !hmaster0_p & v372580e;
assign v3a704b6 = hlock5_p & v3a5c93e | !hlock5_p & v37264cb;
assign v377f298 = hmaster0_p & v3763175 | !hmaster0_p & v3735c5f;
assign v3a6f55b = hbusreq4_p & v3a5fc34 | !hbusreq4_p & v37416c6;
assign v374e4fd = hmaster0_p & v3a63805 | !hmaster0_p & v37684c3;
assign v3742ec5 = hgrant6_p & v8455ab | !hgrant6_p & v3758983;
assign v375b5b4 = hbusreq4_p & v3a57b3c | !hbusreq4_p & v8455ab;
assign v3a70a32 = hbusreq4_p & d23bf8 | !hbusreq4_p & !v1e38224;
assign v3a702da = hmaster2_p & v37480b7 | !hmaster2_p & !v3a6f42a;
assign v3774131 = jx0_p & v360d144 | !jx0_p & v373c72a;
assign v3731fc6 = hbusreq6 & v8455ab | !hbusreq6 & v3a710fc;
assign v3a69555 = hburst1_p & v845605 | !hburst1_p & !v8455ab;
assign v3743156 = hmaster1_p & v37653bf | !hmaster1_p & v3a6fef0;
assign v372ae4f = hlock8_p & v37435f1 | !hlock8_p & v37612d0;
assign v3a6a998 = hmaster2_p & v3774e41 | !hmaster2_p & v8455b3;
assign v3763188 = hmaster3_p & v3a6f710 | !hmaster3_p & v376b6fb;
assign v3a71116 = hbusreq5 & v372c6c4 | !hbusreq5 & v376e0f5;
assign v376a9aa = hbusreq5 & v3a6fc89 | !hbusreq5 & v3764dac;
assign v375aa47 = hlock1 & v3a712a3 | !hlock1 & v3a63621;
assign v374b35e = hmaster2_p & v374d4e6 | !hmaster2_p & v3744df8;
assign v3a58520 = hgrant0_p & v39a4d88 | !hgrant0_p & v2aca784;
assign v3767cfb = hbusreq2 & v3771d77 | !hbusreq2 & v3762502;
assign v3a5a68d = hbusreq4_p & v3a53f42 | !hbusreq4_p & v375b4d8;
assign v3a6f863 = hbusreq8_p & v3729c28 | !hbusreq8_p & v3a62eaa;
assign v3749993 = hmaster0_p & v3745803 | !hmaster0_p & v3a6cf46;
assign v3a69ad3 = hgrant6_p & v3734cb7 | !hgrant6_p & v372afda;
assign v3a6d3c5 = hgrant4_p & v8455ab | !hgrant4_p & v37554a1;
assign v376d6b2 = hlock4 & v376a3bb | !hlock4 & v3a649fd;
assign v375ee2e = hmaster0_p & v372673d | !hmaster0_p & v376d2c6;
assign v373cd5a = hmaster0_p & v3a6ffae | !hmaster0_p & v374d95a;
assign v372cfd2 = hbusreq4 & v3769e3a | !hbusreq4 & v3731230;
assign v3743966 = hmaster2_p & v3a70c39 | !hmaster2_p & v3753329;
assign v3a6f359 = hmaster2_p & v3732dac | !hmaster2_p & v372ec78;
assign v377a751 = hbusreq4 & v37314cb | !hbusreq4 & v8455ab;
assign v3a673fa = hgrant5_p & v3a70e2f | !hgrant5_p & !v8455ab;
assign v372af95 = hmaster1_p & v375047c | !hmaster1_p & v8455ab;
assign v3a70e85 = hbusreq2 & v3743f47 | !hbusreq2 & v8455ab;
assign v373a945 = hbusreq5_p & v3722ad4 | !hbusreq5_p & v3a61246;
assign v376b1aa = jx0_p & v37609c3 | !jx0_p & v3753af9;
assign v376c4ba = hmaster0_p & v9e8a9c | !hmaster0_p & v3760951;
assign v37624b2 = hburst1 & v8455ab | !hburst1 & v3a66464;
assign v35b7769 = hgrant6_p & v8455ab | !hgrant6_p & v3725678;
assign v3730c96 = hmaster0_p & v3a61a7f | !hmaster0_p & v3a64608;
assign v373d081 = hmaster1_p & v375f27b | !hmaster1_p & v1e37349;
assign v37703cb = hgrant5_p & v8455ab | !hgrant5_p & !v3727c6e;
assign v372b2ab = hbusreq0 & v3a711d8 | !hbusreq0 & v3808f45;
assign v3a6b4a2 = hmaster0_p & v3a68426 | !hmaster0_p & v3a5a17f;
assign v37372a1 = hmaster2_p & v374e51a | !hmaster2_p & v374f0f5;
assign v3728085 = jx0_p & v3769fa2 | !jx0_p & v8455ab;
assign v372dbb0 = jx0_p & v3745249 | !jx0_p & v3a56aa0;
assign v3a53bb3 = hbusreq2_p & v3a6fefa | !hbusreq2_p & v374b4a4;
assign v3736058 = hmaster0_p & v375058e | !hmaster0_p & v374a0eb;
assign v376dd91 = hgrant7_p & v8455ab | !hgrant7_p & v373be4d;
assign v372a298 = hlock7 & v377c965 | !hlock7 & v377981a;
assign v3a70ab3 = hbusreq8 & v3a6fb4f | !hbusreq8 & v3734279;
assign v3736785 = hbusreq3_p & v3a61853 | !hbusreq3_p & v8455ab;
assign v37341fd = hbusreq5_p & v3a633c5 | !hbusreq5_p & !v8455ab;
assign v374e5ac = hbusreq2_p & v376fac8 | !hbusreq2_p & !v37520db;
assign v375b34f = hgrant2_p & v3744b27 | !hgrant2_p & v38076a8;
assign v375eb78 = hbusreq1 & v37270d9 | !hbusreq1 & v8455e7;
assign v3a56580 = hbusreq4_p & v3769ad7 | !hbusreq4_p & v23fdeaf;
assign v2acb056 = hbusreq6 & v3723542 | !hbusreq6 & v37280b0;
assign v3760167 = hgrant5_p & v3748cb7 | !hgrant5_p & v37314d7;
assign v3a5fd18 = hbusreq5_p & v372ea02 | !hbusreq5_p & v372b418;
assign v375115e = hlock0 & v376bade | !hlock0 & v37672c8;
assign v8a0a3d = hmaster1_p & v373d091 | !hmaster1_p & v3a6edfb;
assign v3a6f430 = hlock4 & v37445d7 | !hlock4 & v3729a1c;
assign v372807c = hgrant6_p & v375f3e2 | !hgrant6_p & v38063dd;
assign v3a70dcd = hbusreq2 & v376a14f | !hbusreq2 & v8455ab;
assign v3766117 = hlock6 & v376cc1b | !hlock6 & v37474b8;
assign v37576f6 = hlock5 & v3758ff8 | !hlock5 & v3a6dc91;
assign v3732eb2 = hmaster2_p & v3759032 | !hmaster2_p & v376ea4a;
assign v37331df = hbusreq4 & v3a702c2 | !hbusreq4 & v8455ab;
assign v3729173 = hmaster2_p & v374c74f | !hmaster2_p & v372628c;
assign v377bea3 = hgrant4_p & v374880c | !hgrant4_p & v3774a12;
assign v988a3b = hlock8_p & v3764ecd | !hlock8_p & v3a64102;
assign v3a5b807 = hbusreq5 & v3773d27 | !hbusreq5 & v376a04d;
assign v3a6ce52 = hmaster2_p & v3a6f42a | !hmaster2_p & !v375fbbb;
assign v3762be8 = hgrant2_p & v8455ab | !hgrant2_p & !v3a61fd3;
assign v3a64bcf = hmaster1_p & v3761287 | !hmaster1_p & v3a707ab;
assign v37304b3 = hbusreq6_p & v376660c | !hbusreq6_p & v373c96e;
assign v375a67c = hbusreq4_p & v3a6ec04 | !hbusreq4_p & !v8455ab;
assign v3a6f849 = hbusreq0_p & v375803a | !hbusreq0_p & v37747fc;
assign v3a640ff = hbusreq4_p & v374baac | !hbusreq4_p & v3739cda;
assign v374f273 = jx1_p & v3a5e7e8 | !jx1_p & v3772f37;
assign v3767d7c = hbusreq3_p & v37598c6 | !hbusreq3_p & v3722f12;
assign v375da6a = hbusreq5_p & v37280b7 | !hbusreq5_p & v3a6f11e;
assign v3753fea = hgrant6_p & v3a63028 | !hgrant6_p & v376132e;
assign v3a69fe5 = hmaster1_p & v373a4e4 | !hmaster1_p & v3736b19;
assign v3a7014c = hlock0_p & v3725410 | !hlock0_p & v8455b7;
assign v3753163 = hbusreq3 & v375039e | !hbusreq3 & v375da10;
assign v3a6ff7d = hbusreq3 & v39a5381 | !hbusreq3 & v8455ab;
assign v23fd7d9 = hgrant0_p & v374f307 | !hgrant0_p & v3a70e52;
assign v3774416 = hbusreq3_p & v373a3e4 | !hbusreq3_p & v3a5af86;
assign v3747130 = hmaster2_p & v3768495 | !hmaster2_p & v3770bcd;
assign v3a5b1ca = hmaster0_p & v3775dbc | !hmaster0_p & v37301d8;
assign v37331e7 = hbusreq3_p & v3a71263 | !hbusreq3_p & v3a6f1a4;
assign v3809d8b = hbusreq0 & v3763252 | !hbusreq0 & v3a64af7;
assign v3a690a6 = hbusreq7_p & v3763c1f | !hbusreq7_p & v3725be9;
assign v3a6f270 = hbusreq8 & v3a64058 | !hbusreq8 & v3774bad;
assign v374148a = hlock7 & v37692e3 | !hlock7 & v3a6f697;
assign c0d46a = hgrant3_p & v3a6c2b6 | !hgrant3_p & !v374ac2c;
assign v372949c = hgrant3_p & v3733e9e | !hgrant3_p & v37498be;
assign v35772b3 = stateA1_p & v3752b8c | !stateA1_p & v3728b28;
assign v3a6f826 = hlock5_p & v3a56d04 | !hlock5_p & v8455ab;
assign v3808881 = hgrant2_p & v3a55723 | !hgrant2_p & !v3759a88;
assign v3a70b56 = hbusreq6 & v3a6e8d4 | !hbusreq6 & v376c4c5;
assign v3753900 = hmaster1_p & v3a7028a | !hmaster1_p & v373d8c3;
assign v3771d75 = hmaster2_p & v3754df4 | !hmaster2_p & v376d1bb;
assign v3a5db58 = hbusreq7 & v37602c4 | !hbusreq7 & v375da55;
assign v3a70b97 = hmaster0_p & v377d652 | !hmaster0_p & v3774055;
assign v3a5b474 = hbusreq2 & v3731115 | !hbusreq2 & v3a6a4d4;
assign v376c2da = hlock6_p & v3769f88 | !hlock6_p & v8455ab;
assign cff2df = hlock6 & v374d7c1 | !hlock6 & v3a6224d;
assign v375129f = hmaster0_p & v3a69676 | !hmaster0_p & v3a6d897;
assign v372c5a0 = hmaster1_p & v37236b3 | !hmaster1_p & !v3777efb;
assign v372f0ee = hmaster1_p & v3a709ee | !hmaster1_p & v3728a45;
assign v3a661f8 = hmaster1_p & v373a0db | !hmaster1_p & v3765b77;
assign v3779593 = hmaster1_p & v3a635ea | !hmaster1_p & v3a6f9e6;
assign v373fa24 = hlock3_p & v373f1a5 | !hlock3_p & v3726791;
assign v37404bc = hbusreq4 & v376fb50 | !hbusreq4 & v8455ab;
assign v37500db = hmaster1_p & v37356f0 | !hmaster1_p & v37356ec;
assign v375095e = hbusreq7 & v37532f0 | !hbusreq7 & !v3a6fb8f;
assign v3723740 = hmaster2_p & v3a63777 | !hmaster2_p & v37c3782;
assign v3a70a7b = jx2_p & v3a5c317 | !jx2_p & v3a703a9;
assign v3a5fae2 = hmaster0_p & v3a7085e | !hmaster0_p & v3a7163a;
assign v375dd80 = hmaster2_p & v3a6efe8 | !hmaster2_p & v8455bf;
assign v374852b = hbusreq6_p & v37285ad | !hbusreq6_p & v3a5bb64;
assign v374d3d7 = hgrant0_p & v373dc1c | !hgrant0_p & !v8455ab;
assign v3777a9a = hbusreq4 & v3753a06 | !hbusreq4 & v3a70d99;
assign v37766f3 = hbusreq4 & v375c334 | !hbusreq4 & v2092abe;
assign v3a5e2e1 = hgrant6_p & v376e041 | !hgrant6_p & v3731004;
assign v3a704dc = hbusreq4 & v3a6f806 | !hbusreq4 & v37453d7;
assign v375fba5 = hbusreq6_p & v3749ddf | !hbusreq6_p & !v8455ab;
assign v3759749 = hbusreq0 & v3730ae3 | !hbusreq0 & v1e37cd6;
assign v3a70409 = hgrant2_p & v37721cd | !hgrant2_p & v3a6f5da;
assign v3a67f60 = hbusreq4 & v3a6dc08 | !hbusreq4 & adf78a;
assign v37237be = hbusreq2 & v373aed4 | !hbusreq2 & !v3752d10;
assign v3766664 = hlock8_p & v37458a2 | !hlock8_p & !v374f36b;
assign v3734cce = hmaster1_p & v3a635ea | !hmaster1_p & v3a56794;
assign v3a70bec = hmaster2_p & v3a5b289 | !hmaster2_p & v3a65da7;
assign v3a6ec0a = hlock4_p & v3a706d1 | !hlock4_p & v8455b7;
assign v3732f31 = hmastlock_p & v377d8f9 | !hmastlock_p & !v8455ab;
assign v3736003 = hmaster1_p & v8455e7 | !hmaster1_p & v3a6fcb2;
assign v3746824 = hbusreq0_p & v374d836 | !hbusreq0_p & v3743b9e;
assign v380954b = hgrant6_p & v3a69f9e | !hgrant6_p & v3728498;
assign v375b929 = hlock8_p & v3a70ecc | !hlock8_p & v3a6d3bc;
assign v37533ae = hlock6_p & v3730627 | !hlock6_p & v8455b7;
assign v3744aaa = hbusreq5 & v372c6c4 | !hbusreq5 & v23fde69;
assign v3743018 = hmaster0_p & v37640e9 | !hmaster0_p & v374c5c6;
assign v3a63166 = hmaster2_p & v8455ab | !hmaster2_p & v372a20c;
assign v3a6a872 = hbusreq5_p & v8455ab | !hbusreq5_p & v3a6fd62;
assign v37757cb = hbusreq5_p & v3a6e40b | !hbusreq5_p & v372c2da;
assign v3a63197 = hgrant0_p & v3736ab1 | !hgrant0_p & v373f8fb;
assign v375895e = hbusreq0 & v375c608 | !hbusreq0 & v3755744;
assign v3a6d5a8 = hmaster1_p & v376b654 | !hmaster1_p & v3768ae9;
assign v3726460 = hlock0 & v3748797 | !hlock0 & v375eeb0;
assign v3a55b5b = hlock5 & v3768d6c | !hlock5 & v373dde1;
assign v3a6fe6f = hlock5 & v37693a3 | !hlock5 & v3755aca;
assign v3734c05 = hburst0 & v8455ab | !hburst0 & v3734625;
assign v376cd0d = hmaster0_p & v374774d | !hmaster0_p & v3a64bc4;
assign v1e37943 = hmaster1_p & v8455ab | !hmaster1_p & v3725a0b;
assign v376289b = hlock6_p & v377989c | !hlock6_p & v3a6ffca;
assign v376fe90 = hmaster0_p & v8639e9 | !hmaster0_p & v3737ace;
assign v3a6a8c0 = hgrant4_p & v8455c2 | !hgrant4_p & v3771609;
assign v37507a8 = hmaster1_p & v8455ab | !hmaster1_p & !v373335b;
assign v3a670e9 = hbusreq8 & v373804d | !hbusreq8 & v3a6c81d;
assign v3774c1b = hlock0_p & v3759b2f | !hlock0_p & v3a706b0;
assign v3809eb1 = hmaster1_p & v375e037 | !hmaster1_p & v3765dbe;
assign v3a65aba = hgrant6_p & v3a5a258 | !hgrant6_p & v374b697;
assign v377504a = hmaster2_p & v3a635ea | !hmaster2_p & v3a70e98;
assign v23fda46 = jx2_p & v3a708ff | !jx2_p & v3a6261f;
assign v373a0f4 = hgrant5_p & v39a4e19 | !hgrant5_p & v38092f5;
assign v373c728 = hbusreq6 & v3a71416 | !hbusreq6 & !v8455b9;
assign v377306c = hmaster2_p & v3751b37 | !hmaster2_p & v373894d;
assign v37312e3 = hmaster2_p & v3770b26 | !hmaster2_p & v3a70f68;
assign v37590cb = hbusreq4 & v3735d39 | !hbusreq4 & v375f302;
assign v35b85ad = hbusreq5 & v3a6eb1c | !hbusreq5 & v3a6e7ed;
assign v373576f = hmaster0_p & v3740f9c | !hmaster0_p & v37276a8;
assign v3746368 = hbusreq1_p & v377051a | !hbusreq1_p & v3a6f2f2;
assign v376041f = hbusreq6 & v3a70443 | !hbusreq6 & !v8455ab;
assign v23fe142 = hmaster3_p & v372d360 | !hmaster3_p & v2ff8e61;
assign v374c6b8 = hmaster0_p & v373fd94 | !hmaster0_p & v3a6f81b;
assign v37314b5 = hlock2 & v943e48 | !hlock2 & v3a5fb00;
assign v3a68c94 = hmaster2_p & v3759b2f | !hmaster2_p & v375641f;
assign v373f4a5 = hgrant3_p & v377b6ce | !hgrant3_p & v3769157;
assign v373da5b = hgrant0_p & v97ecca | !hgrant0_p & v8455ab;
assign v23fe295 = hmaster2_p & v3771ce2 | !hmaster2_p & !v2acb5a2;
assign v3a5e5d0 = hlock0 & v374d63f | !hlock0 & v3a6b46d;
assign v37443b5 = hbusreq0 & v3759ee4 | !hbusreq0 & v3a67d4a;
assign v3769e50 = hmaster2_p & v3a635ea | !hmaster2_p & v374bb76;
assign v372eaf0 = hlock2 & v38072fd | !hlock2 & v29256ae;
assign v3a6f039 = hmaster0_p & v377bb93 | !hmaster0_p & v8455ab;
assign v377c831 = hbusreq7_p & v3a6f74f | !hbusreq7_p & !v37738b2;
assign v3757272 = hbusreq5_p & v377ee7c | !hbusreq5_p & v3a66e6f;
assign v3775064 = hbusreq5 & v377f4d5 | !hbusreq5 & v3a5d8a9;
assign v3a6ffdd = hgrant5_p & v8455ab | !hgrant5_p & v2acaeee;
assign v3a6fee1 = hgrant6_p & v37304b3 | !hgrant6_p & v374d4ca;
assign v3a6fc19 = hbusreq5_p & v376a799 | !hbusreq5_p & v375636e;
assign v373f497 = hlock8_p & v37231e5 | !hlock8_p & v375e3fd;
assign v3a62ba4 = hgrant5_p & v376a236 | !hgrant5_p & v3a70877;
assign v374d59d = hmaster0_p & v9af7ec | !hmaster0_p & v3750b01;
assign v3a70deb = hgrant5_p & v377d59e | !hgrant5_p & v3724987;
assign v3738745 = hlock4_p & v8455ab | !hlock4_p & v374a97c;
assign v3a647c6 = jx0_p & v3a62f0f | !jx0_p & v377dbdc;
assign v3a5a807 = hbusreq6_p & v373642c | !hbusreq6_p & v8455ab;
assign v3a6c96a = hgrant5_p & v8455ab | !hgrant5_p & v377fc89;
assign v3760af0 = hbusreq1_p & v37547c9 | !hbusreq1_p & !v8455ab;
assign v3a6d569 = hgrant4_p & v3774bad | !hgrant4_p & v3763b0a;
assign v374a9a0 = hbusreq6 & v373a452 | !hbusreq6 & v8455ab;
assign v3809a76 = hgrant3_p & v3a615f7 | !hgrant3_p & v3a71682;
assign v374bab6 = hmaster2_p & v380760a | !hmaster2_p & v3769ba9;
assign v37315a3 = hmaster0_p & v374190f | !hmaster0_p & v3a58b9f;
assign v3a58c79 = hbusreq0_p & ad2d05 | !hbusreq0_p & v377ce66;
assign v3a6e124 = hbusreq5_p & v375888e | !hbusreq5_p & v3a6f5b3;
assign v3a6988c = hbusreq5_p & v3a5d522 | !hbusreq5_p & v3731b41;
assign v3a71241 = jx1_p & v89e294 | !jx1_p & v38076b3;
assign v37559b2 = hmaster0_p & v8455ab | !hmaster0_p & v3a6e432;
assign v3773eee = hmaster0_p & v3a6f443 | !hmaster0_p & v376eaf2;
assign v3739493 = hgrant5_p & v375e035 | !hgrant5_p & v377cf34;
assign v3756465 = hbusreq3 & v3a6f018 | !hbusreq3 & !v3740f3d;
assign v3a6fdd0 = hbusreq3_p & v3778765 | !hbusreq3_p & v3a6a867;
assign v377bcb3 = hmaster0_p & v3a625b1 | !hmaster0_p & v3742cd4;
assign v3766b11 = hbusreq2 & v3770651 | !hbusreq2 & v373c924;
assign v377c2ff = hmaster1_p & v3a66aa4 | !hmaster1_p & v3a71608;
assign v3a67cfe = hbusreq4 & v37307dd | !hbusreq4 & v8455b3;
assign v3a691eb = hgrant4_p & v8455ab | !hgrant4_p & v373abde;
assign v373891b = hgrant4_p & v35b774b | !hgrant4_p & v372cc0a;
assign v3754c5e = hgrant6_p & v3a64e05 | !hgrant6_p & v37401f0;
assign v3756a9e = hmaster2_p & v8455bb | !hmaster2_p & v3a5e7fe;
assign v377b6ce = locked_p & v8455ab | !locked_p & !v35772a6;
assign v3a6fa7e = hbusreq6 & v3740839 | !hbusreq6 & v3748797;
assign v377a968 = hmaster0_p & v8455ab | !hmaster0_p & !v3767631;
assign v3378f5d = hmaster0_p & v3a6bef4 | !hmaster0_p & !v3734b20;
assign v373016b = hbusreq5_p & v3a6b931 | !hbusreq5_p & v377b429;
assign v3a54c77 = hready & v3732eca | !hready & v373fe5e;
assign v375c9ea = hbusreq6 & v3a6006a | !hbusreq6 & v3a7162d;
assign v3a6f911 = hlock7 & v375fda5 | !hlock7 & v377619b;
assign v3744142 = hbusreq6_p & v374513e | !hbusreq6_p & !v37392ad;
assign v3724b5a = hbusreq5_p & v3a5bbbb | !hbusreq5_p & v8455ab;
assign v37237cd = hlock4 & v377e2ae | !hlock4 & v3754422;
assign v3753d9d = hbusreq0 & v376d7c6 | !hbusreq0 & v375bdaf;
assign d138a6 = hbusreq2_p & v37790a9 | !hbusreq2_p & v3756ca5;
assign v3a662f7 = hburst1 & v3a563ad | !hburst1 & v3774ad3;
assign v376a1a3 = hgrant6_p & v3741b28 | !hgrant6_p & v37569ec;
assign v375c924 = hbusreq7 & v3a70f92 | !hbusreq7 & v373c26c;
assign v3737e2e = hmaster2_p & v375501e | !hmaster2_p & v3760513;
assign v325b591 = hbusreq2_p & v3a5e7fe | !hbusreq2_p & !v8455ab;
assign v3775903 = hgrant5_p & v372aaf8 | !hgrant5_p & v3752f8e;
assign v374361e = hmaster1_p & v377b253 | !hmaster1_p & v3762a54;
assign v377d107 = hbusreq4_p & v373014d | !hbusreq4_p & v3a710c1;
assign v377414c = hbusreq4 & v37556ec | !hbusreq4 & v3765e79;
assign v377e0c6 = hbusreq5 & v3a67471 | !hbusreq5 & v8455ab;
assign v3730fbd = hbusreq5 & v3a6a6e1 | !hbusreq5 & v3a7129c;
assign v3a6f33e = hbusreq5_p & v3778ac2 | !hbusreq5_p & v23fd84e;
assign v3742953 = hbusreq0 & v375f98a | !hbusreq0 & v8455ab;
assign v38074aa = hgrant5_p & v8455ab | !hgrant5_p & ad41f9;
assign v3a6f7bf = hbusreq1_p & v3740171 | !hbusreq1_p & v37457fb;
assign v3a66668 = hgrant3_p & v8455ab | !hgrant3_p & !v3768b81;
assign v377a236 = hmaster2_p & v3a6f081 | !hmaster2_p & !v3a7153c;
assign v3738b0c = hbusreq3_p & v3a65cfb | !hbusreq3_p & v8455ab;
assign v375d512 = jx0_p & v3a55cf3 | !jx0_p & v3749535;
assign v3741872 = hmaster1_p & v377c261 | !hmaster1_p & v3a5fd18;
assign v3a703cc = hbusreq0_p & v373e67e | !hbusreq0_p & v8455ab;
assign v373e296 = hlock3 & v376485c | !hlock3 & v37567c7;
assign v3807315 = hbusreq6 & v3a70200 | !hbusreq6 & !v3a5538a;
assign v3737ab4 = jx1_p & v3808cf5 | !jx1_p & v8455ab;
assign v3754e8e = hmaster0_p & v37312e3 | !hmaster0_p & v37565b0;
assign v372b893 = hgrant6_p & v8455ab | !hgrant6_p & v3752b6a;
assign v3739914 = hlock5 & v377c307 | !hlock5 & v376b290;
assign cf6441 = hlock3 & v3809865 | !hlock3 & v3750e9a;
assign v3a6799d = hbusreq5 & a14297 | !hbusreq5 & v3a7005b;
assign v3724b78 = hmaster1_p & v3735e84 | !hmaster1_p & v3755aae;
assign v37581c2 = hgrant6_p & v377f21b | !hgrant6_p & v3a705db;
assign v37584c7 = hgrant6_p & v3a5e24e | !hgrant6_p & v372dcc2;
assign v3a5ceaf = hbusreq5_p & v3a624ec | !hbusreq5_p & !v3745a3b;
assign v3a7039b = hbusreq6 & v373fe5e | !hbusreq6 & v8455e7;
assign v3a70760 = hbusreq8 & v8455e7 | !hbusreq8 & v3739f49;
assign v3771b83 = hmaster2_p & v8455ab | !hmaster2_p & v372e559;
assign v372ed51 = hbusreq1_p & v377e85e | !hbusreq1_p & v8455ab;
assign v37715af = hbusreq6 & v3a68967 | !hbusreq6 & v3a6da8a;
assign v3a2a0f4 = hmaster0_p & v3a633b9 | !hmaster0_p & v23fe28c;
assign v37356aa = hmaster1_p & v376fe45 | !hmaster1_p & v375548b;
assign v37780fd = hmaster2_p & v3a6f443 | !hmaster2_p & v3a6d684;
assign v3a6f3f5 = hmaster2_p & v3a6f92f | !hmaster2_p & !v39a4dbb;
assign v3a60258 = hgrant6_p & v8455c9 | !hgrant6_p & v3768d47;
assign v3a6f496 = hbusreq2_p & v376d1e2 | !hbusreq2_p & v37348ee;
assign v374d4ae = hmaster2_p & v8455bf | !hmaster2_p & !v374b25d;
assign v375d2b1 = hlock7 & v375c924 | !hlock7 & v3a70f92;
assign v3765eee = hbusreq0 & v3a66306 | !hbusreq0 & v37675d5;
assign v3773f27 = hmaster1_p & v3a635ea | !hmaster1_p & v3a6d4f3;
assign v3a60147 = hmaster2_p & v3a6fc9c | !hmaster2_p & v8455ab;
assign v3733664 = hgrant5_p & v3726088 | !hgrant5_p & v3a6f593;
assign v3739774 = hmaster2_p & be54b2 | !hmaster2_p & v3769740;
assign v3a6fb9d = hlock2 & v38072fd | !hlock2 & v3a63a2a;
assign v3739c89 = hbusreq8 & v3778f25 | !hbusreq8 & v376ae9f;
assign v376fa43 = hmaster0_p & v3723dc3 | !hmaster0_p & v3a6e93d;
assign v3769e70 = hlock4 & v3773e77 | !hlock4 & v3752933;
assign v3a5bbeb = hlock4 & v3766727 | !hlock4 & v3a71540;
assign v376a166 = hbusreq6 & v3761362 | !hbusreq6 & v8455ab;
assign v372648f = hbusreq8_p & v3746045 | !hbusreq8_p & v3777995;
assign v3a6f406 = hmaster2_p & v375af43 | !hmaster2_p & v3a67905;
assign v37347cd = hbusreq8 & v3769a16 | !hbusreq8 & v377a27f;
assign v3a70fc0 = hbusreq1_p & v376e00a | !hbusreq1_p & v8455b6;
assign v37571fc = hbusreq7_p & v3763a29 | !hbusreq7_p & v373fd58;
assign v377b209 = hbusreq8_p & v9c8578 | !hbusreq8_p & v376b744;
assign v376eb1f = hbusreq6 & v373f79d | !hbusreq6 & v8455ab;
assign v3773aa9 = hgrant0_p & v8455ab | !hgrant0_p & v3771bb9;
assign v3a6f8b7 = hgrant5_p & v3a6f73f | !hgrant5_p & v3a6f2b7;
assign v372b8fd = hbusreq0 & v3a57ac7 | !hbusreq0 & v374b6ac;
assign v3a56e45 = hbusreq7 & v3758e8d | !hbusreq7 & v3a6f259;
assign v37744e3 = jx1_p & v3a70907 | !jx1_p & v3770362;
assign v374dfe1 = hmaster0_p & v3742dac | !hmaster0_p & v3757ffa;
assign v38068c1 = hmaster1_p & v3a6f327 | !hmaster1_p & !v372fbb1;
assign v3a702de = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a6fc9b;
assign v3a54c12 = hbusreq6_p & v3a64d23 | !hbusreq6_p & v372ef40;
assign v375d288 = hbusreq0_p & v374f307 | !hbusreq0_p & v8455ab;
assign v3a70194 = hmaster1_p & v8455ab | !hmaster1_p & !v3a6f2c6;
assign v38099e8 = hlock3 & v3a6b8a2 | !hlock3 & v23fe0bb;
assign v3a57325 = hlock6_p & v37521ed | !hlock6_p & !v8455ab;
assign v380917f = hlock2 & v2092b23 | !hlock2 & v37415b2;
assign v3757519 = hbusreq8_p & v37647de | !hbusreq8_p & v3761431;
assign v3a6692b = hlock5_p & v37702f3 | !hlock5_p & !v37394b7;
assign v3a70623 = hmaster1_p & v37570f8 | !hmaster1_p & v373d5e7;
assign v3378d8f = hgrant6_p & v39ea76e | !hgrant6_p & v375c265;
assign dacf90 = hbusreq7_p & v37431c0 | !hbusreq7_p & v3a68931;
assign v37233a2 = hmaster2_p & v3a68793 | !hmaster2_p & v3a6039a;
assign v3a70765 = hlock4 & v374e436 | !hlock4 & v373de13;
assign v376c79a = hmaster0_p & v380913f | !hmaster0_p & v376d21d;
assign v3a6b303 = hmaster1_p & v3a68356 | !hmaster1_p & v8455ab;
assign v375a269 = hlock5_p & v23fdadd | !hlock5_p & v3a6abcb;
assign v3a6fec4 = hmaster2_p & v3735fca | !hmaster2_p & v375693b;
assign v3a55cda = hmaster0_p & afdeb4 | !hmaster0_p & v3768495;
assign v372b4c0 = hgrant6_p & v3a62b8d | !hgrant6_p & v3769a36;
assign v3a6f567 = hlock6 & v375534a | !hlock6 & v37642a0;
assign v3735bef = hmaster1_p & v3a71678 | !hmaster1_p & v3767efa;
assign v375c5a8 = hbusreq1_p & v3756bc9 | !hbusreq1_p & v3a6d684;
assign v3a6f6ea = hmaster0_p & v3754ee0 | !hmaster0_p & v3a7026a;
assign v3377c6a = hbusreq4_p & v3740e5a | !hbusreq4_p & v3744dca;
assign v3a556df = hmaster0_p & v8455b0 | !hmaster0_p & v3a6f40d;
assign v8955d0 = hbusreq4_p & v3a66123 | !hbusreq4_p & v372b893;
assign v374a7f2 = hbusreq8 & v3759663 | !hbusreq8 & v3a56918;
assign v37465c7 = hbusreq5_p & v376497a | !hbusreq5_p & !v8455ab;
assign v3a619b8 = hbusreq5 & v3a6fd4e | !hbusreq5 & v3a69ead;
assign v373a415 = hbusreq0 & v3747994 | !hbusreq0 & v8455ab;
assign v3a70ded = hmaster2_p & v8455ab | !hmaster2_p & v3744a0c;
assign v23fe10f = hbusreq6_p & v3748fba | !hbusreq6_p & v377b5c4;
assign v376e0b6 = hmaster0_p & v3a6fe09 | !hmaster0_p & v37315d0;
assign v3a63dbb = hbusreq6_p & adf78a | !hbusreq6_p & v3753dab;
assign v3a67c6d = hgrant5_p & v372e53f | !hgrant5_p & v3753c8c;
assign v3a66811 = hbusreq5_p & v3a70c6c | !hbusreq5_p & cf8423;
assign v3768ae9 = hbusreq5_p & v3755e64 | !hbusreq5_p & !v372b652;
assign v39a4ed6 = hgrant6_p & v8455ab | !hgrant6_p & v374177f;
assign v3735525 = hlock0_p & v375da10 | !hlock0_p & v375588c;
assign v3768bbc = hgrant4_p & v3a6f64e | !hgrant4_p & v3a56b19;
assign v3a6f252 = locked_p & v3a6ef8c | !locked_p & v37566b2;
assign v3724ff0 = hlock5_p & v3a5f9d5 | !hlock5_p & !v3a6fbac;
assign v372d203 = hbusreq3_p & v3a6320d | !hbusreq3_p & v8455ab;
assign v372d748 = hbusreq5_p & v3a6d7cd | !hbusreq5_p & v3a6fb03;
assign v3770aa1 = hmaster0_p & v37645eb | !hmaster0_p & v374953c;
assign v374e92a = hmaster0_p & v377ce1a | !hmaster0_p & v3767e7e;
assign v3727e58 = hmaster2_p & v37696b6 | !hmaster2_p & v375f9df;
assign v375facd = jx0_p & v3a6faed | !jx0_p & v3772e3f;
assign v3a53392 = hgrant5_p & v3a700be | !hgrant5_p & v3765b5c;
assign v3737e2d = hgrant4_p & v3754cf4 | !hgrant4_p & v37704dc;
assign v373e369 = hgrant3_p & v3755b5e | !hgrant3_p & v3a708af;
assign v3a6c0b3 = hlock1 & v3753a3f | !hlock1 & v3778528;
assign v3a57309 = hready & v37386f2 | !hready & v3730cce;
assign v3a5f4ef = hbusreq8_p & v374445b | !hbusreq8_p & v3a70d92;
assign v37759b5 = hbusreq4 & v372cb44 | !hbusreq4 & v3a620d3;
assign v3760ba3 = hbusreq4_p & v3a601a0 | !hbusreq4_p & v375d5ac;
assign c22b44 = hlock3_p & v372c565 | !hlock3_p & v377bdbe;
assign v3749ea2 = hlock3_p & v8455ab | !hlock3_p & v3a5d923;
assign v3a6f459 = jx2_p & v3a6f619 | !jx2_p & v3747d51;
assign v373b0f3 = hbusreq7 & v3772a57 | !hbusreq7 & v3a63ac4;
assign v3a5cfdb = hbusreq1_p & d0a687 | !hbusreq1_p & v8455ab;
assign v372ab70 = hgrant5_p & v8455c6 | !hgrant5_p & v3a70247;
assign v3a703cf = stateA1_p & v3732f31 | !stateA1_p & v372dee5;
assign v3a538b4 = hbusreq6_p & v3769ae2 | !hbusreq6_p & v3a6de90;
assign v3724b74 = hmaster0_p & v37665c5 | !hmaster0_p & v3768c25;
assign v3769ae2 = hbusreq1_p & v3a625ee | !hbusreq1_p & v8455ab;
assign v37747a9 = hbusreq4 & v3729f25 | !hbusreq4 & !v8455ab;
assign v373d7f9 = hbusreq0 & v3a70a2a | !hbusreq0 & v3727347;
assign v3a5c462 = hgrant6_p & v3775293 | !hgrant6_p & v3738602;
assign v3a61f9b = hlock4_p & v3a617b4 | !hlock4_p & v3767437;
assign v3778628 = hbusreq5_p & v3766b26 | !hbusreq5_p & v3731fd2;
assign v3a539ee = stateA1_p & v373c3bd | !stateA1_p & v8455ab;
assign v374ef8d = jx1_p & v8455ab | !jx1_p & v37501a3;
assign v37250fa = hbusreq4 & v3735ea8 | !hbusreq4 & v372cc0a;
assign v376a0e3 = hmaster2_p & v8455ab | !hmaster2_p & !v3a71617;
assign v375d661 = hmaster1_p & v3a556f8 | !hmaster1_p & v37330ca;
assign v374f106 = hlock0_p & v8455ab | !hlock0_p & v3a6f522;
assign v374c6b1 = hbusreq2_p & v376f56d | !hbusreq2_p & v3748c34;
assign v3a7064c = hlock7_p & v37244f3 | !hlock7_p & a792d5;
assign v37625ef = hbusreq0 & v3a60c49 | !hbusreq0 & v3a70d38;
assign v3808db4 = hbusreq8 & v3753ee8 | !hbusreq8 & v3806a1c;
assign v377d8d6 = hlock4_p & v373d825 | !hlock4_p & !v8455ab;
assign v3754237 = hbusreq6 & v37302f1 | !hbusreq6 & !v8455bd;
assign v360bb9f = hbusreq0_p & v375de18 | !hbusreq0_p & !v37282cf;
assign v377190a = hgrant4_p & v37780cc | !hgrant4_p & v8455ab;
assign v377d1ab = hbusreq4 & v37302c5 | !hbusreq4 & v3a6efad;
assign v3a70363 = hbusreq4_p & v3724f5d | !hbusreq4_p & v375a32c;
assign v373de83 = hbusreq8_p & v3808eb8 | !hbusreq8_p & v3770338;
assign v3772d27 = hlock3_p & v3a6f9a8 | !hlock3_p & v374720c;
assign v376ea59 = hmaster2_p & v372c3df | !hmaster2_p & v8455ab;
assign v3a63777 = hbusreq6_p & v3a69de7 | !hbusreq6_p & v3a635ea;
assign v377bbfc = hbusreq8_p & v375c24b | !hbusreq8_p & v374803b;
assign v372a25a = jx0_p & v3a680cd | !jx0_p & v375c525;
assign v373e70e = hmaster0_p & v3a6f3d8 | !hmaster0_p & v3777f6e;
assign v3a59ed6 = hmaster2_p & v372455c | !hmaster2_p & !v376fcc3;
assign v3a5e909 = hlock0 & v377bfc0 | !hlock0 & v375370a;
assign v37728cd = hmaster1_p & v38087e5 | !hmaster1_p & v8a7af6;
assign v3a6f331 = hgrant2_p & v374e5ac | !hgrant2_p & v3733a19;
assign v3a6c09f = hmaster0_p & v3a71195 | !hmaster0_p & v3a6b73c;
assign v3742c6c = hbusreq0 & v37366ed | !hbusreq0 & v37671eb;
assign v3a702b3 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3739bcb;
assign v3a71145 = hbusreq3_p & v3a635ea | !hbusreq3_p & v376bade;
assign v373c423 = hbusreq6_p & v375dc46 | !hbusreq6_p & v37627f9;
assign v3a5eb63 = hgrant5_p & v3a6f07b | !hgrant5_p & v372c09a;
assign v3a70966 = hgrant6_p & v374510e | !hgrant6_p & v373b10f;
assign v37495dc = hbusreq2_p & v3a635ea | !hbusreq2_p & v373081f;
assign v3a6f9c3 = hlock3_p & v373aaa8 | !hlock3_p & !v8455ab;
assign v3a6feca = hlock6_p & v3806f67 | !hlock6_p & v8455ab;
assign v3723635 = hgrant6_p & v8455ab | !hgrant6_p & v3a6f377;
assign v3808ee4 = hgrant2_p & v3742c52 | !hgrant2_p & v375d1fa;
assign v3a70cf6 = hbusreq5 & v373fa8c | !hbusreq5 & v8455b5;
assign v3a6e3d1 = hlock2_p & v377e090 | !hlock2_p & v3761224;
assign v3773f2b = hmaster0_p & v3a5c6d0 | !hmaster0_p & v3769d48;
assign v9f823e = hgrant4_p & v3723430 | !hgrant4_p & v37bfc8c;
assign v377bb56 = hgrant2_p & v8455ab | !hgrant2_p & v377f669;
assign v3774730 = hmaster2_p & baec07 | !hmaster2_p & v8455ab;
assign v3a5b98b = hbusreq5_p & v377cf4f | !hbusreq5_p & v3730145;
assign v373dee0 = hlock7_p & v375e04e | !hlock7_p & v3760a6e;
assign v3728e25 = hbusreq2 & v3a70799 | !hbusreq2 & v8455ab;
assign v3729238 = hmaster0_p & v2092f0f | !hmaster0_p & v375d507;
assign v37509fc = hbusreq5_p & v3a6c5e5 | !hbusreq5_p & v3772200;
assign v375153e = hlock4_p & v372d203 | !hlock4_p & v8455b0;
assign v3a70981 = hbusreq8 & v374350d | !hbusreq8 & v3a6f76b;
assign v372aefc = hlock6 & v373e789 | !hlock6 & v3a705dd;
assign v37440af = hmaster0_p & v37386f5 | !hmaster0_p & v375f87b;
assign v3a5d40d = hbusreq4 & v372936a | !hbusreq4 & v8455ab;
assign v3a705f6 = busreq_p & v376147f | !busreq_p & v374057a;
assign v3744934 = hbusreq4_p & v3755f9b | !hbusreq4_p & !v3a67142;
assign v3757100 = hbusreq5_p & v3735e84 | !hbusreq5_p & v3a715c1;
assign v3a5c653 = hmaster1_p & v37398ac | !hmaster1_p & v373db68;
assign v3a71592 = jx0_p & v3a7041c | !jx0_p & v3752091;
assign v3a6051e = hgrant5_p & v376e66e | !hgrant5_p & v374143e;
assign v3730a73 = hmaster0_p & v3a5c945 | !hmaster0_p & v3a703db;
assign v37625b7 = hlock0_p & v3751b0e | !hlock0_p & v376da28;
assign v3a5a04c = hgrant4_p & v373b295 | !hgrant4_p & !v3a6f6d3;
assign v3733e5a = hmaster1_p & v37249c7 | !hmaster1_p & v3a70516;
assign v3a713b5 = hbusreq5 & v373fa48 | !hbusreq5 & v3a5cb2c;
assign v37339f0 = hbusreq0_p & v3747302 | !hbusreq0_p & v37416b5;
assign v37525c5 = jx0_p & v3a70213 | !jx0_p & v3775622;
assign v3a6b22e = hbusreq7_p & v37387e6 | !hbusreq7_p & v372b7b1;
assign v37318da = hbusreq2 & v37366d0 | !hbusreq2 & v8455ab;
assign v38068b5 = hbusreq2_p & v3a5cc4c | !hbusreq2_p & v37780f6;
assign v374f094 = hmaster1_p & v373e376 | !hmaster1_p & v3a7051d;
assign v3761fd6 = hmaster2_p & v377e089 | !hmaster2_p & v3755dcd;
assign v374217a = hbusreq4 & v3a6dfc9 | !hbusreq4 & v3a70b92;
assign v3a702f0 = hmaster1_p & v3a707ee | !hmaster1_p & v37261b3;
assign v2092c08 = decide_p & v3750012 | !decide_p & v3a5d2f1;
assign v3729385 = jx1_p & v377dadb | !jx1_p & v3a5eecb;
assign c536d5 = hmaster2_p & v376b11a | !hmaster2_p & v3a6910c;
assign v374a543 = hbusreq8 & v3731455 | !hbusreq8 & v3779f0a;
assign v3743057 = hmaster1_p & v3766298 | !hmaster1_p & v3729988;
assign v376110e = hlock6_p & v3a637dd | !hlock6_p & !v8455ab;
assign v3730d6b = hmaster0_p & v3772327 | !hmaster0_p & !v375f664;
assign v377ae0c = hbusreq7 & v3a64ba3 | !hbusreq7 & v3a64293;
assign v3731455 = hlock7 & v3765442 | !hlock7 & v3773a06;
assign v3a71429 = hgrant6_p & v3a5cb5f | !hgrant6_p & v375d707;
assign v3a664b5 = hmaster2_p & v375a1ab | !hmaster2_p & v2ff937f;
assign v3774937 = hmaster0_p & v3755b07 | !hmaster0_p & v3760f64;
assign v3737897 = hbusreq7 & v3a70b26 | !hbusreq7 & v377b735;
assign v3748870 = hgrant2_p & v3a70303 | !hgrant2_p & v3a655a3;
assign v375abaa = hgrant5_p & v3747465 | !hgrant5_p & v3732b3a;
assign v3a548c2 = hmaster2_p & v3a6d684 | !hmaster2_p & v376ea4a;
assign v3a60c49 = hlock4 & v375a92b | !hlock4 & v374178a;
assign v3735aa5 = hmaster1_p & v3a66110 | !hmaster1_p & v3a6f54e;
assign v37796e9 = hbusreq5 & v3a705ba | !hbusreq5 & v8455ab;
assign v2925d03 = hmaster0_p & v3800eea | !hmaster0_p & v3a6f81b;
assign v372d35f = hmaster0_p & v37706e9 | !hmaster0_p & v3776c95;
assign v377aacd = hlock3_p & v376a936 | !hlock3_p & v3a5e91b;
assign v3740083 = hlock0_p & v372391f | !hlock0_p & v37269a2;
assign b539d9 = hmaster3_p & v37597f7 | !hmaster3_p & v3a6f261;
assign v3735859 = hbusreq5_p & v376eed1 | !hbusreq5_p & v376bc8c;
assign v374f3ad = hmaster0_p & v3a635ea | !hmaster0_p & v3a70a6e;
assign v3a55b2d = hlock3 & v377665f | !hlock3 & v37438c9;
assign v373ae2e = hgrant1_p & v376e914 | !hgrant1_p & !v35772a6;
assign v3764aea = hbusreq3_p & v375f462 | !hbusreq3_p & v3747cf5;
assign v3742995 = hgrant4_p & v8455e7 | !hgrant4_p & !v3a5af5c;
assign v37364d2 = hbusreq4_p & v3a6f647 | !hbusreq4_p & v373f8a7;
assign v372c480 = hbusreq4 & v3a6f571 | !hbusreq4 & v3731a5a;
assign v3a7000e = hbusreq3_p & v3a7032d | !hbusreq3_p & v3a70a3c;
assign v3736028 = hlock0_p & v3a635ea | !hlock0_p & !v3a6f1f8;
assign v3744399 = hbusreq5_p & v8455cb | !hbusreq5_p & v3a709fc;
assign v3751cd1 = hbusreq0 & v3a64ca0 | !hbusreq0 & v3a702e5;
assign v375cb51 = hmaster2_p & v377b946 | !hmaster2_p & v374d0e3;
assign v373324d = hmaster0_p & v37435a9 | !hmaster0_p & v375fe03;
assign v37494bb = hbusreq6 & v375dc46 | !hbusreq6 & v3a5b91d;
assign v375d1d9 = hgrant6_p & v372bfa1 | !hgrant6_p & v377ee3c;
assign v37415e4 = jx0_p & v374c885 | !jx0_p & v33790c9;
assign v3768a57 = hgrant6_p & v3a69f9e | !hgrant6_p & v372d1bf;
assign v3769112 = hlock6 & v3768d29 | !hlock6 & v3a56608;
assign v37282ac = hbusreq6_p & v3725bf4 | !hbusreq6_p & v8455ab;
assign v3a701f7 = hlock7 & v3a555a9 | !hlock7 & v3807413;
assign v3766260 = hlock7_p & v3a70367 | !hlock7_p & v3736dfe;
assign v37691d1 = hmaster0_p & v372673d | !hmaster0_p & v373a16b;
assign v37484e0 = hbusreq2_p & v377097a | !hbusreq2_p & v3a62a6d;
assign v377dabc = hgrant3_p & v372ec1c | !hgrant3_p & v3774e8c;
assign v3774a95 = hgrant4_p & v8455b5 | !hgrant4_p & v377e933;
assign v3a62e20 = hgrant5_p & v3a70a54 | !hgrant5_p & v380732c;
assign v3734f70 = hbusreq6 & v3a6f77e | !hbusreq6 & v38072fd;
assign v3a7062d = hmaster2_p & v3a6da5a | !hmaster2_p & v37406e8;
assign v3723501 = hgrant4_p & v3a5f162 | !hgrant4_p & v3a70c5d;
assign v376f455 = stateG10_1_p & v8455e7 | !stateG10_1_p & !v337904e;
assign v3a65335 = jx0_p & v3747b30 | !jx0_p & !v37730df;
assign v3a67905 = hbusreq0 & v37269f4 | !hbusreq0 & v8455ab;
assign v37d8c61 = hbusreq5 & v37454c6 | !hbusreq5 & v3770ea8;
assign v3a606b7 = hmaster2_p & v8455b0 | !hmaster2_p & v3a621cb;
assign v3a5f992 = hmaster2_p & v3729c45 | !hmaster2_p & v372de1e;
assign v3748cd9 = hbusreq5 & v3769f4e | !hbusreq5 & v375e037;
assign v37392e2 = hbusreq5 & v372c6c4 | !hbusreq5 & v3a617a2;
assign v1e37e67 = hbusreq4 & v375cfa5 | !hbusreq4 & v375da82;
assign v37475d9 = hmaster0_p & v376b015 | !hmaster0_p & v3a714d5;
assign v3739e4f = hbusreq8 & v3a6f911 | !hbusreq8 & v376eeb3;
assign v3759be3 = hlock5 & v377fc51 | !hlock5 & v374e843;
assign v37752c8 = hbusreq4 & v3a711e2 | !hbusreq4 & v3756eca;
assign v374f0e7 = hlock3_p & v3724418 | !hlock3_p & v8455b3;
assign v37520db = hbusreq2 & v37282cf | !hbusreq2 & v37674c1;
assign v3727db5 = hgrant4_p & v375c7b9 | !hgrant4_p & v3a29dbd;
assign v372ee98 = hgrant4_p & v374ad81 | !hgrant4_p & !v375b3f0;
assign v375c6cd = hlock7_p & v374704e | !hlock7_p & v3a689d1;
assign v3a5f9ad = hgrant3_p & v372d02d | !hgrant3_p & v3726f97;
assign v377b4c9 = hbusreq0 & v3726229 | !hbusreq0 & !v3733278;
assign v3a70fec = hbusreq4_p & v37404bc | !hbusreq4_p & v8455ab;
assign v3723baf = hbusreq6 & v3a56d0a | !hbusreq6 & v3a6a116;
assign v3747ec5 = hgrant2_p & v8455ab | !hgrant2_p & v3776ca8;
assign v3742121 = hmaster2_p & v3769ae2 | !hmaster2_p & v374f96e;
assign v37611f5 = hbusreq7 & v3a6373e | !hbusreq7 & v8455ab;
assign v3a5ff26 = hmaster2_p & v8455e7 | !hmaster2_p & !v376653d;
assign v37c02a0 = hbusreq2 & adf78a | !hbusreq2 & v3730ffe;
assign v3735d39 = hlock6 & v372e798 | !hlock6 & v3a702bc;
assign v3768a78 = hmaster2_p & v3731b41 | !hmaster2_p & v373b30b;
assign v373f042 = hmaster0_p & v374176c | !hmaster0_p & v8455e7;
assign v3755381 = hbusreq3 & v8455b0 | !hbusreq3 & v3a63805;
assign v2092abe = hbusreq6_p & v8455bf | !hbusreq6_p & v3a6da8a;
assign v376e7bc = hbusreq3_p & v3733e9e | !hbusreq3_p & v1e38224;
assign v373376b = hgrant2_p & v3a56187 | !hgrant2_p & v3768b07;
assign v3a7017d = hmaster0_p & v376ddb6 | !hmaster0_p & v373c3a0;
assign v374ad5f = hlock5_p & v377f2ec | !hlock5_p & v375d1d1;
assign v3a7047c = hgrant4_p & v376a6f1 | !hgrant4_p & v3729e38;
assign v3a5ff81 = stateG2_p & v8455ab | !stateG2_p & v3745b52;
assign v3a594fe = hmaster2_p & v3a635ea | !hmaster2_p & v2ff8bbc;
assign v3a58200 = hbusreq4_p & v3749bf0 | !hbusreq4_p & v3a6bb84;
assign v38064e3 = hbusreq5_p & v3731e50 | !hbusreq5_p & v3a712e9;
assign v3a54ebe = hmaster0_p & v377d107 | !hmaster0_p & v3776914;
assign v373875c = hmaster1_p & v377233c | !hmaster1_p & v3a6da41;
assign v3764c6c = hgrant5_p & v375bf12 | !hgrant5_p & v2ff9397;
assign v373a141 = hbusreq0 & v3a59d65 | !hbusreq0 & v3a67e53;
assign v3774f39 = hmaster1_p & v376c79a | !hmaster1_p & v3a53fb5;
assign v3730789 = hmaster2_p & v3a57384 | !hmaster2_p & v3a707ce;
assign v37354bf = hmaster3_p & v373fe61 | !hmaster3_p & v3a55078;
assign v3a66da0 = hbusreq8 & v377d904 | !hbusreq8 & v8455ab;
assign v3a62a96 = hbusreq3_p & v3a6f9c3 | !hbusreq3_p & !v8455ab;
assign v374270d = hgrant1_p & v375eb78 | !hgrant1_p & v37270d9;
assign v3a58773 = hbusreq0 & v3a702b0 | !hbusreq0 & v8455ab;
assign v374ba57 = hbusreq5_p & v3a6d1ea | !hbusreq5_p & v1e373f8;
assign v3a654fb = hlock2_p & v3a70dcd | !hlock2_p & v3a61a3d;
assign v3a5fa18 = hgrant0_p & v3753e6a | !hgrant0_p & v37356ce;
assign v3a53d04 = hmaster1_p & v37237f1 | !hmaster1_p & v377f264;
assign v3755000 = hgrant4_p & v1e37b99 | !hgrant4_p & !v3755ad5;
assign v3775537 = hbusreq2_p & v3a70d2c | !hbusreq2_p & v8455ab;
assign v3a700d0 = hmaster3_p & v37377f0 | !hmaster3_p & v3a6aa8d;
assign v3a659e5 = hmaster2_p & v3a701c4 | !hmaster2_p & v375444a;
assign v376102a = hlock0_p & v374e35e | !hlock0_p & v376f9d9;
assign dbf06b = hbusreq8 & v3a70819 | !hbusreq8 & v3a60859;
assign v3731cc6 = hmaster1_p & v374502e | !hmaster1_p & c7885c;
assign v3a70cac = hbusreq8 & v23fe312 | !hbusreq8 & v3746b0c;
assign v374143e = hmaster1_p & v3a5e2a3 | !hmaster1_p & v373d3e5;
assign v3755417 = hbusreq4_p & v3732c72 | !hbusreq4_p & v374a86a;
assign v3730d18 = hmaster2_p & v3777311 | !hmaster2_p & v8455ab;
assign v37396de = hbusreq0 & v377bbbd | !hbusreq0 & v3745b60;
assign v3a6f7a1 = hbusreq4_p & v3729e0b | !hbusreq4_p & !v3a70b37;
assign v3a7008c = hgrant2_p & v376495e | !hgrant2_p & v3a703ad;
assign v37793a6 = hmaster2_p & v373f058 | !hmaster2_p & v3a704e5;
assign ce419c = hgrant2_p & v3577306 | !hgrant2_p & ab60dc;
assign v3a6eeb9 = hbusreq7 & v374daa9 | !hbusreq7 & v37258d6;
assign v3774710 = hbusreq3 & v373b7c8 | !hbusreq3 & v8455ab;
assign v3a65ee0 = hmaster0_p & v3a55b91 | !hmaster0_p & !v3a56512;
assign v3732b30 = hbusreq7 & v3779e9b | !hbusreq7 & v3723025;
assign v3a70ff8 = hgrant4_p & v8455ab | !hgrant4_p & v377c41b;
assign v3735ed0 = stateA1_p & v3a6a939 | !stateA1_p & v8455ab;
assign v3731a2e = hbusreq8_p & v372543f | !hbusreq8_p & v3a7011b;
assign v3756304 = hbusreq0 & v374b37d | !hbusreq0 & v372946e;
assign v373d62b = hbusreq2_p & v373449a | !hbusreq2_p & v3a703e0;
assign v37239a5 = hmaster1_p & v375df5a | !hmaster1_p & v3761bd6;
assign v37703c6 = hbusreq0_p & v375323b | !hbusreq0_p & v8455ab;
assign v3a71374 = hmaster2_p & v374c78e | !hmaster2_p & b68bf2;
assign v374679f = hbusreq0 & v3755f4a | !hbusreq0 & v372f570;
assign v3726865 = hgrant6_p & v8455c9 | !hgrant6_p & da4c01;
assign v37787da = hlock0 & v3a60a68 | !hlock0 & v3735e89;
assign v3a700ee = hmaster0_p & v376f0ab | !hmaster0_p & v3764015;
assign v3a700e8 = hmaster3_p & v3a647cd | !hmaster3_p & v3a5af41;
assign v376029a = hbusreq4_p & adf78a | !hbusreq4_p & v3753dab;
assign v3747b3c = hgrant6_p & v8455ab | !hgrant6_p & v373a5b6;
assign v3778355 = hbusreq4 & v3a5a01b | !hbusreq4 & v8455ab;
assign v3763056 = hbusreq4 & v3a6ff9f | !hbusreq4 & v8455ab;
assign bfe049 = hmaster0_p & v3a70fd5 | !hmaster0_p & b20520;
assign v3761c5e = hmaster0_p & v373221a | !hmaster0_p & !v37744d9;
assign v37445b9 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v3778528;
assign ce69d1 = hbusreq6 & v37495dc | !hbusreq6 & v3a635ea;
assign v3774d86 = hmaster2_p & v3a635ea | !hmaster2_p & v377c6b3;
assign v3a7121a = hmaster0_p & v372580e | !hmaster0_p & v3a6eb26;
assign a27bd0 = hbusreq5_p & v3a69f8e | !hbusreq5_p & v37705df;
assign v976f99 = hlock5_p & v377989c | !hlock5_p & v3a6ffca;
assign v3766846 = hbusreq7_p & v3a70510 | !hbusreq7_p & v3a6eef8;
assign v3724e60 = jx0_p & v37326be | !jx0_p & v3a63f57;
assign v375bfd5 = hlock2_p & v3a6219d | !hlock2_p & v3a64d60;
assign v3a6f665 = hbusreq8_p & v3742146 | !hbusreq8_p & v375f0f0;
assign v3a6f76b = hmaster1_p & v3754a25 | !hmaster1_p & v3735a87;
assign v3a6afef = hbusreq4 & v3a710ad | !hbusreq4 & v3755a05;
assign v3a654c1 = hlock6 & v3a6939d | !hlock6 & v3a70f74;
assign v373c3e1 = hbusreq4_p & v3a70fd5 | !hbusreq4_p & v3759749;
assign v3809142 = hgrant5_p & v373ad69 | !hgrant5_p & v3a54b84;
assign v3736141 = hbusreq0_p & v380887a | !hbusreq0_p & v373b288;
assign v377a036 = hbusreq4_p & v373409f | !hbusreq4_p & !v3a70e35;
assign v3a5bcfa = hmaster1_p & v372b8a0 | !hmaster1_p & v37440e4;
assign v375be57 = hmaster1_p & v375b429 | !hmaster1_p & v3a6ee50;
assign v3740839 = hbusreq2_p & v376144f | !hbusreq2_p & v3748797;
assign v376002d = hmaster1_p & v3a5878e | !hmaster1_p & v3747271;
assign v3770f56 = hbusreq7 & v3734cce | !hbusreq7 & v373abcf;
assign v373fe6f = hgrant6_p & v3a5ae1b | !hgrant6_p & v8455ab;
assign v3a71338 = hmaster1_p & v375646d | !hmaster1_p & v3a541ec;
assign v3a5c538 = hmaster2_p & v8455ab | !hmaster2_p & v3a7162d;
assign v3a6cc78 = hmaster0_p & v8455ab | !hmaster0_p & !v3776ca9;
assign v375cdee = hbusreq4_p & v3763d10 | !hbusreq4_p & v1e378da;
assign v37253dc = hbusreq5_p & v3a6ff6f | !hbusreq5_p & v8455ab;
assign v3a6c007 = hlock4 & v3a6d558 | !hlock4 & v3747b3c;
assign v3737ca0 = jx1_p & v3a5eb0f | !jx1_p & v3a5842b;
assign v3768d79 = hbusreq2_p & v375ac70 | !hbusreq2_p & v8455ab;
assign v37359cf = hmaster1_p & v3a56c1f | !hmaster1_p & v37365c6;
assign v3743bc5 = hmastlock_p & v373e5f1 | !hmastlock_p & v8455ab;
assign v3a646f8 = hbusreq0_p & v3a70641 | !hbusreq0_p & v8455e7;
assign v3742358 = hbusreq7_p & v373540f | !hbusreq7_p & !v373bc8f;
assign v372c524 = hbusreq5 & v374b51f | !hbusreq5 & v8455ab;
assign v377b706 = hmaster0_p & v3726699 | !hmaster0_p & v37565ce;
assign v377e181 = hlock6_p & v3a5b68a | !hlock6_p & !v8455ab;
assign v374910b = hbusreq3_p & v3747eef | !hbusreq3_p & v376049c;
assign v37fc910 = hlock6 & v3757ec4 | !hlock6 & v37314b5;
assign v37342ec = hmaster3_p & v3733a4c | !hmaster3_p & v3a5d153;
assign v3724df8 = hbusreq5_p & v3745706 | !hbusreq5_p & v3a711ab;
assign v37744c1 = hlock3 & v3a60f85 | !hlock3 & v374e5e4;
assign v3743efa = hmaster0_p & v37701a0 | !hmaster0_p & v3a64c71;
assign v377913f = stateG10_1_p & v8455ab | !stateG10_1_p & v3752ef1;
assign v3a6a312 = hmaster2_p & v8455b0 | !hmaster2_p & v3776685;
assign v37754ac = jx0_p & v3a6f5ec | !jx0_p & v37c03ff;
assign v377bca1 = hbusreq4 & v3764978 | !hbusreq4 & !v8455ca;
assign v373cae5 = hlock5_p & v374d525 | !hlock5_p & !v375e039;
assign v377241f = hmaster1_p & v375f55e | !hmaster1_p & v3729988;
assign v372fa70 = hgrant6_p & v8455ab | !hgrant6_p & v37439b2;
assign v3a5db8b = hgrant6_p & v3a6eaf4 | !hgrant6_p & !v37317c0;
assign v377d705 = hgrant0_p & v3759d36 | !hgrant0_p & v8455ab;
assign v3a70a34 = hgrant0_p & v3747c3e | !hgrant0_p & v8455ab;
assign v37351a7 = hmaster3_p & v3732df3 | !hmaster3_p & v3a5d176;
assign v3a6e614 = hbusreq7_p & v3a5bbc1 | !hbusreq7_p & v372967b;
assign v375780e = hmaster1_p & v37763bd | !hmaster1_p & v3a6cae3;
assign v3757024 = hlock6_p & v3a676d6 | !hlock6_p & !v373c755;
assign v3a553aa = hmaster2_p & v377c7ae | !hmaster2_p & v35772a6;
assign v3775379 = hgrant7_p & v376ebc7 | !hgrant7_p & !v8455ab;
assign v37299d5 = hbusreq7_p & v3a29760 | !hbusreq7_p & v37525e0;
assign v3727e15 = hmastlock_p & v3a59918 | !hmastlock_p & !v8455ab;
assign v3a66d2e = hbusreq7_p & v377d27f | !hbusreq7_p & v37488cb;
assign v3779fec = hlock0_p & v3a6bddd | !hlock0_p & v372fe5f;
assign v3755ffc = hmaster0_p & v3a70a96 | !hmaster0_p & v3737c3f;
assign v372f357 = hlock7_p & v3764210 | !hlock7_p & !v376c784;
assign v3a5e620 = hmaster2_p & v3a635ea | !hmaster2_p & v3736afd;
assign v1e377bd = hbusreq1 & v373fe5e | !hbusreq1 & !v3753f1a;
assign v3a57037 = hmaster1_p & v372f6d3 | !hmaster1_p & v3723e23;
assign v3a70ec4 = hmaster3_p & v3756fee | !hmaster3_p & v8455ab;
assign v374e692 = hmaster2_p & v8455e7 | !hmaster2_p & v373d825;
assign v3a6f1bf = hmaster0_p & v377598a | !hmaster0_p & v3a61c70;
assign v377ab78 = hmaster1_p & v8455ab | !hmaster1_p & v3a59fbc;
assign v374cab1 = hbusreq5_p & v3753f82 | !hbusreq5_p & !v3764818;
assign v3a600a8 = hmaster1_p & v8455ab | !hmaster1_p & v3a6b29f;
assign v372383a = hlock6_p & v37270d9 | !hlock6_p & v8455e7;
assign v3774ee5 = hbusreq0 & v3754922 | !hbusreq0 & v3a5c6d8;
assign v3749520 = hbusreq7 & v375bc49 | !hbusreq7 & v373340f;
assign v3751ca5 = stateG10_1_p & v3764463 | !stateG10_1_p & !v3806572;
assign v3751719 = hbusreq0 & v372d86a | !hbusreq0 & v377226d;
assign v373c721 = hmaster2_p & v376da22 | !hmaster2_p & a4764c;
assign v375811e = hbusreq6_p & v3748797 | !hbusreq6_p & v3a5cd6c;
assign v374d969 = hlock5 & v3a674c2 | !hlock5 & v374d778;
assign v372a7ae = hgrant2_p & v3a7080a | !hgrant2_p & !v39e9c97;
assign v2acb110 = hbusreq5 & d390f8 | !hbusreq5 & v3760314;
assign v3a6f2e1 = hbusreq6_p & v377cfd9 | !hbusreq6_p & !v372ee7e;
assign v376db07 = stateG10_1_p & v8455ab | !stateG10_1_p & !v3a637dd;
assign v377445c = hbusreq4 & v374eab4 | !hbusreq4 & v37334a3;
assign v3774074 = hburst0 & v372b0cd | !hburst0 & v3752f78;
assign v3755640 = jx0_p & v3a6ba88 | !jx0_p & v376373e;
assign v37761b6 = hbusreq3 & v374cab9 | !hbusreq3 & v37674c1;
assign v3a711a4 = hbusreq6_p & v372a5c8 | !hbusreq6_p & v33790e7;
assign v3a67d3d = hmaster2_p & v8455ab | !hmaster2_p & v3727f14;
assign v3a6bf12 = hgrant6_p & v374852b | !hgrant6_p & v3742a62;
assign v3a65760 = jx0_p & v3767640 | !jx0_p & v37291c7;
assign v375f479 = stateA1_p & v3a6efc9 | !stateA1_p & !v3a71085;
assign v3a71427 = hmaster0_p & v373c076 | !hmaster0_p & v37662e7;
assign a4e409 = jx1_p & v3a7025c | !jx1_p & v3a7061f;
assign v3745d1e = hmaster1_p & v3a635ea | !hmaster1_p & v3a70f0d;
assign v37636e4 = hbusreq2 & v3767f33 | !hbusreq2 & v8455e7;
assign v37398e5 = hmaster2_p & v3764881 | !hmaster2_p & !v3a60f71;
assign v23fe339 = hbusreq4_p & v376e854 | !hbusreq4_p & v3726ae2;
assign v3a5754b = hgrant3_p & v8455ab | !hgrant3_p & v37544fa;
assign v3729792 = hbusreq5_p & v3768e52 | !hbusreq5_p & v8455ab;
assign v3732f54 = hmaster2_p & v37536ae | !hmaster2_p & !v3751510;
assign v3755d20 = hbusreq5 & v376b3d0 | !hbusreq5 & v3a6513d;
assign v3767892 = hbusreq4 & v3a54919 | !hbusreq4 & v37696b6;
assign v375fbc0 = hgrant3_p & v372ad53 | !hgrant3_p & v375ac48;
assign v3a70f62 = hmaster0_p & v3a7076e | !hmaster0_p & v3a6e872;
assign v37625a0 = hlock5_p & v37503c2 | !hlock5_p & v374e210;
assign v3a6667e = hbusreq1 & v372fc81 | !hbusreq1 & !v8455ab;
assign v376a06c = hmaster1_p & v3a69b19 | !hmaster1_p & v376314e;
assign v375559b = hbusreq4 & v8455b0 | !hbusreq4 & v373cc68;
assign v373f3dd = hmaster0_p & v374f307 | !hmaster0_p & v23fdbc1;
assign v372c0f4 = hbusreq3_p & v375a4b3 | !hbusreq3_p & !v373b9a9;
assign d73f1d = hmaster2_p & v3a61517 | !hmaster2_p & v373511d;
assign v3755167 = hgrant6_p & v8455ab | !hgrant6_p & v3742370;
assign v376079a = hmaster3_p & v3a69203 | !hmaster3_p & v37711cd;
assign v376d19f = hmaster2_p & v377bb3a | !hmaster2_p & v8455b0;
assign v3a6856a = hgrant5_p & v376d52a | !hgrant5_p & v3740af7;
assign v375c675 = hbusreq0 & v3a705ad | !hbusreq0 & v8455ab;
assign bb3b0a = hmaster1_p & v376b662 | !hmaster1_p & v3a62ce4;
assign v3a68183 = hgrant5_p & v8455ab | !hgrant5_p & v374dbdf;
assign v376ea5c = hmaster0_p & v373bb6c | !hmaster0_p & v3731d67;
assign v375e5ed = hbusreq5 & v37357d0 | !hbusreq5 & v3a63f9a;
assign v3a714ef = hmaster0_p & v3a7007e | !hmaster0_p & v8455ab;
assign v39eb532 = hbusreq6_p & v3a6f6b6 | !hbusreq6_p & v23fe189;
assign v3726a09 = hbusreq7_p & v3a6b896 | !hbusreq7_p & v37431a0;
assign v3776649 = hbusreq4_p & v380700c | !hbusreq4_p & !v8455ab;
assign v3a5a884 = hlock8 & v377e547 | !hlock8 & v3748299;
assign v3774628 = hbusreq5 & v376702a | !hbusreq5 & v3754c51;
assign v375c54c = hbusreq7_p & v37421c0 | !hbusreq7_p & v372ab1b;
assign v3a5943e = hmaster0_p & v3734967 | !hmaster0_p & v3a692c3;
assign v3723b86 = hbusreq4 & v3a55cf2 | !hbusreq4 & v3737028;
assign v3a6dd29 = hbusreq4_p & v3767b70 | !hbusreq4_p & v375af43;
assign v37651cc = hmaster0_p & v3775303 | !hmaster0_p & v3a5bf75;
assign v3753a06 = hbusreq6_p & v376e89b | !hbusreq6_p & v376b88d;
assign v3763eaa = busreq_p & v3a62a9d | !busreq_p & v8455e1;
assign v3a67fea = hgrant4_p & v3a652de | !hgrant4_p & !v37584c6;
assign v376ebe6 = hgrant6_p & v8455ab | !hgrant6_p & v3a61f3c;
assign v3731e31 = hgrant6_p & v375f2ec | !hgrant6_p & v37674a5;
assign v377081e = hbusreq7 & v3a70b9b | !hbusreq7 & v3734279;
assign v3a71492 = hbusreq8 & v3758b56 | !hbusreq8 & v374d6f6;
assign v3a6f09a = hgrant6_p & v377f09a | !hgrant6_p & !v37663b5;
assign v3a5544e = hmaster1_p & v3a70528 | !hmaster1_p & v3764daf;
assign v37551b8 = hmaster0_p & v3a54c2e | !hmaster0_p & v3a5aaf9;
assign v3733e4f = hmaster0_p & v3a5a01b | !hmaster0_p & v3a63866;
assign v3740762 = hmaster0_p & v376a297 | !hmaster0_p & v376b540;
assign v37745eb = hbusreq5 & v373ec34 | !hbusreq5 & v377c0bd;
assign v23fde6d = hmaster1_p & v3732a75 | !hmaster1_p & b9675e;
assign v8ed2d8 = hbusreq6_p & v3a55630 | !hbusreq6_p & v3a7089f;
assign v377e928 = hbusreq1_p & v8455b6 | !hbusreq1_p & !v375d651;
assign v3a66292 = hmaster2_p & v3a55c0c | !hmaster2_p & v3772935;
assign v3a5d2bc = hlock0 & v3a5f9e6 | !hlock0 & v3a6d500;
assign v375d8f8 = hbusreq8 & v3a5de59 | !hbusreq8 & v3a58723;
assign v3a70f4a = hmaster2_p & v8455ab | !hmaster2_p & !v373ad95;
assign v375792f = hmaster2_p & v8455ab | !hmaster2_p & v3764825;
assign v3742476 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v3a603f3;
assign v373dd82 = hbusreq1 & v3806db7 | !hbusreq1 & v372fba5;
assign v3761019 = hbusreq5_p & v3769740 | !hbusreq5_p & v3731aac;
assign v377b481 = hlock7 & v375c144 | !hlock7 & v3808e88;
assign v37284d5 = hbusreq0 & v3735c51 | !hbusreq0 & v3a6f434;
assign v3a714be = hgrant6_p & v8455ca | !hgrant6_p & v3737075;
assign v37355d8 = hbusreq4_p & v372c84a | !hbusreq4_p & v376871e;
assign v37389db = hbusreq3_p & v3a6ff3c | !hbusreq3_p & v3759947;
assign v3745366 = hgrant6_p & v375f3e2 | !hgrant6_p & v376865d;
assign v3a6b57d = hbusreq7 & v2092ee9 | !hbusreq7 & v3a58723;
assign v3a5d134 = hgrant4_p & v3777f86 | !hgrant4_p & v3a5f9d2;
assign v3a59314 = hbusreq5_p & v374ff84 | !hbusreq5_p & v8455ab;
assign v3730fb9 = hlock7_p & v3742132 | !hlock7_p & v3744751;
assign v3a619a2 = hmaster2_p & v374513e | !hmaster2_p & v3a5e544;
assign v3a7151d = hready & v3775ca5 | !hready & v23fdab8;
assign v372dcaa = hmaster2_p & v376501e | !hmaster2_p & v3a716a0;
assign v376fbd0 = hbusreq6 & v3a6c0f1 | !hbusreq6 & !v8455ab;
assign v372d773 = hbusreq5 & v37690da | !hbusreq5 & v3a7129c;
assign v375bd1f = hbusreq3 & v376d1e2 | !hbusreq3 & v3a69487;
assign v3741c76 = hbusreq0 & v3a59b5f | !hbusreq0 & v9e2dd1;
assign v3a635eb = hmaster3_p & v37374bc | !hmaster3_p & v376bc75;
assign v3761480 = stateA1_p & v373f4d3 | !stateA1_p & v37464c8;
assign v377df1a = hbusreq7 & v373e062 | !hbusreq7 & v372d811;
assign v3a54264 = hmaster0_p & v3a63ea7 | !hmaster0_p & v3a711c0;
assign v377d4a6 = hbusreq6 & v37436bc | !hbusreq6 & v8455ab;
assign v3a6fec6 = hbusreq7 & v3a55491 | !hbusreq7 & v377386a;
assign v3a62dae = hlock7 & v3753fe3 | !hlock7 & v37750a5;
assign v373087b = hbusreq6 & v373c2ec | !hbusreq6 & v375da82;
assign v3a5c0d4 = hbusreq6_p & v3a7093a | !hbusreq6_p & !v8455ab;
assign v374e86a = hbusreq5_p & v372dcac | !hbusreq5_p & v3730be3;
assign v37485e2 = hmaster0_p & v3a70f68 | !hmaster0_p & v376374b;
assign v3755d19 = hmaster0_p & v3772229 | !hmaster0_p & v377312f;
assign v3a6a1b7 = hmaster2_p & v3770754 | !hmaster2_p & v3a7085f;
assign v3a5d93f = hgrant6_p & v3738be9 | !hgrant6_p & v372546e;
assign ca32a1 = hmaster1_p & v2093132 | !hmaster1_p & v3760c32;
assign v376fb50 = hgrant3_p & v3a70ec3 | !hgrant3_p & v377094b;
assign v375b045 = hbusreq6_p & v3a6fc17 | !hbusreq6_p & v37722c4;
assign v376e0cd = hmaster2_p & v3733383 | !hmaster2_p & v3a660f2;
assign v372c00b = hmaster2_p & v8455ab | !hmaster2_p & v376f167;
assign v3a567b7 = hmaster2_p & v3a62826 | !hmaster2_p & v37598ab;
assign v3a5f75a = hbusreq6 & v3a67ec4 | !hbusreq6 & v3a6fdef;
assign v376bf0a = hgrant2_p & v8455ab | !hgrant2_p & v374b690;
assign v372af40 = hbusreq5_p & v1e374d4 | !hbusreq5_p & v373861f;
assign v3a6eaf6 = jx0_p & v374f16d | !jx0_p & v3a65af6;
assign v37630e2 = hlock8 & v373de1d | !hlock8 & v3767be8;
assign v372df69 = hgrant1_p & v90fd44 | !hgrant1_p & v8455ab;
assign v3a70f05 = jx0_p & v3a70cef | !jx0_p & v3767537;
assign v372cb88 = hburst1 & v373d9e5 | !hburst1 & v3a66bdb;
assign v3a70e21 = hbusreq2_p & v372c3d4 | !hbusreq2_p & !v3a5ef5c;
assign v372b33d = hbusreq5 & v3729382 | !hbusreq5 & v3774bad;
assign v3727195 = hmaster1_p & v8455e7 | !hmaster1_p & v37308bc;
assign v3a710dd = hbusreq0 & v377ecd4 | !hbusreq0 & v3776852;
assign v3a712d1 = hlock0 & v3a5aacb | !hlock0 & v3a6f08a;
assign v3a6f843 = hlock8 & v377b7d0 | !hlock8 & v373643b;
assign v3a6b37c = hbusreq6 & v375f317 | !hbusreq6 & v3a6f4bc;
assign v374c3ff = hbusreq5 & v3a709fc | !hbusreq5 & v3a67d83;
assign v372b5ed = hmaster3_p & v3a6ef19 | !hmaster3_p & v3a6e2ec;
assign v372f83b = hbusreq4 & v3a5dd17 | !hbusreq4 & v3a7162d;
assign v3741e56 = hmaster2_p & v3a712c4 | !hmaster2_p & v3a5f7c5;
assign v3778567 = hgrant6_p & v3a57f59 | !hgrant6_p & v3757b0e;
assign v2ff87b0 = hbusreq4_p & v375b26a | !hbusreq4_p & v3778352;
assign v37740e0 = hbusreq3 & v3a6557d | !hbusreq3 & v372cc25;
assign v37558e4 = hbusreq4_p & v374304d | !hbusreq4_p & v373e814;
assign v3739c30 = hgrant3_p & v3772d9a | !hgrant3_p & v2619ae8;
assign v3a6ff30 = hbusreq4_p & v3a704dc | !hbusreq4_p & !v3731de2;
assign v3a7076c = hlock4_p & v2ff9190 | !hlock4_p & v8455ab;
assign v375491e = hlock4 & v3738679 | !hlock4 & v3a6f3da;
assign v37548b3 = hmaster1_p & v3772183 | !hmaster1_p & v377a1dd;
assign v376669c = hmaster2_p & v37320bf | !hmaster2_p & v3a71026;
assign v372809d = hmaster2_p & v373f647 | !hmaster2_p & !v8455ab;
assign v377217c = hbusreq1_p & v3a6e66e | !hbusreq1_p & !v3a6eafc;
assign v3752fbc = hbusreq6_p & v3775bca | !hbusreq6_p & v8455ab;
assign v3724987 = hmaster1_p & v372fc6c | !hmaster1_p & v3a5efc4;
assign v3a7106f = hbusreq3_p & v3a635ea | !hbusreq3_p & v3742b31;
assign v1e37b74 = hmaster2_p & v3736ee0 | !hmaster2_p & v37267a5;
assign v3a6becb = hgrant6_p & v209323b | !hgrant6_p & v374874a;
assign v3746ab6 = hbusreq6_p & v374c33a | !hbusreq6_p & v3737534;
assign v374a950 = hbusreq6_p & v3a62826 | !hbusreq6_p & v35b774b;
assign v3a563ed = hgrant4_p & v8455ab | !hgrant4_p & !v374bda9;
assign v3734041 = hmaster1_p & v3a619c0 | !hmaster1_p & v377ac0f;
assign v3775ad3 = hgrant4_p & v3a7049a | !hgrant4_p & v3a60723;
assign v3731f6b = hbusreq5 & v374314f | !hbusreq5 & v37476b8;
assign v3a6f92f = hbusreq2_p & v3a68c1f | !hbusreq2_p & v3a57f59;
assign v3768904 = hmaster0_p & v360d166 | !hmaster0_p & v374d4d3;
assign v375a3dc = hgrant4_p & v8455ab | !hgrant4_p & v3a5984d;
assign v377516c = hmaster1_p & v3a66110 | !hmaster1_p & v3a6f6a8;
assign v3a70071 = hbusreq5_p & v3730a73 | !hbusreq5_p & v3760e6e;
assign v372a7c2 = hready_p & v3a70c21 | !hready_p & !v8455ab;
assign v3a5cb95 = hmaster1_p & v3806a7b | !hmaster1_p & v3a614d5;
assign v372a8fd = hbusreq7_p & v372f0e0 | !hbusreq7_p & v3a6b9d9;
assign v3a70c35 = hbusreq0 & v375a8ad | !hbusreq0 & v376362f;
assign v375e9c0 = hmaster3_p & v3739d49 | !hmaster3_p & v372a25a;
assign v3770d41 = hbusreq4 & v374ad30 | !hbusreq4 & v373a341;
assign v3727ee4 = hbusreq4 & v372ea48 | !hbusreq4 & v8455ab;
assign v3a67e2e = hgrant1_p & v375d182 | !hgrant1_p & v3a70d71;
assign v3808994 = hbusreq5 & v375609e | !hbusreq5 & v373de86;
assign v3745473 = jx0_p & v97c94a | !jx0_p & v3746cc3;
assign v3a69a1b = hbusreq5_p & v3759bdb | !hbusreq5_p & v3779e72;
assign v3757b16 = hgrant4_p & v8455c2 | !hgrant4_p & v3770161;
assign v372c46e = hmaster2_p & v372e27b | !hmaster2_p & v3a5c33d;
assign v3a6924e = hmaster1_p & v8455ab | !hmaster1_p & v3725d48;
assign v373d139 = hgrant0_p & v8455ab | !hgrant0_p & v3806fbf;
assign v373c991 = hgrant6_p & v3a70193 | !hgrant6_p & v3a593cb;
assign v3a622d0 = hbusreq3 & v375d9f8 | !hbusreq3 & !v3766238;
assign v3772231 = hlock5_p & v372505f | !hlock5_p & !v8455ab;
assign v3a7106b = hmaster2_p & v8455ab | !hmaster2_p & v372a068;
assign v372b4cb = hbusreq4_p & v3770719 | !hbusreq4_p & v3725717;
assign v37446b5 = hbusreq4 & v37482f8 | !hbusreq4 & !v3a7127f;
assign v373a16b = hmaster2_p & v372673d | !hmaster2_p & v3a70374;
assign v3a66088 = hmaster2_p & v3a6823d | !hmaster2_p & v3738d43;
assign v376984d = hmaster2_p & v3a54eae | !hmaster2_p & v3764418;
assign v37337fd = hlock5_p & v3a71194 | !hlock5_p & abd043;
assign v3775bf6 = hbusreq1_p & v376dc21 | !hbusreq1_p & v3774fa8;
assign v373df1f = hmaster0_p & v3775928 | !hmaster0_p & v375058e;
assign v372f02f = hbusreq3_p & v372ec1c | !hbusreq3_p & v3a69487;
assign v373a1b4 = hgrant4_p & v375c697 | !hgrant4_p & v3723ba5;
assign v3a5f592 = hgrant5_p & v8455c6 | !hgrant5_p & v37447e9;
assign v3740b8d = hgrant6_p & v37598ab | !hgrant6_p & v3773a6b;
assign v376581d = hmaster0_p & v3778395 | !hmaster0_p & v8455e7;
assign v3a6f926 = hmaster2_p & v8455e7 | !hmaster2_p & v376f2f8;
assign v3a6ffd0 = hbusreq0 & v3760088 | !hbusreq0 & v3a6f775;
assign v3a6b001 = hgrant7_p & v375e1f6 | !hgrant7_p & v375cf46;
assign v3725717 = hbusreq2_p & v3747302 | !hbusreq2_p & v3743b9e;
assign v3a6dcb9 = hbusreq0 & v3728823 | !hbusreq0 & v3a705e8;
assign v3723df0 = hmaster1_p & v376e605 | !hmaster1_p & v376c1c3;
assign v376d86c = hbusreq4_p & v3744f62 | !hbusreq4_p & v8455ab;
assign v3773796 = hbusreq8_p & v372a1ab | !hbusreq8_p & v3a5df70;
assign v376d0ff = hmaster2_p & v377f734 | !hmaster2_p & v3751491;
assign v373fe5e = locked_p & v376c211 | !locked_p & !v8455ab;
assign v3750c38 = hbusreq6_p & v375a0b3 | !hbusreq6_p & v3a5c5b5;
assign v3a7063c = hlock6_p & v39a4dbb | !hlock6_p & v3736847;
assign v377362f = hbusreq2 & v3a6ab5f | !hbusreq2 & !v2aca977;
assign v373cc9a = hbusreq5_p & v3728fd2 | !hbusreq5_p & !v8455ab;
assign v372d924 = hlock4_p & v380761d | !hlock4_p & v8455ab;
assign v3a6d93d = hbusreq1_p & v8455ab | !hbusreq1_p & !v375bb3a;
assign v375ef27 = hbusreq3_p & v374f609 | !hbusreq3_p & v3a6cacb;
assign v3a67dbc = hlock6 & v374cd10 | !hlock6 & v3727615;
assign v3a70e9f = hgrant0_p & v8455ab | !hgrant0_p & v3752a7e;
assign v372668c = hbusreq5 & v325c90f | !hbusreq5 & v3764761;
assign v3a60013 = hmaster1_p & v3a70101 | !hmaster1_p & v374122a;
assign v3a6e236 = hbusreq3_p & v3a70208 | !hbusreq3_p & v37497b1;
assign v2aca770 = hlock3_p & v3767ed6 | !hlock3_p & v8455b0;
assign v37674c1 = locked_p & v373bdac | !locked_p & v8455ab;
assign v3a70889 = hgrant2_p & v3a680b9 | !hgrant2_p & v377e52f;
assign v3764caf = hbusreq2 & v374ad1e | !hbusreq2 & v37677ee;
assign v3a5bbbb = hbusreq5 & v373d3ec | !hbusreq5 & v8455ab;
assign v3779fbc = hmaster1_p & v377b24b | !hmaster1_p & v377410f;
assign v3806ec4 = hgrant2_p & v8455ab | !hgrant2_p & v3a6c449;
assign v3722b92 = hbusreq4 & v37739f4 | !hbusreq4 & !v3a576d0;
assign v3a6eab0 = hgrant0_p & v8455ab | !hgrant0_p & v37417f6;
assign v37c36b9 = hbusreq7_p & v3763c1f | !hbusreq7_p & v3a6dbec;
assign v3a71637 = hmaster0_p & v3779a06 | !hmaster0_p & !v3741b5e;
assign v3a6f18f = hbusreq6_p & v37308a8 | !hbusreq6_p & !v8455ca;
assign v373e896 = hmaster2_p & v8455ab | !hmaster2_p & v3806dda;
assign v3772773 = hbusreq7_p & v3a70c90 | !hbusreq7_p & bfa92a;
assign v3a67a85 = hbusreq0 & v3a5b70a | !hbusreq0 & v3a55641;
assign v3751491 = hgrant4_p & v8455ab | !hgrant4_p & bae881;
assign v3763acf = hgrant3_p & v8455bd | !hgrant3_p & v374a97f;
assign v372f576 = hgrant1_p & v3a6f8c1 | !hgrant1_p & !v8455ab;
assign v373128b = hlock3 & v377ac8a | !hlock3 & v3a5a3be;
assign v9a88fd = hgrant5_p & v3a5caf4 | !hgrant5_p & !v3a693dc;
assign v3a63717 = hmaster1_p & v3a5e696 | !hmaster1_p & v373519d;
assign v376a7b5 = hbusreq6 & v3750674 | !hbusreq6 & v8455ab;
assign v3a71055 = hmaster1_p & v374a9d0 | !hmaster1_p & v3731088;
assign v374da33 = hgrant5_p & v8455c6 | !hgrant5_p & v3a6fdf9;
assign v3738c99 = hlock0_p & v3753f1a | !hlock0_p & v8455ab;
assign v3742322 = hmaster2_p & v3808ed2 | !hmaster2_p & !v8455ab;
assign v3a70327 = hgrant6_p & v3739884 | !hgrant6_p & v375d715;
assign a9f66a = hbusreq1_p & v3747302 | !hbusreq1_p & v3a71452;
assign v3a66d7e = hlock2_p & v3a63e82 | !hlock2_p & !v35772a6;
assign v374b6ee = hmaster1_p & v377d1dc | !hmaster1_p & v3808fc8;
assign v3a70ccd = hlock5 & v3743d5d | !hlock5 & v377f1ff;
assign v3772dcb = hbusreq8 & v3741863 | !hbusreq8 & v3768734;
assign v3a5d015 = hbusreq5_p & v3732736 | !hbusreq5_p & v3769a60;
assign v3a2abf4 = hbusreq5 & v3a5a2cd | !hbusreq5 & v8455ab;
assign c79715 = hlock5_p & v1e379b9 | !hlock5_p & !v8455ab;
assign v373ac95 = hmaster3_p & v3762363 | !hmaster3_p & v377dc4a;
assign v3a614d5 = hbusreq5_p & v37439a0 | !hbusreq5_p & !v376075c;
assign v3747042 = hbusreq6_p & v3a6ae2d | !hbusreq6_p & v8455ab;
assign v375884e = hgrant6_p & v375fa71 | !hgrant6_p & v3a714ff;
assign v3771a36 = jx1_p & v380a20c | !jx1_p & v3a70d88;
assign v3737672 = jx3_p & v8455ab | !jx3_p & v3a70f5f;
assign v3a6f6d5 = hmaster2_p & v3724270 | !hmaster2_p & v374ab8d;
assign v377bdb8 = hlock2_p & v8455ab | !hlock2_p & v3a6ab5f;
assign v2ff8f0a = hgrant2_p & v3a6f46a | !hgrant2_p & v3a68ad8;
assign v3a711fa = hbusreq6 & v377b4b9 | !hbusreq6 & v372462b;
assign v3728434 = hmaster3_p & v3a6a42a | !hmaster3_p & !v376b1ee;
assign v3808dd8 = hbusreq4 & v3a68f98 | !hbusreq4 & v376e041;
assign v3a6f209 = hmaster2_p & v8455ab | !hmaster2_p & v374a637;
assign v3a6f12b = hbusreq5_p & v3a5ad17 | !hbusreq5_p & v373790d;
assign v375cbe3 = hgrant6_p & v3725230 | !hgrant6_p & v37489ea;
assign v23fe1ca = hmaster1_p & v3a70154 | !hmaster1_p & v37629b0;
assign v3a6fbc9 = hlock8_p & v8455e7 | !hlock8_p & !v3a6ebc6;
assign v3a7124c = hbusreq6_p & v3a5d923 | !hbusreq6_p & v3768931;
assign v3a70f38 = hgrant5_p & v3a633ca | !hgrant5_p & v3a6fb75;
assign v3a6efb9 = hbusreq5_p & v2925cf2 | !hbusreq5_p & v3a7138e;
assign v375dff6 = hmaster0_p & b62443 | !hmaster0_p & v3a5f76b;
assign v377abd6 = hbusreq6_p & v3a6143b | !hbusreq6_p & !v39a4ca8;
assign v375dbf3 = hgrant4_p & v8455ab | !hgrant4_p & v372a5fc;
assign v372c18a = hmaster2_p & v3735512 | !hmaster2_p & v8455ab;
assign v3745039 = hbusreq2 & v23fd923 | !hbusreq2 & v375b9c1;
assign v3759d36 = hlock0_p & v3748797 | !hlock0_p & v372ebaa;
assign v37750a5 = hmaster1_p & v3a5df66 | !hmaster1_p & v374e7fa;
assign v3a6ece9 = hbusreq7_p & v3a69f2b | !hbusreq7_p & v3a70652;
assign v3a6991b = hmaster2_p & v37429a1 | !hmaster2_p & v8fac55;
assign v3a6f91a = hgrant2_p & v8455ab | !hgrant2_p & v3a7047f;
assign v376e7cf = hmaster0_p & v3754fcc | !hmaster0_p & v374e0a9;
assign v3a71650 = jx0_p & v373e86e | !jx0_p & v3758f17;
assign v376b3b0 = hbusreq1_p & v37603f4 | !hbusreq1_p & v3762bbe;
assign v372a738 = hmaster1_p & v37588cf | !hmaster1_p & v377055c;
assign v3a61580 = hlock0 & v3a612af | !hlock0 & d5ffe1;
assign v372e9ef = hmaster2_p & v374743d | !hmaster2_p & v3a68793;
assign v3775931 = hmaster0_p & v9ecbe0 | !hmaster0_p & v3754727;
assign v37438c9 = hbusreq1_p & v377857d | !hbusreq1_p & v373b288;
assign v3737f5f = stateG10_1_p & v39ebac7 | !stateG10_1_p & v3743a2c;
assign v3a7005d = hmaster0_p & v3a5fe3c | !hmaster0_p & v37759ff;
assign v3a70c80 = jx1_p & v3a70b2a | !jx1_p & d7f9ec;
assign v3738457 = hbusreq0 & v380974c | !hbusreq0 & v8455ab;
assign v376cd2f = hbusreq4_p & v3a70c3a | !hbusreq4_p & v3a70393;
assign v3757ec4 = hbusreq6 & v3a6c63e | !hbusreq6 & v3a6c5ee;
assign v3a57fa1 = hlock7_p & v3a6dfec | !hlock7_p & v3773c10;
assign v3a6c2b2 = hbusreq8_p & v3a635ea | !hbusreq8_p & v375c111;
assign v374da92 = hmaster2_p & v372f289 | !hmaster2_p & v376a6f1;
assign v3a674a8 = hgrant8_p & v374020a | !hgrant8_p & v3a7112d;
assign v3a5a980 = hgrant0_p & v8455ab | !hgrant0_p & v3a6fc2e;
assign v3743831 = hmaster1_p & v8455ab | !hmaster1_p & v3775e35;
assign v3a555d7 = hbusreq6 & v374e35e | !hbusreq6 & v8455ab;
assign v3732a95 = hgrant5_p & c8ca6f | !hgrant5_p & v3729f13;
assign v3a702e1 = hgrant6_p & v9ed516 | !hgrant6_p & v3736f3b;
assign v376f47f = hbusreq6 & v37639c6 | !hbusreq6 & v3a5b6de;
assign v8827d7 = hlock4 & v373b51b | !hlock4 & v3a5dd17;
assign v3774ab8 = hbusreq5 & v3a5e4e5 | !hbusreq5 & v374851a;
assign v2ff8e9a = hlock4 & v377870b | !hlock4 & v37611a9;
assign v374aae0 = hmaster2_p & v3a5600a | !hmaster2_p & v3a63659;
assign v3740672 = hbusreq4 & v377f865 | !hbusreq4 & v8455ab;
assign v3a6b32d = hmaster1_p & v37317da | !hmaster1_p & v3723583;
assign v377169f = hbusreq2_p & v37314f2 | !hbusreq2_p & v8455ab;
assign v3a702a7 = hgrant2_p & v3a57959 | !hgrant2_p & v374cba0;
assign v3747598 = hbusreq7 & v3a557d2 | !hbusreq7 & v3728870;
assign v3a7146f = hbusreq0 & v3a70ac7 | !hbusreq0 & v376af2d;
assign v374da4a = hlock2_p & v3743dfc | !hlock2_p & v372c8d1;
assign v376b509 = hlock0_p & v374cab9 | !hlock0_p & v8455ab;
assign v375a455 = jx0_p & v37674fb | !jx0_p & v3774b58;
assign v37586ed = hbusreq7 & v3734aa5 | !hbusreq7 & v8455ab;
assign v3a6572c = hmaster0_p & v377adf5 | !hmaster0_p & !v3a6f92f;
assign v374f12c = jx3_p & v3a70239 | !jx3_p & v377455b;
assign v3a6f382 = hbusreq5_p & v37337fd | !hbusreq5_p & v3a709d1;
assign v3774eed = hmaster1_p & v1e37405 | !hmaster1_p & v3735d84;
assign v3762e54 = hbusreq5 & v3755113 | !hbusreq5 & v3a68356;
assign v376297b = hbusreq8 & v35b70c3 | !hbusreq8 & v375f123;
assign v37573f4 = hbusreq6_p & v374ec8b | !hbusreq6_p & !v8455ab;
assign v3a66ef6 = hgrant2_p & v8455ab | !hgrant2_p & v3757656;
assign v375e9ef = hmaster1_p & v3a7002c | !hmaster1_p & v375c60f;
assign v3a6fe1b = hmaster2_p & v37791a5 | !hmaster2_p & v3754603;
assign v37505a2 = hmaster0_p & v3769ae2 | !hmaster0_p & v37755b2;
assign cfe6df = hlock6_p & v3733ea2 | !hlock6_p & v8455ab;
assign v3739bd5 = hbusreq6 & v3a5b00a | !hbusreq6 & !v8455ab;
assign v3763fdf = hgrant3_p & v3755c31 | !hgrant3_p & v3a6fdb4;
assign v3767429 = hgrant2_p & v374acbe | !hgrant2_p & v3a6f6e7;
assign v37411ca = hmaster1_p & v375058a | !hmaster1_p & v3769d79;
assign v376673b = hmaster1_p & v3724394 | !hmaster1_p & v3a6f9e7;
assign d23562 = hlock7_p & v3747804 | !hlock7_p & v3a6ded8;
assign v3746b4f = hbusreq6_p & v3740171 | !hbusreq6_p & v37457fb;
assign v3a70d71 = locked_p & v8455ab | !locked_p & v3737554;
assign v37626b9 = hbusreq7 & v374ecf9 | !hbusreq7 & v3733b90;
assign v3739dd4 = hgrant6_p & v3a70272 | !hgrant6_p & v3739732;
assign v377661c = hlock6 & v3a6f0b8 | !hlock6 & v3a70ee1;
assign v375cea7 = hbusreq1_p & v37551f2 | !hbusreq1_p & v3753353;
assign v3a7022a = hmaster1_p & v3773ee7 | !hmaster1_p & v376d4f3;
assign v376b795 = hlock6 & v3733360 | !hlock6 & v37344a0;
assign v3724994 = locked_p & v377e976 | !locked_p & v8455ab;
assign v3730c69 = hlock2_p & v3a6219d | !hlock2_p & v372554a;
assign v3a701d9 = hbusreq6 & v3a7008c | !hbusreq6 & v8455ab;
assign v3377aee = hbusreq5 & v3728493 | !hbusreq5 & v374a36b;
assign v3765248 = hmaster1_p & v3769093 | !hmaster1_p & v3742b92;
assign ca095d = hmaster1_p & v3a70209 | !hmaster1_p & v374bb9f;
assign v3a6f8dc = hgrant0_p & v3a70829 | !hgrant0_p & !ad2d05;
assign v376915a = hbusreq0_p & v8455ab | !hbusreq0_p & v3768aaa;
assign v3768196 = hmaster0_p & v3a68a46 | !hmaster0_p & v3a6fc5e;
assign v375cf04 = hmaster0_p & v376fa3e | !hmaster0_p & v37614c1;
assign v375db57 = hmaster2_p & v377234d | !hmaster2_p & v374ab8d;
assign v3a6f121 = hbusreq7_p & v374fe2d | !hbusreq7_p & v3a657d3;
assign v376efaa = hmaster2_p & v3773200 | !hmaster2_p & v377234d;
assign v372543f = hgrant5_p & v8455ab | !hgrant5_p & v3761d2f;
assign v376360a = hbusreq5 & v3a656ca | !hbusreq5 & v8455bf;
assign v3726ef1 = hbusreq3 & v3748900 | !hbusreq3 & !v8455ab;
assign v3a6c0e4 = hgrant0_p & v3731bcf | !hgrant0_p & v3753cc4;
assign v3778345 = hgrant3_p & v374383b | !hgrant3_p & v37711e2;
assign v3743252 = hlock1_p & v8455ab | !hlock1_p & v373cf4e;
assign v375989b = hbusreq6_p & v374e9b8 | !hbusreq6_p & v8455b3;
assign v3a6d74f = hgrant3_p & v373e642 | !hgrant3_p & v3741216;
assign v375f6c7 = hmaster2_p & v3a70c13 | !hmaster2_p & v3a6c004;
assign c9bec3 = hbusreq4_p & v375896e | !hbusreq4_p & !v39a4f17;
assign v3a70e62 = hbusreq6_p & v373f883 | !hbusreq6_p & v3737534;
assign v3a6f2a4 = hgrant6_p & v3a605b5 | !hgrant6_p & v377e582;
assign v373a77b = hgrant5_p & v37400f3 | !hgrant5_p & v3736c8c;
assign v372610a = hbusreq0 & v37419fd | !hbusreq0 & v3a700ac;
assign v376b193 = hbusreq5 & v3a71326 | !hbusreq5 & v3a66632;
assign v374d6f4 = hbusreq3_p & v3a5e24d | !hbusreq3_p & v373b303;
assign v3753233 = hbusreq1_p & v374ed4b | !hbusreq1_p & v8455b6;
assign v3a56069 = hbusreq5_p & v372b9c5 | !hbusreq5_p & v375a4d0;
assign v3757e28 = hlock4_p & v376011a | !hlock4_p & v373c441;
assign v3a71600 = hlock4 & v3751c77 | !hlock4 & v374663d;
assign v376a2de = hmaster0_p & v377bb3a | !hmaster0_p & v374aa46;
assign v37400f3 = hmaster1_p & v377e7ac | !hmaster1_p & !v373a11f;
assign v3a6e318 = hmaster2_p & v3738061 | !hmaster2_p & v37787c1;
assign v3762759 = hmaster2_p & v3a713df | !hmaster2_p & v376d374;
assign v35ba2dd = hgrant2_p & v8455ab | !hgrant2_p & v3a68016;
assign v373024e = hmaster1_p & v376142a | !hmaster1_p & v375f888;
assign v372b2b4 = hbusreq7_p & v3a6fbd3 | !hbusreq7_p & v377583c;
assign v3727472 = hgrant4_p & v37786a6 | !hgrant4_p & v3a5e244;
assign v373216d = hgrant5_p & v373ad69 | !hgrant5_p & v3760690;
assign v3a64c71 = hmaster2_p & v37315c5 | !hmaster2_p & v3760509;
assign v37560c9 = hbusreq5_p & v373f64f | !hbusreq5_p & v3a5b807;
assign v372b6bc = hbusreq4_p & v3a6fc27 | !hbusreq4_p & v8455ab;
assign v3a63688 = hmaster1_p & v3a635ea | !hmaster1_p & v3728d57;
assign v373e5f3 = hbusreq8_p & v3769ba0 | !hbusreq8_p & v374d95f;
assign v3733c53 = hmaster2_p & v3a7142f | !hmaster2_p & v3767848;
assign v3a7026f = hbusreq4 & v3778787 | !hbusreq4 & v3a64af7;
assign v377ad9b = hmaster2_p & adf78a | !hmaster2_p & v3a6f0f6;
assign v3a6fd52 = hmaster0_p & v38087c5 | !hmaster0_p & v373ea19;
assign v3763788 = hgrant1_p & v3732dc6 | !hgrant1_p & v8455ab;
assign v375cf46 = jx1_p & v374b237 | !jx1_p & !v3a704b7;
assign v3a5a510 = hbusreq3_p & v3a5c945 | !hbusreq3_p & v3a57f59;
assign v374352b = hbusreq6_p & v3723abc | !hbusreq6_p & !v3747167;
assign v3a5dd10 = hmaster1_p & v3a708ee | !hmaster1_p & v3727187;
assign v3760353 = hbusreq0 & v37237cd | !hbusreq0 & v37435f7;
assign v3a6f79e = hlock2 & v3a6f418 | !hlock2 & a36a2a;
assign v3727d1e = hlock0_p & v3378ef7 | !hlock0_p & v3744710;
assign v3a61661 = hbusreq7 & v3a71483 | !hbusreq7 & v374f6c0;
assign v377f630 = hmaster1_p & v3a55542 | !hmaster1_p & v373d98d;
assign v372526a = hgrant4_p & v3739896 | !hgrant4_p & v37617de;
assign v376ea4a = hbusreq1_p & v3759032 | !hbusreq1_p & v3733e9e;
assign v375101b = hbusreq8 & v3776084 | !hbusreq8 & v8455ab;
assign v3a6eff3 = hmaster0_p & v3768d11 | !hmaster0_p & v372f9cf;
assign v3724057 = hlock0_p & v377eaf2 | !hlock0_p & v3a710b2;
assign v3a54b5d = hmaster0_p & v3746d89 | !hmaster0_p & v3a56512;
assign v3a6e7ed = hmaster0_p & v376a44f | !hmaster0_p & d54152;
assign v3807513 = hbusreq4 & v3a707ea | !hbusreq4 & v3a685c7;
assign v3807df0 = hbusreq4 & v3a70bea | !hbusreq4 & v375c70c;
assign v3a70856 = hbusreq5_p & v3740885 | !hbusreq5_p & v3a6ff12;
assign v376d34b = hbusreq3 & v372e169 | !hbusreq3 & v3748797;
assign v37578b4 = hgrant6_p & v3744cfe | !hgrant6_p & v3777692;
assign v3770855 = hbusreq2 & v86d3dc | !hbusreq2 & v3757955;
assign v3772c08 = hgrant5_p & v3765e47 | !hgrant5_p & v3a709f7;
assign v3807a23 = hgrant4_p & v376a6f1 | !hgrant4_p & v373270f;
assign v374d4e6 = hgrant4_p & v3a70d99 | !hgrant4_p & v373a972;
assign v3a697f2 = hbusreq0_p & v372dadb | !hbusreq0_p & v3761cec;
assign v372f87b = hbusreq6_p & v3a635ea | !hbusreq6_p & v3762281;
assign v374dd11 = hbusreq8_p & v3732da2 | !hbusreq8_p & v3a6f6c8;
assign v3a71330 = hbusreq4_p & v372ae9d | !hbusreq4_p & v3a6b916;
assign v3a6f410 = hbusreq8 & v377c02f | !hbusreq8 & v8455b3;
assign v375bb6b = hgrant3_p & v374d6f4 | !hgrant3_p & !v374f0a4;
assign v374610e = hbusreq2 & v3a63ff3 | !hbusreq2 & v8455ab;
assign v3a707ee = hmaster0_p & v3a6d098 | !hmaster0_p & v37261b3;
assign v3a7163a = hmaster2_p & a7adce | !hmaster2_p & v3738006;
assign v8455e1 = hmastlock_p & v8455ab | !hmastlock_p & !v8455ab;
assign v3a62bae = hgrant4_p & v372e711 | !hgrant4_p & v3751a9f;
assign v3a6aada = hmaster2_p & v3a5e24e | !hmaster2_p & !v1e38224;
assign v375bcf7 = hbusreq5_p & v3743bde | !hbusreq5_p & v3a66e6f;
assign v376c883 = hlock2 & v3809958 | !hlock2 & v3747704;
assign v3759786 = hbusreq5 & v375aff6 | !hbusreq5 & v374c6b8;
assign v376147a = hlock7_p & v373b6e9 | !hlock7_p & !v8455ab;
assign v3740d32 = hbusreq5 & v374131b | !hbusreq5 & v8455ab;
assign v3731fd2 = hbusreq5 & v3a70f4e | !hbusreq5 & v3771c85;
assign v3a6f591 = hmaster2_p & v8455ab | !hmaster2_p & v3a6f723;
assign v37378d4 = hmaster1_p & v3775dbc | !hmaster1_p & v376fd85;
assign v373859a = hmaster1_p & v376a14f | !hmaster1_p & v3a63004;
assign v37771a2 = stateA1_p & v376faea | !stateA1_p & v8455e1;
assign v377e539 = jx0_p & v3776d4b | !jx0_p & v377a7ee;
assign v373a4ef = hmaster0_p & v376f237 | !hmaster0_p & v3776cbb;
assign v3a56531 = hbusreq6_p & v3749fdc | !hbusreq6_p & v8455ab;
assign v3a5e2c8 = hmaster0_p & dc47a7 | !hmaster0_p & v376df4c;
assign v3a5e2b9 = hbusreq4_p & v3a6b572 | !hbusreq4_p & v3a6c91f;
assign v374f712 = hmaster0_p & v3a63a18 | !hmaster0_p & v375f145;
assign v372a22d = hlock5_p & v8455ab | !hlock5_p & v3a6f03d;
assign a26159 = hgrant4_p & v3a708f2 | !hgrant4_p & v3a70c1f;
assign v3776836 = hlock8 & v3742210 | !hlock8 & v3a705da;
assign v377e298 = hmaster2_p & v3747302 | !hmaster2_p & v3748d67;
assign v37605e6 = hmaster2_p & v372b231 | !hmaster2_p & v3a706f1;
assign v3a70dad = hmaster3_p & v3774a1b | !hmaster3_p & v37607c6;
assign v372dbe7 = hbusreq8 & v37436e6 | !hbusreq8 & v8455bb;
assign v3750a45 = hmaster2_p & v8455ab | !hmaster2_p & v3758133;
assign v37306cd = hbusreq6 & v372c60a | !hbusreq6 & v8455bf;
assign v377535a = hbusreq6 & v372b5f5 | !hbusreq6 & v8455ab;
assign v372e8f2 = hbusreq5_p & v372a27f | !hbusreq5_p & v8455ab;
assign v376cf8c = hbusreq2_p & v3a70272 | !hbusreq2_p & !v3a5b68a;
assign v373c61e = hbusreq4_p & v3729bf3 | !hbusreq4_p & v3a6fd1a;
assign v3a7031c = hmaster0_p & v3758fa8 | !hmaster0_p & v3a58b13;
assign v374312f = hmaster1_p & v8455ab | !hmaster1_p & v3746e10;
assign v372d59d = hmaster1_p & v3742afe | !hmaster1_p & v3a6b90e;
assign v37660f0 = hlock5 & v37786f3 | !hlock5 & v372cf70;
assign v3a70f32 = hgrant4_p & v8455ab | !hgrant4_p & v377e87e;
assign v3752d9f = hmaster1_p & v3757966 | !hmaster1_p & v375d17c;
assign v3808dcb = hmaster1_p & v8455ab | !hmaster1_p & v374677f;
assign v375320f = hlock8 & v3768d56 | !hlock8 & v372c492;
assign v37297cb = hgrant4_p & v374bb76 | !hgrant4_p & v3728625;
assign v3746540 = hgrant4_p & v3735525 | !hgrant4_p & v373484e;
assign v3a63f80 = hbusreq7 & v3a70bfb | !hbusreq7 & v3a60276;
assign v3a59ea2 = hmaster2_p & v373d791 | !hmaster2_p & v376fd4e;
assign v3a71679 = hmaster2_p & v3a635ea | !hmaster2_p & v3735525;
assign v375e22b = hlock3 & v38072fd | !hlock3 & v3a56e5e;
assign v3a6f7b2 = hgrant6_p & v8455ab | !hgrant6_p & !v8455ed;
assign v3732c96 = hgrant5_p & v3a6fa02 | !hgrant5_p & v3a70ed5;
assign v372f71f = hmaster1_p & v3757dd1 | !hmaster1_p & v3722b17;
assign v3a6f700 = hmaster2_p & v3745181 | !hmaster2_p & v37600c0;
assign v37560f1 = hmaster2_p & v3a62caa | !hmaster2_p & v3a6f2cb;
assign v3a7127c = hmaster0_p & v8455ab | !hmaster0_p & !v376a6f1;
assign v3759bd0 = hmaster2_p & v374b887 | !hmaster2_p & v376c4e8;
assign v3a56b19 = hbusreq0 & v3a651b5 | !hbusreq0 & v373e814;
assign v3a6eb22 = hbusreq5 & v3a6e031 | !hbusreq5 & v3378fc3;
assign v3777c59 = hgrant4_p & v3a5a68d | !hgrant4_p & !d648e4;
assign v3747314 = hbusreq0 & v3761006 | !hbusreq0 & v374ee8d;
assign v3744983 = hlock2_p & v373c1d7 | !hlock2_p & v3740fef;
assign v3a54108 = hbusreq2_p & v3a62628 | !hbusreq2_p & v3a658bf;
assign v3732cdc = hbusreq8_p & v3777988 | !hbusreq8_p & v3a64d96;
assign v3a5f05e = hmaster1_p & v372673d | !hmaster1_p & v38076bb;
assign v376e7e4 = hbusreq5 & v3769a00 | !hbusreq5 & !v8455ab;
assign v37408a1 = jx0_p & v3a5a2a4 | !jx0_p & v3729eb8;
assign v37427f8 = hbusreq4 & v3a715d2 | !hbusreq4 & v8455ab;
assign v3a63299 = hlock4 & v37681ed | !hlock4 & v375e0e3;
assign v3754c09 = hgrant5_p & v8455ab | !hgrant5_p & v3a69ed4;
assign v377c2ac = hbusreq1 & v377395f | !hbusreq1 & v8455ab;
assign v376382c = hbusreq0 & v375f504 | !hbusreq0 & v376fa94;
assign v3761006 = hlock4 & v3730451 | !hlock4 & v37590cb;
assign v3752d7a = hgrant7_p & v3741cd4 | !hgrant7_p & v37676b6;
assign v372e3f5 = hlock0 & v3a70b92 | !hlock0 & v375491e;
assign v3a5605f = hmaster0_p & adf78a | !hmaster0_p & v3a70666;
assign v373b0b2 = hmaster1_p & v37736b4 | !hmaster1_p & v3a715cd;
assign v3809e5c = hlock1_p & v376b5ac | !hlock1_p & v37547c9;
assign v3577484 = hmaster0_p & v374bddc | !hmaster0_p & v23fe0c9;
assign v3a6e9fc = hbusreq8 & v8455e7 | !hbusreq8 & v3737700;
assign v3a6fca5 = hgrant3_p & v372f657 | !hgrant3_p & v376a1d7;
assign v37737f9 = hbusreq0_p & v3a5ad13 | !hbusreq0_p & v375d8fb;
assign v377ac1e = hmaster0_p & v37482c7 | !hmaster0_p & v376a6f1;
assign v3736fb1 = jx0_p & v377eed2 | !jx0_p & v3a5803d;
assign v37433b4 = hbusreq2_p & v37797ef | !hbusreq2_p & v372f72b;
assign v3738e3c = hmaster0_p & v3a6f025 | !hmaster0_p & v8d4314;
assign v3a584fd = hmaster0_p & v3807aa1 | !hmaster0_p & v3777cb2;
assign v3778da6 = hbusreq0 & v375ec0b | !hbusreq0 & v3a5acd5;
assign v3a70fa5 = locked_p & v374ee47 | !locked_p & v8455ab;
assign v37422b5 = hlock4_p & v3a70530 | !hlock4_p & !v8455ab;
assign ac69a2 = hbusreq8_p & v373f1ba | !hbusreq8_p & v3a5f1db;
assign v3759842 = hbusreq3_p & v3761181 | !hbusreq3_p & !v8455ab;
assign v376d872 = hgrant5_p & v377dc72 | !hgrant5_p & v3766ed8;
assign v3a6fb3e = hmaster1_p & v374729b | !hmaster1_p & v38097ae;
assign v3a6a435 = hbusreq4_p & v374f677 | !hbusreq4_p & v377b734;
assign v3a70c1d = hmaster1_p & v377380a | !hmaster1_p & !v372bc46;
assign v376d522 = hmaster1_p & v3741d24 | !hmaster1_p & v374122a;
assign v3a58e7f = hgrant6_p & v37517d2 | !hgrant6_p & !v372599c;
assign v3a6c0f1 = hlock6_p & v35b9d52 | !hlock6_p & v3a6ac26;
assign v375c769 = hmaster2_p & v8455ab | !hmaster2_p & v374109e;
assign v3808e3a = hbusreq7 & v37444e7 | !hbusreq7 & v3734279;
assign v3732797 = hgrant6_p & v8455ab | !hgrant6_p & v3a61886;
assign v377d045 = hgrant4_p & v8455ab | !hgrant4_p & v3a5cb6f;
assign v3a66940 = hgrant7_p & v377f7dd | !hgrant7_p & v376513f;
assign v373f1e4 = hgrant2_p & v8455ab | !hgrant2_p & v3751ad8;
assign v3a6f838 = hmaster0_p & v3745181 | !hmaster0_p & v3a6f700;
assign v3a587d6 = hmaster0_p & v3a70030 | !hmaster0_p & v372f260;
assign v375c697 = hbusreq4_p & v1e378da | !hbusreq4_p & v8455ab;
assign v3771f9b = hbusreq6 & v2619b43 | !hbusreq6 & v37443ab;
assign v3763952 = hgrant5_p & v376fe0c | !hgrant5_p & v3a64f54;
assign v377e67a = hlock8 & v3a70662 | !hlock8 & v3743f2c;
assign v3a6eb2e = stateG2_p & v8455ab | !stateG2_p & v3a6e78d;
assign v374dc6d = hlock4_p & v37652a5 | !hlock4_p & v8455b3;
assign v3744835 = hbusreq4_p & v3767561 | !hbusreq4_p & v373f836;
assign v3a70c10 = hbusreq4 & v3a62c49 | !hbusreq4 & v3809ec3;
assign v3a6af5b = hlock8 & v3764955 | !hlock8 & v37408b7;
assign v373913e = hlock2_p & v20d166d | !hlock2_p & v8455ab;
assign ce4d7a = hmaster2_p & v3755dcd | !hmaster2_p & v8455ab;
assign v374f820 = hmaster2_p & v3723211 | !hmaster2_p & v3a71293;
assign v3a5d09b = hmaster2_p & v374b5b6 | !hmaster2_p & v8455ab;
assign v374e55d = hgrant5_p & v37677e2 | !hgrant5_p & v3a6f7a3;
assign v374df63 = hmaster2_p & v3a69444 | !hmaster2_p & v3a54b63;
assign v374875d = hlock6 & v3a714d2 | !hlock6 & v37618ad;
assign v3a6ff5c = hgrant2_p & v3a6b3df | !hgrant2_p & v37693cf;
assign v375a83f = hbusreq6_p & v374d2b3 | !hbusreq6_p & v39eb4a7;
assign v3a708e0 = hmaster2_p & v3768768 | !hmaster2_p & v372f3e8;
assign v37694f9 = hmaster0_p & v37765cf | !hmaster0_p & v37527dc;
assign v372f0bc = hmaster0_p & v37618bf | !hmaster0_p & v3774bdf;
assign v3732931 = hmaster2_p & v3777bd6 | !hmaster2_p & v3a701d7;
assign v3a56bb5 = hmaster1_p & v8455e7 | !hmaster1_p & v376f9ca;
assign v373b30b = hgrant4_p & v8455ab | !hgrant4_p & v376d3e1;
assign v3a71556 = hgrant5_p & v3a64b1e | !hgrant5_p & v3772d0e;
assign v3a71469 = hmaster2_p & v8455ab | !hmaster2_p & v3a56f67;
assign v373a267 = hmaster1_p & v3a6f563 | !hmaster1_p & v3a715d1;
assign v375d3cd = hgrant4_p & v3a6f7a1 | !hgrant4_p & v3a7057a;
assign v37256b3 = hbusreq7 & v3a6f371 | !hbusreq7 & v37782a8;
assign v374e606 = hgrant3_p & v8455be | !hgrant3_p & !v3755e82;
assign v3a703be = hmaster2_p & v3759ad8 | !hmaster2_p & !v37512c0;
assign v3767121 = hmaster2_p & v8455ab | !hmaster2_p & v3a679ae;
assign v3a710bd = hmaster2_p & v37624a2 | !hmaster2_p & v377ef4a;
assign v3a5f6c3 = hbusreq5 & v3a607fa | !hbusreq5 & v3a7122f;
assign v3a70b19 = hmaster0_p & v375214d | !hmaster0_p & !v8455ab;
assign v3a70baf = hbusreq5_p & v3a70f68 | !hbusreq5_p & v3770b26;
assign v375a2ac = hbusreq8 & v3777479 | !hbusreq8 & v3774608;
assign v3a6f7bc = hmaster2_p & v3a6f99b | !hmaster2_p & v3737a5a;
assign v3760bfd = hgrant6_p & v8455ab | !hgrant6_p & v3a56bf0;
assign v2acaff4 = hlock0_p & v373a391 | !hlock0_p & v8455ab;
assign v3a71228 = hbusreq4_p & v372343e | !hbusreq4_p & !v8455ab;
assign v37565d3 = hmaster1_p & v374f9cc | !hmaster1_p & v8455bd;
assign v37435a9 = hmaster2_p & v3a70809 | !hmaster2_p & v3735153;
assign v3770f3a = hbusreq3_p & v3a6f425 | !hbusreq3_p & v23fd7d9;
assign v3777705 = hlock1_p & v3775442 | !hlock1_p & v8455b0;
assign v375f423 = hlock4_p & v3a647e3 | !hlock4_p & v373acc2;
assign v3a71315 = hmaster1_p & v3a714cd | !hmaster1_p & v375134f;
assign v3729c7e = hbusreq4 & v3a70118 | !hbusreq4 & !v8455bd;
assign v377d4dd = hlock8 & v3748059 | !hlock8 & v3a6f09d;
assign v3778eed = hmaster0_p & v374314f | !hmaster0_p & v3766658;
assign v3a70f20 = hlock4_p & v3a653e4 | !hlock4_p & !v8455ab;
assign v38094e9 = hbusreq6 & v3729421 | !hbusreq6 & v8455bd;
assign v3a6fcb8 = hbusreq5_p & v373f247 | !hbusreq5_p & !v3734fa5;
assign v3735907 = hmaster2_p & v376dbdf | !hmaster2_p & v3a696ed;
assign v37395a4 = hlock0_p & v20d166d | !hlock0_p & v8455ab;
assign v3a67e53 = hlock0 & v3725799 | !hlock0 & v373f124;
assign v3765203 = hmaster1_p & v3a635ea | !hmaster1_p & v3a5d21b;
assign v375d0cf = hgrant2_p & v3a5eadd | !hgrant2_p & v3730b5e;
assign v23fe345 = hbusreq7 & v375524c | !hbusreq7 & v374752b;
assign v3722ebc = hmaster0_p & v3a5a807 | !hmaster0_p & v3a5da8f;
assign v376d29a = hbusreq4 & v3a5cd72 | !hbusreq4 & v3a5aacb;
assign b88b06 = hmaster2_p & v8455ab | !hmaster2_p & baea86;
assign v3a65652 = hmaster0_p & v3a65174 | !hmaster0_p & v8455e7;
assign v375a086 = hmaster2_p & v3746745 | !hmaster2_p & v3771dda;
assign v375043c = hmaster2_p & v3a566eb | !hmaster2_p & v3a70464;
assign v3776c44 = hbusreq2_p & v3745451 | !hbusreq2_p & v8455ab;
assign v3a6ff0b = hbusreq8_p & v3779195 | !hbusreq8_p & v3752b90;
assign v3748ded = hmaster2_p & v3a68426 | !hmaster2_p & v8455ab;
assign v372eec5 = hgrant6_p & v372aadd | !hgrant6_p & v3a6ce42;
assign v3a5b576 = hgrant4_p & v8455ab | !hgrant4_p & v3768f5f;
assign v3726994 = jx0_p & v3a6f568 | !jx0_p & v3809e71;
assign v3766048 = hgrant5_p & v8455ab | !hgrant5_p & v3a65a52;
assign v3770ab1 = hlock4 & v37535ae | !hlock4 & v3750ef8;
assign v37247a3 = hgrant4_p & v3744ea3 | !hgrant4_p & !v376cd2f;
assign v3a60e38 = hmaster0_p & v3a6c4e4 | !hmaster0_p & v3761fda;
assign v3a70759 = hlock4_p & v3752d10 | !hlock4_p & v374b25d;
assign v3772c89 = hgrant3_p & v3a5872a | !hgrant3_p & v360d03b;
assign v3725564 = hgrant2_p & v3a6f71a | !hgrant2_p & v3a551e4;
assign v3a56a0d = hmaster1_p & v3a6f92f | !hmaster1_p & v3730c14;
assign be166e = hgrant4_p & v3a6efb6 | !hgrant4_p & v3764370;
assign v3a70104 = hbusreq4_p & v373449c | !hbusreq4_p & v375542d;
assign v3729520 = hlock8 & v3754f72 | !hlock8 & v3a70461;
assign v37416c6 = hbusreq0 & v375d288 | !hbusreq0 & v8455ab;
assign v373766f = hbusreq8 & v3a6fa99 | !hbusreq8 & v3734279;
assign v3a6f7f2 = hmaster1_p & v3758180 | !hmaster1_p & v3a70c28;
assign v375aaca = hbusreq3_p & v377ad9a | !hbusreq3_p & !v8455ab;
assign v3763e46 = hbusreq8 & v3a5e1b7 | !hbusreq8 & v376ae9f;
assign v3a68697 = hgrant4_p & v8455ab | !hgrant4_p & v3a5749f;
assign v3a5cff1 = jx0_p & v374b0eb | !jx0_p & v8455ab;
assign v3a6fcef = hgrant3_p & v375c1d1 | !hgrant3_p & v375018e;
assign v37565ce = hmaster2_p & v373339b | !hmaster2_p & v375c1d9;
assign v376dd15 = hmaster2_p & v372df82 | !hmaster2_p & v3747585;
assign v3a709c3 = hmaster0_p & v377a236 | !hmaster0_p & !b05db7;
assign v3747737 = hmaster2_p & v3a5af94 | !hmaster2_p & !v1e38224;
assign v375b9a0 = hgrant6_p & v8455ab | !hgrant6_p & v3a71458;
assign v37540e2 = hmaster1_p & v37510e5 | !hmaster1_p & v3a70eb0;
assign v3a642c5 = hmaster0_p & v375c4cb | !hmaster0_p & v3a6d897;
assign v3a713c3 = hmaster2_p & v3763fdc | !hmaster2_p & v372ab8d;
assign v39eb4ca = hbusreq4 & v3733df1 | !hbusreq4 & !v8455ab;
assign v3a555f9 = stateA1_p & v8455ab | !stateA1_p & v3727e80;
assign v377d223 = jx0_p & v3a6fd70 | !jx0_p & v8455ab;
assign v375be63 = hmaster2_p & v8455ab | !hmaster2_p & b66167;
assign v372ecad = hmaster3_p & v3a6f15a | !hmaster3_p & v8455ab;
assign v374df50 = hbusreq0 & v3755b94 | !hbusreq0 & v3a6f75e;
assign v372e798 = hbusreq6 & v3a702bc | !hbusreq6 & v3a6fdef;
assign v375ca45 = hmaster1_p & v3a70fe6 | !hmaster1_p & v37474e1;
assign v3a6ff61 = hmaster2_p & v3728c23 | !hmaster2_p & v3a71016;
assign v377ba09 = hgrant4_p & v3a6ff30 | !hgrant4_p & v376a7b2;
assign v3a71460 = hbusreq2_p & v3a714bd | !hbusreq2_p & v3753d60;
assign v3a61f83 = hbusreq5 & v3a6fa62 | !hbusreq5 & v3a6f829;
assign v377a1dd = hmaster0_p & v376cffc | !hmaster0_p & v372626a;
assign v374d8cb = hbusreq2 & v3a5923c | !hbusreq2 & v3a6a4d4;
assign v374c5c5 = hmaster2_p & v3765e03 | !hmaster2_p & v377a3da;
assign v3a624d1 = hmaster2_p & v37432cd | !hmaster2_p & v3777cfc;
assign v376ae69 = hbusreq7_p & v3a29760 | !hbusreq7_p & v3764fe1;
assign v3a6fbe2 = hbusreq2_p & v372ac3a | !hbusreq2_p & v35772a6;
assign v375767e = hgrant3_p & v3a5fb00 | !hgrant3_p & v377844d;
assign v3734200 = hbusreq8 & v959f2d | !hbusreq8 & !v3a6f4b5;
assign v3a5c90c = hbusreq6_p & v3a6f4b2 | !hbusreq6_p & v35772a6;
assign v3746138 = hmaster3_p & v374e55f | !hmaster3_p & v374ae4e;
assign v3754cf4 = hbusreq4_p & v377c2ce | !hbusreq4_p & v373fe10;
assign v3735a87 = hbusreq5_p & v37675f1 | !hbusreq5_p & v3a66e9f;
assign v3a6a1d1 = hmaster0_p & v3a6ffd3 | !hmaster0_p & v373af55;
assign v377bdbe = hbusreq3 & v374b3cf | !hbusreq3 & v8455b3;
assign v376f860 = hlock3_p & v375eef1 | !hlock3_p & !v8455ab;
assign v37299dd = hgrant6_p & v3a6f4e8 | !hgrant6_p & v3768a88;
assign v375318f = hlock2_p & v3728f64 | !hlock2_p & !v8455ab;
assign v3740b82 = hmaster2_p & v37379bb | !hmaster2_p & v373b5f0;
assign v372ef56 = hmaster0_p & v3769093 | !hmaster0_p & v3a6fc28;
assign v3a6823d = hbusreq6_p & v372a0f7 | !hbusreq6_p & !v8455ab;
assign v376dd7a = hmaster1_p & v3a58cfc | !hmaster1_p & v3a56d30;
assign v3735c95 = hbusreq6 & v3a6fa39 | !hbusreq6 & v8455ab;
assign v377fc1f = hgrant4_p & v8455ab | !hgrant4_p & v376b199;
assign v374de25 = hbusreq5 & v3738270 | !hbusreq5 & !v3745239;
assign v3757c7d = hmaster0_p & v375de43 | !hmaster0_p & !v3745704;
assign v37535ae = hbusreq4 & v3750ef8 | !hbusreq4 & v374d63f;
assign v375d10e = hgrant6_p & v372df43 | !hgrant6_p & v8455ab;
assign v3a6e9c0 = hgrant3_p & v8455e1 | !hgrant3_p & !v377ee58;
assign v376c13c = hgrant2_p & v3752a0d | !hgrant2_p & v3a70a1a;
assign v964c47 = hbusreq0_p & v374e35e | !hbusreq0_p & v8455ab;
assign v375a543 = hmaster1_p & v3a68245 | !hmaster1_p & v3a66811;
assign v3a68245 = hlock5 & v3a60755 | !hlock5 & v374c6ff;
assign v3726dfd = hmaster0_p & v37480b7 | !hmaster0_p & v3766669;
assign v3a70e76 = hbusreq5_p & v3a6eb7a | !hbusreq5_p & v3750c08;
assign v37775ce = hmaster0_p & v3758f2e | !hmaster0_p & v3747dd8;
assign bf2cd1 = hbusreq7_p & v375aa44 | !hbusreq7_p & v3a6fec5;
assign v37610f8 = hgrant2_p & v3740110 | !hgrant2_p & v3a5cc4c;
assign v3747a41 = hgrant4_p & v3a5cd53 | !hgrant4_p & v3752523;
assign v376a1c9 = hgrant5_p & v37364a3 | !hgrant5_p & v3a60b0f;
assign v377a68a = hmaster3_p & v372e440 | !hmaster3_p & v375e73a;
assign v3738006 = hbusreq0 & v3a63028 | !hbusreq0 & v8455ab;
assign v3a6fbc5 = hbusreq4 & v375d10e | !hbusreq4 & v373031f;
assign v372fb58 = hmaster2_p & v3769bdb | !hmaster2_p & !v3771c85;
assign v3756471 = hmaster1_p & v8455ab | !hmaster1_p & v3a714ef;
assign v37480ec = hbusreq0 & v3760fab | !hbusreq0 & v3a69ad3;
assign v3731389 = hgrant6_p & v374a664 | !hgrant6_p & v3a6f4dc;
assign v372eb43 = stateG10_1_p & v35772a6 | !stateG10_1_p & v372865e;
assign v3763209 = hbusreq6_p & v3747302 | !hbusreq6_p & v3a6c5ee;
assign v8455e3 = start_p & v8455ab | !start_p & !v8455ab;
assign v377e897 = hmaster2_p & v3a676d6 | !hmaster2_p & v8455e7;
assign v3776150 = hlock5_p & v377098c | !hlock5_p & v377a337;
assign v3a70df4 = hbusreq6 & v3a69544 | !hbusreq6 & v1e378b4;
assign v3737acd = hgrant2_p & v3758472 | !hgrant2_p & !v8455ab;
assign v3747429 = hbusreq7 & v3777586 | !hbusreq7 & v8455ab;
assign v374ed07 = hbusreq3 & v372f85e | !hbusreq3 & v8455ab;
assign v3773078 = hmaster0_p & v3a60a84 | !hmaster0_p & v3748b9d;
assign v3a70252 = hmaster0_p & v3a70c30 | !hmaster0_p & v372b7a3;
assign v3769b3f = hbusreq5_p & v374f345 | !hbusreq5_p & v373bac6;
assign v380913f = hmaster2_p & v3a6dc08 | !hmaster2_p & v3753329;
assign v375e099 = hmaster2_p & v3724394 | !hmaster2_p & v8455c3;
assign v376132e = hgrant2_p & v37605c1 | !hgrant2_p & v3772b2b;
assign v3742b92 = hmaster0_p & v3769093 | !hmaster0_p & v3a71439;
assign v3a6a346 = hbusreq4 & v3a6f20f | !hbusreq4 & v3a60a68;
assign v3a70e6a = hmaster2_p & v373891b | !hmaster2_p & v372a1d6;
assign v374ca8a = hmaster0_p & v374502e | !hmaster0_p & v3a6eb65;
assign v3a625ee = hlock1_p & v8455ab | !hlock1_p & v3771ce2;
assign v375a397 = hgrant4_p & v8455c2 | !hgrant4_p & v3a703b5;
assign v374aa82 = hmaster1_p & v373f042 | !hmaster1_p & v8455e7;
assign v3758e05 = hbusreq4_p & v3a58773 | !hbusreq4_p & v3749eb2;
assign v3a6212b = hgrant2_p & v37745e0 | !hgrant2_p & !v3a712e3;
assign v3a70f92 = hmaster1_p & v8455ab | !hmaster1_p & v3779bde;
assign v3756bd2 = jx1_p & v375d98f | !jx1_p & v37572eb;
assign v3a70bf6 = hmaster2_p & v3744ada | !hmaster2_p & v37350f9;
assign v377b267 = hlock8 & v372946a | !hlock8 & v375d2b1;
assign v37300e3 = hbusreq5_p & v373e587 | !hbusreq5_p & v3a70e47;
assign v373f79d = hlock6_p & v3778ac6 | !hlock6_p & v37531af;
assign v3773856 = hgrant3_p & v9aa8f3 | !hgrant3_p & v37736ad;
assign v374cb21 = hmaster0_p & v3a71182 | !hmaster0_p & !d6aeaf;
assign v3a65f32 = hlock6 & v3727807 | !hlock6 & aef673;
assign v372a4e5 = hmaster1_p & v373fa8c | !hmaster1_p & !v377cb41;
assign v3a7033b = hbusreq6 & v3a71632 | !hbusreq6 & v8455ab;
assign v3725a65 = hgrant5_p & v8455ab | !hgrant5_p & v37726bf;
assign v3724859 = hlock0 & v3a60a68 | !hlock0 & v372e88f;
assign v3a63f27 = hbusreq6 & v39a4ca8 | !hbusreq6 & v8455b5;
assign v3725371 = hmaster0_p & v375121b | !hmaster0_p & v3725e4b;
assign v3763af8 = hlock6 & v373120c | !hlock6 & v373abb7;
assign v376daac = hbusreq8_p & v3740811 | !hbusreq8_p & v37390ec;
assign v373eaee = hgrant6_p & v377b946 | !hgrant6_p & v37447e2;
assign v3766b23 = hlock7_p & v3a5445c | !hlock7_p & v3a5bcfa;
assign v3a70056 = hgrant1_p & v8455ab | !hgrant1_p & !v8455e7;
assign v372d238 = hbusreq6_p & v3769c43 | !hbusreq6_p & v39eb4a7;
assign v3a6fa13 = hmaster2_p & v37583be | !hmaster2_p & !v3a709e2;
assign v3770751 = hgrant3_p & v372ad53 | !hgrant3_p & v3a5d04e;
assign v3a65f3e = hlock0_p & v8455ab | !hlock0_p & v3724112;
assign v9bba04 = hmaster3_p & v8455ab | !hmaster3_p & v37249fe;
assign v3a713ad = hmaster0_p & v3768fb7 | !hmaster0_p & v375bdcc;
assign v3758291 = hmaster1_p & v3a6ef73 | !hmaster1_p & v3a6a64a;
assign v372437d = hmaster1_p & v3771076 | !hmaster1_p & v3742c68;
assign v3761eb6 = hgrant2_p & v3758472 | !hgrant2_p & !v3a6d219;
assign v3778a0a = hbusreq0 & v37522ea | !hbusreq0 & v376e5d2;
assign v377030a = hbusreq5_p & v3a58218 | !hbusreq5_p & v375a10d;
assign v3739d69 = hbusreq8_p & v3806f21 | !hbusreq8_p & v374f48b;
assign v3a605b5 = hbusreq6_p & v3771733 | !hbusreq6_p & v38071a9;
assign v9864a7 = jx0_p & v3a6ff0b | !jx0_p & v37419da;
assign v3a7075c = hbusreq7_p & v3a579da | !hbusreq7_p & v3a65acb;
assign v373abbb = hgrant6_p & v3a6f454 | !hgrant6_p & v23fde98;
assign v3a704a9 = hgrant6_p & v377938d | !hgrant6_p & v3778ac6;
assign v372ac19 = hmaster0_p & v3758cec | !hmaster0_p & v3a6d92f;
assign v373ea29 = hmaster2_p & v8455ab | !hmaster2_p & v3a2975f;
assign v376aa3f = hmaster2_p & v37447e9 | !hmaster2_p & v3769740;
assign v37444d4 = hmaster2_p & v3a70f53 | !hmaster2_p & v3722bca;
assign v3a55c8f = hlock5_p & v3772c95 | !hlock5_p & !v8455ab;
assign v373e0d8 = hmaster0_p & v3a70479 | !hmaster0_p & v375fb03;
assign v3730610 = hbusreq6_p & v35ba2dd | !hbusreq6_p & v3748332;
assign v37762bd = hbusreq4_p & v373f0ee | !hbusreq4_p & v3a69946;
assign v3a70fdb = hgrant4_p & v380911c | !hgrant4_p & v372f3f1;
assign v3a55482 = hbusreq6 & v3745f76 | !hbusreq6 & !v8455ab;
assign v373274f = hbusreq5 & v372d925 | !hbusreq5 & v8455bf;
assign v372a744 = hmaster0_p & v3a5d09b | !hmaster0_p & v3a71614;
assign v3a6f851 = hmaster1_p & v8455ab | !hmaster1_p & v3a2986f;
assign v39ebb7b = hmaster0_p & v373d27f | !hmaster0_p & v3a6581b;
assign v377f34a = hmaster2_p & v3a63172 | !hmaster2_p & v3758539;
assign v372fbb1 = hbusreq5_p & v3a70a82 | !hbusreq5_p & v3738a93;
assign v3806fbf = hbusreq0_p & v3773100 | !hbusreq0_p & v8455ab;
assign v3732fec = start_p & v3746bdb | !start_p & v377f384;
assign v37276eb = hbusreq0_p & v3747302 | !hbusreq0_p & v37496fa;
assign v37419a9 = hlock1_p & v8455ab | !hlock1_p & v3a6ab5f;
assign v3a688f9 = hbusreq7_p & v3a7064c | !hbusreq7_p & !v3755fd4;
assign v3a56130 = hbusreq5_p & v37664c5 | !hbusreq5_p & !v8455ab;
assign v3750f77 = hbusreq5_p & ca2eb2 | !hbusreq5_p & v3a60d50;
assign v372ddf8 = hmaster2_p & v3775eee | !hmaster2_p & v3a600f3;
assign v3755a0f = hlock2 & v37370f8 | !hlock2 & v3a67eec;
assign v3726f97 = hgrant0_p & v3a56ccf | !hgrant0_p & v376e611;
assign v37666bd = hbusreq2 & v3733383 | !hbusreq2 & v8455ab;
assign v375ee68 = hmaster0_p & v374b8fa | !hmaster0_p & v376afb3;
assign v3776b2a = hbusreq0 & v372dd09 | !hbusreq0 & v8455ab;
assign v37621ee = hbusreq1_p & v3758225 | !hbusreq1_p & v375c707;
assign v3777bde = hgrant4_p & v3726f57 | !hgrant4_p & v3255b23;
assign v375ece3 = hbusreq7_p & v3a6cce9 | !hbusreq7_p & v3a550e2;
assign v375d651 = stateG10_1_p & v8455ab | !stateG10_1_p & !v3a5ce2f;
assign v376c4f9 = hbusreq0 & v9fa0b5 | !hbusreq0 & v3751dd7;
assign v3a60b96 = hlock0 & v37519ea | !hlock0 & v3a6dc38;
assign v373d245 = hbusreq5_p & v374c007 | !hbusreq5_p & v372b31a;
assign v3727a6d = hmaster1_p & v3a635ea | !hmaster1_p & v3758b8b;
assign v376b2ab = hmaster0_p & v8a21c4 | !hmaster0_p & v3737721;
assign v9aa32c = hmaster1_p & v3a635ea | !hmaster1_p & v37692dc;
assign v377bdd1 = hmaster1_p & v3a70ea5 | !hmaster1_p & v3a6c38a;
assign v375f87a = hmaster0_p & v372abac | !hmaster0_p & v3750b22;
assign v3756c2e = hbusreq5_p & v372b8da | !hbusreq5_p & v374c9ab;
assign v3731800 = hbusreq8 & v3a6f518 | !hbusreq8 & v375d113;
assign v374c23f = hlock5_p & v377e2b3 | !hlock5_p & v3725a73;
assign v37353c0 = hgrant1_p & v3a70e9a | !hgrant1_p & v37665bf;
assign v3731991 = hbusreq3_p & v3742feb | !hbusreq3_p & v8455ab;
assign v3a70427 = hmaster0_p & v3755002 | !hmaster0_p & v37362ff;
assign v3758ef5 = hgrant1_p & v3a6ec0d | !hgrant1_p & !v8455ab;
assign v3a5a814 = hbusreq8_p & v3a6f7b8 | !hbusreq8_p & v3725688;
assign v37476d9 = hbusreq7 & v372a965 | !hbusreq7 & v375e6fc;
assign v3770a82 = hmaster2_p & v3764881 | !hmaster2_p & !v3766ff7;
assign v3761b5e = hbusreq4_p & v377b24b | !hbusreq4_p & v374b27d;
assign v373d64d = hbusreq7 & v3a5965e | !hbusreq7 & v38064a3;
assign v3765739 = hgrant6_p & v3726bff | !hgrant6_p & v33790e7;
assign v3a70dd0 = hbusreq3 & a9f66a | !hbusreq3 & v375da10;
assign v373d25a = hbusreq7 & v3a53392 | !hbusreq7 & v3749f3b;
assign v3750d09 = hgrant6_p & v377f09a | !hgrant6_p & v372d279;
assign v3a5d4ac = hmaster2_p & v3a6fe4e | !hmaster2_p & v37588a3;
assign v3a66bc6 = hmaster0_p & v8455b0 | !hmaster0_p & v3779f51;
assign v3a68c32 = hbusreq6_p & v3a6f744 | !hbusreq6_p & v3760bd6;
assign v3a60030 = hlock7_p & v3807072 | !hlock7_p & v375fc56;
assign v3a553db = hmaster2_p & v372d435 | !hmaster2_p & v373574c;
assign v3a5a01b = hbusreq6_p & v3a67f8e | !hbusreq6_p & v8455ab;
assign v37262fd = hlock0_p & v3a6f43e | !hlock0_p & v372935c;
assign v374f20c = hbusreq3 & v3775303 | !hbusreq3 & v8455ab;
assign v374ffc1 = hmaster0_p & v377ce1a | !hmaster0_p & v376c85c;
assign v3757ee7 = hbusreq5 & v3742e40 | !hbusreq5 & v8455ab;
assign v1e38260 = hmaster2_p & v3a687be | !hmaster2_p & v377928c;
assign hgrant5 = !v360ba91;
assign v3a6f17b = hlock4 & v3a61a71 | !hlock4 & v3774f4e;
assign v377040f = hmaster2_p & v8455ab | !hmaster2_p & v3758c50;
assign v3a70829 = hlock0_p & v376430b | !hlock0_p & v8455ab;
assign v3a68317 = hbusreq5_p & v3728343 | !hbusreq5_p & v375f742;
assign v3723a2d = hmaster2_p & v8455ab | !hmaster2_p & v37630f1;
assign v376bb27 = hgrant2_p & v8455ab | !hgrant2_p & v3765351;
assign v3735f14 = hlock0_p & v375039e | !hlock0_p & v37277c2;
assign v373083d = jx0_p & v374ce46 | !jx0_p & v373e5f3;
assign v3a644cd = hlock6_p & v3759158 | !hlock6_p & v377b576;
assign v375523d = hmaster0_p & v377bb0e | !hmaster0_p & v3a66292;
assign v3a627a8 = jx2_p & v3a5f8b6 | !jx2_p & v3773613;
assign v3a5d590 = hmaster0_p & v35b77ec | !hmaster0_p & v3a6f3a2;
assign v376bf10 = hbusreq2_p & v39a4e8f | !hbusreq2_p & v37491b7;
assign v375c01d = hgrant3_p & v8455ab | !hgrant3_p & !v376f38d;
assign v3a6f45b = hmaster2_p & v376b4e1 | !hmaster2_p & !v3a5f83e;
assign v3727141 = hmaster2_p & v3a6fe6a | !hmaster2_p & !v3740df7;
assign v375b80e = hlock0_p & v374c936 | !hlock0_p & v1e37ca9;
assign v3a70630 = hmaster2_p & v3a6f8de | !hmaster2_p & v3a5a158;
assign v3a574bf = hbusreq5_p & v375cd8c | !hbusreq5_p & !v3a64b9b;
assign v3a5cf78 = hgrant6_p & v3a5e7c0 | !hgrant6_p & v37375f3;
assign v3a6f8bd = hmaster0_p & v3a712c2 | !hmaster0_p & v3747824;
assign v3a6fc28 = hmaster2_p & v3769093 | !hmaster2_p & v3a6a8ee;
assign v3772567 = hbusreq4 & v3754b98 | !hbusreq4 & v3749d78;
assign v3748126 = hbusreq7 & v377dc20 | !hbusreq7 & !v3723583;
assign v3a6f932 = hbusreq5 & v377d107 | !hbusreq5 & v3742cd4;
assign v372f93c = hmaster0_p & v375ec4e | !hmaster0_p & v8455ab;
assign v372cfec = hlock2_p & v3a70ad2 | !hlock2_p & !v3a712a8;
assign v376887c = hlock1_p & v3738eb6 | !hlock1_p & !v8455ab;
assign v3a64e18 = hbusreq7 & v3763d2c | !hbusreq7 & v374a289;
assign v3a70566 = hgrant6_p & v3a64045 | !hgrant6_p & v3a637ca;
assign v374429f = hgrant2_p & v8455ab | !hgrant2_p & v3a70232;
assign v377dc60 = hlock5 & v3a5e618 | !hlock5 & v376dc6f;
assign v37376dd = hbusreq8 & v374e55d | !hbusreq8 & v8455ab;
assign v3a70dfa = hmaster1_p & v3762e13 | !hmaster1_p & v37486e9;
assign v3745ab5 = hmaster0_p & v37566b2 | !hmaster0_p & v3727af8;
assign v372df9a = hbusreq3_p & v3a5f4b2 | !hbusreq3_p & !v8455ab;
assign v374d926 = hmaster2_p & v374f178 | !hmaster2_p & v3a71455;
assign v3806ec9 = hmaster1_p & v37677b4 | !hmaster1_p & v3a6f33e;
assign v3a70e5b = hgrant6_p & v375987e | !hgrant6_p & v8455ab;
assign v372f1b9 = hlock0 & v3a6f044 | !hlock0 & v3758915;
assign v3749d1d = stateA1_p & v8455ab | !stateA1_p & !v8455ff;
assign v376b5c6 = hbusreq6_p & v374b1ea | !hbusreq6_p & v372bbb3;
assign v375e261 = hbusreq6 & aab2b0 | !hbusreq6 & v8455e7;
assign v37264cb = hmaster0_p & v3763f95 | !hmaster0_p & v3a61cb5;
assign v3778c61 = hmaster2_p & v20930c6 | !hmaster2_p & v3779e95;
assign v3a6eb81 = stateG10_1_p & v8455ab | !stateG10_1_p & !v3a6eb45;
assign v373a9fb = hmaster2_p & v3740d3b | !hmaster2_p & v375c903;
assign v375a6e8 = hbusreq5 & v3722a46 | !hbusreq5 & v28896f0;
assign v377bfc0 = hbusreq2_p & v37496fa | !hbusreq2_p & v3743b9e;
assign v3a6d792 = hbusreq5 & v3a642c5 | !hbusreq5 & v375e512;
assign v3a6d3f3 = hlock2 & v3752c29 | !hlock2 & v3766e5d;
assign v3a5b3f9 = hbusreq8_p & v39a4eaa | !hbusreq8_p & v376f24b;
assign v3a56827 = hbusreq5 & v3a556df | !hbusreq5 & v37476b8;
assign v377ce51 = hgrant2_p & v3731cc3 | !hgrant2_p & v8455ab;
assign v3a6f379 = hmaster2_p & v37773a0 | !hmaster2_p & v3a66822;
assign v3a705a8 = hgrant4_p & v374378e | !hgrant4_p & v3a71474;
assign v33789ef = hmaster0_p & v3733ba7 | !hmaster0_p & v3a6ddea;
assign v375d351 = hgrant5_p & v3a6cbfa | !hgrant5_p & v3a71043;
assign v3742303 = hmaster0_p & v3a635ea | !hmaster0_p & v373d993;
assign v3a6cb96 = hbusreq5_p & v374e5ad | !hbusreq5_p & v372b72d;
assign v3a6fd84 = hbusreq5 & v3759c96 | !hbusreq5 & !v3a715ba;
assign v3743bbe = hgrant4_p & v377c94b | !hgrant4_p & v3a66999;
assign v3a711a9 = hgrant0_p & v8455ab | !hgrant0_p & v3746e79;
assign v3a6fb71 = hbusreq6 & v372383a | !hbusreq6 & v8455ab;
assign v3a6f7c6 = hbusreq7 & v3731f7f | !hbusreq7 & v3a6ec0f;
assign v3765b3c = hmaster2_p & v3767b70 | !hmaster2_p & v375981e;
assign v3a5d365 = hmaster2_p & v373a822 | !hmaster2_p & v3735272;
assign v3a5e496 = hmaster0_p & v3725710 | !hmaster0_p & v373c3a0;
assign v3a6199d = hbusreq6 & v3a6224d | !hbusreq6 & v373b11b;
assign v3737721 = hmaster2_p & v3a58b1f | !hmaster2_p & v373e49f;
assign v3a5a9b3 = hbusreq7_p & v3a6aa9e | !hbusreq7_p & v3743e90;
assign c4d24d = hbusreq5_p & v8455ab | !hbusreq5_p & v373df1f;
assign v3768e37 = hlock8_p & v3a712d5 | !hlock8_p & v3733c7f;
assign v3738f37 = hgrant5_p & v3a713bf | !hgrant5_p & v372a738;
assign v376c687 = hbusreq0 & v3777e0a | !hbusreq0 & v372d967;
assign v373dee7 = hbusreq7_p & v3773940 | !hbusreq7_p & v3764bee;
assign v3731839 = hmaster0_p & v37688bf | !hmaster0_p & v8455ab;
assign v3a7057a = hbusreq4_p & v3772541 | !hbusreq4_p & v3774a1e;
assign v375da52 = hbusreq7 & v377afb7 | !hbusreq7 & v3a572bd;
assign v37567db = hmaster2_p & v8455ab | !hmaster2_p & !v374d648;
assign v3a70ea0 = hbusreq3 & v3760e47 | !hbusreq3 & v37427d3;
assign v3a6505b = hbusreq3_p & v3a6f9ca | !hbusreq3_p & v3725994;
assign v3a6fd86 = jx0_p & v3761497 | !jx0_p & v8455ab;
assign v3758d3f = hbusreq4_p & v375e657 | !hbusreq4_p & !v3a69591;
assign v375a3a8 = hlock0 & v3a635ea | !hlock0 & v3725671;
assign v37423c1 = hbusreq7_p & v3734279 | !hbusreq7_p & v3736779;
assign v372911f = hmaster2_p & v377204f | !hmaster2_p & v3756304;
assign v3750c08 = hmaster0_p & v3757b16 | !hmaster0_p & v23fe217;
assign v3726d94 = hmaster2_p & v8455e7 | !hmaster2_p & v3731859;
assign v3731e50 = hbusreq5 & v3a65911 | !hbusreq5 & v3722fe6;
assign v37490cb = hlock0_p & v376a14f | !hlock0_p & v3763175;
assign v3a5936a = hbusreq5 & v373257d | !hbusreq5 & v37452e7;
assign v3807604 = hbusreq0 & v376a715 | !hbusreq0 & v8455ab;
assign v376c07e = hmaster1_p & v3771646 | !hmaster1_p & !v372e1b6;
assign v3734982 = hmaster2_p & v3730627 | !hmaster2_p & v3a6a261;
assign v3768589 = hgrant4_p & v8455ab | !hgrant4_p & v3a71188;
assign v37412c3 = hbusreq6_p & v373d293 | !hbusreq6_p & v377ab46;
assign v3a6fc7d = hbusreq4_p & v372b6ec | !hbusreq4_p & v8455ab;
assign v3a690c2 = hgrant6_p & v3759e3c | !hgrant6_p & v3a6fdb4;
assign v3778b2a = hmaster1_p & v3735b5a | !hmaster1_p & v3727a10;
assign v376d28f = hgrant0_p & v3a5c945 | !hgrant0_p & v3768ce2;
assign v377b221 = hgrant8_p & v8455bd | !hgrant8_p & v376858c;
assign v3a7159f = hmaster1_p & v3a61a7f | !hmaster1_p & v3a6de83;
assign v3a707d1 = hbusreq3 & v3a5f0cf | !hbusreq3 & v8455ab;
assign v3a6f43b = hlock5_p & v373c916 | !hlock5_p & v8455ab;
assign v3a70030 = hmaster2_p & v3a70374 | !hmaster2_p & v3a6f3e7;
assign v37510d0 = hgrant5_p & v377f630 | !hgrant5_p & !v375ab89;
assign v3a7085e = hmaster2_p & v3a5fc34 | !hmaster2_p & v37541ff;
assign v3a6ef49 = hgrant2_p & v35b8d36 | !hgrant2_p & v3759fe0;
assign v8f6518 = hbusreq4 & v3724621 | !hbusreq4 & v8455ab;
assign v374bff0 = hbusreq5 & v3a61462 | !hbusreq5 & v374c23f;
assign v3a70ee5 = hbusreq4 & v3a713cc | !hbusreq4 & v3a6268c;
assign v3a71135 = hmaster2_p & v3a635ea | !hmaster2_p & v372e83f;
assign v3a6f88b = hbusreq4 & v3735d39 | !hbusreq4 & v3a6fdef;
assign v3730c14 = hmaster0_p & v3a6f92f | !hmaster0_p & v3a6f3f5;
assign v373cc48 = hmaster3_p & v3a5db7b | !hmaster3_p & v3a71650;
assign v373fad7 = hbusreq0 & v374a19d | !hbusreq0 & v8455ab;
assign v3723583 = hbusreq5_p & v377a571 | !hbusreq5_p & v8455ab;
assign d6db19 = hmaster0_p & v3a566eb | !hmaster0_p & v375043c;
assign v375a18e = hbusreq3 & v3a6ab5f | !hbusreq3 & !v2aca977;
assign v377402f = hmaster2_p & v8455ab | !hmaster2_p & v3762cca;
assign v374189f = hgrant2_p & v374306c | !hgrant2_p & v375416d;
assign v3749380 = hgrant3_p & v3a60787 | !hgrant3_p & v3a6acbb;
assign v375345f = hmaster0_p & v3745714 | !hmaster0_p & !v3a56512;
assign v374a95d = hgrant2_p & v3758fa7 | !hgrant2_p & v375978a;
assign v3725392 = hmaster2_p & v3733e9e | !hmaster2_p & v37432c6;
assign v3729ffd = hgrant3_p & v377dd3b | !hgrant3_p & !v8455ab;
assign v373dd7f = hmaster2_p & v3a5971e | !hmaster2_p & v373a3fa;
assign v3a598b7 = hgrant3_p & v8455ab | !hgrant3_p & v372bffc;
assign v373ca3d = hmaster0_p & v1e37d3a | !hmaster0_p & v3a6f2de;
assign v3a6f5ec = hbusreq8_p & v3a68228 | !hbusreq8_p & v3777340;
assign v372c151 = hgrant3_p & v8455bd | !hgrant3_p & v3738fba;
assign v3807754 = hmaster0_p & v37299de | !hmaster0_p & v3762d06;
assign v3a710cc = hmaster1_p & v23fe156 | !hmaster1_p & v3774463;
assign v3a7097d = hmaster2_p & v3743b9e | !hmaster2_p & v376bb26;
assign v3808553 = hlock0_p & v3760f87 | !hlock0_p & v3772af6;
assign v3731230 = hgrant6_p & v8455ab | !hgrant6_p & v3766e4a;
assign v33781d5 = hbusreq4 & v3a5b289 | !hbusreq4 & v8455bb;
assign v3a61604 = hlock6_p & v8455ab | !hlock6_p & !v2acb5a2;
assign v3754025 = hbusreq5_p & v3747de2 | !hbusreq5_p & d03df7;
assign v3733d66 = hmaster1_p & v3a7066c | !hmaster1_p & v374764e;
assign v3a66c12 = hbusreq5 & v3a6f610 | !hbusreq5 & v374e4fa;
assign v37445e6 = hbusreq7_p & v3a6fcf1 | !hbusreq7_p & v2925cef;
assign v3a6a209 = hbusreq0 & v3a5d5e7 | !hbusreq0 & v3a62e01;
assign v3a5b693 = hgrant4_p & v3a53eeb | !hgrant4_p & v3a70cdd;
assign v375024d = hlock0_p & v372dadb | !hlock0_p & v3a697f2;
assign v372e759 = hmaster0_p & v376f576 | !hmaster0_p & !v374c164;
assign v376e562 = hmaster2_p & v376111d | !hmaster2_p & !v3a70131;
assign v3a71102 = hlock0_p & v3a70f6a | !hlock0_p & v3a6f522;
assign v3754ca0 = hgrant8_p & v375f99c | !hgrant8_p & v3a70120;
assign v375b012 = hlock3_p & v3745b07 | !hlock3_p & v8455b0;
assign v3a62443 = hbusreq6 & v3a71453 | !hbusreq6 & !v8455b9;
assign v3750714 = hbusreq2 & v3768eb1 | !hbusreq2 & v8455ab;
assign v3a71415 = hbusreq4 & v3a6773a | !hbusreq4 & v35b774b;
assign v37756f8 = hgrant5_p & v372cdde | !hgrant5_p & v375c65f;
assign v3765901 = hgrant3_p & v376e500 | !hgrant3_p & v373c79c;
assign v3739698 = hmaster2_p & v37625a8 | !hmaster2_p & !v3a6a213;
assign v3a5749f = hgrant6_p & v8455ab | !hgrant6_p & v3766cd5;
assign v3768ba9 = jx1_p & v375c6f5 | !jx1_p & v3a649c2;
assign v37715d9 = hbusreq0 & v3a6ff8f | !hbusreq0 & v377cd7e;
assign v373ee80 = hlock2_p & v3a6672b | !hlock2_p & !v8455ab;
assign v3a6a867 = hgrant0_p & v8455ab | !hgrant0_p & v3735fee;
assign v3740b01 = hbusreq0 & v376e4bd | !hbusreq0 & v8455ab;
assign v3a70a21 = hmaster1_p & v23fd8b2 | !hmaster1_p & v8455ab;
assign v37615a2 = hmaster2_p & v8455ab | !hmaster2_p & v375411b;
assign v374e34d = hbusreq5 & v8455ab | !hbusreq5 & v374ca02;
assign v37482f8 = hburst1 & v373bf7c | !hburst1 & v3a6cfa7;
assign v3a60c38 = hmaster2_p & v377db88 | !hmaster2_p & v3762a49;
assign v3a6a2f3 = hbusreq4_p & v3a58d22 | !hbusreq4_p & !v373325f;
assign v375456e = hmaster0_p & v3a5d8b5 | !hmaster0_p & v379318b;
assign v374f126 = hgrant6_p & v8455ab | !hgrant6_p & v3731478;
assign v372d411 = hlock6_p & v373d825 | !hlock6_p & !v8455ab;
assign v37400d2 = hmaster2_p & v377b423 | !hmaster2_p & !v2678c97;
assign v3772afb = hmaster1_p & v8455e1 | !hmaster1_p & v372fa17;
assign v3a6fb21 = hmaster1_p & v3a6a8ee | !hmaster1_p & v3a714ab;
assign v376b290 = hmaster0_p & v8455ab | !hmaster0_p & v3a61de0;
assign v373e2aa = hmaster1_p & v377c5f8 | !hmaster1_p & v3a61d67;
assign v3743012 = hmaster1_p & v3a700d9 | !hmaster1_p & v372a27f;
assign v376574a = hbusreq0 & v3737220 | !hbusreq0 & v3a6f5e1;
assign v3a67d2f = hgrant4_p & v37286d3 | !hgrant4_p & v3a715a7;
assign v373edf3 = hmaster1_p & v3a635ea | !hmaster1_p & v38064d5;
assign v3771d4f = hbusreq0 & v373059e | !hbusreq0 & v377e11d;
assign v377f611 = hbusreq6 & v374fa0d | !hbusreq6 & v391331d;
assign v3a56eeb = hlock5_p & v8455ab | !hlock5_p & v3728650;
assign v373dc42 = hmaster1_p & v373ef10 | !hmaster1_p & v3a6f7b9;
assign v37662d7 = hmaster3_p & v3722b6f | !hmaster3_p & v375e4d9;
assign v377de41 = hlock1_p & v8455e7 | !hlock1_p & !v374d260;
assign v3a6fe31 = hmaster2_p & v3a653e4 | !hmaster2_p & !v3726139;
assign v373ee17 = hbusreq2_p & v8455e7 | !hbusreq2_p & v374f307;
assign v3a6261b = hlock4 & v374d88f | !hlock4 & d305e8;
assign v373ecae = hbusreq3 & v3a71682 | !hbusreq3 & v8455ab;
assign v3734585 = hmaster2_p & v37c3782 | !hmaster2_p & v3a65762;
assign v3a6c970 = hbusreq4_p & v3726204 | !hbusreq4_p & baccec;
assign v3771cac = hlock7_p & v37232aa | !hlock7_p & v8455b7;
assign v3a70e35 = hbusreq4 & v37282cf | !hbusreq4 & v37674c1;
assign v3a5b545 = hmaster2_p & v3a58cfc | !hmaster2_p & v376d856;
assign v373a331 = hbusreq0 & v3a5a73d | !hbusreq0 & v8455ab;
assign v375ab89 = hmaster1_p & v372625f | !hmaster1_p & v3736ad7;
assign v3a6bdd1 = hgrant6_p & v374bc10 | !hgrant6_p & v3764ca8;
assign v3a69062 = hgrant2_p & v3a6305e | !hgrant2_p & v377b086;
assign v3a713f1 = hbusreq5_p & v377bdec | !hbusreq5_p & v376daf2;
assign v3a70db6 = hbusreq4_p & v3a7163f | !hbusreq4_p & v373bd6c;
assign v3a70a58 = hbusreq8 & v3777e59 | !hbusreq8 & v3778211;
assign v3a709f3 = hbusreq4 & v3748cce | !hbusreq4 & v8455ab;
assign v3727482 = hbusreq2_p & v3741a9b | !hbusreq2_p & v3a7006b;
assign v37232aa = hmaster1_p & v3a64355 | !hmaster1_p & v3a5844c;
assign v373cd16 = hbusreq3_p & v375928d | !hbusreq3_p & v8455ab;
assign v3753e6f = hmaster0_p & v3a70bba | !hmaster0_p & v373af66;
assign v375c9bc = hbusreq5_p & v3742649 | !hbusreq5_p & v3735db2;
assign v3a6ebd8 = hbusreq8 & v373f909 | !hbusreq8 & v8455ab;
assign v3a71261 = hgrant2_p & v375ca6c | !hgrant2_p & v2aca789;
assign v37756ac = hbusreq3_p & v2092ffc | !hbusreq3_p & v37366d2;
assign v3a5ee7d = hbusreq6_p & d4de60 | !hbusreq6_p & v372b2ba;
assign v375b2e5 = hgrant1_p & v373c4e4 | !hgrant1_p & v8455e7;
assign v3a710e9 = hbusreq3_p & v3809282 | !hbusreq3_p & !v3744fa5;
assign v372dd14 = hmaster3_p & v3778a91 | !hmaster3_p & v3773430;
assign v3a620e2 = hlock1_p & v3a562ea | !hlock1_p & v8455b0;
assign v3806e34 = hlock2 & v376f7a7 | !hlock2 & v3a5fb00;
assign v3750b01 = hmaster2_p & v9af7ec | !hmaster2_p & v3774bad;
assign v3a6f4ab = hmaster1_p & v377766c | !hmaster1_p & v374abcc;
assign v376c0dc = jx1_p & v3a58dfb | !jx1_p & v3a6f212;
assign v3735461 = hbusreq6_p & v3768454 | !hbusreq6_p & !v8455ab;
assign v372d149 = hmaster2_p & v3a58cfc | !hmaster2_p & v39a537f;
assign v3a6a7e8 = hmaster1_p & v376984f | !hmaster1_p & v3a66120;
assign v3a70268 = hbusreq3_p & v374ed07 | !hbusreq3_p & v8455ab;
assign v373f11a = hmaster2_p & v3731859 | !hmaster2_p & v8455e7;
assign v3770b04 = hbusreq5_p & v3765bf4 | !hbusreq5_p & fc6f92;
assign v3a6299c = hbusreq7_p & v8455e7 | !hbusreq7_p & !v8455ab;
assign v372ccbb = hbusreq3_p & v3a61392 | !hbusreq3_p & v8455b3;
assign v372ff9a = hlock0 & v3a635ea | !hlock0 & v372c5da;
assign v375bf9a = hbusreq1_p & v3a5a452 | !hbusreq1_p & v8455ab;
assign v3a299ea = hmaster1_p & v3a6cb96 | !hmaster1_p & v8455ab;
assign v2093068 = jx2_p & v3759d98 | !jx2_p & v3773661;
assign v374734d = hbusreq4_p & v374c7f4 | !hbusreq4_p & !v3766bc8;
assign v3577376 = hgrant2_p & v3745f9b | !hgrant2_p & v3771d0f;
assign v3a6ef19 = hbusreq8_p & v3a575d5 | !hbusreq8_p & v3742de5;
assign v3a6f3b5 = hmaster3_p & v374ef97 | !hmaster3_p & v376a662;
assign v3a65934 = hbusreq1_p & v8455eb | !hbusreq1_p & v8455ab;
assign v3746905 = hmaster2_p & v2ff8cfd | !hmaster2_p & v3739c14;
assign v377b8c5 = hgrant5_p & v375bb11 | !hgrant5_p & v3a6fc57;
assign v3723c25 = hbusreq8 & v1e38291 | !hbusreq8 & v3731977;
assign v3762388 = hgrant6_p & v8455ab | !hgrant6_p & v3745b20;
assign v3752215 = hbusreq7 & v3743dce | !hbusreq7 & v3773f27;
assign v373c268 = hbusreq8_p & v3a55290 | !hbusreq8_p & v372f721;
assign v375dd29 = hgrant6_p & v209310e | !hgrant6_p & !v372dab0;
assign v3a700b5 = hbusreq2 & v376f768 | !hbusreq2 & v375da10;
assign v373e941 = hmaster0_p & v3726c61 | !hmaster0_p & v3a5be70;
assign v3768e48 = hlock1_p & v8455ab | !hlock1_p & v8455e7;
assign v377e2e2 = hbusreq2 & v37629e2 | !hbusreq2 & v8455ab;
assign v3a71409 = hgrant3_p & v3778ed4 | !hgrant3_p & !v8455ab;
assign v3761ca6 = hmaster1_p & v3a6f469 | !hmaster1_p & v3a6f78f;
assign v37508b2 = hlock0_p & v2ff9190 | !hlock0_p & v3766438;
assign v3737220 = hlock4 & b04260 | !hlock4 & v3a70514;
assign v3a5cebe = hlock6_p & v3a709e2 | !hlock6_p & v3754aa3;
assign v942053 = hbusreq4_p & v3a635ea | !hbusreq4_p & v375cf36;
assign v2ff8c78 = hburst0 & v3771ce2 | !hburst0 & v3763eaa;
assign v3a71571 = hlock1_p & v3722e5c | !hlock1_p & v35772a6;
assign v37478dd = hbusreq8_p & v375d20f | !hbusreq8_p & v376a0e6;
assign v3a71110 = hbusreq5_p & v37656f7 | !hbusreq5_p & v3a6f2fc;
assign v3a7058a = hbusreq4_p & v8f6518 | !hbusreq4_p & v8455ab;
assign v37306c2 = hbusreq0 & v37678fc | !hbusreq0 & !v8455ab;
assign v380704f = hlock3 & v377ec08 | !hlock3 & v374d59a;
assign v377e16a = hmaster2_p & v3772f85 | !hmaster2_p & v37258b7;
assign v3a6ef2a = hgrant4_p & v37449b3 | !hgrant4_p & v3a7071b;
assign v3a712f6 = hmaster2_p & v376e914 | !hmaster2_p & !v3770559;
assign v2acae91 = hbusreq3_p & v3737c2f | !hbusreq3_p & v3a71102;
assign v376bfb9 = hbusreq5 & v3a65ce7 | !hbusreq5 & v37577cd;
assign v376655b = hgrant2_p & v39a53b3 | !hgrant2_p & v3755aef;
assign v375b776 = hbusreq8_p & v376db98 | !hbusreq8_p & v3a70f40;
assign v374530a = hbusreq6_p & v375a0a1 | !hbusreq6_p & v3a62443;
assign v372c6ce = hlock5_p & v3a65652 | !hlock5_p & !v8455ab;
assign v3778323 = hgrant2_p & v8455ab | !hgrant2_p & !v37433b4;
assign v377b017 = jx0_p & v375f798 | !jx0_p & v374e788;
assign v372dd8e = stateA1_p & v8455ab | !stateA1_p & v8455e1;
assign v3726ddb = hbusreq5 & v3749658 | !hbusreq5 & !v8455ab;
assign v38097db = hgrant6_p & v8455ab | !hgrant6_p & a8afe1;
assign v376b1f6 = hlock4_p & v3775b81 | !hlock4_p & v8455ab;
assign v374f6f9 = hmaster2_p & v374fb8d | !hmaster2_p & v3725578;
assign v376c014 = hmaster0_p & v3753418 | !hmaster0_p & v3a70909;
assign v3740975 = hmaster0_p & v8455ab | !hmaster0_p & v3a71356;
assign v3806f70 = hbusreq4 & v3a6f9c3 | !hbusreq4 & v8455bf;
assign b58331 = hmaster1_p & v373732f | !hmaster1_p & v373f27d;
assign v1e37442 = hbusreq4_p & v3a715b2 | !hbusreq4_p & v3808874;
assign v372e7f8 = hbusreq4_p & v3748797 | !hbusreq4_p & v373dfb4;
assign v3a6c6ce = hmaster2_p & v3a64421 | !hmaster2_p & v373d9e0;
assign v373a5a6 = hbusreq4 & v372bf7f | !hbusreq4 & v3a64af7;
assign v3a5fc61 = hmaster2_p & v373aed4 | !hmaster2_p & v3a5f0b2;
assign v9d97fe = hmaster3_p & v373a560 | !hmaster3_p & v3742fbf;
assign v3a70126 = hlock4 & v3807513 | !hlock4 & v3a707ea;
assign v375591f = hgrant3_p & v3764d17 | !hgrant3_p & v3a6d525;
assign v3724a4b = hgrant2_p & v3742a78 | !hgrant2_p & v376de4e;
assign v3a638fb = hbusreq5_p & v2ff9190 | !hbusreq5_p & v376c902;
assign v3747280 = hmaster1_p & v3769ae2 | !hmaster1_p & v3a6f63a;
assign v3a6cdcd = hmaster1_p & v3a53c87 | !hmaster1_p & v3a68915;
assign v377eee2 = hmaster2_p & v3a70f32 | !hmaster2_p & v3760a1c;
assign v3749004 = hmaster0_p & v3748fe0 | !hmaster0_p & v372fd0a;
assign v3a68871 = hgrant5_p & v8455ab | !hgrant5_p & v377246f;
assign v3a6e708 = hmaster3_p & v8455ab | !hmaster3_p & v33789ca;
assign v3a5524c = hbusreq0 & v373bc30 | !hbusreq0 & v373bd6c;
assign v375c7b0 = hgrant8_p & v37544ab | !hgrant8_p & v376629b;
assign v37612a3 = hmaster1_p & v37286f3 | !hmaster1_p & v3742a61;
assign v3771901 = hlock7_p & v3740777 | !hlock7_p & !v3761916;
assign v3a709cf = hlock2 & v376b018 | !hlock2 & v376e316;
assign v3a67b48 = hbusreq6_p & v3748de3 | !hbusreq6_p & v3a69946;
assign v372339a = hgrant6_p & v377f7e1 | !hgrant6_p & v3a6cd0f;
assign v373d0b2 = hready & v3778528 | !hready & v3a7162d;
assign v374ca2e = hmaster1_p & v377e056 | !hmaster1_p & v3a683c6;
assign v37273d2 = hgrant4_p & v3a5f162 | !hgrant4_p & v3a6f505;
assign v377b8fb = hbusreq5_p & v376cdb7 | !hbusreq5_p & v37775ce;
assign v37626d4 = hbusreq2 & v3733b37 | !hbusreq2 & v8455ab;
assign v37609ab = hgrant4_p & v8455ab | !hgrant4_p & v3769a8e;
assign v37686ea = hmaster2_p & v3777da6 | !hmaster2_p & v3a29850;
assign v3750df3 = hbusreq4 & v373cee7 | !hbusreq4 & v3751d30;
assign v377d9fa = hbusreq8 & v3a5ee7a | !hbusreq8 & a0a219;
assign v3a6f792 = hmaster0_p & v37728b9 | !hmaster0_p & !v35b774b;
assign v3a711ea = hmaster2_p & v375139d | !hmaster2_p & v3752fbc;
assign v3749165 = hgrant5_p & v3a67af1 | !hgrant5_p & v3735fb3;
assign v3756820 = hmaster2_p & v3a709a6 | !hmaster2_p & v37560ff;
assign v3a6e5e8 = hlock0 & v3a6bf41 | !hlock0 & v3778454;
assign v377b0b0 = hmaster0_p & v3a702ee | !hmaster0_p & v3a606b0;
assign v372f6d3 = hbusreq5_p & v2925d03 | !hbusreq5_p & v377e056;
assign v3732817 = hgrant1_p & v374d836 | !hgrant1_p & d8a75b;
assign v380988c = hgrant6_p & v3a6f3aa | !hgrant6_p & v3763004;
assign v3754421 = hbusreq4 & v376e3db | !hbusreq4 & v8455ab;
assign v37521ed = hbusreq3_p & v39a537f | !hbusreq3_p & !v1e38224;
assign v3a5dfad = hlock6_p & v35772b3 | !hlock6_p & v35772a6;
assign v3a6ef38 = hlock8_p & v3a66ba8 | !hlock8_p & v37374e5;
assign v3727d00 = hlock0 & v3a67f97 | !hlock0 & v373f124;
assign v3a70e33 = hbusreq2 & v376b4e1 | !hbusreq2 & !v8455ab;
assign v372a24d = hmaster0_p & v3758fa8 | !hmaster0_p & v3751b37;
assign v3732e59 = hgrant4_p & v377ec59 | !hgrant4_p & v372ac3b;
assign v3735d9e = hmaster3_p & v376978a | !hmaster3_p & v3a61f33;
assign v372ab5a = hgrant0_p & v8455ab | !hgrant0_p & !v3735fee;
assign v3a6fe2d = hbusreq5 & v3a6ac20 | !hbusreq5 & v374e784;
assign v37716c3 = hbusreq2_p & v3a6f3ab | !hbusreq2_p & v8455ab;
assign v375bce2 = hmaster3_p & c8e1cc | !hmaster3_p & v376b1ee;
assign v375bc49 = hmaster1_p & v9bd777 | !hmaster1_p & v372d3b2;
assign v372f520 = hmaster1_p & v373013d | !hmaster1_p & v3728343;
assign v3a554c5 = hbusreq7_p & v373d449 | !hbusreq7_p & v377d521;
assign v3770a8c = hmaster0_p & v3a6ffb6 | !hmaster0_p & v3a661f1;
assign v3a6f774 = hmaster2_p & v3764276 | !hmaster2_p & !v374fb58;
assign v3750e32 = hgrant4_p & v374fb58 | !hgrant4_p & v374e314;
assign v372a068 = hgrant4_p & v8455ab | !hgrant4_p & v37711dd;
assign v373b0e5 = hlock0_p & a38ed7 | !hlock0_p & v374b3e1;
assign v372aa99 = hbusreq3_p & v377b073 | !hbusreq3_p & v377c31a;
assign v3750fc9 = hmaster0_p & v374de0d | !hmaster0_p & v3a6fd53;
assign v3a7003e = hgrant0_p & v3a6b873 | !hgrant0_p & !v3729a9f;
assign v3a68b25 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v3770af6;
assign v3a6e432 = hmaster2_p & v8455ab | !hmaster2_p & v377eaf2;
assign v3a7080a = hbusreq2_p & v3735e39 | !hbusreq2_p & !v3a6d684;
assign v3a6d840 = hlock4 & v3a646ae | !hlock4 & v372456c;
assign v3774276 = hgrant4_p & v380949b | !hgrant4_p & !v3a6f1a5;
assign v3725230 = hlock0_p & v3723430 | !hlock0_p & b9f474;
assign v376784b = hmaster0_p & v3747fdb | !hmaster0_p & v1e37cc1;
assign v3806847 = hlock5 & v3740885 | !hlock5 & v3776454;
assign v37543c2 = hgrant1_p & v3730e71 | !hgrant1_p & v37328bf;
assign v375d84e = hgrant4_p & v8455ab | !hgrant4_p & v3a70ad6;
assign v3a6fe9f = hbusreq6 & v3a70e03 | !hbusreq6 & v8455ab;
assign v3a6bedd = hmaster1_p & v3a563cf | !hmaster1_p & v3a6f6fe;
assign v3a70b60 = hbusreq0_p & v8455ab | !hbusreq0_p & v3a7168a;
assign v372e559 = hbusreq0 & v3a6512b | !hbusreq0 & v37781a8;
assign v3a53a8a = hmaster2_p & v8455ab | !hmaster2_p & v3a6f880;
assign v3779337 = hbusreq6_p & v376803b | !hbusreq6_p & v373a2f2;
assign v373e52d = hgrant4_p & v8455ab | !hgrant4_p & v376ef09;
assign v373fa8c = hmaster0_p & v372f046 | !hmaster0_p & !v3a6bc9a;
assign v3a70806 = hmaster2_p & v8455ab | !hmaster2_p & v3726139;
assign v3a5c945 = locked_p & v8455ab | !locked_p & !v3a619c0;
assign v377e04e = hbusreq7 & v374a60b | !hbusreq7 & v3768734;
assign v3735796 = hmaster2_p & v3747302 | !hmaster2_p & v37320ff;
assign v3a6ca1f = hbusreq4_p & v3a7076c | !hbusreq4_p & v8455ab;
assign v329f8b7 = hready_p & v3769759 | !hready_p & !v3730ab2;
assign v374720c = hbusreq3 & v380974c | !hbusreq3 & v8455b3;
assign v3a62959 = hbusreq7_p & v3741816 | !hbusreq7_p & v374f832;
assign v37425c0 = hlock6_p & v3a67983 | !hlock6_p & v8455b0;
assign v374c78e = hgrant4_p & v8455ab | !hgrant4_p & v3a5864f;
assign v3752e80 = jx0_p & v3738e45 | !jx0_p & v3a6fc81;
assign v376fa38 = hlock3_p & v1e38275 | !hlock3_p & v39a537f;
assign v377ceb5 = hbusreq5_p & v3775064 | !hbusreq5_p & v3a5d8a9;
assign v3729f32 = hlock6_p & v8455ab | !hlock6_p & v39a5265;
assign v37673dd = hbusreq2 & v37274c2 | !hbusreq2 & !v8455b5;
assign v3a70dde = hbusreq6_p & v3763004 | !hbusreq6_p & v3a5edcb;
assign v3a5646d = hbusreq8 & v3745cf8 | !hbusreq8 & v372d071;
assign v3773fd1 = hbusreq6 & v375ac23 | !hbusreq6 & v8455ab;
assign v3807020 = hmaster2_p & v3a71330 | !hmaster2_p & !v3a6eb6e;
assign v3a6f4f0 = hmaster2_p & v3a5a6e6 | !hmaster2_p & v3a6f4ba;
assign v373eb4d = hgrant6_p & v3741f22 | !hgrant6_p & v377cbcb;
assign v376e20f = hmaster1_p & v372d1ae | !hmaster1_p & v3a7055c;
assign v373361a = hbusreq8_p & v3a6d4f8 | !hbusreq8_p & v37654ea;
assign v3a70fcc = hbusreq7_p & v373562f | !hbusreq7_p & v3a64c6b;
assign v375c671 = hbusreq4_p & v3756f06 | !hbusreq4_p & v8455ab;
assign v3a6f054 = hgrant4_p & v3a71164 | !hgrant4_p & v3a701a5;
assign v3a679b5 = hmaster1_p & v3a5f2c0 | !hmaster1_p & !v3a6e0cc;
assign v3a6f312 = hbusreq3_p & v3a70ee7 | !hbusreq3_p & v3733d6e;
assign v3779c8d = hbusreq7_p & v3755e66 | !hbusreq7_p & !v8455ab;
assign v3773430 = jx0_p & v37632c6 | !jx0_p & v3773daf;
assign v37519cb = hmaster2_p & v3a69591 | !hmaster2_p & !v8455ab;
assign aefb3e = hbusreq3 & v37624a2 | !hbusreq3 & v3a7153a;
assign v39a4dd6 = hgrant6_p & v8455ab | !hgrant6_p & v3808fc2;
assign v3762281 = hlock6 & v3a6f659 | !hlock6 & v37574d2;
assign v3a5511c = hlock7 & v373fb42 | !hlock7 & v376592c;
assign v3a70e99 = hbusreq5 & d2afa4 | !hbusreq5 & v374bcb5;
assign v3a6abaa = hgrant0_p & v3a7081c | !hgrant0_p & v374794f;
assign v376c25b = hmaster0_p & v3a6e5f0 | !hmaster0_p & v325b59d;
assign v3774e48 = hgrant5_p & v3a67af1 | !hgrant5_p & v375780e;
assign db86c8 = hbusreq4 & v374179c | !hbusreq4 & !v3a53e0e;
assign v375bff8 = hgrant6_p & v37304b3 | !hgrant6_p & v373abdb;
assign v3a70c94 = hready & v3a70a12 | !hready & v3a635ea;
assign v3731004 = hgrant2_p & v376e041 | !hgrant2_p & v3a5ab6e;
assign v3a633ac = hgrant4_p & v3377c6a | !hgrant4_p & v3a6e8d2;
assign v374ab22 = hgrant4_p & v3738457 | !hgrant4_p & v3a6a48e;
assign v372df47 = hlock0_p & v38072fd | !hlock0_p & v3a70ef2;
assign v23fd7a9 = hmaster2_p & v3a5bf28 | !hmaster2_p & v372ba1c;
assign v374f6a4 = hmaster1_p & v3724e4b | !hmaster1_p & v377e406;
assign v377f5cb = hlock4_p & v3a5f0b2 | !hlock4_p & v3a6f8f5;
assign v373b7be = hmaster0_p & v3a57422 | !hmaster0_p & v3a68cec;
assign v3a6f078 = hmaster3_p & v8455ab | !hmaster3_p & v3737c39;
assign v372ef17 = hmaster0_p & v375fbf2 | !hmaster0_p & v3a70318;
assign v373ad7b = hgrant4_p & v3a6f43a | !hgrant4_p & v3752767;
assign v3747554 = hmaster0_p & v3a706a1 | !hmaster0_p & v3722ae9;
assign v3a6f347 = hlock4_p & v3746063 | !hlock4_p & v8455b0;
assign v372f1e9 = hbusreq5 & v37313e4 | !hbusreq5 & v3a71530;
assign v3a5d48b = hlock0_p & v377eaf2 | !hlock0_p & v37231ed;
assign v37318d7 = hgrant4_p & v3778d9d | !hgrant4_p & v375fdf5;
assign v375c600 = hmaster0_p & v3736eee | !hmaster0_p & !v3746ce0;
assign v37570b7 = hgrant1_p & v3a57445 | !hgrant1_p & v8455e7;
assign v3a5fbcb = hbusreq7 & v374c28e | !hbusreq7 & v3a60276;
assign v3a585d1 = hbusreq4 & v3a6f018 | !hbusreq4 & !v3740f3d;
assign v3725582 = hbusreq2_p & v3a558f6 | !hbusreq2_p & v3a5770d;
assign v376769a = hbusreq5_p & v37384a9 | !hbusreq5_p & v372a20d;
assign v3a6d2df = hbusreq4 & v37447e1 | !hbusreq4 & v3a703c0;
assign v3a712be = stateG3_1_p & v8455ab | !stateG3_1_p & !v845601;
assign v3808c66 = hgrant6_p & v3a6cb16 | !hgrant6_p & v373fcae;
assign v372633a = hbusreq6_p & v37308b0 | !hbusreq6_p & v3a71558;
assign v3a54497 = hgrant4_p & v3a53eeb | !hgrant4_p & v397d85e;
assign v374a08a = hgrant4_p & v3a672e5 | !hgrant4_p & v3737dad;
assign v373ffa9 = hgrant6_p & v3a62c7d | !hgrant6_p & v3a6e159;
assign v3738169 = hgrant4_p & v374e380 | !hgrant4_p & v3763668;
assign v37234d5 = hmaster1_p & v3769a00 | !hmaster1_p & !v376dce5;
assign v3723430 = hready & v8455e7 | !hready & v8455ab;
assign v3a6cdbc = hbusreq3_p & v376442b | !hbusreq3_p & !v8455ab;
assign v3a70b40 = hgrant5_p & v8455ab | !hgrant5_p & v373ec96;
assign v39eb3bd = hgrant2_p & v3a6f20d | !hgrant2_p & v3a54d84;
assign v3a7138d = hbusreq6_p & v377a343 | !hbusreq6_p & !v3777d95;
assign v3809958 = hbusreq2 & v3747704 | !hbusreq2 & v3a70688;
assign v3763046 = hlock7 & v3a6fe10 | !hlock7 & v3a70f4f;
assign v37534a4 = hgrant6_p & v3771b2c | !hgrant6_p & v3748964;
assign v37750bb = hmaster2_p & v3a5b5d3 | !hmaster2_p & !v377b6ce;
assign v3734fa9 = hlock3 & v376485c | !hlock3 & v377857d;
assign v374113f = hbusreq8_p & v3776fec | !hbusreq8_p & v375089b;
assign v3a71659 = hgrant4_p & v8455ab | !hgrant4_p & v3779412;
assign v3747a3f = hmaster2_p & v8455ab | !hmaster2_p & v3776dcd;
assign v3a70777 = hbusreq7 & v373c2e3 | !hbusreq7 & v3a7050a;
assign v3a6a536 = hmaster2_p & v3807f45 | !hmaster2_p & !v3727976;
assign v3a70eff = hbusreq0_p & v37416b5 | !hbusreq0_p & v3743b9e;
assign v98d1dc = hbusreq7 & v373859a | !hbusreq7 & v3a627a1;
assign v37345a5 = hmaster0_p & v8455ab | !hmaster0_p & !v37532c8;
assign v3a6f937 = hbusreq5_p & v3747d82 | !hbusreq5_p & v23fdc4f;
assign v3a55b93 = hbusreq2_p & v37398eb | !hbusreq2_p & v3724f7b;
assign v377efd0 = hgrant2_p & v8455ab | !hgrant2_p & !v37797ef;
assign v3a5d3f6 = hbusreq5_p & v3729933 | !hbusreq5_p & v3255b53;
assign v373c95b = hgrant2_p & v3746dd5 | !hgrant2_p & v3759d5a;
assign v35b773b = hbusreq8 & v374fe49 | !hbusreq8 & v8455bf;
assign v37720ee = hbusreq8 & v374abbf | !hbusreq8 & v8455ab;
assign v374165f = hgrant6_p & v3a635ea | !hgrant6_p & v37406ca;
assign v374d4ca = hgrant2_p & v3a709df | !hgrant2_p & v3753b7d;
assign v3722d8b = hbusreq7 & v377b7e0 | !hbusreq7 & !v3754a25;
assign v3764e69 = hmaster0_p & v37302c7 | !hmaster0_p & v3a71498;
assign v3a587be = hlock5 & v3a5b52c | !hlock5 & v3a2a0f4;
assign v3a64969 = hbusreq6 & v3a5ddea | !hbusreq6 & v372c1cf;
assign v376079e = hmaster3_p & v3a6ebda | !hmaster3_p & v8455ab;
assign v377ea59 = hgrant6_p & v3a6f18f | !hgrant6_p & v3769f0f;
assign v37291c7 = hbusreq8_p & v3a6fc07 | !hbusreq8_p & v372fef2;
assign v37770af = hmaster1_p & v3a675d9 | !hmaster1_p & v377d595;
assign v374e179 = hmaster0_p & v375316c | !hmaster0_p & v377cccb;
assign v3743dae = hbusreq6 & v3a70734 | !hbusreq6 & v3a6687c;
assign v373de47 = jx1_p & v376a2e7 | !jx1_p & v3a5aa8e;
assign v3a7139f = hbusreq0 & v3764de7 | !hbusreq0 & v3750eb8;
assign v373139d = hready_p & v3753a8a | !hready_p & v3a70111;
assign v3729eeb = hgrant4_p & v8455ab | !hgrant4_p & v372320e;
assign v377409c = hbusreq4_p & v3a5bea0 | !hbusreq4_p & v8455ab;
assign v3747d5a = hmaster0_p & v3a6f671 | !hmaster0_p & v373f2a6;
assign v1e378b4 = hbusreq2_p & v3762502 | !hbusreq2_p & v3a5bb64;
assign v380929f = hlock8_p & v376495c | !hlock8_p & b412f3;
assign v3a56eb1 = hlock0_p & v8455ab | !hlock0_p & !v3753f1a;
assign v3765121 = hmaster1_p & v373ff17 | !hmaster1_p & v3731349;
assign v3733df1 = hlock4_p & v374eb89 | !hlock4_p & !v8455ab;
assign v373ab06 = hlock5_p & v3a6eb0d | !hlock5_p & !v8455ab;
assign v372f8d3 = hlock3 & v3748797 | !hlock3 & v374cb4a;
assign v375fda5 = hbusreq7 & v377619b | !hbusreq7 & v372863f;
assign v3734dd8 = hbusreq6 & v372aa55 | !hbusreq6 & v8455ab;
assign v3731d2d = hmaster0_p & v3a709b2 | !hmaster0_p & v374e758;
assign v3a59f8c = hmaster0_p & v3779183 | !hmaster0_p & v3a5db94;
assign v374ed5a = hlock5_p & v3a6e39a | !hlock5_p & v375d152;
assign v3743cd6 = hbusreq6_p & v3756b39 | !hbusreq6_p & v3773d39;
assign v373cff4 = hbusreq0_p & v3732e1b | !hbusreq0_p & v3728e09;
assign v23fd923 = hlock3 & v3a6972b | !hlock3 & v3736028;
assign v3809f27 = hmaster2_p & v375058e | !hmaster2_p & !v3739c94;
assign v3a5acb3 = hlock5 & v3a6f528 | !hlock5 & v3776bdf;
assign v3a6f455 = hmaster0_p & v377bb3a | !hmaster0_p & v3751925;
assign v37497a5 = hgrant5_p & v3764109 | !hgrant5_p & v3808c5f;
assign v3a62986 = hgrant3_p & v8455ab | !hgrant3_p & v372f292;
assign v377bf77 = hbusreq4_p & v3747302 | !hbusreq4_p & v3a538bd;
assign v37384a6 = hbusreq5_p & v3a6f7d0 | !hbusreq5_p & v3a6fa41;
assign v373be73 = hbusreq7 & v97b684 | !hbusreq7 & v372874e;
assign v3723aa8 = hbusreq4 & v3a5e1ab | !hbusreq4 & !v3a60181;
assign v3763846 = hlock5_p & v3746c1d | !hlock5_p & v3746dbf;
assign v3a70f40 = hbusreq7_p & v2092ff6 | !hbusreq7_p & v377ab78;
assign v3a6f243 = hgrant2_p & v8455ab | !hgrant2_p & v3a606e8;
assign v3a7084e = hlock2_p & v373399e | !hlock2_p & !v8455ab;
assign v372d65f = hbusreq0_p & v3a62826 | !hbusreq0_p & v35b774b;
assign v3a59dab = hlock6 & v374ba04 | !hlock6 & v37719f2;
assign v3a5e82d = hbusreq8_p & v3a6f040 | !hbusreq8_p & v8455ab;
assign v37689b5 = hmaster2_p & v3a71330 | !hmaster2_p & !v37389d5;
assign v373b98a = hmaster2_p & v8455ab | !hmaster2_p & !v377a88e;
assign v3a6fd63 = hbusreq6 & v37383c0 | !hbusreq6 & v37470f6;
assign v3a5aa33 = hmaster0_p & a747d7 | !hmaster0_p & v3768616;
assign v376189a = stateA1_p & db20f4 | !stateA1_p & !v3a7147e;
assign v3a5fff6 = hgrant4_p & v37395e8 | !hgrant4_p & v3a5de35;
assign v373fc8a = hgrant2_p & v3a6c5ee | !hgrant2_p & v373c480;
assign v37273be = hgrant3_p & v8455ab | !hgrant3_p & v3a70dc0;
assign v3a6aa59 = hmaster2_p & v8455ab | !hmaster2_p & v3a59178;
assign v3739d51 = hbusreq1 & v3806db7 | !hbusreq1 & v8455ab;
assign v376d251 = hgrant0_p & v3a5b5d3 | !hgrant0_p & v3a2a2fa;
assign v3a6e9b8 = hgrant2_p & v8455ab | !hgrant2_p & !v37611c1;
assign v372cf2e = jx0_p & v3764331 | !jx0_p & v3a5db83;
assign v37419df = hmaster0_p & v3a6b924 | !hmaster0_p & v3a675ad;
assign v372a960 = hbusreq2 & v377b4f2 | !hbusreq2 & v3771e60;
assign v3a674c2 = hbusreq5 & v3a70961 | !hbusreq5 & v3773838;
assign v3736ded = hbusreq2_p & v377419d | !hbusreq2_p & v8455ab;
assign v3a71314 = hbusreq2_p & v374102a | !hbusreq2_p & v8455ab;
assign v377ad57 = hbusreq6_p & v372ec1c | !hbusreq6_p & v3a69487;
assign v37551c4 = hbusreq5 & v3768904 | !hbusreq5 & v3a6ac33;
assign v2ff8ee1 = hgrant7_p & v3a67f5c | !hgrant7_p & v376bded;
assign v37474e8 = hgrant2_p & v37443ab | !hgrant2_p & v3759abe;
assign v3a7038a = hbusreq5 & v3753804 | !hbusreq5 & v3a63f9a;
assign v372f22b = stateG10_1_p & v8455ab | !stateG10_1_p & v37596fd;
assign v373ec83 = hmaster1_p & v37577cd | !hmaster1_p & v372e741;
assign v3a71159 = hmaster0_p & v374048c | !hmaster0_p & v3a70666;
assign v3739bcb = hbusreq0 & v375c3eb | !hbusreq0 & v373cdd5;
assign v3725576 = hmaster1_p & v8455ab | !hmaster1_p & v23fd8a7;
assign v37706bf = hgrant6_p & v3a6ba6a | !hgrant6_p & v3764d9e;
assign v2acaee4 = hmaster1_p & v3809e90 | !hmaster1_p & v3a6e0cc;
assign v3765927 = hmaster0_p & v376285a | !hmaster0_p & v37635de;
assign v376ef4f = hgrant4_p & v8455ab | !hgrant4_p & v3753d9d;
assign v3a631b4 = hbusreq4_p & v373104a | !hbusreq4_p & v374fa4f;
assign v3a6bf04 = hmaster2_p & v3761719 | !hmaster2_p & v3731cf0;
assign v3a70190 = hgrant6_p & v373ba4a | !hgrant6_p & v3a5e1bc;
assign v376311f = hgrant6_p & v372672f | !hgrant6_p & v3769f88;
assign bbbe50 = hbusreq1_p & v377c186 | !hbusreq1_p & !v8455ab;
assign v3769be7 = hbusreq1_p & v3747956 | !hbusreq1_p & v8455ab;
assign ca11a2 = hbusreq5_p & v3a6ec0b | !hbusreq5_p & v376b6d8;
assign v3747d3c = hgrant3_p & v8455ab | !hgrant3_p & !v374d3d7;
assign v3748972 = hbusreq5 & v3a6efa1 | !hbusreq5 & v3a587d6;
assign v376acbb = hbusreq6 & v372989d | !hbusreq6 & v8455ab;
assign v3a6fbd0 = hlock6_p & v3a6ab5f | !hlock6_p & !v8455ab;
assign v3a6ffd8 = hbusreq7 & v3723459 | !hbusreq7 & v3777d70;
assign v37461ac = hbusreq0_p & v375803a | !hbusreq0_p & v375323b;
assign v3762525 = hbusreq6_p & v3a70d7a | !hbusreq6_p & v374ebd1;
assign v3a706b0 = hbusreq0_p & v3759b2f | !hbusreq0_p & v3a6f43e;
assign v3a6f684 = hlock8_p & v3a70063 | !hlock8_p & v8455ab;
assign v374abbf = hmaster1_p & v3a640d1 | !hmaster1_p & v3769ec3;
assign v37488cb = hbusreq7 & v3774f39 | !hbusreq7 & v3a299ea;
assign d03df7 = hmaster0_p & v372c9b0 | !hmaster0_p & v3a6c605;
assign v37298b9 = hbusreq6_p & v3a6ebf1 | !hbusreq6_p & !v8455ab;
assign v37324da = hbusreq5_p & v3a5936a | !hbusreq5_p & v3a68e46;
assign v3751ebd = hlock5_p & v377de29 | !hlock5_p & v3776abb;
assign v374cc2a = hlock1 & v375483e | !hlock1 & v373d0b2;
assign v374fdc8 = hbusreq7_p & v3752b6d | !hbusreq7_p & v376e66e;
assign v373bd6c = hgrant6_p & v8455ab | !hgrant6_p & v3a58102;
assign v943e48 = hbusreq2 & v3a5fb00 | !hbusreq2 & v3a6c5ee;
assign v3a715f9 = hbusreq7 & v3a712bc | !hbusreq7 & v3a6fb20;
assign v376ef3f = hlock0_p & v3a5cfdb | !hlock0_p & v3a71130;
assign v3761825 = hbusreq1 & v375444e | !hbusreq1 & v8455ab;
assign v3730e5d = hgrant2_p & v376defa | !hgrant2_p & !v38068b5;
assign v377329f = hgrant5_p & v377234d | !hgrant5_p & v373578d;
assign v3a6652b = hgrant5_p & v3724718 | !hgrant5_p & !v3724efc;
assign v3763efc = hlock2_p & v8455ab | !hlock2_p & v373e21a;
assign v3724249 = hmaster0_p & v3a6f85a | !hmaster0_p & v372c46e;
assign v3a67dd0 = hbusreq1_p & v373b7f5 | !hbusreq1_p & !v3a630ba;
assign v2925c5b = hgrant4_p & v377b6ce | !hgrant4_p & v3771360;
assign v3a6d48c = hbusreq4_p & v3a7024b | !hbusreq4_p & v376a348;
assign v3a70d90 = hgrant0_p & v37773a9 | !hgrant0_p & v373f8fb;
assign v377504f = hbusreq8_p & v3737695 | !hbusreq8_p & v3728f0a;
assign v3776a5c = hbusreq3 & v375a0ff | !hbusreq3 & v8455ab;
assign v39eb57c = hlock1_p & v3a65f15 | !hlock1_p & !v8455ab;
assign v3a6ecdd = hlock5 & v376f814 | !hlock5 & v376fe90;
assign v376abf6 = hgrant4_p & v8455ab | !hgrant4_p & v375473a;
assign v3a6f2c2 = hmaster0_p & v3767897 | !hmaster0_p & !v3a6607f;
assign c41ef0 = hmaster1_p & v3a6e5f0 | !hmaster1_p & v2acaedd;
assign v3770f46 = hbusreq3_p & v3a57f59 | !hbusreq3_p & !v3a66110;
assign v373f124 = hlock4 & v3732187 | !hlock4 & v37434ce;
assign v3a5ae8d = hmaster0_p & v3735ff7 | !hmaster0_p & v3a57106;
assign v3a702f9 = hbusreq7_p & v3a6f226 | !hbusreq7_p & v3a71664;
assign v372edf6 = hbusreq4_p & v3a6a07b | !hbusreq4_p & v8455ab;
assign v375fd99 = hmaster2_p & v377204f | !hmaster2_p & v37697a3;
assign v23fd804 = hgrant6_p & v3a598a9 | !hgrant6_p & v3a6f331;
assign v377af8e = hmaster1_p & v3a70588 | !hmaster1_p & v375f46d;
assign v373e7c0 = hbusreq6_p & v375135a | !hbusreq6_p & v3a70c02;
assign v3a5ff46 = hbusreq4_p & v3747302 | !hbusreq4_p & v377bfc0;
assign v3a6d3bc = hbusreq8 & v3a7074c | !hbusreq8 & v8455ab;
assign v3a63a21 = hmaster2_p & v374d8ac | !hmaster2_p & v3a7058a;
assign v37538f5 = hlock2_p & v3736913 | !hlock2_p & v8455b0;
assign v23fd9cb = hbusreq7 & v373d239 | !hbusreq7 & v3a60276;
assign v3a61397 = hgrant4_p & v8455ab | !hgrant4_p & v376a65a;
assign v374acbe = hbusreq3_p & v3747302 | !hbusreq3_p & v3a70a88;
assign v3a6094a = hmaster1_p & v8455ab | !hmaster1_p & v91ebb9;
assign v372c051 = hmaster0_p & v37579b8 | !hmaster0_p & !v3776f07;
assign v3752000 = hbusreq2_p & v373014d | !hbusreq2_p & v3a5689e;
assign v3754e78 = hbusreq6_p & v3a5dc35 | !hbusreq6_p & v3743b9e;
assign v3755bbd = hbusreq6 & v3768c2a | !hbusreq6 & v8455ab;
assign v3731bc8 = hbusreq6_p & v377d4a6 | !hbusreq6_p & v8455ab;
assign v39a4d88 = hlock0_p & v3a6f7bf | !hlock0_p & v3751734;
assign v372c565 = hbusreq3 & v37269f4 | !hbusreq3 & v3773ee6;
assign v3a6eb29 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v3a56cdc;
assign v377b49d = hgrant2_p & v3a5f50e | !hgrant2_p & v3a6ca82;
assign v374ceec = hmastlock_p & v3a70a28 | !hmastlock_p & v8455ab;
assign v372fb1b = hbusreq6_p & v37625a8 | !hbusreq6_p & !v2092faa;
assign v3a71582 = hbusreq6 & v372310a | !hbusreq6 & v37496fa;
assign v3a6774e = hbusreq4 & v3a5dc35 | !hbusreq4 & v376f2a7;
assign v3769e4c = hbusreq4 & v3a6fd6a | !hbusreq4 & v1e378b4;
assign v2092f1b = hbusreq8 & v3757fa5 | !hbusreq8 & v38067bb;
assign v374cb24 = hlock5_p & v3a70d07 | !hlock5_p & v3a698ed;
assign v3a71188 = hgrant6_p & v8455ab | !hgrant6_p & v372cb42;
assign v375d102 = hbusreq7 & v3732926 | !hbusreq7 & v3a7129d;
assign v3745315 = hmaster0_p & v3a5e24e | !hmaster0_p & v3776e2b;
assign v8455f1 = hgrant4_p & v8455ab | !hgrant4_p & !v8455ab;
assign v3a6b62d = hgrant6_p & v8455ca | !hgrant6_p & v92141c;
assign v372c3df = hbusreq1_p & v37351bc | !hbusreq1_p & v8455ab;
assign v37690db = stateG2_p & v8455ab | !stateG2_p & v377f108;
assign v3779883 = hmaster0_p & v3a6f92f | !hmaster0_p & v376f6e4;
assign v3745149 = hgrant3_p & v372e48a | !hgrant3_p & !v3a70eec;
assign v3750d61 = hbusreq4_p & v3a5e2e1 | !hbusreq4_p & cecaa5;
assign v3a55e8e = hbusreq2 & v3751734 | !hbusreq2 & v8455ab;
assign v37319d5 = hgrant6_p & v375b912 | !hgrant6_p & v3a70065;
assign b77306 = hmaster0_p & v3733083 | !hmaster0_p & v3a68426;
assign v3734c26 = hbusreq3 & v3806507 | !hbusreq3 & v376d327;
assign v373d34e = hgrant0_p & v3808c39 | !hgrant0_p & a12203;
assign v3747bc9 = hmaster2_p & v3750d37 | !hmaster2_p & !v8455ab;
assign v3a6cf5d = hbusreq2 & v372efbe | !hbusreq2 & v1e3755f;
assign v23fda38 = hbusreq0 & v3a63abb | !hbusreq0 & !v3a70028;
assign v3730d52 = hmaster3_p & v37377f0 | !hmaster3_p & v37760b8;
assign v3a6fac2 = hbusreq4_p & v3a57f59 | !hbusreq4_p & !v3a66110;
assign v37600e9 = hlock0 & v3a635ea | !hlock0 & v375a38e;
assign v377aa2e = hbusreq4 & v3728e09 | !hbusreq4 & !v8455ab;
assign v377eb45 = hbusreq4_p & v37c02a9 | !hbusreq4_p & v372dd0c;
assign v3778484 = hmaster0_p & v3738b4c | !hmaster0_p & v3a710c3;
assign v37623dd = hbusreq6_p & v3a6f9e3 | !hbusreq6_p & v8455ab;
assign v3767d55 = hgrant4_p & v376e914 | !hgrant4_p & !v3a5ef3e;
assign v372b2ef = hmaster2_p & v3739be4 | !hmaster2_p & v3746be0;
assign v1e38305 = hmaster2_p & v8455ab | !hmaster2_p & !v374fa21;
assign v3809d6a = hbusreq6_p & v374d2b3 | !hbusreq6_p & v372bbb3;
assign v3a6fc5c = hbusreq8 & v373d49c | !hbusreq8 & v3a5575e;
assign v37502d4 = hlock2_p & v3733f1c | !hlock2_p & v3a5f292;
assign v3a70e6f = hgrant2_p & v373df0d | !hgrant2_p & v373a181;
assign v3774a13 = hbusreq3 & v2619ae8 | !hbusreq3 & v8455ab;
assign v3806ff6 = hbusreq0 & v37550d4 | !hbusreq0 & v37317f1;
assign v372893a = hlock5_p & v3a606a0 | !hlock5_p & v3746cc1;
assign v37626a9 = hmaster1_p & v372bdc2 | !hmaster1_p & v3743b66;
assign v375d388 = hbusreq8 & c41ef0 | !hbusreq8 & v3a6fde6;
assign v3750f4b = hgrant3_p & v38070c1 | !hgrant3_p & v377bbd1;
assign v3a6fd36 = hmaster1_p & v377e089 | !hmaster1_p & v3a65c31;
assign v37326a0 = hbusreq4_p & v37529d9 | !hbusreq4_p & v8455ab;
assign v3744b27 = hbusreq2_p & v376ef42 | !hbusreq2_p & v1e38224;
assign v3756cea = hbusreq7_p & v3a6fe1c | !hbusreq7_p & v3a70dba;
assign v375460c = hbusreq4_p & v374999b | !hbusreq4_p & v3a6556a;
assign v373930f = hmaster0_p & v3727fcb | !hmaster0_p & v3742851;
assign v3746cbf = hmaster2_p & v375d616 | !hmaster2_p & v375070c;
assign v3a6358e = hlock0 & v3809ec3 | !hlock0 & v3a645b4;
assign v376a094 = hmaster2_p & v3a6f21c | !hmaster2_p & v376d143;
assign v3a5770d = hlock2 & v3775d56 | !hlock2 & v3a6fdc5;
assign v37533ea = hbusreq6_p & v3731004 | !hbusreq6_p & v3a6ed79;
assign v3a7023d = hgrant5_p & v3a62a2d | !hgrant5_p & v373da1b;
assign v3a671f2 = hmaster1_p & v3a61a7f | !hmaster1_p & v3730c96;
assign v3723485 = hmaster2_p & v3a5dfe8 | !hmaster2_p & v3728d9c;
assign v3a5a824 = hlock3_p & v37317ba | !hlock3_p & v3a706b1;
assign v375c718 = hgrant6_p & v37331af | !hgrant6_p & v3a62348;
assign v374b526 = hgrant4_p & v3a6f4c7 | !hgrant4_p & v372efb4;
assign v3737bd8 = hbusreq7_p & v377ecec | !hbusreq7_p & v375fe2b;
assign v374d0e3 = hbusreq6_p & v375da10 | !hbusreq6_p & v376bb26;
assign v3a7133b = hgrant6_p & v8455ab | !hgrant6_p & !v3755a2f;
assign v37487f7 = hbusreq4 & v3a58674 | !hbusreq4 & v373eaee;
assign v373a66b = hmaster1_p & v3a6f222 | !hmaster1_p & v37265f2;
assign v3a5520d = hlock8_p & v375e21d | !hlock8_p & v3a6f681;
assign v3a714ad = hbusreq4_p & v3726d1f | !hbusreq4_p & v374c8ec;
assign v3a6fdbc = hmaster2_p & v9af7ec | !hmaster2_p & v3763c09;
assign v3723021 = hbusreq5_p & v373aaed | !hbusreq5_p & v3a64089;
assign v3748b15 = hmaster0_p & v37570f8 | !hmaster0_p & v3a5d8bc;
assign v3a57e58 = hmaster2_p & v3809ee4 | !hmaster2_p & v37366d0;
assign v3748e81 = hbusreq3_p & v3a65f0f | !hbusreq3_p & !v8455ab;
assign v23fe285 = hbusreq1_p & v8455e7 | !hbusreq1_p & v3a5e8f6;
assign v3a6f563 = hmaster0_p & v20930c9 | !hmaster0_p & !v937864;
assign v377a477 = hmaster2_p & v3777790 | !hmaster2_p & !v3a71016;
assign v3745b02 = hgrant4_p & v8455ab | !hgrant4_p & v372874c;
assign v376366a = hbusreq8 & v3a6022f | !hbusreq8 & v3771933;
assign v3a6f53a = hmaster2_p & v374355f | !hmaster2_p & v3766b48;
assign v372a48e = hbusreq7_p & v3a6fb8b | !hbusreq7_p & v37741f0;
assign v3757818 = hbusreq0 & v377d2ee | !hbusreq0 & v3777e0e;
assign v3749ff9 = hgrant4_p & v3a702c1 | !hgrant4_p & v3730eae;
assign v374c144 = jx2_p & v377e7f8 | !jx2_p & !v3a5e0c9;
assign v37744f5 = hgrant1_p & v8455ab | !hgrant1_p & v3759c90;
assign v37385e9 = hbusreq7 & v3a6fb4a | !hbusreq7 & v3736ded;
assign v3743e3c = hbusreq7_p & v3a5f5ec | !hbusreq7_p & v375b3b7;
assign v3a710f8 = hlock7 & v3a711cf | !hlock7 & v372f2ff;
assign v3a706af = hbusreq4 & v3a70025 | !hbusreq4 & v3a640a0;
assign v37323a2 = hmaster2_p & v3a709ee | !hmaster2_p & v3a5f6d5;
assign v375e93c = hmaster0_p & v3a619c0 | !hmaster0_p & !v3a703db;
assign v37655c5 = hmaster0_p & v3a705e0 | !hmaster0_p & v3a6fd67;
assign v37426bf = hmaster1_p & v3a6e790 | !hmaster1_p & v3770eeb;
assign v3a585fd = hgrant6_p & v8455ab | !hgrant6_p & !v3a6a3e5;
assign v37365fa = hmaster0_p & v3767f36 | !hmaster0_p & v373a246;
assign v37325eb = hlock5 & v35b7153 | !hlock5 & v3a60f21;
assign v3754940 = hgrant2_p & v8455ab | !hgrant2_p & v3a5affd;
assign v3a6add2 = hbusreq5 & v3a712c0 | !hbusreq5 & v374e78a;
assign v377e8e4 = hmaster2_p & v3a66d94 | !hmaster2_p & v3737e2d;
assign v975066 = hbusreq5 & v3759aca | !hbusreq5 & v3765bf4;
assign v39eb452 = hlock4 & v3733bbe | !hlock4 & v3a6f722;
assign v3a66d0e = hlock4_p & v375bff8 | !hlock4_p & v3760854;
assign v3762cdf = hbusreq7_p & v3a6f031 | !hbusreq7_p & v3a57540;
assign v3745717 = hmaster0_p & v8455ab | !hmaster0_p & v8bc7a8;
assign v374aed5 = hbusreq5 & v3a5d45c | !hbusreq5 & v3a6ffd2;
assign v3766298 = hlock5 & v3a58be6 | !hlock5 & v3734fc3;
assign v3745d3f = hmaster3_p & v376c477 | !hmaster3_p & v8455ab;
assign v3a7152f = hbusreq5 & v376d72e | !hbusreq5 & v3754a74;
assign v28e9804 = hready_p & v94c82c | !hready_p & !v8455d9;
assign v95a0a1 = hmaster2_p & v3a6e5f0 | !hmaster2_p & v3a5690e;
assign v374dd61 = hbusreq2 & v3773c69 | !hbusreq2 & v3a70d64;
assign v3776f5e = hbusreq4_p & v3a71617 | !hbusreq4_p & v3a6157d;
assign v3a71599 = hgrant6_p & v3577306 | !hgrant6_p & ce419c;
assign v376dae8 = jx0_p & v37638f9 | !jx0_p & v372459b;
assign v3a5aefc = hbusreq5 & v373f07d | !hbusreq5 & v3763db6;
assign v3759970 = hlock4_p & v37723a2 | !hlock4_p & v3a602d7;
assign v3a6f586 = hbusreq0_p & v37482f8 | !hbusreq0_p & v8455ab;
assign v37638de = hmaster2_p & v372b1dc | !hmaster2_p & !v3771c59;
assign v3734c59 = hmaster3_p & v3733739 | !hmaster3_p & v374adfa;
assign v3776441 = hbusreq2_p & v3740171 | !hbusreq2_p & v37270d9;
assign v376b5f2 = hgrant7_p & v377b679 | !hgrant7_p & v3737ca0;
assign v3a5a4a0 = hbusreq2 & v3a57d40 | !hbusreq2 & !v8455ab;
assign v37508df = hbusreq8 & v3a7051e | !hbusreq8 & v3756ff6;
assign v3a64ca0 = hbusreq2_p & v374fef7 | !hbusreq2_p & v8455ab;
assign v372e351 = hmaster3_p & v3744f37 | !hmaster3_p & !v376b1ee;
assign v3a70276 = hbusreq5_p & v37361a0 | !hbusreq5_p & v37496de;
assign v37510d9 = hbusreq8_p & v3763c1f | !hbusreq8_p & v3a690a6;
assign v3a704d2 = hgrant5_p & v8455ab | !hgrant5_p & !v3769c4c;
assign v372bad7 = jx0_p & v37235f1 | !jx0_p & v8455ab;
assign v3a6fad5 = hmaster2_p & v37360d1 | !hmaster2_p & v3a6f641;
assign v37246b5 = hbusreq5_p & v3751ebd | !hbusreq5_p & v3776abb;
assign v373d5ab = hmaster2_p & v3a70374 | !hmaster2_p & v3765740;
assign v374bd13 = hbusreq8_p & v3a6fbc2 | !hbusreq8_p & !v8455ab;
assign v3a548b2 = hbusreq3 & v3806db7 | !hbusreq3 & v374f87c;
assign v3737c04 = hmaster0_p & v3744a56 | !hmaster0_p & v3a5bcf5;
assign v3a541f5 = hmaster2_p & v3754450 | !hmaster2_p & v8455ab;
assign v3775e66 = hbusreq0_p & v3a635ea | !hbusreq0_p & v37438c9;
assign v3a680cd = hbusreq8_p & v3a6f1ef | !hbusreq8_p & !v8455ab;
assign v3a6c8c0 = hmaster2_p & v3a713df | !hmaster2_p & v3a5f40e;
assign v3a70ea2 = hlock5_p & v3739531 | !hlock5_p & v37626d8;
assign v3a6c549 = hgrant4_p & v372b77b | !hgrant4_p & v374f126;
assign v3766786 = hbusreq5 & v3a69d8f | !hbusreq5 & v8455ab;
assign v3a70eec = hbusreq3_p & v3a6123a | !hbusreq3_p & v37707eb;
assign v3a70fb7 = hlock5 & v377215c | !hlock5 & v374f7cb;
assign b1f7c8 = hbusreq7_p & v3763a29 | !hbusreq7_p & v3a6f00d;
assign v3a6251b = hbusreq3_p & v376e643 | !hbusreq3_p & v377696a;
assign v374d2e5 = hlock0 & v375200e | !hlock0 & v3a57ac7;
assign v3758c4d = hlock7_p & v375a9d7 | !hlock7_p & !v3a704b8;
assign v3a6f757 = hlock1 & v3a70378 | !hlock1 & v3a70459;
assign v37773d6 = hlock5 & v3a5750b | !hlock5 & v3a6caa7;
assign v376dcdc = hbusreq2_p & v3a70f3e | !hbusreq2_p & v8455b7;
assign v3741b6c = hgrant6_p & v374530a | !hgrant6_p & !v3a6bbeb;
assign v373577f = hgrant6_p & v3a65eba | !hgrant6_p & v373261a;
assign v373c3bd = hmastlock_p & v3a5a496 | !hmastlock_p & v8455ab;
assign v374790d = hbusreq1_p & v377217f | !hbusreq1_p & !v37761e4;
assign v377258d = hmaster1_p & v3738253 | !hmaster1_p & v3a6ad93;
assign v3a6fd1a = hgrant6_p & v8455ab | !hgrant6_p & v3730610;
assign v3a5ac5c = hmaster3_p & v2acb5bc | !hmaster3_p & v372e83a;
assign v3743824 = hbusreq3 & v3379037 | !hbusreq3 & v8455ab;
assign v3a715bb = hbusreq5_p & v3a713e2 | !hbusreq5_p & v373dc11;
assign v3a6caa7 = hmaster0_p & v3741343 | !hmaster0_p & v373d076;
assign v1e3778d = hmaster2_p & v8455ab | !hmaster2_p & !v37277a5;
assign v374723b = hbusreq5 & v3747006 | !hbusreq5 & v8455bf;
assign v377a886 = hlock5_p & v3752845 | !hlock5_p & v8455ab;
assign v3a6fa36 = hgrant2_p & v8455ab | !hgrant2_p & v3a626ea;
assign v3a6146a = hbusreq6 & v3756e01 | !hbusreq6 & v3a7081e;
assign v37747db = hbusreq4_p & v376ea4a | !hbusreq4_p & !v3728e09;
assign v3a71014 = hlock1_p & v8455ab | !hlock1_p & v373fe5e;
assign v3754b35 = hgrant4_p & v377b6ce | !hgrant4_p & v373b600;
assign v37308a8 = hbusreq6 & v3a715d2 | !hbusreq6 & v8455ab;
assign v376c27d = hbusreq5_p & v3732736 | !hbusreq5_p & v3a69ef8;
assign v325b5fd = hlock4_p & v3a687be | !hlock4_p & v373f058;
assign v391331d = hgrant2_p & v8455ab | !hgrant2_p & v3778cdd;
assign v3a68057 = hmaster1_p & v37356f0 | !hmaster1_p & v3a5d417;
assign v380971a = hbusreq2 & v35b7808 | !hbusreq2 & v3a67983;
assign v3760251 = jx0_p & v377609a | !jx0_p & v3a70d72;
assign v3722dcd = hmaster0_p & v3a6fab6 | !hmaster0_p & v390071e;
assign v3758c58 = hmaster2_p & v374a950 | !hmaster2_p & v3a6c97d;
assign v373f172 = hbusreq0 & v3746caf | !hbusreq0 & v3752e13;
assign v3738419 = hgrant2_p & v3750d06 | !hgrant2_p & v374cb90;
assign v374283c = hbusreq2_p & v3741cd7 | !hbusreq2_p & v37731c3;
assign v32562a3 = hbusreq4 & v3a6fc43 | !hbusreq4 & v3a63a66;
assign v375d2ff = hlock8 & v374ebbf | !hlock8 & v3749fc1;
assign v360d036 = hmaster2_p & v3a6b6ef | !hmaster2_p & v3772185;
assign v372bffc = hgrant0_p & v8455ab | !hgrant0_p & v360d016;
assign v3731300 = hbusreq3_p & v8455ab | !hbusreq3_p & v3a6255b;
assign v3741e09 = hmaster1_p & ac043d | !hmaster1_p & v3a65388;
assign v374b51f = hlock5_p & v3a70641 | !hlock5_p & v8455ab;
assign v9375a3 = hlock5 & v3a6fe2d | !hlock5 & v3a6ac20;
assign v3a600f3 = hgrant4_p & v3a6e857 | !hgrant4_p & v376f8bf;
assign v3756813 = hmaster0_p & v3a5e696 | !hmaster0_p & v37607af;
assign v374dba6 = hbusreq7 & v3730a90 | !hbusreq7 & v3729370;
assign v3a64a5d = hbusreq8 & v3a6a52c | !hbusreq8 & v3723025;
assign v37482c7 = hmaster2_p & v376a6f1 | !hmaster2_p & v375248f;
assign v3a6c355 = hbusreq3 & v3765e46 | !hbusreq3 & v8455ab;
assign v3747b30 = hmaster1_p & v375a268 | !hmaster1_p & v376a85d;
assign v3767690 = hlock6_p & v3724a4b | !hlock6_p & v3730ffe;
assign v376f468 = jx1_p & v3723447 | !jx1_p & v3739983;
assign v3a6fedb = hbusreq3_p & v3745f4a | !hbusreq3_p & v3754e7b;
assign v3a707b5 = hbusreq4_p & v3a60787 | !hbusreq4_p & v3733d6e;
assign v3a69e18 = hlock0_p & v372fba5 | !hlock0_p & v8455b0;
assign v3a6f5df = hbusreq1 & v376111d | !hbusreq1 & v8455ab;
assign v373f23c = hgrant3_p & v38070c1 | !hgrant3_p & v3a5eac0;
assign v373bc28 = hmaster2_p & v3a70ee7 | !hmaster2_p & v372493b;
assign v377d58d = hbusreq0 & v3a7068a | !hbusreq0 & v3a6002a;
assign v374fa4c = hbusreq6_p & v3a64252 | !hbusreq6_p & v374f8b1;
assign v3a684ee = hmaster1_p & v3a5b23c | !hmaster1_p & !v376ad8c;
assign v375c0cb = hbusreq3 & v37366d0 | !hbusreq3 & v8455ab;
assign v372bb5d = hbusreq7_p & v372b009 | !hbusreq7_p & d62ab4;
assign v3737d48 = hgrant2_p & v8455ba | !hgrant2_p & v377fa89;
assign v372a352 = hbusreq8 & v3a6eeb9 | !hbusreq8 & !v8455ab;
assign v3734625 = stateA1_p & v8455ab | !stateA1_p & !v3a293c5;
assign v372c706 = hgrant6_p & v377f09a | !hgrant6_p & v360d080;
assign v375e167 = hbusreq5 & v3a705b2 | !hbusreq5 & v372b798;
assign v377c9cc = hlock0 & v3a635ea | !hlock0 & v3775e78;
assign v3756109 = hmaster2_p & v372673d | !hmaster2_p & v3a6f442;
assign v3728045 = hmaster2_p & v3a5af94 | !hmaster2_p & !v3a5bf04;
assign v3a70a6e = hmaster2_p & v3a635ea | !hmaster2_p & v3749437;
assign v3747bea = hgrant6_p & v3a68f98 | !hgrant6_p & v3a7103d;
assign v37266c2 = hlock4 & v377dd65 | !hlock4 & v375f302;
assign v373d506 = hgrant3_p & v3a712f0 | !hgrant3_p & v373c6a2;
assign v3777670 = hmaster1_p & v3a6ff69 | !hmaster1_p & c4699e;
assign v375b6d4 = hbusreq5 & v3750fc9 | !hbusreq5 & v3a5fc34;
assign v3758fc4 = hmaster1_p & v3a6a758 | !hmaster1_p & v3a5ceaf;
assign v3757ebc = hmaster1_p & v3726240 | !hmaster1_p & v374e21e;
assign v3a708cd = hgrant7_p & v2093005 | !hgrant7_p & v3740bba;
assign v372f434 = hbusreq7_p & v3a6f5b8 | !hbusreq7_p & !v3a6fd5d;
assign v3751359 = hbusreq0 & v3a2abd2 | !hbusreq0 & v8455ab;
assign v3a6ad46 = hbusreq5_p & v373e474 | !hbusreq5_p & v375607f;
assign v3740de5 = hlock0 & v3778f6c | !hlock0 & v374cd7e;
assign v373c79c = hgrant0_p & v375dab1 | !hgrant0_p & v3770993;
assign v3808e88 = hmaster1_p & v3a635ea | !hmaster1_p & v3a5f6da;
assign v3a70db1 = hmaster0_p & v3766307 | !hmaster0_p & v372c14d;
assign v3a6f8cf = hbusreq7_p & v3763c1f | !hbusreq7_p & v375610e;
assign v89c52e = hbusreq6 & v3a56518 | !hbusreq6 & v372d48d;
assign v3a5e7fe = hlock2_p & v3765e46 | !hlock2_p & !v8455ab;
assign v373a228 = hmaster1_p & v372834d | !hmaster1_p & v3a5d644;
assign v1e37bde = hbusreq5_p & v3a6f7d0 | !hbusreq5_p & v3a68399;
assign v373da11 = jx2_p & v375b031 | !jx2_p & v3a6f3d7;
assign v360d099 = hbusreq8_p & v3a70962 | !hbusreq8_p & v8455ab;
assign v37548a5 = hbusreq5 & v37318e3 | !hbusreq5 & v377e018;
assign v3755b94 = hgrant6_p & v8455ca | !hgrant6_p & v3a65dc4;
assign v372c483 = hmaster0_p & v3730e7d | !hmaster0_p & v3a5c7a3;
assign v3732da2 = hbusreq7_p & v3a70655 | !hbusreq7_p & v3a7013d;
assign v3745484 = hgrant3_p & v375d288 | !hgrant3_p & v373b17c;
assign v37447b9 = hmaster0_p & v3725b69 | !hmaster0_p & v3a6e8d9;
assign v372cb99 = hbusreq0 & v3a704de | !hbusreq0 & v375b3be;
assign v3a70d6d = hbusreq8 & v3779f68 | !hbusreq8 & v3740a94;
assign v861ce0 = hmaster1_p & v8455ab | !hmaster1_p & !v3750519;
assign v377f6a5 = hbusreq7_p & v3727823 | !hbusreq7_p & v37669d0;
assign v3772edc = hbusreq4 & v372a94e | !hbusreq4 & v373484e;
assign v374752b = hmaster1_p & v3739eed | !hmaster1_p & v3a6fd9b;
assign v3a586f1 = hbusreq6 & v3743da3 | !hbusreq6 & v8455ab;
assign v3765474 = hbusreq6_p & v376fe96 | !hbusreq6_p & v3a55d7c;
assign v37386da = hbusreq0 & v375df77 | !hbusreq0 & v8455ab;
assign v3777186 = hbusreq7_p & v376c08d | !hbusreq7_p & v3a6e675;
assign v375e961 = hbusreq8 & v373d97a | !hbusreq8 & v3a5bb57;
assign v3753b80 = hmaster2_p & v3a6d569 | !hmaster2_p & v376954d;
assign v3a70326 = hbusreq2_p & v376ef42 | !hbusreq2_p & v3733e9e;
assign v3741e82 = hbusreq0_p & v3a5ae6d | !hbusreq0_p & v373e8b5;
assign v3a6a093 = hmaster1_p & v3a60974 | !hmaster1_p & v3a70f68;
assign v372b91e = hmaster0_p & v3a5408e | !hmaster0_p & !v373a246;
assign v374f3e3 = hgrant6_p & v3a6f402 | !hgrant6_p & v3a62041;
assign v3a710d3 = hbusreq8 & v3a71610 | !hbusreq8 & v86d727;
assign v37317c0 = hgrant2_p & v3a5c0de | !hgrant2_p & !v3a6f0e3;
assign v375cc17 = hmaster2_p & v376bd43 | !hmaster2_p & v8455ab;
assign v3a60a40 = hbusreq6_p & v3a62041 | !hbusreq6_p & v3759623;
assign v3724345 = hmaster1_p & v3731ca8 | !hmaster1_p & v3a6fab4;
assign v37458dc = hbusreq2 & v373e521 | !hbusreq2 & v37496fa;
assign v23fda78 = hbusreq5_p & v3769023 | !hbusreq5_p & v3a7107f;
assign v3754d88 = hmaster2_p & v3a70364 | !hmaster2_p & v380777f;
assign v3747f5d = hgrant2_p & v3a5f50e | !hgrant2_p & v376e238;
assign v3a7157c = hgrant5_p & v3728876 | !hgrant5_p & v3755423;
assign v374ca88 = hbusreq6_p & v3a70326 | !hbusreq6_p & v3766bc8;
assign v3738c2e = hmaster2_p & v3773262 | !hmaster2_p & v377472b;
assign v3742ec4 = hgrant6_p & v376305b | !hgrant6_p & v3a6fe94;
assign v3a715a4 = hmaster1_p & v3738726 | !hmaster1_p & v8455e7;
assign v374d94e = hmaster0_p & v3751253 | !hmaster0_p & v375355a;
assign v374d480 = hbusreq2 & v3751dc9 | !hbusreq2 & v3a635ea;
assign v3740348 = hbusreq4 & v37386f5 | !hbusreq4 & !v8455b9;
assign v374ec35 = hmaster0_p & v3728d9c | !hmaster0_p & v377ae32;
assign v3a6f645 = hmaster1_p & v3a60bee | !hmaster1_p & v8455ab;
assign v3a5e881 = hbusreq2_p & v884deb | !hbusreq2_p & v373b288;
assign v3a68915 = hbusreq5 & v373a263 | !hbusreq5 & v37694a0;
assign v3776039 = hmaster0_p & v3a635ea | !hmaster0_p & v3725c41;
assign v3764983 = hmaster1_p & v37752be | !hmaster1_p & v3a60b37;
assign v37331a2 = hmaster0_p & v3a62e91 | !hmaster0_p & v3758fa8;
assign v3a5f2c0 = hbusreq5_p & v3a70cb2 | !hbusreq5_p & v372fecd;
assign v375b99c = hmaster1_p & v37403cc | !hmaster1_p & !v3a70f1e;
assign v372f7c6 = hbusreq3_p & v3a6f2dd | !hbusreq3_p & v37455ec;
assign v37343d1 = hgrant5_p & v37308fc | !hgrant5_p & v3a7015e;
assign v375e52f = hmaster2_p & v8455ab | !hmaster2_p & !v3a70385;
assign v3740825 = hlock5_p & v374e745 | !hlock5_p & !v8455ab;
assign v3729308 = hmaster0_p & v377d1dc | !hmaster0_p & v372fa3a;
assign v3a5bd69 = hmaster2_p & v3753f62 | !hmaster2_p & v373f172;
assign v37480c6 = hbusreq5 & v37625a0 | !hbusreq5 & v8455ab;
assign v372b72d = hmaster0_p & v3777ad7 | !hmaster0_p & v8455ab;
assign v3a6f907 = hgrant4_p & v8455ab | !hgrant4_p & v3a5524c;
assign v37665e1 = hmaster2_p & v374ad81 | !hmaster2_p & v3a6eaf4;
assign v3728d9c = hgrant4_p & v8455ab | !hgrant4_p & !v3a6ebf9;
assign v3778765 = hgrant0_p & v8455ab | !hgrant0_p & v372b351;
assign v3746e8b = hmaster2_p & v374b5a8 | !hmaster2_p & v3a621cb;
assign v37393ad = hmaster2_p & v8455ab | !hmaster2_p & v3a6f9ae;
assign v3a612df = hgrant5_p & v3774fee | !hgrant5_p & v3733ee4;
assign v3a60443 = hbusreq7 & v377b8f9 | !hbusreq7 & v374a4cc;
assign dafc4e = hmaster2_p & v3736ee0 | !hmaster2_p & v3a6fd5a;
assign v3746e54 = hmaster3_p & v3378b65 | !hmaster3_p & v2ff8e61;
assign v3a705c0 = hmaster3_p & v3752ed7 | !hmaster3_p & v3a5cf84;
assign v3a70bf7 = hbusreq0 & v3a5f0cf | !hbusreq0 & v3a57f42;
assign v3756b8a = hbusreq0 & v375d445 | !hbusreq0 & v39eb709;
assign v374355d = hbusreq2 & v372d078 | !hbusreq2 & v376e90a;
assign v38097ca = hlock6 & v372eeee | !hlock6 & v37638ee;
assign v372a0e6 = hgrant8_p & v3a66039 | !hgrant8_p & v37788d7;
assign v3a714e8 = hgrant2_p & v8455ab | !hgrant2_p & v3767fa5;
assign v37741bc = hbusreq3 & v376ed91 | !hbusreq3 & v3776fe2;
assign v375a64f = hmaster0_p & v3763b6c | !hmaster0_p & v8455ab;
assign v3772214 = hgrant5_p & v3a5caf4 | !hgrant5_p & !v3807386;
assign v372a80a = hmaster0_p & v3775aa7 | !hmaster0_p & v3809d9e;
assign v3771882 = hmaster0_p & v3a5e747 | !hmaster0_p & v3a66615;
assign v372af6d = jx1_p & v3a6f523 | !jx1_p & v8727d2;
assign v3a61c5e = hgrant8_p & v3a55ec8 | !hgrant8_p & v3765293;
assign v37285eb = hgrant6_p & v8455ab | !hgrant6_p & v3a7011e;
assign v3a5cd72 = hgrant6_p & v3a654c1 | !hgrant6_p & v3a706ed;
assign v37704dc = hbusreq0 & v3a66f0d | !hbusreq0 & v8455ab;
assign v3767797 = hmaster0_p & v376639f | !hmaster0_p & v3735f79;
assign v37615d8 = hgrant6_p & v377cb2b | !hgrant6_p & v374f78c;
assign v376c2e2 = hgrant0_p & v3a70e93 | !hgrant0_p & !v373e5ad;
assign v377e904 = hgrant4_p & v8455ab | !hgrant4_p & v3725d7b;
assign v3763474 = hbusreq7_p & v377ccbf | !hbusreq7_p & v372ee18;
assign v373efdf = hbusreq7 & v374457b | !hbusreq7 & v376ae9f;
assign v3776e2b = hmaster2_p & v3a5e24e | !hmaster2_p & !v3a6d684;
assign v37643e6 = hmaster2_p & v375e53a | !hmaster2_p & v37554b1;
assign v375199a = hbusreq5 & v3a701ec | !hbusreq5 & v3a70cf4;
assign v3a702d3 = hbusreq4_p & v376df24 | !hbusreq4_p & v33782e5;
assign v3a6bc78 = hbusreq1_p & v375ac98 | !hbusreq1_p & v8455b0;
assign v3a70283 = hbusreq6_p & v37456a9 | !hbusreq6_p & v373c728;
assign v377291b = hmaster2_p & v376498f | !hmaster2_p & v3a65d01;
assign v3766a69 = hbusreq8_p & v38079c2 | !hbusreq8_p & v373a41e;
assign v37419d7 = hmaster3_p & v3778a4f | !hmaster3_p & v3768c19;
assign v377a6f2 = hgrant2_p & v3a6fbe2 | !hgrant2_p & v3747dfc;
assign v376ae7f = hlock5 & v3a6a4b9 | !hlock5 & v3a69539;
assign v3a6cfc5 = hmaster2_p & v3a5c945 | !hmaster2_p & !v3735e39;
assign v3778565 = start_p & v8455ab | !start_p & v3a6ff57;
assign v3758b45 = hbusreq5 & v3a7165a | !hbusreq5 & v377edd6;
assign v3724936 = hmaster1_p & v37763b2 | !hmaster1_p & v373a693;
assign v3a6fa99 = hlock7 & v3734279 | !hlock7 & v3808e3a;
assign v3a70291 = jx2_p & v373de47 | !jx2_p & v377e962;
assign v375564e = hbusreq6_p & v8455ab | !hbusreq6_p & v375975b;
assign v3a646f5 = hbusreq2_p & v3a5795e | !hbusreq2_p & v3a6f147;
assign v374bf07 = hmaster2_p & v3723430 | !hmaster2_p & v3a696ed;
assign v23fd98d = hburst1 & v3a6ffa9 | !hburst1 & v3a5a220;
assign v372e711 = hbusreq4_p & v3a635ea | !hbusreq4_p & v373b288;
assign v373f5b1 = hbusreq7_p & v3a7018d | !hbusreq7_p & v3a71030;
assign v373ac71 = hmaster2_p & v3753c2a | !hmaster2_p & v377fc1f;
assign v377d354 = hbusreq4_p & v377eaf2 | !hbusreq4_p & v292555a;
assign v3734256 = hgrant0_p & v3a64c10 | !hgrant0_p & !v3773a9d;
assign v3768f0c = hbusreq4_p & v3747a97 | !hbusreq4_p & v3736f61;
assign v373ddfc = hmaster1_p & v3a6fdd1 | !hmaster1_p & v3a707f3;
assign v3a7012b = hmaster2_p & v3a61a7f | !hmaster2_p & v3a6fdef;
assign v3a6f3bb = hgrant6_p & v8455ab | !hgrant6_p & v373fbca;
assign v37403ef = hmaster2_p & v374314f | !hmaster2_p & b66167;
assign v23fde98 = hgrant2_p & a54211 | !hgrant2_p & v37562f2;
assign v37444c9 = hmaster0_p & v377795a | !hmaster0_p & !v3a706e3;
assign v3a70410 = hbusreq0 & v376a272 | !hbusreq0 & v3a6f9ac;
assign v3a6009a = hmaster1_p & v3a66d94 | !hmaster1_p & v37676c3;
assign v372a20f = hbusreq6_p & v3a6f8f9 | !hbusreq6_p & v3a5c779;
assign v377405e = hmaster0_p & v375b7b0 | !hmaster0_p & v3740d4a;
assign v376eeac = hgrant3_p & v8455ab | !hgrant3_p & v3a5d7bf;
assign v3728e91 = hmaster1_p & v3a635ea | !hmaster1_p & v37c36bf;
assign v3a713b0 = hmaster1_p & v3761d2f | !hmaster1_p & v3761bac;
assign v374fe2d = hlock8_p & v3a58307 | !hlock8_p & v3a7064e;
assign v3a5ef5c = hbusreq1_p & v377a275 | !hbusreq1_p & !v8455ab;
assign v3768985 = hbusreq6 & v3760740 | !hbusreq6 & v8455ab;
assign v3765298 = hbusreq8_p & v372a95a | !hbusreq8_p & !v374ff02;
assign v3a70f8b = hmaster0_p & v377094d | !hmaster0_p & v3726991;
assign v3809d87 = hgrant6_p & v3a653e4 | !hgrant6_p & !v3a6ef50;
assign v376dc16 = hgrant6_p & v8455ab | !hgrant6_p & v3a6ebf8;
assign v38070c1 = hbusreq3_p & v3a59b5c | !hbusreq3_p & !v8455ab;
assign v3769023 = hmaster0_p & v3a6eb72 | !hmaster0_p & v373026e;
assign v377814d = jx1_p & v39eb1dc | !jx1_p & v3764fd5;
assign v3730cde = hmaster2_p & v3760513 | !hmaster2_p & v3a2a13a;
assign v3a571b6 = hlock6 & v377f611 | !hlock6 & v374fa0d;
assign v3760bf8 = hbusreq3_p & v1e379fe | !hbusreq3_p & v374d85e;
assign v37390ec = hbusreq7_p & v3775806 | !hbusreq7_p & v373287a;
assign v372dd98 = hmaster0_p & v3a65b87 | !hmaster0_p & v3757ffa;
assign v3a7129f = hbusreq0 & v377a50f | !hbusreq0 & v372b1e3;
assign v3a714e1 = hlock4 & v3770fbc | !hlock4 & v3a703bb;
assign v37683bf = hmaster1_p & v37570eb | !hmaster1_p & v3a6e844;
assign v3753f62 = hbusreq0 & v3738855 | !hbusreq0 & v375e1a1;
assign v373f7ff = hbusreq4 & v3a5abf4 | !hbusreq4 & !v372fbeb;
assign v3734f7b = hbusreq4_p & v3763d52 | !hbusreq4_p & v3a5f26f;
assign v3a59ffa = hbusreq3_p & v373cdb7 | !hbusreq3_p & v3a61c5a;
assign v3a6f094 = hmaster2_p & v8455b0 | !hmaster2_p & v375ac23;
assign v3774841 = hmaster0_p & v3730e7d | !hmaster0_p & v3a6f15c;
assign v3722dfb = hmaster2_p & v37356f0 | !hmaster2_p & adf78a;
assign v37643ee = start_p & v3a59da9 | !start_p & v3733a6c;
assign v3a70d5f = hmaster0_p & v372b840 | !hmaster0_p & !v8455e7;
assign v3a6f55c = hbusreq8 & v3a5a3d0 | !hbusreq8 & v372d811;
assign v3a702a5 = hbusreq0_p & v375863a | !hbusreq0_p & v373e67e;
assign v373b209 = hbusreq6_p & v3806f68 | !hbusreq6_p & v8455b0;
assign v372e479 = hmaster1_p & v373373d | !hmaster1_p & v37266df;
assign v373af15 = hmaster1_p & v376fa43 | !hmaster1_p & v375d78f;
assign d5bac5 = hmaster2_p & v3a6fa7a | !hmaster2_p & v372b6bc;
assign v3a6ae68 = hbusreq2_p & v3a5a510 | !hbusreq2_p & !v1e382e7;
assign v3a6d71b = hgrant4_p & v3a71128 | !hgrant4_p & v3a6da6b;
assign v37531af = hgrant2_p & v8455ab | !hgrant2_p & v3a6fcd4;
assign v3a6af71 = hlock4_p & v375913f | !hlock4_p & v374b0bc;
assign v3771e6f = hmaster2_p & v8455ab | !hmaster2_p & v3a6fcb0;
assign v374829e = hgrant6_p & v375cfa5 | !hgrant6_p & v3a70f8d;
assign v3a5b660 = hbusreq7_p & v3771cac | !hbusreq7_p & v8455b7;
assign v3a6f7eb = jx0_p & v3737438 | !jx0_p & v376b71f;
assign v372731e = hbusreq2_p & v37765e1 | !hbusreq2_p & v3a6edb9;
assign v3a6581d = hmaster0_p & v3a6ead8 | !hmaster0_p & !v2925cbb;
assign v3a5f292 = hbusreq2 & v374c718 | !hbusreq2 & v8455ab;
assign v374093f = hmaster2_p & v37496fa | !hmaster2_p & v375da10;
assign v3728c5b = hmaster2_p & v3a70893 | !hmaster2_p & v8455ab;
assign v3760fab = hgrant6_p & v3734cb7 | !hgrant6_p & v3a6ccd6;
assign v373fdf0 = hmaster1_p & v3a6ffd3 | !hmaster1_p & v3a6a1d1;
assign v375d0ed = hbusreq6_p & v374cab9 | !hbusreq6_p & v37484df;
assign v3762c26 = hgrant2_p & v374068b | !hgrant2_p & v3725649;
assign v373e98b = hgrant3_p & v8455ab | !hgrant3_p & v3773837;
assign v3a6efe8 = hbusreq3_p & v373afb4 | !hbusreq3_p & v8455ab;
assign v3725872 = hgrant7_p & v8455c1 | !hgrant7_p & v3730712;
assign v3766803 = hmaster0_p & v3807f45 | !hmaster0_p & v3a6a536;
assign v3736a23 = hgrant6_p & v376495e | !hgrant6_p & v3a7008c;
assign v3739a3b = hbusreq4 & v377cdf0 | !hbusreq4 & v3a5f9e6;
assign v374fd12 = hmaster1_p & v3a6fc99 | !hmaster1_p & v3a66c84;
assign v373ee51 = hbusreq4 & v37739f4 | !hbusreq4 & v3734ec1;
assign v3732eaa = hbusreq7 & v374039d | !hbusreq7 & v373e0b1;
assign v3751210 = hmaster1_p & v376832f | !hmaster1_p & v37229e6;
assign v8a94c2 = hmaster2_p & v3a637dd | !hmaster2_p & !v3a6b873;
assign v3727a16 = hbusreq5 & v3a711c6 | !hbusreq5 & v3733d4f;
assign v373f028 = hgrant2_p & v3a6b129 | !hgrant2_p & v3a6f8bb;
assign v3a706a1 = hmaster2_p & v376d268 | !hmaster2_p & v92e6f3;
assign v3a6dfc9 = hlock6 & v3a6b393 | !hlock6 & v3a65827;
assign a33229 = hmaster0_p & v3a71381 | !hmaster0_p & v377f34a;
assign v3a68482 = hmaster2_p & v37386c6 | !hmaster2_p & v3a70374;
assign v37721e3 = hgrant6_p & v8455c9 | !hgrant6_p & v3a7127e;
assign v3761bd1 = hmaster0_p & v3a60395 | !hmaster0_p & v3758d6c;
assign v3a6c0ab = hmaster2_p & v8455bd | !hmaster2_p & !v8455ab;
assign v3a5ddc1 = hgrant4_p & v8455c2 | !hgrant4_p & v3a623ca;
assign v3745b66 = hbusreq5 & v376967e | !hbusreq5 & v3729ee6;
assign v3a5cc17 = hbusreq6_p & v3a5e95a | !hbusreq6_p & v376f48d;
assign v3779075 = hmaster1_p & v372455c | !hmaster1_p & v3724f1d;
assign v377d1cd = hbusreq4 & v3a6fd2d | !hbusreq4 & v39ea0c5;
assign c827f4 = hlock6_p & v8455ab | !hlock6_p & v8455e7;
assign v376460f = hgrant4_p & v3a5bffe | !hgrant4_p & !v3a70731;
assign v3761efb = hgrant3_p & v8455ab | !hgrant3_p & !v3724d93;
assign v3742649 = hmaster0_p & c10173 | !hmaster0_p & v8455ab;
assign v3a70f0d = hmaster0_p & v3a635ea | !hmaster0_p & v374797c;
assign v3a68c1c = hgrant2_p & v3779e45 | !hgrant2_p & v373f5d3;
assign v3752eda = hbusreq6_p & v3a56e7a | !hbusreq6_p & v8455b3;
assign v3762b52 = hlock5_p & v3760681 | !hlock5_p & v8455ab;
assign v375a0ec = hgrant6_p & v3730926 | !hgrant6_p & a6859a;
assign v37690bf = hmaster2_p & v8455ab | !hmaster2_p & v3736806;
assign v3a57444 = hlock5_p & v8455ab | !hlock5_p & v376142a;
assign v3775cb7 = hmaster2_p & v3a70d99 | !hmaster2_p & v3a705c5;
assign v3a62819 = hmaster0_p & v3a635ea | !hmaster0_p & v39e9c98;
assign v3a5ebde = hlock3_p & v3a637dd | !hlock3_p & !v8455ab;
assign v3a6c15c = hmaster1_p & v3a6ffbc | !hmaster1_p & v3759b46;
assign v3a6fda7 = hbusreq2_p & v3a6efce | !hbusreq2_p & !v8455ab;
assign v23fd83f = hbusreq0 & v3a70c7a | !hbusreq0 & v372e863;
assign v3a6f0ca = hmaster1_p & v3748ff3 | !hmaster1_p & v35b77ab;
assign v374f8a5 = hbusreq7 & v372c5a0 | !hbusreq7 & v374837b;
assign v3779283 = hbusreq4 & v375b40c | !hbusreq4 & v8455ab;
assign v3a6d81e = hmaster2_p & v8455ab | !hmaster2_p & v374a877;
assign v37419b2 = hmaster0_p & v375921f | !hmaster0_p & !v3732c95;
assign v376999e = hbusreq6 & v39a5293 | !hbusreq6 & v3377b1b;
assign v374f8f6 = hbusreq5 & v3a65e9d | !hbusreq5 & v3a5fc34;
assign v372bb4b = jx1_p & v37461d8 | !jx1_p & v3a7046a;
assign v3732f8d = hgrant4_p & v37785b8 | !hgrant4_p & v3a671de;
assign v2acae99 = hmaster0_p & v3a6cd8b | !hmaster0_p & v3762ffa;
assign v373b10f = hgrant2_p & v8455ab | !hgrant2_p & v3724a1c;
assign v3a6f4f7 = hbusreq7 & v376e66e | !hbusreq7 & v376e9ed;
assign v376e8e3 = hmaster1_p & v375ba6d | !hmaster1_p & v3739d2a;
assign v3746da7 = hbusreq5_p & v3a5e618 | !hbusreq5_p & v3a5e030;
assign v374e52d = hmaster2_p & v3774bad | !hmaster2_p & v374d54c;
assign v3739ba9 = hbusreq4 & v3750dd3 | !hbusreq4 & v8455bb;
assign v3806ef3 = hbusreq4_p & v23fd8cb | !hbusreq4_p & v3a69946;
assign v3761ac7 = hbusreq6_p & v373ce84 | !hbusreq6_p & v3a7011e;
assign v374bc63 = hbusreq5_p & v373f996 | !hbusreq5_p & v8455ab;
assign v3a6f1fb = hbusreq4_p & v3725799 | !hbusreq4_p & v372a116;
assign v372e305 = hbusreq3 & v3a6d4c2 | !hbusreq3 & v3379037;
assign v372c35a = hlock6_p & v3a7116b | !hlock6_p & !v8455ab;
assign v3741249 = hmaster2_p & v3a67a6f | !hmaster2_p & v37358ab;
assign v374cacb = hmaster0_p & v373b0e7 | !hmaster0_p & v373e15b;
assign v3768dbc = hbusreq5_p & v3807754 | !hbusreq5_p & v3758f02;
assign v3a29520 = hmaster0_p & v3764f60 | !hmaster0_p & v372d42d;
assign v3a66c94 = hmaster1_p & v3742f76 | !hmaster1_p & !v374b0a3;
assign v991591 = hbusreq8 & v3757ab6 | !hbusreq8 & v372e02d;
assign v377ea20 = hgrant4_p & v8455ab | !hgrant4_p & v376513c;
assign v377451f = hlock5 & v3a6d64e | !hlock5 & v3776039;
assign v37612c1 = hmaster0_p & v3a5fabd | !hmaster0_p & v3763b94;
assign v373e782 = hlock2_p & v37625a8 | !hlock2_p & v3a5ace5;
assign v3a70edc = hbusreq1 & v37665bf | !hbusreq1 & v8455ab;
assign v3735bbb = hmaster0_p & v3731724 | !hmaster0_p & v375dfcf;
assign v3757858 = hbusreq8 & v374e05d | !hbusreq8 & !v8455ab;
assign v3744b55 = hbusreq0 & v3a661fe | !hbusreq0 & v3a700b2;
assign v3767258 = hgrant6_p & v3a69146 | !hgrant6_p & v3a63690;
assign v37696fe = hgrant4_p & v1e37996 | !hgrant4_p & v3725bfb;
assign v375d46e = hmaster1_p & v3a6f92f | !hmaster1_p & v3779883;
assign v3a6f79b = hgrant6_p & v8455ab | !hgrant6_p & v3a6abdc;
assign v3a6f600 = hlock7 & v37243ac | !hlock7 & v374be73;
assign v3a555d1 = hbusreq6_p & v373bfea | !hbusreq6_p & v3a629a6;
assign v373ec29 = hbusreq7 & v373dc53 | !hbusreq7 & v3a6fb20;
assign v374f318 = hgrant0_p & v8455ab | !hgrant0_p & !v3776a6e;
assign v372d727 = hgrant4_p & v3a53eeb | !hgrant4_p & v377c34f;
assign v3a6773a = hbusreq3_p & v373997b | !hbusreq3_p & v37738fc;
assign v37697ba = hlock6 & v917087 | !hlock6 & v3a5a7fd;
assign v3756aaa = hmaster2_p & v3a71678 | !hmaster2_p & v37674f6;
assign v3a70fa6 = hgrant4_p & v8455ab | !hgrant4_p & v37558e4;
assign v37bfd3a = hgrant5_p & v375f83b | !hgrant5_p & v373ae02;
assign v3a70052 = hbusreq5_p & v375ebc3 | !hbusreq5_p & v3a6f48e;
assign v3a5dafb = hmaster0_p & v3a6a8ee | !hmaster0_p & v3a70369;
assign v3737c88 = hmaster1_p & v37731ce | !hmaster1_p & v1e374d4;
assign v3729f13 = hmaster1_p & v377accc | !hmaster1_p & v372e2cd;
assign v3725688 = hmaster1_p & v3a57f59 | !hmaster1_p & v3a70dd8;
assign v3762dcf = hmaster2_p & v3778bde | !hmaster2_p & v375352f;
assign v373923a = hlock8_p & v3a70472 | !hlock8_p & v3755d23;
assign v3768995 = hbusreq5_p & v377766c | !hbusreq5_p & v3731857;
assign v3a6123e = hbusreq1_p & v375a842 | !hbusreq1_p & v3732b98;
assign v373c263 = hgrant5_p & v3a67af1 | !hgrant5_p & v374a058;
assign v375fac2 = hmaster1_p & v3729972 | !hmaster1_p & v3a71656;
assign v3a5ca22 = hbusreq8 & v3a6a9d3 | !hbusreq8 & v37776c8;
assign v373499c = hmaster0_p & v377eea3 | !hmaster0_p & v3774a95;
assign v376a149 = hbusreq4 & v375b18e | !hbusreq4 & v373031f;
assign v3756da3 = jx0_p & v3774d9c | !jx0_p & v375e510;
assign v3760a0b = hmaster0_p & v2acafac | !hmaster0_p & v3a6f3cd;
assign v3a6f9a0 = hgrant0_p & v8455ab | !hgrant0_p & v3722be8;
assign v372f694 = stateA1_p & v3a5ff81 | !stateA1_p & v37464c8;
assign v3a6f3cf = hbusreq0_p & v3a6fe6a | !hbusreq0_p & !v8455ab;
assign v3a68d26 = jx1_p & v3734965 | !jx1_p & v3730b5a;
assign v1e37cf9 = hmaster2_p & v3a714fd | !hmaster2_p & v374ab4f;
assign v1e37af3 = hmaster2_p & v3a715c1 | !hmaster2_p & v375a397;
assign v3a6ffc6 = hbusreq4 & v3a7151d | !hbusreq4 & !v8455ab;
assign v3a70c9a = hbusreq4_p & v3739bcd | !hbusreq4_p & v3a70822;
assign v37577b6 = hbusreq4 & v3a654c1 | !hbusreq4 & v375da10;
assign v376cedc = hbusreq4 & v372eaaf | !hbusreq4 & v377395f;
assign v373553c = hbusreq8_p & v3a5bc0a | !hbusreq8_p & v3a6a918;
assign v3a62009 = hbusreq8 & v3a70bc0 | !hbusreq8 & v8455ab;
assign v3a56002 = hmaster2_p & v377f584 | !hmaster2_p & !v8455ab;
assign v3a5ec50 = hbusreq5 & v3749540 | !hbusreq5 & v37363ae;
assign v3760a2c = hbusreq4 & v373a291 | !hbusreq4 & v8455ab;
assign v372545e = hmaster0_p & v3742cd4 | !hmaster0_p & v377f13c;
assign v373dac4 = hmaster0_p & v3a5d548 | !hmaster0_p & v3a59bbd;
assign v3747666 = hmaster2_p & v37422b5 | !hmaster2_p & v3a6f520;
assign v96dd76 = hgrant4_p & v8455c1 | !hgrant4_p & v374586a;
assign v3a70c39 = hlock4_p & v8455b0 | !hlock4_p & !v8455ab;
assign v3a6e699 = hgrant2_p & v3a62826 | !hgrant2_p & v3a5eeb4;
assign v3a6f1d8 = hmaster1_p & v3a635ea | !hmaster1_p & v37710a4;
assign v3a65af6 = hbusreq8_p & v3a578ef | !hbusreq8_p & v37378d4;
assign v373af55 = hmaster2_p & v3a6ffd3 | !hmaster2_p & v3a6fa93;
assign v3a6ff3c = hlock3 & v377cc23 | !hlock3 & v3732715;
assign v3a707ab = hbusreq5_p & v376539b | !hbusreq5_p & !v3a6eb54;
assign v3a711be = hbusreq8 & v3a6f6f2 | !hbusreq8 & a80fe2;
assign v3a5ce2f = hgrant1_p & v8455b6 | !hgrant1_p & !v8455ab;
assign v37351f6 = hmaster1_p & v8455ab | !hmaster1_p & v377c500;
assign v3775da7 = hburst0 & v3757c6f | !hburst0 & v375f479;
assign v37799a0 = hmaster1_p & v3806fc0 | !hmaster1_p & v3768ae9;
assign v375b9c1 = hlock0_p & v3a635ea | !hlock0_p & !v3a5b451;
assign v37690e7 = hmaster1_p & v3a5cdef | !hmaster1_p & v3757a04;
assign v372cd3f = hbusreq6 & v3774b56 | !hbusreq6 & v8455ab;
assign v37298be = hbusreq5_p & v3a638aa | !hbusreq5_p & v3a68525;
assign v372bcd0 = hmaster2_p & v37406d2 | !hmaster2_p & v37796c6;
assign d3b3b2 = hlock0_p & v3a635ea | !hlock0_p & v3779264;
assign v3a706c3 = hbusreq8 & v3755f23 | !hbusreq8 & v372863f;
assign v37609e7 = hbusreq2_p & v3748797 | !hbusreq2_p & v372e30d;
assign v37631a9 = hmaster0_p & v3756f77 | !hmaster0_p & v3a6fec4;
assign b15d44 = jx2_p & v3a6c022 | !jx2_p & v374a526;
assign c8ab71 = hbusreq4_p & v377e934 | !hbusreq4_p & !v3a6830a;
assign v3742582 = hmaster2_p & v3a5c85c | !hmaster2_p & v3a600f3;
assign v3770071 = hmaster0_p & v8455b5 | !hmaster0_p & !v35b774b;
assign v37493c7 = hmaster2_p & v8455ab | !hmaster2_p & !v3a703fc;
assign v373ccde = hbusreq0 & v3a70a18 | !hbusreq0 & v3a6603d;
assign v3756506 = hbusreq0 & v374b3cf | !hbusreq0 & v373e814;
assign v375c76b = hmaster2_p & v37747c0 | !hmaster2_p & v3746e85;
assign v3a61c1f = hmaster2_p & v3747302 | !hmaster2_p & v374d0e3;
assign v3726c20 = hgrant4_p & v3a5a0d2 | !hgrant4_p & v3768af7;
assign v3a5b181 = hbusreq5 & v377b6de | !hbusreq5 & v3760a0b;
assign v377edd6 = hmaster0_p & v3a700e2 | !hmaster0_p & v375ea85;
assign v376049c = hgrant0_p & v3733e9e | !hgrant0_p & v376b3b0;
assign v37744e0 = hmaster2_p & v3725bdc | !hmaster2_p & !v8455ab;
assign v373fdfb = hmaster2_p & v3743bbe | !hmaster2_p & v3779e1b;
assign v3746976 = hbusreq7_p & v375ea88 | !hbusreq7_p & v3a54e0c;
assign v3a6f4d2 = hbusreq2 & v3809b31 | !hbusreq2 & v37450b8;
assign v3a70423 = hlock5 & v3761dda | !hlock5 & v3778857;
assign v3a702fd = jx0_p & v3731a2e | !jx0_p & v377047f;
assign v3a6f656 = hbusreq1_p & v3a690ff | !hbusreq1_p & !v377a018;
assign v3743b62 = hmaster1_p & v8455c2 | !hmaster1_p & v37675f1;
assign v3a70681 = hmaster3_p & v373436a | !hmaster3_p & v3a5cff1;
assign v3750adf = hbusreq0 & v3749008 | !hbusreq0 & v3764c9c;
assign v3774d6e = hbusreq5 & v3770ad8 | !hbusreq5 & v3a635ea;
assign v37472b6 = hgrant7_p & v3a707ff | !hgrant7_p & v3a6ff06;
assign v3728399 = hbusreq0 & v3726905 | !hbusreq0 & !v8455ab;
assign v37684b7 = hmaster0_p & v3770621 | !hmaster0_p & v3756820;
assign v3738a50 = hmaster2_p & v8455e7 | !hmaster2_p & !v8455ab;
assign v374743a = jx2_p & v87f2ea | !jx2_p & v3a59656;
assign v3a6ffbd = hlock0 & v3a6c5ee | !hlock0 & v3a6e50e;
assign v3a60cdb = hbusreq4 & v3a70b1e | !hbusreq4 & !v8455ca;
assign v3a595ba = hlock6 & v373bf4f | !hlock6 & v373f1ac;
assign v3738b0b = hmaster2_p & v9bf1d8 | !hmaster2_p & v377e19d;
assign v376f2c8 = hlock5 & v3a6c64d | !hlock5 & v3809968;
assign v3723698 = hbusreq8 & v3740c94 | !hbusreq8 & v372b61a;
assign v3738adf = hbusreq4_p & v376d41b | !hbusreq4_p & v3757a57;
assign v3a6dac0 = hlock8 & v376fbce | !hlock8 & v3763046;
assign v3807670 = hmaster2_p & v3a6a546 | !hmaster2_p & v3a6f907;
assign v3a57e27 = hlock5_p & v372df76 | !hlock5_p & !v8455ab;
assign v3762815 = hlock1_p & b56d1b | !hlock1_p & v8455b0;
assign v3a6fc3b = hmaster2_p & v3777cfc | !hmaster2_p & v372d2dc;
assign v3a5d405 = hbusreq5 & v377653f | !hbusreq5 & v37383da;
assign v3731499 = hmaster1_p & v376bd43 | !hmaster1_p & v3739e36;
assign v3748caf = hbusreq4_p & b1ca9b | !hbusreq4_p & v377957e;
assign v3808870 = hgrant2_p & v37443ab | !hgrant2_p & v8455ab;
assign v3752f8e = hmaster1_p & v3771076 | !hmaster1_p & v3a58306;
assign v3a5ab9d = hbusreq2 & v3a54c77 | !hbusreq2 & v8455ab;
assign v3741fee = hbusreq8 & v372a6de | !hbusreq8 & v3a647ce;
assign v3a5711b = hmaster2_p & v39a4dbb | !hmaster2_p & !v3a5fdd3;
assign v373d452 = stateA1_p & v39a5381 | !stateA1_p & v8455ab;
assign v373bf1d = hmaster2_p & v377bdc3 | !hmaster2_p & !v372c571;
assign v3a680b9 = hbusreq2_p & v3a5795e | !hbusreq2_p & v3755e35;
assign v3a6c38a = hbusreq5_p & v3755883 | !hbusreq5_p & v377d545;
assign v3a6fbac = hmaster0_p & v3a29d87 | !hmaster0_p & !v3a5ef76;
assign v3a61cb5 = hmaster2_p & v3a6fa7a | !hmaster2_p & v374d8ac;
assign v377b7e0 = hmaster1_p & v3748ac8 | !hmaster1_p & v3729949;
assign v373c2e1 = hmaster1_p & v3a5a01b | !hmaster1_p & v3733e4f;
assign v3a6b5bc = hgrant6_p & v37414b0 | !hgrant6_p & v3a58a8e;
assign v3742034 = hbusreq1 & v374ccb7 | !hbusreq1 & v8455ab;
assign v23fe353 = hbusreq5 & v3a714cd | !hbusreq5 & !v8455ab;
assign v37593a4 = hmaster0_p & v3a6ff15 | !hmaster0_p & v372d42d;
assign v3a71530 = hlock5_p & v35b774b | !hlock5_p & !v3770071;
assign v376b018 = hbusreq2 & v376e316 | !hbusreq2 & v37366b5;
assign v3a6f9f8 = hbusreq3_p & v375082a | !hbusreq3_p & v8455b0;
assign v3760091 = hmaster0_p & v374efb9 | !hmaster0_p & v3a655e9;
assign v372bef4 = hmaster1_p & v373e376 | !hmaster1_p & v3a64e01;
assign v3a6f8d0 = hbusreq0 & v3a5784f | !hbusreq0 & v3775636;
assign v3a61094 = hmaster0_p & v377b429 | !hmaster0_p & v37540d9;
assign v3759a34 = hbusreq4_p & v37450a5 | !hbusreq4_p & !v35772a6;
assign v3740b58 = hbusreq7_p & v376c08d | !hbusreq7_p & v8455cb;
assign v374a891 = hgrant0_p & v3a655c2 | !hgrant0_p & v3a6b2ef;
assign v374aacc = hmaster2_p & v3a635ea | !hmaster2_p & v3760881;
assign v374df88 = hbusreq8 & v3a63fbc | !hbusreq8 & v8455ab;
assign v3776b93 = hbusreq5 & v37350a4 | !hbusreq5 & v38076cf;
assign v3a583dc = hgrant3_p & v373cdbf | !hgrant3_p & v3a6665c;
assign v3a70ff5 = hbusreq4_p & v373f2e2 | !hbusreq4_p & v8455ab;
assign v376c592 = hmaster1_p & v374502e | !hmaster1_p & v3a5bb49;
assign v3741869 = hbusreq5_p & v376e72d | !hbusreq5_p & v360d136;
assign v3a6898d = hbusreq4_p & v3a635ea | !hbusreq4_p & v3769302;
assign v3771e69 = hmaster0_p & v3a71180 | !hmaster0_p & v1e37cc1;
assign v37661b2 = hlock4_p & v372b24d | !hlock4_p & v3a70131;
assign v37784b3 = hbusreq5 & v377b26a | !hbusreq5 & v3a68787;
assign v373759d = hmaster0_p & v8455e7 | !hmaster0_p & v3726d94;
assign v37420de = hbusreq5_p & v373f022 | !hbusreq5_p & v3739a23;
assign v3767183 = hmaster3_p & v3744deb | !hmaster3_p & v3a70424;
assign v372787e = hbusreq5 & v372f235 | !hbusreq5 & v3764dac;
assign v3733557 = hmaster0_p & v8455ab | !hmaster0_p & v3a712d0;
assign v3753921 = hmaster0_p & v3a706a8 | !hmaster0_p & v3777e7d;
assign v3a539af = hlock0 & v3a64af7 | !hlock0 & v3738c75;
assign v3a70a70 = hbusreq0 & v380988c | !hbusreq0 & v3776faf;
assign v374a157 = hmaster0_p & v3a635ea | !hmaster0_p & v3a6f959;
assign v37407cb = hmaster2_p & v374502e | !hmaster2_p & v3a6f018;
assign v376ea50 = hmaster1_p & v375db64 | !hmaster1_p & v3a611cf;
assign v3a7077a = hmaster0_p & v3735907 | !hmaster0_p & v3a6fcab;
assign v20d166d = hmastlock_p & v3760a9d | !hmastlock_p & v8455ab;
assign v3748c3f = hgrant5_p & v373ad69 | !hgrant5_p & v3a6fd77;
assign v3756f21 = jx1_p & v373faf3 | !jx1_p & v372ecad;
assign v3a6fa7a = hbusreq4_p & v3777197 | !hbusreq4_p & v8455ab;
assign v376aa6d = hbusreq3_p & a11f42 | !hbusreq3_p & v8455ab;
assign v3a6be15 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3745de0;
assign v3a7108f = hbusreq0 & v375af36 | !hbusreq0 & v3730a2f;
assign v3729808 = hmaster1_p & v37241db | !hmaster1_p & v374db0f;
assign v37738ae = hmaster0_p & v3a5c473 | !hmaster0_p & v3729004;
assign v3752a7a = hgrant4_p & v3a7133d | !hgrant4_p & v3a70948;
assign v3a689eb = hgrant3_p & v3a55d41 | !hgrant3_p & v376fe30;
assign v3a6b58f = hbusreq7 & v3729d06 | !hbusreq7 & v1e37943;
assign v376fe96 = hbusreq6 & v3a6fbd9 | !hbusreq6 & v3738114;
assign v3a6fab8 = hmaster2_p & v3a6fa4c | !hmaster2_p & v37320ff;
assign v376c12e = hgrant3_p & v3a6d70a | !hgrant3_p & v8455ab;
assign v372f12d = hgrant6_p & v375c7b9 | !hgrant6_p & v3760c90;
assign hgrant6 = !v37bfff7;
assign v374ea29 = hmaster2_p & v3a64349 | !hmaster2_p & !v3a63a7a;
assign v9ccd8a = hbusreq2_p & v3729b37 | !hbusreq2_p & v37764ee;
assign v375a613 = hgrant0_p & v373bd24 | !hgrant0_p & v3a5ae2f;
assign v3a6eb8b = hgrant2_p & v8455ab | !hgrant2_p & v372514f;
assign v3748da1 = hlock7_p & v3761da5 | !hlock7_p & v3761916;
assign v3778a2f = hbusreq5_p & v3774937 | !hbusreq5_p & v3a62cb7;
assign v3751a33 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a63e9e;
assign v3a5762d = hmaster0_p & v374b03c | !hmaster0_p & v372f1d4;
assign v3754176 = hlock0 & v3a641d5 | !hlock0 & v3a68954;
assign v3a6e884 = hmaster1_p & v3757966 | !hmaster1_p & v373198c;
assign v374067c = hbusreq5 & v3a6fd24 | !hbusreq5 & v8455ab;
assign v3a70d4e = hlock7_p & v3768636 | !hlock7_p & v3a5f47b;
assign v3a6ebff = hgrant1_p & v37732c0 | !hgrant1_p & v3809adf;
assign v3a5fd34 = hbusreq2_p & v8455ab | !hbusreq2_p & v376c235;
assign v375ed6f = hbusreq4_p & v3a65da7 | !hbusreq4_p & v377e1f6;
assign v3a6bcf9 = hbusreq4_p & v380956d | !hbusreq4_p & v3759eb6;
assign v377af10 = hbusreq4 & v3a67691 | !hbusreq4 & v3a5e2e1;
assign v377961f = hbusreq3_p & v3a70edb | !hbusreq3_p & v8455ab;
assign v3a6fe3e = hgrant2_p & v3a7156d | !hgrant2_p & v3a6ff3f;
assign v3737b19 = hmaster1_p & v3772f0f | !hmaster1_p & v3a70e99;
assign v1e3737f = hbusreq7_p & v372f03c | !hbusreq7_p & v3a6667c;
assign v37325c5 = hlock5 & v3a5414c | !hlock5 & v3a6fda1;
assign v376d9aa = hlock6 & v3a6f659 | !hlock6 & v884deb;
assign v3a5d63f = hbusreq4 & v374eb89 | !hbusreq4 & v8455ab;
assign v3777226 = hmaster2_p & v8455e7 | !hmaster2_p & v3a7156d;
assign v3a68d2e = hbusreq1_p & v3a635ea | !hbusreq1_p & !v37533b4;
assign v3749a4c = hbusreq5 & v3a70ea1 | !hbusreq5 & v3745458;
assign v3773016 = hgrant1_p & v37467f3 | !hgrant1_p & v377989c;
assign v3a6f571 = hgrant6_p & v3764486 | !hgrant6_p & v8ad83a;
assign v377a89f = hgrant5_p & v3a67acf | !hgrant5_p & v37399f7;
assign v373695f = hbusreq5_p & v3a566eb | !hbusreq5_p & v372647d;
assign v3a6f1f8 = hbusreq0_p & v35772a5 | !hbusreq0_p & !v3770af1;
assign v3734918 = hbusreq6 & v3a6f7bf | !hbusreq6 & v8455e7;
assign v375c366 = hmaster2_p & v37386c6 | !hmaster2_p & v3a70f53;
assign v377b429 = hbusreq4_p & v374e51a | !hbusreq4_p & v375af98;
assign v3a702bd = hmaster2_p & v3a61a7f | !hmaster2_p & v3a6ff99;
assign v3807003 = hbusreq6_p & v3a5fdd3 | !hbusreq6_p & !v3a627cc;
assign v3744bfc = hbusreq6_p & v3a700cd | !hbusreq6_p & !v8455ab;
assign v375798a = hgrant6_p & v8455ab | !hgrant6_p & v3806e35;
assign v3723ac5 = hbusreq1_p & v375d80d | !hbusreq1_p & !v8455ab;
assign v375cd50 = hmaster0_p & v3a5d259 | !hmaster0_p & v372700a;
assign v3752b4b = hgrant3_p & v8455ab | !hgrant3_p & v3a605e8;
assign v3a5ed98 = hbusreq7 & v3a6f4b9 | !hbusreq7 & v377386a;
assign v3729bc6 = hmaster2_p & v3a6162f | !hmaster2_p & v3a71526;
assign v375a4d0 = hmaster0_p & v3770b26 | !hmaster0_p & v377bfc7;
assign v375f8f2 = hmaster0_p & v373a756 | !hmaster0_p & v372f1d4;
assign v3a70e10 = hlock2 & v29256ae | !hlock2 & v3762cc4;
assign v3758bbd = hbusreq4_p & v38072fd | !hbusreq4_p & v3739078;
assign v374089e = hgrant1_p & v3756bc9 | !hgrant1_p & v3a70c07;
assign v376df02 = hbusreq2_p & v377f83c | !hbusreq2_p & v3748d67;
assign v3744ad5 = hbusreq8_p & v3a6fe0c | !hbusreq8_p & v3a71305;
assign v3a6a6c6 = hmaster0_p & v8455b5 | !hmaster0_p & v3a6f5a5;
assign v3725098 = hmaster2_p & v1e38275 | !hmaster2_p & v3a59e87;
assign v3a56d86 = hlock4 & v372f83b | !hlock4 & v3a5dd17;
assign v376bea3 = hlock6 & db903b | !hlock6 & v3a5ef89;
assign v375b265 = hbusreq1 & v35b9d52 | !hbusreq1 & !v8455ab;
assign v3a58c15 = hmaster0_p & v375f2f3 | !hmaster0_p & d26e1e;
assign v3a6f4ec = hgrant6_p & v3a6f18f | !hgrant6_p & v3741401;
assign v3748c75 = hmaster1_p & v37341fd | !hmaster1_p & v3a70c8f;
assign v375c65f = hbusreq5_p & v372a24d | !hbusreq5_p & v375fb9d;
assign v374a454 = hmaster0_p & v3a6bf04 | !hmaster0_p & v3761719;
assign v3726139 = hbusreq1_p & v8455ab | !hbusreq1_p & v374fb58;
assign v376f92c = hlock8_p & v3a7113f | !hlock8_p & v3a6242b;
assign v3a712e4 = hmaster0_p & v3a6f094 | !hmaster0_p & v372f9cf;
assign v3743b9e = locked_p & v8455ab | !locked_p & v3a63621;
assign v3754543 = hgrant2_p & v3a62524 | !hgrant2_p & v3777749;
assign v377d769 = hmaster2_p & v8455e7 | !hmaster2_p & v8455ab;
assign v375a2a3 = hmaster0_p & v8455ab | !hmaster0_p & v3a55f0d;
assign v3726505 = hlock4 & v3750d46 | !hlock4 & v3a539bb;
assign v3745d21 = hlock3_p & v2925c67 | !hlock3_p & v23fdbca;
assign v376f80c = hmaster2_p & v3807f45 | !hmaster2_p & v3a62a6d;
assign v3751261 = hbusreq5 & v3764910 | !hbusreq5 & v3a6d0af;
assign v3a70bc7 = hbusreq2 & adf78a | !hbusreq2 & v8455ab;
assign v375825a = hgrant0_p & v3735f56 | !hgrant0_p & v3a670a1;
assign v3732034 = hbusreq3 & v8455ab | !hbusreq3 & v95d97e;
assign v377ac4c = hgrant6_p & v377f09a | !hgrant6_p & !v3a7062c;
assign v3762223 = hgrant2_p & v3751d98 | !hgrant2_p & v3a57484;
assign v375a03b = hmaster2_p & v8455ab | !hmaster2_p & v3761031;
assign v3750371 = stateA1_p & v3a6efc9 | !stateA1_p & v2acb5a2;
assign v377c4d7 = hbusreq7 & v3749165 | !hbusreq7 & v373c263;
assign v372c84a = hgrant6_p & v8455ab | !hgrant6_p & !v3a635c3;
assign v3a6ac66 = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3a6eba3;
assign v3a6bddd = hlock1 & v3a6891e | !hlock1 & v3a581bd;
assign v375f53a = hbusreq6_p & d78807 | !hbusreq6_p & v373cde8;
assign v3772443 = hbusreq2 & v3a7119e | !hbusreq2 & v8455ab;
assign v373f622 = hgrant3_p & v8455ab | !hgrant3_p & v373d5d6;
assign v3724976 = hmaster3_p & v3a5fd2f | !hmaster3_p & v3a6312c;
assign v372d60f = hbusreq4 & v374cab9 | !hbusreq4 & v37674c1;
assign v376f505 = hbusreq6_p & v377e2f7 | !hbusreq6_p & v3769cd6;
assign v375e574 = hmaster2_p & v3a54c77 | !hmaster2_p & v35772c9;
assign v374749d = hmaster2_p & v377db14 | !hmaster2_p & v3a641d5;
assign v3a6a635 = jx0_p & v375f60e | !jx0_p & v377af48;
assign v374307e = jx0_p & v3255a0f | !jx0_p & v3a5f717;
assign v372e6a1 = hbusreq6_p & v3a6a261 | !hbusreq6_p & v3776751;
assign v3737416 = hgrant2_p & v3a70403 | !hgrant2_p & v3a63b90;
assign v377afaa = hgrant5_p & v376a454 | !hgrant5_p & v3a712a7;
assign v377c9a1 = hmaster2_p & v3a6f9d7 | !hmaster2_p & v8455ab;
assign v3776395 = hlock7 & v3a6ffe9 | !hlock7 & v3730b1c;
assign v375b05e = hbusreq4_p & v3a6f9d1 | !hbusreq4_p & v8455ab;
assign v3748792 = hbusreq2_p & v376d658 | !hbusreq2_p & v375ab6d;
assign v3a71326 = hmaster0_p & v3730789 | !hmaster0_p & v3a6fbd1;
assign v3738f8a = hbusreq7 & v376b28c | !hbusreq7 & v8455ab;
assign v3723134 = hbusreq5_p & v3a5dbd7 | !hbusreq5_p & !v8455ab;
assign v3a6f59e = hmaster0_p & v3a62846 | !hmaster0_p & v3a6e872;
assign v376b57e = hbusreq6_p & v373a2f2 | !hbusreq6_p & v3737534;
assign v3762969 = hmaster0_p & v3725198 | !hmaster0_p & v3808f73;
assign v373cf66 = hbusreq5_p & v3808994 | !hbusreq5_p & v377a60f;
assign v3a715d7 = hmaster0_p & v8455ab | !hmaster0_p & v3a61be2;
assign v3a70b71 = hmaster2_p & v8455b0 | !hmaster2_p & v3a5f40e;
assign v3a6f73c = hbusreq5 & v3a6b462 | !hbusreq5 & v8455ab;
assign v377f401 = hbusreq0 & v3a6f52c | !hbusreq0 & v373185f;
assign v374bdac = hbusreq7 & v3727a6d | !hbusreq7 & v3a6f6e0;
assign v3a658ad = hgrant3_p & v3761b90 | !hgrant3_p & !v8455ab;
assign v375df8e = hmaster2_p & v377c6ce | !hmaster2_p & v3a710c8;
assign v3a7038e = hbusreq6 & v35772a2 | !hbusreq6 & v8455ab;
assign v377f190 = hlock0_p & v3a5ae6d | !hlock0_p & v3741e82;
assign v37711cc = hbusreq6_p & v37776b6 | !hbusreq6_p & v3773fd1;
assign v3a660f2 = hbusreq1_p & v3a70641 | !hbusreq1_p & v3733383;
assign v3769ee7 = hmaster1_p & v37739ed | !hmaster1_p & !v8455ab;
assign v375f67d = hmaster0_p & v380974c | !hmaster0_p & v373908c;
assign v377ecac = hmaster2_p & v372e27b | !hmaster2_p & v8455b3;
assign v375af58 = hbusreq0 & v377e864 | !hbusreq0 & v8455ab;
assign v3773b4b = hbusreq7 & v3a6eb9d | !hbusreq7 & v37761d1;
assign v3a6eb67 = hlock5 & v3774ab8 | !hlock5 & v3a5e4e5;
assign v3a7107e = hmaster0_p & v377b058 | !hmaster0_p & v3769923;
assign v3731172 = hbusreq6 & v374df14 | !hbusreq6 & v3a6da8a;
assign v3a705cb = hmaster0_p & v3a637dc | !hmaster0_p & v3759dfb;
assign v3a6241d = hbusreq3 & v376111d | !hbusreq3 & v8455ab;
assign v3a58287 = hmaster2_p & v375463e | !hmaster2_p & v3739b4c;
assign v373e062 = hmaster1_p & v8455ab | !hmaster1_p & v3771440;
assign v373650c = hbusreq2_p & v372904d | !hbusreq2_p & v3378fb8;
assign v375554d = hbusreq7 & v3577487 | !hbusreq7 & v376382f;
assign v3a690ff = hgrant1_p & v374fb58 | !hgrant1_p & !v3a637dd;
assign v375238e = hbusreq5 & v374f307 | !hbusreq5 & v8455b0;
assign v3769ec3 = hbusreq5_p & v37335ff | !hbusreq5_p & v3756f8c;
assign v3a6b896 = hgrant5_p & v3748eff | !hgrant5_p & v373a228;
assign v3a61323 = hmaster0_p & c86567 | !hmaster0_p & v3769820;
assign v3a70fe9 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3765e79;
assign v3a68793 = hgrant4_p & v3734b97 | !hgrant4_p & v3a70c3a;
assign v3a70d09 = hbusreq5 & v8455ab | !hbusreq5 & !v374066d;
assign v3764f01 = hmaster3_p & v3a5cca9 | !hmaster3_p & v377b017;
assign v3737f89 = hlock3 & v3722f58 | !hlock3 & v37566f4;
assign v373755a = hlock5_p & v8455e7 | !hlock5_p & !v375534d;
assign v3a6b89e = hbusreq6_p & v3761224 | !hbusreq6_p & v3a6557d;
assign v377bb86 = hbusreq3 & v374ea45 | !hbusreq3 & v8455ab;
assign v3a63994 = decide_p & v376233b | !decide_p & v373139d;
assign v375f3ac = hlock5 & v35b77ae | !hlock5 & v374544c;
assign v3745f76 = busreq_p & v3809adf | !busreq_p & !v3748422;
assign v3751c8c = hbusreq4 & v380a0c2 | !hbusreq4 & v37255d9;
assign v374f12d = hbusreq3_p & v3745d21 | !hbusreq3_p & v8455ab;
assign v3764628 = hmaster0_p & v3751c73 | !hmaster0_p & v3761719;
assign v3a71283 = hgrant6_p & v375b01a | !hgrant6_p & v3728a12;
assign v3a5ff7c = hmaster1_p & v3a64eba | !hmaster1_p & v3a6f78f;
assign v373df89 = hbusreq4_p & v3a60a23 | !hbusreq4_p & v374c58c;
assign v37710a4 = hbusreq5_p & v3a6eaf8 | !hbusreq5_p & v3a5f4c6;
assign v37551e3 = hbusreq2 & v372f76a | !hbusreq2 & v374f35a;
assign v372625f = hgrant4_p & v8455e7 | !hgrant4_p & !v3755ad5;
assign v375766c = hbusreq5_p & v360d10b | !hbusreq5_p & !v8455ab;
assign v37272a8 = hbusreq2_p & v3779227 | !hbusreq2_p & v3a6fdf7;
assign v3a6377a = hmaster1_p & v3737415 | !hmaster1_p & v3755ffc;
assign v372fddd = hgrant8_p & v3a6f409 | !hgrant8_p & v376b706;
assign v376d795 = hmaster1_p & v3739d2c | !hmaster1_p & v374e7fa;
assign v3a67ffe = hbusreq6_p & v375b68b | !hbusreq6_p & v375b943;
assign v3a59e74 = hgrant6_p & v377f09a | !hgrant6_p & !v3732939;
assign v375eb79 = hbusreq5_p & v37653ef | !hbusreq5_p & !v3a6491d;
assign v377c5c2 = hbusreq2 & v3a70118 | !hbusreq2 & !v8455bd;
assign v375301b = hlock6_p & v3a6ff5c | !hlock6_p & v3a6dfc6;
assign v377564e = hbusreq4 & c2c2bc | !hbusreq4 & v373eaee;
assign v375a1ab = hgrant4_p & v3732b35 | !hgrant4_p & v3731f7a;
assign v374f89b = hbusreq0 & v3a5f154 | !hbusreq0 & v3a6b18c;
assign v38074c0 = jx0_p & v373e365 | !jx0_p & v3747d0a;
assign v3a658cf = hmaster2_p & v3a53a94 | !hmaster2_p & v3a70272;
assign v3775c0a = hgrant3_p & v8455ab | !hgrant3_p & v3766572;
assign v376d06c = hbusreq8_p & v3779cb5 | !hbusreq8_p & v372c834;
assign v37516ba = hmaster2_p & v377d27a | !hmaster2_p & v8455ab;
assign v37626d8 = hmaster0_p & v3a7114c | !hmaster0_p & v373ad3f;
assign v3a5bd76 = hmaster2_p & v8455b0 | !hmaster2_p & v376ddc6;
assign v3746fcb = hbusreq5_p & v3a6f61a | !hbusreq5_p & !v8455ab;
assign v37494ee = hbusreq2 & v373fe5e | !hbusreq2 & v3a7136f;
assign v9ed0ba = hlock5_p & v3a6602e | !hlock5_p & v372995e;
assign v3757dea = hgrant5_p & v3737f5a | !hgrant5_p & v3a297f5;
assign v37fca9f = hgrant8_p & v8455d2 | !hgrant8_p & a04f67;
assign v3806def = hmaster0_p & v377a366 | !hmaster0_p & v8455ab;
assign v3a6f56c = hbusreq0 & v3a58a1b | !hbusreq0 & v37362b5;
assign v3a5891c = locked_p & v8455ab | !locked_p & !v3809adf;
assign v3750625 = hbusreq4 & v3a70468 | !hbusreq4 & v37686c2;
assign v3a5b875 = hbusreq5 & v376a6f1 | !hbusreq5 & !v3a7127c;
assign v3761433 = hbusreq4_p & v3773fbb | !hbusreq4_p & v375c608;
assign v372562a = hbusreq8 & v3a6b336 | !hbusreq8 & v376ef20;
assign v3a700ea = hmaster0_p & v3a6c4e4 | !hmaster0_p & v375eb29;
assign v37590f4 = hmaster2_p & v3747358 | !hmaster2_p & !v373c111;
assign v3756fba = hgrant3_p & v3757264 | !hgrant3_p & v3a7037c;
assign v3755420 = hgrant6_p & v8455ab | !hgrant6_p & v3a71558;
assign v8455f7 = hgrant7_p & v8455ab | !hgrant7_p & !v8455ab;
assign v3753aa5 = hgrant5_p & v8455ab | !hgrant5_p & !v3a5b070;
assign a61746 = hgrant5_p & v8455c6 | !hgrant5_p & v37587a4;
assign v3a5ed86 = hmaster0_p & v3a635ea | !hmaster0_p & v3745bdc;
assign v3a62b8d = hbusreq6_p & v3a70297 | !hbusreq6_p & v3a708a2;
assign v3a7029f = hbusreq0 & v37574d3 | !hbusreq0 & v372d967;
assign v3768c78 = hbusreq4_p & v3733d6e | !hbusreq4_p & v372ee7e;
assign v375e9a9 = hlock5 & v37602e0 | !hlock5 & v377f26e;
assign v3a5c65d = hgrant5_p & v3a60a56 | !hgrant5_p & v3a601cd;
assign v376b88d = hbusreq2_p & v3a71344 | !hbusreq2_p & v8455ab;
assign v3a6f5a6 = hmaster2_p & v3a5a510 | !hmaster2_p & v3a6d684;
assign v8455ff = stateG2_p & v8455ab | !stateG2_p & !v8455ab;
assign v3a70d86 = hbusreq6 & v372e03f | !hbusreq6 & v8455ab;
assign v3807b40 = hbusreq1_p & v372692d | !hbusreq1_p & v3a70c66;
assign v3a703f1 = hgrant3_p & v3745236 | !hgrant3_p & v3a70d22;
assign v3a6fb62 = hbusreq3 & v375969d | !hbusreq3 & v3a708c2;
assign v3739ac1 = hbusreq6_p & v3a64969 | !hbusreq6_p & v8455b3;
assign v377876f = hbusreq0 & v3733d45 | !hbusreq0 & v3a56372;
assign v377005e = hgrant3_p & v8455e7 | !hgrant3_p & !v3733d5a;
assign v35ba2da = hbusreq4_p & v3768e0c | !hbusreq4_p & v8455ab;
assign v3a60fd6 = hlock6 & v374d3b8 | !hlock6 & v3a709d0;
assign v373c126 = hbusreq8 & v37597fa | !hbusreq8 & v3a6f068;
assign v375f4e8 = hlock6 & v3a6670c | !hlock6 & v3733334;
assign v3a6ad59 = hgrant3_p & v8455ab | !hgrant3_p & v3a5f7f3;
assign v3763299 = hgrant2_p & v37648af | !hgrant2_p & !v37292f4;
assign v374e99f = hmaster0_p & v3730d18 | !hmaster0_p & v3a70666;
assign v1e3825d = hbusreq3_p & v3740ee1 | !hbusreq3_p & v3a66ff2;
assign v3a6db95 = hlock5_p & v3a56ebd | !hlock5_p & v8455ab;
assign v373a6d9 = hmaster0_p & v3a61f4c | !hmaster0_p & v374aa46;
assign v373b012 = hbusreq6_p & v375f326 | !hbusreq6_p & v3a6fe8e;
assign v37480b7 = hbusreq4_p & v375121b | !hbusreq4_p & v8455ab;
assign v372b7e6 = hbusreq8 & v373055b | !hbusreq8 & v3732c96;
assign v3a6f336 = hmaster0_p & v376d9ad | !hmaster0_p & v376a7ac;
assign v37786c6 = hmaster1_p & v3752428 | !hmaster1_p & v3a6fa0a;
assign v372e863 = hlock0 & v3a57959 | !hlock0 & v3a70c7a;
assign v3737c6c = hgrant2_p & v3a54108 | !hgrant2_p & v375e7d6;
assign v3a70434 = hlock7 & v3770f56 | !hlock7 & v3734cce;
assign v37435a0 = hbusreq2_p & v377eaf2 | !hbusreq2_p & v3735512;
assign v3a700d7 = hbusreq5 & v3758561 | !hbusreq5 & v376784b;
assign v3a65c31 = hmaster0_p & v377e089 | !hmaster0_p & v372bd5f;
assign v373bc8f = hmaster1_p & v3730d16 | !hmaster1_p & !v37615d0;
assign v374efb9 = hmaster2_p & v3a655e9 | !hmaster2_p & v3769740;
assign v3a6ec10 = hbusreq8_p & v3a6e7a4 | !hbusreq8_p & v37449d1;
assign v3762bbe = stateG10_1_p & v3a70c07 | !stateG10_1_p & v37603f4;
assign v3a5db7d = hbusreq7 & v3777989 | !hbusreq7 & v3a701bf;
assign v3a5f308 = stateA1_p & v3762fc4 | !stateA1_p & v3807071;
assign v3a5b3e6 = hbusreq5 & v377f298 | !hbusreq5 & v8455ab;
assign v3a5c998 = hmaster0_p & v37686c7 | !hmaster0_p & !v37411c6;
assign v3764ced = hlock0 & v3752cf6 | !hlock0 & v3a70f18;
assign v3a6f7db = jx0_p & v3751440 | !jx0_p & v374a25d;
assign v376d41b = hbusreq0 & a708cc | !hbusreq0 & v377e24d;
assign v3a6b97b = hlock0_p & v3a6f32f | !hlock0_p & v3a70a6d;
assign v374ddef = hmaster1_p & v3724394 | !hmaster1_p & c45930;
assign v372700b = hmaster1_p & v375f159 | !hmaster1_p & v37402ee;
assign v3a5a307 = hmaster1_p & v3757966 | !hmaster1_p & v374b4ef;
assign v37788d6 = hbusreq8 & v3a64f1f | !hbusreq8 & v3a674c4;
assign v374bcac = hbusreq6_p & v373ff4a | !hbusreq6_p & v2092f59;
assign v3752e65 = hbusreq3_p & v374af0d | !hbusreq3_p & v8455ab;
assign v3775557 = hbusreq0_p & v35772c9 | !hbusreq0_p & v8455ab;
assign v3a6fd2a = hbusreq0_p & v35772a5 | !hbusreq0_p & !v376d327;
assign v3777787 = hbusreq1_p & v3a6fc6c | !hbusreq1_p & v3731dc6;
assign v3a5c46a = hgrant5_p & v376ba63 | !hgrant5_p & !v8455ab;
assign v376a847 = hmaster1_p & v374a454 | !hmaster1_p & v3729516;
assign v3a6eb2b = hgrant2_p & v376e1ed | !hgrant2_p & v3730122;
assign v3a6eee3 = hbusreq7_p & v3a57fa1 | !hbusreq7_p & v3740451;
assign v37c02a9 = hbusreq0 & v3775d59 | !hbusreq0 & v8455ab;
assign v3a58e79 = hgrant5_p & v3a714b0 | !hgrant5_p & !v8455ab;
assign v3a6ef50 = hbusreq6_p & v8455ab | !hbusreq6_p & !v3a637dd;
assign v373fe8f = hgrant5_p & v372fef2 | !hgrant5_p & v3769980;
assign v3a6f3c4 = hbusreq4 & v3742ec4 | !hbusreq4 & v380719b;
assign v2889703 = hbusreq2 & v3774c4d | !hbusreq2 & v3a641d5;
assign v3a6f85a = hmaster2_p & v3a6b2c9 | !hmaster2_p & v372e4cf;
assign v372373f = hbusreq1 & v3763175 | !hbusreq1 & v8455ab;
assign v3a7074e = hmaster2_p & v3768a9c | !hmaster2_p & v3a5bb64;
assign v37693a9 = hgrant3_p & v8455ab | !hgrant3_p & v374ac72;
assign v3a6de5e = hgrant7_p & v3737c21 | !hgrant7_p & v372fe43;
assign v377613b = hmaster2_p & v3734967 | !hmaster2_p & !v37625a8;
assign v3731866 = hmaster0_p & v3779060 | !hmaster0_p & v3736d5e;
assign v3749503 = hmaster1_p & v3a61a7f | !hmaster1_p & v360bc74;
assign v3a7002c = hgrant4_p & v3a6ffb6 | !hgrant4_p & v3755928;
assign v3a6f87f = hgrant2_p & v374b72f | !hgrant2_p & !v8455ab;
assign v3a6f047 = hbusreq5 & v3a6f3ef | !hbusreq5 & !v37730ec;
assign v373a4ea = hmaster2_p & v377d1a3 | !hmaster2_p & !v3752fbc;
assign v3a5ee99 = hgrant0_p & v8455ab | !hgrant0_p & v39a4dd4;
assign v373ee66 = hmaster1_p & v3a5f97f | !hmaster1_p & !v3a5cf3c;
assign v3a5378e = hlock4 & v98381a | !hlock4 & v3755a70;
assign v374bfa2 = hbusreq5_p & v39eb4e4 | !hbusreq5_p & v374d9fe;
assign v377e469 = hbusreq6_p & v376ea4a | !hbusreq6_p & !v3728e09;
assign v3a5ead4 = hbusreq5_p & a747d7 | !hbusreq5_p & v37bfc35;
assign v375d00a = hbusreq4 & v376e7e8 | !hbusreq4 & v8455ab;
assign v3739c81 = hgrant6_p & v8455ca | !hgrant6_p & v3725fe5;
assign v374a044 = hgrant0_p & v39a4d88 | !hgrant0_p & v3777fc5;
assign v8e06bc = hmaster2_p & v3a5fc34 | !hmaster2_p & v376ce77;
assign v373dce8 = hmaster3_p & v375ed69 | !hmaster3_p & v376b1ee;
assign v373cba8 = hbusreq8 & v375a8db | !hbusreq8 & v3a56918;
assign v375ef7b = hmaster1_p & v3a57584 | !hmaster1_p & v3a70f33;
assign ad41f9 = hmaster1_p & v376bd43 | !hmaster1_p & v376ab29;
assign v37786f3 = hbusreq5 & v372cf70 | !hbusreq5 & v377de7f;
assign v3a6fadb = hgrant6_p & v377e13b | !hgrant6_p & !v3761d5a;
assign v3767baa = hmaster1_p & v3736b55 | !hmaster1_p & v3a6d2d3;
assign v3753456 = hbusreq6 & v3769bcb | !hbusreq6 & v3a65d01;
assign v375e0cc = hmaster1_p & v3774a7d | !hmaster1_p & v3a661f3;
assign cc4895 = hgrant6_p & v3a70dbe | !hgrant6_p & v37372dd;
assign v3772a9b = hbusreq0 & v3a70beb | !hbusreq0 & v8455ab;
assign v37425ab = hbusreq5_p & v3730526 | !hbusreq5_p & v375a2a3;
assign v373ffa0 = hbusreq6_p & v3a70055 | !hbusreq6_p & v37487a4;
assign v3a6ebc5 = hbusreq5_p & v37293c3 | !hbusreq5_p & !v3a6fdc0;
assign v3733239 = hmaster1_p & v3a6ff25 | !hmaster1_p & v375a878;
assign v377b3cf = hbusreq6 & v3726a38 | !hbusreq6 & !v8455ab;
assign v3744b07 = hbusreq4 & v372cb44 | !hbusreq4 & v377f73c;
assign v99797a = hbusreq5_p & v3a70145 | !hbusreq5_p & !v374729b;
assign v375ab02 = hgrant4_p & v376fc1c | !hgrant4_p & v3a5b541;
assign v3a6fd76 = hgrant5_p & v3a6c3ac | !hgrant5_p & v2acae79;
assign v3a6fef0 = hlock5 & v3768858 | !hlock5 & v376e0b6;
assign v374be5d = hgrant4_p & v8455ab | !hgrant4_p & !v373e827;
assign v3a6b937 = hbusreq7_p & v3751bdd | !hbusreq7_p & v37645da;
assign v3a57378 = hbusreq2 & v3a6e622 | !hbusreq2 & v8455ab;
assign v3a68e71 = hbusreq6_p & v377834b | !hbusreq6_p & v3a6f8de;
assign v37518ac = hmaster1_p & v3a5ead4 | !hmaster1_p & v3743788;
assign v374bf0f = hbusreq5_p & v3755ffc | !hbusreq5_p & v37478bc;
assign v375585e = hmaster0_p & v3a71248 | !hmaster0_p & v373b59f;
assign v1e37996 = hbusreq4_p & v3777a9a | !hbusreq4_p & v3a6fcf3;
assign v3a6f520 = hlock4_p & v377af44 | !hlock4_p & !v8455ab;
assign v372b31a = hbusreq5 & v372f0c7 | !hbusreq5 & v3724733;
assign v3772cab = hmaster1_p & v3a6f8d9 | !hmaster1_p & v3757a04;
assign v3a6fa8f = hmaster0_p & v376efaa | !hmaster0_p & v377234d;
assign v372b46a = hmaster3_p & v3a647c6 | !hmaster3_p & v3775a25;
assign v3a593cb = hbusreq2_p & v3751ecb | !hbusreq2_p & !v8455ab;
assign v375e9b2 = hmaster2_p & v8455ab | !hmaster2_p & v373c612;
assign v37c0294 = hmaster2_p & v8455ab | !hmaster2_p & !v372fb2a;
assign v3a6f8dd = hbusreq0_p & v3770993 | !hbusreq0_p & v3744265;
assign v377ae65 = hgrant0_p & v37600af | !hgrant0_p & v373fc30;
assign v376d817 = hbusreq2 & v37678fc | !hbusreq2 & v8455b3;
assign v377e915 = hbusreq5_p & v3766cfb | !hbusreq5_p & v3a7005b;
assign v37513e6 = hlock7 & v377d15d | !hlock7 & v3a5ab7b;
assign v3a6bc32 = hmaster1_p & v376dea1 | !hmaster1_p & v3728d9c;
assign v377b3c4 = hmaster2_p & v2ff9190 | !hmaster2_p & v37630f1;
assign v375db2a = hlock3_p & v374306c | !hlock3_p & v3a6ffae;
assign v3770578 = hbusreq3_p & v3a58218 | !hbusreq3_p & v373cca3;
assign v3749f78 = hlock6_p & v3a676d6 | !hlock6_p & v377395f;
assign v373e15b = hmaster2_p & v372f349 | !hmaster2_p & v38099c1;
assign v373d0d1 = hbusreq4 & v377e29a | !hbusreq4 & v375da10;
assign v357733c = hgrant6_p & v8455ab | !hgrant6_p & v3a6c636;
assign v376d1e2 = hbusreq0_p & v3740171 | !hbusreq0_p & v8455ab;
assign v376d9c6 = hbusreq4_p & v8455bb | !hbusreq4_p & v3a6573d;
assign v3749529 = hlock0_p & v8455ab | !hlock0_p & v3765b88;
assign v375d0d2 = hmaster2_p & v3a6f42e | !hmaster2_p & v37541ff;
assign v373edc8 = hbusreq3_p & v37697e2 | !hbusreq3_p & v372cc25;
assign v3730986 = hgrant4_p & v3748d67 | !hgrant4_p & cecaa5;
assign v373b287 = jx0_p & v8455cd | !jx0_p & v8455ab;
assign v375ef36 = hlock0_p & v373fe5e | !hlock0_p & !v3739faf;
assign v374006f = hmaster2_p & v3777cfc | !hmaster2_p & v3a5bdd2;
assign v3a6d4f9 = hbusreq6_p & v374faa9 | !hbusreq6_p & v373fc8a;
assign v3a6d64e = hbusreq5 & v3776039 | !hbusreq5 & v3a635ea;
assign v3735fb3 = hmaster1_p & v37763bd | !hmaster1_p & v3746069;
assign v3770c98 = hbusreq8_p & v3727f69 | !hbusreq8_p & v3806dc8;
assign v3747cf5 = hlock0_p & v3a703df | !hlock0_p & v375ecc7;
assign v375f3bc = hgrant7_p & v3a54271 | !hgrant7_p & v374bbca;
assign v375a6a7 = hgrant4_p & v3764049 | !hgrant4_p & v3a5ec7a;
assign v3a66120 = hbusreq5_p & v3775a9f | !hbusreq5_p & v3769740;
assign v3767ea6 = hlock6_p & v3a709ea | !hlock6_p & v3a5db8a;
assign v3a6f169 = hlock0_p & v372dadb | !hlock0_p & v3a6ec06;
assign v37284f3 = hmaster0_p & v3776fb8 | !hmaster0_p & v35b774b;
assign v3739c14 = hgrant4_p & v377b6ce | !hgrant4_p & v372562b;
assign v377cdbe = hlock4 & v38072fd | !hlock4 & v377e2ae;
assign v3a64056 = hgrant6_p & v8455ab | !hgrant6_p & v3769f84;
assign v3757d70 = hbusreq6 & v3756e01 | !hbusreq6 & v372ef16;
assign v3a6814a = hlock4_p & v372391f | !hlock4_p & v375e60f;
assign v374617d = hgrant6_p & v8455ab | !hgrant6_p & v377ce51;
assign v3a70367 = hbusreq7 & v372ad15 | !hbusreq7 & v8455ab;
assign v377c02f = hmaster1_p & v3740a1b | !hmaster1_p & v3727dc9;
assign v3a70143 = hbusreq5_p & v373c372 | !hbusreq5_p & v3a6eb3d;
assign v3a6b475 = hready_p & v3a57b11 | !hready_p & v3146177;
assign v375cbcb = hmaster0_p & v3a6eeb0 | !hmaster0_p & v3a7004b;
assign v37289ee = hlock3 & v3a6ffcf | !hlock3 & v3739b17;
assign v37515a1 = hlock7 & v3a701ee | !hlock7 & v375d95f;
assign v3a704f3 = hbusreq2 & v373a841 | !hbusreq2 & v8455ab;
assign v37236b3 = hmaster0_p & v3a6fa13 | !hmaster0_p & !v37733e3;
assign v3a7162a = hmaster2_p & v8455ab | !hmaster2_p & v3761553;
assign v37674f6 = hgrant4_p & v3a62a6d | !hgrant4_p & v3750c52;
assign v375be54 = hmaster0_p & v3a7157b | !hmaster0_p & v3a6ab7f;
assign v3730568 = hmaster1_p & v3759b20 | !hmaster1_p & v37440e4;
assign v3733b4b = hmaster2_p & v3a70ca8 | !hmaster2_p & v8455ab;
assign v3732c56 = hbusreq8 & v3774bed | !hbusreq8 & v375e958;
assign v3724577 = hgrant2_p & v3730e2e | !hgrant2_p & v3a71061;
assign v373cae8 = hmaster0_p & v376e580 | !hmaster0_p & v8455ab;
assign v3a706e1 = hmaster2_p & baec07 | !hmaster2_p & !v8455ab;
assign v372d764 = hbusreq8_p & v3a5d0d3 | !hbusreq8_p & v8455ab;
assign v372e4b3 = hgrant2_p & v3a6b873 | !hgrant2_p & v3a671a2;
assign v3a5a323 = hgrant5_p & v3a70578 | !hgrant5_p & v373706e;
assign v37263c3 = hlock5_p & v3760eb8 | !hlock5_p & v374fc20;
assign v375139d = hbusreq6_p & v3743d23 | !hbusreq6_p & v8455ab;
assign v373f950 = hbusreq4 & v8455b0 | !hbusreq4 & v375d616;
assign v3a6e3bb = hgrant3_p & v3771d77 | !hgrant3_p & v3749e48;
assign v3a56f2e = jx1_p & v37296ca | !jx1_p & v372e351;
assign v37368c8 = hmaster2_p & v3a7116b | !hmaster2_p & v8455ab;
assign v3a70713 = hbusreq8 & v37379a2 | !hbusreq8 & v3765e47;
assign v376c313 = hbusreq7 & v3737200 | !hbusreq7 & v3a70040;
assign v23fde7b = hbusreq5_p & v3a64a83 | !hbusreq5_p & v8455ab;
assign v3a6efad = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a641d5;
assign v3a6143f = hbusreq4_p & v377e70d | !hbusreq4_p & v377d6f9;
assign v3a70021 = hbusreq5_p & v3766786 | !hbusreq5_p & v8455ab;
assign v37339b7 = hbusreq7 & v37730b3 | !hbusreq7 & v3737808;
assign v9de657 = hmaster2_p & v37406d2 | !hmaster2_p & v3a6f993;
assign v3774859 = hbusreq7 & v3a70eea | !hbusreq7 & !v8455ab;
assign v374f630 = hgrant2_p & v3a680b9 | !hgrant2_p & v3a71231;
assign v3a5ada2 = jx2_p & v3735468 | !jx2_p & v3a56a52;
assign v37777ba = hgrant6_p & v3a6f5d2 | !hgrant6_p & v86d306;
assign v37434eb = hgrant5_p & v8455ab | !hgrant5_p & v3a705ea;
assign v3755a96 = hmaster0_p & v3a7050e | !hmaster0_p & !v375f664;
assign v37656be = hmaster0_p & v37717ea | !hmaster0_p & v3723be4;
assign v3a6fe18 = hgrant4_p & v8455ab | !hgrant4_p & v3757772;
assign v3a63b7a = hbusreq5 & v37229e0 | !hbusreq5 & v375d9df;
assign v376d9d4 = hbusreq3 & v3a63bbc | !hbusreq3 & v8455ab;
assign v3a566c1 = hbusreq5_p & v3a71118 | !hbusreq5_p & v3a70924;
assign v373de8a = hgrant6_p & v2acaf72 | !hgrant6_p & !v3761b75;
assign d3af9c = hbusreq0_p & v373997b | !hbusreq0_p & v37738fc;
assign v37494ce = hmaster0_p & v3a70dd9 | !hmaster0_p & v3757ffa;
assign v3763252 = hlock0 & v3a64af7 | !hlock0 & v3a7002a;
assign v376aa57 = hmaster2_p & v376a6f1 | !hmaster2_p & v375058e;
assign v3754fac = hbusreq6 & v377961f | !hbusreq6 & v8455ab;
assign v3a6cab1 = hbusreq2 & v37453d8 | !hbusreq2 & v3773ee6;
assign v3a5d80f = hbusreq4 & v3738745 | !hbusreq4 & v8455ab;
assign v373e1a6 = hgrant3_p & v374551a | !hgrant3_p & v8455ab;
assign v373d8e4 = jx0_p & v376cab5 | !jx0_p & v376a74a;
assign v3a709b4 = hmaster2_p & v3a63777 | !hmaster2_p & v3747302;
assign v3757740 = hmaster2_p & v3a66dc0 | !hmaster2_p & !v8455ab;
assign v3761f74 = hbusreq7_p & v3a6b4db | !hbusreq7_p & v3a571e5;
assign v3770b73 = hbusreq5_p & v37432cd | !hbusreq5_p & v37320bf;
assign v3766f30 = jx0_p & v3a658d5 | !jx0_p & v3a5b642;
assign v374e056 = hlock6_p & v37395e6 | !hlock6_p & v8455e7;
assign v37729bf = hmaster2_p & v3a70059 | !hmaster2_p & !v3760700;
assign v3a70257 = hgrant2_p & v3758472 | !hgrant2_p & !v3742cde;
assign v376a052 = hbusreq5 & v377682b | !hbusreq5 & v3756737;
assign v37667e4 = hbusreq7_p & v3733e5a | !hbusreq7_p & v377974f;
assign v373db25 = hbusreq7 & v3a6eb9e | !hbusreq7 & v376bc9b;
assign v3779736 = hgrant4_p & v3a695c9 | !hgrant4_p & !v3778464;
assign v374dbf7 = hlock5 & v3a5dc67 | !hlock5 & v37548f5;
assign v3a7132e = hmaster1_p & v3a5bf5f | !hmaster1_p & v3738dc0;
assign v3a71373 = hbusreq5_p & v374326f | !hbusreq5_p & v3a6f537;
assign v3777bfc = hmaster0_p & v3a567b7 | !hmaster0_p & v3758c58;
assign v3770e30 = hbusreq6 & v3a70fd2 | !hbusreq6 & v3a7162d;
assign v3a53ae0 = hmaster0_p & v3a6f942 | !hmaster0_p & v3727889;
assign v3766a64 = hbusreq5_p & v3a70796 | !hbusreq5_p & v2acb068;
assign v3a6addc = hbusreq7 & v3745d0a | !hbusreq7 & v8455ab;
assign v376419b = hlock8_p & v3a558dc | !hlock8_p & v8455ab;
assign v3a70101 = hmaster0_p & v37365ce | !hmaster0_p & v3a70f9c;
assign v3778354 = jx0_p & v375efe8 | !jx0_p & v372fe64;
assign v3a68789 = hbusreq7 & v3a5f5db | !hbusreq7 & v3a7006e;
assign v3a6fcaa = hlock0_p & v8455ab | !hlock0_p & v3a6900c;
assign v3724c9c = hmaster2_p & v3a619c0 | !hmaster2_p & v376d856;
assign v372e611 = hbusreq8 & v3a71119 | !hbusreq8 & v3a710bb;
assign v3a6f2b7 = hmaster1_p & v3a6e581 | !hmaster1_p & v376704f;
assign v3807a4a = hlock5 & v372c863 | !hlock5 & v3a5ddaa;
assign v1e37b48 = hmaster1_p & v3a62a6d | !hmaster1_p & v375750d;
assign v3a6f3ac = hmaster0_p & v3747a36 | !hmaster0_p & v375449f;
assign v375c2e6 = hbusreq8_p & v374726f | !hbusreq8_p & v3a6fba2;
assign v3729263 = hmaster0_p & v3774b2b | !hmaster0_p & v375d3fd;
assign v3a6a1e9 = hbusreq2_p & v3755aef | !hbusreq2_p & v373bb0f;
assign v3a5902d = hbusreq7_p & v3767704 | !hbusreq7_p & v3a6bde4;
assign v37672c8 = hlock4 & v3a5c127 | !hlock4 & v374bc27;
assign v3a7165e = hbusreq8 & v3a6a084 | !hbusreq8 & v37305e3;
assign v37659e4 = hmaster2_p & v3725198 | !hmaster2_p & v3736ded;
assign v3733c82 = hmaster1_p & v376ee65 | !hmaster1_p & v3a67524;
assign v2acb5a2 = hmastlock_p & v37464c8 | !hmastlock_p & v8455ab;
assign v373f7ef = hmaster0_p & v3a6992f | !hmaster0_p & !v3a64977;
assign v3746641 = hgrant4_p & v3a70912 | !hgrant4_p & v372a3af;
assign v373f0d2 = hmaster1_p & v37737b9 | !hmaster1_p & v37709ec;
assign v375f69e = hmaster2_p & v3a61a7f | !hmaster2_p & v3723b5b;
assign v2092a68 = hmaster0_p & v3a63ee6 | !hmaster0_p & v3a6f3b9;
assign v3750b8c = hmaster2_p & v372e443 | !hmaster2_p & v3a655e9;
assign v37542d8 = hbusreq5_p & v37720f9 | !hbusreq5_p & v3749004;
assign v3767b88 = hbusreq4_p & v3a58b8f | !hbusreq4_p & v3763b0a;
assign v376b561 = hmaster2_p & v3a709ee | !hmaster2_p & v35772a6;
assign v3a7037c = hlock0_p & v37757e0 | !hlock0_p & v8455b0;
assign v3a607fa = hmaster0_p & v8455b0 | !hmaster0_p & v3729360;
assign v3a7088d = hgrant6_p & v374a664 | !hgrant6_p & v3773a45;
assign v37652eb = hbusreq0 & v37746ea | !hbusreq0 & v377c31d;
assign v3a70a3c = hbusreq3 & v3a63805 | !hbusreq3 & v8455ab;
assign v3a5eb8f = hbusreq5_p & v3736ad7 | !hbusreq5_p & v373d42f;
assign v3a60276 = hgrant5_p & v3740052 | !hgrant5_p & v3722fb7;
assign v3731737 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3a69bfd;
assign v37710c7 = hgrant4_p & v375e99f | !hgrant4_p & v37435a8;
assign v3775721 = hmaster2_p & v375a67c | !hmaster2_p & !v3a70fec;
assign v37775dd = hbusreq5 & v372f202 | !hbusreq5 & v3738ea9;
assign v37280c8 = hbusreq2_p & v3a705ad | !hbusreq2_p & !v37450cb;
assign v377dcbc = hgrant3_p & v8455bd | !hgrant3_p & v3769806;
assign v375d2ee = hmaster1_p & v3a5d327 | !hmaster1_p & v3748b0e;
assign v375a7bd = stateG10_1_p & v35772a6 | !stateG10_1_p & v3762453;
assign v374ac2e = hmaster0_p & be181b | !hmaster0_p & v38087ba;
assign v3734b20 = hmaster2_p & v3a5e291 | !hmaster2_p & !v375fd29;
assign v3a570a0 = jx1_p & v3a60ef2 | !jx1_p & v3760317;
assign v3a70945 = hready_p & v377b221 | !hready_p & v39378d6;
assign v3765e46 = hbusreq1_p & v8455ab | !hbusreq1_p & v3a6a939;
assign v8cdbc1 = hgrant6_p & v3a598a9 | !hgrant6_p & v373621d;
assign v3778464 = hbusreq4_p & v377594d | !hbusreq4_p & v373d72e;
assign v3a6ff56 = hbusreq7_p & v37546c9 | !hbusreq7_p & v374df25;
assign v377ea3c = hbusreq5 & v375fbf2 | !hbusreq5 & !v374e0f6;
assign v3731b53 = hmaster1_p & v3a6d7f2 | !hmaster1_p & v3a5c816;
assign v3a70f25 = jx1_p & v3767c03 | !jx1_p & v3a70ec4;
assign v3767b5a = hmaster1_p & v3a635ea | !hmaster1_p & v3a6d0af;
assign v3a6c7ef = hbusreq0 & v3750002 | !hbusreq0 & c7355c;
assign v3738251 = hgrant4_p & v1e37b99 | !hgrant4_p & v3a68607;
assign v3a6f37c = hbusreq2 & v3a6dc08 | !hbusreq2 & adf78a;
assign v374f6c0 = hgrant5_p & v3745fd1 | !hgrant5_p & v372da7e;
assign v1e3795b = hgrant6_p & v3a696ed | !hgrant6_p & v3774b56;
assign v3a6fdc3 = hbusreq6_p & v37272ed | !hbusreq6_p & !v372df2a;
assign c0b4d9 = hbusreq3_p & v3a6f748 | !hbusreq3_p & v373132b;
assign v1e37ca9 = hbusreq0_p & v374c936 | !hbusreq0_p & v373b710;
assign v37650e4 = hmaster1_p & v374b7f6 | !hmaster1_p & v375b400;
assign v3a6b4de = hlock8 & v376b44a | !hlock8 & v3a5511c;
assign v3a6f8a9 = hbusreq5 & v374f359 | !hbusreq5 & v3a6fa7c;
assign v3a7076d = hbusreq4_p & v3a5dde7 | !hbusreq4_p & v38097a9;
assign v372f59c = hmaster2_p & v374b3f8 | !hmaster2_p & v3722c80;
assign v376b199 = hgrant6_p & v8455ab | !hgrant6_p & v37753da;
assign v3a5efb8 = hbusreq4_p & v3a7020e | !hbusreq4_p & v3a713c8;
assign v377f2bb = hmaster1_p & v374f0c1 | !hmaster1_p & v3a58761;
assign v374f9ce = hbusreq0 & v37513bc | !hbusreq0 & v3777e0e;
assign v375a288 = hlock0_p & v37738fc | !hlock0_p & !v39a4ca8;
assign v376eeb3 = hlock7 & v3a70de5 | !hlock7 & v374a79e;
assign v3a6869d = hmaster1_p & v3a6373e | !hmaster1_p & v3729ca6;
assign v3747193 = hlock0 & v37285eb | !hlock0 & v3778cdb;
assign v37450a5 = hlock4_p & v3a63e82 | !hlock4_p & !v35772a6;
assign v38064a2 = hbusreq6 & v3777a6c | !hbusreq6 & v375da95;
assign v3724bdd = hbusreq7_p & v3a6effd | !hbusreq7_p & v3738aa6;
assign v3a6e40f = hbusreq7_p & v3a67182 | !hbusreq7_p & v3a5aff3;
assign v374ecd5 = hbusreq4_p & v8455ab | !hbusreq4_p & v3a6a939;
assign v374ab76 = hlock8_p & v3a70f15 | !hlock8_p & !v8455ab;
assign v37399d4 = hmaster1_p & v3a6ccc4 | !hmaster1_p & v3a7055c;
assign v3a5ba7f = hmaster2_p & v8455ab | !hmaster2_p & v374036a;
assign v373dafc = hgrant0_p & v372b931 | !hgrant0_p & v375323b;
assign v3736d87 = hbusreq8_p & v372e0fc | !hbusreq8_p & v374897d;
assign v3806b35 = hgrant3_p & v38070c1 | !hgrant3_p & v37508a4;
assign v373690a = hbusreq4_p & v3739f0e | !hbusreq4_p & cecaa5;
assign v3a5e9d3 = hlock1 & v8c0e15 | !hlock1 & v3a593ee;
assign ad187c = hmaster1_p & v375c791 | !hmaster1_p & v3753542;
assign v3a5ac8b = hbusreq5 & v3a6a990 | !hbusreq5 & v8455ab;
assign v3a54fb2 = hburst0_p & v8455ab | !hburst0_p & !v8455d7;
assign v37787c1 = hgrant4_p & v372f346 | !hgrant4_p & v37756ab;
assign v3730d6c = hmaster2_p & v375069a | !hmaster2_p & v37284d5;
assign v3a69ead = hmaster0_p & v372a966 | !hmaster0_p & v8455ab;
assign v375ea13 = hmaster0_p & v3772775 | !hmaster0_p & v2678bee;
assign v375bdcc = hmaster2_p & v375166c | !hmaster2_p & v372a85f;
assign v3a6f2ba = hmaster0_p & v3758b78 | !hmaster0_p & v37733e3;
assign v3a706be = hmaster0_p & v3a58218 | !hmaster0_p & v3a6f249;
assign v375dc63 = hbusreq8_p & v372c4cd | !hbusreq8_p & v3a5a807;
assign v373a759 = hmaster2_p & v3747b15 | !hmaster2_p & v373e38a;
assign v3741816 = hlock7_p & v372bb35 | !hlock7_p & v374f832;
assign v374b0c1 = hbusreq3 & v3773b23 | !hbusreq3 & v8455ab;
assign v372ba1c = hgrant4_p & v8455c2 | !hgrant4_p & v3a70a81;
assign v3a6f255 = hmaster2_p & v3766484 | !hmaster2_p & v375199d;
assign v2acaedd = hmaster0_p & v3a6e5f0 | !hmaster0_p & v3a7004f;
assign v37429c2 = hmaster2_p & v3751913 | !hmaster2_p & v8455ab;
assign v3a70e19 = hbusreq4 & v372d336 | !hbusreq4 & v37519ea;
assign v373cb9c = stateG2_p & v3a5a496 | !stateG2_p & v37643ee;
assign v374c75e = hbusreq4_p & v3757f01 | !hbusreq4_p & v377ceea;
assign v3a6fa5d = hmaster0_p & v37430c6 | !hmaster0_p & v374ba88;
assign v3a63f66 = hbusreq5 & v3a57444 | !hbusreq5 & v8455ab;
assign v375a412 = hmaster0_p & v8455ab | !hmaster0_p & v3a70f4a;
assign v373d0e1 = stateG10_1_p & v3a6e7b3 | !stateG10_1_p & v3a69a06;
assign v376085a = hbusreq0 & v377910a | !hbusreq0 & v3a572e9;
assign v376b015 = hmaster2_p & v377097a | !hmaster2_p & v8455ab;
assign v372f478 = hlock5_p & v3761071 | !hlock5_p & v377843d;
assign v377b205 = hbusreq7 & v373e07e | !hbusreq7 & v3746f9d;
assign v89a0d1 = hbusreq0 & v3a6b41e | !hbusreq0 & v3a7149e;
assign v3a71008 = hgrant5_p & v3a6a872 | !hgrant5_p & v372f89e;
assign v376d7a5 = hmaster2_p & v373a4e4 | !hmaster2_p & v3a70fb2;
assign v3a5d2f1 = hready_p & v3a62615 | !hready_p & v374151e;
assign v372ba66 = hmaster0_p & v375eee3 | !hmaster0_p & v374c78e;
assign v3776be5 = hmaster1_p & v3725198 | !hmaster1_p & v3a63e68;
assign v3751f46 = hbusreq6 & v373ee80 | !hbusreq6 & v8455ab;
assign v377a291 = hbusreq2_p & v3748797 | !hbusreq2_p & v3724069;
assign v38092b4 = hlock6_p & v3a5b5d3 | !hlock6_p & v3a658bf;
assign v376fc77 = hlock4 & v3a707aa | !hlock4 & v3a5af1e;
assign v376c69d = hlock7 & v373b0f3 | !hlock7 & v3772a57;
assign v3807113 = hbusreq0 & v373b14a | !hbusreq0 & v3a60b96;
assign v3a711b4 = hbusreq8 & v375be90 | !hbusreq8 & v376382f;
assign v374c3d0 = hgrant6_p & v2ff9348 | !hgrant6_p & v8455ab;
assign v3752dd0 = hbusreq4_p & v37339c8 | !hbusreq4_p & v8455ab;
assign v377d97d = hlock7 & v375fc73 | !hlock7 & v3a70727;
assign v3764978 = hbusreq6 & v3a57325 | !hbusreq6 & v8455ab;
assign v3774161 = hmaster2_p & v380760a | !hmaster2_p & v3a6fac9;
assign v3a57891 = hbusreq5_p & a2a6f3 | !hbusreq5_p & v373346a;
assign v3733f28 = hbusreq4 & v3a6dc08 | !hbusreq4 & v3730ffe;
assign v3728738 = hmaster0_p & v3760513 | !hmaster0_p & v3738e6e;
assign v3759f4c = hlock3_p & v3a70f80 | !hlock3_p & v3a6eb83;
assign v376f0c1 = hbusreq3_p & v374af6a | !hbusreq3_p & v37410d9;
assign v373d8d8 = hmaster0_p & v3750c50 | !hmaster0_p & v373da59;
assign v372d3e8 = hbusreq2_p & v3723676 | !hbusreq2_p & v3a63bdb;
assign v3a6eed1 = hbusreq7_p & v3767dd2 | !hbusreq7_p & v377c487;
assign v3757e2f = hgrant4_p & v3a6ff32 | !hgrant4_p & v374f1ae;
assign v3a60bbf = hbusreq6_p & v3a70a92 | !hbusreq6_p & v3753317;
assign v3731df6 = hbusreq2 & v374b70d | !hbusreq2 & v8455ab;
assign v3724c55 = hbusreq4_p & v8455ab | !hbusreq4_p & v37665bf;
assign v376d306 = hbusreq4_p & v376ac74 | !hbusreq4_p & v8455ab;
assign v3a6fd53 = hmaster2_p & v374b992 | !hmaster2_p & v374ac60;
assign v376f261 = hgrant7_p & v372d8bd | !hgrant7_p & v373917f;
assign v372ebc8 = hmaster0_p & v372c18a | !hmaster0_p & v8455ab;
assign v3744806 = hmaster0_p & v8455ab | !hmaster0_p & v373165b;
assign v373e267 = hmaster2_p & v3a704c7 | !hmaster2_p & v377edba;
assign v374aec2 = hgrant4_p & v3a7024f | !hgrant4_p & v3a6b51f;
assign v3a66584 = hbusreq6_p & v3a69df1 | !hbusreq6_p & v37728d3;
assign v37627ec = hbusreq5_p & v3739904 | !hbusreq5_p & v377ea20;
assign v376c4a9 = hbusreq4_p & v372f3f1 | !hbusreq4_p & v23fd96e;
assign v3763c0a = hbusreq0 & v3756018 | !hbusreq0 & v3a5acd5;
assign v3776337 = hmaster1_p & v373013d | !hmaster1_p & v3a68317;
assign v376a867 = hgrant2_p & v8455ab | !hgrant2_p & v3744796;
assign v3a6073f = hmaster0_p & v3a708c3 | !hmaster0_p & v3773e17;
assign v3a7136a = hlock4 & v3770d41 | !hlock4 & v374ad30;
assign v376b99f = hgrant6_p & v3750d06 | !hgrant6_p & v377903f;
assign v3746265 = hbusreq2_p & v3751734 | !hbusreq2_p & v3a59409;
assign v3a6f641 = hgrant4_p & v8455ab | !hgrant4_p & v373e814;
assign v3a63368 = hgrant5_p & v37492d2 | !hgrant5_p & v376c31d;
assign v3725310 = hbusreq0_p & v37376c8 | !hbusreq0_p & v8455ab;
assign v375ede6 = hmaster0_p & v3a6e4ec | !hmaster0_p & v37458ca;
assign v3751862 = hbusreq4 & v3730ba6 | !hbusreq4 & !v3a640a0;
assign v372e244 = hbusreq6_p & v3a654c1 | !hbusreq6_p & v376bb26;
assign v37280b7 = hbusreq5 & v373324d | !hbusreq5 & v3758ee1;
assign v3772c8e = hmaster1_p & v3a700d9 | !hmaster1_p & v3a70606;
assign v374a9fa = hgrant5_p & v375c67c | !hgrant5_p & v3728d28;
assign v3748d17 = hgrant2_p & v8455ab | !hgrant2_p & v3a533ae;
assign v377903c = hburst0 & v372fe05 | !hburst0 & v376acf0;
assign v2889709 = hmaster2_p & v3777da6 | !hmaster2_p & v3773fc7;
assign v37799ca = hmaster2_p & v37bfc35 | !hmaster2_p & v3a6908b;
assign v3a66b26 = hgrant0_p & v37368d3 | !hgrant0_p & !v3776a6e;
assign v377085b = hlock0 & v3a5f9e6 | !hlock0 & v374a297;
assign v3726eea = hmaster0_p & v372c064 | !hmaster0_p & v8455ab;
assign v374b8ad = hgrant2_p & v377182c | !hgrant2_p & v37721b2;
assign v3a6f5a5 = hmaster2_p & v8455b5 | !hmaster2_p & v37c0382;
assign v3a70b08 = hgrant0_p & v3a6fcaa | !hgrant0_p & v374037a;
assign v8455d1 = hbusreq8_p & v8455ab | !hbusreq8_p & !v8455ab;
assign v37233d2 = hbusreq4 & v3a6db1a | !hbusreq4 & v3a64af7;
assign v3747465 = hmaster1_p & v376bd2c | !hmaster1_p & v3a70071;
assign v3a5f485 = hbusreq2_p & v3729991 | !hbusreq2_p & v375c1d1;
assign v3a6ab69 = hlock6 & v3760d8d | !hlock6 & v376cad6;
assign v3a65e17 = hmaster2_p & v373561e | !hmaster2_p & v3778091;
assign v374fcde = hgrant5_p & v375d7bc | !hgrant5_p & v3a714da;
assign v373ec72 = hlock6_p & v37681fa | !hlock6_p & v3a7092a;
assign v3a70f9a = hmaster0_p & v3748db2 | !hmaster0_p & v3732938;
assign v373ab9e = hgrant6_p & v3a57b60 | !hgrant6_p & v3a6fff9;
assign v3745075 = hbusreq0_p & v3a63805 | !hbusreq0_p & v8455b0;
assign v3a6999c = hlock3_p & v37396eb | !hlock3_p & !v8455ab;
assign v3773200 = hbusreq4_p & v37504eb | !hbusreq4_p & v8455ab;
assign v372601c = hmaster0_p & v3777b00 | !hmaster0_p & v3a70f41;
assign v374b21a = hbusreq6 & v3723430 | !hbusreq6 & v8455ab;
assign v37273f4 = hmaster1_p & v37438ba | !hmaster1_p & v3754025;
assign v372ad15 = hgrant5_p & v3767852 | !hgrant5_p & v37400fe;
assign v3765d94 = jx0_p & v3a57f18 | !jx0_p & v375d34f;
assign v3a715c5 = hmaster2_p & v8455ab | !hmaster2_p & v3a5a01b;
assign v3a70bf0 = hmaster1_p & v374a8e2 | !hmaster1_p & v8455ab;
assign v3a70923 = hbusreq3_p & v3a70eb6 | !hbusreq3_p & v3a63621;
assign v374cda0 = hgrant6_p & v8455ab | !hgrant6_p & v3a6ad04;
assign v3a711dd = hgrant2_p & v3a62a6d | !hgrant2_p & v375af3c;
assign v377f883 = hbusreq8 & v3774641 | !hbusreq8 & v3a55e3c;
assign v37375e4 = hgrant6_p & v8455ca | !hgrant6_p & v3730fb0;
assign v376c80f = hbusreq4 & v39eb4cb | !hbusreq4 & v3a5b6de;
assign v3a70b53 = stateA1_p & v8455ab | !stateA1_p & !v37314db;
assign v3a6fc2f = hbusreq6_p & v8455bf | !hbusreq6_p & v374c163;
assign v3a5980d = hbusreq1_p & v3a6fde8 | !hbusreq1_p & v8455ab;
assign v3a6eefe = stateG10_1_p & v8455ab | !stateG10_1_p & v3745b36;
assign v375e8d2 = hmaster1_p & v3a57584 | !hmaster1_p & v374d8c9;
assign v3a6ccd6 = hbusreq6_p & v373cdb0 | !hbusreq6_p & v37311de;
assign v3a6450a = hmaster1_p & v3739702 | !hmaster1_p & v8455e7;
assign v3748256 = hgrant5_p & v8455ab | !hgrant5_p & v3738263;
assign v3731749 = hbusreq6 & v3a6f806 | !hbusreq6 & v37453d7;
assign v3744693 = hlock0_p & v3758cec | !hlock0_p & !v3744710;
assign v3723aea = hgrant1_p & v372a837 | !hgrant1_p & v37665bf;
assign v3743910 = hmaster2_p & v377234d | !hmaster2_p & v3773200;
assign v3a6e844 = hbusreq5_p & v3773340 | !hbusreq5_p & v3a708d6;
assign v3a56ccf = hlock0_p & v37457fb | !hlock0_p & !v39a5381;
assign v3739e0d = hgrant7_p & v8455ab | !hgrant7_p & v3766126;
assign v3770993 = hbusreq1_p & v3a70c73 | !hbusreq1_p & !v9dc858;
assign v3727960 = hbusreq5 & v292554f | !hbusreq5 & v376784b;
assign v372cb77 = hbusreq6 & v373081f | !hbusreq6 & v3723e1f;
assign v372cd65 = hbusreq5 & v3a57ebf | !hbusreq5 & v3a55eda;
assign v3769e01 = hbusreq5_p & v376fbff | !hbusreq5_p & v8455ab;
assign v3757afc = hmaster1_p & v374ffd5 | !hmaster1_p & !v3a64641;
assign v373e2f9 = hmaster2_p & v3a68426 | !hmaster2_p & v3725410;
assign v3a6fad0 = stateA1_p & v3a6efc9 | !stateA1_p & v1e37481;
assign v3809399 = hgrant2_p & v3778ed4 | !hgrant2_p & !v8455ab;
assign v376dd8b = hbusreq8_p & v3a7067d | !hbusreq8_p & v3a6ef96;
assign v37257c8 = hbusreq2_p & v3a6106c | !hbusreq2_p & v374e606;
assign v3748a16 = hmaster0_p & v372cf1f | !hmaster0_p & v8455ab;
assign v376486a = hbusreq5_p & v3727c3c | !hbusreq5_p & v23fd799;
assign v8455ef = hgrant3_p & v8455ab | !hgrant3_p & !v8455ab;
assign v1e37d35 = hbusreq5 & v2acaf4f | !hbusreq5 & v8455ab;
assign v3a6f290 = hmaster1_p & v3749ba6 | !hmaster1_p & !v37421bd;
assign v3a6ff82 = hbusreq0 & v373a90e | !hbusreq0 & v3a709d2;
assign v3a6f032 = hbusreq3_p & v375bdd4 | !hbusreq3_p & v3744f35;
assign v3a5e2a9 = hbusreq5 & v37534c6 | !hbusreq5 & v8455ab;
assign v376144f = hbusreq2 & v3723c0d | !hbusreq2 & v3748797;
assign v3759886 = hbusreq4 & v8455e7 | !hbusreq4 & v8455ab;
assign v37429e5 = hbusreq4_p & v3747302 | !hbusreq4_p & v37485ce;
assign v373f488 = hbusreq4_p & v3746683 | !hbusreq4_p & v3a68d49;
assign v376e9c5 = hbusreq6 & v3a67967 | !hbusreq6 & v8455ab;
assign v3746d49 = hmaster2_p & v373d27f | !hmaster2_p & v3746641;
assign v3a6452e = hmaster2_p & v374f9c6 | !hmaster2_p & v37716ca;
assign v3758f6d = hgrant3_p & v35b7299 | !hgrant3_p & v37619b8;
assign v3a5923c = hgrant3_p & v94ea62 | !hgrant3_p & v8455ab;
assign v3a5b451 = hbusreq0_p & v35772a5 | !hbusreq0_p & !v377c6b3;
assign c4dd17 = hlock5_p & v3a705f5 | !hlock5_p & v3a6fdee;
assign v3a6e47f = hlock3_p & v3740349 | !hlock3_p & v3a6c355;
assign v3725e33 = hmaster1_p & v373b7be | !hmaster1_p & b52e7d;
assign ae60a0 = hbusreq8 & v3a6f5e9 | !hbusreq8 & v373ea00;
assign v3a6f78f = hbusreq5_p & v3736e12 | !hbusreq5_p & v3a5e9e9;
assign be145a = hmaster2_p & v3a71678 | !hmaster2_p & v8455ab;
assign v3746cc0 = hbusreq4_p & v3748797 | !hbusreq4_p & v3749655;
assign v3749f94 = hmaster0_p & v37548c4 | !hmaster0_p & b0e59c;
assign v3a55ba9 = hgrant3_p & v8455ab | !hgrant3_p & v3733e88;
assign v3a6f03e = hlock0 & v3731230 | !hlock0 & v376b5ad;
assign v3761497 = hbusreq8_p & v3755ab8 | !hbusreq8_p & v3a6a87d;
assign v373f63e = hgrant2_p & v3a6b3df | !hgrant2_p & v37538e4;
assign v3770bd5 = hgrant4_p & v3766ff1 | !hgrant4_p & v3a61739;
assign v325c94d = hbusreq5_p & v375398e | !hbusreq5_p & v372545e;
assign v3a5eaa1 = hbusreq2_p & v374a70f | !hbusreq2_p & v8455ab;
assign v375820a = hbusreq5 & v37263c3 | !hbusreq5 & v8455ab;
assign v3734062 = hgrant4_p & v3a6bcf9 | !hgrant4_p & v3a705b9;
assign v377598f = hlock0 & v3a708cf | !hlock0 & v3a64cfa;
assign v3761909 = hgrant3_p & v3733dd4 | !hgrant3_p & v3a6fedb;
assign v3726d0c = hbusreq7_p & v376fed4 | !hbusreq7_p & !v377478a;
assign v3a6e4de = hbusreq6_p & a8afe1 | !hbusreq6_p & v3a6fa28;
assign v3a6fff0 = hbusreq6_p & v3a6bf6d | !hbusreq6_p & v8455b7;
assign v375b974 = hgrant3_p & v35b774b | !hgrant3_p & v3a6ebb1;
assign v372b10b = hlock5_p & v377c35c | !hlock5_p & v3779797;
assign v3728c23 = hbusreq6_p & v377ec28 | !hbusreq6_p & v8455ab;
assign v375d149 = hgrant6_p & v3a635ea | !hgrant6_p & aac430;
assign v3764eb2 = hbusreq0 & v375b9e1 | !hbusreq0 & v375564e;
assign v37234c3 = hbusreq2_p & v374fbcf | !hbusreq2_p & !v8455ab;
assign v374dad0 = hmaster2_p & v372c2bf | !hmaster2_p & v37607a7;
assign v3a5bcf5 = hmaster2_p & v3a6f05e | !hmaster2_p & v377df9c;
assign v3a6ebb7 = hready & v3a63621 | !hready & v3a635ea;
assign v3a6bf6d = hbusreq6 & v37533ae | !hbusreq6 & v3a5efb2;
assign v373c239 = hmaster1_p & v37469c4 | !hmaster1_p & v375e9c8;
assign v376d9ed = hbusreq8 & v3a6d401 | !hbusreq8 & v375aa07;
assign v9bbda1 = hbusreq4 & v3767561 | !hbusreq4 & v8455bb;
assign v3a69267 = hmaster0_p & v3731415 | !hmaster0_p & v37420b6;
assign v3772ad5 = hbusreq2 & v3a5600a | !hbusreq2 & v373b3fb;
assign v3a593b0 = hmaster1_p & v376e1fb | !hmaster1_p & v8455ab;
assign v373b667 = hlock7 & v3738087 | !hlock7 & v374fa18;
assign v375166c = hgrant4_p & v373b7c5 | !hgrant4_p & v3a6ef22;
assign v3776e9c = hbusreq4 & v372640f | !hbusreq4 & v8455ab;
assign v375af3c = hgrant3_p & v8455ab | !hgrant3_p & v3a70268;
assign v3a6fc07 = hmaster1_p & v37782c9 | !hmaster1_p & v375bc70;
assign v3727dc9 = hbusreq5_p & v3771971 | !hbusreq5_p & v3764539;
assign v3a70c52 = hbusreq0 & v372c91d | !hbusreq0 & v3a6f817;
assign v3a70fcf = hmaster2_p & v3a56b60 | !hmaster2_p & v37364cf;
assign v372f657 = hbusreq3_p & v375db2a | !hbusreq3_p & v3a6ffae;
assign v37540e7 = hbusreq6 & v3773b7b | !hbusreq6 & v3a635ea;
assign v375c1a7 = hlock8 & v3737808 | !hlock8 & v377f694;
assign v373d11f = hbusreq4_p & v3a6f43e | !hbusreq4_p & v372935c;
assign v373580a = hgrant6_p & v377f21b | !hgrant6_p & v3a70e8d;
assign v3740473 = hgrant3_p & v377dd3b | !hgrant3_p & v372846c;
assign v3a2981b = hgrant3_p & v3759032 | !hgrant3_p & v3a5e02b;
assign v37618e0 = hbusreq3 & v374f307 | !hbusreq3 & v8455b0;
assign v3754b66 = hbusreq0 & v37674c1 | !hbusreq0 & !v8455ab;
assign v3768857 = hbusreq4_p & v1e379d2 | !hbusreq4_p & v3a70cfe;
assign v37670db = hmaster2_p & v3a635ea | !hmaster2_p & v3a6c5ee;
assign v3a5eac0 = hgrant0_p & v3745b32 | !hgrant0_p & v3a5ef59;
assign v372a1ab = hmaster1_p & v3a5fc34 | !hmaster1_p & v377b9a2;
assign v3724c46 = hmaster1_p & v3a61397 | !hmaster1_p & v3773b0f;
assign v37362e9 = hmaster2_p & v3a6fa7a | !hmaster2_p & v376dc26;
assign v37611df = hmaster1_p & v3753eb2 | !hmaster1_p & v1e3733c;
assign v373e748 = hgrant2_p & v3a5c945 | !hgrant2_p & v3a70f19;
assign v3726f76 = hbusreq7_p & v37382ee | !hbusreq7_p & !v3a5a06e;
assign v37392ae = hmaster2_p & v37356b4 | !hmaster2_p & v373ae83;
assign v376f2a5 = hbusreq4_p & v3751acf | !hbusreq4_p & v374f028;
assign v373daac = hlock6_p & v375ef36 | !hlock6_p & !v8455ab;
assign v3774463 = hbusreq5_p & v8455b7 | !hbusreq5_p & v3a5bb85;
assign v3a6acab = hbusreq3_p & v374fa0a | !hbusreq3_p & v3728ca9;
assign v3a707a1 = hbusreq5_p & v3a706be | !hbusreq5_p & v3a573a7;
assign v37520a9 = hbusreq6_p & v372adc8 | !hbusreq6_p & v8455ab;
assign v3a70ecf = locked_p & v3a5e24e | !locked_p & v3a66110;
assign v3a5c127 = hbusreq4 & v374bc27 | !hbusreq4 & v376bade;
assign v3759007 = hgrant4_p & v3a602a4 | !hgrant4_p & v3a6face;
assign v3a6c6ec = hmaster2_p & v3a71416 | !hmaster2_p & v3a71453;
assign v1e37370 = hgrant4_p & v375c7b9 | !hgrant4_p & v377762d;
assign v374835b = hbusreq8 & v3a631d0 | !hbusreq8 & !v373d081;
assign v3a6b372 = hmaster3_p & v376c9a5 | !hmaster3_p & v8455ab;
assign v3732ef8 = jx1_p & v3759ff9 | !jx1_p & v3a708ed;
assign v3736d51 = hbusreq0_p & v37376c8 | !hbusreq0_p & v373f8fb;
assign v3a6fb66 = hbusreq6 & v3a5b037 | !hbusreq6 & v8455ab;
assign v373fe39 = hmaster1_p & v372ca6e | !hmaster1_p & v3743f5b;
assign v372cac6 = hgrant4_p & v3a60c86 | !hgrant4_p & v3a5ec7a;
assign v375444e = hready & v3726dfa | !hready & !v3761480;
assign v376a40c = hbusreq5_p & v3a7115c | !hbusreq5_p & v3a70e16;
assign v3a66aa4 = hbusreq1_p & v3809e5c | !hbusreq1_p & v8455ab;
assign v37625a8 = hlock0_p & v37502b7 | !hlock0_p & v3754b6c;
assign v373abde = hgrant6_p & v8455ab | !hgrant6_p & v3a6687c;
assign v3a65100 = hbusreq7_p & v3a71039 | !hbusreq7_p & v35b708c;
assign v3a71551 = hmaster1_p & v3a6fd19 | !hmaster1_p & !v3a64641;
assign v3a5921b = hbusreq7_p & v3a6dca6 | !hbusreq7_p & v376fe7d;
assign v3739ab4 = hbusreq4_p & v376f56d | !hbusreq4_p & v373df7f;
assign v375f708 = hmaster0_p & v3a58ca1 | !hmaster0_p & !v3733767;
assign v2ff87d3 = hbusreq5_p & v3750a6f | !hbusreq5_p & c2b7ee;
assign v3736dfe = hbusreq7 & a72a7c | !hbusreq7 & v3a703f6;
assign v3730ab2 = hmaster3_p & v373eef9 | !hmaster3_p & v8455dd;
assign v37711e1 = hbusreq2 & v37699f2 | !hbusreq2 & v3a70c74;
assign v3a65436 = hbusreq3_p & v3730cda | !hbusreq3_p & v3777962;
assign v375c8e6 = hbusreq4_p & v376e89b | !hbusreq4_p & v376b88d;
assign v3a6be07 = hbusreq7_p & v374d972 | !hbusreq7_p & v8455d3;
assign v3a6f223 = hbusreq7_p & v373a7f7 | !hbusreq7_p & !v372c335;
assign v3a6080b = hbusreq5 & v3a68904 | !hbusreq5 & v373f14d;
assign v3777fc5 = hbusreq1_p & v375b2e5 | !hbusreq1_p & v3a6e9a4;
assign v376afb3 = hmaster2_p & v374b8fa | !hmaster2_p & v3a59c65;
assign v376f277 = hbusreq2_p & v3a606e8 | !hbusreq2_p & v377affd;
assign v375f777 = hmaster1_p & v3761719 | !hmaster1_p & v3729381;
assign v3768573 = hgrant2_p & v37523f4 | !hgrant2_p & v372fa02;
assign v3745053 = hlock0_p & v3776fa4 | !hlock0_p & v8455ab;
assign v3a713ee = hbusreq2_p & v3743eda | !hbusreq2_p & v37573b9;
assign v374ac72 = hbusreq3_p & v3737c13 | !hbusreq3_p & v3a640c5;
assign v375aca9 = hlock3_p & v374ae3d | !hlock3_p & v37720e5;
assign v37648cd = hlock0 & v37651c2 | !hlock0 & v376ba89;
assign v377e089 = hbusreq3_p & v3751f56 | !hbusreq3_p & v8455ab;
assign a64c20 = hbusreq8_p & v3a709eb | !hbusreq8_p & v37631bf;
assign v3a5a210 = hmaster1_p & v3377b0f | !hmaster1_p & v8b1055;
assign v37723fb = hmaster1_p & v8455d9 | !hmaster1_p & !v8455ab;
assign v3a69391 = hbusreq7 & v375ceb9 | !hbusreq7 & v3740a94;
assign v377546d = hgrant5_p & v8455c6 | !hgrant5_p & v3756091;
assign v3770ff4 = hmaster2_p & v8455ab | !hmaster2_p & v373aa3d;
assign v3a6f20c = hmaster1_p & v375e8d9 | !hmaster1_p & v37242b9;
assign v3a70c2c = hmaster2_p & v377fada | !hmaster2_p & v3a616ad;
assign v3a6f4c3 = hgrant4_p & c51aa0 | !hgrant4_p & v3a6becb;
assign v3739514 = hmaster2_p & v3a66aa4 | !hmaster2_p & v37738fc;
assign v3775b81 = locked_p & aca3c3 | !locked_p & v8455ab;
assign v95151c = hlock6 & v3a6ec52 | !hlock6 & v3a71078;
assign v3726a2b = hmaster1_p & v3a5a45e | !hmaster1_p & v3a62a6d;
assign v375640f = hbusreq6 & v37482f8 | !hbusreq6 & !v3a6fe6a;
assign v3739dfa = hmaster1_p & v2925d03 | !hmaster1_p & v3a6fa7c;
assign v3a6f6b6 = hgrant2_p & v37603a3 | !hgrant2_p & v3a71335;
assign v373c480 = hgrant3_p & v3a6c5ee | !hgrant3_p & bdda12;
assign v3a63690 = hbusreq6_p & v3730bf5 | !hbusreq6_p & v3776f7f;
assign v374838d = hmaster2_p & v376b4e5 | !hmaster2_p & v3730a3d;
assign v3762230 = hbusreq7 & v374705f | !hbusreq7 & v3a7071f;
assign v3a6574d = hbusreq5_p & v3775508 | !hbusreq5_p & v37620b4;
assign v3778a82 = hlock8_p & v8455e7 | !hlock8_p & !v8455ab;
assign v3a6ead6 = hbusreq4 & v3a70d04 | !hbusreq4 & v3a635ea;
assign v3746061 = hmaster0_p & v3a606b7 | !hmaster0_p & v3a6f379;
assign v3767437 = hlock0_p & v3a6a939 | !hlock0_p & !v8455ab;
assign v376c26e = hbusreq0 & v3a6b92c | !hbusreq0 & v377763c;
assign v3a621cb = hbusreq6_p & v3a59ee0 | !hbusreq6_p & v8455ab;
assign v3a67e79 = hgrant6_p & v3a645ca | !hgrant6_p & v3a70a43;
assign v37350f0 = hmaster2_p & v8455ab | !hmaster2_p & v3758d56;
assign v31461d5 = decide_p & v3a6b475 | !decide_p & v3a57b11;
assign v376c99e = hbusreq4_p & v3a66ea9 | !hbusreq4_p & v3a6f374;
assign v373aaf0 = hbusreq8 & v37505e1 | !hbusreq8 & v37545b7;
assign v37313e5 = hbusreq0 & v3729864 | !hbusreq0 & v3a6211e;
assign v3725ef7 = hgrant1_p & v337947a | !hgrant1_p & v3743690;
assign v37490ae = hbusreq5_p & v377bdec | !hbusreq5_p & v3733b46;
assign v3a6f6f0 = hbusreq8_p & v3a643ef | !hbusreq8_p & v38071c7;
assign v376bc6b = hbusreq5 & v39a53eb | !hbusreq5 & v8455ab;
assign v23fe101 = hlock6 & v375b7e1 | !hlock6 & v3a5dcfc;
assign v3a6fb83 = hlock0 & v3a635ea | !hlock0 & v3738937;
assign v374448e = hgrant4_p & v3735cb3 | !hgrant4_p & v3a5ca44;
assign v3a6f3d7 = jx3_p & v3724bbf | !jx3_p & v373bafb;
assign v373c627 = hbusreq1_p & v3768e48 | !hbusreq1_p & !v8455ab;
assign v3a702d9 = hmaster2_p & v374c5b2 | !hmaster2_p & v3a6ac60;
assign v3764979 = hbusreq3 & d44200 | !hbusreq3 & v8455ab;
assign v3a6dcf0 = hbusreq6 & v37482f8 | !hbusreq6 & !v3a703df;
assign v37418f3 = hbusreq8_p & v3a6aa9e | !hbusreq8_p & v3a5a9b3;
assign v3762f98 = hbusreq6_p & v37535e7 | !hbusreq6_p & v3a5ee12;
assign v3a5bb4f = hgrant6_p & v375564e | !hgrant6_p & v37548e6;
assign v37382ee = hlock7_p & v3740f78 | !hlock7_p & !v3a5a06e;
assign v3769e46 = hbusreq8_p & v3771502 | !hbusreq8_p & v376e663;
assign v3a6b17e = hmaster0_p & v376a91d | !hmaster0_p & v376ebc6;
assign v3a5fae3 = hgrant6_p & v3a6e31f | !hgrant6_p & v377815b;
assign v37462ae = hmaster0_p & v375bacc | !hmaster0_p & v3729173;
assign v37748b2 = hbusreq4 & v376c863 | !hbusreq4 & v8455ab;
assign v3762145 = hbusreq5_p & v373d5df | !hbusreq5_p & v374f52f;
assign v377b4fa = jx3_p & v3763b09 | !jx3_p & v3a708cd;
assign v376d48b = hmaster0_p & v3a5ab05 | !hmaster0_p & v8455ab;
assign v37265f2 = hmaster0_p & v3a66778 | !hmaster0_p & !v3728739;
assign v37241fd = hbusreq1_p & v3a63057 | !hbusreq1_p & v8455ab;
assign v377c5f4 = hmaster2_p & v3a6f240 | !hmaster2_p & v3a71631;
assign v376096f = hbusreq6 & v3a5b68a | !hbusreq6 & !v8455ab;
assign v3743e4a = hmaster1_p & a568f8 | !hmaster1_p & v3778fab;
assign v3766924 = hbusreq6_p & v377c07a | !hbusreq6_p & v374ec91;
assign v372be9b = hbusreq0_p & v3722e5c | !hbusreq0_p & v35772a6;
assign v3a70bc0 = hmaster1_p & v37596de | !hmaster1_p & v3724798;
assign v375a311 = hbusreq5_p & v3a5f2bd | !hbusreq5_p & v3a678de;
assign v3746806 = hbusreq6_p & v8455ab | !hbusreq6_p & v374fb58;
assign v3a55d78 = hbusreq5_p & v8d2bbf | !hbusreq5_p & !v3a68bdb;
assign v3774e5a = hbusreq5 & v374980f | !hbusreq5 & v3776cb6;
assign v37499a4 = hbusreq7_p & v374e8c3 | !hbusreq7_p & v3a70498;
assign v377c5de = hmaster2_p & v3a62caa | !hmaster2_p & v373bd76;
assign v37c048c = hgrant4_p & v375cc1b | !hgrant4_p & v3a5e55e;
assign v3a6d5b3 = hbusreq1 & v3a5ef54 | !hbusreq1 & v3a635ea;
assign v3754b79 = hbusreq4 & v375a938 | !hbusreq4 & !v3a70759;
assign v372316a = hbusreq5 & v373da33 | !hbusreq5 & v8455ab;
assign v375f852 = hbusreq5_p & v3a67d66 | !hbusreq5_p & v3a6f97b;
assign v3a6f58f = hlock8 & v37281be | !hlock8 & v3a704fb;
assign v3768eac = hbusreq4 & v3a7001d | !hbusreq4 & v3a5741c;
assign v3735ae4 = hbusreq8 & v373f1d4 | !hbusreq8 & v3755cc3;
assign v3a66476 = hgrant0_p & v3745b32 | !hgrant0_p & v23fe03a;
assign v3a69ef8 = hbusreq5 & v3a62cb7 | !hbusreq5 & v3728738;
assign v3a5fa4c = hlock5 & v3775526 | !hlock5 & v3724023;
assign v3725325 = hmaster1_p & v374db8d | !hmaster1_p & v3722b6c;
assign v3779c5d = hmaster1_p & v3806f0b | !hmaster1_p & v3a6f8c7;
assign v374e345 = hbusreq0 & v37451ad | !hbusreq0 & v3770c96;
assign v3257329 = hgrant2_p & v3730e2a | !hgrant2_p & v373c387;
assign v3a6f2f5 = hmaster2_p & v3a6fd81 | !hmaster2_p & v376d374;
assign v3740161 = hgrant4_p & v8455ab | !hgrant4_p & v3779070;
assign v3760f64 = hbusreq6_p & v8455bb | !hbusreq6_p & v3a65da7;
assign v377c0d5 = hlock5_p & v375415d | !hlock5_p & v3a69547;
assign v3773d82 = hgrant2_p & v374f307 | !hgrant2_p & v374ad1e;
assign v37292df = hgrant6_p & v3a6f312 | !hgrant6_p & v3754d8a;
assign v3758c64 = hlock1_p & v3a637dd | !hlock1_p & !v8455ab;
assign v3a635b9 = hmaster1_p & v3a61e95 | !hmaster1_p & v372661f;
assign v3a56570 = hlock7 & v3734279 | !hlock7 & v377aaa9;
assign v37541c6 = hmaster0_p & v3a59aa1 | !hmaster0_p & v376305d;
assign v374d153 = hbusreq0 & v372ab46 | !hbusreq0 & v373e814;
assign v3760073 = hlock3_p & v3a70020 | !hlock3_p & v2acaf74;
assign v3a5c511 = hlock5_p & v3770f96 | !hlock5_p & v376142a;
assign v375fbf2 = hbusreq4_p & v3a70209 | !hbusreq4_p & v3730ba6;
assign v3a666bb = hmaster0_p & v3a6c4e4 | !hmaster0_p & v373e484;
assign v3a70e73 = hbusreq7_p & v376ce17 | !hbusreq7_p & v376cd0a;
assign v3a6fc6a = hlock6 & v374668c | !hlock6 & v372dd89;
assign v3a615f5 = hbusreq8 & v374dabc | !hbusreq8 & v3a671f2;
assign v374b4d6 = hbusreq1_p & v8455eb | !hbusreq1_p & !v375bb3a;
assign v3a6b8aa = hbusreq0 & v3730755 | !hbusreq0 & v8455ab;
assign v373f503 = hlock1_p & v3a70a24 | !hlock1_p & !v8455ab;
assign v3a5d6aa = hmaster2_p & v3766b95 | !hmaster2_p & v3775688;
assign v372450e = hmaster1_p & v377fbd5 | !hmaster1_p & v377f264;
assign v376ebdd = hlock1_p & v3736a37 | !hlock1_p & !v8455ab;
assign v3752977 = hmaster0_p & v3727d7e | !hmaster0_p & v37243fe;
assign v3a67629 = hbusreq2 & v37457fb | !hbusreq2 & v8455e7;
assign v373ad68 = hgrant4_p & v3a62d48 | !hgrant4_p & v373d5dc;
assign v374d59a = hbusreq3 & v3a71452 | !hbusreq3 & v37416b5;
assign v3a70a03 = hlock4 & v374c61d | !hlock4 & v375d1ae;
assign v3a71503 = hbusreq0 & v8455b0 | !hbusreq0 & v3a59461;
assign v3a5be15 = hgrant4_p & v3734a92 | !hgrant4_p & v374ab4f;
assign v373d4f7 = hbusreq7_p & v373d09a | !hbusreq7_p & !v377516c;
assign v3a70974 = hbusreq2_p & v375d774 | !hbusreq2_p & v8455ab;
assign v3a6639e = hmaster1_p & v9243ac | !hmaster1_p & v37558f2;
assign v3777d39 = hbusreq0 & v3727d00 | !hbusreq0 & v3a67e53;
assign v3743da0 = hlock0_p & v3806db7 | !hlock0_p & v377378e;
assign v373628e = hbusreq6_p & v3a614cb | !hbusreq6_p & v373b288;
assign v3a69674 = hmaster0_p & v3763175 | !hmaster0_p & v3a6fdbf;
assign v3a5b0f5 = hlock8_p & v374215e | !hlock8_p & v374c6de;
assign v373e789 = hbusreq6 & v39eb3bd | !hbusreq6 & v3731004;
assign v38076b3 = hmaster3_p & v37599b8 | !hmaster3_p & v37511f6;
assign v3a637dc = stateA1_p & v8455e1 | !stateA1_p & v372fc17;
assign v3a5e544 = hbusreq3_p & v377fb9d | !hbusreq3_p & v8455ab;
assign a13040 = hgrant5_p & v3a6ffc3 | !hgrant5_p & v3a7135e;
assign v374d6ff = hbusreq5_p & v3a70ae8 | !hbusreq5_p & v3a6ecdd;
assign v377ed8e = hlock6_p & v8455e1 | !hlock6_p & !v8455ab;
assign v377ce66 = hbusreq1_p & v37570b7 | !hbusreq1_p & !v8455ab;
assign v374113d = hbusreq6 & v3a5d3af | !hbusreq6 & v3742f28;
assign aca3c3 = hmastlock_p & v3a6fa4f | !hmastlock_p & v8455ab;
assign v3a687e0 = hbusreq0 & v372f759 | !hbusreq0 & v376ab01;
assign v375da10 = hbusreq1_p & v3747302 | !hbusreq1_p & v37496fa;
assign v3777498 = hbusreq5_p & v37514e4 | !hbusreq5_p & v372e4ac;
assign v372e99c = hmaster1_p & v3a60332 | !hmaster1_p & v3776923;
assign v3733a0e = hbusreq7 & bb3b0a | !hbusreq7 & v3a29814;
assign v3752ee5 = hmaster2_p & v3a5e24e | !hmaster2_p & v39a537f;
assign v377d27a = hbusreq0 & v3779008 | !hbusreq0 & dbc26f;
assign v3750da4 = jx0_p & v3766246 | !jx0_p & v37573c5;
assign v373bb2f = hmaster1_p & v8455ab | !hmaster1_p & v375c9bc;
assign v3a54d84 = hlock2 & v3a6c8dc | !hlock2 & v3a64703;
assign v3a6f69c = jx1_p & v375c2e2 | !jx1_p & v8455ab;
assign v209310e = hbusreq2_p & v8455ab | !hbusreq2_p & !v3a637dd;
assign v373bf09 = hmaster0_p & v3772696 | !hmaster0_p & v3a71133;
assign v37727f9 = hmaster1_p & v35b774b | !hmaster1_p & v3a70620;
assign v380a1a6 = hbusreq2 & c61447 | !hbusreq2 & v3761ad0;
assign v3751981 = jx0_p & v3a6f834 | !jx0_p & !v3a594e8;
assign v3745b71 = hbusreq5 & v3a6aaed | !hbusreq5 & !v8455ab;
assign v2ff87db = decide_p & v23fd910 | !decide_p & v377a6c4;
assign v373d434 = hgrant0_p & v8455ab | !hgrant0_p & !v3a71287;
assign v23fe329 = hgrant6_p & v3748194 | !hgrant6_p & !v3a54c12;
assign v3749a12 = busreq_p & v3749d1d | !busreq_p & !v8455fd;
assign v23fd910 = hready_p & v2ff9353 | !hready_p & v3726c99;
assign v3a6744e = hmaster2_p & v8455ab | !hmaster2_p & v3a704cc;
assign v3a70bfb = hgrant5_p & v3a6fc98 | !hgrant5_p & v3748ab9;
assign v37656f7 = hbusreq5 & v377bd77 | !hbusreq5 & v8455ab;
assign v374f52a = hmaster0_p & v3a58cfc | !hmaster0_p & v3a5b545;
assign v376d256 = hbusreq2 & v3a7104b | !hbusreq2 & !v8455ab;
assign v375a02d = hbusreq3_p & v3730cda | !hbusreq3_p & v37244e7;
assign v37592d6 = hbusreq2 & v377ba55 | !hbusreq2 & v8455ab;
assign v373ce86 = hgrant4_p & v8455c2 | !hgrant4_p & v374df50;
assign v3a656b6 = hbusreq0 & v38097db | !hbusreq0 & v3725ec4;
assign v3a713bb = hmaster1_p & v3a5e24e | !hmaster1_p & v9b81ab;
assign v375b878 = hgrant6_p & v37379fc | !hgrant6_p & v3748fba;
assign v3a6d098 = hmaster2_p & v37261b3 | !hmaster2_p & v8455ab;
assign v37310be = hgrant6_p & v3a645b0 | !hgrant6_p & v3a6a1fd;
assign v3a58615 = hmaster2_p & v376641b | !hmaster2_p & !v3a71453;
assign v373d32e = hbusreq5_p & v376ce6f | !hbusreq5_p & v3a6f809;
assign v3a71354 = hgrant2_p & v3a5b5d3 | !hgrant2_p & !v373f4a5;
assign v376b8f1 = hlock4_p & v8455ab | !hlock4_p & v39a5265;
assign v3a6dbf0 = hgrant6_p & v37293f6 | !hgrant6_p & v3a6ba77;
assign v3741ef3 = hgrant6_p & v8455ab | !hgrant6_p & v37532a6;
assign v374f31d = hmaster2_p & v3747042 | !hmaster2_p & v3a5a01b;
assign v3771d56 = hmaster1_p & v3a56cfd | !hmaster1_p & v372e749;
assign v3729d1a = hbusreq3_p & v39a537f | !hbusreq3_p & !v3a63bbc;
assign v377d596 = hmaster2_p & v3736847 | !hmaster2_p & v3a627cc;
assign v8d9a96 = hbusreq6 & v376f56d | !hbusreq6 & !v8455ab;
assign v375210d = hmaster0_p & v376aa57 | !hmaster0_p & v3757c5c;
assign v372810e = hbusreq4 & v3a6ec2a | !hbusreq4 & v8455ab;
assign v375f15c = hmaster2_p & v374e28f | !hmaster2_p & !v37369b2;
assign v3a5d065 = hbusreq8_p & v3a70578 | !hbusreq8_p & v3758bcd;
assign v94ce87 = hbusreq3 & v37482f8 | !hbusreq3 & !v372b24d;
assign v3734abe = hbusreq6 & v37564e4 | !hbusreq6 & !v8455bd;
assign a7e544 = jx0_p & v375ab8e | !jx0_p & v3a62f8e;
assign v3a57f41 = hlock0_p & v3768ac7 | !hlock0_p & v3744710;
assign v3725626 = hmaster1_p & v3a628cf | !hmaster1_p & v3a6eb7d;
assign v3a54e0c = hgrant5_p & v8455ab | !hgrant5_p & v3752ebb;
assign v374612b = hlock4_p & v20d166d | !hlock4_p & v8455ab;
assign v3a571fa = hmaster2_p & v372348c | !hmaster2_p & v3a6efea;
assign v372fa0f = hbusreq6 & v3763175 | !hbusreq6 & v8455ab;
assign v377f46d = hbusreq6_p & v3a6324b | !hbusreq6_p & v8455bb;
assign v376f979 = hmaster0_p & v377851b | !hmaster0_p & v373e267;
assign v372e4e1 = hmaster0_p & v8455ab | !hmaster0_p & v37656e5;
assign v3779e70 = stateG10_1_p & v2aca977 | !stateG10_1_p & v3748900;
assign v3a70d04 = hlock6 & ce69d1 | !hlock6 & v37495dc;
assign v3a6f529 = hmaster2_p & v3a63777 | !hmaster2_p & v377b946;
assign v377104a = hbusreq5_p & v3723d73 | !hbusreq5_p & !v8455ab;
assign v375fcb7 = hbusreq4 & v373c4c2 | !hbusreq4 & !v8455bd;
assign v3a6c4bb = hbusreq7 & b0015f | !hbusreq7 & v377e30e;
assign v3741d24 = hmaster0_p & v3741d52 | !hmaster0_p & v3a70f9c;
assign v3a5b25f = hmaster0_p & v3745714 | !hmaster0_p & v3a61c70;
assign v3a5f626 = hgrant5_p & v8455ab | !hgrant5_p & v375e074;
assign v3746559 = jx1_p & v377c8c8 | !jx1_p & v377aed3;
assign v377b951 = hmaster1_p & v3768995 | !hmaster1_p & v3a5a5c8;
assign v3772229 = hmaster2_p & v3a70ecb | !hmaster2_p & v8455ab;
assign v3755d8e = hlock7_p & v37716b0 | !hlock7_p & v3a7087f;
assign v377ab46 = hlock6 & v373b6c0 | !hlock6 & v3a6f9b9;
assign v372d1f0 = hmaster0_p & v3768495 | !hmaster0_p & v23fdebb;
assign a1bc5b = hmaster2_p & v3a6a8c0 | !hmaster2_p & v3769740;
assign v37719a9 = hmaster0_p & v375b5ce | !hmaster0_p & v3736ded;
assign v37527dc = hmaster2_p & v37705c0 | !hmaster2_p & v376fad7;
assign v377eada = hmaster0_p & v373e625 | !hmaster0_p & v375ec23;
assign v3a70761 = hmaster2_p & v3a635ea | !hmaster2_p & v377ca49;
assign v3a56b7c = hmaster2_p & v3a6f91e | !hmaster2_p & v372a071;
assign v37372dd = hlock6 & v3762c73 | !hlock6 & b4f73f;
assign v3a5d7f7 = hgrant5_p & v373471a | !hgrant5_p & !v8455ab;
assign v3a6eb09 = hmaster1_p & v3a58cfc | !hmaster1_p & v3745a3b;
assign v37584c6 = hbusreq0 & v377ac4c | !hbusreq0 & b3f461;
assign v3767b2e = hbusreq7 & v375dd92 | !hbusreq7 & v3776f7d;
assign v3773f26 = hmaster2_p & dc5fea | !hmaster2_p & v3775e81;
assign v373dcd2 = hlock3 & v37254c0 | !hlock3 & v3734c26;
assign v397d860 = decide_p & v37666b4 | !decide_p & v376a25e;
assign v375e346 = hmaster2_p & v3777790 | !hmaster2_p & !v376b4ad;
assign v3a6f9c7 = hlock4 & v3808dd8 | !hlock4 & v3a68f98;
assign v3a7039c = jx1_p & v377d414 | !jx1_p & v377f7dd;
assign v377cf4f = hmaster0_p & v377b24b | !hmaster0_p & v8bc1c0;
assign v3a6d0a1 = hgrant2_p & v3a55b61 | !hgrant2_p & v3a65d4e;
assign v3a5f0f0 = jx0_p & v376fe68 | !jx0_p & v3730f97;
assign v3770fb7 = hmaster2_p & v37261b3 | !hmaster2_p & v8f695f;
assign v377f4e5 = hgrant6_p & v376e0fa | !hgrant6_p & v3768ec4;
assign v376d766 = hmaster0_p & v8455e7 | !hmaster0_p & v375ace5;
assign v3a70d57 = hgrant2_p & v377182c | !hgrant2_p & v374f485;
assign v3a574d6 = hbusreq5 & v375a5e3 | !hbusreq5 & v8455ab;
assign v3a6fae2 = hlock0_p & v37682c6 | !hlock0_p & v375589b;
assign v373ea50 = jx0_p & v37386d3 | !jx0_p & v8455ab;
assign v37327fe = hmaster0_p & v3a693b7 | !hmaster0_p & v3740e4c;
assign v372cb36 = hbusreq8 & v3a60223 | !hbusreq8 & v377386a;
assign v3a672c9 = hbusreq1_p & v376d45f | !hbusreq1_p & v3a5bf04;
assign v3a70242 = hmaster1_p & v372317f | !hmaster1_p & v3a6fb0e;
assign v37717ee = hlock5 & v3a5aefc | !hlock5 & v373f07d;
assign v3770a5a = hmaster0_p & v3764a6c | !hmaster0_p & v377cccb;
assign v377d945 = hmaster2_p & v8455ab | !hmaster2_p & v372e821;
assign v3746f37 = hgrant1_p & v3a65c29 | !hgrant1_p & v8455ab;
assign v373c342 = hgrant5_p & v3a6bd0f | !hgrant5_p & v375c4c7;
assign v375c05f = hbusreq4 & v373014d | !hbusreq4 & v8455bf;
assign v373b11b = hlock2 & v3740fe0 | !hlock2 & v376bb88;
assign v376a7ac = hmaster2_p & v376d9ad | !hmaster2_p & v374362e;
assign v37430db = hbusreq8_p & v372e611 | !hbusreq8_p & v37742f4;
assign v3a6ab5f = stateA1_p & v8455e1 | !stateA1_p & !v3757c6f;
assign v37435a8 = hbusreq0 & v3a54ba5 | !hbusreq0 & v373bfd9;
assign v3a6051a = hlock0_p & v37401f0 | !hlock0_p & v3a5df94;
assign v376e491 = hmastlock_p & v3a6affa | !hmastlock_p & !v8455ab;
assign v3736fdd = hgrant0_p & v8455ab | !hgrant0_p & v3a703cc;
assign v3743ef0 = hbusreq0 & v377dfec | !hbusreq0 & v8455ab;
assign v3770fff = hbusreq7 & v3a6fa70 | !hbusreq7 & v3a5f3f0;
assign v3740233 = hlock5_p & v3a7066b | !hlock5_p & v3748446;
assign v3a6ec01 = hgrant5_p & v3a6f5a4 | !hgrant5_p & v2092ac1;
assign v3740c5f = hmaster0_p & v3a635ea | !hmaster0_p & v3750ad1;
assign v3a5c842 = hgrant5_p & v3740ed1 | !hgrant5_p & v3a573bb;
assign v37372eb = hlock5 & v3754ba1 | !hlock5 & v375129f;
assign v3a6fc76 = hbusreq7_p & v3767c92 | !hbusreq7_p & v3a6242b;
assign v373f0c7 = hbusreq7_p & v3727b7f | !hbusreq7_p & v37470de;
assign v3753804 = hmaster0_p & v372ed5f | !hmaster0_p & v8455ab;
assign v3736b57 = hbusreq4 & v3750f8f | !hbusreq4 & v3748797;
assign v37347b2 = hbusreq5 & v372afe7 | !hbusreq5 & v375b0ad;
assign v3769a34 = hmaster0_p & v376111d | !hmaster0_p & v3736b1d;
assign v3a7146b = hbusreq0 & v3765dda | !hbusreq0 & v8455ab;
assign v3764462 = hbusreq6_p & v3775de3 | !hbusreq6_p & v3a5f315;
assign v377d607 = hbusreq7_p & v377ab40 | !hbusreq7_p & v3a7054d;
assign v3a6e123 = hbusreq4_p & v3a63805 | !hbusreq4_p & v8455b0;
assign v376dffd = hbusreq8 & v375e439 | !hbusreq8 & v37624e5;
assign v3a5d0b6 = hgrant3_p & v372f657 | !hgrant3_p & v3a6fff6;
assign v377d52e = hgrant3_p & v8455ab | !hgrant3_p & v3a70a34;
assign v3745529 = hlock4_p & v8455ab | !hlock4_p & v373fe5e;
assign v377538f = stateG10_1_p & v3a635ea | !stateG10_1_p & v373a8d6;
assign v3a69d78 = hmaster1_p & v3a6f9a1 | !hmaster1_p & !v35b77ab;
assign v3a58fe9 = hbusreq7_p & v3746d75 | !hbusreq7_p & v3a618ea;
assign aa5556 = hbusreq6 & v3a5600a | !hbusreq6 & v8455ab;
assign v376293b = hbusreq8 & v372809b | !hbusreq8 & v3723e62;
assign v3a713cd = hmaster0_p & v8455ab | !hmaster0_p & v35ba1c6;
assign v376641b = hbusreq2_p & v3a6fbef | !hbusreq2_p & !v8455ab;
assign v3a705ee = hmaster1_p & v373e01f | !hmaster1_p & v8455ab;
assign v3a6f051 = hlock5_p & v373bbd0 | !hlock5_p & v37404c5;
assign v3a6fcfa = hmaster0_p & v374c5e2 | !hmaster0_p & v3a7031b;
assign v375a7d3 = hlock4 & v3a63da7 | !hlock4 & v3777eed;
assign v375b42e = hbusreq4_p & v3747302 | !hbusreq4_p & v3a7063e;
assign v374fb51 = hgrant6_p & v8455ca | !hgrant6_p & v373fee1;
assign v3a6fe61 = hbusreq7 & v3a702e3 | !hbusreq7 & v3759284;
assign v374f547 = hbusreq6_p & v377b3cf | !hbusreq6_p & !v8455ab;
assign v3a70466 = hlock2 & v2889703 | !hlock2 & v3774c4d;
assign v374faa9 = hgrant2_p & v3747302 | !hgrant2_p & v37765e1;
assign v377ed2d = hbusreq5_p & v37556c1 | !hbusreq5_p & v3a63966;
assign v3a6f9cd = hmaster2_p & v3764881 | !hmaster2_p & !v374a2cc;
assign v3748cb7 = hmaster1_p & v8455ab | !hmaster1_p & v3a6ceb0;
assign v3a57cd0 = hbusreq6_p & v3a594a5 | !hbusreq6_p & v3a704ee;
assign v374b40e = hmaster1_p & v8455e7 | !hmaster1_p & v3a55aa3;
assign v376b540 = hmaster2_p & v37429e5 | !hmaster2_p & v3a5bb64;
assign v377f09a = hbusreq6_p & v3a6fce6 | !hbusreq6_p & !v8455ab;
assign v374d13c = hbusreq2 & v3a55e7f | !hbusreq2 & v3a713e3;
assign v3a64e2a = hlock0 & v3a635ea | !hlock0 & v376ffbf;
assign v3a7029b = hbusreq3_p & v380704f | !hbusreq3_p & v3743b9e;
assign v3739acd = hmaster0_p & v3a70463 | !hmaster0_p & !v3750088;
assign v374fcac = hbusreq8 & v3a7043d | !hbusreq8 & !v8455ab;
assign v375e320 = hmaster1_p & v3738ca1 | !hmaster1_p & v3a70f68;
assign v23fde66 = hbusreq7_p & v3750254 | !hbusreq7_p & v3a69bdc;
assign v37384cb = hmaster3_p & v3724579 | !hmaster3_p & v3a713e8;
assign v3a70a79 = hmaster2_p & v375a94a | !hmaster2_p & !v8455ab;
assign v3769090 = hmaster2_p & v374f5e0 | !hmaster2_p & v3a5e070;
assign v3763104 = hlock4_p & v377b774 | !hlock4_p & v8455bf;
assign v3a6fa49 = hgrant2_p & v8455ab | !hgrant2_p & !v3770919;
assign v3769323 = hmaster1_p & v376c7f9 | !hmaster1_p & v28896cd;
assign v3a68607 = hgrant6_p & v374a664 | !hgrant6_p & v37765fb;
assign v2acaeb7 = hgrant3_p & v376ace9 | !hgrant3_p & v376fa80;
assign v3774d2a = hbusreq8 & v3747429 | !hbusreq8 & v372e2eb;
assign v3a71124 = hbusreq7 & v3a6375b | !hbusreq7 & v3a5a807;
assign v3a66910 = hbusreq4_p & v3a6f59d | !hbusreq4_p & !v8455ab;
assign v3a5eaaf = hgrant4_p & v8455ab | !hgrant4_p & v374617d;
assign baccec = hbusreq6_p & v3a6fd5c | !hbusreq6_p & !v372df2a;
assign v3a709d5 = hbusreq7_p & v376d872 | !hbusreq7_p & v375ddaf;
assign v3a5d834 = hbusreq7_p & v3a70d4e | !hbusreq7_p & v3a5f47b;
assign v376a1d7 = hbusreq3_p & v3a5fa18 | !hbusreq3_p & v3a7145b;
assign v3a5acc7 = hmaster2_p & v8455ab | !hmaster2_p & !v3753ccf;
assign v3806a6f = hbusreq2 & v37645a8 | !hbusreq2 & v3a70b92;
assign v3a70b9e = hbusreq6_p & v3757ec8 | !hbusreq6_p & v37375bc;
assign v376139f = hmaster1_p & v375d387 | !hmaster1_p & v3779931;
assign v3a704cd = jx0_p & v2ff87d7 | !jx0_p & v373150d;
assign v374ebc5 = hbusreq0 & v374096a | !hbusreq0 & v8455ab;
assign v3a6eef6 = hbusreq0_p & v3a64ee3 | !hbusreq0_p & !v37583be;
assign v3773afc = hmaster1_p & v3749f94 | !hmaster1_p & v3773dc6;
assign v377542e = hbusreq2 & v3725c68 | !hbusreq2 & v3a635ea;
assign v3751e7c = hbusreq7 & v3809b0a | !hbusreq7 & v376ae9f;
assign v374ee76 = jx1_p & v3756d56 | !jx1_p & v3a701f0;
assign v372526e = hgrant3_p & v3a69c6f | !hgrant3_p & v3757f9b;
assign v3a6f343 = hbusreq2 & v3a70385 | !hbusreq2 & !v3378ef7;
assign v3a5ab33 = hbusreq0 & v3a571fd | !hbusreq0 & v3a70876;
assign v375cab0 = hbusreq2_p & v37273c2 | !hbusreq2_p & v375d161;
assign v3755d10 = hmaster1_p & v3a70b35 | !hmaster1_p & v376e441;
assign v3729ddd = hmaster0_p & v3a6fa97 | !hmaster0_p & !v372a450;
assign v376b65a = hmaster2_p & v374aec2 | !hmaster2_p & v3730986;
assign v3a6fcda = hbusreq0 & v376dba6 | !hbusreq0 & v3a6c717;
assign v3738d54 = hmaster3_p & v373b9e9 | !hmaster3_p & !v3a681f5;
assign v377ce7d = hgrant6_p & v375b7bd | !hgrant6_p & v3a71265;
assign v3a714fe = jx0_p & v3808ceb | !jx0_p & v372e9b1;
assign v376bd2c = hbusreq5_p & v3a5c945 | !hbusreq5_p & v3a57f59;
assign v3a70278 = hburst1 & v3a6ffa9 | !hburst1 & v37739c7;
assign v3778176 = hlock1_p & v8455ab | !hlock1_p & v39a5265;
assign v372976e = hgrant4_p & v8455ab | !hgrant4_p & v3756b8a;
assign v3a70d4a = hgrant8_p & v8455ab | !hgrant8_p & v37629db;
assign v3a58a1b = hlock4 & v376a3bb | !hlock4 & v3a63fc5;
assign v374472d = hbusreq5_p & v374b362 | !hbusreq5_p & v37518e7;
assign v3a714ac = hbusreq2_p & v3764a16 | !hbusreq2_p & v375bc5b;
assign v375ccc3 = hbusreq4 & v3a5b121 | !hbusreq4 & v8455bf;
assign v372c016 = hmaster1_p & v3736d47 | !hmaster1_p & v374de43;
assign v3779dae = hbusreq3_p & v375c7f8 | !hbusreq3_p & !c17897;
assign v3a5b01c = hmaster1_p & v3a57f59 | !hmaster1_p & v3a60836;
assign v3a705e1 = hlock1_p & v8455ab | !hlock1_p & !v376430b;
assign v3728b47 = hbusreq8_p & v3756343 | !hbusreq8_p & v8455ab;
assign v374cb90 = hgrant3_p & v3750d06 | !hgrant3_p & !v3a5a798;
assign v3a6cc9a = hmaster2_p & v3a5600a | !hmaster2_p & v3754c5e;
assign v3a6fac9 = hbusreq4_p & v37501e1 | !hbusreq4_p & v8455b3;
assign v372a0cb = hbusreq7 & v3a70f38 | !hbusreq7 & v3730f6f;
assign v373217b = stateG10_1_p & v372fc51 | !stateG10_1_p & v37393f0;
assign v374e43a = hbusreq4 & v3a61901 | !hbusreq4 & v372e83f;
assign v3752e8e = hlock0_p & v8455ab | !hlock0_p & v3a70b60;
assign v3a549f5 = jx1_p & v3763e6c | !jx1_p & v3a7132c;
assign v3a715b2 = hbusreq0 & v3a5b4be | !hbusreq0 & v8455ab;
assign v3724710 = stateG10_1_p & v8455ab | !stateG10_1_p & v374ed4b;
assign c47a78 = hbusreq8 & v373f3ac | !hbusreq8 & v374312f;
assign v376ed30 = hbusreq6_p & v376803b | !hbusreq6_p & v374e26d;
assign v3a6fc30 = hbusreq2_p & v3a6f99d | !hbusreq2_p & !v8455ab;
assign v3727a12 = hbusreq8 & v372a298 | !hbusreq8 & v375bfc4;
assign v3770c2a = hmaster1_p & v3a6a872 | !hmaster1_p & v37331d1;
assign v3a5ddef = hmaster1_p & v38063ce | !hmaster1_p & v37474e1;
assign v37390ff = hbusreq3 & v37482f8 | !hbusreq3 & !v3a7104b;
assign v3a6f7fb = hbusreq2_p & v3a70cd3 | !hbusreq2_p & v3763acf;
assign v37374bc = jx0_p & v3a6a81f | !jx0_p & v3a64a7b;
assign v3a6c793 = hbusreq5_p & v3a70d97 | !hbusreq5_p & v8455b0;
assign v37435b7 = hmaster1_p & v3762f27 | !hmaster1_p & v3759c8c;
assign v3a7123c = hgrant8_p & v8455d2 | !hgrant8_p & v372b69c;
assign v373fd50 = hlock0 & v3735525 | !hlock0 & v37729db;
assign v372e268 = hmaster1_p & v3a6f563 | !hmaster1_p & v374554d;
assign v3a6f758 = hbusreq5 & v374f077 | !hbusreq5 & v37583f0;
assign v3a6b129 = hbusreq2_p & v3725252 | !hbusreq2_p & v3a71379;
assign v372ff0a = hgrant4_p & v3a70aeb | !hgrant4_p & v3a70b7c;
assign v3764539 = hmaster0_p & v3741b59 | !hmaster0_p & v3737f8d;
assign v3808952 = hlock4 & v3a71037 | !hlock4 & v3a5715d;
assign v374d138 = hmaster2_p & v3769093 | !hmaster2_p & v37325a2;
assign v3a5bc4f = hmaster1_p & v8455ab | !hmaster1_p & v3a6fbc7;
assign v3724696 = hbusreq5 & v3a58c07 | !hbusreq5 & v37476b8;
assign v3a6fb7f = hmaster0_p & v3a635ea | !hmaster0_p & v372cea0;
assign v3726d1f = hgrant6_p & v3747302 | !hgrant6_p & v374faa9;
assign v3a6e33a = hlock8 & v3746312 | !hlock8 & v3749544;
assign v3a57c78 = hbusreq5 & v3774a7d | !hbusreq5 & v8455ab;
assign v3a5af68 = hmaster1_p & v373014d | !hmaster1_p & v37307a7;
assign v376a1dd = hgrant4_p & v37604e9 | !hgrant4_p & v3a680e3;
assign v3a6fbdb = hbusreq5 & v3740681 | !hbusreq5 & v3767e7f;
assign v37496d3 = hlock6_p & v3a5f0b2 | !hlock6_p & v3a6f8f5;
assign v375355a = hmaster2_p & v3a6f4f8 | !hmaster2_p & v3a5b037;
assign v373e4c0 = hlock0 & v374e768 | !hlock0 & v39eb452;
assign v376e7a5 = hmaster2_p & v39a5265 | !hmaster2_p & v3a714aa;
assign v377efdc = hbusreq3_p & v377caa3 | !hbusreq3_p & !v8455ab;
assign v3731320 = hbusreq4_p & v3754fc8 | !hbusreq4_p & v375af57;
assign v3736da4 = hgrant3_p & v376ea4a | !hgrant3_p & v28896c8;
assign v37325cf = hbusreq6_p & v374eac6 | !hbusreq6_p & v3725717;
assign v3a6f629 = hbusreq5_p & v375d577 | !hbusreq5_p & !v3a70cf6;
assign v37343bd = hbusreq8 & v3737298 | !hbusreq8 & v8455ab;
assign v3a700ff = hbusreq7_p & v37249fe | !hbusreq7_p & v3a5d646;
assign v377e29a = hlock6 & v3774aa2 | !hlock6 & v3738d0b;
assign v372713b = hmaster0_p & v3a635ea | !hmaster0_p & v376a480;
assign v375e00a = hbusreq6 & v3763a20 | !hbusreq6 & v8455bf;
assign v3a60b88 = hgrant4_p & v9ed516 | !hgrant4_p & v3a7005f;
assign v3a5f3a1 = hmaster2_p & v37731ce | !hmaster2_p & v37745c3;
assign v3a57b00 = hgrant5_p & v8455ab | !hgrant5_p & !v37348f5;
assign v3a703d7 = hmaster0_p & v38073bb | !hmaster0_p & v376132a;
assign v3779f67 = hlock6_p & v8455ab | !hlock6_p & v375d5ac;
assign v3723e5d = hlock4 & v3745b0f | !hlock4 & v3775a92;
assign v3a55078 = jx0_p & v376d3a6 | !jx0_p & v37630e2;
assign v375ac50 = hgrant4_p & v3a6fe35 | !hgrant4_p & v3a702d3;
assign v3725d73 = hbusreq6 & v374e056 | !hbusreq6 & v8455ab;
assign v37306bb = hbusreq1 & v3a63621 | !hbusreq1 & v3a635ea;
assign v3741d83 = hmaster0_p & v20d166d | !hmaster0_p & v3a70c98;
assign v373deb5 = stateA1_p & v8455e1 | !stateA1_p & v8455ab;
assign v3a6f118 = hbusreq8 & v3732632 | !hbusreq8 & v3a707e5;
assign v372e474 = hbusreq0_p & v3a635ea | !hbusreq0_p & v3a6edab;
assign v373d551 = hgrant2_p & v3a59bb4 | !hgrant2_p & v377abb1;
assign v3a675b9 = hmaster1_p & v3733cfb | !hmaster1_p & v377b6ce;
assign v376ecc8 = hbusreq6_p & v3764978 | !hbusreq6_p & v8455ab;
assign v3769d3d = jx1_p & v8455ab | !jx1_p & v3767183;
assign v373f0e6 = hbusreq0 & v3a6f8fd | !hbusreq0 & v3726381;
assign v372396a = hgrant3_p & v360d1cb | !hgrant3_p & v372c577;
assign v3745e1f = hgrant6_p & v3a6ba6a | !hgrant6_p & v373e09c;
assign v3a54484 = jx0_p & v3747b4c | !jx0_p & v373b647;
assign v3765f99 = hlock5_p & v3a609da | !hlock5_p & v8455cb;
assign v3a67f49 = hmaster1_p & v3a65a0f | !hmaster1_p & v3a5a807;
assign v372b627 = hbusreq8 & dc571e | !hbusreq8 & v8455ab;
assign v3a5f853 = hbusreq7_p & v3a71161 | !hbusreq7_p & v3750c57;
assign v37355db = hgrant0_p & v8455ab | !hgrant0_p & v3726bb8;
assign v3762cff = hlock0_p & v372c3df | !hlock0_p & v3a5996e;
assign v3749544 = hlock7 & v3740c73 | !hlock7 & v3770e77;
assign v3a711e6 = hmaster0_p & v380760a | !hmaster0_p & !v3762e85;
assign d4d3bb = hmaster2_p & v3730ddd | !hmaster2_p & v3a71228;
assign v3731b90 = hmaster2_p & v3a5979b | !hmaster2_p & v3760700;
assign v3735936 = hlock5_p & v3a5d527 | !hlock5_p & v8455ab;
assign v3734fa5 = hbusreq5 & v8455ab | !hbusreq5 & v3a6fd4a;
assign v3a61246 = hbusreq5 & v3807183 | !hbusreq5 & !v3a6c5e5;
assign v373da95 = hgrant4_p & v8455ab | !hgrant4_p & v3779f1c;
assign v3763793 = hbusreq1 & v37583be | !hbusreq1 & !v8455ab;
assign v3a6f428 = hready & v3740415 | !hready & v38072fd;
assign v3a5b71a = hlock0_p & v8455e7 | !hlock0_p & v8455ab;
assign v3762034 = hbusreq4_p & v3742e30 | !hbusreq4_p & !v8455ab;
assign v3722a7e = hgrant6_p & v377f09a | !hgrant6_p & v3a5e363;
assign v373d5ac = hbusreq5_p & v3a57486 | !hbusreq5_p & v3776da7;
assign v373e2b7 = hgrant5_p & v3741e09 | !hgrant5_p & v3742d2a;
assign v3a667cf = hmaster2_p & v3753c73 | !hmaster2_p & v1e37523;
assign v373f1aa = hgrant5_p & v8455ab | !hgrant5_p & !v3a6f64d;
assign v373d9a2 = hmaster2_p & v377a3bd | !hmaster2_p & v3a56b60;
assign v37503ce = hgrant5_p & v373fe39 | !hgrant5_p & v37717ed;
assign v372d732 = hmaster1_p & v372ca6e | !hmaster1_p & v374610d;
assign v37530e8 = hmaster1_p & v3a6eb67 | !hmaster1_p & v37300e3;
assign v376c5f3 = hbusreq4_p & v3a70a7d | !hbusreq4_p & v37551ec;
assign v3a6f2d8 = hmaster0_p & v3a635ea | !hmaster0_p & v23fd9f9;
assign v377e172 = hgrant6_p & v377618a | !hgrant6_p & v3778151;
assign v3759b9a = hgrant0_p & v3a655c2 | !hgrant0_p & v37376c8;
assign v376af8e = hlock7 & a0a219 | !hlock7 & v37297f9;
assign v3a5df66 = hlock5 & v3a713d5 | !hlock5 & v373e219;
assign v3732bb6 = hmaster0_p & v376d1b3 | !hmaster0_p & v37411c6;
assign v3730451 = hbusreq4 & v3740a38 | !hbusreq4 & v3a6fdef;
assign v37706dd = hbusreq4_p & v3a711e7 | !hbusreq4_p & v3730d6a;
assign v37776f0 = hlock5 & v3a6d792 | !hlock5 & v3a642c5;
assign v3730c0b = hmaster1_p & v1e379c4 | !hmaster1_p & v375523e;
assign v377bbbb = hbusreq2 & v3778251 | !hbusreq2 & v3748797;
assign v377222a = hgrant6_p & v3a6f3a1 | !hgrant6_p & v37341b2;
assign v377638d = hlock5 & v375aa18 | !hlock5 & v374518e;
assign v3754227 = hbusreq3_p & v375ea58 | !hbusreq3_p & !v8455ab;
assign b6ae10 = hbusreq4_p & v375b878 | !hbusreq4_p & v2acafdf;
assign v3a700e9 = hmaster0_p & v3a70987 | !hmaster0_p & v3a62079;
assign v3a711c1 = hbusreq6_p & v3776e85 | !hbusreq6_p & v3736439;
assign v1e37bf6 = hgrant6_p & v8455ab | !hgrant6_p & v2092baa;
assign v1e37ca4 = hbusreq0 & v3a6243f | !hbusreq0 & bf29af;
assign v3a6f809 = hbusreq5 & v3a7045d | !hbusreq5 & v375d152;
assign v3a62a53 = hgrant2_p & v3a710e1 | !hgrant2_p & v3a56bd5;
assign v375c7c4 = hbusreq7_p & v3a6799a | !hbusreq7_p & !v3742360;
assign v3a70000 = hbusreq5 & v3728ced | !hbusreq5 & v3a68787;
assign v3a62015 = hgrant4_p & v8455ab | !hgrant4_p & v3758b89;
assign v375e06b = hmaster0_p & v376501e | !hmaster0_p & v376196f;
assign v3a7036a = hgrant3_p & v37c1a6f | !hgrant3_p & v376bc4b;
assign v375329c = hmaster0_p & v3a71135 | !hmaster0_p & v3727e58;
assign v3755e23 = hbusreq6_p & v3a56582 | !hbusreq6_p & !v3a6f897;
assign v376596c = hbusreq8_p & v3a70d59 | !hbusreq8_p & v8455ab;
assign v3727662 = hgrant6_p & v8455ab | !hgrant6_p & v3a6f767;
assign v374a637 = hbusreq3_p & v3a7162d | !hbusreq3_p & v3778528;
assign v3747787 = hgrant4_p & v3a70bd6 | !hgrant4_p & v373cf60;
assign v3727bd4 = hbusreq5_p & v3769edd | !hbusreq5_p & v375671a;
assign v3764c4c = hlock2_p & v8455ab | !hlock2_p & v3771ce2;
assign v3a6f782 = hbusreq2 & v3a6ab5f | !hbusreq2 & !v3a6ee22;
assign v3a70d3f = hmaster2_p & v37737aa | !hmaster2_p & v373366b;
assign v3a70d7f = hbusreq4_p & v374550d | !hbusreq4_p & v373b671;
assign v377371c = hbusreq7_p & v372c470 | !hbusreq7_p & v37304a0;
assign v3728cb3 = hgrant5_p & v372c4cd | !hgrant5_p & v373fde1;
assign v375a26b = jx0_p & v3a715c4 | !jx0_p & v3779fdf;
assign v3a6fcf1 = hlock7_p & v3a6427b | !hlock7_p & v37257e5;
assign v3752957 = hbusreq6_p & v38093aa | !hbusreq6_p & v372c37f;
assign v3776779 = hmaster1_p & v3a635ea | !hmaster1_p & v3a7138c;
assign v3730be3 = hmaster0_p & v374a6ce | !hmaster0_p & v3a6ef7f;
assign v3a63b56 = hgrant1_p & v37470eb | !hgrant1_p & !v37457fb;
assign v3760d83 = hgrant1_p & v8455ab | !hgrant1_p & !v3a7057b;
assign v3a70cfe = hbusreq4 & v3a70530 | !hbusreq4 & v8455ab;
assign v3769df4 = hbusreq1 & v39a5265 | !hbusreq1 & !v3a6fd79;
assign v3a5e7dc = hmaster2_p & v3778e28 | !hmaster2_p & !v2678c97;
assign v3a54c8b = hmaster2_p & v3a66d43 | !hmaster2_p & v37229f0;
assign v3772374 = hbusreq5_p & v374ab4b | !hbusreq5_p & v376c335;
assign v3761d4e = hbusreq2 & v3745f76 | !hbusreq2 & !v8455ab;
assign v2acaeda = hbusreq4 & v3a2a33d | !hbusreq4 & v3a6134b;
assign ca50c0 = hlock5 & v372afcc | !hlock5 & v3754379;
assign v373c965 = hlock6_p & v3736ded | !hlock6_p & v8455bb;
assign v3747346 = hgrant3_p & v3a6f22b | !hgrant3_p & v3773871;
assign v3a70200 = hlock6_p & v39a5265 | !hlock6_p & !v8455ab;
assign v3807174 = hlock8 & v3a55076 | !hlock8 & v3735d01;
assign v3745801 = hgrant1_p & v8455ab | !hgrant1_p & v3a7162d;
assign v3a6f581 = hgrant3_p & v8455ab | !hgrant3_p & v3a6fea3;
assign v3766f8a = hmaster3_p & v372a8d9 | !hmaster3_p & v3a70eb8;
assign v3767902 = hlock7_p & v376d6b9 | !hlock7_p & !v8455ab;
assign v3a61714 = hmaster0_p & v377be72 | !hmaster0_p & v3a70476;
assign v3a58b3f = hgrant2_p & v8455bd | !hgrant2_p & v39378d6;
assign v3a58673 = hmaster1_p & v8455ab | !hmaster1_p & v3a63dba;
assign v375cf11 = hmaster0_p & v3750faa | !hmaster0_p & !v3a539bf;
assign v3a6f5c0 = hgrant1_p & v8455ab | !hgrant1_p & v376045b;
assign v3a6ecd1 = hlock7_p & v3a5cb92 | !hlock7_p & v3a6eb91;
assign v3a6f75d = hmaster2_p & v3730dc4 | !hmaster2_p & v3763fdc;
assign v37504f9 = hmaster2_p & v37430e7 | !hmaster2_p & v3757da6;
assign v3806fe2 = hmaster0_p & v1e3786e | !hmaster0_p & v373e62a;
assign v3a54811 = hlock0 & v3a5fc82 | !hlock0 & v3724715;
assign v3a665dd = hbusreq2 & v3a6fff7 | !hbusreq2 & v8455ab;
assign v377728d = hgrant2_p & v8455ab | !hgrant2_p & v3a5f5bb;
assign v3743f7a = hmaster0_p & v37760f9 | !hmaster0_p & v3a705e6;
assign v3774829 = hmaster2_p & v1e3824a | !hmaster2_p & v3a63a7a;
assign v3a64089 = hmaster0_p & v3a659d0 | !hmaster0_p & v3a70ad3;
assign v3759031 = hbusreq2_p & v3a654fb | !hbusreq2_p & v8455ab;
assign v37350a4 = hlock5_p & v3a703a7 | !hlock5_p & !v3759265;
assign v372c91d = hlock0_p & v8455ab | !hlock0_p & v3a5d923;
assign v3a5b51d = hmaster1_p & v374b8fa | !hmaster1_p & v376f942;
assign v3731399 = hbusreq3 & v3779fec | !hbusreq3 & v3a6fdef;
assign v3757601 = hgrant2_p & v3750269 | !hgrant2_p & v372834c;
assign v3748ae2 = hbusreq3 & v373adae | !hbusreq3 & v8455ab;
assign v1e379f7 = hgrant2_p & v372aacd | !hgrant2_p & v3a701cd;
assign v372b689 = jx0_p & v8455ab | !jx0_p & v3a5fa09;
assign v3a70cfc = hgrant4_p & v3724e30 | !hgrant4_p & v376cbb7;
assign v39ed7e4 = hgrant5_p & v8455ab | !hgrant5_p & v8455c5;
assign v37554cd = hmaster0_p & v3727f3b | !hmaster0_p & v3a7094f;
assign v377dc15 = hgrant1_p & v376dbdf | !hgrant1_p & !v8455ab;
assign v3a656bd = hgrant5_p & v8455c6 | !hgrant5_p & v375a397;
assign v3746c1d = hmaster0_p & v3765b3c | !hmaster0_p & v375d3fd;
assign v375aaf3 = hbusreq6_p & v3a712d6 | !hbusreq6_p & v3a65e52;
assign v3755dcd = hbusreq3_p & v375a7cd | !hbusreq3_p & v8455ab;
assign v2092b0b = hmaster2_p & v377ea86 | !hmaster2_p & !v8455ab;
assign v37531b1 = hlock4_p & v376430b | !hlock4_p & v8455ab;
assign v3734868 = hmaster1_p & v3a635ea | !hmaster1_p & v375c8c8;
assign v375ed69 = jx0_p & v373765a | !jx0_p & v37510d9;
assign v374d8c9 = hmaster0_p & v3a57584 | !hmaster0_p & v3a6f84c;
assign v372acab = hlock4_p & v3a6fc30 | !hlock4_p & v3a70e4f;
assign v3754565 = hbusreq0 & v3747c90 | !hbusreq0 & b96080;
assign v3766160 = hmaster0_p & v3751dba | !hmaster0_p & v3735f79;
assign v376b1d4 = hbusreq8_p & v3759569 | !hbusreq8_p & v372acd3;
assign v3a6fbcb = hmaster2_p & v3a663b9 | !hmaster2_p & v3a65762;
assign v3a56688 = hbusreq0 & v375e47e | !hbusreq0 & v3a708dd;
assign v28896b4 = hmaster2_p & v8455ab | !hmaster2_p & v3a70e4b;
assign v373e877 = hlock0_p & v8455ab | !hlock0_p & v3a6f776;
assign v3769617 = jx3_p & v377e896 | !jx3_p & v3a67880;
assign v3773575 = hgrant6_p & v37409f4 | !hgrant6_p & v8455ab;
assign v38065f1 = hbusreq5_p & v3775687 | !hbusreq5_p & v3a66632;
assign v3755608 = hbusreq6_p & v3753f1a | !hbusreq6_p & !v8455ab;
assign v3a665d5 = hmaster2_p & v37483ff | !hmaster2_p & v8455ab;
assign v3a6efb6 = hbusreq4_p & v3734067 | !hbusreq4_p & !v3a68b49;
assign v375ff4e = hmaster2_p & v37795d3 | !hmaster2_p & v375a1ab;
assign v3731596 = hbusreq4 & v39a537f | !hbusreq4 & !v8455ab;
assign v3807b9c = jx3_p & v3746559 | !jx3_p & v376c010;
assign v3a712c6 = hbusreq5 & v3a70a37 | !hbusreq5 & v8455ab;
assign v3255a16 = hbusreq6 & v3740171 | !hbusreq6 & v8455ab;
assign v376bb88 = hbusreq3_p & v3751dc9 | !hbusreq3_p & v373b288;
assign v373f401 = hgrant6_p & v8455c9 | !hgrant6_p & v3760aa7;
assign v372c353 = jx0_p & v375cd3f | !jx0_p & v3766a69;
assign v374948b = hbusreq5_p & v3768fba | !hbusreq5_p & v8455ab;
assign v3a68f62 = locked_p & v376189a | !locked_p & !v8455ab;
assign v3a70c67 = hmaster1_p & v3739c6f | !hmaster1_p & v3a5c41b;
assign v3753dbd = hmaster0_p & v3a5bcfd | !hmaster0_p & v375a086;
assign v3a6a52b = hmaster2_p & v377db88 | !hmaster2_p & v3a70c3e;
assign v377b9fd = hmaster0_p & v37567db | !hmaster0_p & v8455ab;
assign v37682c6 = hbusreq1_p & v376e00a | !hbusreq1_p & v3739166;
assign v3a59ba9 = hbusreq6_p & v3a70f78 | !hbusreq6_p & v372bf9f;
assign v3725088 = hbusreq7_p & v2ff8bb1 | !hbusreq7_p & !v3737bfe;
assign v372826c = jx1_p & v37419d7 | !jx1_p & v3727de3;
assign v99aa13 = hmaster2_p & v3a6f92f | !hmaster2_p & v3a70326;
assign v3a701a0 = hgrant6_p & v3a6cb16 | !hgrant6_p & v373f704;
assign v3a70e07 = hbusreq6_p & v372d5bb | !hbusreq6_p & v372b22b;
assign v3a6fea9 = hbusreq4_p & v1e3787a | !hbusreq4_p & !v3a703c3;
assign v3a6f4bc = hgrant2_p & v8455ab | !hgrant2_p & v375c31a;
assign v3a6eb1c = hmaster0_p & v3776865 | !hmaster0_p & v3a59bbd;
assign v3735891 = hmaster2_p & v3a70147 | !hmaster2_p & v37631d9;
assign v3a6fcd4 = hgrant3_p & v8455ab | !hgrant3_p & v3759570;
assign v380760a = hbusreq4_p & v3a5f21c | !hbusreq4_p & !v8455ab;
assign v3a55f0d = hmaster2_p & v8455ab | !hmaster2_p & !v3a63559;
assign v37498be = hgrant0_p & v3733e9e | !hgrant0_p & v3a6f4fc;
assign v376ed58 = hmaster1_p & v8455ab | !hmaster1_p & v3a70712;
assign v375fb71 = hbusreq7_p & v3a6501d | !hbusreq7_p & v3a55c44;
assign v3769c47 = hgrant4_p & v3a602a4 | !hgrant4_p & v3771fbb;
assign v3a6f02f = hbusreq2_p & v3756149 | !hbusreq2_p & v376306b;
assign v375f664 = hmaster2_p & v373164a | !hmaster2_p & !v3a63559;
assign v37406ca = hbusreq6_p & v374faa9 | !hbusreq6_p & v3377b1b;
assign v377c931 = hbusreq0 & v3a6e7d8 | !hbusreq0 & v37713fe;
assign v3747d0e = hlock5 & v3779b31 | !hlock5 & v37496fc;
assign v3a5d06d = hbusreq4 & v3764ca0 | !hbusreq4 & v374e768;
assign v3740352 = hmaster0_p & v3a5cd4c | !hmaster0_p & v3a610f8;
assign v37433f5 = hmaster2_p & v3a6a8ee | !hmaster2_p & v373de4b;
assign v377852a = hbusreq2 & v373a27c | !hbusreq2 & v8455ab;
assign v37384a3 = hmaster2_p & v377bea3 | !hmaster2_p & v372edd9;
assign v3741d52 = hmaster2_p & v3a71377 | !hmaster2_p & v377f32e;
assign v3a706a8 = hmaster2_p & v3763295 | !hmaster2_p & v374e855;
assign v3a59883 = hlock0_p & v377217c | !hlock0_p & v3a70b72;
assign v37642a0 = hlock2 & v3739743 | !hlock2 & v3757ae7;
assign v3759c48 = hgrant5_p & v3756ba5 | !hgrant5_p & v3764d3e;
assign v376bc98 = hbusreq7_p & v3a57e1a | !hbusreq7_p & a5c619;
assign v3753445 = hbusreq8_p & v3a70d60 | !hbusreq8_p & v37258d0;
assign v3a58ef3 = hmaster2_p & v3806db7 | !hmaster2_p & v3a70641;
assign v37393e8 = jx1_p & v37354bf | !jx1_p & v374e1f0;
assign v2aca264 = hbusreq0 & v3760bfd | !hbusreq0 & v377e639;
assign v372eb5c = hmaster2_p & v3a63805 | !hmaster2_p & v8455ab;
assign v3a6ef3e = hlock7_p & v373a58c | !hlock7_p & !v8455ab;
assign v374f87c = hready & v3a690ec | !hready & v376c211;
assign v3a5dd17 = hlock6 & v375c9ea | !hlock6 & v3a6006a;
assign v3732eca = stateA1_p & v8455ab | !stateA1_p & v372b7fb;
assign v3a6d897 = hmaster2_p & v3776323 | !hmaster2_p & v374b0cb;
assign v373ec80 = hbusreq7_p & v3777d70 | !hbusreq7_p & v3762c4c;
assign v3741384 = hgrant4_p & v3a5e63b | !hgrant4_p & v3a70e69;
assign v3a6d874 = hmaster0_p & v3a6f8a7 | !hmaster0_p & !v3a539bf;
assign v3764ca0 = hgrant6_p & v3760a55 | !hgrant6_p & v377868e;
assign dac328 = hbusreq4_p & v3763d52 | !hbusreq4_p & v375ebe9;
assign v3a6fb4b = hmaster1_p & v3a5e0b8 | !hmaster1_p & v3727187;
assign v3a6f240 = hbusreq0 & v3767437 | !hbusreq0 & !v8455ab;
assign v3730828 = hmaster1_p & v373e474 | !hmaster1_p & v3a61a2d;
assign v37258b4 = hmaster0_p & v360d136 | !hmaster0_p & v372309d;
assign v3768048 = hmaster1_p & v3a6c5e5 | !hmaster1_p & v8455ca;
assign v374673a = hgrant6_p & v8455ab | !hgrant6_p & v3773bc6;
assign v3a7087f = hbusreq8 & v3a6ec28 | !hbusreq8 & v3740380;
assign v3809cc0 = hmaster0_p & v3753825 | !hmaster0_p & v376d21d;
assign v3a581fb = hbusreq8 & v380987d | !hbusreq8 & v8455ab;
assign v376121f = hbusreq2 & v375d009 | !hbusreq2 & v3757955;
assign v3746a45 = hbusreq8 & v3a5740f | !hbusreq8 & v8455ab;
assign v3746888 = hgrant3_p & v377f76a | !hgrant3_p & !v2092f20;
assign v376e68d = hbusreq7 & v3a6ff0e | !hbusreq7 & v3a6f1d8;
assign v3a70df8 = hbusreq7 & v3731555 | !hbusreq7 & !v8455b9;
assign v3776da7 = hmaster0_p & v3769ad5 | !hmaster0_p & v3a6f3b9;
assign v3a6facd = hmaster2_p & v8455ab | !hmaster2_p & v374ca62;
assign v3a5445c = hbusreq7 & v374cff2 | !hbusreq7 & v3730568;
assign v3743366 = hbusreq3 & v3a6f77c | !hbusreq3 & v3725cbf;
assign v3a71066 = hmaster2_p & v3a6d590 | !hmaster2_p & v374ab8d;
assign v3a71276 = hgrant4_p & v8455ab | !hgrant4_p & v3a6fd5e;
assign v3a6fc7a = hbusreq4_p & v37250fa | !hbusreq4_p & v3a702e1;
assign v3a7167d = hmaster2_p & v3754dd0 | !hmaster2_p & v3730a3d;
assign v3a6b463 = stateG3_2_p & v8455ab | !stateG3_2_p & !v845601;
assign v3757956 = hgrant4_p & v375da82 | !hgrant4_p & v3775999;
assign v376189d = hmaster2_p & v3753837 | !hmaster2_p & v3a70d85;
assign v374ef4a = hbusreq5_p & v3a70f2d | !hbusreq5_p & !v375b342;
assign v3732a04 = hbusreq8 & v373b17e | !hbusreq8 & v3774eed;
assign v373d27f = hgrant4_p & v372cab6 | !hgrant4_p & v3a6f9c4;
assign v3756202 = hgrant5_p & v373bdd9 | !hgrant5_p & v3a6f8b9;
assign v375e6ed = hgrant6_p & v3807003 | !hgrant6_p & v37450ff;
assign v376d542 = hgrant5_p & v3a70578 | !hgrant5_p & v3a6f70b;
assign v3a704c3 = jx0_p & v3a53cc2 | !jx0_p & v3769e46;
assign v3a62cb7 = hmaster0_p & v3742035 | !hmaster0_p & v3a56002;
assign v8455fd = stateA1_p & v8455ab | !stateA1_p & !v8455ab;
assign v3a6e91d = hlock2 & v3a6f613 | !hlock2 & v3a70eb6;
assign v3a6eaba = hmaster0_p & v3a619c0 | !hmaster0_p & v3724c9c;
assign v375b0d4 = hmaster2_p & v372615f | !hmaster2_p & v3258762;
assign v377abbe = jx0_p & v8455ab | !jx0_p & v374888e;
assign v372c09e = hbusreq8 & v375d3bb | !hbusreq8 & !v376053b;
assign v372ee5a = hbusreq5_p & v3749242 | !hbusreq5_p & v3746008;
assign v374304d = hbusreq0 & v37554d5 | !hbusreq0 & v374052a;
assign v377754d = hgrant2_p & v376e914 | !hgrant2_p & v373f4a5;
assign v3a6e6fa = hbusreq0 & v377c079 | !hbusreq0 & v3a67833;
assign v3a6eb52 = hbusreq2 & v37482f8 | !hbusreq2 & !v3a703df;
assign v23fdc46 = hgrant2_p & v8455ab | !hgrant2_p & v38063c6;
assign v3a6844c = jx0_p & v3729113 | !jx0_p & v3728a4a;
assign v3777b84 = hgrant5_p & v3739239 | !hgrant5_p & v3734129;
assign v373c387 = hgrant3_p & v3a70c36 | !hgrant3_p & v376c1cc;
assign v1e382dc = hgrant7_p & v3a614df | !hgrant7_p & v3a6c40d;
assign v3a6f726 = hmaster0_p & v37240a4 | !hmaster0_p & v3770fa1;
assign v3761d38 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f2d1;
assign v3a6f29c = hbusreq0 & v373f401 | !hbusreq0 & v3726865;
assign v377f83c = hlock2 & v3752fb7 | !hlock2 & v3769c81;
assign v374ab03 = hmaster0_p & v3a70bba | !hmaster0_p & v3746a7e;
assign b4ac83 = hbusreq0 & v3757ecc | !hbusreq0 & v3a70062;
assign v373ec96 = hmaster1_p & v3a67577 | !hmaster1_p & v3a70a01;
assign v3a6fe06 = hgrant2_p & v3758472 | !hgrant2_p & !v3768d79;
assign v3734658 = hbusreq5_p & v377535e | !hbusreq5_p & v3a70a99;
assign v3a63331 = hlock4 & v3a70525 | !hlock4 & v3768349;
assign v3a70961 = hmaster0_p & v3753a2e | !hmaster0_p & v376b540;
assign v3a65ae2 = hmaster1_p & v3745181 | !hmaster1_p & v377b0a3;
assign v3770db3 = hmaster2_p & v3a6937a | !hmaster2_p & v372f100;
assign v375ceee = hmaster2_p & v377a3bd | !hmaster2_p & v374a08a;
assign v3726d97 = hbusreq2 & v372da76 | !hbusreq2 & v3a6fdef;
assign v3777602 = hbusreq7 & v376f1d0 | !hbusreq7 & v3737808;
assign v374ac6d = hmaster1_p & v3a672e6 | !hmaster1_p & !v8455ab;
assign v372ec65 = hmaster0_p & v38097ee | !hmaster0_p & v3779f51;
assign v3762790 = hbusreq5 & v3809f61 | !hbusreq5 & v8455ab;
assign v377c2ba = hgrant1_p & v8455e7 | !hgrant1_p & !v8455ab;
assign v3a6a2f8 = hmaster2_p & v8455e7 | !hmaster2_p & v376dbdf;
assign v377773f = hlock2_p & v377814b | !hlock2_p & v3a6ef74;
assign v3a6f6c0 = hmaster0_p & v3766d0a | !hmaster0_p & v3777da6;
assign v3727c74 = hmaster1_p & v3a635ea | !hmaster1_p & v37579f7;
assign v3762617 = hmaster1_p & v37411ab | !hmaster1_p & v3a5f869;
assign v3a6f90a = hbusreq2_p & v3a70635 | !hbusreq2_p & v374d479;
assign v3a622c0 = hbusreq1 & v37328bf | !hbusreq1 & v8455ab;
assign v375588c = hbusreq0_p & v375da10 | !hbusreq0_p & v376bb26;
assign v374b07a = hbusreq3 & v3a7045c | !hbusreq3 & v8455ab;
assign v3764b3f = hbusreq2_p & v3a70e85 | !hbusreq2_p & v8455ab;
assign v3a70c7a = hlock4 & v3a7056c | !hlock4 & v3727713;
assign v380777f = hbusreq4_p & v3750dd3 | !hbusreq4_p & v3a5f984;
assign v377113b = hlock8 & v3a6fa20 | !hlock8 & v3a5faf0;
assign v3773e17 = hmaster2_p & v3a66ade | !hmaster2_p & v37c048c;
assign v3a71566 = hlock4 & v3a7005e | !hlock4 & v3739635;
assign v3a6f902 = hbusreq4 & v3a5b68a | !hbusreq4 & !v8455ab;
assign v37760f9 = hmaster2_p & v3a70374 | !hmaster2_p & v3a5b7db;
assign v376fd32 = hmaster0_p & v3a706dc | !hmaster0_p & v3a6fcab;
assign v3751c12 = start_p & v3730a0f | !start_p & v8455ab;
assign v38072bd = hmaster2_p & v3a635ea | !hmaster2_p & v3a6f2cb;
assign v3a6fdbf = hmaster2_p & v376a14f | !hmaster2_p & v3733383;
assign v3a6bc65 = hbusreq2_p & v372cedb | !hbusreq2_p & !v8455ab;
assign v375e30b = hlock5 & v3736fb4 | !hlock5 & v3a7114a;
assign v3a65aa5 = hbusreq5_p & v3778a97 | !hbusreq5_p & v372834d;
assign v37651c2 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3a63621;
assign v3a5899d = hlock4 & v3773e77 | !hlock4 & v376bea3;
assign v376b903 = hbusreq6_p & v3a70409 | !hbusreq6_p & v3a59517;
assign v3a53a94 = hbusreq4_p & v3759032 | !hbusreq4_p & v3733e9e;
assign v3774247 = hmaster2_p & v3a635ea | !hmaster2_p & v377d58d;
assign v3a6ef62 = hbusreq3_p & v376f56d | !hbusreq3_p & v377f200;
assign v377c065 = hmaster2_p & v3769d48 | !hmaster2_p & v3a6f4ba;
assign v374fc17 = hbusreq5_p & v374aed5 | !hbusreq5_p & v375a187;
assign v3a6f36d = hmaster2_p & v372d905 | !hmaster2_p & v377955b;
assign v35ba1a5 = hbusreq2_p & v3a5a035 | !hbusreq2_p & v8455ab;
assign v376c422 = hmaster0_p & v37688d1 | !hmaster0_p & v3a7114b;
assign v8455cb = hlock6_p & v8455ab | !hlock6_p & !v8455ab;
assign v3735350 = jx0_p & v3a7084f | !jx0_p & v37716e1;
assign v3753942 = hbusreq8 & v2092a89 | !hbusreq8 & v3733173;
assign v376ad77 = hmaster2_p & v375058e | !hmaster2_p & !v8455ab;
assign v377f669 = hgrant3_p & v8455ab | !hgrant3_p & v377f27f;
assign v376305b = hbusreq6_p & v3a67729 | !hbusreq6_p & v37306cd;
assign v3749ec6 = hmaster2_p & v3779060 | !hmaster2_p & v375c5a8;
assign v3a68a46 = hmaster2_p & v3a6fc5e | !hmaster2_p & v3769740;
assign v3767e55 = hmaster2_p & v3a71133 | !hmaster2_p & v3772696;
assign v3a70893 = hbusreq3_p & v924b19 | !hbusreq3_p & v8455ab;
assign v3a6765d = hmaster2_p & v377f734 | !hmaster2_p & v3774647;
assign v373e85a = hgrant0_p & v3a5b5d3 | !hgrant0_p & !v374790d;
assign v3a70b5b = hbusreq5_p & v372d891 | !hbusreq5_p & v3a6fc77;
assign v373026e = hmaster2_p & v3a64a09 | !hmaster2_p & v3a708c2;
assign v376b962 = hready_p & v3732f65 | !hready_p & v3a7124f;
assign v37270a2 = hmaster2_p & v376bd43 | !hmaster2_p & !v8455ab;
assign v372650c = hgrant4_p & v37579c1 | !hgrant4_p & !v8455ab;
assign v3a6b2ef = hbusreq1_p & v37362ea | !hbusreq1_p & v3a6d922;
assign v3736ae6 = hmaster1_p & v3a71343 | !hmaster1_p & v377f264;
assign v23fdf1b = hmaster2_p & v3732e59 | !hmaster2_p & v360d0fd;
assign v3a57cb4 = hgrant0_p & v3a696ed | !hgrant0_p & ccdd71;
assign v3a5d55b = hbusreq8 & v3a70e4a | !hbusreq8 & v3759284;
assign v373b747 = hbusreq5_p & v3a71557 | !hbusreq5_p & v8455ab;
assign v3764015 = hmaster2_p & v3770abd | !hmaster2_p & v3745b02;
assign v3775606 = hmaster0_p & v372ad5d | !hmaster0_p & v3a6ff97;
assign v3730b63 = hgrant6_p & v8455ab | !hgrant6_p & v3a6a95e;
assign v37324c0 = hmastlock_p & v376282b | !hmastlock_p & v8455ab;
assign v3a6bedb = hgrant6_p & v3752957 | !hgrant6_p & v3749bef;
assign v376a752 = hmaster0_p & v37566b2 | !hmaster0_p & v3a5d994;
assign v37494a9 = hgrant4_p & v8455ab | !hgrant4_p & v3768538;
assign v37474dc = hlock0 & v372f1b8 | !hlock0 & v23fe175;
assign v3742360 = hmaster1_p & v377adf5 | !hmaster1_p & v3a6fb9b;
assign v3a5797b = hgrant3_p & v8455be | !hgrant3_p & v374ce92;
assign v3a6ebae = hlock0 & v3a7164a | !hlock0 & v3a603ad;
assign v375082a = hbusreq3 & v23fd7d9 | !hbusreq3 & v8455b0;
assign v37266bd = hbusreq8_p & v3a6f7b8 | !hbusreq8_p & v3736dfd;
assign v37634cf = hmaster0_p & v3a6f475 | !hmaster0_p & v3a71614;
assign v3727bc6 = hmaster0_p & v23fe20d | !hmaster0_p & v3a70a2b;
assign v3a6b0a1 = hmaster1_p & v8455ab | !hmaster1_p & v3a6f039;
assign v3a6f6ca = hmaster1_p & v376aa54 | !hmaster1_p & v3a6fcbe;
assign v3a6582d = jx0_p & v373738e | !jx0_p & v8455ab;
assign v373de4b = hbusreq4_p & v3a64dc2 | !hbusreq4_p & v8455ab;
assign v3a6180b = hgrant6_p & v37658d7 | !hgrant6_p & v3a61482;
assign v372c5da = hlock4 & v372a39d | !hlock4 & v376d9aa;
assign v3a6196d = hbusreq5 & v3a5b719 | !hbusreq5 & c7ae7d;
assign v3a7152c = hgrant2_p & v3779060 | !hgrant2_p & v372fd97;
assign v3a5417e = hbusreq4_p & v373109c | !hbusreq4_p & v3a5c50b;
assign v3a6c688 = hlock2_p & v375a99b | !hlock2_p & v3a669ae;
assign v3a71664 = hbusreq8 & v3737711 | !hbusreq8 & v3a6f4f7;
assign v974eb9 = hbusreq5_p & v37366d5 | !hbusreq5_p & v3a60d50;
assign v377abcb = hbusreq0 & v3775e78 | !hbusreq0 & v377c9cc;
assign v376f39f = hbusreq7_p & v375ae3d | !hbusreq7_p & v3a6e33a;
assign v3a6ff46 = hmaster2_p & v8455ab | !hmaster2_p & !b62916;
assign v3a5cc79 = hmaster0_p & v3a70743 | !hmaster0_p & v8455e7;
assign v374e538 = hmaster1_p & v3a56b92 | !hmaster1_p & v374776b;
assign v3a579da = hbusreq8 & v376dacb | !hbusreq8 & v8455b3;
assign v377346e = hmaster2_p & v3770f96 | !hmaster2_p & v8455ab;
assign v3745b51 = hbusreq7_p & v2acaeaa | !hbusreq7_p & v3a70eb7;
assign v3a64190 = hbusreq0 & v374c6e1 | !hbusreq0 & v3757b55;
assign v3a7114a = hbusreq5 & v376e74b | !hbusreq5 & v3762a76;
assign v3a54f85 = hbusreq6 & v3766b81 | !hbusreq6 & v3a635ea;
assign v3a701ec = hmaster0_p & v3a66ade | !hmaster0_p & v3a71667;
assign v3a69203 = hgrant5_p & v8455ab | !hgrant5_p & v377ea20;
assign ae0bd0 = hmaster0_p & v37350f0 | !hmaster0_p & v372b3f6;
assign v373d338 = hgrant2_p & v3731b33 | !hgrant2_p & v377b983;
assign v3a58cd5 = hmastlock_p & v3727fe3 | !hmastlock_p & v8455ab;
assign v3a70995 = hbusreq6 & v377aa23 | !hbusreq6 & v3a70a88;
assign v372bbab = hmaster1_p & v3727d4c | !hmaster1_p & v374a7b4;
assign v1e37519 = hgrant4_p & v37466cb | !hgrant4_p & v3771913;
assign v377ea73 = hbusreq3 & v39a5265 | !hbusreq3 & !v3a6b6f3;
assign v924b19 = hbusreq3 & v3a70641 | !hbusreq3 & v8455ab;
assign v3742de5 = hbusreq7_p & v3a575d5 | !hbusreq7_p & v375bc6f;
assign v3a5fee0 = hmaster2_p & v3806db0 | !hmaster2_p & v3a7106c;
assign v377246f = hmaster1_p & v35b7169 | !hmaster1_p & v3731826;
assign v3774908 = hbusreq6_p & v37494bb | !hbusreq6_p & v3a5b91d;
assign v3756fee = jx0_p & v3a62e99 | !jx0_p & v38074ed;
assign v37270ad = hmaster0_p & v3a6dfb2 | !hmaster0_p & v37559b4;
assign v3806640 = decide_p & v376b3a9 | !decide_p & v3903ee6;
assign v3746f84 = hlock0_p & v3773b23 | !hlock0_p & v8455b0;
assign v38076bb = hlock5 & v3779a9c | !hlock5 & v37565a6;
assign v3733392 = jx0_p & v374431a | !jx0_p & v3766a7d;
assign v3a70fda = hgrant4_p & v3741925 | !hgrant4_p & !v8455ab;
assign v3744202 = hbusreq7_p & v3a59a60 | !hbusreq7_p & !v3747141;
assign v3725bb3 = hmaster1_p & v375b429 | !hmaster1_p & v3738ed2;
assign v3a711db = hmaster2_p & v3744b55 | !hmaster2_p & v37425c6;
assign v376d327 = hlock1 & v3a712a3 | !hlock1 & v3a6ebb7;
assign v3768da7 = hmaster0_p & v3735c06 | !hmaster0_p & v8455ab;
assign v23fe159 = hbusreq2_p & v377eaf2 | !hbusreq2_p & v3778528;
assign v3727b10 = hmaster0_p & v376166b | !hmaster0_p & v3807a26;
assign v375361a = hbusreq2 & v3a63805 | !hbusreq2 & v3755791;
assign v3757407 = hlock0 & v372348c | !hlock0 & v3a710eb;
assign v3a5a647 = hbusreq0_p & v3a71452 | !hbusreq0_p & v3743b9e;
assign v3a70254 = hbusreq7_p & v374727f | !hbusreq7_p & !v373580c;
assign v37366d2 = hgrant0_p & v3743b9e | !hgrant0_p & v3a706c7;
assign v3a57ec9 = hlock4 & v3a71569 | !hlock4 & cc4895;
assign v3773165 = hlock8_p & v3806a7a | !hlock8_p & !v8455ab;
assign v37612f7 = hgrant6_p & v3734967 | !hgrant6_p & v3749d74;
assign v3a6b908 = hbusreq2_p & v3752201 | !hbusreq2_p & v380854b;
assign v374df4b = hbusreq4 & v373a755 | !hbusreq4 & !v3a640a0;
assign v377c8ca = hmaster1_p & v8455ab | !hmaster1_p & v372b48a;
assign v374baea = hlock0 & v3a708c2 | !hlock0 & v3a64cfa;
assign v37551df = hgrant2_p & v3771696 | !hgrant2_p & !d138a6;
assign v373c7af = hgrant5_p & v37465c7 | !hgrant5_p & !v8455ab;
assign v3750c9f = hlock4_p & v373b36c | !hlock4_p & v3722a7e;
assign v3a70892 = hbusreq8 & v37551eb | !hbusreq8 & v8455ab;
assign v3a710cb = hbusreq6_p & v375bdd4 | !hbusreq6_p & v375dbd4;
assign v3a67971 = hmaster0_p & v3a5c7be | !hmaster0_p & v3750088;
assign v3764601 = hlock0 & v373031f | !hlock0 & v3a7073b;
assign dac346 = hgrant3_p & v8455ab | !hgrant3_p & v3a6831c;
assign v3a57db8 = hbusreq4_p & v374b32b | !hbusreq4_p & v3a701e9;
assign v3731eb5 = hbusreq6 & v377ed8e | !hbusreq6 & v8455cb;
assign v377c023 = hlock4 & v3748797 | !hlock4 & v3a6eb1b;
assign v3a711f0 = hgrant1_p & v377de41 | !hgrant1_p & !v3727a6c;
assign v373505c = hmaster2_p & v373f6ee | !hmaster2_p & v376a056;
assign v3752091 = hbusreq8_p & v3a6a40b | !hbusreq8_p & v3765395;
assign v3a5db94 = hmaster2_p & v3779183 | !hmaster2_p & v37674f6;
assign v3a705aa = hbusreq7 & v373f2d2 | !hbusreq7 & v376ae9f;
assign v372b982 = stateA1_p & v2aca977 | !stateA1_p & !v38073d4;
assign v3a5f38a = hbusreq6 & v3a70180 | !hbusreq6 & v3765e79;
assign v373a4a8 = hmaster1_p & v3a5fc34 | !hmaster1_p & v3753bb4;
assign v3a6eba5 = hlock6 & v3a5fbb0 | !hlock6 & v3759c6c;
assign v3a68b74 = hbusreq2_p & v3a6eb6b | !hbusreq2_p & v37305cc;
assign v3a7167c = hgrant5_p & v37751bb | !hgrant5_p & v3776d42;
assign v3a6f2b6 = hbusreq4 & v374282f | !hbusreq4 & v376fcc3;
assign v3a70a4f = hbusreq4 & v374ffb7 | !hbusreq4 & v373785d;
assign v375bdf0 = hgrant3_p & v3726139 | !hgrant3_p & v3a63135;
assign v37643af = hgrant6_p & beb1cf | !hgrant6_p & v374d183;
assign v375d559 = hlock6 & v3770e30 | !hlock6 & v3a6006a;
assign v375ac98 = hlock1_p & v3a651b8 | !hlock1_p & v8455b0;
assign v3a65e3c = hbusreq0 & v37660dd | !hbusreq0 & v8455ab;
assign v377047f = hbusreq8_p & v3763086 | !hbusreq8_p & v373c30e;
assign v3773a5b = hbusreq6 & v3732706 | !hbusreq6 & v3765261;
assign v37486e9 = hmaster0_p & v3762e13 | !hmaster0_p & v374a0ae;
assign v3742259 = hbusreq0_p & v3a70641 | !hbusreq0_p & v8455ab;
assign v3a70cdf = hgrant0_p & v8455ab | !hgrant0_p & v3a6b297;
assign v3a5aa5c = hbusreq5 & v38073e8 | !hbusreq5 & v3764dac;
assign v377b626 = hbusreq5_p & v3a53f85 | !hbusreq5_p & v375aceb;
assign v376e643 = hbusreq3 & v3740171 | !hbusreq3 & v8455e7;
assign v3741920 = hbusreq8 & v8455e7 | !hbusreq8 & v374757c;
assign v37291ce = hlock0_p & v3a6f018 | !hlock0_p & !v8455ab;
assign v3a6da5a = hgrant4_p & v3731c6f | !hgrant4_p & v3a5de8f;
assign v37781ac = hbusreq6_p & v375685b | !hbusreq6_p & v3775d1d;
assign v3738aa6 = hbusreq7 & v376a9f5 | !hbusreq7 & v377a2b2;
assign v37623b8 = hbusreq6_p & v3748797 | !hbusreq6_p & v376d4ca;
assign bb70de = hmaster0_p & v3750b02 | !hmaster0_p & v372f260;
assign v374e8c3 = hlock8_p & v3a713b4 | !hlock8_p & v35772a6;
assign v374cd6b = hmaster1_p & v372cb06 | !hmaster1_p & v3a6f62f;
assign v3a6fc05 = hmaster2_p & v3762a9f | !hmaster2_p & v37683c2;
assign v3a6e543 = hbusreq0 & v3760f4e | !hbusreq0 & v8455ab;
assign v373e62a = hmaster2_p & v1e3786e | !hmaster2_p & v8455ab;
assign v372ccc4 = hbusreq4 & v35b7808 | !hbusreq4 & v375a16d;
assign v3a5a81d = hmaster0_p & v375be63 | !hmaster0_p & v375c76b;
assign v3a697e4 = hlock4 & v373ff1c | !hlock4 & v3a7024c;
assign v3a70f28 = hlock0 & v3a70126 | !hlock0 & v3764270;
assign v3a6a57c = hmaster0_p & v377a3bd | !hmaster0_p & v375ceee;
assign v373997b = hbusreq1_p & v3a711b7 | !hbusreq1_p & v8455ab;
assign v372ab80 = hmaster0_p & v376d81c | !hmaster0_p & v3745704;
assign v37442e1 = hbusreq0 & v1e374ce | !hbusreq0 & v373c856;
assign v3a71398 = jx0_p & v3726a78 | !jx0_p & v3767cc0;
assign v37307dd = hbusreq6_p & v8455b3 | !hbusreq6_p & v3767437;
assign v3a67ab5 = hmaster2_p & v37356f0 | !hmaster2_p & v3a6dc08;
assign v3763c0d = hmaster1_p & v373732f | !hmaster1_p & v375918d;
assign v2093083 = hmaster2_p & v3a635ea | !hmaster2_p & v3a6efea;
assign v3a6a4d4 = hgrant3_p & v3a704bd | !hgrant3_p & v8455ab;
assign v3a6f6bf = hlock5 & v37707db | !hlock5 & v3a703aa;
assign v37763b2 = hmaster0_p & v376c644 | !hmaster0_p & v373665b;
assign v3741ba8 = hmaster0_p & v2acae60 | !hmaster0_p & !v3752281;
assign v3a64ee3 = hburst1 & v39a537f | !hburst1 & v375c69e;
assign v3723701 = hbusreq4_p & v3764381 | !hbusreq4_p & v3731e31;
assign v3729cfa = hmaster0_p & v3a29da0 | !hmaster0_p & v37509a9;
assign v375a5a1 = hmaster2_p & v8455ab | !hmaster2_p & !v3a5cebb;
assign v3a6973f = hmaster1_p & v3754c02 | !hmaster1_p & v3a6fcbe;
assign v373fd7b = hbusreq5_p & v372feea | !hbusreq5_p & v8455ab;
assign v372af35 = hbusreq7_p & v373a8be | !hbusreq7_p & v3779015;
assign v3a6f9ed = hmaster2_p & v376aa76 | !hmaster2_p & v376d1bb;
assign v3a66c5b = hmaster2_p & v3747302 | !hmaster2_p & v37716ca;
assign v3a685ee = hgrant5_p & v3a69714 | !hgrant5_p & v3a712cc;
assign v3a6c55a = hlock0_p & v3a5980d | !hlock0_p & v3770187;
assign v3a63ac4 = hmaster1_p & v3a703d7 | !hmaster1_p & v3a6f4da;
assign v3a704f1 = hbusreq6 & adf78a | !hbusreq6 & v8455ab;
assign v3a66d3e = hmaster2_p & v3778a0a | !hmaster2_p & v8455ab;
assign v3738fba = hbusreq3_p & v3743f94 | !hbusreq3_p & v3a5cd20;
assign v37627a2 = hmaster0_p & v3770c59 | !hmaster0_p & v3779a60;
assign v3a6e3f0 = hbusreq6 & v3a69488 | !hbusreq6 & v37554c0;
assign v374e9ac = hgrant2_p & v35b774b | !hgrant2_p & v373bff4;
assign v372ce94 = hlock7 & v3a6fec6 | !hlock7 & v3a55491;
assign v374446c = hgrant4_p & v8455ab | !hgrant4_p & v3a70432;
assign v37429c5 = hmaster1_p & v3764e58 | !hmaster1_p & v373d5ac;
assign v3732588 = hbusreq2 & v3a6eab3 | !hbusreq2 & v8455ab;
assign v374d751 = hlock4_p & v3730627 | !hlock4_p & v8455b7;
assign v3772021 = hbusreq5 & v374d13d | !hbusreq5 & v373790d;
assign v3767018 = hbusreq6 & v3a70200 | !hbusreq6 & !v37238b1;
assign v37338d8 = hbusreq2_p & v3a65da7 | !hbusreq2_p & !v8455ab;
assign v3a6fcb0 = hbusreq4_p & v380881d | !hbusreq4_p & v3758e7b;
assign v375588a = hlock5_p & v377bd17 | !hlock5_p & v372d925;
assign v377cbf0 = hmaster1_p & v372ec9f | !hmaster1_p & v3773ee7;
assign v3a6002a = hlock0 & v374d0e3 | !hlock0 & v3a7068a;
assign v375eb29 = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v3a5b7c2;
assign v3739aa6 = hgrant6_p & v37436bc | !hgrant6_p & v3a6f431;
assign v3743172 = hgrant7_p & v3a6e0bf | !hgrant7_p & v37367ba;
assign v373fd72 = hbusreq0 & v374f3e3 | !hbusreq0 & v373e814;
assign v3771026 = hgrant3_p & v3a67b5e | !hgrant3_p & !v37649ee;
assign v375983d = hgrant6_p & v375c7b9 | !hgrant6_p & v37458a3;
assign v3774b58 = hbusreq8_p & v374f838 | !hbusreq8_p & v3735113;
assign v3a6f388 = hmaster0_p & v3734062 | !hmaster0_p & v37698a1;
assign v372de3b = hgrant4_p & v8455ab | !hgrant4_p & v374ce71;
assign v3a66a86 = hmaster3_p & v3751981 | !hmaster3_p & !v3732cf6;
assign v3a676ce = hbusreq4_p & v3a5d80f | !hbusreq4_p & v8455c9;
assign v3a6f951 = hbusreq7_p & v3755d8e | !hbusreq7_p & v37289b0;
assign v3a67dab = hmaster2_p & v373366b | !hmaster2_p & v3758133;
assign v3728e09 = hbusreq1_p & v39a537f | !hbusreq1_p & !v1e38224;
assign v37334fc = hmaster2_p & v377766c | !hmaster2_p & !v37536ae;
assign v33782e5 = hbusreq0 & v3a67b28 | !hbusreq0 & v37734f8;
assign v9864ec = hbusreq8 & v37592d5 | !hbusreq8 & v3744b11;
assign v373446a = hbusreq4_p & v377b0f7 | !hbusreq4_p & v374877e;
assign v3777140 = jx0_p & v376bc5b | !jx0_p & v8455ab;
assign v37524c6 = start_p & v3746bdb | !start_p & v37794be;
assign v3a6f86a = hlock5 & v372a460 | !hlock5 & v9ae4c2;
assign v375c463 = hgrant2_p & v375c55a | !hgrant2_p & v3a7036a;
assign v374663d = hgrant6_p & v8455ab | !hgrant6_p & v374a096;
assign v377e6f5 = hmaster2_p & v3a6f018 | !hmaster2_p & v3754aa3;
assign v37431bb = hmaster0_p & v3a70538 | !hmaster0_p & v3722caa;
assign v374dafa = hgrant2_p & v3a5f50e | !hgrant2_p & v375c6c7;
assign v3a704cc = hbusreq4 & v3a70c39 | !hbusreq4 & v8455ab;
assign v3a64608 = hmaster2_p & v3a61a7f | !hmaster2_p & v3a70a88;
assign v3738114 = hlock6_p & v375bf9a | !hlock6_p & v3755791;
assign v374a8da = hmaster0_p & v377f5e0 | !hmaster0_p & v8455ab;
assign v3a55395 = hgrant4_p & v8455ab | !hgrant4_p & v39a4dd6;
assign v3755a02 = hbusreq4_p & v374550d | !hbusreq4_p & v3a6fdcc;
assign v37740ec = hgrant6_p & v3773044 | !hgrant6_p & v3a70ce6;
assign v3778dd7 = hbusreq4 & v3762312 | !hbusreq4 & v3a5cd72;
assign v3a5987a = hlock0 & v3756eca | !hlock0 & v23fe175;
assign v3a67133 = jx1_p & v3a6deec | !jx1_p & v373dce8;
assign v372e9f3 = hbusreq2_p & v3747302 | !hbusreq2_p & v372310a;
assign v3730bae = hmaster0_p & v374b077 | !hmaster0_p & v377bbf7;
assign v3762613 = hbusreq5_p & v8455ab | !hbusreq5_p & v3a6dd22;
assign v374cf20 = hbusreq2_p & v3755026 | !hbusreq2_p & v3745484;
assign v375eeb0 = hlock4 & v3748797 | !hlock4 & v3a71197;
assign v37501fd = hgrant3_p & v8455ab | !hgrant3_p & c32250;
assign v3a702e9 = hmaster2_p & v3759a34 | !hmaster2_p & v2ff8e1f;
assign v3a63057 = hgrant1_p & v3755791 | !hgrant1_p & !v375b737;
assign v3a704c4 = hlock7_p & v3a70f2e | !hlock7_p & v3773076;
assign v3771696 = hbusreq2_p & v372391f | !hbusreq2_p & !v375c5a8;
assign v3732d3e = hmaster2_p & v3a6ff25 | !hmaster2_p & v3731210;
assign v37654e1 = hmaster1_p & v8455ab | !hmaster1_p & !v3757490;
assign v3779015 = hlock8_p & v377e031 | !hlock8_p & v8455cf;
assign v375d9a7 = hbusreq6 & v37353b5 | !hbusreq6 & v8455ab;
assign v3736d97 = hmaster0_p & v9b63b0 | !hmaster0_p & v3778277;
assign v375aea8 = hgrant5_p & v377673f | !hgrant5_p & v3779d6b;
assign v3762072 = hlock4_p & v3725410 | !hlock4_p & v8455b7;
assign v3a6194e = hmaster1_p & v8455ab | !hmaster1_p & v3a6f1f5;
assign v3a70cd3 = hlock2_p & v3a55844 | !hlock2_p & v3734465;
assign v3750134 = hgrant2_p & v372d3e8 | !hgrant2_p & v3a6fc7b;
assign v3a5acd5 = hgrant6_p & v3771b2c | !hgrant6_p & v3757601;
assign v373945c = hlock8 & v3a64a5d | !hlock8 & d3a24d;
assign v3a635c3 = hgrant2_p & v8455e7 | !hgrant2_p & !v8455ab;
assign v37565c3 = hmaster2_p & v3a5b5d3 | !hmaster2_p & v3770559;
assign v3768b80 = hbusreq5 & v3731e16 | !hbusreq5 & v3745871;
assign v375a71d = hbusreq7_p & v3a70d60 | !hbusreq7_p & v37548be;
assign v37737c9 = hgrant2_p & v374bf8a | !hgrant2_p & v3a5b539;
assign v3808dd0 = hmaster0_p & v3a7128b | !hmaster0_p & v37614c1;
assign v374c297 = hgrant5_p & v3a68707 | !hgrant5_p & v3a56855;
assign v374ad30 = hbusreq6_p & v3a635ea | !hbusreq6_p & v37445f1;
assign v3a7136f = locked_p & v3763ad3 | !locked_p & !v8455ab;
assign v3a5986c = hbusreq4_p & v3a71513 | !hbusreq4_p & v372c219;
assign v3a70180 = hbusreq2_p & v37701cf | !hbusreq2_p & v373b288;
assign v37521ff = hbusreq1 & v3a581bd | !hbusreq1 & v3a70a12;
assign v3770c99 = hmaster0_p & v3a6c6ec | !hmaster0_p & v372fba0;
assign v3732701 = hbusreq4_p & v373330f | !hbusreq4_p & v8455ab;
assign v3a70c06 = hbusreq7 & v3746746 | !hbusreq7 & v3a6639e;
assign v3a5a035 = hlock2_p & v8455ab | !hlock2_p & v39a5265;
assign v3a709e5 = hgrant4_p & v3735cb3 | !hgrant4_p & v3a58d63;
assign v373fe0d = hlock7 & v372c3c0 | !hlock7 & v3739f1d;
assign v3a711b5 = hbusreq4 & v3a6f7fd | !hbusreq4 & v8455ab;
assign v3a625c9 = hbusreq4 & v3723903 | !hbusreq4 & v3a635ea;
assign v3a6a64a = hbusreq5_p & v37400ba | !hbusreq5_p & v37775dd;
assign v3736a75 = hmaster2_p & v3a5d678 | !hmaster2_p & v377ca49;
assign v3a6267f = hbusreq2_p & v3773ee6 | !hbusreq2_p & v3a617b4;
assign v38063dd = hgrant2_p & v3732d55 | !hgrant2_p & v377d8eb;
assign v3746fce = hbusreq1_p & v3734f9f | !hbusreq1_p & !v8455ab;
assign v3a6f53e = jx0_p & v3771431 | !jx0_p & v3a71227;
assign v377b4b9 = hgrant2_p & v37639c6 | !hgrant2_p & v3a709cf;
assign v374f832 = hbusreq7 & v1e3780d | !hbusreq7 & v8455ab;
assign v35b9d52 = stateA1_p & v376a35c | !stateA1_p & v3757c6f;
assign v3731666 = hbusreq2 & v3a63805 | !hbusreq2 & v8455ab;
assign v3737ac8 = hbusreq3_p & v3a6d1a4 | !hbusreq3_p & v37485f0;
assign v3752cc4 = hbusreq7_p & v37503ce | !hbusreq7_p & v376ab0f;
assign v3762502 = hlock0_p & v3747302 | !hlock0_p & v37276eb;
assign cb8cbb = hmaster1_p & v377e442 | !hmaster1_p & v3762100;
assign v3755451 = hgrant6_p & v3a5b89b | !hgrant6_p & v3a6488f;
assign v3758526 = hmaster1_p & v375f8f2 | !hmaster1_p & v376abdf;
assign v3770735 = hgrant2_p & v23fe159 | !hgrant2_p & v8455ab;
assign v3a56318 = hgrant6_p & v373cc95 | !hgrant6_p & v3745b15;
assign d39337 = hgrant0_p & v3a6ffb6 | !hgrant0_p & v373c428;
assign v376df24 = hbusreq0 & v3a6fb8c | !hbusreq0 & v3736db8;
assign v373483e = hbusreq5 & v8455ab | !hbusreq5 & v3a58c07;
assign v3756a05 = hmaster2_p & v8455ab | !hmaster2_p & v3774f24;
assign v377df2e = hgrant4_p & v3751f34 | !hgrant4_p & v3a709e2;
assign v3a634b9 = jx0_p & v3a70ab8 | !jx0_p & v3747897;
assign v3a2a766 = stateA1_p & v8455ab | !stateA1_p & v376e491;
assign v3732f65 = jx2_p & v37751b2 | !jx2_p & v377311c;
assign v3775709 = hlock8 & v37388f6 | !hlock8 & v3776c6e;
assign v372e88f = hlock4 & v3a6a346 | !hlock4 & v3723bac;
assign v3a57ef6 = hbusreq8 & v377a855 | !hbusreq8 & v373db25;
assign v90b307 = hgrant5_p & v372773c | !hgrant5_p & !v8455ab;
assign v2acafdd = jx0_p & v374113f | !jx0_p & !v376a74a;
assign v3763b0a = hbusreq0 & v8455ab | !hbusreq0 & v373e814;
assign v375978a = hgrant3_p & v3754227 | !hgrant3_p & v3a618b7;
assign v2925cbb = hmaster2_p & v376f4b2 | !hmaster2_p & v3765d74;
assign v3a668ec = hlock3_p & v3378fca | !hlock3_p & v8455b0;
assign v376d72e = hmaster0_p & v3a6f676 | !hmaster0_p & v372f07d;
assign v3a70f30 = hmaster1_p & v372e91a | !hmaster1_p & v3a64879;
assign v357748a = decide_p & v3a700ab | !decide_p & v3a6086a;
assign v3a705bf = hbusreq6_p & v3759032 | !hbusreq6_p & !v39a537f;
assign v375b6fe = hbusreq8_p & v3778a82 | !hbusreq8_p & !v8455ab;
assign v373c82f = hbusreq8 & v3777216 | !hbusreq8 & v8455ab;
assign v3a6f993 = hbusreq3_p & v37406d2 | !hbusreq3_p & v3753dab;
assign v3a6eef5 = hmaster2_p & v374eab4 | !hmaster2_p & v3a71016;
assign v3a705de = hlock6_p & v37625a8 | !hlock6_p & v3a5ace5;
assign v3a69fcf = hbusreq5_p & v372490a | !hbusreq5_p & !v3a70ce5;
assign v3a713f0 = hmaster2_p & v3740171 | !hmaster2_p & v3767f33;
assign v3a712a2 = hmaster2_p & v3a6f081 | !hmaster2_p & !v3730a3d;
assign v37518f0 = jx0_p & v3774372 | !jx0_p & v3a6fb0a;
assign v375604f = hgrant6_p & v374a3db | !hgrant6_p & v3a6fd47;
assign v3a59ddc = hmaster1_p & v869938 | !hmaster1_p & v38065f1;
assign v374c425 = hbusreq2_p & v3a64b41 | !hbusreq2_p & v3a6f0a9;
assign v3759ac1 = hbusreq5_p & v2093037 | !hbusreq5_p & v372601c;
assign v3a5803d = hbusreq8_p & v3a6f5ff | !hbusreq8_p & v3740f78;
assign v377c47d = stateA1_p & v3a7091d | !stateA1_p & v37324c0;
assign v3a6c580 = hbusreq2_p & v3a714bd | !hbusreq2_p & v374d479;
assign v3a5af1e = hlock6 & v3a6e21a | !hlock6 & v3755665;
assign v375cbe2 = hmaster2_p & v8455ab | !hmaster2_p & !v3773fdc;
assign v3746d92 = jx0_p & v3a70f55 | !jx0_p & v23fdbfc;
assign v374156a = hmaster0_p & v375d76b | !hmaster0_p & v8455c2;
assign v3749437 = hbusreq0 & v39eb56c | !hbusreq0 & v375c728;
assign v377e710 = hmaster3_p & v3777140 | !hmaster3_p & v373ae27;
assign v372d3e5 = hgrant2_p & v3a71164 | !hgrant2_p & v2ff8be4;
assign v37346c5 = jx2_p & v3752a05 | !jx2_p & v3a68391;
assign v3a6eecd = hbusreq3 & v377857d | !hbusreq3 & v3a635ea;
assign v3770075 = hbusreq2_p & v3746a2b | !hbusreq2_p & v3a63621;
assign v3a7003d = hbusreq8_p & v8455ab | !hbusreq8_p & v3734473;
assign v3a61f3c = hgrant2_p & v8455ab | !hgrant2_p & v3a71437;
assign v375ac70 = hbusreq2 & v375d161 | !hbusreq2 & v8455ab;
assign v374523b = hbusreq0 & v3725671 | !hbusreq0 & v375a3a8;
assign v3758adb = hgrant3_p & v374383b | !hgrant3_p & v372618d;
assign v3a6ef00 = hbusreq4 & aab2b0 | !hbusreq4 & v8455e7;
assign v3a64f1f = hmaster1_p & v8455ab | !hmaster1_p & v3a625ac;
assign v2acafac = hmaster2_p & v3a635ea | !hmaster2_p & v3745f9b;
assign v3a700e0 = hmaster2_p & v37646e1 | !hmaster2_p & v37631d9;
assign v3776b61 = hgrant0_p & v3768062 | !hgrant0_p & v3a6123e;
assign v377f397 = hbusreq6_p & v3a635ea | !hbusreq6_p & ac9d0d;
assign v373b6e4 = hgrant7_p & v377f7dd | !hgrant7_p & v37368d0;
assign v374177d = hmaster0_p & v37795d3 | !hmaster0_p & v375ff4e;
assign v3807ac3 = hlock6 & v3a57214 | !hlock6 & v3a70f43;
assign v37643b5 = hbusreq0 & v3a710aa | !hbusreq0 & v3732b1e;
assign v3a62965 = hmaster2_p & v3747302 | !hmaster2_p & v3a6f4c7;
assign v3a652a6 = hgrant2_p & v8455ab | !hgrant2_p & v3a5af82;
assign v377f2ec = hmaster0_p & v1e38260 | !hmaster0_p & v377a985;
assign v3a58674 = hgrant6_p & v3754e78 | !hgrant6_p & v3a675bc;
assign v3777763 = hmaster0_p & v373a1b4 | !hmaster0_p & v3a70a42;
assign v3740885 = hbusreq5 & v3776454 | !hbusreq5 & v3a6ff12;
assign v3770891 = jx0_p & v37617d8 | !jx0_p & v3734397;
assign v37790a6 = hbusreq5 & v372f0bc | !hbusreq5 & v3757ad8;
assign v3766df9 = hgrant3_p & v3754227 | !hgrant3_p & v373d7fe;
assign v3937409 = decide_p & v3a70945 | !decide_p & v377b221;
assign v3766b26 = hbusreq5 & v377faae | !hbusreq5 & v37357ce;
assign v3727f86 = hgrant1_p & v3732f00 | !hgrant1_p & !v8455ab;
assign v3764df7 = hgrant2_p & v375a268 | !hgrant2_p & v375da17;
assign v3a68c7d = hmaster0_p & v3748451 | !hmaster0_p & v377a577;
assign v3a71361 = hbusreq7 & v373a0e2 | !hbusreq7 & v372beb6;
assign v360d03f = hlock1 & v373dd8a | !hlock1 & v3743b9e;
assign v373eecc = hlock6 & v37559ea | !hlock6 & v374956a;
assign v3a5df87 = hlock6 & v38072fd | !hlock6 & v3734f70;
assign v360d136 = hbusreq4_p & v376e72d | !hbusreq4_p & v37252c2;
assign v3a6f56b = hmaster0_p & v372e712 | !hmaster0_p & v373f2a6;
assign v376533e = hbusreq6 & v3a6eead | !hbusreq6 & v3762502;
assign v377ca8e = hgrant6_p & v3741f22 | !hgrant6_p & v37381eb;
assign v374c5fc = hmaster0_p & v377a369 | !hmaster0_p & v1e37cc1;
assign v38088e1 = hmaster2_p & v3752cc5 | !hmaster2_p & v3a54497;
assign v3752767 = hgrant6_p & v3a6f43a | !hgrant6_p & v3806f19;
assign v3770415 = hbusreq2_p & v377bdb8 | !hbusreq2_p & v8455ab;
assign v3764f39 = hgrant5_p & v375ed60 | !hgrant5_p & v374a849;
assign v372c9b0 = hmaster2_p & v3753dab | !hmaster2_p & v3732c51;
assign v3722e5c = locked_p & v35772a5 | !locked_p & v35772a6;
assign v37430c6 = hlock2_p & v3755002 | !hlock2_p & !v8455ab;
assign v3a70a42 = hmaster2_p & v373a1b4 | !hmaster2_p & !v8455ab;
assign v37332dd = hbusreq2 & v372df9a | !hbusreq2 & v377957e;
assign v3a6bb47 = hbusreq7 & v377d428 | !hbusreq7 & v3743a4c;
assign v3a6f13e = hmaster2_p & v8455ab | !hmaster2_p & v3a6fd91;
assign v3771ae3 = hburst1 & v373d9e5 | !hburst1 & v3a703d1;
assign v373642c = hbusreq6 & v8455e7 | !hbusreq6 & v8455ab;
assign v376583c = hmaster0_p & v3771fb7 | !hmaster0_p & v3a7004b;
assign v37337f1 = hbusreq5 & v3779aa8 | !hbusreq5 & !v3a5398c;
assign v376af8c = hlock5_p & v372750b | !hlock5_p & v3a701f2;
assign v3a5a72a = hbusreq4 & v3747042 | !hbusreq4 & v8455ab;
assign v373681a = hbusreq2_p & v376f5ef | !hbusreq2_p & !v8455ab;
assign v3759570 = hgrant0_p & v8455ab | !hgrant0_p & v375e459;
assign v374ad81 = hbusreq6_p & v3a70ee7 | !hbusreq6_p & v3733d6e;
assign v3733fad = hbusreq4 & v3723614 | !hbusreq4 & v3763104;
assign v3a6f95b = hbusreq7 & v3a711c8 | !hbusreq7 & v373fe8f;
assign v374ccb7 = hburst1 & v37295fe | !hburst1 & v325b5ea;
assign v3a6f049 = hlock7_p & v3a6ddb3 | !hlock7_p & !v3a6146c;
assign v928541 = hlock0 & v373abde | !hlock0 & v377723a;
assign v3738397 = hgrant0_p & v23fe0bb | !hgrant0_p & v3761cec;
assign v373f224 = hbusreq6_p & v39eb536 | !hbusreq6_p & v8455ab;
assign v372cfeb = hbusreq6_p & v376110e | !hbusreq6_p & v3a637dd;
assign v3a707c4 = hbusreq1_p & v37585e6 | !hbusreq1_p & !v8455ab;
assign v377cf34 = hmaster1_p & v3a635ea | !hmaster1_p & v3743a8a;
assign v37511f6 = jx0_p & v3767e38 | !jx0_p & v3745f63;
assign v3737d38 = hbusreq6_p & v37367f1 | !hbusreq6_p & v8455ab;
assign v3759232 = hbusreq8 & v3a6ebfc | !hbusreq8 & v374757c;
assign v37247b5 = hmaster0_p & v3734c5c | !hmaster0_p & v3a6fa45;
assign v373c617 = hbusreq8 & v380909f | !hbusreq8 & v3779f1e;
assign v3a61c70 = hmaster2_p & v376d285 | !hmaster2_p & v3758166;
assign v38087c5 = hgrant4_p & v3a70104 | !hgrant4_p & v3a56688;
assign v3729b4c = hbusreq4_p & v3a58907 | !hbusreq4_p & v3a6ebf2;
assign v375a59f = hbusreq7_p & v375b15b | !hbusreq7_p & v8455ab;
assign v3a63bd4 = hmaster0_p & v37430c6 | !hmaster0_p & v3751d6f;
assign v3728c08 = hgrant4_p & v8455ab | !hgrant4_p & v37771ca;
assign v376c30b = hmaster0_p & v8455ab | !hmaster0_p & v37764f7;
assign v3a5f02e = hgrant4_p & v376a6f1 | !hgrant4_p & v372cac5;
assign v3a7113a = hbusreq0 & v3a712c5 | !hbusreq0 & v8455ab;
assign v3a639a1 = hgrant5_p & v375afbf | !hgrant5_p & v3a7047b;
assign v377b2b6 = hbusreq6 & v3733c46 | !hbusreq6 & v8455ab;
assign v3a6d1fa = hlock0 & v3730695 | !hlock0 & v3742723;
assign v3a70bf2 = hgrant4_p & v8455ab | !hgrant4_p & v3a55785;
assign v374c34d = hbusreq5_p & v377abe1 | !hbusreq5_p & v3a7143d;
assign v38070ea = hmaster0_p & v3a700b2 | !hmaster0_p & v3a6eae9;
assign v3735d01 = hlock7 & v3a63f80 | !hlock7 & v3a70bfb;
assign v3a6eb7f = hmaster1_p & v3759cc1 | !hmaster1_p & v8455ab;
assign v374476d = hmaster2_p & v373abdd | !hmaster2_p & v373e1d0;
assign v3a6eaf3 = hbusreq4_p & v3a7139c | !hbusreq4_p & aca44a;
assign v37251f6 = hbusreq3_p & v3733ba1 | !hbusreq3_p & v37366d2;
assign v3779852 = hmaster1_p & v37524cf | !hmaster1_p & v3a60e4c;
assign v3749091 = hbusreq5_p & v3a70675 | !hbusreq5_p & v23fd7e1;
assign v3a568ac = hgrant1_p & v3a637dc | !hgrant1_p & v3a7048a;
assign v37647de = hgrant5_p & v37244f1 | !hgrant5_p & !v3a6f796;
assign v37290af = hlock2_p & v377b8ee | !hlock2_p & !v8455ab;
assign v377d99d = hbusreq3 & v3748ca3 | !hbusreq3 & v373006f;
assign v3a6fc50 = hmaster0_p & v3a63de8 | !hmaster0_p & d95e20;
assign v3745202 = hmaster0_p & v3a63777 | !hmaster0_p & v3a60649;
assign v373a188 = hbusreq2 & v3a6f993 | !hbusreq2 & v8455ab;
assign v3a61988 = stateG2_p & v8455ab | !stateG2_p & !v376f693;
assign v1e37762 = hgrant6_p & v8455ab | !hgrant6_p & v373f1e4;
assign v374e5ab = hbusreq7 & v33782fe | !hbusreq7 & !v8455ca;
assign v372fff3 = hbusreq4 & v3731eff | !hbusreq4 & v37775f9;
assign v3746259 = hbusreq0 & v374c0e4 | !hbusreq0 & v3770eb9;
assign v3a66d7b = hgrant3_p & v8455ab | !hgrant3_p & v37714e6;
assign v3a6a393 = hgrant3_p & v3a70a88 | !hgrant3_p & v3726006;
assign v3741280 = hmaster0_p & v374bf07 | !hmaster0_p & v3a6fcab;
assign v3a615bb = hlock2 & v38072fd | !hlock2 & v377b27b;
assign v374d612 = hmaster1_p & v3a635ea | !hmaster1_p & cbfab3;
assign v3760317 = hmaster3_p & v3776311 | !hmaster3_p & !v376b1ee;
assign v3a629fb = jx1_p & v376079a | !jx1_p & v3a69957;
assign v3761719 = hgrant4_p & v8455ab | !hgrant4_p & v375ce35;
assign v372d866 = hmaster2_p & v377c6b3 | !hmaster2_p & v376e90a;
assign v372fdfd = hmaster1_p & v373fd7b | !hmaster1_p & v373e055;
assign v3a5ac38 = hmaster2_p & v38073be | !hmaster2_p & v374686d;
assign v3577318 = hbusreq5_p & v9fc6a0 | !hbusreq5_p & v3a6498e;
assign v375b03c = hmaster1_p & v3769a71 | !hmaster1_p & v37638ef;
assign v3767a7b = hbusreq3 & v39a4e5f | !hbusreq3 & v37317a9;
assign v3739368 = hbusreq7 & v3a561f0 | !hbusreq7 & v37670dd;
assign v373cd8f = hmaster2_p & v3a58cfc | !hmaster2_p & !v3a5bf04;
assign v3a67cff = hbusreq6_p & v3747302 | !hbusreq6_p & v37496fa;
assign v3766852 = hbusreq8 & v372a4e5 | !hbusreq8 & v3773536;
assign v3a7137f = hlock0 & v374f35a | !hlock0 & v3a5c25e;
assign v376a88b = hbusreq6_p & v376b600 | !hbusreq6_p & !v3a5bf04;
assign v3742005 = hmaster1_p & v8455ab | !hmaster1_p & v3a710de;
assign v3a62caa = hbusreq0 & v375a38e | !hbusreq0 & v37600e9;
assign v3a704d1 = hmaster1_p & v373ad69 | !hmaster1_p & v375ac12;
assign v3a6f4ef = hgrant2_p & v375e7cc | !hgrant2_p & v3a5bb98;
assign v377e545 = hgrant2_p & v3774c1b | !hgrant2_p & v3a6f6f4;
assign v3777d7c = hmaster0_p & v3a6953d | !hmaster0_p & !v3a70386;
assign b5da28 = hmaster0_p & v377e31b | !hmaster0_p & v373a822;
assign v3809a6a = hgrant4_p & v8455ab | !hgrant4_p & v374d859;
assign v3a5e686 = hgrant3_p & v3752a0d | !hgrant3_p & v3745dac;
assign v3a70317 = hbusreq4 & v377a1d3 | !hbusreq4 & v374d0f9;
assign d950cb = hbusreq8 & v37629fc | !hbusreq8 & v3734279;
assign v3750f4c = hmaster2_p & v375bb51 | !hmaster2_p & v3a6eb7b;
assign v3a67471 = hmaster0_p & v3754f93 | !hmaster0_p & v8455e7;
assign v3807107 = hgrant0_p & v8455e7 | !hgrant0_p & v373e67e;
assign v375fe83 = hlock5 & v372def9 | !hlock5 & v3a7102f;
assign v3807c0c = hlock0_p & v3806507 | !hlock0_p & v3a70cd2;
assign v3768dd8 = hmaster0_p & v3765265 | !hmaster0_p & v3a5fde5;
assign v372b3ca = hbusreq5_p & v374bc9c | !hbusreq5_p & v3767e79;
assign v372ff75 = hbusreq7_p & v1e38301 | !hbusreq7_p & v3a5e19b;
assign v3a6015c = hlock5 & v3a59085 | !hlock5 & v3727c07;
assign v374b6ba = hbusreq4_p & v373a303 | !hbusreq4_p & v372d19a;
assign v37697f0 = hbusreq5_p & v37349f9 | !hbusreq5_p & v375b0ad;
assign bee241 = hgrant2_p & v8455ab | !hgrant2_p & v3773137;
assign v3a70bc4 = hbusreq7 & v376543b | !hbusreq7 & v3a5f218;
assign v373ab12 = hlock4_p & v373ad95 | !hlock4_p & v8455ab;
assign v37700b9 = hbusreq2 & v3749907 | !hbusreq2 & v8455ab;
assign v373d4fc = hgrant2_p & v8455ab | !hgrant2_p & v3752e71;
assign v3a5f67d = hbusreq2_p & v8455bf | !hbusreq2_p & v3770b6e;
assign v3773098 = hmaster1_p & v3a6614b | !hmaster1_p & v3777527;
assign v9b03cc = hbusreq0 & v37672c8 | !hbusreq0 & v375115e;
assign v3773f70 = hbusreq8_p & v3746acf | !hbusreq8_p & v3a7090b;
assign v37502f1 = hmaster0_p & v374074a | !hmaster0_p & v3774438;
assign v37738ca = hbusreq5 & v374153d | !hbusreq5 & v8455ab;
assign v3733be0 = hlock0_p & v3a5f8d0 | !hlock0_p & v3a63805;
assign v3725be8 = hmaster3_p & v3765962 | !hmaster3_p & v374bb74;
assign v3a6f77b = hgrant7_p & v3a58792 | !hgrant7_p & v3a6bb4b;
assign v37781d4 = hbusreq5 & v372c6c4 | !hbusreq5 & v373ab06;
assign v377e57f = hbusreq4_p & v3a6f043 | !hbusreq4_p & v3a5db41;
assign v3726bff = hbusreq6_p & ca1199 | !hbusreq6_p & !v3a6fdae;
assign v3733da3 = hgrant3_p & v3a64f9b | !hgrant3_p & v3a6f748;
assign v3a65a2e = jx1_p & v373c0a8 | !jx1_p & v376a70f;
assign v375d6b4 = hmaster2_p & v37737aa | !hmaster2_p & b66167;
assign v3a7160f = hgrant4_p & v372b77b | !hgrant4_p & v377b0a0;
assign v3a6df51 = hbusreq7_p & v377113b | !hbusreq7_p & v37263d2;
assign v374f359 = hmaster0_p & v3740953 | !hmaster0_p & v3a59bbd;
assign v3733f1c = hbusreq2 & v37693cf | !hbusreq2 & v8455ab;
assign v373d5f0 = hbusreq5_p & v3742649 | !hbusreq5_p & v37bfc97;
assign v3a6ff10 = hlock0 & v374165f | !hlock0 & v377150c;
assign v375d849 = hgrant5_p & v3807b27 | !hgrant5_p & v3772a4f;
assign v35b776e = hbusreq8 & v3766048 | !hbusreq8 & v377435f;
assign v3751253 = hmaster2_p & v3777311 | !hmaster2_p & v377961f;
assign v3a53f00 = hbusreq6_p & v38093aa | !hbusreq6_p & v37786bb;
assign v3738910 = hgrant2_p & v8455ab | !hgrant2_p & v37452d5;
assign v3a7093f = hmaster1_p & v3a6f224 | !hmaster1_p & v3778c14;
assign v3a5520a = hmaster0_p & v3723211 | !hmaster0_p & v374f820;
assign v376a94b = hbusreq8 & v3a55bfa | !hbusreq8 & v3737808;
assign v380949b = hbusreq4_p & v37632f8 | !hbusreq4_p & !v3737860;
assign v39ea0c2 = hbusreq5 & v3767a85 | !hbusreq5 & v3a6c09f;
assign v3750ce8 = hgrant6_p & v8455ab | !hgrant6_p & v372eaf3;
assign v3731dc1 = hmaster0_p & v374f857 | !hmaster0_p & v372a696;
assign v3a62f59 = hgrant7_p & v3768b2d | !hgrant7_p & v375fb86;
assign v3a64da2 = hmaster1_p & v3742dfb | !hmaster1_p & v3a6eec3;
assign v3744e62 = hgrant5_p & v37408e4 | !hgrant5_p & v377312b;
assign v375dbc6 = hgrant1_p & v3a7069e | !hgrant1_p & !v3a6e9b1;
assign v376646a = hlock6 & v375fbb7 | !hlock6 & v37616e0;
assign v37750c2 = hgrant6_p & v8455ab | !hgrant6_p & v3750b85;
assign v3768fc7 = hmaster2_p & v37674c1 | !hmaster2_p & v8455ab;
assign v375473a = hgrant6_p & v373f0a3 | !hgrant6_p & v8455ab;
assign v3744410 = hbusreq8 & v372cb2c | !hbusreq8 & v8455ab;
assign v373264f = hmaster1_p & v3777d7c | !hmaster1_p & v8455ca;
assign v376d2b7 = hbusreq4_p & v3759837 | !hbusreq4_p & v3740348;
assign v37481bf = hmaster2_p & v3728685 | !hmaster2_p & v3a6f2d9;
assign v397fb7c = hmaster1_p & v3743efa | !hmaster1_p & v39eb519;
assign v373ad86 = hmaster0_p & v3a6e31f | !hmaster0_p & v3730876;
assign v372ff68 = hbusreq0 & v37721e3 | !hbusreq0 & v372594c;
assign v3730043 = hlock4 & v1e379ef | !hlock4 & v3a6f567;
assign v375b752 = hbusreq8_p & v375a71d | !hbusreq8_p & v37258d0;
assign v3722bfc = hmaster1_p & v3a5a01b | !hmaster1_p & v373676d;
assign v3a6fb42 = hbusreq7_p & v37723ed | !hbusreq7_p & !v374dba6;
assign v3740fc3 = hbusreq5 & v376f07c | !hbusreq5 & v8455ab;
assign v3a5f495 = hmaster2_p & v3a63dbb | !hmaster2_p & v3734af2;
assign v373824d = hgrant5_p & v8455ab | !hgrant5_p & v376296b;
assign v372eab1 = hbusreq4_p & v3737d38 | !hbusreq4_p & v3a6efc8;
assign dc47a7 = hmaster2_p & v3a5fc34 | !hmaster2_p & v3a63a7a;
assign v374bb16 = hbusreq8 & v3742a4d | !hbusreq8 & v3a6fba3;
assign v3a6f94e = hbusreq4_p & v375da9d | !hbusreq4_p & v372ff68;
assign v3a6fb65 = hmaster2_p & v376926f | !hmaster2_p & v3755b56;
assign v3722a9c = hgrant4_p & v3739896 | !hgrant4_p & v373f10d;
assign v3a71459 = hmaster0_p & v3759279 | !hmaster0_p & !v372362a;
assign v337902c = hmaster2_p & v3743f3c | !hmaster2_p & v3a69946;
assign v3773697 = hbusreq5_p & v3765f99 | !hbusreq5_p & v8455cb;
assign v3a7045f = hlock0 & v3731230 | !hlock0 & v3a71600;
assign v373aa91 = hmaster0_p & v3738a2b | !hmaster0_p & v3747bfe;
assign v3a70d3d = hmaster1_p & v3a70856 | !hmaster1_p & v37697f0;
assign v3a6ffb1 = jx1_p & v3a5e65e | !jx1_p & v3a6f407;
assign v374aa71 = hgrant4_p & v376ea4a | !hgrant4_p & v3a63d3c;
assign b2271d = hbusreq6 & v375cdd7 | !hbusreq6 & v8455ab;
assign v37614fa = hlock8_p & v3a5d8e8 | !hlock8_p & v990999;
assign v3744f1e = jx1_p & v374b228 | !jx1_p & v3a68f22;
assign v3a6935c = hgrant4_p & v8455ab | !hgrant4_p & aba148;
assign v3a581f1 = hmaster1_p & v3726eea | !hmaster1_p & v377a571;
assign v373580c = hmaster1_p & v1e382e7 | !hmaster1_p & v3a7115d;
assign v8c9ea7 = hgrant5_p & v3748c75 | !hgrant5_p & v376f9d3;
assign v3a57750 = hlock0 & v3809ec3 | !hlock0 & v374fc57;
assign v360d140 = hmaster0_p & v37480b7 | !hmaster0_p & v3a702da;
assign v376654b = hmaster2_p & v35b9d52 | !hmaster2_p & v8455ab;
assign v376d6d9 = hgrant5_p & v8455e7 | !hgrant5_p & v3a6f225;
assign v3a70cd5 = stateA1_p & v8455ab | !stateA1_p & !v3745b85;
assign v3a6fc6c = hgrant1_p & v377eaf2 | !hgrant1_p & v8455ab;
assign v375144b = hgrant4_p & v3a6d809 | !hgrant4_p & v3a67ee6;
assign v3a6f539 = hlock3_p & v374c2b4 | !hlock3_p & !v8455be;
assign v3a54bcd = stateG10_1_p & v8455b0 | !stateG10_1_p & !v377ed8c;
assign v3a70fa3 = hbusreq5_p & v380a170 | !hbusreq5_p & v3778aa6;
assign v3a710ae = hgrant5_p & v3730019 | !hgrant5_p & v3737c88;
assign v3a59351 = hgrant0_p & v8455ab | !hgrant0_p & v39eaa47;
assign v3a6b4f6 = hgrant0_p & v8455ab | !hgrant0_p & v3a6fd57;
assign v375b787 = hbusreq5 & v3a61de8 | !hbusreq5 & v3765cd5;
assign v376f321 = hmaster0_p & v3a5fc34 | !hmaster0_p & v3730e43;
assign v375aa0d = hlock5_p & v3a711a8 | !hlock5_p & v8455ab;
assign v3a54b31 = hmaster2_p & v8455ab | !hmaster2_p & v3723b00;
assign v37677ee = hgrant3_p & v8455b0 | !hgrant3_p & v3743e56;
assign v376755f = hmaster1_p & v3745e51 | !hmaster1_p & v3758ee1;
assign v3a62b09 = hbusreq5 & v3a5a2c6 | !hbusreq5 & v3a5bf21;
assign v375e1de = hmaster1_p & v373014d | !hmaster1_p & v3a5732f;
assign v39a4f35 = decide_p & v375c6d6 | !decide_p & v37330d6;
assign v8455d3 = hlock8_p & v8455ab | !hlock8_p & !v8455ab;
assign v3730d34 = hlock0 & v3a70a7f | !hlock0 & v3759f23;
assign v37342f2 = hgrant4_p & v8455ab | !hgrant4_p & v3738491;
assign v3a70212 = hbusreq0 & v373e21a | !hbusreq0 & !v372e30c;
assign v37574f8 = hlock0_p & v3769ae2 | !hlock0_p & v373453a;
assign v37248fd = hgrant4_p & v3747ac9 | !hgrant4_p & v3a56d2d;
assign v376c6fb = hmaster0_p & v3a715b7 | !hmaster0_p & v372dcf7;
assign v37c3782 = hbusreq0 & v3a70e77 | !hbusreq0 & v37508c2;
assign v3a70a55 = hbusreq2_p & v3a6fa15 | !hbusreq2_p & v8455ab;
assign v377af89 = hmaster1_p & v3776864 | !hmaster1_p & v373f27d;
assign v3a71411 = hbusreq6_p & v3a2978d | !hbusreq6_p & v3a53f2b;
assign v3807a8d = hgrant6_p & v3a6f61e | !hgrant6_p & !v372b795;
assign v3a5b20c = hmaster0_p & v37432cd | !hmaster0_p & v3a5e7c4;
assign v3766792 = hmaster0_p & v37652d4 | !hmaster0_p & v3a70c2c;
assign v3a66161 = hmaster0_p & v3a707d0 | !hmaster0_p & v37527dc;
assign v3749fd7 = hbusreq4 & v3a58f20 | !hbusreq4 & v8455ab;
assign v3730060 = hmaster2_p & v377bf71 | !hmaster2_p & v374355e;
assign v3a6995c = hbusreq0 & v3723e64 | !hbusreq0 & v3736a23;
assign v3743613 = hmaster0_p & v3a6f5c8 | !hmaster0_p & v379318b;
assign v3a6ef63 = hgrant5_p & v8455ab | !hgrant5_p & v375e320;
assign v375c044 = hmaster2_p & v8455ab | !hmaster2_p & v37609ab;
assign v39eb033 = hlock5_p & v377c7c0 | !hlock5_p & v373014d;
assign v376e65d = hbusreq0 & v3749e5a | !hbusreq0 & v374edff;
assign v3738d86 = hbusreq7_p & v37497a5 | !hbusreq7_p & v3a5c65d;
assign v376a877 = hgrant6_p & v377f09a | !hgrant6_p & v936e47;
assign v3a7145f = hgrant2_p & v3a646f5 | !hgrant2_p & v37316b7;
assign v3a70932 = hbusreq5 & v374801c | !hbusreq5 & v8455bb;
assign v3a70386 = hmaster2_p & v8455ab | !hmaster2_p & !v8455ca;
assign v3a6ef74 = hgrant3_p & v377dd3b | !hgrant3_p & v37509c7;
assign v3a5d830 = hgrant6_p & v3723012 | !hgrant6_p & v8455ab;
assign v3a6fad6 = hmaster2_p & v3778e28 | !hmaster2_p & !v23fe339;
assign v3a716a6 = hlock4_p & v8455ab | !hlock4_p & !v3753f1a;
assign v3a70d23 = hmaster1_p & v37560c9 | !hmaster1_p & v3727387;
assign v377d69c = hgrant4_p & v3a70bd6 | !hgrant4_p & v375ea89;
assign v992750 = hmaster1_p & v3769ae2 | !hmaster1_p & v37505a2;
assign v3a6dc91 = hmaster0_p & v3a5bbc2 | !hmaster0_p & v37520ad;
assign v3a6909a = hbusreq4_p & v373fe5e | !hbusreq4_p & v8455e7;
assign v3a60134 = hlock7 & v37758de | !hlock7 & v3776066;
assign v374b4ef = hmaster0_p & v3a5c5e5 | !hmaster0_p & v3757966;
assign v3a700a8 = hmaster2_p & v3773c36 | !hmaster2_p & v3760c3c;
assign v3a6ebac = hmaster2_p & v3a6a2f3 | !hmaster2_p & v3a667e7;
assign v37532a6 = hgrant2_p & v8455ab | !hgrant2_p & !v373c853;
assign v374055c = hmaster0_p & v3a5c945 | !hmaster0_p & v3808e82;
assign v377dd3b = hbusreq3_p & v3a674ac | !hbusreq3_p & !v8455ab;
assign v37493b9 = hbusreq2_p & v3740f70 | !hbusreq2_p & v3767cd6;
assign v3731678 = hlock0_p & v375e657 | !hlock0_p & v3a5fdab;
assign v3a5c80e = hgrant6_p & v3807f45 | !hgrant6_p & v3a5ff5a;
assign v375f938 = hmaster1_p & v374db8d | !hmaster1_p & v3a70ba1;
assign v37281ca = hmaster0_p & v3772c5a | !hmaster0_p & v3729004;
assign v3740247 = hbusreq8 & v373f909 | !hbusreq8 & v376e66e;
assign v375c4f9 = hmaster0_p & v37483ff | !hmaster0_p & v3a665d5;
assign v373d8c0 = stateG10_1_p & v90a00a | !stateG10_1_p & !v3a714e6;
assign v373c924 = hgrant3_p & v8455ab | !hgrant3_p & v376a6d7;
assign v37300a5 = hbusreq4_p & v374d6dd | !hbusreq4_p & v37759b6;
assign v3a61038 = hmaster0_p & v372ba1c | !hmaster0_p & v373cfbd;
assign v372bcd3 = hbusreq5 & v37713e8 | !hbusreq5 & v3a70f0d;
assign v3a71304 = hbusreq6_p & v3a62d18 | !hbusreq6_p & !v3a672c9;
assign v3728ea6 = hlock1 & v375483e | !hlock1 & v3778528;
assign v3a66a4f = jx0_p & v3a61132 | !jx0_p & v3a6f625;
assign v376e532 = hlock4_p & v3a707b7 | !hlock4_p & v373127e;
assign v3a70a88 = hlock0_p & v37496fa | !hlock0_p & v3a706df;
assign v376a7da = hmaster1_p & v375c6c1 | !hmaster1_p & v2acb110;
assign v37559ec = hmaster2_p & v3a53dbb | !hmaster2_p & v3768889;
assign v3a66e4c = hbusreq6_p & v3a67729 | !hbusreq6_p & v375fe5b;
assign v372c03b = hmaster2_p & v8455b0 | !hmaster2_p & v3a63659;
assign v3a70b76 = hbusreq6 & v37554c0 | !hbusreq6 & v23fd967;
assign v3a6810b = hmaster0_p & v377e897 | !hmaster0_p & v8455e7;
assign v3a6b297 = hlock0_p & v3a6f316 | !hlock0_p & v377bf0d;
assign v37652a5 = hlock0_p & v8455ab | !hlock0_p & v3a6ab5f;
assign v3765e47 = hmaster1_p & v8455ab | !hmaster1_p & v3a7122f;
assign v3a6f45c = hmaster0_p & v37610e5 | !hmaster0_p & v3759584;
assign v377adf5 = hbusreq2_p & v3807bf8 | !hbusreq2_p & v3a66110;
assign v37366b5 = hgrant3_p & v3a5b6de | !hgrant3_p & v3749629;
assign v3a7140f = hmaster0_p & v3a6fa69 | !hmaster0_p & v3a6fb52;
assign v37418ab = hmaster1_p & v374f307 | !hmaster1_p & v377f579;
assign v372f739 = hmaster1_p & v377b626 | !hmaster1_p & v375da6a;
assign v2092be1 = hbusreq4_p & v3726d1f | !hbusreq4_p & v372b847;
assign v3749f49 = hmaster3_p & v3a69203 | !hmaster3_p & v3a7168c;
assign v3a5f2bd = hlock5_p & v372ab0f | !hlock5_p & v3a678de;
assign v3754aa3 = hbusreq3_p & v3756465 | !hbusreq3_p & !v8455ab;
assign v3779f92 = hmaster1_p & v8455c2 | !hmaster1_p & v374b497;
assign v37390ed = hgrant0_p & v8455e7 | !hgrant0_p & !v376f178;
assign v37721e6 = hlock1_p & v3a70010 | !hlock1_p & !v8455ab;
assign v3724a1c = hbusreq2_p & v374fd8d | !hbusreq2_p & v8455ab;
assign v3776d42 = hmaster1_p & v3a70557 | !hmaster1_p & v3a70adb;
assign v3767b62 = hmaster0_p & v374006f | !hmaster0_p & v3740e4c;
assign v3a6ff74 = hlock4_p & v372a00b | !hlock4_p & v3a6fb2b;
assign v23fd89c = hbusreq5_p & v3731aaf | !hbusreq5_p & v3756737;
assign v3a69390 = hbusreq5_p & v3765f99 | !hbusreq5_p & v374c3ff;
assign v374888e = hbusreq7_p & v3a5f714 | !hbusreq7_p & !v3749ed5;
assign v377b456 = hbusreq5_p & v37725d6 | !hbusreq5_p & v8455ab;
assign v373c4a7 = hmaster1_p & v8455ab | !hmaster1_p & v3739914;
assign v37709d2 = hbusreq2_p & v376dbdf | !hbusreq2_p & !v372fc81;
assign v3751c87 = hbusreq1_p & v8455e7 | !hbusreq1_p & !v3752648;
assign v3764d3e = hmaster1_p & v37294a9 | !hmaster1_p & v375652a;
assign v33790e4 = hbusreq6_p & v37535e7 | !hbusreq6_p & v3a6f7a0;
assign v374fe7b = hbusreq2_p & v3a635ea | !hbusreq2_p & v377d41d;
assign v375bc5b = hgrant3_p & v3754e5a | !hgrant3_p & v3730693;
assign v3737a76 = hlock4_p & v3726077 | !hlock4_p & v8455ab;
assign v375a4fa = hbusreq2_p & v39a537f | !hbusreq2_p & !v39a5381;
assign v373c8bb = hgrant5_p & v3774063 | !hgrant5_p & v376d3e2;
assign v3a6b18a = hbusreq1_p & v372456f | !hbusreq1_p & v374a63c;
assign v375e948 = hgrant2_p & v377e867 | !hgrant2_p & v373e369;
assign v3766ed8 = hmaster1_p & v3a6b60d | !hmaster1_p & v3774b16;
assign v377dd0d = hbusreq5_p & v3a708f7 | !hbusreq5_p & v8455ab;
assign v3761727 = hbusreq7_p & v8455b7 | !hbusreq7_p & v3a710cc;
assign v374b522 = hmaster2_p & v3757966 | !hmaster2_p & v3760453;
assign v3728333 = hmaster1_p & v8455ab | !hmaster1_p & v3a55672;
assign v3a70443 = hlock6_p & v37439ad | !hlock6_p & v3a6f744;
assign v3738d63 = hlock0_p & v3a7162d | !hlock0_p & v37457c1;
assign c7ba89 = hmaster0_p & v37261b3 | !hmaster0_p & v3770fb7;
assign v3758e73 = hmaster1_p & v8455ab | !hmaster1_p & v3a715d7;
assign v37539bc = hgrant6_p & v3765474 | !hgrant6_p & v3741f3c;
assign v377fbeb = hbusreq7 & v3a64dbb | !hbusreq7 & v37305e3;
assign v39ebb5d = hbusreq7_p & v374b7ea | !hbusreq7_p & v372fb53;
assign v376e2fb = hbusreq5 & v372e031 | !hbusreq5 & v3768828;
assign v3740922 = hbusreq7 & v3a6094a | !hbusreq7 & v3a67312;
assign v3a6bfb5 = jx0_p & v3739808 | !jx0_p & v3727194;
assign v37606f0 = hmaster2_p & v37453d7 | !hmaster2_p & v8455ab;
assign v3a70533 = hbusreq8_p & v37751bb | !hbusreq8_p & v3734579;
assign v3759501 = hbusreq5_p & v374326f | !hbusreq5_p & v8455cb;
assign v3755bb4 = hmaster1_p & v374c522 | !hmaster1_p & v3747271;
assign v376c902 = hbusreq4_p & v2ff9190 | !hbusreq4_p & v39a53f3;
assign v3765b28 = hlock2_p & v3a5fa25 | !hlock2_p & v3723747;
assign v376fa3e = hmaster2_p & v3a567ec | !hmaster2_p & v3771d4f;
assign v3755c3f = hmaster1_p & v3a6f9d3 | !hmaster1_p & v3a6b78f;
assign v3772140 = hmaster0_p & v3a58218 | !hmaster0_p & v3773a25;
assign v3a5c687 = hmaster1_p & v8455ab | !hmaster1_p & v376d9f8;
assign v372d685 = hgrant7_p & v8455ce | !hgrant7_p & v374158f;
assign v8a7f7e = hbusreq1_p & v3a5c5ae | !hbusreq1_p & !v37606c7;
assign v3a6f9ae = hgrant4_p & v8455ab | !hgrant4_p & v373ea10;
assign v373b3fb = hready & v3726dfa | !hready & !v372f694;
assign v35b7044 = hgrant6_p & v37381bb | !hgrant6_p & !v3a70ece;
assign v3a640fd = hbusreq5_p & v3378992 | !hbusreq5_p & !v373644e;
assign v377714d = hlock0_p & b0c091 | !hlock0_p & !v3744710;
assign v373243e = hbusreq2_p & v37693cf | !hbusreq2_p & v3743698;
assign v377e2f7 = hgrant2_p & v3a6ceb7 | !hgrant2_p & !v3a64b41;
assign v3a6f234 = hmaster1_p & v3768e52 | !hmaster1_p & !v3a70924;
assign v3748b2c = hmaster0_p & v374502e | !hmaster0_p & v374328c;
assign v3736969 = hmaster2_p & v3a70b17 | !hmaster2_p & v3a5cfac;
assign v3769806 = hbusreq3_p & v3a70bd0 | !hbusreq3_p & v3a5cd20;
assign v3a6546f = hgrant6_p & v3a6f2d4 | !hgrant6_p & v375a579;
assign v375ec1d = hbusreq7 & v37313a7 | !hbusreq7 & v8455ab;
assign v3a6f1b9 = hmaster1_p & v39a4e99 | !hmaster1_p & v3757a04;
assign v3731be6 = hbusreq2 & v376b21a | !hbusreq2 & !v8455ab;
assign v3a57fa3 = hmaster1_p & v3809439 | !hmaster1_p & v3a590d1;
assign v3a6b4ae = hbusreq1_p & v3a5e3d3 | !hbusreq1_p & v3745801;
assign v37252ee = hlock5_p & v3a5a01b | !hlock5_p & v374e402;
assign v3a71245 = hmaster0_p & v3a70103 | !hmaster0_p & v8455e7;
assign v3771e8d = hlock2 & v3742cfe | !hlock2 & v3a712b6;
assign v3724a15 = hbusreq8_p & v3a70c57 | !hbusreq8_p & v3a709cb;
assign v374d7ce = hgrant3_p & v3768726 | !hgrant3_p & v3a71402;
assign v37286bb = hgrant1_p & v3a626a1 | !hgrant1_p & v3751fa8;
assign v3a299f3 = hmaster1_p & v3750375 | !hmaster1_p & v374975c;
assign v372e93d = hbusreq1 & v3a676d6 | !hbusreq1 & v8455ab;
assign v3a70182 = hbusreq3 & v3a619c0 | !hbusreq3 & !v8455ab;
assign v23fd9af = hbusreq7_p & v372641e | !hbusreq7_p & v3a54952;
assign v3a70b83 = hgrant6_p & v8455ca | !hgrant6_p & v37451f8;
assign v3a5c4e1 = hbusreq5 & v3a70149 | !hbusreq5 & v8455ab;
assign v3a6eebd = hmaster2_p & v3a70a88 | !hmaster2_p & v3735525;
assign v373ae02 = hmaster1_p & v373d27f | !hmaster1_p & bf5753;
assign v376ea51 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3a70a7f;
assign v37432e1 = hgrant8_p & v3748c4c | !hgrant8_p & v3730097;
assign v372e94f = hmaster2_p & v3a6fa93 | !hmaster2_p & v373698e;
assign v3a66819 = hbusreq7_p & v375070a | !hbusreq7_p & v3741c39;
assign v3a6ecee = hmaster3_p & v3a70ae5 | !hmaster3_p & v3774131;
assign v3744dc6 = hbusreq6_p & v3725786 | !hbusreq6_p & v3a70257;
assign v377435f = hgrant5_p & v8455ab | !hgrant5_p & v3741c3d;
assign v377d74d = hbusreq0_p & v376f73c | !hbusreq0_p & v376ea4a;
assign v3776516 = hlock0 & v3a5741c | !hlock0 & v372fecf;
assign v2ff9190 = hmastlock_p & v3a6eb2e | !hmastlock_p & v8455ab;
assign v374e1f6 = hbusreq5_p & v3760b46 | !hbusreq5_p & v3a58c07;
assign c1a4f5 = hbusreq1_p & v3762453 | !hbusreq1_p & v375a7bd;
assign v376bad8 = hbusreq3 & v3731258 | !hbusreq3 & v37359d8;
assign v3a6da8a = hbusreq2_p & v8455bf | !hbusreq2_p & v375c1d1;
assign v3726c61 = hgrant4_p & v3a6e31f | !hgrant4_p & v3a5fae3;
assign v3a6f130 = hgrant4_p & v1e37b99 | !hgrant4_p & !v3a5af5c;
assign v37444b4 = hbusreq4_p & v3779734 | !hbusreq4_p & v3a67f60;
assign v3727943 = hbusreq0 & v375370a | !hbusreq0 & v3a5e909;
assign v8455db = hmaster1_p & v8455ab | !hmaster1_p & !v8455ab;
assign v3a637dd = stateA1_p & v8455e1 | !stateA1_p & !v8455ab;
assign v372a1f6 = hgrant5_p & v8455ab | !hgrant5_p & !v374b6ee;
assign v374f9f5 = hlock0_p & v3a5614c | !hlock0_p & v373a696;
assign v3759b2f = hbusreq1_p & v3a5891c | !hbusreq1_p & v3759032;
assign v3a6f555 = hmaster1_p & v372b3dd | !hmaster1_p & v3768774;
assign v3729830 = hmaster0_p & v377d1dc | !hmaster0_p & v2092ef2;
assign v3759f77 = hlock5_p & v3a669bc | !hlock5_p & !v8455ab;
assign v37466cb = hbusreq6_p & v3a6fa50 | !hbusreq6_p & v8455ab;
assign v3a7147e = hmastlock_p & v3a5fcfc | !hmastlock_p & !v8455ab;
assign v37755b2 = hmaster2_p & v3769ae2 | !hmaster2_p & v8455b7;
assign v376f42c = hbusreq8 & v376c8f2 | !hbusreq8 & v3a70040;
assign v3771428 = hmaster1_p & v3a2a911 | !hmaster1_p & v374b074;
assign v39a4ce0 = jx2_p & v3a6b368 | !jx2_p & v376662b;
assign v376cc45 = hmaster1_p & v373425d | !hmaster1_p & v8455ab;
assign v373186a = hbusreq0 & adf78a | !hbusreq0 & v3730ffe;
assign v3755e82 = hbusreq3_p & c511c2 | !hbusreq3_p & v372ab5a;
assign v375dd84 = hgrant5_p & v377d146 | !hgrant5_p & v3a6f3f8;
assign v3730f5d = hmaster1_p & v3a6fc5a | !hmaster1_p & v8455e7;
assign v3a6f9a4 = hmaster2_p & v377e904 | !hmaster2_p & v3777da6;
assign v3a60340 = hbusreq0 & v3751c8c | !hbusreq0 & !v1e37cd6;
assign v3a713ef = hbusreq5_p & v373e72e | !hbusreq5_p & v3a60e38;
assign v3a6f1c5 = hbusreq3_p & v2092ffc | !hbusreq3_p & v3a70376;
assign v3a62481 = hmaster0_p & v3a707d0 | !hmaster0_p & v37390c9;
assign v37534c6 = hmaster0_p & v3722de8 | !hmaster0_p & v2092ec6;
assign v372626a = hmaster2_p & v37c033d | !hmaster2_p & v3a5b693;
assign v3a53873 = hlock0 & v3a70a88 | !hlock0 & v3754a42;
assign v375c358 = hbusreq7_p & v377fab4 | !hbusreq7_p & v8455ab;
assign v3737478 = hgrant4_p & v3a624da | !hgrant4_p & v3a712b2;
assign v37286f3 = hmaster0_p & v37372a1 | !hmaster0_p & v3757765;
assign v37639a1 = hbusreq8_p & v373a4a8 | !hbusreq8_p & v3a5fc34;
assign v372f3a4 = hbusreq7 & v3772a15 | !hbusreq7 & v3a6f45d;
assign v3769630 = hbusreq4_p & v3a5fdd3 | !hbusreq4_p & !v3a627cc;
assign v3a71265 = hgrant2_p & v375b7bd | !hgrant2_p & v3745c8f;
assign v3a7092f = hmaster1_p & v3750b5b | !hmaster1_p & v3a588e5;
assign v373abb7 = hgrant2_p & v37565a5 | !hgrant2_p & v377e26b;
assign v373cdb0 = hgrant2_p & v8455ab | !hgrant2_p & v3a58dac;
assign v3767385 = hlock4 & v3770fbc | !hlock4 & v3a55838;
assign v3757772 = hgrant6_p & v8455ab | !hgrant6_p & v3a6f83c;
assign v3732415 = hbusreq2_p & v3729c6b | !hbusreq2_p & v8455ab;
assign v372bfcc = hmaster2_p & v8455ab | !hmaster2_p & v376b21a;
assign v3a6e7a4 = hlock8_p & v375408d | !hlock8_p & v3771804;
assign v3a70e6b = hbusreq0 & v377c3ad | !hbusreq0 & v373bd6c;
assign v37430e7 = hbusreq0 & v8455b3 | !hbusreq0 & !v8455ab;
assign v372fe57 = hmaster1_p & v2ff9190 | !hmaster1_p & v3752ab6;
assign v375259d = hbusreq8_p & v3725a65 | !hbusreq8_p & v3763832;
assign v37463a6 = hgrant2_p & v3779e45 | !hgrant2_p & v37773fa;
assign v376454b = hgrant3_p & v3a5e485 | !hgrant3_p & !v3738ce7;
assign v3764e52 = hbusreq4 & v3769160 | !hbusreq4 & v8455ab;
assign v375e074 = hmaster1_p & v373a1b4 | !hmaster1_p & v372535d;
assign v3764210 = hmaster1_p & v3a65b2b | !hmaster1_p & v37605ab;
assign v374b199 = hmaster1_p & v37795d3 | !hmaster1_p & v374177d;
assign v37728d0 = hlock1_p & v3728608 | !hlock1_p & v8455ab;
assign v3739417 = hbusreq3 & v3a6dc08 | !hbusreq3 & v8455b0;
assign v39e9c6f = hgrant1_p & v3a70f83 | !hgrant1_p & v8455ab;
assign v373eedf = hbusreq1_p & v3a71476 | !hbusreq1_p & v8455ab;
assign v375c19b = hmaster2_p & v3a635ea | !hmaster2_p & v374f9c6;
assign v3761611 = stateG10_1_p & v37328bf | !stateG10_1_p & v37275a7;
assign v375ec4e = hmaster2_p & v8455ab | !hmaster2_p & !v3a57012;
assign v3776ace = hgrant6_p & v8455ab | !hgrant6_p & v377bb56;
assign v372d279 = hgrant2_p & v3a5f50e | !hgrant2_p & v3a606ee;
assign v375534d = hmaster0_p & v8455ab | !hmaster0_p & !v8455e7;
assign d4044f = hmaster1_p & v37730d2 | !hmaster1_p & v3741a07;
assign v3a573af = hbusreq5 & v3a6802f | !hbusreq5 & v3a7098f;
assign v3765ef0 = hbusreq4 & v380974c | !hbusreq4 & v8455b3;
assign v3a6fb1f = hbusreq6 & v376641b | !hbusreq6 & v376728e;
assign v3a6ebbc = hlock3_p & v374b57c | !hlock3_p & v8455b7;
assign v3778afd = hgrant4_p & v372f3e0 | !hgrant4_p & b4ac83;
assign v37682c0 = hbusreq2_p & v3a635ea | !hbusreq2_p & v375408a;
assign v377987e = hbusreq7_p & v3747079 | !hbusreq7_p & v3752da9;
assign v376f768 = hlock3 & v3753163 | !hlock3 & v375039e;
assign v37313fa = hmaster0_p & v377c7ae | !hmaster0_p & v3a553aa;
assign v3737ea9 = hlock4_p & v8455ab | !hlock4_p & v2092ab0;
assign v3a6ba91 = hmaster0_p & v37673fe | !hmaster0_p & v3808e2e;
assign v3a6f578 = hgrant5_p & v3730587 | !hgrant5_p & v3727d77;
assign v3a71039 = hlock7_p & v3a6f118 | !hlock7_p & v3a6f154;
assign v3a5eefd = hmaster1_p & v3769f23 | !hmaster1_p & v3730c86;
assign v3768f7f = hbusreq4 & v37578d4 | !hbusreq4 & v35b774b;
assign v3a5b7db = hgrant4_p & v376af6a | !hgrant4_p & v377d367;
assign v3730a8b = hmaster2_p & v3a70957 | !hmaster2_p & v374aa71;
assign v3a548a0 = hmaster0_p & v35b70ee | !hmaster0_p & v8455ab;
assign v376dc26 = hbusreq4_p & v3722f65 | !hbusreq4_p & v8455ab;
assign v375993d = hbusreq5_p & v37784a0 | !hbusreq5_p & !v3a71637;
assign v3779195 = hbusreq7_p & v376dffd | !hbusreq7_p & v3a5fa09;
assign v373abae = hlock6 & v3757254 | !hlock6 & v3a61d2e;
assign v37510a5 = hbusreq4_p & v3a5f69c | !hbusreq4_p & v3a6f5a0;
assign v376d955 = hlock3_p & v8455ab | !hlock3_p & v373fe5e;
assign v37243ac = hbusreq7 & v374be73 | !hbusreq7 & v376ae9f;
assign v3749e13 = hlock0 & v372e83f | !hlock0 & v3a54455;
assign v374b7d8 = hlock5 & v374b4f8 | !hlock5 & v373794a;
assign v3a62f0b = hlock6_p & v373389a | !hlock6_p & !v374b25d;
assign v3a6f914 = hbusreq6 & v374956a | !hbusreq6 & v37574d2;
assign v3768ec7 = hmaster2_p & v2925c39 | !hmaster2_p & v3a62abc;
assign v3738336 = hmaster2_p & v3a6422d | !hmaster2_p & v8455ab;
assign v373a7a6 = stateG10_1_p & v8455ab | !stateG10_1_p & v37233a4;
assign v377b7d0 = hbusreq8 & v373643b | !hbusreq8 & v3a6f1c8;
assign v28896f0 = hmaster0_p & v38072bd | !hmaster0_p & v3a6a9d7;
assign v3769e94 = hbusreq4_p & v3a6ac2e | !hbusreq4_p & v3764898;
assign v376cd09 = hbusreq5 & v376c422 | !hbusreq5 & v37333de;
assign v374a8a5 = hbusreq0 & v372437c | !hbusreq0 & v375564e;
assign v37284f8 = hlock6_p & v8455ab | !hlock6_p & !v3753f1a;
assign v3732302 = hlock0_p & v8455b7 | !hlock0_p & v374e61f;
assign v3807bf8 = busreq_p & v3809adf | !busreq_p & !v3751094;
assign v3743d58 = hgrant2_p & v3759b2f | !hgrant2_p & v37790a9;
assign v3a6f63c = hmaster2_p & v3a603a1 | !hmaster2_p & v8455ab;
assign v3a71352 = hready_p & v3742ed3 | !hready_p & v39ed7e4;
assign d1e3dd = hgrant4_p & v3807f45 | !hgrant4_p & v37740fd;
assign db0673 = hbusreq1 & v374f307 | !hbusreq1 & v8455ab;
assign v3a65b10 = hgrant5_p & v374d7a7 | !hgrant5_p & v377fb50;
assign v373512b = hlock4_p & v3a5b5d3 | !hlock4_p & v3a658bf;
assign v3738270 = hlock5_p & v3a6f726 | !hlock5_p & !v3724325;
assign v3a70bee = hbusreq5_p & v3774e5a | !hbusreq5_p & v3a66514;
assign v3748cce = hbusreq6_p & v37406d2 | !hbusreq6_p & v3753dab;
assign v3a55c48 = jx0_p & v372664e | !jx0_p & !v376ff42;
assign v3774103 = hlock5_p & v375e444 | !hlock5_p & v3a6fe3d;
assign v3730145 = hmaster0_p & v3761b5e | !hmaster0_p & v3770331;
assign v37443ab = hbusreq2_p & v8455bb | !hbusreq2_p & !v8455ab;
assign v373f9df = hmaster2_p & v8455ab | !hmaster2_p & v3a55959;
assign v374b0a3 = hbusreq5_p & v373100d | !hbusreq5_p & v3731994;
assign v3a6f449 = hbusreq5_p & v37493b4 | !hbusreq5_p & v37512c1;
assign v3a6e8a4 = hgrant2_p & v8455ab | !hgrant2_p & v37753f2;
assign aa5585 = jx1_p & v3754aa8 | !jx1_p & v37451db;
assign v3a7130b = hmaster0_p & v374314f | !hmaster0_p & v3740c92;
assign v3a54789 = hmaster3_p & v3a5e687 | !hmaster3_p & v3a6f731;
assign v375b777 = hbusreq8_p & v3a70c90 | !hbusreq8_p & v3768c98;
assign v3806e35 = hgrant2_p & v8455ab | !hgrant2_p & !v3a658ad;
assign v3a6673e = hbusreq7 & v3a704f5 | !hbusreq7 & v3733483;
assign v37276a0 = hmaster1_p & v3a61149 | !hmaster1_p & v374e21e;
assign v375ec23 = hmaster2_p & v373e625 | !hmaster2_p & v37447e9;
assign v37515e1 = hgrant5_p & v3774dcd | !hgrant5_p & v37684e6;
assign v373e055 = hbusreq5_p & v3727385 | !hbusreq5_p & v8455ab;
assign v3744c5e = hmaster1_p & v3722b21 | !hmaster1_p & !v374975c;
assign v372b4a0 = hbusreq4_p & v3a6aa9f | !hbusreq4_p & v8455ab;
assign v3728f25 = hgrant4_p & v8455c1 | !hgrant4_p & v3766f14;
assign v3a65671 = hmaster2_p & v377c931 | !hmaster2_p & v23fd83f;
assign v3729435 = hmaster0_p & v3a6ff5b | !hmaster0_p & v3745d9c;
assign v3743ff2 = hgrant4_p & v37782c9 | !hgrant4_p & v373350e;
assign v376634b = hgrant7_p & v373a2cc | !hgrant7_p & !v3a71461;
assign v3a65b39 = hlock5_p & v3762fdb | !hlock5_p & v8455ab;
assign v376e568 = hgrant0_p & d70af8 | !hgrant0_p & v8455ab;
assign v373e86e = hbusreq7_p & v3a59c73 | !hbusreq7_p & v372fdfd;
assign v373339c = hbusreq0_p & v3a635ea | !hbusreq0_p & v37567c7;
assign v37385fc = hlock8_p & v37654bc | !hlock8_p & v992750;
assign v3a6d003 = hmaster2_p & v3775303 | !hmaster2_p & v3a5f8d0;
assign v3775544 = jx0_p & v37565d3 | !jx0_p & !v376cef0;
assign v373665b = hmaster2_p & v3735272 | !hmaster2_p & v373f911;
assign v3748bb1 = hgrant1_p & v3a6f4d3 | !hgrant1_p & v3a6f252;
assign v3758b89 = hbusreq4_p & v376b8f8 | !hbusreq4_p & v375a677;
assign v3a70fcd = hmaster1_p & v3776864 | !hmaster1_p & v375918d;
assign v377926d = hmaster2_p & v3a706a0 | !hmaster2_p & v374b6ba;
assign v372311c = hmaster0_p & v3a68426 | !hmaster0_p & v373e2f9;
assign v3a64792 = hbusreq4 & v373a27c | !hbusreq4 & v8455ab;
assign v3756764 = hmaster2_p & v375a268 | !hmaster2_p & !v377b6ce;
assign v3767cd6 = hgrant3_p & v35b7299 | !hgrant3_p & !bd3213;
assign v3a6cf15 = hbusreq8 & v373adf1 | !hbusreq8 & v8455bb;
assign v3a5fa09 = hgrant5_p & v376e66e | !hgrant5_p & v3a6367f;
assign v3a5a853 = hbusreq6_p & v376803b | !hbusreq6_p & v3737534;
assign v374ebb6 = hmaster2_p & v372ff0a | !hmaster2_p & v375d3cd;
assign v376a822 = hgrant2_p & v3a5b5d3 | !hgrant2_p & v3a6f842;
assign c7355c = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a711da;
assign v375a38b = hlock4_p & v3a6ff67 | !hlock4_p & v8455cb;
assign v3a6b29f = hmaster0_p & v8455ab | !hmaster0_p & v376c22c;
assign v3a576a4 = hmaster2_p & v3758fa8 | !hmaster2_p & v3735272;
assign v372f76c = hlock0 & v3752cf6 | !hlock0 & v3a6d840;
assign v373e49f = hbusreq0 & v37302ea | !hbusreq0 & v377c0fe;
assign v3722e59 = hmaster2_p & v3758cec | !hmaster2_p & v8455ab;
assign v37526a5 = hmaster2_p & v377ea20 | !hmaster2_p & v3a6bb45;
assign v37456a9 = hbusreq6 & v376e89b | !hbusreq6 & v3a70d99;
assign v37235f9 = hgrant6_p & v3a66e4c | !hgrant6_p & v38072fb;
assign v372beb8 = hlock0_p & v3a68426 | !hlock0_p & v8455b7;
assign v377d41d = hlock2 & v3773043 | !hlock2 & v3a5eafa;
assign v37470f6 = hgrant2_p & v8455ab | !hgrant2_p & v375b93d;
assign v373b5b8 = hgrant6_p & v375d877 | !hgrant6_p & v373342f;
assign v372790e = hbusreq5_p & v3742649 | !hbusreq5_p & v37723b7;
assign v373b48c = hmaster2_p & v3a62a6d | !hmaster2_p & v8455ab;
assign v373f1ac = hbusreq6 & v3778fec | !hbusreq6 & v3a6eead;
assign v37712f8 = hbusreq0 & v376d935 | !hbusreq0 & v3a6180b;
assign v3764e3f = hbusreq8 & v3741cc4 | !hbusreq8 & v3a60276;
assign v3a6fa7c = hmaster0_p & v377ce3f | !hmaster0_p & d54152;
assign v3a6c7f2 = jx1_p & v8455ab | !jx1_p & v37522e8;
assign v374b3bf = hlock0_p & v37757e0 | !hlock0_p & v3a67d6f;
assign v3a5b57a = hbusreq0 & v372d816 | !hbusreq0 & v3746fd4;
assign v3a6a1b9 = hbusreq2 & v376a8d5 | !hbusreq2 & v3a57309;
assign v373cb54 = hbusreq6 & v3a70bc8 | !hbusreq6 & v8455ab;
assign v3806c70 = hmaster1_p & v3a713ad | !hmaster1_p & v375bcf7;
assign v375da9f = hmaster2_p & v35772a6 | !hmaster2_p & v3770559;
assign v3a6ff5e = hbusreq7_p & v3759421 | !hbusreq7_p & v3a7033f;
assign v373dc68 = hbusreq0 & v3767b66 | !hbusreq0 & v3775b30;
assign v3a60395 = hmaster2_p & v377834b | !hmaster2_p & v8455ab;
assign v3a705c7 = hmaster0_p & afdeb4 | !hmaster0_p & v23fdebb;
assign v375dc5f = hmaster2_p & v376111d | !hmaster2_p & !v376b4e1;
assign v3808531 = hmaster0_p & v3a5af94 | !hmaster0_p & v37441fb;
assign v3746351 = hbusreq4_p & v3763104 | !hbusreq4_p & v8455bf;
assign v3a613cc = hbusreq0 & v3806e7b | !hbusreq0 & v375314d;
assign v3a70672 = hlock1_p & v2925c39 | !hlock1_p & !v8455ab;
assign v3a706c2 = hbusreq5_p & v374cbc3 | !hbusreq5_p & v8455ab;
assign v375463f = hgrant0_p & v8455ab | !hgrant0_p & v37245d9;
assign v3a6877a = hbusreq7_p & v373f8c4 | !hbusreq7_p & v3a6652b;
assign v3742a4e = hmaster1_p & v3a538ba | !hmaster1_p & v3730c86;
assign v3726a78 = hbusreq7_p & v3a6178e | !hbusreq7_p & !v375c041;
assign v1e37a35 = hmaster1_p & v3737928 | !hmaster1_p & !v376ad8c;
assign v374ad16 = hbusreq6_p & v3723430 | !hbusreq6_p & v8455e7;
assign v3736894 = hmaster0_p & v375e574 | !hmaster0_p & v3a6ab7f;
assign v3a61e10 = hbusreq2_p & v377eb2d | !hbusreq2_p & v8455b0;
assign v9d35e2 = hmaster2_p & v35772a6 | !hmaster2_p & v3a64ded;
assign v3a5d356 = hgrant0_p & v375d690 | !hgrant0_p & v377b673;
assign v3a626bd = hmaster1_p & v93ca8c | !hmaster1_p & !v37702c5;
assign v3a702ff = hgrant2_p & v374a6fc | !hgrant2_p & v3748f48;
assign v373d119 = jx1_p & v380700f | !jx1_p & v3a532f2;
assign v37576af = hbusreq7_p & v3733cf4 | !hbusreq7_p & v3a65ea7;
assign v3a61149 = hlock5 & v3a70d2a | !hlock5 & v3770a5a;
assign v376df43 = start_p & v3a5a496 | !start_p & v377f384;
assign v3a5f375 = jx1_p & v8455ab | !jx1_p & !v3a5ef0d;
assign v3773e34 = hbusreq6 & v3776441 | !hbusreq6 & v8455e7;
assign v3a59918 = stateG2_p & v8455ab | !stateG2_p & v3a6cd1b;
assign v3a6d80d = hbusreq7_p & v3a70623 | !hbusreq7_p & v3807550;
assign v3a5a5a7 = hbusreq5 & v3767797 | !hbusreq5 & v3770ad8;
assign v3a705df = hbusreq5 & v3a5aac9 | !hbusreq5 & v8455ab;
assign v3a6feee = hgrant4_p & v3a53eeb | !hgrant4_p & v3739bcd;
assign v3a5a06e = hmaster1_p & v3a5af94 | !hmaster1_p & v37552cb;
assign v3a6fdd7 = hbusreq8 & v373fe0d | !hbusreq8 & v3734ba4;
assign v3a60711 = hbusreq3 & v8455ab | !hbusreq3 & v3776aa8;
assign v3a5bd9c = hmaster1_p & v376b743 | !hmaster1_p & v376a40c;
assign v3766a74 = hlock6_p & v372d203 | !hlock6_p & v8455b0;
assign v3a62d56 = hgrant2_p & v37664d0 | !hgrant2_p & v8455ab;
assign v3768616 = hmaster2_p & a747d7 | !hmaster2_p & v3a6890e;
assign v3a57d41 = hmaster2_p & v3a7033d | !hmaster2_p & !v8455ab;
assign v3a6f765 = hmaster2_p & v373325f | !hmaster2_p & !v374e542;
assign v3a6e159 = hbusreq6_p & v373fb30 | !hbusreq6_p & v3a69b5c;
assign v3733c70 = jx0_p & v3733ac0 | !jx0_p & v37418f3;
assign v37625a7 = hmaster0_p & v3761719 | !hmaster0_p & v3a60a24;
assign v3756bd8 = hmaster2_p & v9b03cc | !hmaster2_p & v376bb26;
assign v37436cf = hgrant6_p & v3a6c7fe | !hgrant6_p & v373374d;
assign v372f58a = jx3_p & v3a6c7f2 | !jx3_p & v8455ab;
assign v373d825 = hbusreq3_p & v373fe5e | !hbusreq3_p & v8455e7;
assign v3a65155 = hbusreq5_p & v3772140 | !hbusreq5_p & v3776a2e;
assign v3a703ac = hbusreq2 & v373fe5e | !hbusreq2 & !v3753f1a;
assign b4444b = hbusreq3 & v3a70e9f | !hbusreq3 & v8455ab;
assign v372700e = jx0_p & v376e4c5 | !jx0_p & v3a6de3a;
assign v377070e = hbusreq0 & v37680af | !hbusreq0 & v375924f;
assign v37660dd = hbusreq6_p & v3a69487 | !hbusreq6_p & v375d288;
assign v374c9ab = hbusreq5 & v8455b0 | !hbusreq5 & v8455ab;
assign v37277ab = hbusreq8_p & v3a635ea | !hbusreq8_p & v372552c;
assign v376ee08 = jx2_p & v3734ef4 | !jx2_p & v3a674a8;
assign v3a71309 = hmaster1_p & v3745ced | !hmaster1_p & v37658d9;
assign v3a61d2e = hbusreq2_p & v374a430 | !hbusreq2_p & v3a68d2e;
assign v37784d0 = hmaster0_p & v3a6dafc | !hmaster0_p & v3a713a7;
assign v373cf9c = hbusreq0 & v3a68310 | !hbusreq0 & v9a2413;
assign v3a70267 = hmaster2_p & v374ab22 | !hmaster2_p & v3771c85;
assign v375a023 = hmaster2_p & v372433d | !hmaster2_p & v3768ba1;
assign v375aeb3 = hgrant5_p & v8455ab | !hgrant5_p & v374e663;
assign v374544f = hmaster2_p & v3a704cc | !hmaster2_p & v8455ab;
assign v3a5a63c = hbusreq6_p & v37601d6 | !hbusreq6_p & v376bc6a;
assign v23fd83c = hmaster2_p & v3a70fda | !hmaster2_p & v377d1dc;
assign v3769039 = hbusreq0_p & v3779324 | !hbusreq0_p & v373da69;
assign v3a53d98 = hmaster1_p & v3a6f51e | !hmaster1_p & v3a706f4;
assign v3a6ef0e = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a70a7f;
assign v3a625d8 = hgrant6_p & v3766b5e | !hgrant6_p & v377a6f2;
assign v3a70819 = hlock7 & v373b1bb | !hlock7 & v376e20f;
assign v3769c43 = hbusreq6 & v374d2b3 | !hbusreq6 & v3a703d3;
assign v3a6f501 = hbusreq4_p & v3a635ea | !hbusreq4_p & v37651c2;
assign v3729cbe = hbusreq6_p & v377c068 | !hbusreq6_p & v377b860;
assign v375add1 = hmaster0_p & v3745589 | !hmaster0_p & v377d1dc;
assign v3762949 = hgrant2_p & v8455ab | !hgrant2_p & v3745dc7;
assign v3a625a1 = hmaster2_p & v8455ab | !hmaster2_p & v3a70c39;
assign v3a621e7 = hgrant4_p & v374acbe | !hgrant4_p & v375c70c;
assign v37467be = hmaster2_p & v3a61a7f | !hmaster2_p & v377204f;
assign v375449f = hmaster2_p & v373f647 | !hmaster2_p & !v3768a41;
assign a2a6f3 = hbusreq5 & v375874f | !hbusreq5 & v3753576;
assign v3a5e922 = hlock6_p & v3a568f7 | !hlock6_p & v373c755;
assign v3724e14 = hmaster1_p & v3a669c6 | !hmaster1_p & v375ecd4;
assign v3a70929 = hbusreq4_p & v3743b98 | !hbusreq4_p & v37759b6;
assign v3747452 = hbusreq5 & v373c005 | !hbusreq5 & v3764dac;
assign v3750b85 = hgrant2_p & v8455ab | !hgrant2_p & v377d6e5;
assign v372d071 = hmaster1_p & v3a6f6bc | !hmaster1_p & v373f4dd;
assign v2092ff6 = hmaster1_p & v8455ab | !hmaster1_p & v3773107;
assign v3a714cf = hgrant4_p & v8455ab | !hgrant4_p & v376ef46;
assign v3750d37 = locked_p & v2925c39 | !locked_p & !v8455ab;
assign v377c0f5 = hgrant0_p & v8455ab | !hgrant0_p & v3748bb7;
assign v3733360 = hbusreq6 & v37344a0 | !hbusreq6 & v3765261;
assign d70cde = hbusreq7_p & v373d687 | !hbusreq7_p & v376604d;
assign v374fad3 = hgrant0_p & v375f3f0 | !hgrant0_p & !v3771728;
assign v37400ba = hbusreq5 & v373e28c | !hbusreq5 & v376de5c;
assign v3748400 = hbusreq5 & v374cb0f | !hbusreq5 & v376a3f7;
assign v3a6f4fd = hbusreq4 & v3a5ab85 | !hbusreq4 & v373bd6c;
assign v377e24d = hbusreq4 & v373b1cb | !hbusreq4 & v8455ab;
assign v37497b1 = hgrant0_p & v3a637dc | !hgrant0_p & b8006a;
assign v3a60a23 = hbusreq0 & v3a6bedb | !hbusreq0 & v377c31d;
assign v3728dd0 = hbusreq5 & v3755e1f | !hbusreq5 & v8455ab;
assign v3770fb6 = hbusreq0_p & v377ba55 | !hbusreq0_p & v8455ab;
assign v3806572 = hgrant1_p & v8455ab | !hgrant1_p & !v3764463;
assign v3806912 = hgrant0_p & v8455ab | !hgrant0_p & v37619dc;
assign v3a63002 = hlock4 & v3778454 | !hlock4 & v374d28d;
assign v374b88a = jx0_p & v3a5921b | !jx0_p & a5f27e;
assign v3a6ef95 = hgrant4_p & v3a6c970 | !hgrant4_p & v3726204;
assign aa3e48 = hgrant3_p & v8455ab | !hgrant3_p & v3740060;
assign v3750c57 = hmaster1_p & v3a584be | !hmaster1_p & v39ebb63;
assign v375c3b0 = hlock1_p & v2ff9362 | !hlock1_p & v3a63bb0;
assign v372d1a4 = hbusreq2_p & v376fbcd | !hbusreq2_p & v3a6b6d2;
assign v2aca83b = hbusreq8_p & v3a5bf56 | !hbusreq8_p & v376ec1d;
assign v3a6bf3c = hmaster0_p & v8455ab | !hmaster0_p & v373fd4c;
assign v3a70cb4 = hgrant5_p & v3727d4c | !hgrant5_p & v374b8fa;
assign v3a65b0a = hmaster0_p & v37797d5 | !hmaster0_p & v3761c61;
assign v3a6dfc6 = hgrant2_p & v375318f | !hgrant2_p & v8455ab;
assign v3a7085f = hgrant4_p & v8455ab | !hgrant4_p & v3a66545;
assign v3726240 = hlock5 & v37380be | !hlock5 & v374e179;
assign v37280a3 = hlock5 & v3727c91 | !hlock5 & v3a5e2eb;
assign v373eb05 = hmaster3_p & v3724579 | !hmaster3_p & v3737f16;
assign v3761db0 = hmaster0_p & v375351d | !hmaster0_p & v3a7004b;
assign v377b48b = hmaster0_p & v380714f | !hmaster0_p & !v3a71505;
assign v3a702b6 = hbusreq0 & v3754b83 | !hbusreq0 & v3755305;
assign v3a6f05e = hgrant4_p & v3a6feb3 | !hgrant4_p & v375f9ec;
assign v3a61482 = hbusreq6_p & v3743338 | !hbusreq6_p & v3750b9e;
assign v374bace = hbusreq5 & v3a68232 | !hbusreq5 & v8455ab;
assign v373f492 = hgrant2_p & v8455ab | !hgrant2_p & v377ba5a;
assign v3807026 = hbusreq6_p & v3a6fa49 | !hbusreq6_p & v3762be8;
assign v375fe02 = hmaster0_p & v372b390 | !hmaster0_p & v3775219;
assign v3746fe7 = hgrant5_p & v8455ab | !hgrant5_p & v3a6947c;
assign baec07 = hbusreq4_p & v376f56d | !hbusreq4_p & v374cbe3;
assign v376ce37 = hbusreq2 & v3a6f32f | !hbusreq2 & !v3a5614c;
assign v3779070 = hbusreq4_p & v375d00a | !hbusreq4_p & v8455ab;
assign v3722da3 = hgrant2_p & v3a61e10 | !hgrant2_p & v8455ab;
assign v376011a = hgrant6_p & v377938d | !hgrant6_p & v3a712d6;
assign v376c3fd = hmaster0_p & v373a1d7 | !hmaster0_p & v3a5bd69;
assign v375e9c8 = hmaster0_p & v37469c4 | !hmaster0_p & v3a577de;
assign v3758c5e = hgrant5_p & v373dc42 | !hgrant5_p & v3a63930;
assign v3a64b9b = hbusreq5 & v8455ab | !hbusreq5 & v3774b12;
assign v3a6c63e = hlock2 & v376f7a7 | !hlock2 & v38099e8;
assign v3a5a2d4 = hmaster1_p & v3577306 | !hmaster1_p & v376b03d;
assign v375cdb1 = hbusreq3_p & v37720d8 | !hbusreq3_p & v8455ab;
assign v374f4ae = hgrant7_p & v8455ab | !hgrant7_p & v3754c09;
assign v375316c = hmaster2_p & v35b7092 | !hmaster2_p & v3756304;
assign v3a6403e = hgrant6_p & v8455ab | !hgrant6_p & v37470f6;
assign v37417f6 = hbusreq1_p & v37543c2 | !hbusreq1_p & v3761611;
assign v376bf69 = hbusreq3 & v35b7808 | !hbusreq3 & v377eb9d;
assign v3a5d41e = hbusreq7_p & v37bfd3a | !hbusreq7_p & v31c3043;
assign v3724db7 = hbusreq6 & v377b9ab | !hbusreq6 & v8455ab;
assign v372e05a = hmaster2_p & v373dfec | !hmaster2_p & v3728f25;
assign v3726efb = hbusreq6 & v3a6847c | !hbusreq6 & v8455ab;
assign v376d7ee = hbusreq2_p & v3a5b2fd | !hbusreq2_p & v3724f7b;
assign v3a5cc14 = hmaster0_p & v3a6e09b | !hmaster0_p & !v373a246;
assign v37358ae = hmaster1_p & v3a62542 | !hmaster1_p & v3a6fb2f;
assign v37777d1 = hmaster1_p & v3a635ea | !hmaster1_p & v3a5982a;
assign v37582e7 = hmaster1_p & v3a7079a | !hmaster1_p & v374c8b8;
assign v39748fd = hbusreq7_p & v375eb37 | !hbusreq7_p & v3723089;
assign v3a70b8f = hbusreq5_p & v3a6fd66 | !hbusreq5_p & v372f0bb;
assign v3746a7e = hmaster2_p & v3738d51 | !hmaster2_p & v377d69c;
assign v37262ab = hbusreq5_p & v3762dc3 | !hbusreq5_p & v372294a;
assign v3751291 = hlock4 & v372a9a6 | !hlock4 & v3a6f79b;
assign v374ac57 = hmaster1_p & v3740bb7 | !hmaster1_p & v8e42b4;
assign v373a3c3 = hbusreq5_p & v3773340 | !hbusreq5_p & v3773015;
assign d973ae = hbusreq7 & v3a5ddef | !hbusreq7 & v374d163;
assign v375811b = hmaster3_p & v3a5e2fa | !hmaster3_p & v377d223;
assign v377831d = hlock0_p & v37718fb | !hlock0_p & v3a67d6f;
assign v37774b6 = hlock8 & v374132e | !hlock8 & v3a6ebee;
assign v3a60f21 = hmaster0_p & v8455ab | !hmaster0_p & v3724779;
assign v376618c = hgrant4_p & v377b6ce | !hgrant4_p & !v3757727;
assign v3734bc3 = hlock3_p & v3738e79 | !hlock3_p & !v8455ab;
assign a747d7 = hgrant4_p & v3739190 | !hgrant4_p & v3a70554;
assign v37431ce = hbusreq7 & v3a713ea | !hbusreq7 & v3771933;
assign v3770fbc = hbusreq4 & v3a55838 | !hbusreq4 & v373f3b5;
assign v3a6f8b9 = hmaster1_p & v209312a | !hmaster1_p & v373a791;
assign v3754f5d = hlock2 & v374d40b | !hlock2 & v23fdf85;
assign v3a697a5 = hmaster0_p & v3740212 | !hmaster0_p & v3a594ab;
assign v3a650e9 = hmaster2_p & v35772a6 | !hmaster2_p & v3778b8c;
assign v377bcf5 = hmaster2_p & v3a58cfc | !hmaster2_p & !v1e38224;
assign v3a5f602 = hbusreq5_p & v375d417 | !hbusreq5_p & v37541c6;
assign v28896e3 = hbusreq0 & v3777666 | !hbusreq0 & v3a71660;
assign v3a7010d = hmaster0_p & v372f3b1 | !hmaster0_p & v88d9b8;
assign v37395f5 = hgrant6_p & v377f09a | !hgrant6_p & a69e17;
assign v377123e = hgrant2_p & v8455ab | !hgrant2_p & a17325;
assign v375a4f6 = hmaster1_p & v376aaee | !hmaster1_p & v373ed57;
assign v376f38d = hbusreq3_p & v374d3d7 | !hbusreq3_p & v3724d93;
assign v3725710 = hmaster2_p & v3747302 | !hmaster2_p & v3a687a7;
assign v3a71588 = hmaster0_p & v3743b64 | !hmaster0_p & v3758d6c;
assign v3a637fd = hlock7 & v3738259 | !hlock7 & v37475f4;
assign v374a526 = hgrant8_p & v3a6f7d4 | !hgrant8_p & v3a7092b;
assign v372e2eb = hbusreq7 & v3a64868 | !hbusreq7 & v8455ab;
assign v3752b8c = hmastlock_p & v377f108 | !hmastlock_p & !v8455ab;
assign v3a6f080 = hmaster1_p & v374a9d0 | !hmaster1_p & v3a707b9;
assign v3779a60 = hmaster2_p & v3731caa | !hmaster2_p & v3770bcd;
assign v377d23c = hbusreq7_p & v3a6fa57 | !hbusreq7_p & v376af81;
assign v3a7164f = hmaster1_p & v3729238 | !hmaster1_p & v3728040;
assign v377dfe2 = hgrant0_p & v3a64c10 | !hgrant0_p & !bbbe50;
assign v3a59c5e = hlock5 & v3a63f9a | !hlock5 & v3a7038a;
assign v3a5a76b = hbusreq2 & v3724e8e | !hbusreq2 & v377b774;
assign v3a6fe94 = hbusreq6_p & v337897a | !hbusreq6_p & v3a5988f;
assign v3a63545 = hbusreq6 & v3a704d5 | !hbusreq6 & v8455ab;
assign v377ba78 = hmaster2_p & v3a6ffb6 | !hmaster2_p & v9ed516;
assign v3760be5 = hmaster2_p & v375b429 | !hmaster2_p & v3730e98;
assign v373a013 = hbusreq6_p & v3777a52 | !hbusreq6_p & v3774cee;
assign v3a540a4 = hbusreq4 & v3a712ac | !hbusreq4 & v37283bb;
assign v3a60ab2 = hmaster2_p & v3a635ea | !hmaster2_p & v3770e95;
assign v376397d = hmaster2_p & v3a70374 | !hmaster2_p & v3a53e66;
assign v37629ba = jx0_p & v3a710d8 | !jx0_p & v377a0f2;
assign v3a6f7a2 = hbusreq4_p & v8455b7 | !hbusreq4_p & v37476fd;
assign v37622aa = hbusreq8 & v3a68b25 | !hbusreq8 & v3768500;
assign v3735fd1 = hmaster1_p & v37483ff | !hmaster1_p & v375c4f9;
assign v375dd92 = hmaster1_p & v376a9f7 | !hmaster1_p & v3a6fd9b;
assign v1e37c3e = hlock0_p & v376b4e1 | !hlock0_p & v8455ab;
assign v3a70d45 = hbusreq4 & v3a57506 | !hbusreq4 & v3a58a90;
assign v375a312 = hbusreq6_p & v3735f0b | !hbusreq6_p & v3a70cb6;
assign v3a56372 = hbusreq4 & v3724273 | !hbusreq4 & v8455ab;
assign v3a713b7 = hmaster2_p & v3774bad | !hmaster2_p & v8455b3;
assign v3a6924d = hbusreq7 & v3a700b9 | !hbusreq7 & v8455ab;
assign v372b551 = hmaster0_p & v37782c9 | !hmaster0_p & v3a71645;
assign v3a69a06 = hgrant1_p & v3757568 | !hgrant1_p & v3a6e7b3;
assign a75a41 = hbusreq6 & d44200 | !hbusreq6 & v8455ab;
assign v375fabf = hbusreq3_p & v8455e9 | !hbusreq3_p & v374f318;
assign v3731c1c = hbusreq6 & v374bc3e | !hbusreq6 & v377ce51;
assign v37771ca = hgrant6_p & v8455ab | !hgrant6_p & v37591da;
assign v373ed70 = hburst0 & v1e38224 | !hburst0 & !v8455e1;
assign v375a3dd = hmaster2_p & v377cfd9 | !hmaster2_p & v373e8ad;
assign v3a56c18 = hbusreq7 & v37352dc | !hbusreq7 & v3a62a6d;
assign v3a70649 = hbusreq6 & v3a70893 | !hbusreq6 & v8455ab;
assign v3737c52 = hgrant8_p & v3a70f25 | !hgrant8_p & v377d45b;
assign v3a6fc67 = hmaster0_p & v376e72d | !hmaster0_p & v3a7032a;
assign v209312a = hgrant4_p & v3735cb3 | !hgrant4_p & v3a6f75c;
assign v376fd7a = hlock4_p & v3725198 | !hlock4_p & v3a5b289;
assign v3a5f69c = hbusreq4 & v376e532 | !hbusreq4 & v3763104;
assign v3735049 = hbusreq7 & v37649e9 | !hbusreq7 & v8455ab;
assign v37536c3 = hbusreq0 & v3a708f6 | !hbusreq0 & v8455ab;
assign v38074a8 = hmaster0_p & v374e409 | !hmaster0_p & !v375c7b9;
assign v373087c = jx0_p & d9fd79 | !jx0_p & v3a54d04;
assign v377c0fa = jx0_p & v8455ab | !jx0_p & v37366b7;
assign v3a708a0 = hbusreq5 & v37252ee | !hbusreq5 & v8455ab;
assign v3a6a213 = hbusreq3_p & v3a60787 | !hbusreq3_p & v3733d6e;
assign v376da21 = hlock8_p & v3a70760 | !hlock8_p & !v8455ab;
assign v3a6ef30 = hmaster0_p & v376cebe | !hmaster0_p & v3a6e4cd;
assign v3a6ef8c = hburst1 & v3a5815e | !hburst1 & v3a713b2;
assign v37667d3 = hlock7 & v377cd41 | !hlock7 & v377a422;
assign v376d4ca = hlock6 & v3748797 | !hlock6 & v37326a5;
assign v37753da = hgrant2_p & v8455ab | !hgrant2_p & v376693b;
assign v3a712bc = hmaster1_p & v8455ab | !hmaster1_p & v3747d0e;
assign v3a568e4 = hgrant6_p & v373b209 | !hgrant6_p & v375a312;
assign v376358f = hbusreq4_p & v3742c6c | !hbusreq4_p & v3a68d2e;
assign v3a65612 = hmaster2_p & v3739ab4 | !hmaster2_p & v8455ab;
assign v372bc78 = jx1_p & v3773881 | !jx1_p & v8455ab;
assign v375fc56 = hbusreq7 & v3724c8c | !hbusreq7 & v8455bb;
assign v35b7805 = hmaster0_p & v37462ed | !hmaster0_p & v8455ab;
assign v37460cd = hmaster2_p & v375ced2 | !hmaster2_p & v3a6152c;
assign v357742d = hlock5_p & v3767b70 | !hlock5_p & v3771c85;
assign v37470d6 = hbusreq3_p & v3737ada | !hbusreq3_p & v8455ab;
assign v3727fd0 = hbusreq3 & v37282cf | !hbusreq3 & v37674c1;
assign v37346fe = hmaster1_p & v3a574bf | !hmaster1_p & v3771b8a;
assign v37693fe = hbusreq5_p & v3756683 | !hbusreq5_p & v3741435;
assign v3a2a144 = hgrant0_p & v377ba55 | !hgrant0_p & v8455ab;
assign v37453dd = hmaster2_p & v3737e2d | !hmaster2_p & v3a290f9;
assign v3a6e591 = hbusreq1 & v37566b2 | !hbusreq1 & !v8455ab;
assign v3a6fd21 = hmaster1_p & v372b219 | !hmaster1_p & v3769ec3;
assign v3a6de83 = hlock5 & v3a62403 | !hlock5 & v3763364;
assign v3a6c1ac = hbusreq2 & v373aecf | !hbusreq2 & !v8455ab;
assign v3a594a5 = hgrant2_p & v37676b8 | !hgrant2_p & v3747346;
assign v376afb1 = hmaster2_p & v376111d | !hmaster2_p & !v8455e1;
assign v3a6ae2d = hbusreq6 & v3a70641 | !hbusreq6 & v8455ab;
assign v3a61796 = jx3_p & v373fa73 | !jx3_p & aa5585;
assign v92a8d7 = hbusreq8 & v3727195 | !hbusreq8 & v374aa67;
assign v37410dc = hbusreq5 & v3a63306 | !hbusreq5 & v37316cb;
assign v373be25 = hbusreq1_p & v3809adf | !hbusreq1_p & v39a537f;
assign v372d525 = hbusreq7_p & v3763952 | !hbusreq7_p & v37286e7;
assign v374819d = hbusreq5 & v375808f | !hbusreq5 & v8455ab;
assign v3a6f91b = hbusreq8 & v3a579e2 | !hbusreq8 & v3728870;
assign v3762e7a = hbusreq8_p & v3737808 | !hbusreq8_p & v3a652db;
assign v372e34d = locked_p & v8455ab | !locked_p & !v3a580a0;
assign v3a539c3 = hgrant5_p & v8455ab | !hgrant5_p & v3757996;
assign v37733d9 = hbusreq5_p & v374055c | !hbusreq5_p & v3a70dd8;
assign v3a6de3a = hmaster1_p & v8455ab | !hmaster1_p & !v3759c80;
assign v376fc98 = hlock2 & v3752e46 | !hlock2 & v375d51e;
assign v3724f24 = hbusreq3_p & v372842d | !hbusreq3_p & v37366d2;
assign v3771507 = hgrant4_p & v8455ab | !hgrant4_p & v3777178;
assign v373cdb4 = stateA1_p & v3a67241 | !stateA1_p & v8455ab;
assign v375c0f1 = hbusreq5_p & v3a63def | !hbusreq5_p & !v376ea13;
assign v2ff9391 = hmaster2_p & v37247a3 | !hmaster2_p & !v373c07d;
assign v3725678 = hgrant2_p & v8455ab | !hgrant2_p & v3766d04;
assign v3a6ff57 = stateG3_2_p & v8455ab | !stateG3_2_p & !v373aaca;
assign v3768070 = hmaster2_p & v3771076 | !hmaster2_p & v373d9e0;
assign v373fb71 = hbusreq0 & v37291ce | !hbusreq0 & !v3760bd6;
assign v3a6bd87 = hbusreq1_p & v2aca977 | !hbusreq1_p & v3779e70;
assign v3a712e6 = hbusreq3_p & v3a5e24d | !hbusreq3_p & v3a54bc5;
assign v37477cb = hbusreq5_p & v37384a9 | !hbusreq5_p & v3a68c26;
assign v3a57593 = hgrant4_p & v8455ab | !hgrant4_p & v377a4c1;
assign v374b95f = hmaster0_p & v375b534 | !hmaster0_p & v376fd9a;
assign v372b7b7 = hlock3 & v3a70e84 | !hlock3 & v376d327;
assign v372a71e = hbusreq4_p & v3a635ea | !hbusreq4_p & v3753b6a;
assign v3779b95 = hbusreq2_p & v37309cf | !hbusreq2_p & !v8455ab;
assign v3a68954 = hlock4 & v37371b2 | !hlock4 & v376bea3;
assign v3a70083 = hgrant4_p & v3a630b7 | !hgrant4_p & v3a691f2;
assign a5f27e = hmaster1_p & v3726cd4 | !hmaster1_p & v8455ab;
assign v373769f = hbusreq6_p & v9f9402 | !hbusreq6_p & v37443ab;
assign v3a705ba = hmaster0_p & v3a6f094 | !hmaster0_p & v3763c9c;
assign v372b646 = hbusreq8 & v3a60223 | !hbusreq8 & v372ce94;
assign v3738e6e = hmaster2_p & v3760513 | !hmaster2_p & !v8455ab;
assign v3a6ff68 = jx0_p & v8455b5 | !jx0_p & !v3a63de8;
assign v3779fb2 = hbusreq2 & v3a7051c | !hbusreq2 & v8455ab;
assign v3747276 = hgrant2_p & v8455ab | !hgrant2_p & v3741d51;
assign v377f13c = hmaster2_p & v3a6f57c | !hmaster2_p & v3a70e46;
assign v376af98 = hlock4 & v3a6e793 | !hlock4 & v373e154;
assign v3736c94 = hbusreq0_p & v3a707de | !hbusreq0_p & v3a706c7;
assign v375c351 = hgrant4_p & v8455ab | !hgrant4_p & v3776ace;
assign v3a706b8 = hmaster1_p & v3a70cb2 | !hmaster1_p & !v372f9b4;
assign v3a6f371 = hmaster1_p & v8455b0 | !hmaster1_p & v3a68821;
assign v3772c57 = hbusreq2_p & v39ea273 | !hbusreq2_p & v374b8cb;
assign v3773661 = jx3_p & v3a70abd | !jx3_p & v377814d;
assign v3a7106e = hbusreq4_p & v3773bbc | !hbusreq4_p & v377aa2e;
assign v3a70117 = hmaster2_p & v37745a0 | !hmaster2_p & v37380c4;
assign v3a67b5e = hbusreq3_p & v372391f | !hbusreq3_p & !v375c5a8;
assign v376cdb7 = hmaster0_p & v3777467 | !hmaster0_p & v3747dd8;
assign v3773340 = hbusreq5 & v23fe37e | !hbusreq5 & v372cd37;
assign v373f92e = hbusreq6_p & v3773ee6 | !hbusreq6_p & v3a617b4;
assign v3a5f5b3 = hbusreq6_p & v3728f87 | !hbusreq6_p & v3756ec2;
assign v3762ac3 = hmaster1_p & v3a5acb3 | !hmaster1_p & v37705ec;
assign v3a6f610 = hmaster0_p & v37345aa | !hmaster0_p & v3769923;
assign v372ed34 = hbusreq4_p & v375c845 | !hbusreq4_p & v3a6f639;
assign v2ff8f1e = hbusreq3_p & v3752ec0 | !hbusreq3_p & v3a5903a;
assign v372ec32 = hmaster0_p & v1e38305 | !hmaster0_p & !v3a66088;
assign v3a6f7e2 = hgrant5_p & v37418ab | !hgrant5_p & v3768727;
assign v377c551 = hbusreq6 & v377123e | !hbusreq6 & v380730d;
assign v3770e2d = hgrant6_p & v375564e | !hgrant6_p & v376b576;
assign v3a6fc2d = hmaster2_p & v375ad1d | !hmaster2_p & v37310c2;
assign v3733886 = hmaster1_p & v376d66b | !hmaster1_p & v28896cd;
assign v3a6fa04 = hmaster0_p & v37741f1 | !hmaster0_p & v372e5fb;
assign v372aafb = hgrant4_p & v3a70401 | !hgrant4_p & !v3a71232;
assign v376f51c = hmaster0_p & v3a6e4ec | !hmaster0_p & v3764a7d;
assign v3a7094a = hlock0_p & v3a670a1 | !hlock0_p & v3772dd1;
assign v3a5f066 = hbusreq5 & v3a715df | !hbusreq5 & v8455ab;
assign v3741e80 = hgrant3_p & v37647e7 | !hgrant3_p & v37617d4;
assign v375bc6e = hgrant0_p & v8455e7 | !hgrant0_p & !v3725310;
assign v373a2f2 = hgrant2_p & v8455ab | !hgrant2_p & v3757fcc;
assign v375e510 = hbusreq7_p & v3725dd5 | !hbusreq7_p & v3738f37;
assign v3a6bddf = hmaster2_p & d99853 | !hmaster2_p & v8455e7;
assign v3806f0b = hbusreq5_p & v376f56d | !hbusreq5_p & v3a702ee;
assign v3a6f6cf = hmaster2_p & v3767d55 | !hmaster2_p & !v376888c;
assign v377ec1c = hgrant6_p & v3a6efa4 | !hgrant6_p & v8455ab;
assign v374e288 = hmaster2_p & v3763327 | !hmaster2_p & v3761ed2;
assign v3a70731 = hbusreq4_p & v372f37d | !hbusreq4_p & v37711c5;
assign v37726b0 = hgrant7_p & v3771a36 | !hgrant7_p & v372ef62;
assign v376b7ff = hbusreq7 & v3a63daa | !hbusreq7 & v377f80c;
assign v3a5d0d3 = hlock8_p & v337904a | !hlock8_p & v8455ab;
assign v375808f = hbusreq0 & v3a58218 | !hbusreq0 & v8455ab;
assign v3741216 = hgrant0_p & v8455ab | !hgrant0_p & v3758f3c;
assign v2093037 = hmaster0_p & v37795d3 | !hmaster0_p & v3a6fd45;
assign v3759c1f = hbusreq4_p & v372b88d | !hbusreq4_p & v8455ab;
assign v3a701ac = hmaster1_p & v3757966 | !hmaster1_p & v3761071;
assign v37659c5 = hbusreq5_p & v375b046 | !hbusreq5_p & v23fe316;
assign v8ac439 = hbusreq8 & v3773b4b | !hbusreq8 & v8455ab;
assign v37639c3 = hgrant6_p & v8455e7 | !hgrant6_p & v373ac39;
assign v3758c15 = hmaster0_p & v377b3c4 | !hmaster0_p & v374523d;
assign v373449a = hgrant3_p & ae7027 | !hgrant3_p & v372f747;
assign v372dd89 = hgrant2_p & v3778fec | !hgrant2_p & v3760343;
assign v377419a = hlock4 & b21e3c | !hlock4 & v3723635;
assign v3a7064e = hlock7_p & v3723d31 | !hlock7_p & !v8455ab;
assign v3774346 = hgrant3_p & v8455ab | !hgrant3_p & !v3a65532;
assign v37558eb = hbusreq0 & v3a6f8fb | !hbusreq0 & v8455ab;
assign v3725786 = hgrant2_p & v8455e7 | !hgrant2_p & !v3742cde;
assign v3a71684 = hbusreq0 & v3a71566 | !hbusreq0 & v3a6f0f2;
assign v3a710b4 = hmaster2_p & v8455b0 | !hmaster2_p & v3a63805;
assign v3a5b27f = hmaster2_p & v3724af9 | !hmaster2_p & v37386da;
assign v39eb4ab = hgrant4_p & v3775b81 | !hgrant4_p & v8455ab;
assign v37276d6 = hbusreq5 & v3732c0a | !hbusreq5 & v3a64f63;
assign v3775d59 = hbusreq2_p & v377144d | !hbusreq2_p & v3a6a0b0;
assign v3722f8e = hbusreq7_p & v375b929 | !hbusreq7_p & v3a694a5;
assign v3740f5d = hgrant4_p & v3a6e2d0 | !hgrant4_p & !v3a5e96b;
assign v3778fb2 = hbusreq3_p & v3759dd9 | !hbusreq3_p & v8455ab;
assign v3723e77 = hgrant6_p & v377f09a | !hgrant6_p & !v3a71563;
assign v3a56a52 = hgrant8_p & v8455ab | !hgrant8_p & v3a5e394;
assign v3728813 = hmaster2_p & v3756ef1 | !hmaster2_p & v377db88;
assign v3a58c95 = hbusreq7_p & v3775729 | !hbusreq7_p & v3765406;
assign v35b6dae = hbusreq7_p & v3a565bc | !hbusreq7_p & v37256b3;
assign v3a6f949 = hgrant3_p & v375da10 | !hgrant3_p & v3733c39;
assign v3a6f682 = hmastlock_p & v37493ce | !hmastlock_p & !v8455ab;
assign v3a70064 = jx1_p & v3a6fea0 | !jx1_p & v3a6f543;
assign v3a6ef07 = hlock8 & c47a78 | !hlock8 & v3a6fa1d;
assign v3a5bbaa = hmaster1_p & v3a5c75c | !hmaster1_p & v3a5c41b;
assign v3a67315 = hmaster0_p & v3a6e31f | !hmaster0_p & v38068ec;
assign v375590f = hbusreq6_p & v8455bf | !hbusreq6_p & v3a5f67d;
assign v3752648 = stateG10_1_p & v8455ab | !stateG10_1_p & !v377c2ba;
assign v376e0f5 = hlock5_p & v3a67471 | !hlock5_p & !v8455ab;
assign v1e38282 = hbusreq4 & v3a6fd37 | !hbusreq4 & v8455ab;
assign v3a6f59d = hbusreq4 & v39a5381 | !hbusreq4 & !v8455ab;
assign v37674a3 = hbusreq4 & v373ab15 | !hbusreq4 & v3a6b53f;
assign v37730ec = hlock5_p & v376d48b | !hlock5_p & v8455ab;
assign v372324a = hbusreq2 & v37251cc | !hbusreq2 & v8455ab;
assign v3759c9c = stateG10_1_p & v37457fb | !stateG10_1_p & !v3a63b56;
assign v37741f1 = hmaster2_p & v377c6b3 | !hmaster2_p & v3a68d2e;
assign v3731478 = hbusreq6_p & v376803b | !hbusreq6_p & v8455ab;
assign v3809ec3 = hgrant6_p & v8455ab | !hgrant6_p & v3765261;
assign v3765f60 = hgrant6_p & v8455ab | !hgrant6_p & v37240e6;
assign v37271fd = hgrant5_p & v376a8c8 | !hgrant5_p & v3a6f7d2;
assign v3a70074 = hgrant2_p & v8455ab | !hgrant2_p & v3744c9d;
assign v3a70585 = hmaster2_p & v3730e7d | !hmaster2_p & v3a6f8de;
assign v3746ab7 = hmaster0_p & v1e382e7 | !hmaster0_p & v3764d6b;
assign v3a5e7e0 = hlock7_p & v3754fc6 | !hlock7_p & !v3a6f58f;
assign v3a711e7 = hgrant6_p & v8455ab | !hgrant6_p & v37729c7;
assign v374b5da = hgrant6_p & v2acaf72 | !hgrant6_p & !c6598e;
assign v3a7102b = hlock0 & v3a635ea | !hlock0 & v3726505;
assign v3a55d2f = hbusreq3_p & v377aacd | !hbusreq3_p & v8455ab;
assign v3759ca7 = hbusreq6 & v37537ef | !hbusreq6 & v37372c9;
assign v1e373f8 = hmaster0_p & v3a620f1 | !hmaster0_p & v3a6fdbd;
assign v376d8d1 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v3a7162d;
assign v373bfea = hlock6 & v3a67b86 | !hlock6 & v3a6e3f0;
assign v39a5380 = hmaster2_p & v3a6890e | !hmaster2_p & v3778b19;
assign v3722eaf = hlock0_p & v372391f | !hlock0_p & v3729880;
assign v37620eb = hlock4 & v3748797 | !hlock4 & v3a6f2ad;
assign v3a570c0 = jx2_p & v3a59fd0 | !jx2_p & v3a7123c;
assign v3778e2d = hmaster1_p & v3734967 | !hmaster1_p & v3a5943e;
assign v375ecd5 = hbusreq2_p & v3737053 | !hbusreq2_p & !v8455ab;
assign v3800eea = hmaster2_p & v37496fa | !hmaster2_p & v376e041;
assign v3733a4c = jx0_p & v373e2f2 | !jx0_p & v3a5d065;
assign v377c723 = hgrant2_p & v3a709df | !hgrant2_p & v3777417;
assign v374eb9c = hbusreq8_p & v377f0fb | !hbusreq8_p & v3a6393d;
assign v376a662 = hbusreq8_p & v3a5b0f5 | !hbusreq8_p & v8455ab;
assign v3a5c5fc = hbusreq6_p & v3733e9e | !hbusreq6_p & v1e38224;
assign v37607d2 = hbusreq6_p & v3743d58 | !hbusreq6_p & v37609a6;
assign v3a6f3ad = hbusreq3 & v3730946 | !hbusreq3 & v3a70a88;
assign v3755019 = hburst1 & v3a64235 | !hburst1 & v3a6edfa;
assign v3724c25 = hbusreq4 & v3757c7f | !hbusreq4 & v3a5a807;
assign v3768f71 = hlock7_p & v37751bb | !hlock7_p & !v3736d1d;
assign v373e858 = hgrant6_p & v3a6f61e | !hgrant6_p & !v373228a;
assign v372b923 = hbusreq5 & v3a5565d | !hbusreq5 & v3a70f0d;
assign v3730a7b = hmaster1_p & v3a582ea | !hmaster1_p & v374bba3;
assign v374dbdf = hmaster1_p & v3771507 | !hmaster1_p & v3a543c5;
assign v376967e = hmaster0_p & v377f170 | !hmaster0_p & !v3a634eb;
assign v3760750 = hmaster2_p & v3a6f018 | !hmaster2_p & v374044c;
assign v3778d07 = hgrant6_p & v3a67403 | !hgrant6_p & v3a644ab;
assign v37710fb = hmaster2_p & v2acb5a2 | !hmaster2_p & !v3773fdc;
assign v3a6fe1c = hgrant5_p & v37575fd | !hgrant5_p & v377da41;
assign v374f768 = hmaster1_p & v377e089 | !hmaster1_p & v3765a1d;
assign v3765268 = hlock8_p & v3a6fc42 | !hlock8_p & v3a575e5;
assign v372a20b = hmaster2_p & v8455b0 | !hmaster2_p & v3a702c2;
assign v3a70364 = hbusreq4_p & v8455bb | !hbusreq4_p & v377e1f6;
assign v3a70172 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a641d5;
assign v3a71282 = hmaster2_p & v8455ab | !hmaster2_p & v3a603a1;
assign v3a5fc82 = hbusreq6_p & v3a635ea | !hbusreq6_p & v372348c;
assign v3749fc1 = hlock7 & v376daa7 | !hlock7 & v374f272;
assign v3a70393 = hgrant6_p & v37572df | !hgrant6_p & v3744458;
assign v3a6eb55 = hgrant0_p & v3a57f41 | !hgrant0_p & v3776a6e;
assign v3a56bd5 = hbusreq2_p & v374c671 | !hbusreq2_p & v8455b0;
assign v373c01a = hlock6_p & v372546e | !hlock6_p & v3773a45;
assign v3a5c3ba = hmaster2_p & v374813d | !hmaster2_p & v3752869;
assign c5b5f4 = hlock8_p & v2ff9190 | !hlock8_p & v372fe57;
assign v3757506 = hbusreq8 & v3a69910 | !hbusreq8 & v3766dc8;
assign v3725a06 = hgrant3_p & v3a6efc6 | !hgrant3_p & v3a6123a;
assign v37424a9 = hbusreq5_p & v37266df | !hbusreq5_p & !v375a2ff;
assign v373a7ab = hmaster0_p & v375eee3 | !hmaster0_p & v3a6c03d;
assign v3a5f030 = hmaster2_p & v8455ab | !hmaster2_p & !v3a56864;
assign v3a63d55 = hbusreq0 & v375df77 | !hbusreq0 & v37604b3;
assign v3a6fe76 = hmaster3_p & v3764099 | !hmaster3_p & v372ff96;
assign v3a6b2ea = hbusreq8_p & v3752248 | !hbusreq8_p & v3a70dfd;
assign v3745b5b = hgrant5_p & v372c0de | !hgrant5_p & !v373a4b2;
assign v3766a7d = hbusreq8_p & v374ef62 | !hbusreq8_p & v376d88f;
assign v37693ce = hmaster2_p & v8455ab | !hmaster2_p & !v3754aa3;
assign v3756b5c = hbusreq5 & v372b316 | !hbusreq5 & v3378fc3;
assign v374e9b8 = hbusreq6 & v8455cb | !hbusreq6 & v8455b3;
assign v3a60b37 = hbusreq5_p & v375d455 | !hbusreq5_p & v3761065;
assign v3764dda = hmaster0_p & v372edf8 | !hmaster0_p & v3a66e30;
assign v3a69bdc = hgrant5_p & v1e37daf | !hgrant5_p & v3a5b58e;
assign v373f684 = hmaster1_p & v37662ac | !hmaster1_p & v3728d9c;
assign v20930c2 = hgrant6_p & v91cdff | !hgrant6_p & v3a65e52;
assign v376b4d4 = hlock7 & v23fd9cb | !hlock7 & v373d239;
assign v3a6f9e6 = hlock5 & v3a7026d | !hlock5 & v3766acb;
assign v3a6e790 = hmaster0_p & v377c125 | !hmaster0_p & v37653d1;
assign v3a6b1d4 = hgrant4_p & v375c7b9 | !hgrant4_p & v375983d;
assign v37425a8 = hbusreq7 & v3a701fe | !hbusreq7 & a0a219;
assign v37772c0 = hbusreq5_p & v3766e62 | !hbusreq5_p & v8455e7;
assign v374bb9f = hmaster0_p & v3a70209 | !hmaster0_p & v3a70137;
assign v3756ce5 = hlock8 & v3a5e8ac | !hlock8 & v3a67d7b;
assign v3a70ffe = jx0_p & v3a6eafe | !jx0_p & v3749dc2;
assign v3a6f3f8 = hmaster1_p & v37795d3 | !hmaster1_p & v2093037;
assign v3a67c13 = hbusreq3_p & v3745f76 | !hbusreq3_p & v3a6fe90;
assign v377c17f = hbusreq1_p & v37598e6 | !hbusreq1_p & !v3a593e0;
assign c32250 = hbusreq3_p & v3752943 | !hbusreq3_p & v8455ab;
assign v374cbc4 = hmaster2_p & v3a70809 | !hmaster2_p & v37571c0;
assign v3771bb9 = hlock0_p & b254e2 | !hlock0_p & v375c541;
assign v3a5def7 = hmaster1_p & v3a608b8 | !hmaster1_p & v8455ab;
assign v3756577 = hbusreq5 & v373e6bc | !hbusreq5 & v8455ab;
assign v3754018 = hmaster0_p & v373ecb2 | !hmaster0_p & v94e9e0;
assign v372def9 = hbusreq5 & v3a7102f | !hbusreq5 & v360bc74;
assign v372b44a = hlock6 & v3a70ba7 | !hlock6 & v3a70ee1;
assign v373ae83 = hbusreq0 & v37522ff | !hbusreq0 & v376663a;
assign v3a70511 = hbusreq4 & v3a5c462 | !hbusreq4 & v373d10f;
assign v374bd4a = hbusreq5_p & v3752321 | !hbusreq5_p & v37404d0;
assign v3760a52 = hmaster2_p & v3a70374 | !hmaster2_p & v3a621e7;
assign v3a6f710 = hbusreq8_p & v3a6f7a6 | !hbusreq8_p & v8455ab;
assign v3738855 = hbusreq6_p & v3a70279 | !hbusreq6_p & v3a6a910;
assign v3a6fcb7 = hmaster0_p & v3735d6f | !hmaster0_p & !v3a70386;
assign v3771fb3 = hbusreq6_p & v3a6d951 | !hbusreq6_p & v372fa0f;
assign v3a670d6 = hbusreq3 & v3779fec | !hbusreq3 & v3a6ca99;
assign v3761fc1 = hbusreq2_p & v372e88a | !hbusreq2_p & v3a6f0a9;
assign v3759a88 = hgrant3_p & v3a6f53d | !hgrant3_p & !v3a5e09d;
assign v376b576 = hbusreq6_p & v3a5706c | !hbusreq6_p & v377894b;
assign v376e3db = hlock4_p & v3a7020b | !hlock4_p & v3a6fac6;
assign v3735906 = hbusreq6_p & v3727bca | !hbusreq6_p & v3737a29;
assign v375eff3 = hbusreq2 & v3a6fa5e | !hbusreq2 & v8455ab;
assign v373a101 = hbusreq2_p & v377abb1 | !hbusreq2_p & v373b42b;
assign v375f28d = hlock7 & v3a70676 | !hlock7 & v3a70c06;
assign v376348c = hbusreq6 & v3a70200 | !hbusreq6 & !v37413fc;
assign v373dd77 = hbusreq6_p & v3a70641 | !hbusreq6_p & v8455e7;
assign v37350b7 = hbusreq4_p & v3a5c945 | !hbusreq4_p & !v3a66110;
assign v373dc2f = stateG10_1_p & v376ba47 | !stateG10_1_p & v375cec6;
assign v3772c0a = hmaster0_p & v3a6e584 | !hmaster0_p & v8455e7;
assign v3a557a1 = hbusreq5_p & v373adaa | !hbusreq5_p & v374f533;
assign v3a6dae2 = hbusreq6_p & v374a4a0 | !hbusreq6_p & v375d22f;
assign v376158d = hgrant4_p & v35b774b | !hgrant4_p & v3735ea8;
assign v3725a2e = hbusreq5_p & v3a58016 | !hbusreq5_p & !v3744d2a;
assign v3748fde = hmaster2_p & afdeb4 | !hmaster2_p & v374bfcf;
assign v3a6b2e5 = hgrant2_p & v3a70403 | !hgrant2_p & v3756bb9;
assign v37777d2 = hbusreq3 & v3a58520 | !hbusreq3 & v8455ab;
assign v372a0f7 = hbusreq6 & v3a6fbd0 | !hbusreq6 & !v3a5538a;
assign v3750d46 = hbusreq4 & v3a539bb | !hbusreq4 & v3a635ea;
assign v3759a67 = hmaster0_p & v377234d | !hmaster0_p & v3743910;
assign v37524a6 = hbusreq2 & v3a6440f | !hbusreq2 & v3a6fefa;
assign v3a66ade = hgrant4_p & v3a5690d | !hgrant4_p & v3a6f647;
assign v372b0ac = hgrant1_p & v3a57445 | !hgrant1_p & v374e78f;
assign v3723fb3 = hmaster3_p & v375f1db | !hmaster3_p & v3a6f86f;
assign v376f718 = hmaster1_p & v3758cec | !hmaster1_p & v372ac19;
assign v3a6f1db = hbusreq7 & v90b307 | !hbusreq7 & v373556f;
assign v3758672 = hmaster2_p & v3749437 | !hmaster2_p & v3a6f4c7;
assign v3763668 = hbusreq2_p & v3745014 | !hbusreq2_p & !v8455ab;
assign v3775d04 = hlock6 & v372a6c2 | !hlock6 & v377aa23;
assign v375d924 = hbusreq4_p & v3a70488 | !hbusreq4_p & v3a64af7;
assign v3a68ef7 = hgrant4_p & v3a53eeb | !hgrant4_p & v37395f5;
assign v3a70e0f = hbusreq4 & v3a608b9 | !hbusreq4 & !v376b6c8;
assign v3739e21 = hbusreq8 & v3765b9b | !hbusreq8 & v37723c6;
assign v37536bf = hgrant4_p & v8455ab | !hgrant4_p & v3a70f11;
assign v377e9b0 = hlock5 & v377bb38 | !hlock5 & v37397ba;
assign v3809194 = hbusreq0 & v376a149 | !hbusreq0 & v3a67cd1;
assign v3726845 = hlock0_p & v3751734 | !hlock0_p & !v8455ab;
assign v3740db1 = hgrant6_p & v209310e | !hgrant6_p & !v1e37a26;
assign v372516b = hbusreq4_p & v3762f76 | !hbusreq4_p & v8455ab;
assign v372f006 = hmaster2_p & v3a6dfb2 | !hmaster2_p & v373be25;
assign v3a5398c = hmaster0_p & v3a60cd0 | !hmaster0_p & !v3771e23;
assign v3770769 = hbusreq6_p & v37406d2 | !hbusreq6_p & v372d0ad;
assign db3b98 = hgrant2_p & v8455b9 | !hgrant2_p & v375f0af;
assign v3778787 = hgrant6_p & v8455ab | !hgrant6_p & v3a62465;
assign v38099a4 = hmaster0_p & a1b632 | !hmaster0_p & v376df4c;
assign v3a708bc = jx0_p & v3a70acb | !jx0_p & v3776691;
assign v38093aa = hbusreq6 & v375911a | !hbusreq6 & v3a69487;
assign v375023c = jx3_p & v3a5f375 | !jx3_p & !v3808db7;
assign v3a6ff4f = hgrant6_p & v37722e5 | !hgrant6_p & v3a704ee;
assign v3a53e46 = jx1_p & v3a635eb | !jx1_p & v377c72c;
assign v3732187 = hbusreq4 & v37434ce | !hbusreq4 & v3725799;
assign v3744838 = hbusreq5 & v3761334 | !hbusreq5 & v3743fc1;
assign v372ab19 = hmaster2_p & v3a635ea | !hmaster2_p & v3a6f4c7;
assign v373195f = hgrant4_p & v8455ab | !hgrant4_p & v373869b;
assign v33789ca = hmaster1_p & v374a8da | !hmaster1_p & v8455ab;
assign v3758c50 = hgrant4_p & v8455ab | !hgrant4_p & v3a703d9;
assign v3730946 = hlock0_p & v3a5e9d3 | !hlock0_p & v372a399;
assign v3a6a5e6 = hmaster2_p & v3776649 | !hmaster2_p & !v8455ab;
assign v3a5df33 = hgrant5_p & v8455ab | !hgrant5_p & v377e904;
assign v3748656 = hmaster0_p & v3a62a68 | !hmaster0_p & v38088e1;
assign v8455d9 = hmaster0_p & v8455ab | !hmaster0_p & !v8455ab;
assign v372969d = jx1_p & v23fe142 | !jx1_p & v3746e54;
assign v3a6e81d = hmaster0_p & v373a0d6 | !hmaster0_p & v372f59c;
assign v37717d0 = hmaster0_p & v375808f | !hmaster0_p & v3a6ff25;
assign v373b1bb = hbusreq7 & v376e20f | !hbusreq7 & v3a60859;
assign v3a5c6f9 = hbusreq6_p & v3a7084e | !hbusreq6_p & v3732564;
assign v3a6d695 = hmaster1_p & v373014d | !hmaster1_p & v372d925;
assign v3a55fc6 = hbusreq6_p & v3a65241 | !hbusreq6_p & !v8455ab;
assign v3735354 = hbusreq3_p & v375da09 | !hbusreq3_p & !v8455ab;
assign v3a6f5a2 = hmaster0_p & v373b203 | !hmaster0_p & v3a5b071;
assign v3a58c00 = hlock7_p & v8455e7 | !hlock7_p & !v8455ab;
assign v35b708c = hbusreq8 & v3765a2e | !hbusreq8 & v3a6bb56;
assign v3806498 = hbusreq5 & v3764c7c | !hbusreq5 & v3730b15;
assign v3a71235 = hbusreq5 & v37246d9 | !hbusreq5 & v8455ab;
assign v3a5bc72 = hgrant5_p & v8455c6 | !hgrant5_p & v3765590;
assign v374c7f4 = hbusreq2_p & v3809adf | !hbusreq2_p & v39a537f;
assign v3723add = hmaster0_p & v3a6953d | !hmaster0_p & v8455ca;
assign v373f3b5 = hgrant6_p & v377bfc0 | !hgrant6_p & v3767266;
assign v373691d = hbusreq6 & v376f2f8 | !hbusreq6 & v8455ab;
assign v375647b = hmaster2_p & v376111d | !hmaster2_p & v37482f8;
assign v37638ef = hbusreq5_p & v3756beb | !hbusreq5_p & v37283c8;
assign v3a61d5b = hmaster0_p & v3a700b2 | !hmaster0_p & v376db27;
assign v374a0c5 = hbusreq4_p & v3738e72 | !hbusreq4_p & !v377586c;
assign v377559f = hbusreq5 & v3760bc2 | !hbusreq5 & !v3a64862;
assign v372f289 = hbusreq4_p & v37294d3 | !hbusreq4_p & !v3a62a13;
assign v373e76a = hlock0 & v3a6403e | !hlock0 & v372b858;
assign v374cb05 = hlock2 & v375021b | !hlock2 & v37383f6;
assign v374cb9e = hgrant4_p & v3726f57 | !hgrant4_p & v3755ec0;
assign v3a7012e = hbusreq0 & v3a6f6b4 | !hbusreq0 & !v375be12;
assign v3750a17 = hbusreq8_p & v373bca5 | !hbusreq8_p & v3a715f8;
assign v3729996 = hgrant4_p & v37604e9 | !hgrant4_p & v3a6fe21;
assign v376a14f = hready & v3a5d532 | !hready & v8455e7;
assign v377bd77 = hlock5_p & v3746c51 | !hlock5_p & v3a6a557;
assign v374e7b5 = hlock7_p & v3752348 | !hlock7_p & v3a5f439;
assign v375eb37 = hlock7_p & v375dbda | !hlock7_p & v377e5a6;
assign v37293c2 = hready_p & v3a6f459 | !hready_p & !v3776fae;
assign v3764809 = hbusreq0 & v3a67e79 | !hbusreq0 & v8455ab;
assign v37314fc = hgrant4_p & v8455ab | !hgrant4_p & v3a651fb;
assign v374ffd5 = hmaster0_p & v3736be5 | !hmaster0_p & !v373197c;
assign v3a65755 = hmaster1_p & v3a635ea | !hmaster1_p & v3733e1f;
assign v3a6efce = hlock2_p & v37494ee | !hlock2_p & !v8455ab;
assign v376196f = hmaster2_p & v376501e | !hmaster2_p & v3754dd0;
assign v377e004 = hmaster2_p & v38074c2 | !hmaster2_p & v3a56e63;
assign v374a23b = hbusreq4 & v3a63805 | !hbusreq4 & v8455ab;
assign v3775a8e = hbusreq5_p & v3742649 | !hbusreq5_p & v3729544;
assign v3a706ea = hmaster1_p & v3a61a7f | !hmaster1_p & v3761b23;
assign v3a709a6 = hbusreq6_p & v376e1c4 | !hbusreq6_p & v8455bf;
assign v37257f8 = hgrant0_p & v8455ab | !hgrant0_p & !v37398f3;
assign v3a651fb = hbusreq0 & v3a645b4 | !hbusreq0 & v3a6358e;
assign v37695c7 = hmaster0_p & v3a696a7 | !hmaster0_p & v372b7a8;
assign v375b5d6 = hbusreq8 & v3779c5d | !hbusreq8 & v373e4a7;
assign v3767dc1 = hlock5_p & v8455e7 | !hlock5_p & v3a672e6;
assign v3751dcc = hlock5 & v3a63f9a | !hlock5 & v3751e62;
assign v3755502 = hbusreq5_p & v3a70264 | !hbusreq5_p & !v3731fab;
assign v3739f84 = hgrant2_p & v37598dc | !hgrant2_p & !v3734f09;
assign v3a62654 = hbusreq2_p & v3a5561b | !hbusreq2_p & v3a5d0b6;
assign v37591f3 = hlock0 & v3a6c5ee | !hlock0 & v3a64b90;
assign v374c61d = hbusreq4 & v3771ab9 | !hbusreq4 & v376e041;
assign v3a67c50 = hmaster0_p & v376285a | !hmaster0_p & v3a7096f;
assign v37520ad = hmaster2_p & v376ef4f | !hmaster2_p & v1e37523;
assign v3768d6c = hbusreq5 & v373dde1 | !hbusreq5 & v373790d;
assign v3751f28 = hgrant3_p & v372ffd2 | !hgrant3_p & v3734256;
assign v3a63cf3 = hbusreq7 & v37470fc | !hbusreq7 & v8455ab;
assign v3807a93 = hmaster1_p & v8455ab | !hmaster1_p & v3a706da;
assign v377be72 = hmaster2_p & v373f6ee | !hmaster2_p & v3757c7f;
assign v375e70f = hlock7_p & v3764ca7 | !hlock7_p & !v8455ab;
assign v374d5fa = hmaster1_p & v372b9c5 | !hmaster1_p & v3a70f68;
assign v3768288 = hbusreq4 & v377e29a | !hbusreq4 & v3a654c1;
assign v3735444 = hbusreq4 & v3a627a7 | !hbusreq4 & v374d63f;
assign v3a676a9 = hgrant2_p & v3a6c63e | !hgrant2_p & v3a708b9;
assign v37313a7 = hgrant5_p & v38073ff | !hgrant5_p & v373da6d;
assign v375c7a9 = hbusreq4 & v3765ab2 | !hbusreq4 & v3737028;
assign v373150d = hbusreq8_p & v3759569 | !hbusreq8_p & v3750b64;
assign v374d80f = hlock4 & v377414c | !hlock4 & v37556ec;
assign v377aa06 = hgrant6_p & v8455c9 | !hgrant6_p & v3a5cbd8;
assign v374d183 = hbusreq6_p & v377cdee | !hbusreq6_p & v3a6fc54;
assign v3734fba = hbusreq5 & v3a63699 | !hbusreq5 & v3a63f9a;
assign stateG3_1 = !v2092c08;
assign v374d669 = hlock7_p & v3755066 | !hlock7_p & v3a70652;
assign v374d33d = hlock0 & v3749bf0 | !hlock0 & v3727c62;
assign v37420e2 = hlock4 & v3a6f69f | !hlock4 & v3731eff;
assign v3744b1b = hbusreq4_p & v372eafa | !hbusreq4_p & v3731596;
assign v37738be = hbusreq5 & v3a6512d | !hbusreq5 & v3775931;
assign v3a5bf56 = hbusreq7_p & v3a6beff | !hbusreq7_p & v8455ab;
assign v3a5c2d7 = hbusreq4 & v373399e | !hbusreq4 & v8455ab;
assign v94e000 = hgrant2_p & v3a53f43 | !hgrant2_p & v372d59e;
assign v3a56230 = hmaster0_p & v3a707cf | !hmaster0_p & v37653d1;
assign v376fb92 = hbusreq8 & v377d671 | !hbusreq8 & v8455c3;
assign v374a1f5 = hgrant4_p & v8455c2 | !hgrant4_p & v373ae0a;
assign v374335b = hbusreq8_p & v3a6ebdc | !hbusreq8_p & v3a70170;
assign v374c9c2 = hmaster0_p & v376b5a4 | !hmaster0_p & !v3739ea5;
assign v377312f = hmaster2_p & v3a5bd58 | !hmaster2_p & v3740dc6;
assign v376aaee = hlock5 & v3a70a89 | !hlock5 & v376d172;
assign v372f89e = hbusreq5_p & v37278fd | !hbusreq5_p & v3777f01;
assign v37244f3 = hmaster1_p & v37285fa | !hmaster1_p & v3a66a3a;
assign v377437d = hbusreq4_p & v37570f8 | !hbusreq4_p & v3a6fd3e;
assign v377e9bb = hbusreq0 & v3728f3a | !hbusreq0 & v374a3b8;
assign v374eb71 = hlock4_p & v3a703fc | !hlock4_p & !v8455ab;
assign v372342b = hbusreq0 & v37233a7 | !hbusreq0 & v3726739;
assign v3a5bda1 = hbusreq6_p & v3737d48 | !hbusreq6_p & v3a5bf99;
assign v3a6512d = hmaster0_p & v37564a2 | !hmaster0_p & v3754727;
assign v3a71072 = hbusreq5 & v3a6ef2c | !hbusreq5 & v380760a;
assign v3727f67 = hmaster0_p & v8455e7 | !hmaster0_p & v3743c45;
assign v37564d1 = hmaster2_p & v37651c2 | !hmaster2_p & v373a341;
assign v3a58eed = hgrant4_p & v23fde7c | !hgrant4_p & v3763c0a;
assign v377055c = hbusreq5_p & v23fd817 | !hbusreq5_p & v3770aa1;
assign v3731258 = hgrant0_p & v1e3791d | !hgrant0_p & v374a45c;
assign v3a698ab = hbusreq5 & v28896f0 | !hbusreq5 & v375d417;
assign v3756930 = hbusreq0 & v373577f | !hbusreq0 & v37718de;
assign v376071e = hbusreq2_p & v377de0d | !hbusreq2_p & v8455ab;
assign v3729187 = hmaster2_p & v3a70059 | !hmaster2_p & !v3a70fec;
assign v374dc13 = hgrant4_p & v372a71e | !hgrant4_p & v3a6d09c;
assign v3a6faac = hlock0_p & v3a54c77 | !hlock0_p & !v8455ab;
assign v37231ed = hbusreq0_p & v37787ec | !hbusreq0_p & v3a7162d;
assign v374880c = hbusreq4_p & v3738fe2 | !hbusreq4_p & v3742dce;
assign v372faf1 = hgrant0_p & v373dc1c | !hgrant0_p & ad2d05;
assign v372348c = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a63621;
assign v3732b98 = stateG10_1_p & v3a63621 | !stateG10_1_p & v3a7148d;
assign v375e993 = hmaster2_p & v3742f64 | !hmaster2_p & v8455ab;
assign v3724e98 = hgrant2_p & v8455ab | !hgrant2_p & v372a406;
assign v3a714f1 = hlock5 & v3a6c044 | !hlock5 & v374a157;
assign v3726c36 = hbusreq0_p & v3747302 | !hbusreq0_p & v3a71452;
assign v3776d97 = hbusreq6_p & v3777a52 | !hbusreq6_p & v372abc8;
assign v3728c14 = hmaster2_p & v376bade | !hmaster2_p & v376bb26;
assign v3778fa0 = hgrant6_p & v3a6eb39 | !hgrant6_p & v3749c91;
assign v3a6eb46 = hlock5 & v3a70c4b | !hlock5 & v372c3d7;
assign v3a710bc = hlock3_p & v376a4c0 | !hlock3_p & v2093059;
assign v3749dad = busreq_p & v3745536 | !busreq_p & v8455ff;
assign v3751c00 = jx1_p & v377a308 | !jx1_p & v375a2a7;
assign v372e27f = hgrant3_p & v9ed516 | !hgrant3_p & v37441b5;
assign v37481c3 = hmastlock_p & v3760ef5 | !hmastlock_p & !v8455ab;
assign v3a5a7c6 = hbusreq3_p & v3a6fe6a | !hbusreq3_p & v3a703df;
assign v3a647e3 = hgrant6_p & v37418ac | !hgrant6_p & v3754e70;
assign v3a703d1 = hburst0 & v373d9e5 | !hburst0 & v377ac6f;
assign v374333e = hlock5 & v372b923 | !hlock5 & v3a5565d;
assign v3731e7b = hbusreq2_p & v3a70641 | !hbusreq2_p & v8455e7;
assign v1e37583 = decide_p & v3a70069 | !decide_p & v3732aab;
assign v38090f4 = hgrant6_p & v8455b0 | !hgrant6_p & v3a56dd5;
assign v3a7082d = hgrant4_p & v3a6a22c | !hgrant4_p & v3a6fd34;
assign v3a5988f = hgrant2_p & v3a5b12c | !hgrant2_p & v376278c;
assign v3740e8d = hlock8_p & v376297b | !hlock8_p & v375c99d;
assign v3a5e667 = hlock0 & v3748797 | !hlock0 & v3736b57;
assign v375ecf5 = hbusreq6_p & v3749586 | !hbusreq6_p & v3a60882;
assign v3a58a3b = hbusreq7 & v375372b | !hbusreq7 & v3772cab;
assign v377e442 = hbusreq5_p & v8455bf | !hbusreq5_p & v377bcb3;
assign v374f003 = hbusreq8_p & v3a62959 | !hbusreq8_p & v3752552;
assign v3a617b4 = hlock0_p & v37665bf | !hlock0_p & v8455e7;
assign v3a70957 = hgrant4_p & v3733e9e | !hgrant4_p & v3a71012;
assign v3766e62 = hbusreq5 & v37308bc | !hbusreq5 & v8455e7;
assign v3a63def = hlock5_p & v376fd33 | !hlock5_p & v37767d7;
assign v374ffb7 = hbusreq6_p & v3a635ea | !hbusreq6_p & v377629f;
assign v3779cb7 = hbusreq2_p & v377b1db | !hbusreq2_p & v8455ab;
assign v3a6540f = hmaster1_p & v375ac26 | !hmaster1_p & v3a6ec22;
assign v3806dc8 = hbusreq7_p & v37295a5 | !hbusreq7_p & !v1e37759;
assign v373c334 = hmaster1_p & v3a705d4 | !hmaster1_p & v3a6dcf3;
assign v3a566c0 = hbusreq5_p & v3740614 | !hbusreq5_p & v3a58c07;
assign v373d7ea = hlock0 & v3768751 | !hlock0 & v3a70ff1;
assign v375eef1 = hbusreq3 & v39a5265 | !hbusreq3 & !v376f665;
assign v3a70655 = hlock7_p & v374cb02 | !hlock7_p & v3a6cc5f;
assign v3753198 = hmaster3_p & v37350e9 | !hmaster3_p & v3766830;
assign v375ee2a = hgrant6_p & v3a6ab8c | !hgrant6_p & ce82b0;
assign v3809fbb = hbusreq7 & v3773098 | !hbusreq7 & v3a6fc5d;
assign v37316f2 = hbusreq5_p & v3756012 | !hbusreq5_p & v3a6eb21;
assign v3a5bf21 = hlock5_p & v8455ab | !hlock5_p & !v3a63d83;
assign v3a6fdcc = hbusreq0 & v3758ff4 | !hbusreq0 & v377c31d;
assign v23fe189 = hgrant2_p & v37691fa | !hgrant2_p & v3a70624;
assign v3a6a0c4 = hbusreq7 & v3755f2d | !hbusreq7 & v8455ab;
assign v3a6f4bd = hmaster2_p & v8455ab | !hmaster2_p & v3a703c5;
assign v374b73b = hbusreq6 & v3732564 | !hbusreq6 & v37443ab;
assign v375b676 = hbusreq8 & v375f848 | !hbusreq8 & v373c7af;
assign v3744a56 = hmaster2_p & v3a5fe9e | !hmaster2_p & v3a67d2f;
assign v3a6fc41 = hmaster0_p & v3a6fd7e | !hmaster0_p & !v3a634eb;
assign v3a655a3 = hbusreq2_p & v3723f24 | !hbusreq2_p & v37c0077;
assign v3724e45 = hmaster2_p & v377169f | !hmaster2_p & v3732415;
assign v376fe45 = hmaster0_p & v37774d3 | !hmaster0_p & d8c443;
assign v3a70cc2 = hgrant2_p & v3a6ec1e | !hgrant2_p & v8455ab;
assign v3a6f908 = hlock4 & v3a6a346 | !hlock4 & v3a6f20f;
assign v377dbdc = hbusreq8_p & v3a6fbc4 | !hbusreq8_p & v3a59c72;
assign v373ab3d = hlock8_p & v8455ab | !hlock8_p & v372667b;
assign v3a696a7 = hgrant4_p & v3a637dc | !hgrant4_p & v37373af;
assign v372879d = hmaster2_p & v3a62a6d | !hmaster2_p & v377097a;
assign v3728f66 = hmaster1_p & v8455ab | !hmaster1_p & v3748829;
assign v3a6fa77 = hmaster0_p & v3773708 | !hmaster0_p & v37341d3;
assign v3a6eedf = hmaster1_p & v3765008 | !hmaster1_p & v8455ab;
assign v3a702bc = hlock2 & v373e962 | !hlock2 & v3742d54;
assign v3764efe = hbusreq2 & v374f307 | !hbusreq2 & v8455ab;
assign v3773ca3 = hmaster2_p & v3a6abf7 | !hmaster2_p & v377047a;
assign v377b94f = hbusreq6_p & v3725947 | !hbusreq6_p & v8455ab;
assign v3727fe3 = stateG2_p & v8455ab | !stateG2_p & v3738cfc;
assign v3a6f39b = hbusreq6 & v3809ebc | !hbusreq6 & v3738510;
assign v3741abc = hmaster1_p & v3a6f868 | !hmaster1_p & v8455ab;
assign v3a61280 = hmaster0_p & v373eba7 | !hmaster0_p & v3776c95;
assign v3a65b79 = hbusreq5_p & v375c4e0 | !hbusreq5_p & v375a688;
assign v3a70aa6 = hmaster1_p & v2093252 | !hmaster1_p & !v376256f;
assign v3a70feb = hbusreq5 & v3a58527 | !hbusreq5 & v3758661;
assign v374ac60 = hbusreq0 & v3a6f496 | !hbusreq0 & v8455ab;
assign v3761300 = hmaster2_p & v372625f | !hmaster2_p & v3772e0c;
assign v3732bd2 = hbusreq0 & v37652f1 | !hbusreq0 & v3775725;
assign v3729544 = hlock5 & v3735ac0 | !hlock5 & v376fbe3;
assign v39a4e99 = hbusreq5_p & v377a18b | !hbusreq5_p & v377e056;
assign v3a6f2d4 = hbusreq6_p & v376c6ed | !hbusreq6_p & v3771f9b;
assign v372d70c = hmaster1_p & v374db48 | !hmaster1_p & v3a6fcb8;
assign v37318e2 = hlock0 & v3808952 | !hlock0 & v3a57ac7;
assign v3a7048d = hbusreq4 & v372b5f5 | !hbusreq4 & v8455ab;
assign v375898f = hlock0_p & v35772b3 | !hlock0_p & v35772a6;
assign v3a6fd48 = hgrant3_p & v3a70544 | !hgrant3_p & v3a623c7;
assign v374b4c5 = hmaster1_p & v3a55466 | !hmaster1_p & v8455ab;
assign v376e9ed = hgrant5_p & v376e66e | !hgrant5_p & v3a62fc9;
assign v3a5a5c4 = hmaster1_p & v372c0cc | !hmaster1_p & v376d896;
assign v3a6fc3f = hmaster2_p & v3a6fc74 | !hmaster2_p & v3754b03;
assign v23fe20c = hbusreq5_p & v3a705df | !hbusreq5_p & v3a57c78;
assign v375dcf5 = hgrant6_p & v8455ca | !hgrant6_p & v3739460;
assign v1e37916 = hbusreq8 & v3747917 | !hbusreq8 & v376ae9f;
assign v3a6f83b = hbusreq7 & v373c4a7 | !hbusreq7 & v3737808;
assign v376498f = hbusreq6_p & v3747302 | !hbusreq6_p & v3a70a88;
assign v3a67c3b = hmaster2_p & v3a635ea | !hmaster2_p & v375cf36;
assign v375e47e = hgrant6_p & v3777996 | !hgrant6_p & v37786a4;
assign v3a6e7ce = hbusreq5_p & v3a6d874 | !hbusreq5_p & v375dd02;
assign v3a70a0e = hbusreq6 & v37485c0 | !hbusreq6 & v373c965;
assign v37664f6 = hlock1_p & v8455ab | !hlock1_p & !v2acb5a2;
assign v3a70ad0 = hmastlock_p & v3a6e78d | !hmastlock_p & v8455ab;
assign v372f49f = hmaster1_p & v3a70528 | !hmaster1_p & v3754025;
assign v3766315 = hgrant2_p & v8455ba | !hgrant2_p & v375ebdd;
assign v3a6f07f = hmaster0_p & v37720ce | !hmaster0_p & !v3a6ebac;
assign v37645a8 = hbusreq3_p & v3a67eec | !hbusreq3_p & v3743b9e;
assign v373b88a = hgrant6_p & v374c70d | !hgrant6_p & v3769010;
assign v372864a = hbusreq6 & v3737075 | !hbusreq6 & v3776e85;
assign v37356d4 = hbusreq0_p & v8455b0 | !hbusreq0_p & v8455ab;
assign v3a70463 = hmaster2_p & v3755252 | !hmaster2_p & !v373c21c;
assign v3a5c85c = hgrant4_p & v376c484 | !hgrant4_p & v37686f3;
assign v3753429 = hbusreq4_p & v3755f9b | !hbusreq4_p & !v3752c4d;
assign v3a54e47 = hgrant5_p & v37463ef | !hgrant5_p & v3a71093;
assign v3736257 = hbusreq7 & v3a6e552 | !hbusreq7 & v3748c3f;
assign v372c713 = hbusreq6 & v373e9a5 | !hbusreq6 & v3a716a3;
assign v3726b90 = hmaster2_p & v376142a | !hmaster2_p & v8455ab;
assign v376314e = hbusreq5_p & v372c0fd | !hbusreq5_p & v3a6fac1;
assign v37314db = hmastlock_p & v373d2e0 | !hmastlock_p & !v8455ab;
assign v3a6500c = hgrant0_p & v3a6ebf6 | !hgrant0_p & v374059d;
assign v3751dc9 = hlock3 & v3a6eecd | !hlock3 & v377857d;
assign v375401a = hbusreq0_p & v8455ab | !hbusreq0_p & v3a6f656;
assign v372f5e5 = hbusreq8 & v3722bfc | !hbusreq8 & v3808dcb;
assign v3a70ff4 = hmaster0_p & v377234d | !hmaster0_p & v1e37bb4;
assign v3756c83 = hbusreq4 & v373fe6f | !hbusreq4 & v373031f;
assign v376005f = hgrant2_p & v3808ed4 | !hgrant2_p & v376441d;
assign v373804d = hlock7 & v37487a6 | !hlock7 & v3a6f1b9;
assign v372e440 = jx0_p & v8455ab | !jx0_p & v3a6f72e;
assign v373e6f1 = hbusreq6_p & v377e2f7 | !hbusreq6_p & v38095b2;
assign v3a7066c = hgrant4_p & v374306c | !hgrant4_p & v37297f4;
assign v373a54d = hmaster2_p & v375121b | !hmaster2_p & v3745a5f;
assign v3a6f9b4 = hlock7 & v373dd40 | !hlock7 & v3a63688;
assign v372fb2a = hbusreq4_p & v3728ee0 | !hbusreq4_p & !v8455ab;
assign v373a26b = hbusreq5_p & v37276d6 | !hbusreq5_p & !v3a706c1;
assign v3a6f437 = hbusreq7 & v3a6ecb7 | !hbusreq7 & v3809142;
assign v372bf87 = hgrant3_p & v3a68aa8 | !hgrant3_p & v376bad8;
assign v3a613f4 = hbusreq4_p & v3a6431f | !hbusreq4_p & !v3772827;
assign v3a6fa6e = hbusreq3 & v3725410 | !hbusreq3 & v3a706d1;
assign v37c033d = hgrant4_p & v8455e7 | !hgrant4_p & v375c845;
assign v3a59c21 = hbusreq5 & v374fde8 | !hbusreq5 & !v373bcdd;
assign v375c2d0 = hmaster1_p & v8455ab | !hmaster1_p & !v3746fcb;
assign v3a57c2a = hgrant2_p & v3773e41 | !hgrant2_p & !v3a660e9;
assign v37283c0 = hmaster2_p & v3725410 | !hmaster2_p & v8455ab;
assign v3730b8c = hbusreq5_p & v373a7ab | !hbusreq5_p & v3a6c09f;
assign v373bd3d = hmaster0_p & v37245f8 | !hmaster0_p & v3745186;
assign v376a4dd = hgrant2_p & v37443ab | !hgrant2_p & v3757fcc;
assign v3a58057 = hbusreq6_p & v372c614 | !hbusreq6_p & v8455ab;
assign v3765021 = hlock4 & v3a6fd4b | !hlock4 & v37659e2;
assign v376230d = hbusreq8 & v374d03f | !hbusreq8 & v3a6b798;
assign v3a560b8 = hmaster2_p & v372391f | !hmaster2_p & !v375641f;
assign v3770bed = hbusreq4 & v3774000 | !hbusreq4 & v8455ab;
assign v3728b10 = hlock5 & v377d491 | !hlock5 & v3a6f6ea;
assign v3770ee9 = hmaster2_p & v37737aa | !hmaster2_p & v8455ab;
assign v3722f37 = start_p & v8455d5 | !start_p & !v8455ab;
assign v373fb1a = hmaster1_p & v3a635ea | !hmaster1_p & v373f6cf;
assign v374c190 = hbusreq5 & v3722dcd | !hbusreq5 & v3a70971;
assign v3a5fa29 = hmaster1_p & v3752428 | !hmaster1_p & v3727bd4;
assign v373933b = hgrant6_p & v3a6ab8c | !hgrant6_p & v3a702ff;
assign v372c503 = hbusreq2 & v373399e | !hbusreq2 & v8455ab;
assign d5e2c2 = hmaster1_p & v3779060 | !hmaster1_p & v3731866;
assign v3a70446 = hgrant4_p & v3749c4b | !hgrant4_p & !v3a6d096;
assign v3a5c42c = hbusreq5_p & v372e443 | !hbusreq5_p & v3757b16;
assign v3a7166e = hbusreq5_p & v3726ddb | !hbusreq5_p & !v8455ab;
assign v374cdc4 = hmaster2_p & v3807aa1 | !hmaster2_p & !v3a70059;
assign v3774629 = hmaster3_p & v3769f60 | !hmaster3_p & !v374c63d;
assign v373b5d8 = hbusreq2_p & v3a70893 | !hbusreq2_p & v373cd16;
assign v3a7050a = hmaster1_p & v375841a | !hmaster1_p & v8455ab;
assign a94d63 = hmaster0_p & v3760592 | !hmaster0_p & v8455ab;
assign v376428f = hbusreq4_p & v3768076 | !hbusreq4_p & !v374c0e3;
assign v3770234 = hgrant6_p & v3745f9b | !hgrant6_p & v3577376;
assign v3a56e5e = hbusreq3 & v3a66e91 | !hbusreq3 & v38072fd;
assign v372f37d = hgrant6_p & v3759032 | !hgrant6_p & v3a70970;
assign v375fbbb = hbusreq4_p & v3777a00 | !hbusreq4_p & v8455ab;
assign v3767cc9 = hbusreq4_p & v3a6499e | !hbusreq4_p & !v8455ab;
assign v3a53ffa = hgrant6_p & v376e914 | !hgrant6_p & v3a6c835;
assign v374e0a4 = hmaster0_p & v37560b4 | !hmaster0_p & v3a68848;
assign v3a69430 = hbusreq4 & v377abd6 | !hbusreq4 & !v8455b5;
assign v373ad3c = hbusreq1_p & v3747302 | !hbusreq1_p & v3740646;
assign v3a6e6e1 = hbusreq6 & v37626a4 | !hbusreq6 & v3739da7;
assign v37689be = hmaster0_p & v377e16a | !hmaster0_p & v3a6eebb;
assign v376faf6 = hmaster0_p & v3a67899 | !hmaster0_p & !v8455bf;
assign v374478f = hmaster0_p & v3a70407 | !hmaster0_p & v3a6be79;
assign v3736fb6 = hmaster2_p & v374ab22 | !hmaster2_p & v376fb60;
assign v375918d = hbusreq5_p & v3744efc | !hbusreq5_p & v3a55d64;
assign v3a650bb = hbusreq0 & v3762a9c | !hbusreq0 & !v37740f9;
assign v3726e48 = hmaster0_p & v8455ab | !hmaster0_p & v3767985;
assign v3806882 = hmaster2_p & v39eb4ab | !hmaster2_p & v375995f;
assign v3a5d74e = hburst1 & v376c211 | !hburst1 & v3a65a34;
assign v375fcac = hbusreq7_p & v3a71254 | !hbusreq7_p & v37262ec;
assign v3759664 = jx3_p & v3760912 | !jx3_p & v3a6ff62;
assign v375c903 = hgrant4_p & v376e041 | !hgrant4_p & v3a5e2e1;
assign v37733f9 = hbusreq0 & v3760a2c | !hbusreq0 & v3727347;
assign v3741435 = hbusreq5 & v3763f95 | !hbusreq5 & v8455ab;
assign v372cb9d = hmaster2_p & v3a619c0 | !hmaster2_p & v375de18;
assign v3738d43 = hgrant6_p & v376a3ca | !hgrant6_p & v3757ec8;
assign v3758915 = hlock4 & v3a70c7f | !hlock4 & v373b78b;
assign v3a70936 = hmaster0_p & v3732f54 | !hmaster0_p & !v375f664;
assign v3779a80 = hbusreq5 & v3a70dd3 | !hbusreq5 & v3a6edb5;
assign v375f0f0 = hmaster1_p & v3a5e24e | !hmaster1_p & v3774542;
assign v3a62a51 = hgrant6_p & v8455ab | !hgrant6_p & v3747552;
assign v374dfad = hlock5_p & v3779477 | !hlock5_p & v372dd98;
assign v3a6faed = hmaster1_p & v8455ab | !hmaster1_p & !v1e37d14;
assign stateA1 = !v1e37583;
assign v3772b2b = hbusreq2_p & v377dabc | !hbusreq2_p & v3a6ef1f;
assign v3a6ec1f = hgrant6_p & v3a70b74 | !hgrant6_p & v8455ab;
assign v3745df8 = hbusreq6_p & v3726d2a | !hbusreq6_p & v373867c;
assign v952f44 = hbusreq5 & v8455ab | !hbusreq5 & v3733174;
assign v90a00a = locked_p & v8455ab | !locked_p & !v39ebac7;
assign v376fddd = hmaster3_p & v3730e4c | !hmaster3_p & v3a57311;
assign v37685f1 = hgrant5_p & v3809af2 | !hgrant5_p & v3a70419;
assign v373d9aa = hgrant0_p & v8455ab | !hgrant0_p & !v37682c6;
assign v3731d69 = hbusreq3_p & v377eaf2 | !hbusreq3_p & v3778528;
assign v3778572 = hbusreq4 & v39a4f09 | !hbusreq4 & v372ae6a;
assign v3725dd5 = hbusreq7 & v3749106 | !hbusreq7 & v3a6b31c;
assign v377a4e5 = hmaster1_p & v3a6ef47 | !hmaster1_p & v373c437;
assign v377e05a = hbusreq2_p & v372f012 | !hbusreq2_p & !v8455ab;
assign v375994d = hgrant5_p & v3755786 | !hgrant5_p & !v8455ab;
assign v373b11a = hgrant4_p & v8455ab | !hgrant4_p & v3762d6e;
assign cc809f = hbusreq1 & v37674c1 | !hbusreq1 & !v8455ab;
assign v3a7018b = hmaster2_p & v8455ab | !hmaster2_p & v3728e09;
assign v376fdd4 = hmaster1_p & v374e4fa | !hmaster1_p & v3a6f4da;
assign v37360d1 = hgrant4_p & v3772b7e | !hgrant4_p & v3763e44;
assign v3755aae = hmaster0_p & v3735e84 | !hmaster0_p & be0e1a;
assign v3764a2c = hmaster0_p & v3730553 | !hmaster0_p & v3a6f291;
assign v3722f3b = hgrant2_p & v372493b | !hgrant2_p & v374cc7f;
assign v3a7110d = hmaster0_p & v374d313 | !hmaster0_p & v8455ab;
assign v3a6d9a6 = hmaster0_p & v3731857 | !hmaster0_p & v38071bb;
assign v375571d = hbusreq4_p & v9684f8 | !hbusreq4_p & v8455e7;
assign v3a6b478 = hgrant8_p & v3741fea | !hgrant8_p & v377e89a;
assign v375a16a = hbusreq5 & v3a6ba91 | !hbusreq5 & v377326a;
assign v3773048 = hbusreq2_p & d44200 | !hbusreq2_p & !v3a7151d;
assign v3759bdb = hmaster0_p & v3a6f6ec | !hmaster0_p & !v373aec4;
assign v3726905 = hbusreq4 & v3767437 | !hbusreq4 & v8455b3;
assign v377cc27 = hlock2 & v3a712da | !hlock2 & v3a66d50;
assign v2ff8e74 = hbusreq5 & v3745202 | !hbusreq5 & v374e016;
assign v3a59a2b = hmaster0_p & v8455ab | !hmaster0_p & !v374f820;
assign v374c6de = hbusreq8 & v3806f1f | !hbusreq8 & v8455ab;
assign v3763d79 = hbusreq4_p & v3778921 | !hbusreq4_p & v3769945;
assign v3727171 = jx1_p & v375bce2 | !jx1_p & v3a7154d;
assign v372de6f = hmaster0_p & v372647d | !hmaster0_p & v374bd2c;
assign v3a6fdd6 = hbusreq2_p & v372e6ee | !hbusreq2_p & v8455ab;
assign v37390d6 = hmaster2_p & v3a635ea | !hmaster2_p & v3a70c74;
assign v372a6c8 = hmaster0_p & v37771ed | !hmaster0_p & v374000d;
assign v3a6fafd = hbusreq4_p & v3a62a6d | !hbusreq4_p & v3a70b17;
assign v3a6ec03 = hgrant6_p & v8455ab | !hgrant6_p & v3778962;
assign v375c278 = hmaster2_p & v3a5f413 | !hmaster2_p & v374cbc0;
assign v375603c = hgrant2_p & v37346be | !hgrant2_p & !v377cc25;
assign v3747e1f = hmaster2_p & v377955b | !hmaster2_p & v372d905;
assign v3766b48 = hbusreq4_p & v3a6fb2b | !hbusreq4_p & v3a6c9ab;
assign v375016d = hbusreq5 & v374fde8 | !hbusreq5 & !v3a6f40a;
assign v3767059 = hmaster1_p & v8455ab | !hmaster1_p & v375f354;
assign v3730398 = hmaster2_p & v3a70ab0 | !hmaster2_p & v8455ab;
assign v377652b = hbusreq6 & v3a5e7fe | !hbusreq6 & v8455bb;
assign v377a681 = hmaster1_p & v3731beb | !hmaster1_p & v3761bd6;
assign v3a60dd5 = hmaster0_p & v3807f45 | !hmaster0_p & v376eaf1;
assign v3a6b7e9 = hbusreq4_p & v3a70778 | !hbusreq4_p & v3a6c2a9;
assign v375469c = hmaster2_p & v3a55773 | !hmaster2_p & v8455ab;
assign v376d8fd = hlock5_p & v375ac09 | !hlock5_p & !v3757cd1;
assign v37435f6 = hbusreq3_p & v37311d6 | !hbusreq3_p & !v8455e9;
assign v374ac78 = hbusreq5 & v3a57baa | !hbusreq5 & v375f906;
assign v372386d = hgrant4_p & v3a65e3c | !hgrant4_p & v3751359;
assign v3762640 = hmaster1_p & v375ce8d | !hmaster1_p & v3a70601;
assign v1e37dcd = hmaster0_p & v3a6a516 | !hmaster0_p & !v3a70cab;
assign v3777573 = hgrant6_p & v37346be | !hgrant6_p & v375603c;
assign v373ec4c = jx1_p & v380a20c | !jx1_p & v3a56abc;
assign v37430f5 = hmaster0_p & v372b1dc | !hmaster0_p & v37638de;
assign v372b29d = hbusreq5_p & v8455e7 | !hbusreq5_p & !v8455ab;
assign v3a2a0e9 = hbusreq8 & v374fdeb | !hbusreq8 & v3779e29;
assign v3a663dd = hmaster1_p & v372998e | !hmaster1_p & !v3779ac0;
assign v3a53f1c = hmaster3_p & v376ba96 | !hmaster3_p & v3a705d0;
assign v3727a6b = hbusreq8_p & v3a65ce5 | !hbusreq8_p & v375c7c4;
assign v373588a = hbusreq3 & v37348ee | !hbusreq3 & v3a69487;
assign v3759387 = hgrant4_p & v3739ddf | !hgrant4_p & v3a70e0c;
assign v375f30d = hgrant0_p & v8455ab | !hgrant0_p & v3760af0;
assign v375f2f2 = hmaster2_p & v3a6f07d | !hmaster2_p & v3a70a51;
assign v37402d8 = hmaster2_p & v3a70a88 | !hmaster2_p & v374acbe;
assign v3a636d9 = hbusreq6 & v37496d3 | !hbusreq6 & v3a56e79;
assign v3740ab8 = hmaster2_p & v37367a0 | !hmaster2_p & !v376e854;
assign v3734c16 = hbusreq8_p & v3759569 | !hbusreq8_p & v3a6af5b;
assign v374608b = hmaster1_p & v3a63ea7 | !hmaster1_p & v373abd0;
assign v2acaeee = hmaster1_p & v3a66667 | !hmaster1_p & v3728d9c;
assign v3a5948f = hlock5_p & v373862e | !hlock5_p & v3a67471;
assign v3a715eb = hgrant5_p & v3a6f55a | !hgrant5_p & v3725269;
assign v372bd2b = hbusreq5_p & v3807dc9 | !hbusreq5_p & v8455ab;
assign v3a56642 = hbusreq3_p & v3a5a5ec | !hbusreq3_p & v8455ab;
assign v3a6f6bc = hbusreq5_p & v8455ab | !hbusreq5_p & v3a5f41b;
assign v37688bf = hmaster2_p & v375bf9a | !hmaster2_p & v8455ab;
assign v377a352 = hmaster2_p & v3741384 | !hmaster2_p & v37273d2;
assign v372b7e5 = hbusreq3_p & v3776615 | !hbusreq3_p & v37447bf;
assign v37353c6 = stateA1_p & v37440c3 | !stateA1_p & !v38073d4;
assign v3a5c0ac = hgrant6_p & v376a88b | !hgrant6_p & !v374c801;
assign v3726357 = hmaster0_p & v3731b90 | !hmaster0_p & v373197c;
assign v374d1ad = hgrant5_p & v3a62a2d | !hgrant5_p & v372f71f;
assign v3a56ebd = hmaster0_p & v374216a | !hmaster0_p & v8455ab;
assign v3a6f526 = hmaster1_p & v3a5877f | !hmaster1_p & v3a6c38a;
assign v375648e = hbusreq4_p & v3754aa3 | !hbusreq4_p & v375aaca;
assign v360d03b = hgrant0_p & v376969b | !hgrant0_p & v3a5ca02;
assign v37596a6 = hlock7 & v375f0de | !hlock7 & v3a6f873;
assign v374c2aa = hmaster1_p & v3a62a6d | !hmaster1_p & v3a6fd2f;
assign v3a6c390 = hbusreq2_p & v3a70cd3 | !hbusreq2_p & v3757fcc;
assign v37609a8 = hmaster2_p & v8455ab | !hmaster2_p & v372a4c1;
assign v3742b9d = hmaster2_p & v3759031 | !hmaster2_p & v3a687be;
assign v376e74b = hmaster0_p & v3763b5d | !hmaster0_p & v372f59c;
assign v376999f = hbusreq4_p & v3769ae2 | !hbusreq4_p & v3a538b4;
assign v3a70207 = hmaster3_p & v8455ab | !hmaster3_p & v377d51d;
assign v3a70096 = hgrant4_p & v3a5e544 | !hgrant4_p & v3776d7d;
assign v377073b = hmaster1_p & v3a5dbd7 | !hmaster1_p & v3a70924;
assign v377e0d2 = hmaster2_p & v3a539ae | !hmaster2_p & v3a5fff6;
assign v3a64d8f = hbusreq5 & v3a64082 | !hbusreq5 & v375240c;
assign v372dd77 = hmaster1_p & v3a5fae2 | !hmaster1_p & v3743f5b;
assign v374b0a9 = hbusreq6_p & v3a5b7b5 | !hbusreq6_p & v3732cb4;
assign v3a66c6c = hlock4 & v3a6fd4b | !hlock4 & v374ad67;
assign v3750ae0 = hmaster0_p & v3722dfe | !hmaster0_p & v372f997;
assign v374b972 = hmaster1_p & v372be74 | !hmaster1_p & v8455ab;
assign v3a706a3 = hlock8 & v3741fee | !hlock8 & v372a6de;
assign v3a654c4 = hgrant3_p & v37331e7 | !hgrant3_p & v372ae0b;
assign v373a438 = hmaster1_p & v3a5bf28 | !hmaster1_p & v376d89f;
assign v39ebaee = hlock7 & v376e68d | !hlock7 & v3a6ff0e;
assign v3a6fd4f = hlock5 & v3732b92 | !hlock5 & v1e37cba;
assign v376e9e9 = hgrant4_p & v8455ab | !hgrant4_p & v3779f43;
assign v3a65540 = hbusreq5_p & v3726594 | !hbusreq5_p & !v3a619c0;
assign v373f1ba = hgrant5_p & v8455ab | !hgrant5_p & !v3a70e2d;
assign v375bd0e = hgrant6_p & v8455ab | !hgrant6_p & v3a5b6c5;
assign v375af98 = hbusreq0 & v3729022 | !hbusreq0 & !v8455ab;
assign v3a5a1ff = hgrant3_p & v3a682b1 | !hgrant3_p & v3a70b08;
assign v372538e = hbusreq3_p & v375d7b6 | !hbusreq3_p & v37504b9;
assign a53cf9 = hbusreq4 & v375e12d | !hbusreq4 & v3765e79;
assign v3809f65 = hbusreq3_p & v3a5e591 | !hbusreq3_p & v8455b3;
assign v3768726 = hbusreq3_p & v37528b9 | !hbusreq3_p & v3a6f1a4;
assign v3a6cb50 = hlock3_p & v375c0cb | !hlock3_p & v3a59b5c;
assign v37624a2 = hbusreq1_p & v2acaef3 | !hbusreq1_p & v8455ab;
assign v373da69 = hbusreq1_p & v3766452 | !hbusreq1_p & !v37606c7;
assign d44200 = hready & v3a68f62 | !hready & v8455ab;
assign v3a70749 = hgrant6_p & v3a69de7 | !hgrant6_p & v3a635ea;
assign v374e0b8 = hmaster0_p & v377d1dc | !hmaster0_p & v3765dbc;
assign v3773b0f = hmaster0_p & v3a61397 | !hmaster0_p & v37377c8;
assign v3750ff0 = hlock5 & v3a64e3e | !hlock5 & v3a6d2d7;
assign c61b3c = hlock6_p & v3750d37 | !hlock6_p & !v8455ab;
assign v376a464 = hbusreq4 & v372e8cc | !hbusreq4 & v374617d;
assign v959f2d = hmaster1_p & v3a70fd5 | !hmaster1_p & v3735050;
assign v373e0d0 = hbusreq5_p & v37641b8 | !hbusreq5_p & v372cd61;
assign v3a71435 = hbusreq5 & v375121b | !hbusreq5 & !v8455c2;
assign v3a56e79 = hlock6_p & v377b774 | !hlock6_p & v8455bf;
assign v373d1bb = hbusreq6_p & v376c635 | !hbusreq6_p & v372b22b;
assign v3a62d82 = hmaster2_p & v377d142 | !hmaster2_p & v3730e98;
assign v23fdbe3 = hmaster0_p & v3a5865e | !hmaster0_p & v3742f25;
assign v3a559f0 = hgrant0_p & v375039e | !hgrant0_p & v37769ee;
assign v3740646 = hlock1 & v375bd8a | !hlock1 & v3a593ee;
assign v3a65e55 = hmaster0_p & v3a635ea | !hmaster0_p & v3741f67;
assign v3751b37 = hgrant4_p & v8455ab | !hgrant4_p & v3a6fadc;
assign v3a5b585 = hmastlock_p & v376bcad | !hmastlock_p & !v8455ab;
assign v372ef3e = hbusreq5_p & v3a6fd75 | !hbusreq5_p & !v3732c0d;
assign v376e1d4 = hbusreq5 & v3735b0b | !hbusreq5 & v3a6d4f3;
assign v3a69da8 = hmaster1_p & v3a6ff31 | !hmaster1_p & v3a5744d;
assign v3a6fdae = hbusreq6 & v39a5381 | !hbusreq6 & v8455ab;
assign v377c700 = hbusreq4 & v374616d | !hbusreq4 & v8455ab;
assign v3733dd8 = hbusreq6 & v3a70466 | !hbusreq6 & v3a641d5;
assign v3745f63 = hbusreq8_p & v3750797 | !hbusreq8_p & v3a6f4e0;
assign v3766126 = jx1_p & v3749f49 | !jx1_p & v376cb9d;
assign v373081f = hlock2 & v37548d8 | !hlock2 & v3a70eb6;
assign v3a60e4c = hbusreq5_p & v37745eb | !hbusreq5_p & v375e486;
assign v3a7083c = hmaster0_p & v3a70d3e | !hmaster0_p & v37660f2;
assign v3a5f20c = hbusreq0_p & v8455ab | !hbusreq0_p & v3a6d4c2;
assign v3a70f9f = hbusreq4 & v374eb71 | !hbusreq4 & !v3746303;
assign v375a56b = hbusreq8_p & v375d98c | !hbusreq8_p & v376d52a;
assign v3a70507 = hbusreq0 & v373e21a | !hbusreq0 & !v3737423;
assign v374270e = hgrant6_p & v373f8f8 | !hgrant6_p & v3a70f26;
assign v375f44a = hbusreq5 & v376ca9f | !hbusreq5 & v3a637a1;
assign v3770653 = hmaster0_p & v37666f6 | !hmaster0_p & v373f1db;
assign v3739f75 = hmaster2_p & v374f307 | !hmaster2_p & d44200;
assign v376a20e = hbusreq3 & v3a5d469 | !hbusreq3 & v3a69487;
assign v3a551e2 = hmaster1_p & fc6f92 | !hmaster1_p & v3a707a7;
assign v37294a9 = hlock5 & v3731b28 | !hlock5 & v377aed1;
assign v372b6b9 = hlock8 & v374e8f7 | !hlock8 & v376c6b3;
assign v3a70706 = hlock5_p & v3741ba8 | !hlock5_p & v3a698ed;
assign v3a705e6 = hmaster2_p & v3a62bae | !hmaster2_p & v3a701a2;
assign v3756afd = hmaster1_p & v373395b | !hmaster1_p & v3727dc9;
assign v373935b = hlock4_p & v3a700c7 | !hlock4_p & v3a702c2;
assign v37c36cb = hmaster2_p & v3768202 | !hmaster2_p & !v8455b3;
assign v3759f61 = hlock3 & v37605bb | !hlock3 & v3729d8d;
assign v375796c = hgrant4_p & v3a6ad1f | !hgrant4_p & v3a6d4b7;
assign v376fb6e = hmaster3_p & v3743fee | !hmaster3_p & v3769a63;
assign v3a61de0 = hmaster2_p & v8455ab | !hmaster2_p & v3753ee0;
assign v372de63 = hlock8 & v372b4d8 | !hlock8 & v37508df;
assign v3a71203 = hmaster0_p & v372f4ea | !hmaster0_p & v372acd0;
assign v3754b61 = hgrant2_p & v3a70a50 | !hgrant2_p & v3771e8d;
assign v373e376 = hbusreq5_p & v375238e | !hbusreq5_p & v8455b0;
assign v3a704e3 = hmaster0_p & v37368ce | !hmaster0_p & v3a59a05;
assign v3a5fc05 = hmaster0_p & v3732ecb | !hmaster0_p & !v3733767;
assign d68a4d = hbusreq4_p & v3a6143b | !hbusreq4_p & !v39a4ca8;
assign v3773ad7 = hbusreq7_p & v3751406 | !hbusreq7_p & v3a6f843;
assign v3755898 = hmaster3_p & v8455ab | !hmaster3_p & v374ae67;
assign v373698e = hgrant4_p & v376ea4a | !hgrant4_p & v3a55640;
assign v374db0f = hbusreq5_p & v37738ca | !hbusreq5_p & v375ee43;
assign v372cf51 = hgrant5_p & v3736b12 | !hgrant5_p & v3764811;
assign v376e25b = hbusreq2_p & v3a62bce | !hbusreq2_p & v8455ab;
assign v376e860 = jx1_p & v35772dd | !jx1_p & v3a6ef55;
assign v3a715a7 = hbusreq0 & v373b5b8 | !hbusreq0 & v3722f10;
assign v376cf03 = hbusreq7_p & v3a65587 | !hbusreq7_p & v377ab78;
assign v375076f = jx0_p & v3a5e660 | !jx0_p & v3a5f592;
assign v3722f65 = hbusreq4 & v3a70641 | !hbusreq4 & v8455ab;
assign v3a6fe4e = hbusreq0 & v3a6dc08 | !hbusreq0 & v8455ab;
assign v3a6665c = hgrant0_p & v3a6eeb5 | !hgrant0_p & v374c936;
assign v373ef28 = hbusreq8 & v3a6ccc6 | !hbusreq8 & v3a60276;
assign v374f645 = hlock8_p & v3768502 | !hlock8_p & v376fb92;
assign v37308fc = hmaster1_p & v373664d | !hmaster1_p & v37316f2;
assign v3774c4d = hbusreq3_p & v373dcd2 | !hbusreq3_p & v3a63621;
assign v3a703e2 = hmaster1_p & v37331a2 | !hmaster1_p & v3a7031c;
assign v372707d = hgrant4_p & v3763b9b | !hgrant4_p & v3a5b7e7;
assign v3777cae = hgrant2_p & v8455ab | !hgrant2_p & v3756559;
assign v377a5d4 = jx0_p & v8455ab | !jx0_p & v376778a;
assign v3765968 = hgrant3_p & v373e642 | !hgrant3_p & v3a6b4f6;
assign v3a7114c = hmaster2_p & v39a537f | !hmaster2_p & v3a59e87;
assign v3a6dd4d = hmaster1_p & v3756810 | !hmaster1_p & v3a62ad8;
assign v3776fae = jx2_p & v3733bed | !jx2_p & v3734c75;
assign v375822b = hmaster1_p & v375c791 | !hmaster1_p & v376f09b;
assign v374b32b = hgrant6_p & v37483dd | !hgrant6_p & v3a70d7a;
assign v3a710a2 = hlock2 & v3a7150e | !hlock2 & v374212e;
assign v373519d = hmaster0_p & v3a5e696 | !hmaster0_p & v373c1a0;
assign v3750ebc = hlock2_p & v2925c39 | !hlock2_p & !v8455ab;
assign v376b934 = hgrant8_p & v3a53e46 | !hgrant8_p & v3758cc6;
assign v3a632aa = hbusreq4_p & v3a6ff82 | !hbusreq4_p & v373b7c5;
assign v3a63203 = hbusreq6_p & v372aefc | !hbusreq6_p & v3a6ed79;
assign v3750d27 = hbusreq4_p & v3a711b5 | !hbusreq4_p & v8455ab;
assign v3a6fb86 = hbusreq0 & v3771d2d | !hbusreq0 & v372b388;
assign v3a56847 = hbusreq5_p & v3774df5 | !hbusreq5_p & !v373822e;
assign v376bc4b = hgrant0_p & v3808c39 | !hgrant0_p & v376e364;
assign v37429b9 = hgrant2_p & v8455ab | !hgrant2_p & v376dc15;
assign v37577e7 = hlock4_p & v375a116 | !hlock4_p & v373b0be;
assign v37505cd = hbusreq7_p & v3725a38 | !hbusreq7_p & v374ac6d;
assign v3773dc6 = hbusreq5_p & v373c22e | !hbusreq5_p & v3a70f4d;
assign v3a5c823 = hbusreq2_p & v3a62329 | !hbusreq2_p & v372af67;
assign v373539e = jx0_p & v3a71009 | !jx0_p & v8455ab;
assign v3a69dc1 = hbusreq4 & v3a70e5a | !hbusreq4 & v3755820;
assign v377dc72 = hmaster1_p & v3a6a758 | !hmaster1_p & v3a650a7;
assign v3a705ef = hbusreq0 & v3a70562 | !hbusreq0 & v1e37cd6;
assign v3731fd8 = hgrant4_p & v376a6f1 | !hgrant4_p & v3757b58;
assign v3722e52 = jx0_p & v3a6af23 | !jx0_p & v374c05b;
assign b09623 = stateA1_p & v3a6841c | !stateA1_p & v3777ff3;
assign v3761431 = hbusreq7_p & v37510d0 | !hbusreq7_p & v3a6fbb5;
assign v3739a53 = hbusreq6_p & v2619ae8 | !hbusreq6_p & v2acaff4;
assign v377034f = hbusreq7 & v375caa2 | !hbusreq7 & v3756200;
assign v372b034 = hmaster1_p & v3a65ee0 | !hmaster1_p & !v376a3f5;
assign v3a6f749 = hmaster0_p & v3765109 | !hmaster0_p & v3748179;
assign v374620b = hmaster1_p & v3a5b05d | !hmaster1_p & v375c003;
assign v3a29850 = hgrant4_p & v8455ab | !hgrant4_p & v37315c8;
assign v373ca17 = hbusreq7_p & v3a58c00 | !hbusreq7_p & !v8455ab;
assign v39a4e12 = hbusreq3_p & v376f73c | !hbusreq3_p & !v3732e1b;
assign v3727194 = hbusreq8_p & v374d726 | !hbusreq8_p & v3a709d5;
assign v1e3755f = hgrant3_p & v8455e7 | !hgrant3_p & v3807107;
assign v374e9c0 = hbusreq6_p & v374f35a | !hbusreq6_p & v3a68d2e;
assign v3762245 = hbusreq4_p & v373f10d | !hbusreq4_p & v3a2a14e;
assign v375bf93 = hgrant4_p & v3730e2a | !hgrant4_p & v37297e4;
assign v3a711b9 = hgrant6_p & v3744cfe | !hgrant6_p & v3752222;
assign v3753838 = hmaster1_p & v8455ab | !hmaster1_p & v3a6fc1c;
assign v3a6f2f8 = hgrant5_p & v8455ab | !hgrant5_p & !v375c099;
assign v377957e = hbusreq3_p & v2acadfb | !hbusreq3_p & !v8455ab;
assign v375818a = hbusreq5 & v8455ab | !hbusreq5 & v3a70682;
assign v3a6a73a = hbusreq5_p & v3a65d33 | !hbusreq5_p & v3a6daed;
assign v39a5382 = hgrant1_p & v3a5dbb7 | !hgrant1_p & v8455ab;
assign v375a345 = hbusreq4 & v3a6c9ab | !hbusreq4 & v2092abe;
assign v3731826 = hbusreq5_p & v3a5b45b | !hbusreq5_p & v377f734;
assign v374f21c = hbusreq5 & v37798b9 | !hbusreq5 & v3a61f85;
assign v3737a21 = hmaster1_p & v3a54b5d | !hmaster1_p & v376a3f5;
assign v377a0cb = hgrant5_p & v37621c1 | !hgrant5_p & v3746b22;
assign v3725403 = hmaster1_p & v374b564 | !hmaster1_p & v3a6574d;
assign v3a54b46 = hgrant4_p & v8455c1 | !hgrant4_p & v373446a;
assign v37384fa = hlock0_p & v3a70641 | !hlock0_p & !v8455ab;
assign v3a6a1d9 = hbusreq8 & v372bebe | !hbusreq8 & v3a635ea;
assign v37769d5 = hgrant7_p & v375f862 | !hgrant7_p & v373cedb;
assign v3a6488f = hgrant2_p & v372479c | !hgrant2_p & v3a5cc3c;
assign c0990a = hgrant4_p & v374a0c5 | !hgrant4_p & v3a61753;
assign v37377fd = hlock5 & v3741d11 | !hlock5 & v3726013;
assign v3a5c75a = hmaster2_p & v37570f8 | !hmaster2_p & v3736f61;
assign v375a4ea = hmaster2_p & v375c791 | !hmaster2_p & v3a62968;
assign v3a68116 = hmaster1_p & v374d451 | !hmaster1_p & v3a6f08c;
assign v375941a = hmaster2_p & v3a6ff25 | !hmaster2_p & v3a70da3;
assign v3748360 = hmaster2_p & v3757a88 | !hmaster2_p & v376856b;
assign v37416f0 = hbusreq0_p & a9f66a | !hbusreq0_p & v376bb26;
assign v375aae9 = hlock0_p & cf3b5d | !hlock0_p & v3a65bb5;
assign v373f836 = hbusreq6_p & v3767561 | !hbusreq6_p & v3729700;
assign v3a70cc0 = hbusreq3_p & v3749a89 | !hbusreq3_p & !v8455ab;
assign v373c1a2 = hmaster1_p & v3a661fe | !hmaster1_p & v376486a;
assign v3a5ee7a = hlock7 & a0a219 | !hlock7 & v376abcc;
assign v3763813 = hgrant5_p & v372f55a | !hgrant5_p & v3767938;
assign v23fd8b7 = hmaster1_p & v3a5af94 | !hmaster1_p & v3779288;
assign v376e794 = hbusreq2_p & v3752c04 | !hbusreq2_p & v372ea9a;
assign v3a66999 = hbusreq0 & v3a63f3d | !hbusreq0 & v39ebb74;
assign v3a6f5e1 = hlock0 & v3775999 | !hlock0 & v3737220;
assign v23fdf30 = hlock4 & v209300d | !hlock4 & v377a1d3;
assign v3a612a3 = hbusreq2_p & v3763efc | !hbusreq2_p & v8455b3;
assign v373d440 = hgrant3_p & v37655d3 | !hgrant3_p & v3a7045c;
assign v373b785 = hbusreq7 & v3773712 | !hbusreq7 & v3a5b93f;
assign v3a707cf = hmaster2_p & v3a65dcf | !hmaster2_p & v377b030;
assign v3a5e747 = hmaster2_p & v3806db0 | !hmaster2_p & v3a5c30f;
assign v3776c9c = hmaster2_p & v3a5b8b9 | !hmaster2_p & v377f526;
assign v374249a = hmaster2_p & v372455c | !hmaster2_p & !v374282f;
assign v373852b = hmaster1_p & v3a7158e | !hmaster1_p & v373d32e;
assign v3a705da = hlock7 & v373ec29 | !hlock7 & v373dc53;
assign v3a655c2 = hlock0_p & v3740171 | !hlock0_p & v39a537f;
assign v372d0db = hgrant8_p & v37544ab | !hgrant8_p & v3808904;
assign v377c671 = hbusreq6 & v3767437 | !hbusreq6 & v8455b3;
assign v3807a2e = hlock0 & v3a70a88 | !hlock0 & v375cb14;
assign v374f5a1 = hbusreq5_p & v37624a5 | !hbusreq5_p & !v3a6f6a8;
assign v374fb30 = hmaster0_p & v3a5dba4 | !hmaster0_p & v37341d3;
assign v3a6fb06 = hbusreq5 & v3a6eece | !hbusreq5 & v3a6fa7c;
assign v3a299d4 = hbusreq1_p & v37757e0 | !hbusreq1_p & v37732a0;
assign v377536e = hbusreq3_p & v3748797 | !hbusreq3_p & v3a603e0;
assign v37bfc97 = hmaster0_p & v372862a | !hmaster0_p & v8455ab;
assign v3a6e0cc = hbusreq5_p & v3769d07 | !hbusreq5_p & !v376c789;
assign v37251cc = hgrant3_p & v373197e | !hgrant3_p & v3a6f0ee;
assign v3a53e66 = hgrant4_p & v23fd83f | !hgrant4_p & v3733a5f;
assign v373a7dc = hbusreq8 & v375571e | !hbusreq8 & a0a219;
assign v375e486 = hmaster0_p & v3a6effc | !hmaster0_p & v37766fb;
assign v3727ed2 = hlock0 & v3a5f9e6 | !hlock0 & v3729030;
assign v3807723 = hmaster1_p & v3772bff | !hmaster1_p & !v377cf71;
assign v3a6f962 = hgrant6_p & v8455ca | !hgrant6_p & v3a6887f;
assign v377c842 = hbusreq4 & v37592f8 | !hbusreq4 & v8455ab;
assign cb89d9 = hbusreq3 & v375c4a1 | !hbusreq3 & v8455ab;
assign v3a5567a = hbusreq7_p & v3a6f414 | !hbusreq7_p & v3743fea;
assign v376c854 = hmaster2_p & v3a6f781 | !hmaster2_p & v3a70147;
assign v3748560 = hlock4 & v3748797 | !hlock4 & v372a04c;
assign v372a116 = hgrant6_p & v3a5bb64 | !hgrant6_p & v376dab5;
assign v375f8b1 = hbusreq7_p & v377c4bf | !hbusreq7_p & v377c9f3;
assign v374e61f = hbusreq1_p & v8455b7 | !hbusreq1_p & !v8455ab;
assign v3a70a2d = hmaster1_p & v3a573af | !hmaster1_p & v374de3d;
assign v3a6926b = hmaster1_p & v375b659 | !hmaster1_p & v375b812;
assign v3762d26 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3a6d434;
assign v376004c = hbusreq2_p & v1e37932 | !hbusreq2_p & !v8455ab;
assign v372cac5 = hbusreq4_p & v377349f | !hbusreq4_p & v3a6a1df;
assign v3770163 = hbusreq4 & v373ee80 | !hbusreq4 & v8455ab;
assign v37770c9 = hgrant6_p & v8455e7 | !hgrant6_p & v3732cb4;
assign v372e571 = hbusreq5_p & v3a5f6da | !hbusreq5_p & v3a5f4c6;
assign v3a5d217 = hmaster2_p & v372348c | !hmaster2_p & v3a6efad;
assign v39eb709 = hlock0 & v3a5741c | !hlock0 & v375d445;
assign v3a7124f = jx2_p & v3a6f04f | !jx2_p & v3a7099f;
assign v3727b4a = hbusreq6_p & v3a635ea | !hbusreq6_p & d57388;
assign v3a6cd0f = hbusreq6_p & v3a6f91a | !hbusreq6_p & v3a7057f;
assign v377fab4 = hlock7_p & v3a6fb23 | !hlock7_p & v3a6addc;
assign v37606e1 = hmaster2_p & v3a61517 | !hmaster2_p & v3722bca;
assign v3a70d6f = stateG10_1_p & v8455ab | !stateG10_1_p & !v8455e7;
assign v37792d9 = hbusreq6_p & v3750d37 | !hbusreq6_p & !v3732dc6;
assign v373e12b = hbusreq5 & v376f56d | !hbusreq5 & !v37682ce;
assign v3806b87 = hbusreq2_p & v373e369 | !hbusreq2_p & ac438c;
assign v2092bfc = hbusreq8_p & v3809b53 | !hbusreq8_p & v3778211;
assign v37732a0 = stateG10_1_p & v37757e0 | !stateG10_1_p & v3773b23;
assign v3a65b5d = hbusreq6_p & v375178f | !hbusreq6_p & v8455ab;
assign v372b57a = hgrant5_p & v3a6afcd | !hgrant5_p & v372e74c;
assign v35b71ca = hbusreq2 & v376dbdf | !hbusreq2 & v8455ab;
assign v3724b20 = hbusreq5 & v374fde8 | !hbusreq5 & !v3a6f43b;
assign v3751dd7 = hlock0 & v3748797 | !hlock0 & v9fa0b5;
assign v37501e1 = hbusreq4 & v8455c3 | !hbusreq4 & v8455b3;
assign v374e7e6 = hbusreq4_p & v37733f9 | !hbusreq4_p & v3a60258;
assign v3a6ec56 = hgrant6_p & v374bc10 | !hgrant6_p & v38095b2;
assign v3727aa3 = hlock3 & v3747c93 | !hlock3 & v3a6c0b3;
assign v3a6e82d = hmaster1_p & v374cfd8 | !hmaster1_p & v373e30f;
assign v372d593 = hgrant1_p & v3a658bf | !hgrant1_p & v35772a6;
assign v3a70a41 = hbusreq6_p & v374d674 | !hbusreq6_p & !v8455ab;
assign v99b6f5 = hmaster2_p & v3a661fe | !hmaster2_p & v8455b0;
assign v374ef3e = hbusreq7 & v377b647 | !hbusreq7 & v3749f3b;
assign v374c870 = hmaster0_p & v3773f88 | !hmaster0_p & v3a6fcab;
assign v376597e = hlock8 & v3a6fdd7 | !hlock8 & v373fe0d;
assign v37257e5 = hbusreq7 & v3a6d695 | !hbusreq7 & v8455bf;
assign v3a6fbca = hbusreq0 & v3a61895 | !hbusreq0 & v3a5e4f4;
assign v373a693 = hmaster0_p & v376c644 | !hmaster0_p & v3746a62;
assign v3731c27 = hmaster1_p & v373e5c8 | !hmaster1_p & v3a715ea;
assign a04f67 = jx3_p & v3a6df62 | !jx3_p & v372d685;
assign v39eaae4 = hbusreq7 & v3774e7b | !hbusreq7 & v3749503;
assign v3a71207 = hmaster2_p & v3a566eb | !hmaster2_p & v375bfdf;
assign v37420b6 = hmaster2_p & v376abf6 | !hmaster2_p & v3a69169;
assign v3a6bc0e = hmaster2_p & v8455ab | !hmaster2_p & v374284d;
assign v3a6570f = hbusreq5_p & v3a624d7 | !hbusreq5_p & v372316a;
assign a7f6c5 = hgrant3_p & v8455ab | !hgrant3_p & v3749408;
assign v3761bac = hbusreq5_p & v373c372 | !hbusreq5_p & v1e37b76;
assign v3a5bb49 = hmaster0_p & v374502e | !hmaster0_p & v3771b63;
assign v3a60f85 = hbusreq3 & v374e5e4 | !hbusreq3 & v3a635ea;
assign v3a582c5 = hgrant4_p & v374306c | !hgrant4_p & v375c883;
assign v3761947 = hmaster2_p & v380881d | !hmaster2_p & v8455ab;
assign v37322a9 = hmaster2_p & v8455ab | !hmaster2_p & v2acb5a2;
assign v37366da = hmaster1_p & v8455ca | !hmaster1_p & v377672d;
assign v372b48a = hbusreq5_p & v377de7f | !hbusreq5_p & v3a6107c;
assign v3a6fc7f = hgrant4_p & v377b330 | !hgrant4_p & v3a5c65e;
assign v3a6f94c = hmaster2_p & v3a6f4ba | !hmaster2_p & v1e37519;
assign v375d41f = hmaster3_p & v3a6bfb5 | !hmaster3_p & v3750e8a;
assign v375e459 = hbusreq1_p & v8455eb | !hbusreq1_p & !v8455ab;
assign v3726a7e = hmaster0_p & v374f75e | !hmaster0_p & v374ac24;
assign v375b828 = hbusreq0 & v8455b0 | !hbusreq0 & v3722e7a;
assign v372d5e5 = hmaster1_p & v3a6f417 | !hmaster1_p & v3a5f602;
assign v3770648 = jx1_p & v1e37e04 | !jx1_p & v3a6f078;
assign v3a70eba = hmaster2_p & v8455ab | !hmaster2_p & v3778a0a;
assign v3a6f86f = jx0_p & v1e37c6e | !jx0_p & v3744ad5;
assign v374ad82 = hgrant6_p & v3770559 | !hgrant6_p & v375538a;
assign v3768ac7 = hbusreq1_p & v3753f1a | !hbusreq1_p & !v8455ab;
assign v3a7117d = hlock7 & v3749ae8 | !hlock7 & v3743798;
assign v3a6fbaf = hbusreq5_p & v3a6fde5 | !hbusreq5_p & v3a6f6a8;
assign v3a5ee6b = hmaster2_p & v37430c6 | !hmaster2_p & v377de7b;
assign v3a6f42e = hbusreq0 & v37261df | !hbusreq0 & v8455ab;
assign v3776aa8 = hbusreq1_p & v95d97e | !hbusreq1_p & v3a6a9cf;
assign v37713e8 = hmaster0_p & v3a635ea | !hmaster0_p & v376456d;
assign v37332eb = hbusreq7 & v37399d4 | !hbusreq7 & v3a5666f;
assign v3742db5 = hbusreq4_p & v374da7f | !hbusreq4_p & v3753940;
assign v3a5a0d2 = hbusreq0 & v375afc7 | !hbusreq0 & v3761ba8;
assign v3755a84 = hbusreq4 & v37467da | !hbusreq4 & v3806e7b;
assign v3a703b5 = hbusreq4_p & v3753001 | !hbusreq4_p & v380919d;
assign v3739e4c = hbusreq1_p & v374f0c1 | !hbusreq1_p & v3577306;
assign v374125a = hgrant3_p & v3724f9c | !hgrant3_p & v3a5ee99;
assign v3808d48 = hmaster2_p & v3a6f43e | !hmaster2_p & v375641f;
assign v37609c3 = hbusreq8_p & v377b233 | !hbusreq8_p & !v374fcfe;
assign v372346b = hbusreq4_p & v37747a9 | !hbusreq4_p & !v8455ab;
assign v3775dfb = hmaster0_p & v375e346 | !hmaster0_p & !v3729793;
assign v3733bbe = hbusreq4 & v3a6f722 | !hbusreq4 & v374e768;
assign v3a63f3d = hgrant6_p & v3a69ae7 | !hgrant6_p & v373530a;
assign v3a6feb3 = hbusreq4_p & v3768f7f | !hbusreq4_p & v3a69430;
assign v3a6f6d3 = hbusreq0 & v3a710f6 | !hbusreq0 & v3741f5e;
assign v3a56cdc = hmaster0_p & v3a6c4e4 | !hmaster0_p & v3728fcd;
assign v376fff8 = hgrant5_p & v375b9a3 | !hgrant5_p & v37371be;
assign v3725c02 = hgrant0_p & v3a69ac0 | !hgrant0_p & v3746e79;
assign v376964a = hbusreq5_p & v3727a16 | !hbusreq5_p & v3a6efc0;
assign v3a60f71 = hbusreq6_p & v3a6f2c0 | !hbusreq6_p & v8455ab;
assign v377b4bf = hmaster0_p & v377b774 | !hmaster0_p & v3774524;
assign v375cfe0 = hbusreq5_p & v372d75d | !hbusreq5_p & v373ea8d;
assign v375f9e9 = hgrant4_p & v3a6f4c7 | !hgrant4_p & v3732bd2;
assign v3778ab3 = hmaster0_p & v37721cb | !hmaster0_p & v373cddc;
assign v3a5457f = hbusreq6 & v376a006 | !hbusreq6 & v3a5b91d;
assign v3a61e9f = hmaster0_p & v8455ab | !hmaster0_p & !v3763fec;
assign v3765442 = hbusreq7 & v3773a06 | !hbusreq7 & v3779f0a;
assign v35772c9 = hbusreq1_p & v3a70641 | !hbusreq1_p & v8455e7;
assign v372620f = hmaster0_p & v38068c8 | !hmaster0_p & v376ff64;
assign v3742140 = hbusreq6 & v3a70118 | !hbusreq6 & !v8455bd;
assign v375d059 = hgrant4_p & v374ed52 | !hgrant4_p & v372d9b0;
assign v376079d = hlock7 & v3a715b8 | !hlock7 & v377e071;
assign v37250b1 = hmaster1_p & v8455ab | !hmaster1_p & v372da0b;
assign v3a6f49e = hbusreq2_p & v3747302 | !hbusreq2_p & v373bd77;
assign v377ed18 = hmaster0_p & v3a5d2f9 | !hmaster0_p & v3a59bbd;
assign v3a6f775 = hlock0 & v3a635ea | !hlock0 & v3760088;
assign v3a6fee4 = jx0_p & v377b6ce | !jx0_p & !v8455ab;
assign v3a6767d = hbusreq6 & v373b759 | !hbusreq6 & v3767266;
assign v3768064 = hmaster0_p & v377c7c0 | !hmaster0_p & v37625f2;
assign v372424e = hgrant4_p & v3769bec | !hgrant4_p & v3748858;
assign v3734129 = hmaster1_p & v37593a4 | !hmaster1_p & v3a69a1b;
assign v37735ba = hmaster1_p & v3a640e3 | !hmaster1_p & v376314e;
assign v37251f1 = hmaster0_p & v8455bf | !hmaster0_p & v377bbf7;
assign v3755a10 = hlock0_p & v37376c8 | !hlock0_p & v3756a09;
assign v3a6be38 = hlock7 & v376374e | !hlock7 & v374067b;
assign v3806e88 = hbusreq6_p & v3a5a36d | !hbusreq6_p & v8455ab;
assign v376a297 = hmaster2_p & v3747302 | !hmaster2_p & v37697a3;
assign v377d7db = hbusreq6 & v37406d2 | !hbusreq6 & v8455ab;
assign v374a00a = hbusreq0 & v37416e1 | !hbusreq0 & v8455ab;
assign v3739a23 = hmaster0_p & v3736048 | !hmaster0_p & v3726434;
assign v3a579d1 = hmaster1_p & v8455ab | !hmaster1_p & v375485b;
assign v377f35c = hmaster1_p & v3a6fbac | !hmaster1_p & !v3a70bee;
assign v3766cfc = hlock5_p & v3a5cb4c | !hlock5_p & !v3769b75;
assign v3a68848 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3a6f94e;
assign v377d256 = hbusreq4 & v3a70209 | !hbusreq4 & !v8455ca;
assign v3a6a478 = hmaster0_p & v372baa1 | !hmaster0_p & !v3a6e8d9;
assign v3a700fe = hgrant2_p & v8455e7 | !hgrant2_p & v377d67a;
assign v3745b39 = hbusreq5_p & v3728b10 | !hbusreq5_p & v3745510;
assign v3729ed5 = hbusreq5_p & v375be54 | !hbusreq5_p & v3a652a2;
assign v373bac2 = hmaster2_p & v375649e | !hmaster2_p & v374d54c;
assign v3733727 = hlock2 & v376144f | !hlock2 & v3723c0d;
assign v377584f = hmaster1_p & v375777d | !hmaster1_p & v377055c;
assign v3a70d7e = hmaster1_p & v3a635ea | !hmaster1_p & v375e349;
assign v37564e4 = hbusreq3_p & v3a70cfb | !hbusreq3_p & v8455ab;
assign v3a7129c = hmaster0_p & v3a635ea | !hmaster0_p & v3764bf2;
assign v37564a2 = hmaster2_p & v8455b0 | !hmaster2_p & v3766202;
assign v3a6fefd = hbusreq8_p & v3751bdd | !hbusreq8_p & v3a6b937;
assign v3a608b8 = hlock5 & v3724547 | !hlock5 & v3769325;
assign v374b393 = hbusreq5 & v3a6fbee | !hbusreq5 & v8455ab;
assign v3a71353 = hbusreq6_p & v3a5b5c4 | !hbusreq6_p & v3a6da8a;
assign v3751154 = hbusreq7_p & v3737de9 | !hbusreq7_p & v3a5e998;
assign v3741cfb = hbusreq0 & v3736b57 | !hbusreq0 & v3a5e667;
assign v3764d0b = hgrant4_p & v37449b3 | !hgrant4_p & v376382c;
assign v3750254 = hgrant5_p & v39eb44e | !hgrant5_p & v3a65ae2;
assign v3a639a2 = hmaster2_p & v35b774b | !hmaster2_p & v3730e2a;
assign v325c957 = hmaster1_p & v3779fd2 | !hmaster1_p & v3a566c1;
assign v373d136 = hbusreq6_p & v3a69a04 | !hbusreq6_p & v8455b0;
assign v373d79e = hbusreq5_p & v3772183 | !hbusreq5_p & v374f4d4;
assign v3a6178c = hlock5_p & v3753418 | !hlock5_p & v374ab22;
assign v3723f1a = hbusreq2 & v3a7028d | !hbusreq2 & v8455ab;
assign v3775498 = hbusreq7_p & v3746fe7 | !hbusreq7_p & v3735b3d;
assign v3743580 = hmaster0_p & v3806c9a | !hmaster0_p & v3a5c645;
assign v377f104 = hlock0 & v3a70d64 | !hlock0 & v375c4ac;
assign v375cdf8 = hmaster2_p & v3a663c3 | !hmaster2_p & v37651b4;
assign a18d54 = hmaster1_p & v3a548a0 | !hmaster1_p & v8455ab;
assign v3a70a2a = hbusreq4 & v3a6c437 | !hbusreq4 & v8455ab;
assign v376defa = hbusreq2_p & v373de66 | !hbusreq2_p & !v3a5bf04;
assign v374fa8c = hmaster0_p & v38097ee | !hmaster0_p & v373c545;
assign v377edba = hbusreq2_p & v3a60787 | !hbusreq2_p & v3733d6e;
assign v3770cd8 = hbusreq1_p & v37234e7 | !hbusreq1_p & !v3728df3;
assign v3a68f3d = hmaster2_p & v3a614b1 | !hmaster2_p & !v8455ab;
assign v373e67e = hbusreq1_p & v8455e7 | !hbusreq1_p & !v3a70d6f;
assign v3a6aaaa = hbusreq0 & v377b0a0 | !hbusreq0 & v3750ce8;
assign v375635b = hgrant0_p & v3746404 | !hgrant0_p & v8455ab;
assign v3a708f2 = hbusreq4_p & v3a68004 | !hbusreq4_p & !v3a5ef5c;
assign v374e768 = hgrant6_p & v3a65d01 | !hgrant6_p & v3a6a116;
assign v3730a34 = hmaster0_p & v3a6ad22 | !hmaster0_p & v3a54c8b;
assign v3a6f918 = hbusreq3_p & v3776996 | !hbusreq3_p & !v8455ab;
assign v37479ee = hmaster3_p & v3722f50 | !hmaster3_p & !v376b1ee;
assign v377ba55 = hready & v3732eca | !hready & v376c211;
assign v3731977 = hmaster1_p & v3a57584 | !hmaster1_p & v3a59431;
assign v3738259 = hbusreq7 & v37475f4 | !hbusreq7 & v3768734;
assign d893c7 = hmaster2_p & c7d478 | !hmaster2_p & v8455ab;
assign v374decf = hmaster0_p & v3a66fd9 | !hmaster0_p & v3777536;
assign v3769141 = hmaster1_p & v375a397 | !hmaster1_p & v37401c2;
assign v375f2b3 = hmaster0_p & v37782c9 | !hmaster0_p & v3a70994;
assign v377618a = hbusreq6_p & v3a5c945 | !hbusreq6_p & !v3a619c0;
assign v374727f = hlock7_p & v3734579 | !hlock7_p & !v373580c;
assign v3a71368 = hmaster2_p & v3a635ea | !hmaster2_p & v23fd83f;
assign v376a47b = hmaster0_p & v3a62eee | !hmaster0_p & v3a6fb52;
assign v3a5e38d = hbusreq5 & v3a6f674 | !hbusreq5 & v8455bb;
assign v3a5a5d1 = hbusreq6_p & v376005f | !hbusreq6_p & v3762223;
assign v3a6f8b2 = hbusreq8_p & v3a64ef2 | !hbusreq8_p & v376a74a;
assign v37348e5 = jx0_p & v3767091 | !jx0_p & !v377c9b3;
assign v372f4f1 = hgrant2_p & v3a6fd27 | !hgrant2_p & v375591f;
assign v3a69796 = hbusreq0 & v373ff4a | !hbusreq0 & v3725ba8;
assign v3a70213 = hbusreq7_p & v374a89b | !hbusreq7_p & v3a58d6b;
assign v377433b = hbusreq6_p & v374b1ea | !hbusreq6_p & v3a55349;
assign v373eef7 = busreq_p & v372dd8e | !busreq_p & v8455e1;
assign v374ed51 = hbusreq3_p & v376b8e9 | !hbusreq3_p & v3a6fb84;
assign v3773137 = hbusreq2_p & v3747d3c | !hbusreq2_p & v3761efb;
assign v3a59275 = hbusreq2 & v3a70893 | !hbusreq2 & v8455ab;
assign v374287d = hmaster2_p & v374b5a8 | !hmaster2_p & v3a5f40e;
assign v3726668 = hbusreq3_p & v3a6665c | !hbusreq3_p & v39a4dd7;
assign v3a660c0 = hmaster2_p & v3806db7 | !hmaster2_p & v3a660f2;
assign v372d1bf = hgrant2_p & v3a5b12c | !hgrant2_p & v3a62986;
assign v3a5e221 = hbusreq2_p & v372f73c | !hbusreq2_p & v374a4ea;
assign v376775d = hgrant5_p & v3a64b55 | !hgrant5_p & v3733b02;
assign v37697a3 = hbusreq0 & v37729db | !hbusreq0 & v373fd50;
assign v373c219 = hlock6 & v3744adf | !hlock6 & v37662d3;
assign v3739ddd = hbusreq7_p & v374fddd | !hbusreq7_p & v374ac6d;
assign v3775526 = hbusreq5 & v3724023 | !hbusreq5 & v37bfc97;
assign v3a69e22 = hmaster2_p & v372ec6d | !hmaster2_p & v373384b;
assign v3729720 = hmaster1_p & v3a613e6 | !hmaster1_p & v3769948;
assign v37439c2 = hbusreq6 & v3751215 | !hbusreq6 & v8455ab;
assign v3764ba8 = hgrant1_p & v374a5a9 | !hgrant1_p & !v8455ab;
assign v372ed89 = hbusreq5_p & v3a6f70f | !hbusreq5_p & v8455ab;
assign v375104f = hgrant1_p & v8455b6 | !hgrant1_p & v3741e12;
assign v375e3a5 = hbusreq7_p & v3753f71 | !hbusreq7_p & v373aec3;
assign v3a5adfd = hbusreq2_p & v3745a0a | !hbusreq2_p & v372f9c3;
assign v3a64eac = hmaster0_p & v376501e | !hmaster0_p & v372b3b0;
assign v3a6a0e4 = hlock7 & v377df1a | !hlock7 & v373e062;
assign v360d109 = hbusreq2_p & v377109d | !hbusreq2_p & v3a63ff3;
assign v37739ba = hlock8_p & v3725d14 | !hlock8_p & v37622aa;
assign v3739395 = hgrant4_p & v3773e5f | !hgrant4_p & v376ddc6;
assign v373ec38 = hmaster2_p & v374e35e | !hmaster2_p & v3723b00;
assign v3733b46 = hbusreq5 & v3a70cd6 | !hbusreq5 & !v8455ca;
assign v37255d9 = hbusreq6_p & v376b4e1 | !hbusreq6_p & v374fc8e;
assign v37752af = hlock5 & v377d302 | !hlock5 & v3764306;
assign v3725b4f = hbusreq3_p & v37283a8 | !hbusreq3_p & !v3a5bf04;
assign v372410a = hbusreq4_p & v3749f51 | !hbusreq4_p & v374b07c;
assign v3a6fd17 = hgrant0_p & v3a5d822 | !hgrant0_p & v3755a10;
assign v3a714ab = hmaster0_p & v3a6a8ee | !hmaster0_p & v3a63f29;
assign v3730288 = hmaster2_p & v3806f67 | !hmaster2_p & v8455ab;
assign v3a7154e = hgrant3_p & v3739018 | !hgrant3_p & v3730452;
assign v3a6fbc7 = hlock5 & v3a5a47b | !hlock5 & v3a5b9d6;
assign v37402b8 = hmaster1_p & v3a6eb46 | !hmaster1_p & v374e21e;
assign v3a5acca = hbusreq6 & v3a55ecf | !hbusreq6 & v8455ab;
assign v375e62f = hbusreq5_p & v374fc3b | !hbusreq5_p & v8455ab;
assign v376e364 = hlock0_p & v375803a | !hlock0_p & v37461ac;
assign v374e5e4 = hlock0_p & v3a635ea | !hlock0_p & v372dfbe;
assign v3806ec2 = hlock2 & v3a5b474 | !hlock2 & v3731115;
assign v3a70cda = hbusreq4_p & v3a70b1e | !hbusreq4_p & v3a5fe39;
assign v3a6fa37 = hgrant6_p & v3a68c32 | !hgrant6_p & v3a6f744;
assign v3a71036 = hmaster0_p & v3a61397 | !hmaster0_p & v3a6416b;
assign v373413c = hbusreq2 & v3725c68 | !hbusreq2 & v3751dc9;
assign v3a5d4e9 = hbusreq8 & v376dcf6 | !hbusreq8 & v3776f7d;
assign dc5fea = hgrant4_p & v8455ab | !hgrant4_p & v3741dee;
assign v374fcfe = hmaster1_p & v3a6dfb2 | !hmaster1_p & v376980f;
assign v3258d68 = hbusreq3_p & v37757e0 | !hbusreq3_p & v3773b23;
assign v372c702 = hbusreq8_p & v3a70efb | !hbusreq8_p & v8455ab;
assign v3a61410 = hmaster2_p & v3809ebc | !hmaster2_p & v8455ab;
assign v3a65aca = hbusreq4_p & v37733f9 | !hbusreq4_p & v3a70315;
assign d320a7 = hmaster1_p & v37790c8 | !hmaster1_p & v3a683c6;
assign v374b1ea = hgrant2_p & v8455ab | !hgrant2_p & v372673b;
assign v3760eb8 = hmaster0_p & v374bc02 | !hmaster0_p & v3752281;
assign v3a6909f = hbusreq7_p & v3776445 | !hbusreq7_p & v8455ab;
assign v37297f4 = hgrant6_p & v374306c | !hgrant6_p & v374189f;
assign v3a6ff47 = hmaster2_p & v373f647 | !hmaster2_p & !v37750f7;
assign v372692d = hgrant1_p & v3a626a1 | !hgrant1_p & v3a57330;
assign v3a6c9aa = hmaster2_p & v3a6dc83 | !hmaster2_p & v375463e;
assign v3765219 = hlock4 & v3731f08 | !hlock4 & v3a6ab69;
assign v37640ff = hmaster0_p & v380974c | !hmaster0_p & v3a6eb98;
assign v3726c8c = hmaster0_p & v3728d9c | !hmaster0_p & v3a5491d;
assign v3738d51 = hgrant4_p & c51aa0 | !hgrant4_p & v3756aea;
assign v373aec4 = hmaster2_p & v373cd0c | !hmaster2_p & !v380951e;
assign v3a6ff4b = hbusreq5 & v3777647 | !hbusreq5 & !v3a715ba;
assign v37616e1 = stateG10_1_p & v8455ab | !stateG10_1_p & v3747398;
assign v377135e = hgrant6_p & v8455ab | !hgrant6_p & v37623dd;
assign v3a6fb3f = hmaster1_p & v3807aa1 | !hmaster1_p & v23fde6a;
assign v3723d31 = hbusreq8 & v37635a4 | !hbusreq8 & v8455ab;
assign v377211f = hmaster2_p & v372475d | !hmaster2_p & v3a6f4eb;
assign v3742f4c = hbusreq2 & v3771d77 | !hbusreq2 & v375d689;
assign v375c041 = hbusreq7 & v373bd8b | !hbusreq7 & v3807723;
assign v376c208 = hmaster2_p & v3a58261 | !hmaster2_p & !v8455ab;
assign v360be60 = hbusreq0 & v3764de7 | !hbusreq0 & v377bf9f;
assign v3760337 = hbusreq8_p & v3a714b7 | !hbusreq8_p & v3a63cf5;
assign v3729d8d = hbusreq3 & v3809093 | !hbusreq3 & v37438c9;
assign v3765f0a = hmaster1_p & v3a6c4e4 | !hmaster1_p & v376ff46;
assign v1e3757b = hgrant0_p & v3749c27 | !hgrant0_p & !v8455ab;
assign v3a706ef = hbusreq8_p & v3762363 | !hbusreq8_p & v3732586;
assign v3765b30 = hlock0_p & v3a653e4 | !hlock0_p & !v374c9ee;
assign v372b5c0 = hbusreq7 & v375ff99 | !hbusreq7 & v3a60276;
assign v3a6fcae = hbusreq4_p & v37558eb | !hbusreq4_p & v3a57122;
assign v3a63135 = hgrant0_p & v3726139 | !hgrant0_p & !v372a9bd;
assign v377e81a = hmaster2_p & v8455ab | !hmaster2_p & v3778528;
assign v3769302 = hbusreq0 & v373029d | !hbusreq0 & v3743f54;
assign c46b05 = hbusreq5_p & v376f4c5 | !hbusreq5_p & v3a6c31f;
assign v375b6c3 = hlock5_p & v3730a73 | !hlock5_p & !v375e93c;
assign v3a60787 = hlock0_p & v3a5891c | !hlock0_p & v3758c0d;
assign v3771160 = hmaster2_p & v2ff8c74 | !hmaster2_p & dc5fea;
assign v3a6f942 = hgrant4_p & v37609d7 | !hgrant4_p & v374c88a;
assign v3746444 = hlock8 & v92391b | !hlock8 & v3a6eee7;
assign v3768091 = hgrant4_p & v8455ab | !hgrant4_p & v375798a;
assign v3a5dc82 = hlock6 & v37761cb | !hlock6 & v37621ea;
assign v37291f8 = jx0_p & v8455ab | !jx0_p & v3a6f9be;
assign v3754f93 = hmaster2_p & v8455ab | !hmaster2_p & v8455e7;
assign v37367ba = jx1_p & v377596e | !jx1_p & v3728434;
assign v2acaff1 = hmaster1_p & v8455ab | !hmaster1_p & b1feb1;
assign v360bc74 = hmaster0_p & v3a61a7f | !hmaster0_p & v3a7012b;
assign v3747c0b = hgrant2_p & v8455ab | !hgrant2_p & v8c890d;
assign v3a713ae = hgrant6_p & v372aadd | !hgrant6_p & v375ff98;
assign v3a6a1af = hmaster2_p & v3a6dd29 | !hmaster2_p & v8455ab;
assign v3a7120c = hbusreq4 & v376e25b | !hbusreq4 & v3a70d99;
assign v3a70d38 = hlock0 & v3a635ea | !hlock0 & v3a60c49;
assign v3748d8c = stateG10_1_p & v376ba47 | !stateG10_1_p & !v38071c1;
assign v3a71660 = hgrant6_p & v3750c38 | !hgrant6_p & v377cdea;
assign v375d5f3 = hlock1_p & v377ce00 | !hlock1_p & v8455b0;
assign v373f6c9 = hbusreq3_p & v3a6b691 | !hbusreq3_p & v3a640c5;
assign v37724ca = hbusreq1 & d44200 | !hbusreq1 & v8455ab;
assign v3724efc = hmaster1_p & v373e0d0 | !hmaster1_p & v3752b5c;
assign v372874c = hgrant6_p & v8455ab | !hgrant6_p & !v3a6f804;
assign v3a58e15 = hmaster1_p & v3756cf2 | !hmaster1_p & v3752913;
assign v3752e1b = hbusreq4_p & v37539fc | !hbusreq4_p & v3a60d86;
assign v3779f1c = hgrant6_p & v8455ab | !hgrant6_p & v3a6fd50;
assign v3736dc2 = hmaster2_p & v374a6a5 | !hmaster2_p & v375d5ac;
assign v3806f1f = hgrant5_p & v3a6cf91 | !hgrant5_p & v3a69036;
assign v37592f8 = hgrant6_p & v91cdff | !hgrant6_p & v3a5da57;
assign v3a62ce4 = hbusreq5_p & v3a6c6ac | !hbusreq5_p & v8455ab;
assign v37444ae = jx0_p & v376d81a | !jx0_p & v1e37ae9;
assign v3a70b17 = hbusreq3_p & v3a710b5 | !hbusreq3_p & v8455ab;
assign v8e4471 = hgrant5_p & v3723f0c | !hgrant5_p & v3a708b6;
assign b66167 = hgrant4_p & v3723b00 | !hgrant4_p & v374616d;
assign v3755806 = hlock3_p & v3a60711 | !hlock3_p & v8455ab;
assign v373744b = hbusreq2_p & v3809ebc | !hbusreq2_p & !v3727976;
assign v9243ac = hlock5 & v373a4cd | !hlock5 & v37373bb;
assign v372c903 = hbusreq2_p & v3753b5e | !hbusreq2_p & v38072fd;
assign v3764834 = hgrant1_p & v8455b6 | !hgrant1_p & v3723430;
assign v3a6f02e = hgrant3_p & v37522bc | !hgrant3_p & v3a6f1c5;
assign v3a611bd = hmaster2_p & v375dcac | !hmaster2_p & v37551b9;
assign v3769404 = hbusreq3 & v3738397 | !hbusreq3 & bdda12;
assign v3a56aeb = hbusreq3_p & v373cdb7 | !hbusreq3_p & v3732302;
assign v3726023 = hmaster2_p & v373a7a5 | !hmaster2_p & v3a71134;
assign v377b838 = hlock5 & v377de7f | !hlock5 & v372a309;
assign v3747804 = hbusreq7 & v3772098 | !hbusreq7 & v37297ac;
assign v3733542 = hgrant6_p & v37414b0 | !hgrant6_p & v3a70a95;
assign v377faae = hlock5_p & v3734419 | !hlock5_p & v373c04a;
assign v37582c2 = hmaster2_p & v377437d | !hmaster2_p & v37430e7;
assign v3a5fb90 = hmaster1_p & v23fdac1 | !hmaster1_p & v8455b9;
assign v3a6cd89 = hmaster3_p & v372facf | !hmaster3_p & v372cf2e;
assign v3734dd6 = hmaster2_p & v375d800 | !hmaster2_p & v376358f;
assign v3a584be = hbusreq5_p & v3724394 | !hbusreq5_p & v372b902;
assign v3a6f80b = hmaster1_p & v3772904 | !hmaster1_p & v3a68289;
assign v375e75d = hbusreq4_p & v3758636 | !hbusreq4_p & v3809240;
assign v373b4ce = hbusreq3_p & v2aca977 | !hbusreq3_p & v3a6fd79;
assign v376935b = hbusreq4_p & v3a704c7 | !hbusreq4_p & !v3a6f2e1;
assign v8455b1 = hbusreq0_p & v8455ab | !hbusreq0_p & !v8455ab;
assign v3a6ffeb = hbusreq8_p & v3731202 | !hbusreq8_p & v376fbe5;
assign v3a64a09 = hbusreq4_p & v3747302 | !hbusreq4_p & v3a6c5ee;
assign v374071d = hbusreq7_p & v894fb9 | !hbusreq7_p & v3a6fcd8;
assign v373f5fc = jx0_p & v3740d9e | !jx0_p & v374f243;
assign v372e169 = hlock1 & v3727507 | !hlock1 & v374e2a1;
assign v325b5e0 = hgrant2_p & v3a71460 | !hgrant2_p & v37671ad;
assign v3a712d6 = hgrant2_p & v377182c | !hgrant2_p & v37538e4;
assign v3807413 = hbusreq7 & v3a6f474 | !hbusreq7 & v3a55491;
assign v3a6c4a4 = hmaster0_p & v3a6f7dd | !hmaster0_p & v377c065;
assign v3a6f506 = hmaster0_p & v3746cbf | !hmaster0_p & v3769f01;
assign v3a694b9 = hmaster0_p & v3a5711b | !hmaster0_p & !v37654c4;
assign v3a6fe75 = hbusreq5 & v37655c5 | !hbusreq5 & v373755a;
assign v3768383 = hlock6 & v374af2f | !hlock6 & v3a70b56;
assign v377a855 = hgrant5_p & v3a6fc07 | !hgrant5_p & v3a7079d;
assign v372d035 = hmaster0_p & v372de68 | !hmaster0_p & v376aaef;
assign v376093b = hmaster2_p & v37583be | !hmaster2_p & !v37388ce;
assign v375afbf = hmaster1_p & v3744280 | !hmaster1_p & v372ef3e;
assign v3a6cfa1 = hgrant5_p & b58331 | !hgrant5_p & v374ac57;
assign v3a6f457 = hgrant2_p & v8455ab | !hgrant2_p & v8455ef;
assign v380761c = hgrant3_p & v377abd1 | !hgrant3_p & v37402f0;
assign v3a68bb1 = hbusreq6 & v3a5d3af | !hbusreq6 & v3a69c05;
assign v374ac8a = hmaster3_p & v8455ab | !hmaster3_p & v377cc72;
assign v377119f = hgrant5_p & v8455ab | !hgrant5_p & v377894f;
assign v3a7052e = hmaster2_p & v3747302 | !hmaster2_p & v3779cf9;
assign v3a70425 = hbusreq6 & v3724aaf | !hbusreq6 & v8455ab;
assign v3754871 = hbusreq2 & v3751734 | !hbusreq2 & !v8455ab;
assign v374d99a = hgrant6_p & v3725fe1 | !hgrant6_p & v9644fd;
assign v3772e0a = hbusreq2_p & v380761c | !hbusreq2_p & v3a71547;
assign v3a702ec = hgrant2_p & v8455ba | !hgrant2_p & v3737a30;
assign v375ecff = hbusreq4_p & v372a3af | !hbusreq4_p & v3a7029f;
assign v3a2a2fa = hlock0_p & v37682a8 | !hlock0_p & v3764f8a;
assign v3a61b45 = hbusreq5 & v374e1fd | !hbusreq5 & v8455ab;
assign v372988e = hgrant4_p & v372dffe | !hgrant4_p & v3767a93;
assign v3747243 = hmaster2_p & v3a6a939 | !hmaster2_p & v3765e46;
assign v3751ab7 = hbusreq0 & v377d86e | !hbusreq0 & v1e37cd6;
assign v3773daf = hbusreq7_p & v3a7137d | !hbusreq7_p & !v37797f4;
assign v372d6e5 = hbusreq3_p & v3a6fcf9 | !hbusreq3_p & v3a71644;
assign v37302c7 = hmaster2_p & v3747302 | !hmaster2_p & v3a6f71a;
assign v374a556 = hbusreq5_p & v374f0c1 | !hbusreq5_p & v23fe061;
assign v377b612 = hbusreq2_p & v3a713e3 | !hbusreq2_p & v3a701b3;
assign v3a6fe0a = hgrant3_p & v8455ab | !hgrant3_p & v3a71378;
assign v3a5b4bd = hmaster0_p & v373f911 | !hmaster0_p & v3746a62;
assign v3755136 = hmaster2_p & v8455ab | !hmaster2_p & v3772715;
assign v37764b1 = hbusreq1 & v37386a9 | !hbusreq1 & v3a635ea;
assign v37671ad = hbusreq2_p & v3a56f66 | !hbusreq2_p & v3a6a1f4;
assign v3a58836 = stateG10_1_p & v3a700a5 | !stateG10_1_p & !bda6d5;
assign v3a5e363 = hgrant2_p & v373681a | !hgrant2_p & v35b70e6;
assign v3756d56 = hmaster3_p & v3a70fde | !hmaster3_p & v8455ab;
assign v3734827 = hgrant4_p & v1e37b99 | !hgrant4_p & v3749686;
assign v3775688 = hgrant4_p & v8455ab | !hgrant4_p & v377e698;
assign v37529d6 = hlock7 & v9fecca | !hlock7 & v372d2cd;
assign v3759f09 = hbusreq0 & v375c0c4 | !hbusreq0 & v3760b79;
assign v3a710bf = hmaster1_p & v3a679e2 | !hmaster1_p & v376a411;
assign v3a6f235 = hmaster0_p & v3a6f475 | !hmaster0_p & v3732938;
assign v3a62d59 = hbusreq6 & v372310a | !hbusreq6 & v3755a0f;
assign v3a70b26 = hmaster1_p & v8455ab | !hmaster1_p & !v3768a11;
assign v3a703d3 = hgrant2_p & v8455ab | !hgrant2_p & v3761efb;
assign v373fb32 = hmaster3_p & v8455ab | !hmaster3_p & v376fe7d;
assign v3749b37 = hbusreq2 & v3731ffc | !hbusreq2 & v3a70a88;
assign v3a58307 = hlock7_p & v8ac439 | !hlock7_p & v375c648;
assign v376223b = hbusreq2 & v3a5600a | !hbusreq2 & v3766ea9;
assign v373bd5e = hgrant5_p & v3809e97 | !hgrant5_p & v3a5d97a;
assign v375a8d5 = hmaster1_p & v377d077 | !hmaster1_p & v37650d7;
assign v3a6b23f = hgrant2_p & v375c7b9 | !hgrant2_p & v3a65f4c;
assign v3a59e1c = hbusreq0 & v8455b0 | !hbusreq0 & v3a54c2e;
assign v3a70d77 = hlock6_p & v374b3bf | !hlock6_p & v37406d2;
assign v3759fe0 = hbusreq2_p & v3725a06 | !hbusreq2_p & v3a5cc4c;
assign v37745e0 = hbusreq2_p & v37432c6 | !hbusreq2_p & !v37521ed;
assign v3a66c5c = hbusreq2_p & v3a6eb6b | !hbusreq2_p & v3742d37;
assign v3a57f64 = hbusreq8 & v37255a2 | !hbusreq8 & !v3772cc3;
assign v375e5bb = hmaster2_p & v3775303 | !hmaster2_p & v8455ab;
assign v3a62e42 = hmaster2_p & v3a70cec | !hmaster2_p & v376112d;
assign v3a70568 = hgrant3_p & v3744dd2 | !hgrant3_p & v3756943;
assign v373f94e = hbusreq4_p & v8455ab | !hbusreq4_p & v3a5e239;
assign v374638c = hgrant6_p & v37711cc | !hgrant6_p & v3a58b28;
assign v3a5d2f9 = hmaster2_p & v377b330 | !hmaster2_p & v37786a6;
assign v3761031 = hgrant4_p & v8455ab | !hgrant4_p & v3a6fe8a;
assign v372a414 = hbusreq3 & v3a6e438 | !hbusreq3 & v8455ab;
assign v3a70371 = hgrant4_p & v8455c1 | !hgrant4_p & v3a67257;
assign v377e867 = hbusreq2_p & v376c569 | !hbusreq2_p & v3a6f4c5;
assign v376e90a = hbusreq3_p & v3a635ea | !hbusreq3_p & v377c6b3;
assign v3a6f133 = stateG10_1_p & v8455ab | !stateG10_1_p & v3763788;
assign v3729b33 = hbusreq2 & v8455ab | !hbusreq2 & v95d97e;
assign v377e071 = hgrant5_p & v3760989 | !hgrant5_p & v3768e14;
assign v1e374cc = hbusreq6 & v3740171 | !hbusreq6 & v8455e7;
assign v376508b = hmaster0_p & v3a6facd | !hmaster0_p & v3a708e0;
assign v3a5b826 = hbusreq0 & v3a6f102 | !hbusreq0 & v3a6f0d3;
assign v3a5b90b = hbusreq2_p & v3776b18 | !hbusreq2_p & !v8455ab;
assign v3a6f04c = hgrant6_p & v8455ab | !hgrant6_p & v3775a4f;
assign v3a58964 = hlock0_p & v3a5891c | !hlock0_p & !v37528b0;
assign v377180a = jx0_p & v3770c98 | !jx0_p & v8455ab;
assign v376c6ed = hbusreq6 & v3726c5b | !hbusreq6 & v373c965;
assign v37431ec = hgrant4_p & v3771d4f | !hgrant4_p & v3768e7e;
assign v377c29f = hgrant3_p & v360d1cb | !hgrant3_p & v3a711a9;
assign v37331af = hbusreq6_p & v3731fc6 | !hbusreq6_p & v3a57ed1;
assign v3a56fcd = hbusreq3_p & v376a20e | !hbusreq3_p & v3757e0b;
assign v3a5c7ca = hmaster1_p & v3745b71 | !hmaster1_p & !v3a2abf4;
assign v3755ec0 = hbusreq0 & v373ffa9 | !hbusreq0 & v8455ab;
assign v3733083 = hmaster2_p & v372ab21 | !hmaster2_p & v8455ab;
assign v3a57d2f = hgrant6_p & v8455ab | !hgrant6_p & v377c258;
assign v3a6bb4b = hmaster3_p & v376fe00 | !hmaster3_p & v3a62e20;
assign v375c31a = hlock2 & v374d8cb | !hlock2 & v3a5923c;
assign v377f5ca = hmaster1_p & v3a635ea | !hmaster1_p & v3806599;
assign v375076a = hbusreq5 & v3808e6b | !hbusreq5 & v3a6fe91;
assign v372f05b = hbusreq8 & v372f23a | !hbusreq8 & v376d85d;
assign v3a6a22c = hbusreq4_p & v3a7012f | !hbusreq4_p & v35772a6;
assign v372e374 = hgrant5_p & v3a70578 | !hgrant5_p & v3762ca6;
assign v37519a8 = hmaster0_p & v3747892 | !hmaster0_p & v3a6e93d;
assign v375bc6f = hgrant5_p & v8455ab | !hgrant5_p & v3726448;
assign v3769c7f = hbusreq0 & v3a70322 | !hbusreq0 & v372b8d7;
assign v3a71677 = hmaster0_p & v3a6ef5a | !hmaster0_p & v374d8ea;
assign v37578f3 = hbusreq4 & v3a66aa4 | !hbusreq4 & v35b774b;
assign v3a6a910 = hbusreq6 & v8455b0 | !hbusreq6 & adf78a;
assign v373fecb = hlock8_p & v3378f5b | !hlock8_p & v3a70e5c;
assign v3808d68 = hgrant5_p & v8455ab | !hgrant5_p & v3378b6c;
assign v3a714b1 = hbusreq6_p & v35772a2 | !hbusreq6_p & v3a70cc3;
assign v3742f25 = hmaster2_p & v3757765 | !hmaster2_p & v8455ab;
assign v373e5c8 = hbusreq5_p & v3730389 | !hbusreq5_p & v3761f78;
assign v377b074 = hgrant7_p & v8455ab | !hgrant7_p & v3a5a260;
assign v3776125 = hbusreq6 & v3755a0f | !hbusreq6 & v37496fa;
assign v376d57d = hmaster1_p & v3745939 | !hmaster1_p & v374bf0f;
assign v3765758 = hbusreq0 & v3773fbb | !hbusreq0 & v375dd2b;
assign v374a25d = hmaster1_p & v8455ab | !hmaster1_p & v374dcfb;
assign v3a71617 = hbusreq0 & v375bdd4 | !hbusreq0 & !v3a6ebf1;
assign v3762de5 = hmaster1_p & v373013d | !hmaster1_p & v3a5f0d0;
assign v3755738 = hmaster2_p & v3a635ea | !hmaster2_p & v3a6fa4c;
assign v375f78f = hmaster2_p & v37556fd | !hmaster2_p & v373e209;
assign v3778754 = hbusreq4_p & v374998d | !hbusreq4_p & v37285eb;
assign v3a6fe07 = hbusreq8 & v3741418 | !hbusreq8 & v375b801;
assign v3752b8f = hmaster2_p & v3a59217 | !hmaster2_p & !v3a7141c;
assign v3a5ab6e = hgrant3_p & v3a635ea | !hgrant3_p & v3a57b0d;
assign v377abd1 = hbusreq3_p & v3a5c945 | !hbusreq3_p & !v3a66110;
assign v373c26c = hmaster1_p & v8455ab | !hmaster1_p & v374e78a;
assign v373c2a2 = hgrant4_p & v372b77b | !hgrant4_p & v2aca264;
assign v37432c6 = hbusreq3_p & v3759032 | !hbusreq3_p & v3733e9e;
assign v373e16b = hmaster2_p & v3a5fc82 | !hmaster2_p & v372348c;
assign v3a5cb45 = hbusreq6_p & v374113d | !hbusreq6_p & v3725dc4;
assign v3a70f8d = hlock6 & v3a70b76 | !hlock6 & v37554c0;
assign v373f537 = hgrant5_p & v3761ca6 | !hgrant5_p & v397fb7c;
assign v8455b7 = hlock1_p & v8455ab | !hlock1_p & !v8455ab;
assign v37796ee = hbusreq6_p & v3735fc0 | !hbusreq6_p & v3748d67;
assign v3a6efb7 = hbusreq8 & v3a69d78 | !hbusreq8 & !v8455ab;
assign v3a5a37a = hmaster0_p & v3a65e17 | !hmaster0_p & v3a68b7d;
assign v3a7144a = hbusreq6 & v3770e35 | !hbusreq6 & v375f9df;
assign v372fbeb = hlock4_p & v39a535f | !hlock4_p & v8455ab;
assign v3a7068f = hmaster1_p & v3751e0a | !hmaster1_p & v3735859;
assign v3a708f0 = hgrant2_p & v3a62a6d | !hgrant2_p & v37c0077;
assign v380733a = hbusreq3 & v3768062 | !hbusreq3 & v3a6c5ee;
assign v3a6fa86 = hbusreq4 & v3a70468 | !hbusreq4 & v374af92;
assign v3a6f5d2 = hbusreq6_p & v375306b | !hbusreq6_p & v3a6dcdc;
assign v374e033 = hbusreq5_p & v3745abb | !hbusreq5_p & v8455ab;
assign v3739791 = hbusreq4_p & v376107b | !hbusreq4_p & v8455e7;
assign v37c028b = hmaster1_p & v3a5e24e | !hmaster1_p & v3a70a31;
assign v372dcff = hmaster2_p & v373e6d2 | !hmaster2_p & v372424e;
assign v3729fa0 = hlock4 & v37411bc | !hlock4 & v3762385;
assign v3752e24 = hgrant6_p & v372493b | !hgrant6_p & v3744d18;
assign v37737b9 = hbusreq5_p & v3727f68 | !hbusreq5_p & !v3a69dbd;
assign v373c5ea = hmaster1_p & v3809af2 | !hmaster1_p & v3a6f974;
assign v37618dc = hburst0 & v3a6f776 | !hburst0 & v3763eaa;
assign v377a92d = hmaster0_p & v3a58cfc | !hmaster0_p & !v3a6f443;
assign v3a709ba = hbusreq4 & v374291b | !hbusreq4 & v37519ea;
assign v3752f2e = hgrant6_p & v3a605b5 | !hgrant6_p & v3a65605;
assign v3764203 = hmaster2_p & v3765e79 | !hmaster2_p & v3a6f71a;
assign v3a70c13 = hgrant4_p & v375380a | !hgrant4_p & v3749686;
assign v37766b2 = hmaster3_p & v3a622a9 | !hmaster3_p & v3a70122;
assign v3a6f0e3 = hbusreq2_p & v3758dfe | !hbusreq2_p & v3a6eee6;
assign v376662b = jx3_p & v3751fde | !jx3_p & v38096d8;
assign v3729d06 = hmaster1_p & v8455ab | !hmaster1_p & v373c8ac;
assign v3a573ec = hbusreq7_p & v37249fe | !hbusreq7_p & v3764383;
assign v3a54466 = hmaster0_p & v3726023 | !hmaster0_p & v3764ed7;
assign v373144a = hmaster0_p & v3a6a54d | !hmaster0_p & v3759584;
assign v3a664ed = hbusreq7 & v3a6fb6f | !hbusreq7 & v8455ab;
assign v374943a = hlock5_p & v373ad86 | !hlock5_p & !v38098bf;
assign v377ea64 = hmaster0_p & v37640e9 | !hmaster0_p & v3a6f495;
assign v376dba6 = hgrant6_p & v3739d45 | !hgrant6_p & v375ecf5;
assign v3a5952d = hbusreq1_p & v3763793 | !hbusreq1_p & !v8455ab;
assign v37381c2 = hmaster0_p & v8455ab | !hmaster0_p & v374a46d;
assign v3a5db06 = hmaster0_p & v377a865 | !hmaster0_p & v3a7017e;
assign v37753f2 = hgrant3_p & v3747c3e | !hgrant3_p & v8455ab;
assign v373869b = hbusreq4_p & v3777ce4 | !hbusreq4_p & v372c84a;
assign v373447d = hbusreq3_p & v3728c46 | !hbusreq3_p & !v8455ab;
assign v3a532f2 = hmaster3_p & v8455ab | !hmaster3_p & v372700e;
assign v3a5cb4c = hmaster0_p & v3779060 | !hmaster0_p & v37500e0;
assign v373a27c = locked_p & v8455ab | !locked_p & v37566b2;
assign v972988 = hmaster0_p & v3a6f1b7 | !hmaster0_p & v3a5f992;
assign v37565af = hmaster2_p & v3a6e31f | !hmaster2_p & !v3735e39;
assign v372b7cc = hgrant6_p & v3a71389 | !hgrant6_p & v3a6b2e5;
assign v3a6a557 = hmaster0_p & v37356f0 | !hmaster0_p & v3746c51;
assign v375931f = hbusreq5 & v3a70936 | !hbusreq5 & v3730d6b;
assign v2092f59 = hbusreq2_p & v373ff4a | !hbusreq2_p & bdc54c;
assign v3a69de7 = locked_p & v3750fc8 | !locked_p & v3a635ea;
assign v3727f9c = hbusreq5_p & v3773340 | !hbusreq5_p & v88e7d1;
assign v3a70f6a = hburst1 & v3a6f8df | !hburst1 & v3a6f02c;
assign v372dd0c = hbusreq0 & v375e91f | !hbusreq0 & v8455ab;
assign v37735ec = hgrant0_p & v3a66492 | !hgrant0_p & v8455ab;
assign v3771d0f = hbusreq2_p & v3a5ab6e | !hbusreq2_p & v377002f;
assign v3764132 = hbusreq4_p & v375c4e6 | !hbusreq4_p & v8455ab;
assign v373ec1f = hlock5_p & v3a70d5f | !hlock5_p & v8455ab;
assign v1e37e66 = hready & v37779ea | !hready & v8455ab;
assign v37520ee = hmaster2_p & v37297d0 | !hmaster2_p & v374fe54;
assign v375cfd7 = hbusreq6 & v377e60e | !hbusreq6 & v373c965;
assign v376abd3 = hbusreq5_p & v374bd38 | !hbusreq5_p & !v8455ab;
assign v375084d = hlock6 & v3729e5f | !hlock6 & v3a6b37c;
assign v3758f2e = hmaster2_p & v3a70326 | !hmaster2_p & v3748609;
assign v3a620f2 = hmaster1_p & v3774db3 | !hmaster1_p & v3761e97;
assign v3764c4a = hbusreq7_p & v3a6aa15 | !hbusreq7_p & v3807029;
assign v37286e7 = hgrant5_p & v376ee65 | !hgrant5_p & v3a5dd70;
assign v376ac08 = hbusreq6_p & v374b21a | !hbusreq6_p & v8455ab;
assign v37783ba = hmaster0_p & v8455ab | !hmaster0_p & v37434e1;
assign v37504b9 = hgrant0_p & v3735f56 | !hgrant0_p & v3a7094a;
assign v3a5dd62 = hbusreq4 & v3a59264 | !hbusreq4 & v3752767;
assign v3a709f8 = hbusreq0 & v3765ef0 | !hbusreq0 & v8455ab;
assign v3745452 = hbusreq6 & v2acaf41 | !hbusreq6 & v3746efb;
assign v1e37b99 = hbusreq4_p & v8455e7 | !hbusreq4_p & !v8455ab;
assign v3758c07 = hmaster0_p & v8455b0 | !hmaster0_p & v376b86f;
assign v376da8d = jx0_p & v9c9e05 | !jx0_p & v3a70ed8;
assign v3768180 = hmastlock_p & v3a5a496 | !hmastlock_p & !v8455ab;
assign v3a583b0 = hmaster2_p & v8455ab | !hmaster2_p & v376c1de;
assign v37463e5 = hgrant6_p & v3a5e7c0 | !hgrant6_p & v3a5757f;
assign v3a70347 = hmaster0_p & v373dd7f | !hmaster0_p & v3779988;
assign v3a56cca = hlock4 & v376b2a2 | !hlock4 & v373abae;
assign v3a6f2af = hgrant4_p & v8455ab | !hgrant4_p & v3a6f3af;
assign v3a670a1 = hbusreq1_p & v3a64566 | !hbusreq1_p & !v373e16a;
assign v3a6f22c = hbusreq2_p & v3754202 | !hbusreq2_p & v8455ab;
assign v376f24b = hbusreq7_p & v39a4eaa | !hbusreq7_p & v3a537c5;
assign v3a703ad = hgrant3_p & v376495e | !hgrant3_p & v375c4a1;
assign v37667eb = hbusreq8 & v3760e1b | !hbusreq8 & v3a6ec0f;
assign v3a7078d = hbusreq7 & v376924d | !hbusreq7 & v3808914;
assign v377c15d = hbusreq5_p & v3a5c3a0 | !hbusreq5_p & v373e474;
assign v3a60976 = hmaster2_p & v3a635ea | !hmaster2_p & v3764418;
assign v3745aff = hbusreq3 & v1e37e76 | !hbusreq3 & v8455ab;
assign v3755774 = hmaster2_p & v37325a2 | !hmaster2_p & d5f283;
assign v3a712dd = hgrant4_p & v372d1d7 | !hgrant4_p & !v8455ab;
assign v372d816 = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a6ff58;
assign v372ba4d = hbusreq3 & v3749435 | !hbusreq3 & v8455ab;
assign v3755199 = hgrant6_p & v8455ca | !hgrant6_p & v3774908;
assign v377f6c3 = hmaster0_p & v3726c61 | !hmaster0_p & v3a6f49f;
assign v373b759 = hgrant2_p & v377cd0d | !hgrant2_p & v3a658b0;
assign v3779860 = hlock4_p & v37718fb | !hlock4_p & v3a57309;
assign v3a56608 = hlock2 & v2092f5e | !hlock2 & v3a6b560;
assign v3a6f579 = hgrant6_p & v8455c9 | !hgrant6_p & v376ed30;
assign v3a63df4 = hgrant4_p & v37716ca | !hgrant4_p & v373dfb5;
assign v37371df = hlock5_p & a94d63 | !hlock5_p & v373a327;
assign v3a6f4e3 = hmaster0_p & v3a5fabd | !hmaster0_p & v3766df8;
assign v3a65088 = hlock5_p & v3775651 | !hlock5_p & v35772a6;
assign v3735675 = hmaster0_p & v3771ce2 | !hmaster0_p & v3760c1b;
assign v3734583 = hlock5 & v37711ec | !hlock5 & v3a69758;
assign v377de92 = hgrant2_p & v375ca6c | !hgrant2_p & v375e551;
assign v917443 = hmaster1_p & v374ab4b | !hmaster1_p & v373c437;
assign v3727cec = hlock7_p & v3a6681e | !hlock7_p & v3769310;
assign v380951e = hgrant4_p & v3a70272 | !hgrant4_p & v3776ea4;
assign v3773390 = hbusreq6_p & v3a5457f | !hbusreq6_p & v3a5b91d;
assign v3a67c36 = hbusreq4_p & v377789d | !hbusreq4_p & !v8455ab;
assign v377f3af = hburst1_p & v8455ab | !hburst1_p & !v3730383;
assign v3a6fd6f = hgrant1_p & v3a71571 | !hgrant1_p & v35772a6;
assign v3a7130e = hlock5_p & v377115d | !hlock5_p & v8455cb;
assign v3a2aed2 = hbusreq5_p & v3a71132 | !hbusreq5_p & v3a659f5;
assign v375ca08 = hbusreq3 & v2acaff4 | !hbusreq3 & v8455ab;
assign v376e17a = hbusreq4_p & v374d970 | !hbusreq4_p & v3744792;
assign v374990a = hbusreq8 & v3a710f8 | !hbusreq8 & v3a6fe04;
assign v3763d20 = hgrant4_p & v3751e76 | !hgrant4_p & v3778281;
assign v3750b04 = hlock2_p & v3722e5c | !hlock2_p & v35772a6;
assign v376fc23 = hbusreq7_p & v3a6eefa | !hbusreq7_p & v37658de;
assign v2ff87d2 = hmaster0_p & v8455ab | !hmaster0_p & !v377f424;
assign v37444e7 = hmaster1_p & v3a7067e | !hmaster1_p & v8455ab;
assign v3a6fa93 = hgrant4_p & v3759032 | !hgrant4_p & v372f37d;
assign v3755b5c = hmaster0_p & v3730bd8 | !hmaster0_p & v375820e;
assign v3a5baf5 = hmaster1_p & v374e99f | !hmaster1_p & v3774399;
assign v372d4eb = hlock5 & v372354b | !hlock5 & v374d255;
assign v37662e7 = hmaster2_p & v3a5f1d4 | !hmaster2_p & v3a6f138;
assign v3a69036 = hmaster1_p & v3a6fce0 | !hmaster1_p & v372c8d0;
assign v377b058 = hmaster2_p & v3a6fa4c | !hmaster2_p & v3a6eb7b;
assign v37736c4 = hbusreq7 & v377e071 | !hbusreq7 & v372f1a8;
assign v1e37acb = hmaster1_p & v3753418 | !hmaster1_p & v376c014;
assign v3a5f358 = hbusreq8 & v37529d6 | !hbusreq8 & v3a6cf88;
assign v3727540 = hmaster0_p & v37430c6 | !hmaster0_p & v3a5ee6b;
assign v373cc68 = hlock1_p & v3755791 | !hlock1_p & !v8455ab;
assign v372e1b6 = hbusreq5_p & v376bfa7 | !hbusreq5_p & !v37627f6;
assign v3a64703 = hgrant3_p & v3a7106f | !hgrant3_p & v372b9c6;
assign v375e50f = hmaster1_p & v377b3bd | !hmaster1_p & v373ed57;
assign v377a018 = stateG10_1_p & v3a637dd | !stateG10_1_p & !v3a690ff;
assign v3a5b541 = hbusreq4_p & v3728127 | !hbusreq4_p & v3724368;
assign v3746be0 = hgrant4_p & v8455ab | !hgrant4_p & v922f0a;
assign v372c433 = hlock5_p & v377086c | !hlock5_p & v3738f35;
assign v3758df6 = hgrant4_p & v3a5bb64 | !hgrant4_p & v372a116;
assign v373ff4a = hlock0_p & v3730627 | !hlock0_p & v8455b7;
assign v377e39f = hbusreq2 & v3a59409 | !hbusreq2 & !v8455ab;
assign v3808f2f = hbusreq7 & v360d0fb | !hbusreq7 & v37582e7;
assign v374d402 = hgrant6_p & v375f3e2 | !hgrant6_p & v3779081;
assign v3774391 = hmaster0_p & v3775dbc | !hmaster0_p & v3742f52;
assign v3a7156a = hlock0 & v374a637 | !hlock0 & v37232a6;
assign v3a63ece = hmaster0_p & v37793e4 | !hmaster0_p & v37293e0;
assign v372b870 = hgrant5_p & v3762de5 | !hgrant5_p & v37289bc;
assign v3723404 = hlock6 & v3a6ec52 | !hlock6 & v373cb58;
assign v3730712 = hgrant5_p & v8455c1 | !hgrant5_p & v3793188;
assign v3a582d8 = hbusreq0 & v1e38288 | !hbusreq0 & v3a6180b;
assign v37256c0 = jx0_p & v3a648f6 | !jx0_p & v3807174;
assign v373d964 = hmaster0_p & v3a6bce0 | !hmaster0_p & v3736d58;
assign v3a71138 = hgrant6_p & v3759b6f | !hgrant6_p & v37576d1;
assign v1e37c38 = hmaster2_p & v3732f8d | !hmaster2_p & v3738c0a;
assign v3a71541 = hmaster0_p & v3a712c8 | !hmaster0_p & !v3a6cf7f;
assign v3777ff7 = stateA1_p & v8455ab | !stateA1_p & !aa6771;
assign v37548d8 = hbusreq2 & v3a70eb6 | !hbusreq2 & v3a635ea;
assign v3761cd5 = hbusreq4_p & v3722f65 | !hbusreq4_p & !v8455c2;
assign v3a6eb3c = hgrant3_p & v374d42c | !hgrant3_p & !v8455ab;
assign v3745020 = hbusreq0_p & v3a5d673 | !hbusreq0_p & v8455b5;
assign v3a5ff4b = hmaster2_p & b68bf2 | !hmaster2_p & v3a711ed;
assign v3a6aea2 = hmaster3_p & v375c32d | !hmaster3_p & v8455ab;
assign v377845d = hbusreq5_p & v3745e51 | !hbusreq5_p & v37c014f;
assign v3a6f474 = hmaster1_p & v3a6f9ff | !hmaster1_p & v374b0a3;
assign v3743dfc = hbusreq2 & v3a660f2 | !hbusreq2 & v8455ab;
assign v374c885 = hbusreq8_p & v8455ab | !hbusreq8_p & v380731d;
assign v3770f17 = hmaster0_p & v372707d | !hmaster0_p & v3761ae0;
assign v3752943 = hbusreq3 & v373dafc | !hbusreq3 & v8455ab;
assign v3a5ee7e = hbusreq8_p & v3a631f7 | !hbusreq8_p & v373ec80;
assign v373bfd3 = hmaster1_p & v3744280 | !hmaster1_p & v376abdf;
assign v375038a = hbusreq8_p & v3a60125 | !hbusreq8_p & v373042a;
assign v375dea9 = hgrant5_p & v372349f | !hgrant5_p & v3a6f389;
assign v3a57f8b = hgrant2_p & v8455ab | !hgrant2_p & v3766e8b;
assign v374e7f2 = hmaster3_p & v8455e1 | !hmaster3_p & !v375c7b9;
assign v373aec3 = hgrant5_p & v8455c6 | !hgrant5_p & v3a6f80b;
assign v3774cde = hgrant4_p & v3726139 | !hgrant4_p & v3a5e6b2;
assign v37413b6 = hbusreq6_p & v3a5408c | !hbusreq6_p & v3a5bb64;
assign v375789e = hmaster2_p & v3a6f8de | !hmaster2_p & v8455ab;
assign v3a6f7cd = hbusreq5_p & v3a62949 | !hbusreq5_p & !v3731d87;
assign v37392ad = hbusreq3_p & aadac1 | !hbusreq3_p & !v8455ab;
assign v3761136 = hbusreq0 & v3739ac1 | !hbusreq0 & v8455c9;
assign v3378a2d = hmaster2_p & v3a5e24e | !hmaster2_p & v3735e39;
assign v37470de = hgrant5_p & v8455ab | !hgrant5_p & v374bba3;
assign v373af5d = hbusreq6 & v37650bd | !hbusreq6 & v3377b1b;
assign v376efcc = hmaster0_p & v3a5f41b | !hmaster0_p & v37354da;
assign v3a60e6d = hbusreq8_p & v373951e | !hbusreq8_p & v8455ab;
assign v3a67458 = hgrant4_p & v3743c89 | !hgrant4_p & v373f94e;
assign v3761b24 = hmaster0_p & v37564a2 | !hmaster0_p & v3736d58;
assign v37617a9 = hbusreq6 & v3a70a23 | !hbusreq6 & v380701a;
assign v373a4f7 = hbusreq6 & v3a6fe3e | !hbusreq6 & v8455ab;
assign v2619ad7 = hbusreq5_p & v372da2f | !hbusreq5_p & v372bc6c;
assign v374fddd = hlock7_p & v3a66c34 | !hlock7_p & v374ac6d;
assign v3a6f60d = hmaster2_p & v3a635ea | !hmaster2_p & v373df13;
assign v3a70f67 = hgrant6_p & v3a2a8f2 | !hgrant6_p & v374aca8;
assign v37388aa = hmaster0_p & v374c582 | !hmaster0_p & v37559ec;
assign v38063c6 = hgrant3_p & v8455ab | !hgrant3_p & v377c0f5;
assign v3731f08 = hbusreq4 & v3a6ab69 | !hbusreq4 & v376bade;
assign v3a70a5f = hbusreq8_p & v3a5df33 | !hbusreq8_p & v375f97d;
assign v3a712a1 = jx3_p & v3a5f375 | !jx3_p & !v3a6eaea;
assign v3736439 = hgrant2_p & v8455ba | !hgrant2_p & v377b612;
assign v377a1ef = hbusreq5_p & v377beba | !hbusreq5_p & v8455ab;
assign v375b0e8 = hbusreq2 & v3a6c7c6 | !hbusreq2 & v3a70688;
assign v374cd48 = hbusreq2 & v377825c | !hbusreq2 & v374a637;
assign v3a5d882 = hbusreq4 & v3741afa | !hbusreq4 & v373abde;
assign v376e1ed = hbusreq2_p & v3730122 | !hbusreq2_p & v376cc20;
assign v3a5ae76 = hmaster2_p & v37416c6 | !hmaster2_p & v3a63a7a;
assign v3737ace = hmaster2_p & v8639e9 | !hmaster2_p & v8455ab;
assign v3764585 = hmaster2_p & v374c107 | !hmaster2_p & !v373c07d;
assign v373bfab = hbusreq0 & v3a6f7c7 | !hbusreq0 & v8455ab;
assign v37c0339 = hmaster1_p & v8455ab | !hmaster1_p & v373ccbc;
assign v376a272 = hlock4 & v3a625c9 | !hlock4 & v3723903;
assign v3a6430c = hbusreq1_p & v37748e5 | !hbusreq1_p & v38072fd;
assign v3746745 = hbusreq4_p & v377506b | !hbusreq4_p & v8455bb;
assign v376e611 = hbusreq1_p & v374473f | !hbusreq1_p & v376f455;
assign v376df25 = hmaster2_p & v3722e5c | !hmaster2_p & v3770559;
assign v3768633 = hbusreq6_p & v3a70a0e | !hbusreq6_p & v3738f5a;
assign v37233f1 = hlock5_p & v3a70b97 | !hlock5_p & v3a66514;
assign v3a70359 = hbusreq5 & v376a6f1 | !hbusreq5 & v373d35d;
assign v374176c = hmaster2_p & v373fe5e | !hmaster2_p & v8455e7;
assign v376b829 = hlock7_p & v3a70898 | !hlock7_p & !v8455ab;
assign v3764114 = hgrant2_p & v3a5baaf | !hgrant2_p & !v375e7d6;
assign v3777c9b = hbusreq7 & v375b56c | !hbusreq7 & v3a635ea;
assign v374f048 = jx1_p & v3a66039 | !jx1_p & v37479ee;
assign v3757955 = hgrant3_p & v3a708c2 | !hgrant3_p & v377ad8f;
assign v373d357 = hburst0 & v2aca977 | !hburst0 & v3a65f1f;
assign v3a70eea = hmaster1_p & v3725bdc | !hmaster1_p & v377b3ff;
assign v37335a5 = hgrant5_p & v8455c6 | !hgrant5_p & v37302fb;
assign v3a5d25d = hgrant5_p & v375e9ca | !hgrant5_p & v3a6f080;
assign v3a61a71 = hbusreq4 & v3a5f7d7 | !hbusreq4 & v3765e79;
assign v3a6c60e = hbusreq3_p & v3773ee6 | !hbusreq3_p & v3a617b4;
assign v3740380 = hbusreq7 & v3726e7b | !hbusreq7 & v376746b;
assign bdc54c = hbusreq3_p & v373ff4a | !hbusreq3_p & v37232bd;
assign v3766bbb = hbusreq7_p & v2092eb6 | !hbusreq7_p & v3a6f191;
assign v377eac7 = hgrant4_p & v374cd18 | !hgrant4_p & v37432d3;
assign v372e775 = jx1_p & v37474c1 | !jx1_p & v2092fa9;
assign v3a6ce42 = hgrant2_p & v3a6db06 | !hgrant2_p & v374ac3f;
assign v3a56338 = hgrant2_p & v3a6c80b | !hgrant2_p & v37300b7;
assign v37390c9 = hmaster2_p & v3a61b9c | !hmaster2_p & v3a57d9f;
assign v3a61d5f = hbusreq2_p & v374d13c | !hbusreq2_p & v3a53dbf;
assign v3a64eba = hbusreq5_p & v3727a16 | !hbusreq5_p & v3730fab;
assign v375582f = hbusreq4_p & v374d6dd | !hbusreq4_p & v37476fd;
assign v377795a = hmaster2_p & v35772a6 | !hmaster2_p & !v3761ad8;
assign v3737d23 = hgrant5_p & v3a7093f | !hgrant5_p & v372ddbc;
assign v37311fa = hmaster2_p & v3769ae2 | !hmaster2_p & v3730627;
assign v377eba4 = hgrant2_p & v3742c52 | !hgrant2_p & v3732bc0;
assign v3751b35 = hmaster2_p & v3743851 | !hmaster2_p & v375796c;
assign v3a70418 = hbusreq3_p & v3a551d6 | !hbusreq3_p & v3a640c5;
assign v3809b44 = hbusreq3 & v37407b3 | !hbusreq3 & v3733c39;
assign v373c590 = hlock8_p & v3734ed6 | !hlock8_p & v375e3fd;
assign v372475a = hbusreq0_p & v377c3fb | !hbusreq0_p & v8455ab;
assign v3732355 = hlock4 & v3807df0 | !hlock4 & v3a70bea;
assign v3a6f7c7 = hbusreq4 & v375911a | !hbusreq4 & v3a69487;
assign v373e10c = hgrant2_p & v377182c | !hgrant2_p & v373d440;
assign v3a70c55 = hlock4 & v3a6de95 | !hlock4 & v374cda0;
assign v3775f4f = hgrant6_p & v3a635ea | !hgrant6_p & v3809a8b;
assign v377c6d0 = hbusreq4_p & v3764702 | !hbusreq4_p & v37310be;
assign v3a6f1ab = hbusreq6_p & v3a70d99 | !hbusreq6_p & v2ff9314;
assign v376c652 = hmaster0_p & v3a6efcd | !hmaster0_p & v37374a1;
assign v3740a1b = hmaster0_p & v377c5f4 | !hmaster0_p & v373fc36;
assign v3761916 = hmaster1_p & v3a678de | !hmaster1_p & v35772a6;
assign v3749a46 = hbusreq7 & v3a6eace | !hbusreq7 & v373f537;
assign v373f9bf = hmaster2_p & v372c3df | !hmaster2_p & v3a6773a;
assign v3730a0f = hburst0_p & v8455ab | !hburst0_p & v845605;
assign v376c03e = hlock0_p & v3a5891c | !hlock0_p & !v3809adf;
assign v374bd09 = hbusreq4_p & v3762502 | !hbusreq4_p & v3a5bb64;
assign v3733dd4 = hbusreq3_p & v3739d22 | !hbusreq3_p & v376bb26;
assign v3a63e9b = hmaster0_p & v3759aeb | !hmaster0_p & v37481bf;
assign v377577b = hbusreq7_p & v375c1a7 | !hbusreq7_p & v3737808;
assign v373602d = hgrant1_p & v3743745 | !hgrant1_p & v8455ab;
assign v3743285 = hbusreq6_p & v3730bf5 | !hbusreq6_p & v3a70b55;
assign v3733fd8 = hgrant3_p & v3750d06 | !hgrant3_p & !v39eb517;
assign v37296f5 = hmaster0_p & v377bf37 | !hmaster0_p & v3760f64;
assign v377c71d = hmaster2_p & v3a59e1c | !hmaster2_p & v375d4e5;
assign v375e3d1 = hbusreq4_p & v374679f | !hbusreq4_p & v3a5e96b;
assign v372834d = hmaster0_p & v3a70967 | !hmaster0_p & dcb1a9;
assign v372c577 = hgrant0_p & v3a69ac0 | !hgrant0_p & v3a6d0ef;
assign v3a70924 = hbusreq5 & v3577324 | !hbusreq5 & !v3a5b955;
assign v3a6e089 = hbusreq4 & v3755dcd | !hbusreq4 & !v8455bd;
assign v3a6f291 = hmaster2_p & v37307dd | !hmaster2_p & v372ab46;
assign v3a5d6a6 = hgrant2_p & v374f617 | !hgrant2_p & v372a786;
assign v3a71196 = hmaster0_p & v3a61a7f | !hmaster0_p & v3807b28;
assign v37425a1 = hbusreq6_p & v374fe73 | !hbusreq6_p & v3779f13;
assign v8455d2 = hbusreq8 & v8455ab | !hbusreq8 & !v8455ab;
assign v3a70645 = hbusreq2_p & v3a5e7a5 | !hbusreq2_p & v3a6124f;
assign v3a616f0 = hbusreq7_p & v374e7b5 | !hbusreq7_p & v3a5f439;
assign v39ebb31 = hbusreq5 & v3746e94 | !hbusreq5 & v373a7ab;
assign v3a705f5 = hmaster0_p & v3a6f5c8 | !hmaster0_p & v3a296d8;
assign v3a67fd0 = hmaster1_p & v3a7119d | !hmaster1_p & v37702c5;
assign v375ed5a = hgrant0_p & v8455ab | !hgrant0_p & !v373b31d;
assign v374b320 = hgrant6_p & v8455ab | !hgrant6_p & v375f4e8;
assign v3769bdb = hgrant4_p & v373aca2 | !hgrant4_p & v3739815;
assign v3a60f18 = hbusreq0 & v373b548 | !hbusreq0 & v8455ab;
assign v373bb3a = hbusreq8 & v373763f | !hbusreq8 & v3a55e3c;
assign v3760da6 = hgrant5_p & v8455ab | !hgrant5_p & !v3723a94;
assign v3a70ca7 = hgrant6_p & v3a2a8f2 | !hgrant6_p & v3735134;
assign v3a6d8af = hmaster3_p & v373cb82 | !hmaster3_p & v372c7b7;
assign v375e21e = hbusreq5_p & v3770717 | !hbusreq5_p & v37723ce;
assign v373c897 = hmaster2_p & v373b30b | !hmaster2_p & v3a681ed;
assign v372cd1f = hmaster1_p & v374514e | !hmaster1_p & v376508b;
assign v372a2e4 = hbusreq7 & v376e66e | !hbusreq7 & v8455ab;
assign v3a5f891 = hbusreq5 & v38075cd | !hbusreq5 & v375495e;
assign v374f593 = hbusreq1 & v376430b | !hbusreq1 & v376653d;
assign v373fbc7 = hgrant3_p & v8455ab | !hgrant3_p & v377c31a;
assign v3a6eee7 = hlock7 & v3a5db58 | !hlock7 & v3736ae5;
assign v3378f5b = hbusreq8 & v3a7091e | !hbusreq8 & v3724665;
assign v37558f2 = hbusreq5_p & v3a70dbb | !hbusreq5_p & v3a65847;
assign v3a7157e = hgrant6_p & v8455ab | !hgrant6_p & v3731e3a;
assign v3a6f237 = hbusreq5 & v3759efd | !hbusreq5 & v3a7088b;
assign v3a6ebaa = hbusreq4 & v3757e28 | !hbusreq4 & v8455ab;
assign v3a6f786 = hmaster1_p & v8455ab | !hmaster1_p & v373a902;
assign v3760d59 = stateG2_p & v3a5a496 | !stateG2_p & v3a6446a;
assign v1e378a8 = hlock8 & v374a543 | !hlock8 & v3731455;
assign v3753dd4 = hgrant6_p & v373b687 | !hgrant6_p & v3a6d0a1;
assign v3a6006a = hlock2 & v3a670fe | !hlock2 & a36a2a;
assign v3764238 = hmaster1_p & v3776db0 | !hmaster1_p & v3762a54;
assign v3743eae = hbusreq6_p & v375e01c | !hbusreq6_p & !v8455ca;
assign v3a710c2 = hbusreq3 & v37317a9 | !hbusreq3 & v374f35a;
assign v376740b = hgrant5_p & v8455ab | !hgrant5_p & v3a70f06;
assign v3a5f714 = hmaster1_p & v3a67bce | !hmaster1_p & v3734d9a;
assign v372cedb = hbusreq2 & v39a5381 | !hbusreq2 & !v8455ab;
assign v376f01b = jx0_p & v373827a | !jx0_p & v376dd8b;
assign v3736e7c = hbusreq7 & v3731159 | !hbusreq7 & v8455bf;
assign v3a63c15 = hbusreq4_p & v3726d1f | !hbusreq4_p & v3749bf0;
assign v374d525 = hmaster0_p & v3a5c945 | !hmaster0_p & c60fa0;
assign v3745e29 = hbusreq8 & v3a55e75 | !hbusreq8 & v8455ab;
assign v3729dfc = hbusreq4_p & v3a65aeb | !hbusreq4_p & v9bbda1;
assign v3a68228 = hbusreq7_p & v374650b | !hbusreq7_p & v37434eb;
assign v3a70385 = hbusreq1_p & v39a5265 | !hbusreq1_p & v8455e1;
assign v3760e13 = jx0_p & v8455ab | !jx0_p & v3759628;
assign v380702c = hgrant5_p & v3a70746 | !hgrant5_p & v3a6da59;
assign v3728164 = hmaster2_p & v377ba55 | !hmaster2_p & v8455ab;
assign v3a70fdf = hbusreq6 & v3a6143b | !hbusreq6 & !v8455b5;
assign v376f167 = hgrant4_p & v8455ab | !hgrant4_p & v3a70f6b;
assign v37234e7 = hgrant1_p & v3759032 | !hgrant1_p & !v3809adf;
assign v3a68407 = hbusreq0 & v3722e90 | !hbusreq0 & v37248c1;
assign v37660f2 = hmaster2_p & v376eea3 | !hmaster2_p & v372a9c7;
assign v3a69892 = hmaster2_p & v3809ebc | !hmaster2_p & v3a5cfac;
assign c17a4a = hbusreq5 & v3728abd | !hbusreq5 & v8455ab;
assign v374eddc = hbusreq5 & v3740a1b | !hbusreq5 & v8455b3;
assign v3a6fb9f = hlock5_p & v376d9ad | !hlock5_p & v8455e7;
assign v3a6f2d9 = hgrant4_p & v8455e7 | !hgrant4_p & !v372516b;
assign v37312e2 = hbusreq2 & v3756bb9 | !hbusreq2 & v8455ab;
assign v3a60c77 = hbusreq1 & v3a54c77 | !hbusreq1 & v8455ab;
assign v377c348 = hgrant5_p & v8455ab | !hgrant5_p & v37294c5;
assign v37592d5 = hmaster1_p & v375b429 | !hmaster1_p & v37355c9;
assign v377c923 = hbusreq6_p & v37244a0 | !hbusreq6_p & v377efd0;
assign v3a65f15 = hbusreq1 & v39a5265 | !hbusreq1 & !v3a6ac2a;
assign v3a6fec1 = hmaster0_p & v3a71368 | !hmaster0_p & v375d2b3;
assign v3a5984d = hbusreq0 & v376c6a8 | !hbusreq0 & v3a64af7;
assign v3a5e357 = hbusreq0_p & v3807bf8 | !hbusreq0_p & v3a66110;
assign v37743e0 = hmaster2_p & v375808f | !hmaster2_p & v380881d;
assign v3727e10 = hgrant4_p & v8455ab | !hgrant4_p & v8455f5;
assign v3a6b4e8 = hmaster2_p & v377190a | !hmaster2_p & v3a56122;
assign v3a62072 = hgrant3_p & v3a6fab5 | !hgrant3_p & v35b9d52;
assign v3728493 = hmaster0_p & v3a617a6 | !hmaster0_p & v3764a7d;
assign v3773c13 = hlock7 & v3779097 | !hlock7 & v3727c74;
assign v3760592 = hmaster2_p & v3a2975f | !hmaster2_p & v8455ab;
assign v3a57384 = hbusreq0 & v3769e70 | !hbusreq0 & v3806f08;
assign v3a5edcb = hgrant2_p & v2092ac0 | !hgrant2_p & v37725f6;
assign v3743486 = hmaster2_p & v8455b2 | !hmaster2_p & v3754b66;
assign v375c7a3 = hbusreq8 & v3a6fbf6 | !hbusreq8 & v3734279;
assign v3a70a1a = hgrant3_p & v3752a0d | !hgrant3_p & v3777ca9;
assign v3a6ebdc = hbusreq7_p & v380910e | !hbusreq7_p & v3a70a46;
assign v3772409 = hbusreq5_p & v3a71097 | !hbusreq5_p & v3a5d644;
assign v3a6f40c = hlock0_p & ad2d05 | !hlock0_p & v3a58c79;
assign v37388f6 = hbusreq8 & v3776c6e | !hbusreq8 & a0a219;
assign v3772f85 = hgrant4_p & v3a56d26 | !hgrant4_p & v3a5e239;
assign v375abdb = hmaster0_p & v373dd7f | !hmaster0_p & v3a715c3;
assign v3a700a3 = hmaster0_p & v373bded | !hmaster0_p & v3a6ddea;
assign v3a57ac7 = hlock4 & v3a71037 | !hlock4 & v37285ad;
assign v37457c1 = hbusreq0_p & v3a7162d | !hbusreq0_p & v3778528;
assign v375e5d4 = hgrant3_p & v8455b0 | !hgrant3_p & dc6ea3;
assign v37566b2 = busreq_p & v39a537f | !busreq_p & !v3730dea;
assign v3757d20 = hbusreq3_p & v373128b | !hbusreq3_p & v373b288;
assign v3766c8c = hbusreq0_p & v3a70641 | !hbusreq0_p & v3733383;
assign v372919a = hbusreq0_p & v3a696ed | !hbusreq0_p & v8455ab;
assign v3728d14 = hbusreq0 & v3757559 | !hbusreq0 & !v1e37cd6;
assign v3a700e5 = hbusreq4 & v377d10c | !hbusreq4 & v3749bf0;
assign d0a687 = hlock1_p & v8455ab | !hlock1_p & v374e78f;
assign v3a6fdd2 = hlock4_p & v8455ab | !hlock4_p & v3a6ab5f;
assign v3a6c40f = hlock2_p & v3a7143c | !hlock2_p & v3739bb2;
assign v372fe58 = hmaster0_p & v37473af | !hmaster0_p & v3a6fd67;
assign v375ca6c = hbusreq2_p & v3a70dcd | !hbusreq2_p & v3a71567;
assign v3a707c2 = busreq_p & v3775476 | !busreq_p & !v372b3cf;
assign v3a62f8e = hlock8 & v3753942 | !hlock8 & v2092a89;
assign v3a70b35 = hmaster0_p & v2ff8ce3 | !hmaster0_p & v37341d3;
assign v37300c9 = hgrant3_p & v8455ab | !hgrant3_p & v3a6da33;
assign v3756cf0 = hgrant6_p & v3a700ae | !hgrant6_p & v3a701a9;
assign v37751ae = hmaster3_p & v3729440 | !hmaster3_p & v8455ab;
assign v3a6f46a = hbusreq2_p & v37700b9 | !hbusreq2_p & v372d490;
assign v37629d2 = jx1_p & v3a53a43 | !jx1_p & v37383bb;
assign v3a57fff = hbusreq6_p & v377803a | !hbusreq6_p & v37597a4;
assign v372a96f = hmaster2_p & v376a6f1 | !hmaster2_p & !v3776f5e;
assign v3a71424 = hbusreq1 & v39a537f | !hbusreq1 & v8455ab;
assign v3a55838 = hgrant6_p & v372879a | !hgrant6_p & v3777cb9;
assign v376d92b = hbusreq0 & v377c023 | !hbusreq0 & v3a5621f;
assign v374e248 = hlock0_p & v374f0c1 | !hlock0_p & v377f6ff;
assign v372b840 = hmaster2_p & v376653d | !hmaster2_p & !v8455e7;
assign v375e3fd = hmaster1_p & v3a6ffae | !hmaster1_p & v373cd5a;
assign v374677f = hmaster0_p & v8455ab | !hmaster0_p & v3737d2f;
assign v3733d45 = hbusreq4 & v372b7cc | !hbusreq4 & v8455ab;
assign v3724069 = hlock2 & v3748797 | !hlock2 & v377bbbb;
assign v3a70620 = hmaster0_p & v35b774b | !hmaster0_p & v3773b18;
assign v3735da7 = hmaster1_p & v372d24a | !hmaster1_p & v3a2abf4;
assign v3a5e6b2 = hgrant6_p & v3726139 | !hgrant6_p & v3725bea;
assign v3779412 = hgrant6_p & v8455ab | !hgrant6_p & v3724e98;
assign v3778b48 = hbusreq5_p & v37286f3 | !hbusreq5_p & v377b429;
assign v3724fe7 = hgrant6_p & v3a5c5fc | !hgrant6_p & v3808eaa;
assign v374d03f = hmaster1_p & v8455ab | !hmaster1_p & v376f4a6;
assign v373fcbf = hmaster0_p & v372ed51 | !hmaster0_p & v376a40d;
assign v3753542 = hmaster0_p & v375c791 | !hmaster0_p & v373d7e9;
assign v37581c0 = hlock3_p & v3a6c467 | !hlock3_p & v8455b0;
assign v37554d5 = hbusreq4 & v376489a | !hbusreq4 & v8455ab;
assign v37690ea = hlock6 & v3773a5b | !hlock6 & v3732706;
assign v3754c51 = hmaster0_p & v37295e7 | !hmaster0_p & v3a70d99;
assign v373d69f = hmaster2_p & v3a712c4 | !hmaster2_p & v376112d;
assign v3733940 = hmaster2_p & v37306c2 | !hmaster2_p & v3a71631;
assign bef73a = hbusreq1_p & v374ed4b | !hbusreq1_p & !v3a54bcd;
assign v3a68b34 = hbusreq6 & v3a6910c | !hbusreq6 & v8455ab;
assign v3a5f8b6 = hgrant8_p & v8455ab | !hgrant8_p & v376dd91;
assign v3a6ec20 = hmaster0_p & v37386c6 | !hmaster0_p & v3a68482;
assign ae317f = hbusreq6 & v374b65e | !hbusreq6 & !v8455ab;
assign v3a5ef89 = hlock2 & v3a65da2 | !hlock2 & v3a70923;
assign v3a65a19 = hbusreq4 & v3746b4f | !hbusreq4 & v8455e7;
assign bbba6b = hmaster2_p & v3a714fd | !hmaster2_p & v3a5be15;
assign v3a6bf86 = hbusreq2_p & v376e238 | !hbusreq2_p & v3a7052a;
assign v3a704b4 = hmaster2_p & v3a5e24e | !hmaster2_p & !v3759032;
assign v375cd3f = hbusreq8_p & v92aebd | !hbusreq8_p & v376c712;
assign v3a61132 = hbusreq7_p & v3a70307 | !hbusreq7_p & v373eb03;
assign v3a6fc77 = hbusreq5 & v3a60691 | !hbusreq5 & aa9893;
assign v376773f = hbusreq4_p & v3a709e1 | !hbusreq4_p & v8455ab;
assign v3745d14 = hbusreq5 & v3768429 | !hbusreq5 & !v372c051;
assign v3a63659 = hgrant4_p & v3a5a03f | !hgrant4_p & v374ebb0;
assign v3a6ef5a = hgrant4_p & v8455c2 | !hgrant4_p & v376269a;
assign v3a637a5 = hgrant5_p & v37712fa | !hgrant5_p & v376b1b7;
assign v374c8b8 = hbusreq5_p & v3a6be05 | !hbusreq5_p & v37511c6;
assign v373fd51 = hbusreq8_p & v37380d5 | !hbusreq8_p & !v376c4fd;
assign v3763832 = hbusreq7_p & v3752aa3 | !hbusreq7_p & v37470de;
assign v3730f7e = hmaster2_p & v3756f10 | !hmaster2_p & !v374cb97;
assign v374f968 = hgrant4_p & v3735cb3 | !hgrant4_p & v3a6ad00;
assign v3740f70 = hgrant3_p & v8455e7 | !hgrant3_p & !bd3213;
assign v3730601 = hmaster2_p & v3a637dc | !hmaster2_p & !v8455ab;
assign v3733bfc = hbusreq5_p & v374a1f5 | !hbusreq5_p & v3a53c18;
assign v3774dcd = hmaster1_p & v3577306 | !hmaster1_p & v3a700a6;
assign v3759119 = hbusreq4_p & v37259cc | !hbusreq4_p & v374dce0;
assign v377b59e = hmaster2_p & v3740161 | !hmaster2_p & v3a7106c;
assign v3a64ff4 = hmaster0_p & v377ce1a | !hmaster0_p & v3a6dd80;
assign v3a67fb5 = jx0_p & v3a70df5 | !jx0_p & v37490d7;
assign v3a6817f = hmaster2_p & v3736d47 | !hmaster2_p & v37297cb;
assign v3733739 = hbusreq8_p & v3a606d2 | !hbusreq8_p & v3746976;
assign v3a6f9ab = hmaster2_p & v3a619c0 | !hmaster2_p & !v37282cf;
assign v3a67d6f = hbusreq0_p & v3a57309 | !hbusreq0_p & v8455ab;
assign v374e409 = hmaster2_p & v8455e1 | !hmaster2_p & !v375c7b9;
assign v3762079 = hbusreq5 & v3a66bc6 | !hbusreq5 & v3a60594;
assign v3a6f151 = hgrant2_p & v8455ab | !hgrant2_p & v3774346;
assign v372b02f = hbusreq4_p & v3768e70 | !hbusreq4_p & v3a66ac0;
assign v3a5fe39 = hbusreq6_p & v3a70b1e | !hbusreq6_p & v8455ab;
assign v3746b22 = hmaster1_p & v3a7002c | !hmaster1_p & v2acafb4;
assign v3a6f48e = hbusreq5 & v3a6f87e | !hbusreq5 & v8455ab;
assign v3a66615 = hmaster2_p & v3776715 | !hmaster2_p & v376f409;
assign v376fbe0 = hgrant4_p & v3729dfc | !hgrant4_p & v37511a1;
assign v37790a9 = hgrant3_p & v3759b2f | !hgrant3_p & v3a6edb1;
assign v374a0ac = hmaster0_p & v37572d0 | !hmaster0_p & v3a6ef24;
assign v375fb86 = jx1_p & v3776e23 | !jx1_p & v3724976;
assign v3740cd2 = hmaster1_p & v3a60dfb | !hmaster1_p & v3731349;
assign v3809561 = hbusreq5 & v374fb30 | !hbusreq5 & v372e885;
assign v372cb42 = hgrant2_p & v8455ab | !hgrant2_p & v3a5ce6f;
assign v3a7073b = hlock4 & v376a149 | !hlock4 & v375b18e;
assign v3730370 = hmaster0_p & v3727e69 | !hmaster0_p & v3767e71;
assign v37577d8 = hlock3 & v3a5a985 | !hlock3 & v3a670d6;
assign v35b710e = hlock4_p & v3a568f7 | !hlock4_p & v373c755;
assign v3a5df70 = hmaster1_p & v3a5fc34 | !hmaster1_p & v376f321;
assign v372dab1 = locked_p & v380775e | !locked_p & v3a6ffae;
assign v3a6e7a7 = hlock0_p & v3a70fc0 | !hlock0_p & v3a6ae99;
assign v3a5ddee = hlock2_p & v3772ad5 | !hlock2_p & v8455b0;
assign v376a480 = hmaster2_p & v3a635ea | !hmaster2_p & v375e854;
assign v376e663 = hlock8 & v3772d2f | !hlock8 & v3765f12;
assign v3a5a3d0 = hlock7 & v3a59eab | !hlock7 & v3a587a1;
assign v3768d47 = hbusreq6_p & v3736a9a | !hbusreq6_p & v3a5ee12;
assign v3a701e7 = hgrant3_p & v37331e7 | !hgrant3_p & v373be9e;
assign v37785b8 = hbusreq4_p & v37506d6 | !hbusreq4_p & !v8455ab;
assign v37479c3 = hgrant5_p & v3765e47 | !hgrant5_p & v3a63717;
assign v3a71392 = jx1_p & v373c071 | !jx1_p & v3759ff9;
assign v3a55cd6 = hbusreq3_p & v3a6143b | !hbusreq3_p & !v39a4ca8;
assign v373d932 = hbusreq3_p & v3a54344 | !hbusreq3_p & v3a5cd20;
assign v3755783 = hmaster1_p & v3763f95 | !hmaster1_p & v3a70820;
assign v377c8fd = hmaster0_p & v3a6ffb6 | !hmaster0_p & v3a5ace8;
assign v37331ef = hgrant3_p & v37669b4 | !hgrant3_p & v3777962;
assign v3a6f4e8 = hbusreq6_p & v3768a88 | !hbusreq6_p & v3779d86;
assign v3760bc2 = hmaster0_p & v375725f | !hmaster0_p & v3776b20;
assign v37369d7 = hmaster2_p & v37590a2 | !hmaster2_p & v3756304;
assign v3a71305 = hbusreq7_p & v8455cb | !hbusreq7_p & v375830c;
assign v3724048 = hbusreq4 & v37281e7 | !hbusreq4 & v23fdaed;
assign v3750ba3 = hlock5 & v37437cf | !hlock5 & v3a568ee;
assign v3751094 = stateA1_p & v8455ab | !stateA1_p & v3a6efc4;
assign v3a6f43a = hbusreq6_p & v375da82 | !hbusreq6_p & v3725717;
assign v3a5aaca = hbusreq5_p & v3748400 | !hbusreq5_p & v373c688;
assign v377bfc7 = hmaster2_p & v3770b26 | !hmaster2_p & v3745b02;
assign v377a7ee = hbusreq7_p & a0a219 | !hbusreq7_p & v377696e;
assign v3a704de = hlock4 & v38072fd | !hlock4 & v3a6cb62;
assign v3752707 = hbusreq4 & v376e89b | !hbusreq4 & v3a70d99;
assign v375792c = hmaster0_p & v8455ab | !hmaster0_p & v375f6c7;
assign v3a703a9 = jx3_p & v376b5f2 | !jx3_p & d5c12b;
assign v3a6ff71 = hmaster0_p & v3a5af94 | !hmaster0_p & !v3a6ef21;
assign v3734dc5 = jx0_p & v374edb8 | !jx0_p & v3762bdf;
assign v373d9d3 = hgrant6_p & v37304b3 | !hgrant6_p & v3a548f2;
assign v3a640a0 = hbusreq6_p & v8455ca | !hbusreq6_p & !v8455ab;
assign v3741cd4 = jx1_p & v377e0a4 | !jx1_p & v37705be;
assign v3a605f1 = hlock6 & v3723baf | !hlock6 & v3a56d0a;
assign v39a53a4 = hgrant6_p & v373c81c | !hgrant6_p & v3a6f4ef;
assign v372aaf8 = hmaster1_p & v3a635ea | !hmaster1_p & v372d4eb;
assign v1e37481 = hmastlock_p & v3a62251 | !hmastlock_p & v8455ab;
assign v3766809 = jx1_p & v374bf69 | !jx1_p & v3a5a25a;
assign v3766e5d = hgrant3_p & v3a61cbf | !hgrant3_p & v376a7fc;
assign v37432e2 = hmaster2_p & v376111d | !hmaster2_p & !v37583be;
assign v376c490 = hgrant6_p & v377f09a | !hgrant6_p & !be2682;
assign v37474df = hbusreq5 & v376d76c | !hbusreq5 & v3756996;
assign v3768c98 = hbusreq7_p & v3a70c90 | !hbusreq7_p & v372cf51;
assign v376a2c0 = hgrant4_p & v3757568 | !hgrant4_p & v37753e0;
assign v37617ed = hmaster2_p & v8455ab | !hmaster2_p & v377a9a1;
assign v376e3a0 = hmaster0_p & v3757f09 | !hmaster0_p & v3a6f13e;
assign v372c23f = jx0_p & v3750e4f | !jx0_p & v37322d8;
assign v3a6d2ae = hbusreq6 & v3a7151d | !hbusreq6 & !v8455ab;
assign v3768358 = hmaster2_p & v372cac6 | !hmaster2_p & v374448e;
assign v372bc4c = hbusreq5_p & v3a6be05 | !hbusreq5_p & v3745734;
assign v3734b15 = hbusreq2 & v3a69d81 | !hbusreq2 & v37360b3;
assign v3a6600c = hbusreq6 & v3a7045b | !hbusreq6 & v8455ab;
assign v3765fcf = hbusreq6_p & v3a6f3a8 | !hbusreq6_p & !v3a658bf;
assign v377bdc3 = hgrant4_p & v3739791 | !hgrant4_p & !v8455ab;
assign v375d707 = hgrant2_p & v375c55a | !hgrant2_p & v3a6fd82;
assign v37634d0 = hbusreq5 & v372ab6c | !hbusreq5 & v3730370;
assign v3730722 = hbusreq5 & v3a5ed86 | !hbusreq5 & v3a5584b;
assign v3742a8b = hmaster0_p & v3764276 | !hmaster0_p & v3a6f774;
assign v3774af1 = hgrant7_p & v3a60ac5 | !hgrant7_p & v376f468;
assign v376ca61 = hmaster1_p & v3a71585 | !hmaster1_p & v377d080;
assign v37503e7 = hgrant7_p & v8455ab | !hgrant7_p & v37556ce;
assign v37438b9 = hbusreq6_p & v3722d81 | !hbusreq6_p & v8455ab;
assign v3a6c0c1 = hmaster1_p & v376eed8 | !hmaster1_p & v377a27c;
assign v3a691ca = hbusreq7_p & v3737456 | !hbusreq7_p & v3a71094;
assign v3767c03 = hmaster3_p & v3742825 | !hmaster3_p & v8455ab;
assign v376d1b4 = hbusreq5_p & v375820a | !hbusreq5_p & v8455ab;
assign v3a61298 = hgrant3_p & v8455e7 | !hgrant3_p & !v3a70524;
assign v373e30f = hbusreq5_p & v3a5f453 | !hbusreq5_p & !v8455ab;
assign v376cfc1 = hmaster2_p & v3a70f1c | !hmaster2_p & v3758f19;
assign v3a7161b = hmaster0_p & v3a7022c | !hmaster0_p & v373185b;
assign v373fbca = hgrant2_p & v8455ab | !hgrant2_p & v37249f1;
assign v37348f5 = hmaster1_p & v3a63d77 | !hmaster1_p & v376b27a;
assign v3743792 = hmaster0_p & v375e6a0 | !hmaster0_p & v37691e2;
assign v3a6f1eb = hmaster1_p & v377d1dc | !hmaster1_p & v374e0b8;
assign v373a246 = hmaster2_p & v3744981 | !hmaster2_p & v3a5b68a;
assign v3a5a24b = hgrant4_p & v3577306 | !hgrant4_p & v3a71599;
assign v37510e0 = hlock4 & v3a6f88b | !hlock4 & v3735d39;
assign v3749cdf = hbusreq0 & v3723b86 | !hbusreq0 & v8455ab;
assign v376e2ac = hbusreq6 & v374704d | !hbusreq6 & v8455ab;
assign v372fc6c = hmaster0_p & v377e630 | !hmaster0_p & v377b556;
assign v3768264 = hbusreq3_p & v3752ec0 | !hbusreq3_p & v3a66b26;
assign v373b599 = hmaster2_p & v3a6fe0d | !hmaster2_p & !v3a5e817;
assign v3738766 = hbusreq2_p & v3a29842 | !hbusreq2_p & v3a5759a;
assign v3765576 = hbusreq4_p & v3745241 | !hbusreq4_p & v3745ce8;
assign v376d081 = hgrant2_p & v3a65827 | !hgrant2_p & v3754f5d;
assign v3742e54 = hmaster1_p & v3746c51 | !hmaster1_p & v3750d8e;
assign v375745a = hmaster3_p & v373a494 | !hmaster3_p & v3761912;
assign v375185f = hgrant2_p & v37543d8 | !hgrant2_p & v37725f6;
assign v377cdee = hbusreq6 & v3776db6 | !hbusreq6 & v1e37a04;
assign v3a6f737 = hbusreq7_p & v3a565bc | !hbusreq7_p & v3a6f3dc;
assign v3a663c7 = hgrant2_p & v375ca6c | !hgrant2_p & v2acaeb7;
assign v3a69677 = hbusreq7 & v3a6bedd | !hbusreq7 & v372f464;
assign v375f2ec = hbusreq6_p & v375306b | !hbusreq6_p & v3756b48;
assign v3a5818a = hbusreq4_p & v373510a | !hbusreq4_p & v8455ab;
assign b6057e = hmaster1_p & v3a6f443 | !hmaster1_p & v3a694b4;
assign v3a6f417 = hbusreq5_p & v3a635ea | !hbusreq5_p & v374457a;
assign v373f4cf = hmaster1_p & v372ed89 | !hmaster1_p & v3a6f601;
assign v3a6bde4 = hbusreq8 & v3754eb4 | !hbusreq8 & v8455ab;
assign v377ee58 = hgrant0_p & v375c7b9 | !hgrant0_p & v3a635ff;
assign v845765 = hmaster1_p & v3759031 | !hmaster1_p & v3a6fb8d;
assign v372f236 = hgrant6_p & v3a61e59 | !hgrant6_p & v3a705fb;
assign v3a674b3 = hmaster0_p & v3748360 | !hmaster0_p & v37281fb;
assign ab60dc = hgrant3_p & v3577306 | !hgrant3_p & v3747cdb;
assign v3a56114 = jx1_p & v3a5aa42 | !jx1_p & v372d417;
assign v3731685 = hbusreq4 & v376c87d | !hbusreq4 & v3756eca;
assign v372cb8c = hmaster0_p & v3729bc6 | !hmaster0_p & v3a70c2c;
assign v3a6fe10 = hbusreq7 & v23fe0ff | !hbusreq7 & v3a6fd20;
assign v1e37523 = hgrant4_p & v8455ab | !hgrant4_p & v3731230;
assign v3a689e5 = hmaster0_p & v37393ad | !hmaster0_p & v3a6fe1b;
assign v3767d4e = hbusreq3 & v3a6ab5f | !hbusreq3 & !v3a6ac2a;
assign v372871c = hgrant5_p & v372c334 | !hgrant5_p & v3776352;
assign v374fe49 = hmaster1_p & cfaa3a | !hmaster1_p & v3735bbc;
assign v3a711e4 = hmaster2_p & v37745a0 | !hmaster2_p & v373698e;
assign v1e37a06 = hmaster0_p & v3a62fc6 | !hmaster0_p & v376730a;
assign v3a6f6de = hbusreq1_p & v374fc6c | !hbusreq1_p & v8455b0;
assign v3740dcd = hbusreq2 & v37468ea | !hbusreq2 & v372e83f;
assign v37491b7 = hgrant3_p & v8455bd | !hgrant3_p & v375b65b;
assign v37315da = hbusreq6_p & v3a5ff09 | !hbusreq6_p & v8455ab;
assign v3727517 = hlock0_p & v3759b2f | !hlock0_p & !v373be25;
assign v3a70d72 = hbusreq8_p & v37546a4 | !hbusreq8_p & v37334ff;
assign v3779d96 = hmaster1_p & v8455ab | !hmaster1_p & v373e60c;
assign v37725f6 = hbusreq2_p & v3760279 | !hbusreq2_p & v376c747;
assign v376bce3 = hbusreq8_p & v374bc20 | !hbusreq8_p & v372f434;
assign v372ff09 = hmaster2_p & v3a6fc7f | !hmaster2_p & v3727472;
assign v377881b = hlock3 & v3a711fb | !hlock3 & v37774c7;
assign v376dd64 = hlock5 & v3806498 | !hlock5 & v3764c7c;
assign v37378e5 = hbusreq4 & v373127e | !hbusreq4 & v8455bf;
assign v3a647e2 = hbusreq6 & v8455b0 | !hbusreq6 & v3a63805;
assign v3775165 = hgrant2_p & v3750269 | !hgrant2_p & v37306d8;
assign v372c2da = hbusreq5 & v37566b2 | !hbusreq5 & !v8455ab;
assign v3a65260 = hbusreq5_p & v377eada | !hbusreq5_p & v3a71677;
assign v3377b1b = hgrant2_p & v37496fa | !hgrant2_p & v3a6fefa;
assign v3a70f2c = hmaster3_p & v375076f | !hmaster3_p & v3a6ae54;
assign aeaf7c = hmaster1_p & v3a5e24e | !hmaster1_p & v374083d;
assign v3a613e6 = hbusreq5_p & v377efe1 | !hbusreq5_p & v37577ab;
assign v37377df = hmaster2_p & v3728c23 | !hmaster2_p & v376b4ad;
assign v3a5b945 = jx3_p & v37645aa | !jx3_p & v372b3b6;
assign v3757863 = hgrant4_p & v376f0fb | !hgrant4_p & v377d60e;
assign v3a6ebe8 = hlock8_p & v3730b84 | !hlock8_p & v3a6bde4;
assign v373172e = hmaster1_p & v8455e7 | !hmaster1_p & v377a975;
assign v3723fce = hgrant6_p & v8455ab | !hgrant6_p & v37412c3;
assign c3d672 = hgrant6_p & v3a5cb45 | !hgrant6_p & v377459d;
assign v37301dd = hmaster0_p & v374ac8c | !hmaster0_p & v374f397;
assign v3752c61 = hbusreq2 & v374ed4f | !hbusreq2 & v3770751;
assign v377d6d3 = hbusreq4 & v376b57f | !hbusreq4 & v373bd6c;
assign v3723299 = hbusreq4_p & c7d127 | !hbusreq4_p & v373683d;
assign v3756fbd = hmaster0_p & v37685c3 | !hmaster0_p & v3a7026a;
assign v3a70abb = hgrant5_p & v8455c6 | !hgrant5_p & b9f306;
assign v3a6a322 = hbusreq6 & v374d8bb | !hbusreq6 & v377c6b3;
assign v3a7032a = hmaster2_p & v376e72d | !hmaster2_p & v8455cb;
assign v37251c9 = hbusreq5 & v3732f19 | !hbusreq5 & v375b0ad;
assign v37435f7 = hlock0 & v38072fd | !hlock0 & v37237cd;
assign v3755f23 = hlock7 & v3748d3c | !hlock7 & v3771633;
assign v3a70235 = hmaster2_p & v8455ab | !hmaster2_p & v377a657;
assign v374efee = hbusreq3_p & v3768b81 | !hbusreq3_p & v3a627d8;
assign v3a6d2d3 = hmaster0_p & v375fb93 | !hmaster0_p & v8455b5;
assign v3a6fde6 = hbusreq7 & v3a656dd | !hbusreq7 & v3724e14;
assign v35b7808 = hready & v8455ab | !hready & v3730cce;
assign v376aeae = hlock2 & v376121f | !hlock2 & v375d009;
assign v3a675b2 = hmaster3_p & v37303aa | !hmaster3_p & v372c353;
assign v3a55271 = stateG10_1_p & v8455ab | !stateG10_1_p & a9f810;
assign v3742cde = hbusreq2_p & v376c63d | !hbusreq2_p & v8455ab;
assign v377700a = hmaster2_p & v377c9bd | !hmaster2_p & v3a5a807;
assign v3753386 = hbusreq1_p & v377b24b | !hbusreq1_p & v3577306;
assign v3774f3b = hbusreq4 & v39a4ca8 | !hbusreq4 & v8455b5;
assign v3743eb5 = hbusreq3_p & v3749b84 | !hbusreq3_p & v377c31a;
assign v3a6f687 = hbusreq6_p & v3769f88 | !hbusreq6_p & v3a5da57;
assign v3739531 = hmaster0_p & v3725098 | !hmaster0_p & v373ad3f;
assign v3a7075d = hbusreq8 & v3a70080 | !hbusreq8 & v3a703ba;
assign v3773804 = hmaster2_p & v8455ab | !hmaster2_p & !v377ea86;
assign v374bf59 = hgrant6_p & v380649c | !hgrant6_p & v3a55630;
assign v373296d = hmaster2_p & v3a70557 | !hmaster2_p & v3a6fa93;
assign v377acae = hlock4_p & v3a709ea | !hlock4_p & v3a70131;
assign v377234d = hbusreq4_p & v3759886 | !hbusreq4_p & v8455ab;
assign v3a66f3e = hbusreq0 & v37321c2 | !hbusreq0 & v372d48a;
assign v3a5f1db = hbusreq7_p & v373f1ba | !hbusreq7_p & v376b70a;
assign v372ee0e = hbusreq6_p & v3a59424 | !hbusreq6_p & !v8455ab;
assign v3a6f856 = hbusreq4 & v37739f4 | !hbusreq4 & !v37531b1;
assign v3767651 = jx3_p & v3a6756b | !jx3_p & v3a70e5f;
assign v3a5bcc4 = hmaster1_p & v3a566eb | !hmaster1_p & d6db19;
assign v3748645 = hbusreq2 & v3748e81 | !hbusreq2 & v8455ab;
assign v377ee3c = hbusreq6_p & v8455ab | !hbusreq6_p & v3724577;
assign v3732e09 = hmaster2_p & v3a6854c | !hmaster2_p & v3a6ea66;
assign v3742370 = hgrant2_p & v8455ab | !hgrant2_p & v3a66d7b;
assign v3a6facb = hmaster2_p & v377234d | !hmaster2_p & v3724270;
assign v3741863 = hlock7 & v3a6f92d | !hlock7 & v374c297;
assign v3a5b05d = hbusreq5_p & v372834d | !hbusreq5_p & v35ba1cf;
assign v373cd0c = hgrant4_p & v37585bf | !hgrant4_p & !v37541d3;
assign v3a71654 = hmaster2_p & v3769740 | !hmaster2_p & be54b2;
assign v374fef8 = stateG10_1_p & v3751fa8 | !stateG10_1_p & v3a610e9;
assign v35b70ed = hmaster1_p & v3769093 | !hmaster1_p & v372ef56;
assign v3a68391 = hgrant8_p & v8455ab | !hgrant8_p & !v3742441;
assign v373dcb0 = hgrant1_p & v3771ee8 | !hgrant1_p & v3740171;
assign v372452c = hbusreq0 & v1e37a72 | !hbusreq0 & v3a6ebae;
assign v3806f21 = hbusreq7_p & v375ec1d | !hbusreq7_p & v8455ab;
assign v3735f30 = hgrant5_p & v8455ab | !hgrant5_p & v3a70b13;
assign v3a70d99 = hbusreq2_p & v3a61a3d | !hbusreq2_p & v8455ab;
assign v372642c = hbusreq4_p & v373ee51 | !hbusreq4_p & !v8455ab;
assign v377b68e = hgrant6_p & v377938d | !hgrant6_p & v374b8ad;
assign v3a6ef70 = hbusreq8 & v3772aaf | !hbusreq8 & v3773c40;
assign v3a66e30 = hmaster2_p & v372edf8 | !hmaster2_p & v3a5c562;
assign v3750bc4 = hmaster1_p & v372b4b4 | !hmaster1_p & v3a7152a;
assign v372dbf1 = hbusreq3 & v3746f84 | !hbusreq3 & v8455ab;
assign v3a70fea = hlock7 & v377c2bc | !hlock7 & v377f5ca;
assign v3a71024 = hbusreq0 & v3a70b83 | !hbusreq0 & v37644e0;
assign v3762e13 = hgrant4_p & v8455ab | !hgrant4_p & v3a5818a;
assign v3a70381 = hmaster0_p & v23fe361 | !hmaster0_p & v3730930;
assign v373fb40 = hbusreq7_p & v375d849 | !hbusreq7_p & v3a61bef;
assign stateG10_6 = !v3985143;
assign v3755c31 = hbusreq3_p & v3a6fdb4 | !hbusreq3_p & v372ade8;
assign v2889706 = hbusreq5 & v3a5cd4c | !hbusreq5 & v8455ab;
assign v3746caf = hbusreq2_p & v3730c69 | !hbusreq2_p & v372554a;
assign v3753f1d = hmaster0_p & v372d866 | !hmaster0_p & v3769820;
assign v3741736 = hmaster1_p & v8455ab | !hmaster1_p & v360d00f;
assign v375e1b0 = hmaster2_p & v3a635ea | !hmaster2_p & v37786a6;
assign v373ad8b = hlock5_p & v3a6ff3e | !hlock5_p & v3761472;
assign v3760c90 = hgrant2_p & v375c7b9 | !hgrant2_p & v373bb2d;
assign v3a6c2d4 = hgrant3_p & v8455ab | !hgrant3_p & v3737f89;
assign v3733ec6 = hlock1_p & v8455ab | !hlock1_p & !v8455b6;
assign v3a6eafe = hbusreq7_p & v37249fe | !hbusreq7_p & v3a6054b;
assign v3a7105f = hbusreq5 & v3745aae | !hbusreq5 & v3a61b59;
assign v3a56f9d = hlock5_p & v3a70099 | !hlock5_p & v3757cd1;
assign v3740bcb = hmaster2_p & v3774f38 | !hmaster2_p & !v8455ab;
assign v37455ec = hgrant0_p & v37262fd | !hgrant0_p & v374288a;
assign v3735112 = hgrant6_p & v3764486 | !hgrant6_p & v37376c1;
assign v37777a2 = hbusreq3_p & v3733d6e | !hbusreq3_p & v372ee7e;
assign v3a71166 = hlock0 & v3a6f71a | !hlock0 & v3729fa0;
assign v373d0a3 = hmaster2_p & v3a5600a | !hmaster2_p & v37685bb;
assign v3774452 = hgrant5_p & v3a6f1d8 | !hgrant5_p & v3727a04;
assign v3a70f5f = jx1_p & v374b237 | !jx1_p & v8455ab;
assign v3776ada = hgrant4_p & v8455ab | !hgrant4_p & v3763b0a;
assign v3a6f718 = hbusreq2_p & v377cece | !hbusreq2_p & v376bb26;
assign v375455d = hmaster1_p & v377766c | !hmaster1_p & v3756bde;
assign v3a61b59 = hmaster0_p & v3a7074d | !hmaster0_p & v37789ca;
assign v376b15b = hbusreq6_p & v3a5b289 | !hbusreq6_p & v2619b43;
assign v3a2976c = hmaster0_p & v2093018 | !hmaster0_p & v3a71498;
assign v3a6fd5e = hbusreq4_p & v37315c8 | !hbusreq4_p & v3756918;
assign v94335e = hbusreq7 & v3a5d25d | !hbusreq7 & v3774452;
assign v3a678de = hmaster0_p & v373bdd1 | !hmaster0_p & v35772a6;
assign v8455c2 = hbusreq4 & v8455ab | !hbusreq4 & !v8455ab;
assign v3738826 = hbusreq5_p & v3a70252 | !hbusreq5_p & v37435fd;
assign dab321 = hbusreq3_p & v375bd1f | !hbusreq3_p & v377696a;
assign v3a6818c = hbusreq7 & v3747b55 | !hbusreq7 & c5ed52;
assign v3a7046b = hlock4 & v3724e2a | !hlock4 & v374dffc;
assign v3769e7f = hbusreq4_p & v3765370 | !hbusreq4_p & v38072fd;
assign v374fedc = hmaster0_p & v3a6fc3a | !hmaster0_p & !v3775f27;
assign v37797a3 = hlock2_p & v8455ab | !hlock2_p & v373fe5e;
assign v3760eeb = hbusreq4_p & v3740171 | !hbusreq4_p & v37457fb;
assign v375acae = hmaster1_p & v3a61397 | !hmaster1_p & v3a71036;
assign v372fef2 = hmaster1_p & v37782c9 | !hmaster1_p & v375f2b3;
assign v373b4c8 = hbusreq8_p & v3a665b4 | !hbusreq8_p & v3745498;
assign v373e284 = hgrant5_p & v3a6f6af | !hgrant5_p & v37660d9;
assign v3a712f5 = hbusreq7 & v3779593 | !hbusreq7 & v372fdd0;
assign v3a704b8 = hmaster1_p & v913004 | !hmaster1_p & !v374cab1;
assign v3a7111f = stateG3_2_p & v8455ab | !stateG3_2_p & v3725f3b;
assign v3778277 = hmaster2_p & v372aafb | !hmaster2_p & !v3750b61;
assign v374b962 = hbusreq0_p & v8455ab | !hbusreq0_p & !v3a637dd;
assign v3765c49 = hlock5 & v3751ffd | !hlock5 & v37572af;
assign v3a6ffbc = hbusreq5 & v373568b | !hbusreq5 & v376c5b2;
assign v377aed1 = hmaster0_p & v37571c8 | !hmaster0_p & v3a6d897;
assign v3a6ef24 = hmaster2_p & v37256d2 | !hmaster2_p & v373a303;
assign v3a65ce7 = hmaster0_p & v3a614a1 | !hmaster0_p & v376cd84;
assign v372e25b = hbusreq4_p & v373a141 | !hbusreq4_p & v372a116;
assign v3769980 = hmaster1_p & v3a7028a | !hmaster1_p & v3779958;
assign v3a715ea = hbusreq5_p & v3775393 | !hbusreq5_p & c7658c;
assign v375e349 = hlock5 & v3744c08 | !hlock5 & v374f3ad;
assign v3772b81 = hmaster1_p & v3a635ea | !hmaster1_p & v377e355;
assign v376af1a = hmaster0_p & v3a6f765 | !hmaster0_p & !v3a6ebac;
assign v37520c4 = hgrant4_p & v374bd6a | !hgrant4_p & v375409b;
assign v373812a = jx3_p & v3a5f375 | !jx3_p & !v37500e2;
assign v376ff85 = hmaster2_p & v374734d | !hmaster2_p & v3747623;
assign v3741f4b = hbusreq0 & v3a63805 | !hbusreq0 & v373cc68;
assign v3a6f4b6 = hbusreq0_p & v3770993 | !hbusreq0_p & v3a670a1;
assign v3a6a8b4 = hmaster1_p & v3a635ea | !hmaster1_p & v375427c;
assign v3a5aa9d = hgrant2_p & v3748609 | !hgrant2_p & v3773b55;
assign v377df7d = hmaster2_p & v3755252 | !hmaster2_p & !v37541ff;
assign v3746a2b = hlock2 & v37548d8 | !hlock2 & v374868d;
assign v373fa73 = jx1_p & v3a66349 | !jx1_p & v373e11e;
assign v3a62cb5 = hmaster1_p & v3a6cc78 | !hmaster1_p & v8455ab;
assign v3745b32 = hlock0_p & v377ba55 | !hlock0_p & !v8455ab;
assign v3736a59 = hmaster1_p & v37302a2 | !hmaster1_p & v3a6cd87;
assign v3a5c3c4 = hmaster1_p & v3a70ac4 | !hmaster1_p & v8455ab;
assign v3724325 = hmaster0_p & v3776767 | !hmaster0_p & !v3770fa1;
assign v9ac541 = hbusreq7 & v372a06a | !hbusreq7 & v3726a2b;
assign v3a64c32 = hgrant7_p & v8455ab | !hgrant7_p & v3a629fb;
assign v375bed5 = hlock8_p & v375e961 | !hlock8_p & !v3a70f70;
assign v3763f8b = hbusreq1 & v39a5265 | !hbusreq1 & !v3733ea2;
assign v3757dee = hbusreq5_p & v37795d3 | !hbusreq5_p & v3777b00;
assign v3763c20 = hmaster1_p & v3a5e24e | !hmaster1_p & v3745315;
assign v373b0d2 = hbusreq4_p & v3747302 | !hbusreq4_p & v3733da4;
assign v37547c9 = hbusreq1 & v8455e7 | !hbusreq1 & v8455ab;
assign v377857d = hlock1 & v3770db8 | !hlock1 & v373b288;
assign v3758fc7 = hgrant2_p & v8455ba | !hgrant2_p & v3a6f67e;
assign v3a5f78a = hmaster2_p & v3a635ea | !hmaster2_p & v3a6162f;
assign v373ff58 = hgrant3_p & v377b6ce | !hgrant3_p & !v373e85a;
assign v3a6f470 = hbusreq8 & v375e8c1 | !hbusreq8 & v8455ab;
assign v372552c = hlock8 & v3a706c3 | !hlock8 & v3739e4f;
assign v374f3a3 = hgrant4_p & v3a6f32d | !hgrant4_p & v3a6aefd;
assign v377e493 = hmaster1_p & v37263bf | !hmaster1_p & v3a660e6;
assign v3738762 = hbusreq6_p & v377efd0 | !hbusreq6_p & v3778323;
assign v3a5beb8 = hmaster0_p & v3758cec | !hmaster0_p & v8455e7;
assign v3a70d85 = hgrant4_p & v380911c | !hgrant4_p & v376c4a9;
assign v3747897 = hbusreq8_p & v3a70d9b | !hbusreq8_p & v372fc7e;
assign v3757651 = hgrant2_p & v8455ab | !hgrant2_p & v3737ce6;
assign v3a6fc46 = hgrant6_p & v3734067 | !hgrant6_p & !v37551df;
assign v375ff95 = hlock1_p & v372e93d | !hlock1_p & v377c2ac;
assign v3742241 = hbusreq4_p & v37fca8d | !hbusreq4_p & v372cbdb;
assign v372fecd = hmaster0_p & v37424df | !hmaster0_p & v375449f;
assign v3a5408c = hlock6 & v376533e | !hlock6 & v3a6eead;
assign v3772098 = hmaster1_p & v3a71140 | !hmaster1_p & v372e749;
assign v3752d2c = hbusreq4_p & v376ac08 | !hbusreq4_p & v3a5a807;
assign v3a71186 = hmaster2_p & v3724270 | !hmaster2_p & v375f61e;
assign v374f1c3 = hgrant3_p & v37243d7 | !hgrant3_p & v3a6f2dd;
assign v3a6eece = hmaster0_p & v375e1b0 | !hmaster0_p & v3a59bbd;
assign v3a5918c = hmaster2_p & v3761719 | !hmaster2_p & v3773fc7;
assign v9181c9 = hbusreq3_p & v39a5381 | !hbusreq3_p & v3a63bbc;
assign adf1da = hbusreq4_p & v1e3771d | !hbusreq4_p & v3a7154f;
assign v3a6b102 = hbusreq4 & v3757575 | !hbusreq4 & v8455ab;
assign v373a291 = hlock4_p & v3a6f1e6 | !hlock4_p & v3a62550;
assign v3a537c5 = hgrant5_p & v8455ab | !hgrant5_p & v3a669dc;
assign v3a6f818 = hmaster2_p & v3a5b8b9 | !hmaster2_p & v3a6fcb0;
assign v375f61e = hbusreq4_p & v3725819 | !hbusreq4_p & v8455ab;
assign v37626ae = hlock8_p & v3744410 | !hlock8_p & v3a5b4a0;
assign v3a705d7 = hlock3_p & v372a958 | !hlock3_p & !v3a558c2;
assign v3731b88 = hlock0_p & v3770993 | !hlock0_p & v3a6f8dd;
assign v374d04b = hlock2_p & v3a6ebb0 | !hlock2_p & v3a6f9f6;
assign v374af22 = hbusreq0 & v3724715 | !hbusreq0 & v3a54811;
assign v3a6f1e6 = hgrant6_p & v3771b2c | !hgrant6_p & v3a575d6;
assign v3a6f954 = hbusreq5 & v3773a00 | !hbusreq5 & v3746e10;
assign v3733d5a = hbusreq3_p & v37684cf | !hbusreq3_p & v8455ab;
assign v3a6bc47 = hbusreq2 & v376c235 | !hbusreq2 & v8455ab;
assign v3a705ce = hgrant2_p & v8455b9 | !hgrant2_p & v3725f02;
assign v372ba40 = hmaster2_p & v374a1f5 | !hmaster2_p & v3a6fc5e;
assign v3746303 = hlock4_p & v375045d | !hlock4_p & v8455ab;
assign v3746487 = hbusreq5_p & v20d166d | !hbusreq5_p & v3750c50;
assign v3a6220e = hmaster0_p & v3a70117 | !hmaster0_p & v372c1fc;
assign v37676cd = hlock5_p & v37719a9 | !hlock5_p & !v3746ae3;
assign v3a6000d = hgrant6_p & v377f09a | !hgrant6_p & !v3a53c50;
assign v3737e04 = hlock6 & v3a640ab | !hlock6 & v3a70e10;
assign v372ff79 = hbusreq8_p & v3a709e8 | !hbusreq8_p & v376753a;
assign v374212e = hlock3 & v373184e | !hlock3 & v374f76a;
assign v3a6fd0c = hmaster0_p & v3751631 | !hmaster0_p & v35b71da;
assign v3a702e0 = hbusreq8 & v3a5d99f | !hbusreq8 & v3a5f218;
assign v3a68ad7 = hmaster1_p & v37419b4 | !hmaster1_p & v3a6a33a;
assign v3a70654 = hbusreq3_p & v372b74c | !hbusreq3_p & v3a6eb55;
assign v3770a68 = hmaster2_p & v374a6a5 | !hmaster2_p & v3a601a0;
assign v3a6f82c = hmaster2_p & v3a66110 | !hmaster2_p & v39a537f;
assign v37518fa = hbusreq3 & v3770af1 | !hbusreq3 & v377c6b3;
assign v3767be8 = hlock7 & v377e04e | !hlock7 & v374a60b;
assign v3a6972b = hbusreq3 & v3736028 | !hbusreq3 & v375b9c1;
assign v3a614cb = hlock6 & v3729f05 | !hlock6 & v37574d2;
assign v3740b8c = hbusreq7_p & v37240c0 | !hbusreq7_p & v373cba8;
assign v37606ba = hbusreq6 & v37672a5 | !hbusreq6 & v374acbe;
assign v375af57 = hbusreq0 & v37247f2 | !hbusreq0 & v8455ab;
assign v3a71327 = jx0_p & v3a6eaee | !jx0_p & v3742ecd;
assign v3a6f5c8 = hmaster2_p & v3a68838 | !hmaster2_p & v3776685;
assign v3a6be44 = hbusreq3_p & v3727215 | !hbusreq3_p & !v8455ab;
assign v37546c9 = hmaster1_p & v3a53e30 | !hmaster1_p & v23fde7b;
assign v37604e1 = hbusreq7_p & v375b22c | !hbusreq7_p & v375c652;
assign v3731d87 = hmaster0_p & v3a712c8 | !hmaster0_p & v372a696;
assign v376d4ee = hbusreq2 & v373502a | !hbusreq2 & v3a66051;
assign v3a5690d = hbusreq4_p & v376e033 | !hbusreq4_p & v33781d5;
assign v3773613 = hgrant8_p & v376abd1 | !hgrant8_p & v3769617;
assign v3a70261 = hlock4 & v377338f | !hlock4 & v3a6eb1e;
assign v377cef3 = hbusreq5 & v3726dfd | !hbusreq5 & !v37358ab;
assign v3775476 = stateA1_p & v8455ab | !stateA1_p & !v3a6ffe0;
assign v3a6fb0a = hlock8 & v374952b | !hlock8 & v3809ab5;
assign v3774f1e = hmaster1_p & v37316cb | !hmaster1_p & !v375d417;
assign v374bbcc = hbusreq0 & v3a59ba9 | !hbusreq0 & v8455ab;
assign v3a6fc97 = hbusreq7_p & v3a6f76d | !hbusreq7_p & v3a68871;
assign v3a545a7 = hmaster0_p & v37710c7 | !hmaster0_p & v3746f11;
assign v375bb3a = stateG10_1_p & v8455ab | !stateG10_1_p & !v8455eb;
assign v3a709d1 = hmaster0_p & v3744af9 | !hmaster0_p & !v372a696;
assign v376d4b7 = hgrant3_p & v8455be | !hgrant3_p & !v3728506;
assign v37445d7 = hbusreq4 & v3729a1c | !hbusreq4 & v373a341;
assign v3736b12 = hbusreq5_p & v3765cd5 | !hbusreq5_p & !v8455ab;
assign v3727c1d = hbusreq4 & v373f6ee | !hbusreq4 & v3a5a807;
assign v376a715 = hgrant6_p & v3a69487 | !hgrant6_p & v3729f6a;
assign v3773e52 = hmaster3_p & v374cd37 | !hmaster3_p & v8455ab;
assign v3a5cef4 = hbusreq2 & v372777c | !hbusreq2 & v377ba5a;
assign v3a708ad = hbusreq0 & v3765053 | !hbusreq0 & v8455ab;
assign v373e27e = hbusreq5_p & v377a13b | !hbusreq5_p & v377ef58;
assign v3a61ceb = hbusreq8_p & v3a5a323 | !hbusreq8_p & v3748494;
assign v3a5f6c2 = hmaster2_p & v3a6dc08 | !hmaster2_p & v3a6f993;
assign v3750c0d = hbusreq6 & v3a56e63 | !hbusreq6 & !v8455ab;
assign v37281e7 = hgrant6_p & v8455ca | !hgrant6_p & v375dc46;
assign v375bce7 = hmaster2_p & v3a63621 | !hmaster2_p & v3a641d5;
assign v3a5836e = hbusreq6_p & v3a651fc | !hbusreq6_p & v376bb26;
assign v3751e0a = hbusreq5_p & v3a619c0 | !hbusreq5_p & v3a66110;
assign v3a63bdb = hbusreq2 & v3767437 | !hbusreq2 & v8455b3;
assign v3755c8b = hgrant2_p & v3750269 | !hgrant2_p & v3770751;
assign v3a660a5 = hbusreq8_p & v373754d | !hbusreq8_p & v8455ab;
assign v373712d = hbusreq2 & v35b7808 | !hbusreq2 & v377eb9d;
assign v373a5b6 = hlock6 & v3a633a7 | !hlock6 & v377028b;
assign v3a695b7 = hmaster0_p & v3779060 | !hmaster0_p & v3749ec6;
assign v3a5d717 = hgrant3_p & v3a709c1 | !hgrant3_p & v3a71400;
assign v3723023 = hmaster2_p & v377989c | !hmaster2_p & v8455ab;
assign v3a6f31e = hbusreq7 & v3739493 | !hbusreq7 & v37775c7;
assign v3726077 = hgrant6_p & v3760ba8 | !hgrant6_p & v95d97e;
assign v3754b98 = hgrant6_p & v37697ba | !hgrant6_p & v3748353;
assign v3750883 = hmaster2_p & v8455ab | !hmaster2_p & v3778993;
assign v37406d2 = hlock0_p & v8455b0 | !hlock0_p & !v8455ab;
assign v372f475 = hbusreq6 & v3a711dd | !hbusreq6 & v3a708f0;
assign v1e378ce = jx0_p & v37592c9 | !jx0_p & v3a5b333;
assign v376489b = hbusreq0 & v374d80f | !hbusreq0 & v3749ec0;
assign v3a710f9 = hbusreq2_p & v3739b40 | !hbusreq2_p & v8455e7;
assign v376c635 = hgrant2_p & v3a6ceb7 | !hgrant2_p & !v377bc89;
assign v3773c40 = hbusreq7 & v3772aaf | !hbusreq7 & v37358f3;
assign v376804b = hlock6 & v375068a | !hlock6 & v3a6bf60;
assign v3a6f321 = hlock5_p & v3726339 | !hlock5_p & v3752a43;
assign v3a70eb7 = hgrant5_p & v37289bb | !hgrant5_p & v3768c2e;
assign v377fb81 = hmaster2_p & v3a70209 | !hmaster2_p & !v372ae9d;
assign v375d70e = hmaster2_p & v3a5f6d5 | !hmaster2_p & v3a62a08;
assign v3a70378 = hbusreq1 & v3a70459 | !hbusreq1 & v3a635ea;
assign v3732dc6 = locked_p & v3759ca5 | !locked_p & v8455ab;
assign v3a70f3d = hgrant6_p & v8455ab | !hgrant6_p & v3777a66;
assign v3a59649 = hmaster2_p & v37651c2 | !hmaster2_p & v3a5fc82;
assign v3a6d4c2 = hbusreq1 & v3749cea | !hbusreq1 & v3379037;
assign v3a70111 = jx2_p & v377e7f8 | !jx2_p & !v3a55352;
assign v37672aa = hgrant4_p & v8455ab | !hgrant4_p & v3a6fec9;
assign v3739896 = hbusreq4_p & v374d6dd | !hbusreq4_p & v8455b7;
assign v373af6f = hmaster0_p & v3a6ffca | !hmaster0_p & v3a572d0;
assign v375db64 = hbusreq5_p & v3a6fbec | !hbusreq5_p & v8455ab;
assign v37668e9 = hbusreq4_p & v377416d | !hbusreq4_p & v8455ab;
assign v376db98 = hbusreq7_p & v2092ff6 | !hbusreq7_p & v3a65587;
assign v3729991 = hlock2_p & v3a6e94b | !hlock2_p & v3750775;
assign v376e113 = hbusreq7_p & v3a6fdb1 | !hbusreq7_p & v8455ab;
assign v38094b8 = hlock5 & v3a7166f | !hlock5 & v37583f0;
assign v374aa90 = hbusreq4 & v3762388 | !hbusreq4 & v3809ec3;
assign v3a6e916 = hbusreq5 & v374fde8 | !hbusreq5 & !v3a65b39;
assign v3759aeb = hmaster2_p & v37297d0 | !hmaster2_p & v3770027;
assign v37775eb = hlock6 & v3759ca7 | !hlock6 & v37440a8;
assign v3a5cf28 = hgrant5_p & v8455ab | !hgrant5_p & !v373b887;
assign v3765615 = hbusreq7_p & v37697d0 | !hbusreq7_p & v375d2cf;
assign v3747b4c = hbusreq8_p & v3737808 | !hbusreq8_p & v374fa1e;
assign v3741401 = hgrant2_p & v37699a0 | !hgrant2_p & v3806b35;
assign v3a60130 = hgrant2_p & v3a70e21 | !hgrant2_p & v375964f;
assign v3776483 = hburst0_p & v8455ab | !hburst0_p & v3746c8d;
assign v3731e8c = hbusreq1_p & v372f5e7 | !hbusreq1_p & v3a5e8f6;
assign v3a6dc38 = hlock4 & v3a70e19 | !hlock4 & v372d336;
assign v3a68d49 = hbusreq0 & v3766b27 | !hbusreq0 & v3768a57;
assign v3774882 = hmaster2_p & v8455ab | !hmaster2_p & !v37356cc;
assign v3768de8 = hmaster0_p & v374729b | !hmaster0_p & !v3734967;
assign v3a701a5 = hbusreq0 & v372d8c9 | !hbusreq0 & v37331c0;
assign v3a5757f = hgrant2_p & v3a66671 | !hgrant2_p & v377a039;
assign v3a53fa4 = hbusreq6_p & v3775fb0 | !hbusreq6_p & v3a6f38c;
assign v3737223 = hbusreq6_p & v376dbdf | !hbusreq6_p & !v372fc81;
assign v376639f = hmaster2_p & v3a62caa | !hmaster2_p & v3a70410;
assign v3733b65 = locked_p & v3a5e24e | !locked_p & v3a61254;
assign v3a70e7d = hmaster2_p & v3a635ea | !hmaster2_p & v376aa76;
assign v3a6542a = hmaster0_p & v372984e | !hmaster0_p & v3a6f3cd;
assign v37711c8 = hbusreq2 & v3a54c77 | !hbusreq2 & v377ba55;
assign v375194a = hmaster1_p & v3734a4f | !hmaster1_p & v3a7055c;
assign v3a65a34 = hburst0 & v376c211 | !hburst0 & v3a555f9;
assign v376b7db = hgrant2_p & v3a6eead | !hgrant2_p & v37398eb;
assign v3734ca9 = hlock5 & v377de7f | !hlock5 & v3777b5f;
assign v3a621ea = hgrant6_p & v375b142 | !hgrant6_p & v372570c;
assign v360cfe2 = hbusreq3 & v3a59351 | !hbusreq3 & v8455ab;
assign v3a58604 = hmaster1_p & v375d387 | !hmaster1_p & v3a6fc4a;
assign v373cc82 = hbusreq5 & v3a6fdd1 | !hbusreq5 & v8455b3;
assign v3a64417 = hbusreq6_p & v373b10f | !hbusreq6_p & v374a84c;
assign v37585bf = hbusreq4_p & v37625a8 | !hbusreq4_p & !v2092faa;
assign v3a6fe50 = hlock5 & v3a71525 | !hlock5 & v37604fe;
assign v3730fab = hbusreq5 & cfaa3a | !hbusreq5 & v8455bf;
assign v35b7160 = hbusreq3_p & v3a5810a | !hbusreq3_p & v8455ab;
assign v372d30b = hmaster0_p & v3762e13 | !hmaster0_p & v3a6f54c;
assign v3a6607f = hmaster2_p & v37594c5 | !hmaster2_p & v3779eea;
assign v373cc51 = hgrant6_p & v91cdff | !hgrant6_p & v3743b79;
assign v3764ef1 = hmaster1_p & v37797c2 | !hmaster1_p & v373adb9;
assign v3a6f55d = hgrant5_p & v373bb2f | !hgrant5_p & v37710ad;
assign v37593a1 = hgrant4_p & v3746351 | !hgrant4_p & v3746683;
assign v3a6f4f5 = hmaster2_p & v377a801 | !hmaster2_p & v373a496;
assign v3a61ab0 = hmaster2_p & v3a70fd5 | !hmaster2_p & !v37367a0;
assign v376b18f = jx0_p & v3a63383 | !jx0_p & v3a70497;
assign v3a6b336 = hbusreq7 & v37685f1 | !hbusreq7 & v376ef20;
assign v372abf1 = hgrant6_p & v8455ab | !hgrant6_p & v372633a;
assign v3a71498 = hmaster2_p & v3a5ff46 | !hmaster2_p & v1e378b4;
assign v3a6e793 = hbusreq4 & v3754b2c | !hbusreq4 & v375da82;
assign v374fbcf = hbusreq2 & v372fc81 | !hbusreq2 & !v8455ab;
assign v375384f = hmaster0_p & v3a560b8 | !hmaster0_p & !v3a6cf7f;
assign v37484de = hbusreq1_p & v376b0fd | !hbusreq1_p & v8455ab;
assign v37606dc = hgrant4_p & v8455ab | !hgrant4_p & v3a6ef90;
assign v3a680e3 = hgrant6_p & v37604e9 | !hgrant6_p & v376a822;
assign v3806798 = hbusreq0 & v373b748 | !hbusreq0 & v3a70210;
assign v374b873 = hmaster1_p & v3a6f629 | !hmaster1_p & v3755502;
assign v3a6f621 = hbusreq5 & v3755c19 | !hbusreq5 & v373790d;
assign v373aecf = locked_p & v377a2e4 | !locked_p & !v8455ab;
assign v3a61cb0 = hmaster0_p & v3729b75 | !hmaster0_p & d4d3bb;
assign v374bec2 = hmaster1_p & v8455ab | !hmaster1_p & v3a675bb;
assign v3808db7 = jx1_p & v380a20c | !jx1_p & v3a5a2d0;
assign v3744577 = hburst0 & v2aca977 | !hburst0 & v375161a;
assign v3764881 = hbusreq4_p & v3a5b7c2 | !hbusreq4_p & v377a376;
assign v3747b81 = hmaster2_p & v374b8fa | !hmaster2_p & v3a68ef7;
assign v37747b4 = hgrant3_p & v374383b | !hgrant3_p & v8455ab;
assign v3a6b8cc = hmaster2_p & v376b0f2 | !hmaster2_p & v374c900;
assign v37591bc = hmaster0_p & v3a67447 | !hmaster0_p & v375355a;
assign v3a5524f = hmaster2_p & v375646d | !hmaster2_p & v8455ab;
assign v3a70a16 = hlock7 & v3755ae2 | !hlock7 & v375e9ca;
assign v3771667 = hbusreq6_p & v37404da | !hbusreq6_p & v3727db9;
assign v373a1a4 = hlock8_p & v3a57eae | !hlock8_p & !v3a59a60;
assign v37587fa = hmaster2_p & v3a7002c | !hmaster2_p & v3764dc0;
assign v3a66c20 = hgrant4_p & v3760ba3 | !hgrant4_p & v3a601a0;
assign v37258d0 = hmaster1_p & v8455ab | !hmaster1_p & v373d2e3;
assign v375d4de = hmaster2_p & v3a6162f | !hmaster2_p & v3a70891;
assign v3a5dbb7 = hbusreq1 & v3753dab | !hbusreq1 & v8455ab;
assign v375977c = hmaster0_p & v3725770 | !hmaster0_p & v3a6f53a;
assign v376c010 = jx1_p & v3a62f68 | !jx1_p & v3a5881c;
assign v3743c84 = hgrant5_p & v37359cf | !hgrant5_p & v3a7140b;
assign v3768b99 = hbusreq2_p & v3763f48 | !hbusreq2_p & v3a6600a;
assign v3a71555 = hgrant4_p & v8455ab | !hgrant4_p & v376ea99;
assign v96ab98 = hbusreq7_p & v3a712b5 | !hbusreq7_p & v3a6b4de;
assign v372658a = hmaster2_p & v8455bb | !hmaster2_p & v37522d3;
assign ca01e4 = hbusreq2_p & v373fbb4 | !hbusreq2_p & v8455ab;
assign v3a706eb = hbusreq5_p & v3a5936a | !hbusreq5_p & v3754981;
assign v3a6fa0a = hbusreq5_p & v374c679 | !hbusreq5_p & v372c85e;
assign v3739112 = hbusreq5_p & v375add1 | !hbusreq5_p & v376dd48;
assign v3a71054 = hbusreq4 & v3763fb5 | !hbusreq4 & v3a5b6de;
assign v3a53ed2 = hmaster0_p & v37386c6 | !hmaster0_p & v375c366;
assign v3a569a9 = hbusreq0 & v376cc23 | !hbusreq0 & v3a704a9;
assign v3775c0b = hbusreq4 & v377f73c | !hbusreq4 & v3a620d3;
assign v3a6f3d8 = hmaster2_p & v39a537f | !hmaster2_p & v3751734;
assign v373ff04 = hgrant4_p & v8455c2 | !hgrant4_p & v3752c73;
assign v37372c9 = hgrant2_p & v3a70a88 | !hgrant2_p & v3a6a393;
assign v23fe316 = hmaster0_p & v376d780 | !hmaster0_p & v3a6ff47;
assign v3a706b5 = hbusreq3_p & v372f747 | !hbusreq3_p & v374e418;
assign v3a6fd68 = hgrant6_p & v373c81c | !hgrant6_p & v372cede;
assign v3a632d8 = hgrant4_p & v3a70272 | !hgrant4_p & v3739dd4;
assign v3a54b2b = hmaster1_p & db1dc4 | !hmaster1_p & v3a5ad83;
assign v3a53f4c = hlock0_p & v20d166d | !hlock0_p & v3a66447;
assign v3a60618 = hlock2_p & v3a6cab1 | !hlock2_p & v37521af;
assign v3751f56 = hbusreq3 & v37566b2 | !hbusreq3 & v8455ab;
assign v3a5a8e6 = hmaster1_p & v3a5cff8 | !hmaster1_p & v37474e1;
assign v3751b9a = hbusreq5_p & v3a56a79 | !hbusreq5_p & v3a5dffe;
assign v3727eb2 = hbusreq0_p & v8455e7 | !hbusreq0_p & v374f307;
assign v3a58ca1 = hmaster2_p & v8455ab | !hmaster2_p & !v3757aa1;
assign v3a678d2 = hlock4_p & v3724a4b | !hlock4_p & adf78a;
assign v3a6333a = hbusreq5 & v375dd02 | !hbusreq5 & v3772200;
assign v3a70248 = hlock4_p & v3806db7 | !hlock4_p & v3a54c77;
assign v3a6eb0b = hlock3 & v3731afc | !hlock3 & d435c2;
assign v38072f4 = hbusreq2_p & v3a707cd | !hbusreq2_p & !v37521ed;
assign v37299de = hmaster2_p & v3740f5d | !hmaster2_p & v3a67fea;
assign v373c921 = hmaster1_p & v372cdde | !hmaster1_p & v3a5c860;
assign v3a55419 = hgrant4_p & v376d1bb | !hgrant4_p & v3728963;
assign v8ebe6e = hmaster0_p & v377bb3a | !hmaster0_p & v376d19f;
assign v3a6f51e = hmaster0_p & v3a57ccf | !hmaster0_p & v3726991;
assign v37289f0 = hgrant4_p & v8455c2 | !hgrant4_p & v3a67ff8;
assign v373cf73 = hbusreq7_p & v373dee0 | !hbusreq7_p & v3760a6e;
assign v3a58687 = hmaster0_p & v3771076 | !hmaster0_p & v3778d73;
assign v3a67965 = hmaster0_p & v374eab3 | !hmaster0_p & v376b540;
assign v3761b75 = hbusreq6_p & c6598e | !hbusreq6_p & v3a6fe06;
assign v3743e56 = hgrant0_p & v8455b0 | !hgrant0_p & v3a714c9;
assign v377b159 = hlock1_p & v3747c3e | !hlock1_p & v8455ab;
assign v3a704bd = hbusreq3_p & v377eaf2 | !hbusreq3_p & v3a7162d;
assign v373d27a = hbusreq0 & v376aad2 | !hbusreq0 & v372d967;
assign v3a5e5ec = hlock7_p & v3765b5a | !hlock7_p & v376e9e1;
assign v3743aee = hgrant1_p & v372a837 | !hgrant1_p & v8455ab;
assign v375427c = hlock5 & v1e3751e | !hlock5 & v3a6ae14;
assign v3733b77 = hbusreq0 & v3753526 | !hbusreq0 & v3a6eb0a;
assign v377052f = hbusreq3_p & v377eaf2 | !hbusreq3_p & v3738d63;
assign v3769c70 = hmaster2_p & v37482f8 | !hmaster2_p & v3a709e2;
assign v37437bb = hgrant5_p & v37626a9 | !hgrant5_p & v3771fea;
assign v3754ee0 = hmaster2_p & v3a635ea | !hmaster2_p & v376d1bb;
assign v3a562ea = hbusreq1 & v3a5600a | !hbusreq1 & v375444e;
assign v3a5f7d7 = hlock6 & v3740232 | !hlock6 & v3a5e881;
assign v37678fc = hlock0_p & v3379037 | !hlock0_p & !v8455ab;
assign v3772e90 = stateA1_p & v3762fc4 | !stateA1_p & !v3777ff3;
assign v376e033 = hbusreq4 & v376fd7a | !hbusreq4 & v3a63a66;
assign v3a709ce = jx1_p & v3723d16 | !jx1_p & v376f2f4;
assign v3a6d9c6 = stateG10_1_p & v35772a5 | !stateG10_1_p & !v3a635ea;
assign v3a6f5b3 = hbusreq5 & v3727fa7 | !hbusreq5 & v8455ab;
assign v374bf36 = hmaster2_p & v3759dda | !hmaster2_p & v3a713c9;
assign v37596d5 = hbusreq4 & v373e2c3 | !hbusreq4 & v8455e7;
assign v3a66998 = hbusreq8_p & v3747b78 | !hbusreq8_p & v3738b0f;
assign v3748609 = hbusreq2_p & v376f73c | !hbusreq2_p & v376ea4a;
assign v3a6afe8 = hlock6 & v3751e5e | !hlock6 & v376f501;
assign v37765fe = hbusreq3_p & v3a60132 | !hbusreq3_p & v8455ab;
assign v3a54455 = hlock4 & v375ad94 | !hlock4 & v3a5b7b9;
assign v3743745 = hbusreq1 & v3379037 | !hbusreq1 & v8455ab;
assign v3a712b1 = hgrant6_p & v3a5c0d4 | !hgrant6_p & !v8455ab;
assign v376ae9f = hmaster1_p & v8455ab | !hmaster1_p & v373790d;
assign v3a6f191 = hmaster1_p & v374a556 | !hmaster1_p & v3763bc4;
assign v37433e6 = hmaster2_p & v3754e5e | !hmaster2_p & v8455ab;
assign v3809f0e = hmaster0_p & v3761d7d | !hmaster0_p & !v377211f;
assign v3757e93 = hbusreq5 & v372713b | !hbusreq5 & v3806636;
assign v3769870 = hlock8 & v3a6fe07 | !hlock8 & v3741418;
assign v3a6546b = hmaster0_p & v3740aa7 | !hmaster0_p & v3747666;
assign v1e37cab = hbusreq6 & v374c163 | !hbusreq6 & v3a6da8a;
assign v373e5e7 = hgrant5_p & v8455ab | !hgrant5_p & da7312;
assign v3756a5f = hmaster0_p & v3741249 | !hmaster0_p & !v3a70da2;
assign v377ee7c = hmaster0_p & v2ff8e5c | !hmaster0_p & v3a6f90c;
assign v3733cd1 = hmaster2_p & v3a61bfd | !hmaster2_p & !v3744c10;
assign v38093c2 = hmaster0_p & v3750e23 | !hmaster0_p & v3a58d68;
assign v37364af = hmaster2_p & v8455b3 | !hmaster2_p & v37430e7;
assign v3732170 = hmastlock_p & v376f693 | !hmastlock_p & !v8455ab;
assign v3a6eaf7 = jx1_p & v37576ec | !jx1_p & v35b7768;
assign v375b943 = hbusreq6 & v3a701e4 | !hbusreq6 & !v8455ab;
assign v3a70794 = hbusreq3 & v3778765 | !hbusreq3 & v37447bf;
assign v374409a = hbusreq4_p & v37629cf | !hbusreq4_p & !v374e28f;
assign v373ff17 = hmaster0_p & v3751c1c | !hmaster0_p & v3a70476;
assign v3747ced = hbusreq8_p & v3737808 | !hbusreq8_p & v375fecf;
assign v37665f9 = hmaster1_p & v3a704bf | !hmaster1_p & v3a70499;
assign v374f1e9 = hbusreq5_p & v3774ae5 | !hbusreq5_p & !v3777825;
assign v37539fc = hgrant6_p & v3775234 | !hgrant6_p & v3a6ef49;
assign v37356b4 = hbusreq0 & v375ef49 | !hbusreq0 & v37346e8;
assign v3a5e8a0 = hgrant4_p & v3741609 | !hgrant4_p & !v3a7146f;
assign v2ff8d08 = hgrant4_p & v8455c9 | !hgrant4_p & v3985138;
assign v3a6ec29 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3724f05;
assign v37586d3 = hmaster0_p & v375d7fc | !hmaster0_p & v3a5bcf5;
assign v375ff5c = hlock2_p & v3a665dd | !hlock2_p & v3760f1e;
assign v3a70712 = hlock5 & v3a6f954 | !hlock5 & v3773a00;
assign v3a710a3 = hmaster0_p & v3764276 | !hmaster0_p & v3771be4;
assign v377c470 = hbusreq6 & v8455b0 | !hbusreq6 & v375d616;
assign v376e41a = hgrant0_p & v3a5c945 | !hgrant0_p & v3734c60;
assign v3a59a60 = hmaster1_p & v377439e | !hmaster1_p & v3a67e97;
assign v38099a1 = hbusreq4 & v3727b4a | !hbusreq4 & v3a635ea;
assign v3747797 = hmaster2_p & v374cab9 | !hmaster2_p & !v3751734;
assign v3764bd6 = hlock4 & v373b92c | !hlock4 & v3378e07;
assign v3769982 = hmaster0_p & v3a5d32a | !hmaster0_p & v3a5f992;
assign v375dd02 = hmaster0_p & v3730d1e | !hmaster0_p & !v3a6bbc6;
assign v3a71092 = hgrant6_p & v8455ab | !hgrant6_p & a2e8c8;
assign v37363da = hmaster0_p & v374d4e6 | !hmaster0_p & v3a6dded;
assign v374b7ea = hgrant5_p & v37429a7 | !hgrant5_p & v3738aa2;
assign v37325f4 = hgrant4_p & v377b6ce | !hgrant4_p & v3744e11;
assign v3a6d367 = hmaster2_p & v372aed1 | !hmaster2_p & v3a6ef2a;
assign v373556f = hgrant5_p & v3a6f253 | !hgrant5_p & !v8455ab;
assign v3a69ba1 = hmaster1_p & v37638fe | !hmaster1_p & v3a563c1;
assign v3809386 = hlock7_p & v3770c0d | !hlock7_p & !v8455ab;
assign v1e379fe = hlock0_p & v3a6ac26 | !hlock0_p & v8455ab;
assign v372abd8 = hlock0_p & v3722e5c | !hlock0_p & v372be9b;
assign v374554d = hbusreq5_p & d7e38d | !hbusreq5_p & v3766bdf;
assign v377d3e4 = hbusreq3 & v37359d8 | !hbusreq3 & v8455ab;
assign v3768b3d = hbusreq0 & v3778637 | !hbusreq0 & c7355c;
assign v3749a29 = hmaster3_p & v8455ab | !hmaster3_p & v3768d1d;
assign v3a6f7b3 = hmaster0_p & v3764684 | !hmaster0_p & v373c3a0;
assign v374bce5 = hbusreq7_p & v3a6b896 | !hbusreq7_p & v3a71546;
assign v3a6e7e1 = hbusreq1 & v373006f | !hbusreq1 & v8455ab;
assign v372e59e = hbusreq3 & v8455b0 | !hbusreq3 & v373cc68;
assign v374c58c = hbusreq0 & v374fd8a | !hbusreq0 & c7355c;
assign v9381f3 = hbusreq8_p & v3769712 | !hbusreq8_p & v3a6fc6d;
assign v3757663 = hbusreq3 & v3751734 | !hbusreq3 & !v8455ab;
assign v3772541 = hbusreq0 & v3760b17 | !hbusreq0 & v3a6ec56;
assign v3755fd4 = hmaster1_p & v376480b | !hmaster1_p & !v3a66a3a;
assign v374b912 = hlock5 & v3769cc4 | !hlock5 & v3a5b89a;
assign v3a70f43 = hgrant2_p & v8455ab | !hgrant2_p & v374283c;
assign v1e382c4 = hmaster2_p & v8455ab | !hmaster2_p & v37615d8;
assign v375e6ff = hmaster2_p & v3a67577 | !hmaster2_p & v8455ab;
assign v37352fa = hmaster3_p & v3a704c3 | !hmaster3_p & v37751c3;
assign v3756b48 = hbusreq2_p & v8455b7 | !hbusreq2_p & v374d479;
assign v3a6939d = hbusreq6 & v3a70f74 | !hbusreq6 & v375da10;
assign v37450cb = hbusreq0_p & v3a7151d | !hbusreq0_p & !v8455ab;
assign v3a7138a = hbusreq4 & v3a6af1d | !hbusreq4 & v3a5741c;
assign v3738f35 = hmaster0_p & v3779c38 | !hmaster0_p & v373594b;
assign v3a715ba = hmaster0_p & v3a6604e | !hmaster0_p & !v8455ab;
assign v3a70588 = hbusreq5_p & v377011b | !hbusreq5_p & v374e0a4;
assign v3a5e999 = hmaster2_p & v3a705f2 | !hmaster2_p & v3767b70;
assign v3a70876 = hlock0 & v374165f | !hlock0 & v3a571fd;
assign v37276a5 = hgrant2_p & v372f02f | !hgrant2_p & v3a703f1;
assign v3a6febd = hlock0_p & v3732e1b | !hlock0_p & v373cff4;
assign v3776225 = jx2_p & v376be82 | !jx2_p & v3a70762;
assign v373449d = hmaster0_p & v37507d6 | !hmaster0_p & v3a6f3b9;
assign v375e29c = hmaster3_p & v3752e80 | !hmaster3_p & v373ba93;
assign v375d8fb = hbusreq1_p & v3745b36 | !hbusreq1_p & v3a6eefe;
assign v3746f11 = hmaster2_p & v37710c7 | !hmaster2_p & v3775eee;
assign v3a6f106 = hlock5_p & v360d0c7 | !hlock5_p & !v8455ab;
assign v3a6897b = jx1_p & v35b7096 | !jx1_p & v377b0fb;
assign v373e28c = hmaster0_p & v3735ed2 | !hmaster0_p & v3a708e7;
assign v3a6294e = hmaster0_p & v3a6fa7a | !hmaster0_p & d5bac5;
assign v377bfb6 = hgrant2_p & v8455b9 | !hgrant2_p & v37690af;
assign v3a6f6c5 = hmaster2_p & v8455bd | !hmaster2_p & v3a6be44;
assign v372cec6 = hmaster2_p & v3a6c5ee | !hmaster2_p & v376bb26;
assign v372ab1b = hbusreq8 & v3737c1c | !hbusreq8 & v3762396;
assign v3a5a8c3 = hgrant2_p & v37721eb | !hgrant2_p & v8455ab;
assign v3738dca = hlock2_p & v8455e7 | !hlock2_p & !v8455ab;
assign v3a6da9c = hbusreq1_p & v2ff9190 | !hbusreq1_p & v8455ab;
assign v3735a77 = hbusreq8_p & v37284b7 | !hbusreq8_p & v37604e1;
assign v374ebac = hbusreq8_p & v376f62e | !hbusreq8_p & v3a70b2d;
assign v374abf3 = hbusreq0_p & v376d856 | !hbusreq0_p & !v3a5bf04;
assign v8c4a86 = hbusreq2_p & v376b141 | !hbusreq2_p & v8455bf;
assign v3a66750 = hbusreq2_p & v3a5ddee | !hbusreq2_p & v8455b0;
assign v373042a = hbusreq7_p & v3a691ea | !hbusreq7_p & v3752e82;
assign v3a6ab8d = hgrant3_p & v3a68aa8 | !hgrant3_p & v3740e49;
assign v375f123 = hbusreq7 & v3746f58 | !hbusreq7 & v372b870;
assign v375a16d = hlock4_p & v375d4e5 | !hlock4_p & v8455b0;
assign v3732968 = hbusreq0 & v23fdc13 | !hbusreq0 & v3a6464f;
assign v3749e4b = hbusreq5 & v1e37c22 | !hbusreq5 & v373de86;
assign v374eb89 = hbusreq6 & v372b304 | !hbusreq6 & v3379037;
assign v3728270 = hmaster0_p & v375fa7a | !hmaster0_p & v3a59905;
assign v372f151 = hgrant4_p & v8455c1 | !hgrant4_p & v372ed55;
assign v3778492 = hbusreq4 & v3776441 | !hbusreq4 & v8455e7;
assign v3a5be0b = hmaster0_p & v39ea76e | !hmaster0_p & v3724734;
assign v3768e0c = hbusreq4 & v3a63eaf | !hbusreq4 & v8455ab;
assign v3a56494 = hlock0 & v373bd6c | !hlock0 & v376ae41;
assign v376bcaa = hbusreq4_p & v3740171 | !hbusreq4_p & v37270d9;
assign v3a6f84a = hmaster2_p & v3a58d22 | !hmaster2_p & v374e542;
assign v37509f2 = hmaster0_p & v37237e8 | !hmaster0_p & v376ff85;
assign v3a60767 = hmaster0_p & v8455ab | !hmaster0_p & !v3a68f3d;
assign v374be73 = hmaster1_p & v8455ab | !hmaster1_p & v3734583;
assign v37685bf = hbusreq5_p & v3a71097 | !hbusreq5_p & v3809388;
assign v376c4ef = hbusreq5_p & v3774f56 | !hbusreq5_p & v375929c;
assign v3a5fde5 = hmaster2_p & v3765265 | !hmaster2_p & v3a70f1c;
assign v372b351 = hbusreq1_p & v374ed4b | !hbusreq1_p & v3724710;
assign v3a71524 = hlock6_p & v3a619c0 | !hlock6_p & !v8455ab;
assign v377bd9b = hlock5 & v377d4e1 | !hlock5 & v3762a76;
assign v3745510 = hlock5 & v375076a | !hlock5 & v3753a1d;
assign v3735bbc = hbusreq5_p & v373f940 | !hbusreq5_p & v3a6f012;
assign v3a7057f = hgrant2_p & v8455ab | !hgrant2_p & v3a67bff;
assign v3775341 = hbusreq0_p & v3a67dd0 | !hbusreq0_p & v3a59720;
assign v3778d9d = hbusreq4_p & v3a7033a | !hbusreq4_p & v37247f2;
assign v37397f0 = hgrant6_p & v3a70bd6 | !hgrant6_p & v3a705a5;
assign v3a56da3 = hbusreq4_p & v37761fe | !hbusreq4_p & v377e698;
assign v3a68f05 = hgrant8_p & v377f0e7 | !hgrant8_p & v3a5ba95;
assign v3a55a19 = hlock3_p & v372391f | !hlock3_p & v375e60f;
assign v3763ca5 = hbusreq8_p & v37730cd | !hbusreq8_p & v3777d70;
assign v37333de = hmaster0_p & d73f1d | !hmaster0_p & v3a63d22;
assign v3a6f7ef = hlock5_p & v3724e64 | !hlock5_p & v37296f5;
assign v3775120 = hbusreq8_p & v3a69427 | !hbusreq8_p & !v3758ab3;
assign v374d8ac = hbusreq4_p & v3a7033a | !hbusreq4_p & v8455ab;
assign v3757aa1 = hbusreq1_p & v375af00 | !hbusreq1_p & !v8455ab;
assign v3a70d29 = hlock8_p & v3a5e4e3 | !hlock8_p & v3767704;
assign v374e08e = hbusreq7_p & v3755d8e | !hbusreq7_p & v3a7087f;
assign v380887a = hlock1 & v357732f | !hlock1 & v3a70a12;
assign v375b97a = hmaster0_p & v3725932 | !hmaster0_p & v375c621;
assign v373409f = hbusreq4 & v374362e | !hbusreq4 & !v35b710e;
assign v3a6f891 = hmaster1_p & v3a696a7 | !hmaster1_p & bde868;
assign v372eb00 = hmaster2_p & v377329c | !hmaster2_p & !v8455ab;
assign v374c01f = hlock0_p & v37665bf | !hlock0_p & v3a6a939;
assign v3775a29 = hgrant4_p & v8455ab | !hgrant4_p & !v3a57c0b;
assign v3a6f467 = hlock5 & v3a6ae23 | !hlock5 & v3a6b768;
assign v3a6e02d = hbusreq6 & v37429b9 | !hbusreq6 & v377728d;
assign v376d85d = hmaster1_p & v8455bb | !hmaster1_p & v3743e7b;
assign v3a61964 = hlock8 & v373e4ca | !hlock8 & v37355e3;
assign v3769f61 = hbusreq4_p & v3779060 | !hbusreq4_p & !v3a6dfb2;
assign v3a53dff = hgrant3_p & v8455ab | !hgrant3_p & v3a65245;
assign v372298c = hbusreq4_p & v3749cdf | !hbusreq4_p & v37274ef;
assign v376480c = hlock4 & v3a6dd7e | !hlock4 & v3a5b8e4;
assign v373a0ea = hmaster2_p & v8455ab | !hmaster2_p & !v39a5265;
assign v3a71512 = hbusreq7 & v3a6f5aa | !hbusreq7 & v3733b90;
assign v3733e9e = locked_p & v8455ab | !locked_p & v1e38224;
assign v3a71156 = hgrant7_p & v377997c | !hgrant7_p & v3a71241;
assign v3577344 = hbusreq7 & v37665c9 | !hbusreq7 & v376c07e;
assign v3750dd3 = hlock2_p & v373aaa8 | !hlock2_p & !v8455ab;
assign v376e4bd = hgrant6_p & v372f02f | !hgrant6_p & v37276a5;
assign v37577db = hbusreq6 & v377d41d | !hbusreq6 & v375cf36;
assign v3774075 = hbusreq0 & v39a52e6 | !hbusreq0 & v372ee41;
assign v3745eb8 = hlock5 & v3749840 | !hlock5 & v376747e;
assign v3771da0 = hmaster3_p & v3a56dff | !hmaster3_p & v3726994;
assign v373bf74 = hmaster2_p & v372b6db | !hmaster2_p & !v8455ab;
assign v377ed4b = hmaster1_p & v3a5459f | !hmaster1_p & !v376ca02;
assign v3777243 = hmaster3_p & v3775e46 | !hmaster3_p & v3a69091;
assign v377265b = hmaster1_p & v3a6ff8c | !hmaster1_p & v376256f;
assign v377653f = hmaster0_p & v377429c | !hmaster0_p & v3a6e872;
assign v37661db = hbusreq0 & v372bdd9 | !hbusreq0 & v377349f;
assign v373b18b = hmaster2_p & v3a6fd81 | !hmaster2_p & v3a5f40e;
assign v3a70d5c = hmaster3_p & v8455ab | !hmaster3_p & v376c3f8;
assign v3a70ffb = hbusreq2_p & v375ff5c | !hbusreq2_p & v8455ab;
assign v3752845 = hmaster0_p & v3738336 | !hmaster0_p & v8455ab;
assign v3a6f5ae = hlock5 & v3a5cb0e | !hlock5 & v37680a7;
assign v374ebd1 = hgrant2_p & v3a6ae68 | !hgrant2_p & v3772e0a;
assign v3740c73 = hbusreq7 & v3a6eb97 | !hbusreq7 & v3776859;
assign v37672af = hgrant4_p & v3729031 | !hgrant4_p & v8455ab;
assign v3a5a573 = hbusreq4 & v3754f6b | !hbusreq4 & v8455ab;
assign v3728526 = hbusreq6_p & v3769f88 | !hbusreq6_p & v376b1bf;
assign v3a6c6ac = hbusreq5 & v373f88a | !hbusreq5 & v8455ab;
assign v375a250 = hgrant0_p & v376dfed | !hgrant0_p & v376bf8d;
assign v3a6f00d = hmaster1_p & v380a170 | !hmaster1_p & v3777527;
assign v3776fec = hbusreq8 & v8455ab | !hbusreq8 & v3765e47;
assign v3a7119e = hgrant3_p & v37579a9 | !hgrant3_p & v377320c;
assign v3756091 = hmaster1_p & v3733bfc | !hmaster1_p & v3740c13;
assign v375af0b = hbusreq5_p & v3760bfa | !hbusreq5_p & v3a71072;
assign v375d3e2 = hmaster1_p & v8455ab | !hmaster1_p & v3766c68;
assign v3a6a129 = hlock4_p & v373a841 | !hlock4_p & v8455e7;
assign v374bcfb = hbusreq6 & v3723493 | !hbusreq6 & v8455ab;
assign v3a6fa10 = hbusreq8_p & v3a635ea | !hbusreq8_p & v2092f2c;
assign v3733334 = hgrant2_p & v8455ab | !hgrant2_p & v3378a03;
assign v3a5bf75 = hmaster2_p & v3775303 | !hmaster2_p & v3a6c23b;
assign v3737456 = hgrant5_p & v8455c6 | !hgrant5_p & v3a5f894;
assign v3a7000f = hmaster2_p & v3a70bf4 | !hmaster2_p & v376f903;
assign v37582e1 = hmaster0_p & v37640e9 | !hmaster0_p & v373d55f;
assign v3a6a95a = hbusreq7 & v37351f6 | !hbusreq7 & !v8455ab;
assign v3763716 = hbusreq5_p & v374c9c2 | !hbusreq5_p & v376ee82;
assign v376bade = hbusreq1_p & v3a635ea | !hbusreq1_p & v373b288;
assign v3a6f6f8 = hbusreq8_p & v376ae9f | !hbusreq8_p & v373b241;
assign v3a63daa = hmaster1_p & v35b7168 | !hmaster1_p & v3760c3d;
assign v3a60125 = hgrant5_p & v376dfc9 | !hgrant5_p & v3a64fee;
assign v375e373 = stateA1_p & v3a5ff81 | !stateA1_p & v3a5cf0b;
assign v3808ed4 = hbusreq2_p & v3744983 | !hbusreq2_p & v3740fef;
assign v3757254 = hbusreq6 & v3a61d2e | !hbusreq6 & v3a6efea;
assign v37771ed = hmaster2_p & v372424e | !hmaster2_p & v8455ab;
assign v3747ad6 = hlock0 & v375b9c1 | !hlock0 & v376fc77;
assign v37597fa = hlock7 & v37591f2 | !hlock7 & v375a543;
assign v8639e9 = hgrant4_p & v8455ab | !hgrant4_p & v3742af4;
assign v3a700d4 = hmaster1_p & v39a4df7 | !hmaster1_p & v8455bd;
assign v3741c39 = hbusreq8 & v3774757 | !hbusreq8 & v3742476;
assign v3a6ad1f = hbusreq4_p & v37536c3 | !hbusreq4_p & v3a705ef;
assign v3a69409 = hmaster1_p & v3a62a25 | !hmaster1_p & v376046c;
assign v3a55033 = hbusreq2_p & v376d256 | !hbusreq2_p & !v8455ab;
assign v3a54560 = hbusreq0 & v37474dc | !hbusreq0 & v3a5987a;
assign v373e587 = hlock5 & v3a6fb06 | !hlock5 & v3a6eece;
assign v3a70e7b = hbusreq4_p & v375524f | !hbusreq4_p & !v8455ab;
assign v3a6d219 = hbusreq2_p & v3732588 | !hbusreq2_p & v8455ab;
assign v3a70c28 = hbusreq5_p & v3768c08 | !hbusreq5_p & v3768dd8;
assign v3769696 = hmaster2_p & v3a635ea | !hmaster2_p & v377bfc0;
assign v3a55ee6 = hbusreq0 & v37307dd | !hbusreq0 & !v8455ab;
assign v3a702c6 = hgrant3_p & v3a5a510 | !hgrant3_p & v3a71270;
assign v3a66373 = hgrant5_p & v373f260 | !hgrant5_p & v3a5dd10;
assign v37503c2 = hmaster0_p & v3759031 | !hmaster0_p & v3a5ce54;
assign v37259e6 = hgrant6_p & v3a6b873 | !hgrant6_p & v372e4b3;
assign bf3e2b = hgrant3_p & v8455ab | !hgrant3_p & v3749b84;
assign v3a64f54 = hmaster1_p & v373899b | !hmaster1_p & v3765c1f;
assign v3752f9b = hmaster0_p & v3a6de93 | !hmaster0_p & v374e51a;
assign v372e3ea = hbusreq4_p & v3809194 | !hbusreq4_p & v373031f;
assign v374aa67 = hbusreq7 & v3727195 | !hbusreq7 & v3736003;
assign v3771dd8 = hmaster3_p & v3a6f9bf | !hmaster3_p & v372d49e;
assign v377a356 = hgrant4_p & v3769630 | !hgrant4_p & v375e6ed;
assign v3756031 = hbusreq5 & v3a700e9 | !hbusreq5 & v3a64624;
assign v3a7017e = hmaster2_p & v377a865 | !hmaster2_p & v8455ab;
assign v376f1d0 = hmaster1_p & v8455ab | !hmaster1_p & v3769753;
assign v879494 = hmaster0_p & v8455ab | !hmaster0_p & !v3740bcb;
assign v3731b11 = hbusreq3_p & v3a5d356 | !hbusreq3_p & v374e03d;
assign v3a68f5f = hbusreq5_p & v373d27f | !hbusreq5_p & v3734062;
assign v372f2b7 = hbusreq0 & v3a7062e | !hbusreq0 & v375bcf2;
assign v372493b = hlock0_p & v376f73c | !hlock0_p & v377d74d;
assign v3a5c2f5 = hbusreq7 & v3758c5e | !hbusreq7 & v37437bb;
assign v377da41 = hmaster1_p & v3a566eb | !hmaster1_p & v37555b4;
assign v3a29814 = hbusreq5_p & v3a6fe4a | !hbusreq5_p & v8455ab;
assign v3a59656 = jx3_p & v3a53962 | !jx3_p & v375c6cc;
assign v37250a3 = hlock3 & v376be2c | !hlock3 & v372c134;
assign v374b4da = hgrant2_p & v3a5718e | !hgrant2_p & v8455ab;
assign v374803b = hbusreq7_p & v3a5a4c0 | !hbusreq7_p & v3a56929;
assign v373e0b1 = hmaster1_p & v375eefe | !hmaster1_p & v376ad8c;
assign v3a70e38 = hmaster1_p & v3729d0b | !hmaster1_p & !v375c0f1;
assign v3763b5d = hmaster2_p & v3a70374 | !hmaster2_p & v3764a2d;
assign v3723809 = hbusreq8_p & v3765615 | !hbusreq8_p & v3a70d41;
assign v37697fc = hbusreq2_p & v376f56d | !hbusreq2_p & v3a6ef62;
assign v3a5cebb = hbusreq0 & v3a6fc17 | !hbusreq0 & !v3765b09;
assign v3a6f9a1 = hmaster0_p & v3742698 | !hmaster0_p & !v2092ec6;
assign v37370b9 = hgrant2_p & v37234e0 | !hgrant2_p & !a6f1de;
assign v37230ec = hmaster2_p & v377e419 | !hmaster2_p & v3730b6c;
assign v3735486 = hmaster2_p & v3a7142f | !hmaster2_p & v3744df8;
assign v3746a87 = hmaster2_p & v3769740 | !hmaster2_p & v37289f0;
assign v376c2b7 = hgrant4_p & v3a5bffe | !hgrant4_p & !v3a71170;
assign v375d690 = hlock0_p & v3759032 | !hlock0_p & !v39a537f;
assign v37654b9 = hgrant6_p & v8455ca | !hgrant6_p & v37252d0;
assign v3748851 = hready_p & v3773bd7 | !hready_p & v374743a;
assign v3a58017 = hmaster0_p & v3746b7f | !hmaster0_p & v3764683;
assign v374e61c = hbusreq8_p & v3737bd8 | !hbusreq8_p & v3723fa6;
assign v3764219 = hmaster0_p & v377038e | !hmaster0_p & v3767121;
assign v3a706df = hbusreq0_p & v37496fa | !hbusreq0_p & v3743b9e;
assign v3a5fa45 = hbusreq7 & v372b57a | !hbusreq7 & v3a6e721;
assign v3776faf = hgrant6_p & v3a6f3aa | !hgrant6_p & v3743338;
assign v2acaf72 = hbusreq6_p & v3a70cd1 | !hbusreq6_p & !v3a65562;
assign v3762ffa = hmaster2_p & v8455ab | !hmaster2_p & v3a5f371;
assign v3a66bdb = hburst0 & v373d9e5 | !hburst0 & v8455ab;
assign v3723d79 = hmaster1_p & v3a635ea | !hmaster1_p & v3a7129c;
assign v377e431 = hgrant5_p & v3a6fa8b | !hgrant5_p & v373b08f;
assign v3a564a8 = hbusreq2 & v3a6c60e | !hbusreq2 & v3773ee6;
assign v375f317 = hgrant2_p & v8455ab | !hgrant2_p & v3806ec2;
assign v3a6cf44 = hgrant5_p & ca32a1 | !hgrant5_p & v3a64b87;
assign v37385d3 = hmaster1_p & v37773d6 | !hmaster1_p & v37705ec;
assign v3a573bb = hmaster1_p & v3745bee | !hmaster1_p & v376b2f4;
assign v3733cf4 = hgrant5_p & v8455ab | !hgrant5_p & !v377d1dc;
assign v3a59517 = hgrant2_p & v373a25b | !hgrant2_p & v377add5;
assign v3729d65 = hbusreq6_p & v2aca977 | !hbusreq6_p & v3a6fd79;
assign v3a6fdf5 = hmaster1_p & v3725380 | !hmaster1_p & v374b074;
assign v33789f3 = hlock8_p & v8455ab | !hlock8_p & v3a6f681;
assign v372be16 = hgrant4_p & v8455ab | !hgrant4_p & v3a5b903;
assign v3759cb9 = hbusreq5_p & v37507dc | !hbusreq5_p & v3a6f5a2;
assign v3727703 = hbusreq2 & v3a6ad59 | !hbusreq2 & v3a6a82a;
assign v3770754 = hgrant4_p & v35b724a | !hgrant4_p & v8455ab;
assign v3a6affa = stateG2_p & v3a5a496 | !stateG2_p & v8455ab;
assign v3809da1 = hlock3_p & v20d166d | !hlock3_p & v8455ab;
assign v3745b9c = hmaster2_p & v374ad16 | !hmaster2_p & v37436bc;
assign v3a64b55 = hmaster1_p & v337905c | !hmaster1_p & v3723e23;
assign v377f548 = hgrant4_p & v3a708f2 | !hgrant4_p & v3a6fc7a;
assign v3756234 = hbusreq8_p & v373f497 | !hbusreq8_p & v375e3fd;
assign v3a5ab84 = hgrant6_p & v3a605b5 | !hgrant6_p & v3a558c5;
assign v37300ba = hmaster0_p & v3a637dc | !hmaster0_p & v3730601;
assign v3a57486 = hbusreq5 & v2092a68 | !hbusreq5 & v3744abe;
assign v377843d = hmaster0_p & v37617dd | !hmaster0_p & v3757966;
assign v3773506 = hbusreq4_p & v375b2e2 | !hbusreq4_p & v377bf71;
assign v3a53f42 = hbusreq4 & v376a056 | !hbusreq4 & v3a5a807;
assign v3a6d096 = hbusreq4_p & v374bf59 | !hbusreq4_p & v3a58db9;
assign v3747afb = hmaster2_p & v373a27c | !hmaster2_p & v3740171;
assign v3730dc4 = hbusreq0 & v8455b0 | !hbusreq0 & v3755791;
assign v377d8b7 = hbusreq6_p & v375c06a | !hbusreq6_p & !v8455ab;
assign v3737571 = hbusreq6_p & v3a60f22 | !hbusreq6_p & v3806f24;
assign v3732515 = hgrant6_p & v3728d84 | !hgrant6_p & v3a69ada;
assign v37639b1 = hbusreq0 & v3a714fc | !hbusreq0 & v3a5b1a3;
assign v3759020 = start_p & v37688a5 | !start_p & v8455ab;
assign v37355ce = hbusreq4 & v3a6c1ec | !hbusreq4 & v38072fd;
assign v1e37d14 = hbusreq5_p & v3725804 | !hbusreq5_p & !v8455ab;
assign v3730a22 = hlock8_p & v8455ab | !hlock8_p & v374e3c1;
assign v376a454 = hmaster1_p & v8455ab | !hmaster1_p & v373e48c;
assign v374c576 = hlock7 & v3a6130e | !hlock7 & v3a6fd76;
assign v375a28e = hmaster2_p & v372e711 | !hmaster2_p & v37716ca;
assign ab638b = hlock3_p & v8455ab | !hlock3_p & v8455e7;
assign v3a60b90 = hmaster2_p & v375c791 | !hmaster2_p & a96343;
assign v37271e7 = hbusreq4_p & v3a708a2 | !hbusreq4_p & v8455b0;
assign v375efc9 = hbusreq2 & v3a64703 | !hbusreq2 & v37275ef;
assign v3a5e7fd = hlock1 & v374197c | !hlock1 & v37521ff;
assign v3a70616 = hmaster0_p & v3a5d6aa | !hmaster0_p & v3a65752;
assign v3a6e0f4 = hbusreq0 & v39a52e6 | !hbusreq0 & v3a6f746;
assign v2acae79 = hmaster1_p & v3a6deea | !hmaster1_p & v373fb22;
assign v2092eb7 = hgrant4_p & v377b6ce | !hgrant4_p & v37229b8;
assign v3773336 = hbusreq5_p & v3a6fbbd | !hbusreq5_p & !v360d0c7;
assign v376226e = hbusreq5 & v376e115 | !hbusreq5 & v373755a;
assign v3761f39 = hgrant3_p & v3759512 | !hgrant3_p & !v3751364;
assign v373f9ad = hlock0 & v38072fd | !hlock0 & v3763186;
assign v373402f = hgrant5_p & v375478f | !hgrant5_p & v3a70d3d;
assign v37485ce = hbusreq0 & v3a6d03c | !hbusreq0 & v3726979;
assign v3a58fe2 = hmaster0_p & v37434c6 | !hmaster0_p & v8455b3;
assign v3727293 = hbusreq3_p & v3731e0f | !hbusreq3_p & v8455ab;
assign v374d5c0 = hlock6_p & v3740df7 | !hlock6_p & v3757aa1;
assign v3768ef1 = hlock2 & v372eae4 | !hlock2 & v3a55b2d;
assign v3a70bc8 = hlock6_p & v8455ab | !hlock6_p & v3771ce2;
assign v376ffbf = hlock4 & v3a62197 | !hlock4 & v375b349;
assign v373b6e9 = hbusreq8 & v3a698b7 | !hbusreq8 & v8455ab;
assign v37757e0 = hready & v3726dfa | !hready & !v373dceb;
assign v3768c2a = hlock6_p & v37407f5 | !hlock6_p & v3a6f4dc;
assign v3a61519 = hmaster1_p & v3754a54 | !hmaster1_p & v375e120;
assign v3a71540 = hgrant6_p & v8455ab | !hgrant6_p & v3a571b6;
assign v376d4d9 = hbusreq8 & v375cfd9 | !hbusreq8 & v373a8a1;
assign v375e94c = hlock5_p & v3a70d43 | !hlock5_p & v8455cb;
assign v3a560d9 = hbusreq8 & v3733b9a | !hbusreq8 & v373adea;
assign v3a6bbed = hgrant3_p & v8455ab | !hgrant3_p & v37470d6;
assign d0b9d7 = hgrant3_p & v8455e7 | !hgrant3_p & v37598c6;
assign v373e88f = hmaster1_p & v37430c6 | !hmaster1_p & v3a70c12;
assign v23fe0bb = hbusreq1_p & v37416b5 | !hbusreq1_p & v3743b9e;
assign v372294a = hmaster0_p & v3a6ff5b | !hmaster0_p & v375afe9;
assign v373bdd9 = hmaster1_p & v3761915 | !hmaster1_p & v3a70052;
assign v374c9d9 = hbusreq7 & v3a5c5e1 | !hbusreq7 & v3737808;
assign v3a70f3e = hlock2_p & v3a715e2 | !hlock2_p & v8455b7;
assign v3732086 = hlock0 & v3749bf0 | !hlock0 & v37544cb;
assign v373e09c = hgrant2_p & v3757c37 | !hgrant2_p & v380749d;
assign v37283ff = hbusreq0 & v37291ce | !hbusreq0 & !v3a6fa37;
assign v3a60e7e = hbusreq6_p & v3a60cbd | !hbusreq6_p & v8455ab;
assign v372ca2a = hlock4_p & v3a660f2 | !hlock4_p & v35772c9;
assign v3a70fc4 = hmaster0_p & ab0224 | !hmaster0_p & v37614c1;
assign v3a6b73b = hmaster0_p & v3a5473a | !hmaster0_p & v3747971;
assign v3a6f396 = hmaster1_p & v8cd321 | !hmaster1_p & v3745b39;
assign v3750f72 = hgrant2_p & v3a635ea | !hgrant2_p & v3a5a29e;
assign v3a70222 = hmaster2_p & v377bb3a | !hmaster2_p & v372d203;
assign v3763183 = hmaster0_p & v3a6f9cd | !hmaster0_p & !v3746ce0;
assign v372ad2c = hmaster1_p & v3a5c3d6 | !hmaster1_p & v39ebb8a;
assign v37374a1 = hmaster2_p & v8455ab | !hmaster2_p & v8455bb;
assign v3761178 = hmaster2_p & v375f94a | !hmaster2_p & v3747d68;
assign v376f73c = hbusreq1_p & v3a5891c | !hbusreq1_p & v376ef42;
assign v37635ab = hmaster2_p & v3a70a5c | !hmaster2_p & v373de4b;
assign v377d545 = hbusreq5 & v3a6f0f5 | !hbusreq5 & v372a744;
assign v3765395 = hbusreq7_p & v372ea2d | !hbusreq7_p & v3a6e0ab;
assign v375c806 = hgrant0_p & v37773a9 | !hgrant0_p & v377c3fb;
assign v374037a = hlock0_p & v3a70e52 | !hlock0_p & v37531ff;
assign v3768130 = hgrant2_p & v8455ab | !hgrant2_p & v375a6e6;
assign v3752684 = hmaster2_p & v3772b00 | !hmaster2_p & v3759506;
assign v3755e97 = hbusreq0 & v3745f8d | !hbusreq0 & v8455ab;
assign v380909f = hlock7 & v376f536 | !hlock7 & v374a0ab;
assign v3758ab3 = hmaster1_p & v377adf5 | !hmaster1_p & v374b879;
assign v3723bf9 = hbusreq8_p & v374a510 | !hbusreq8_p & v3771ea2;
assign v3a627b3 = hlock4 & v376d2dc | !hlock4 & v3762a2a;
assign v373c1ff = hmaster0_p & v377e27e | !hmaster0_p & v375f2f2;
assign v3756ef4 = hmaster2_p & v373891b | !hmaster2_p & v375bf93;
assign v38097c4 = hbusreq7_p & v377ce96 | !hbusreq7_p & v3a6fb7b;
assign v3a5a36d = hbusreq6 & v3a6113b | !hbusreq6 & v8455ab;
assign v37434b2 = hmaster2_p & v3a5e817 | !hmaster2_p & !v3a55cd6;
assign v3a70406 = jx0_p & v37739a8 | !jx0_p & v3760167;
assign v37415c3 = hbusreq5_p & v37497ce | !hbusreq5_p & !v376a4ba;
assign v376e7f5 = hmaster2_p & v376a31b | !hmaster2_p & v3762870;
assign v3a575d5 = hgrant5_p & v8455ab | !hgrant5_p & v376cdc4;
assign v3760e75 = hbusreq6_p & v37329e1 | !hbusreq6_p & !v8455ab;
assign v3a58f20 = hlock4_p & v374caab | !hlock4_p & v373399e;
assign v372f071 = hbusreq6 & v3a70131 | !hbusreq6 & !v8455ab;
assign v3741bd4 = jx0_p & v3724bdd | !jx0_p & v3760ca3;
assign v3737c39 = jx0_p & v3a700ff | !jx0_p & v373ff40;
assign v375f77f = hmaster0_p & v3a5a6e6 | !hmaster0_p & v372421d;
assign v3727347 = hbusreq4 & v37784cc | !hbusreq4 & v8455ab;
assign v373b687 = hbusreq2_p & v3747302 | !hbusreq2_p & v3a70b92;
assign v373228a = hbusreq6_p & v377c3ea | !hbusreq6_p & v375f326;
assign v376a8c8 = hmaster1_p & v3a715bb | !hmaster1_p & v3731123;
assign v3a6f27d = hbusreq4_p & v3a635ea | !hbusreq4_p & v377c6b3;
assign v373ff99 = locked_p & v3a617fa | !locked_p & !v8455ab;
assign v373b7dd = hbusreq5_p & v3a65402 | !hbusreq5_p & !v372bb0f;
assign v377b92f = hgrant4_p & v3a53eeb | !hgrant4_p & v3a56d78;
assign v377c7b2 = hbusreq2 & v374b3cf | !hbusreq2 & v8455b3;
assign v37675f4 = hgrant3_p & v3759842 | !hgrant3_p & v376f148;
assign v3756683 = hbusreq5 & v3a6fc35 | !hbusreq5 & v8455ab;
assign v3a703ba = hbusreq7 & v372588c | !hbusreq7 & cb8cbb;
assign v3a646fb = hbusreq2_p & v373081f | !hbusreq2_p & v3a63621;
assign v3774618 = hgrant7_p & v8455ab | !hgrant7_p & v23fdea8;
assign v3738aa2 = hmaster1_p & v3770538 | !hmaster1_p & v3a6db03;
assign v3a6202c = hbusreq8_p & v377a522 | !hbusreq8_p & d5e2c2;
assign v3768873 = hmaster2_p & v3a70cc3 | !hmaster2_p & v3a67967;
assign v376c351 = hgrant2_p & v372fd12 | !hgrant2_p & v37406a7;
assign v3a6ebd2 = hmaster0_p & v377e5ac | !hmaster0_p & v372c1fc;
assign v3a553bc = hmaster1_p & v377e156 | !hmaster1_p & v374e8a2;
assign v373142a = hbusreq6 & v37348ee | !hbusreq6 & v3a69487;
assign v3767dd2 = hlock7_p & v375a475 | !hlock7_p & v377c487;
assign v3751a94 = hbusreq5_p & v37278f5 | !hbusreq5_p & v376c652;
assign v372e821 = hbusreq0 & v372539e | !hbusreq0 & v3a700b6;
assign v374a7c3 = hgrant7_p & v373d81e | !hgrant7_p & v372e775;
assign v3722f12 = hgrant0_p & v37773a9 | !hgrant0_p & v3a6f40c;
assign v374f138 = hbusreq4_p & v3a70f9f | !hbusreq4_p & !v8455ab;
assign v3747800 = hbusreq4_p & v376acee | !hbusreq4_p & v3a6c7ef;
assign v374d6f6 = hmaster1_p & v375329c | !hmaster1_p & v375523e;
assign v37676a5 = hbusreq7_p & v374b2c2 | !hbusreq7_p & v3734810;
assign v3a60723 = hbusreq4_p & v3a7165d | !hbusreq4_p & v3a6ff26;
assign v37625d5 = jx0_p & v37261a6 | !jx0_p & v3a6731d;
assign v3a6fa30 = hbusreq3_p & v37720d8 | !hbusreq3_p & v3a5cd20;
assign v37462ee = hmaster2_p & v3a6fdd1 | !hmaster2_p & v3a6f240;
assign v3a6fafe = hmaster2_p & v3a70d99 | !hmaster2_p & v37369b2;
assign v3765222 = hmaster1_p & v377d1dc | !hmaster1_p & v3723923;
assign ce7a16 = hbusreq7_p & v3727cec | !hbusreq7_p & v37419fa;
assign v3758a11 = hmaster3_p & v37390ca | !hmaster3_p & v372ab45;
assign v3a702fe = hlock2 & v37379d7 | !hlock2 & v372600f;
assign v3a63cce = hmaster1_p & v372faf3 | !hmaster1_p & v377cb0b;
assign v3766645 = hbusreq7 & v3745dae | !hbusreq7 & v3770ecc;
assign v377b5aa = hmaster3_p & v3a55c48 | !hmaster3_p & !v377463d;
assign v37589e1 = hmaster0_p & v3732eb2 | !hmaster0_p & v3a658cf;
assign v37577b7 = hbusreq4_p & v3a6f12a | !hbusreq4_p & v373c4d4;
assign v3759519 = hmaster2_p & v3a710c6 | !hmaster2_p & v37716c3;
assign v377b038 = hgrant4_p & v3742241 | !hgrant4_p & v3a5bc04;
assign v3a700db = hmaster2_p & v3a62bae | !hmaster2_p & v3758df6;
assign v373bac6 = hmaster0_p & v375fdc9 | !hmaster0_p & v373931a;
assign v3a554a6 = hbusreq6 & v3a619c0 | !hbusreq6 & !v8455ab;
assign v3a64f7e = hbusreq0 & v374b3bf | !hbusreq0 & v8455ab;
assign v3741e9d = hbusreq1 & v3a63621 | !hbusreq1 & v3a6ebb7;
assign v374dffc = hgrant6_p & v8455ab | !hgrant6_p & v3a6efd2;
assign v37274c2 = hlock0_p & v3a6143b | !hlock0_p & v376b2e9;
assign v3725e12 = hlock8_p & v3a545c8 | !hlock8_p & v3731d66;
assign v37644e0 = hgrant6_p & v8455ca | !hgrant6_p & v3a662fe;
assign v3a6f9c4 = hbusreq0 & v3741ae7 | !hbusreq0 & v373e814;
assign v372a7c1 = hbusreq7 & v37639fa | !hbusreq7 & v377da29;
assign v3a6ff89 = hmaster1_p & d38ecb | !hmaster1_p & v377b3b0;
assign v3a6f64d = hmaster1_p & v373b887 | !hmaster1_p & v3a5a162;
assign v377cece = hlock2 & v376195f | !hlock2 & v3748755;
assign v3729eb8 = hbusreq8_p & v3a6738e | !hbusreq8_p & v376c8a4;
assign v3725a39 = hmaster1_p & v373ce2b | !hmaster1_p & v37702c5;
assign v3a6a6e1 = hmaster0_p & v3a635ea | !hmaster0_p & v3751a97;
assign v3776fe2 = hbusreq1_p & v3a70607 | !hbusreq1_p & v8455ab;
assign v376a0fc = hlock0 & v373f0ee | !hlock0 & d5ffe1;
assign v3757b39 = hbusreq5_p & v3756012 | !hbusreq5_p & v372eb90;
assign v2acaeeb = hmaster1_p & v3a60888 | !hmaster1_p & v3a299f8;
assign v3740374 = hgrant2_p & v39a53b3 | !hgrant2_p & v3a6a1e9;
assign v3a5ed64 = jx0_p & v23fde7f | !jx0_p & v3728b1d;
assign v373d029 = hmaster0_p & v372b1dc | !hmaster0_p & v3a641ea;
assign v9a07a5 = hgrant2_p & v8455ab | !hgrant2_p & v375feb1;
assign v3737860 = hbusreq6_p & v373be25 | !hbusreq6_p & !v372935c;
assign v3a66e91 = hlock1 & v37748e5 | !hlock1 & v3a6f428;
assign v374294f = hbusreq7 & v3a60131 | !hbusreq7 & v3a62ba4;
assign v372bf7f = hgrant6_p & v8455ab | !hgrant6_p & v3a6eba5;
assign v3746683 = hbusreq0 & v3a6fd11 | !hbusreq0 & v374a407;
assign v37717a4 = hbusreq4 & v8455b0 | !hbusreq4 & v3770769;
assign v3a580ca = hmaster0_p & v37386f5 | !hmaster0_p & v3a71299;
assign v37664d0 = hbusreq2_p & v377eaf2 | !hbusreq2_p & v3738d63;
assign v3722caa = hmaster2_p & v3762807 | !hmaster2_p & v3a70272;
assign v37630d9 = hlock2_p & v376e914 | !hlock2_p & !v3a658bf;
assign v3a6aef7 = hmaster2_p & v3774bad | !hmaster2_p & v372e4cf;
assign v3a575dc = hmaster0_p & v37355ea | !hmaster0_p & !v375449f;
assign v372b4d8 = hbusreq8 & v377d97d | !hbusreq8 & v3749503;
assign v37688df = hbusreq6 & v3742905 | !hbusreq6 & v375b044;
assign v3a712cc = hmaster1_p & v3a562b7 | !hmaster1_p & bfae74;
assign v377e5a6 = hbusreq7 & v3a5740f | !hbusreq7 & v3a70bf0;
assign v374b57c = hbusreq3 & v3730627 | !hbusreq3 & v3a5980d;
assign v3a70682 = hmaster0_p & v8455ab | !hmaster0_p & !v3a5a226;
assign v37454a8 = hlock4_p & v373e209 | !hlock4_p & v8455e7;
assign v3731b02 = hbusreq4 & v3a6f347 | !hbusreq4 & v3763f6f;
assign v374376b = hbusreq6 & v373b11b | !hbusreq6 & v3a70a7f;
assign v37400aa = hmaster2_p & v3757966 | !hmaster2_p & v3a6f2af;
assign v3a64968 = hbusreq6_p & v3a6f243 | !hbusreq6_p & v377ca3b;
assign v3749caf = hbusreq6_p & v377a461 | !hbusreq6_p & v8455ab;
assign v3a6f4ce = hmaster0_p & a568f8 | !hmaster0_p & v3747586;
assign v3a63e87 = hbusreq6 & v3a5dbc7 | !hbusreq6 & v375de7f;
assign v3a5979b = hbusreq4_p & v37c007b | !hbusreq4_p & v8455ab;
assign v3753fb7 = hmaster0_p & v3a711df | !hmaster0_p & v3764b6e;
assign v37329ec = hgrant4_p & v3776e5b | !hgrant4_p & v37364d2;
assign v376f62e = hlock8_p & v37369df | !hlock8_p & v3a70b2d;
assign v3a713b4 = hmaster1_p & v3775651 | !hmaster1_p & v3762145;
assign v3a710bb = hmaster1_p & v372b1dc | !hmaster1_p & v3a5db5f;
assign v3a6c8b0 = hlock5 & v376b193 | !hlock5 & v377d004;
assign v3768add = hbusreq0_p & v377b24b | !hbusreq0_p & v3753386;
assign v374b42b = hmaster0_p & v8455ab | !hmaster0_p & v3a65e71;
assign v3a683f9 = hmaster1_p & v375d337 | !hmaster1_p & v373ebac;
assign v37500c2 = hgrant6_p & v37346be | !hgrant6_p & v37762b6;
assign v3a6fb27 = hlock4_p & v8455ab | !hlock4_p & !v373c978;
assign v374b00b = hlock8_p & v37720ee | !hlock8_p & v3767c92;
assign v37274ef = hbusreq0 & v372cb28 | !hbusreq0 & v8455ab;
assign v374c0e3 = hbusreq4 & v376641b | !hbusreq4 & v376728e;
assign v3a701d8 = hgrant6_p & v37792d9 | !hgrant6_p & !v8455ab;
assign v3a6b078 = hmaster1_p & v3735b5a | !hmaster1_p & v3a7127d;
assign v375a319 = hbusreq5_p & v375b8a2 | !hbusreq5_p & v37729fa;
assign v374b589 = hbusreq8_p & v3737808 | !hbusreq8_p & v3737143;
assign v374a565 = hbusreq7 & v373852b | !hbusreq7 & v3a572ee;
assign v3a6f4d5 = hmaster1_p & v3738944 | !hmaster1_p & v3761719;
assign v373a36a = hlock8 & v377aa4d | !hlock8 & ac8c4a;
assign v3a70482 = hbusreq7 & v376a1c9 | !hbusreq7 & v3774bc0;
assign v3774109 = hlock1_p & v3a6f574 | !hlock1_p & v8455ab;
assign v3a5ab7b = hmaster1_p & v3a635ea | !hmaster1_p & v3a56687;
assign v3a655d2 = hmaster1_p & v37784d0 | !hmaster1_p & v3a6f33e;
assign v3a6224d = hlock2 & v3736901 | !hlock2 & v3757d20;
assign v372c834 = hbusreq7_p & v374db33 | !hbusreq7_p & v8455ab;
assign v37292f4 = hgrant3_p & v3a653e4 | !hgrant3_p & !v375c5cf;
assign v374f397 = hmaster2_p & v3a71410 | !hmaster2_p & v374f968;
assign v3a676c6 = hlock5 & v3a6624e | !hlock5 & v3775606;
assign v375f452 = hgrant4_p & v8455ab | !hgrant4_p & v3767b88;
assign v3a5c026 = hmaster2_p & v3757e2f | !hmaster2_p & v8455ab;
assign v39eb4cb = hlock6 & v3a58cf7 | !hlock6 & v3806c41;
assign v3a7082a = hbusreq3_p & v3a635ea | !hbusreq3_p & bba7f1;
assign v374f48b = hbusreq7_p & v20930fa | !hbusreq7_p & v8455ab;
assign v377984a = hmaster0_p & v377caa3 | !hmaster0_p & v377bbf7;
assign v374297b = hgrant4_p & v8455ab | !hgrant4_p & v377640c;
assign v3751285 = hmaster0_p & v3727d4d | !hmaster0_p & v37399d0;
assign v3771ce8 = hbusreq5_p & v3756577 | !hbusreq5_p & v373edd6;
assign v372562b = hgrant6_p & v377b6ce | !hgrant6_p & v377184d;
assign v374caa8 = hmaster1_p & v377a1ee | !hmaster1_p & v3752caa;
assign v377789d = hbusreq4 & v3743a4d | !hbusreq4 & !v376a246;
assign v374e519 = hmaster2_p & v3a65369 | !hmaster2_p & v377f61e;
assign v373325b = hgrant6_p & v372bfa1 | !hgrant6_p & v3a664ba;
assign v376ecae = hmaster1_p & v37793e4 | !hmaster1_p & v37717ee;
assign v375bb11 = hmaster1_p & v375527f | !hmaster1_p & v3a57891;
assign v3761ed2 = hbusreq0 & v3a5f0cf | !hbusreq0 & v3a5dd7f;
assign v3760e47 = hgrant0_p & v3a69b5f | !hgrant0_p & v3a6f169;
assign v3a67729 = hbusreq6 & v2092aba | !hbusreq6 & v3a62f0b;
assign v37234f5 = hlock0_p & v3a7104b | !hlock0_p & v375ecc7;
assign v376543b = hmaster1_p & v8cd321 | !hmaster1_p & v376314e;
assign v3a70863 = hmaster1_p & v3a67e13 | !hmaster1_p & v3728d9c;
assign v376cbb7 = hbusreq0 & v3a63f06 | !hbusreq0 & v374db32;
assign v3768ce2 = hbusreq1_p & v3726570 | !hbusreq1_p & !v377baa6;
assign v3776c04 = hbusreq4_p & v373bfab | !hbusreq4_p & v3a70d01;
assign v3a5e245 = hmaster1_p & v37386f5 | !hmaster1_p & v3a580ca;
assign v3a6f568 = hbusreq8_p & v377244a | !hbusreq8_p & v3a6ff5e;
assign v3753030 = hbusreq0 & v3a70f18 | !hbusreq0 & v3764ced;
assign v372efb1 = hmaster2_p & v8455ab | !hmaster2_p & v374caab;
assign v3775fae = hgrant2_p & v3a6f02f | !hgrant2_p & v3748bf9;
assign v94c82c = hgrant8_p & v8455ab | !hgrant8_p & !b8cdcc;
assign v3a6de4f = hmaster2_p & v3a635ea | !hmaster2_p & v373a341;
assign v376910a = hgrant5_p & v3a6f396 | !hgrant5_p & v3a5bd9c;
assign v3a6ccc6 = hbusreq7 & v3744657 | !hbusreq7 & v3a60276;
assign v3779958 = hbusreq5 & v3a6f79f | !hbusreq5 & v3764dda;
assign v3a6fb20 = hmaster1_p & v8455ab | !hmaster1_p & aac06c;
assign v372fcfc = hbusreq7 & v375194a | !hbusreq7 & v37750a5;
assign v3751e76 = hbusreq4_p & v3729ed7 | !hbusreq4_p & v3739ba9;
assign v3a66b88 = hbusreq6 & v3778fda | !hbusreq6 & v3739da7;
assign v3731f3c = hmaster0_p & v8455ab | !hmaster0_p & !v377d769;
assign v375da55 = hmaster1_p & v374c5fc | !hmaster1_p & v23fd89c;
assign v3768af7 = hbusreq0 & v374ba61 | !hbusreq0 & v3a6632a;
assign v372b881 = hgrant4_p & v37476bd | !hgrant4_p & v3a70c72;
assign v37260af = hgrant5_p & v8455c6 | !hgrant5_p & v3752edc;
assign v3a61a15 = hmaster0_p & v3a54aa0 | !hmaster0_p & v3749f86;
assign v3757966 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f3bb;
assign v377d785 = hgrant6_p & v3729214 | !hgrant6_p & v376a399;
assign v372a536 = hlock4_p & v3730de2 | !hlock4_p & v3777a8c;
assign v3a6cef4 = hbusreq3 & v373d78b | !hbusreq3 & v8455ab;
assign v3a6a236 = hlock6 & v38072fd | !hlock6 & v3a715ae;
assign v372fe10 = hgrant6_p & v3751c68 | !hgrant6_p & v2aca977;
assign v3a5687e = hmaster2_p & v3a635ea | !hmaster2_p & v373bd76;
assign v373366b = hgrant4_p & v8455e7 | !hgrant4_p & v37770c9;
assign v375034b = hbusreq6_p & v3a64252 | !hbusreq6_p & v3752f21;
assign v37465d4 = hbusreq8 & v37586d1 | !hbusreq8 & v3768734;
assign v3752e63 = hbusreq2_p & v3777412 | !hbusreq2_p & v8455ab;
assign v3778aac = hbusreq5_p & v3773340 | !hbusreq5_p & v372b33d;
assign v37476b8 = hmaster0_p & v3a700e2 | !hmaster0_p & v3a6f40d;
assign v3777ac3 = hmaster2_p & v9af7ec | !hmaster2_p & v375649e;
assign v377c7ce = hgrant6_p & v3779060 | !hgrant6_p & v3a7152c;
assign v3a293c5 = hmastlock_p & v3745b85 | !hmastlock_p & !v8455ab;
assign v3743ea8 = hbusreq6 & v372c3d4 | !hbusreq6 & v3760f87;
assign v3a701cb = hmaster1_p & v3748a16 | !hmaster1_p & v8455ab;
assign v3741a71 = hmaster2_p & v3a635ea | !hmaster2_p & v3769ecf;
assign v3757082 = hbusreq1_p & v375dbc6 | !hbusreq1_p & !v8455ab;
assign v376f5ed = hbusreq8 & v375c735 | !hbusreq8 & v3768734;
assign v37554a1 = hbusreq4_p & v3a6f044 | !hbusreq4_p & v3a713c8;
assign v3771fea = hmaster1_p & v3a62f70 | !hmaster1_p & ae4185;
assign v380649c = hbusreq6_p & v3759b2f | !hbusreq6_p & !v373be25;
assign v372fc81 = hready & v3a70fa5 | !hready & v3a713e1;
assign v3743def = hlock8 & v3a6f551 | !hlock8 & v3a595fd;
assign v377228d = hgrant2_p & v375afc1 | !hgrant2_p & v8455ab;
assign v377c9b1 = hmaster2_p & v3a6f22c | !hmaster2_p & v372a0b0;
assign v373399e = hbusreq3_p & v8455ab | !hbusreq3_p & v3a6a939;
assign v372475d = hbusreq4_p & v375f169 | !hbusreq4_p & !v3a70af5;
assign v3a6f2ee = hmaster0_p & v376d9c6 | !hmaster0_p & v3738e6e;
assign v3a66c14 = hgrant5_p & v3731c27 | !hgrant5_p & v3724345;
assign v3a570f5 = hlock6_p & v3776441 | !hlock6_p & v8455e7;
assign v3752b5c = hbusreq5_p & v3a63628 | !hbusreq5_p & v3741ab9;
assign v372e02c = hbusreq7 & c80162 | !hbusreq7 & v375ab92;
assign v3738087 = hbusreq7 & v374fa18 | !hbusreq7 & v373a8a1;
assign v3777749 = hgrant3_p & ae7027 | !hgrant3_p & v3a65546;
assign v373c631 = hbusreq2 & v37665bf | !hbusreq2 & v8455ab;
assign v3a5ca02 = hlock0_p & v3a6b2ef | !hlock0_p & v3757811;
assign v3757888 = hmaster2_p & v37782c9 | !hmaster2_p & v3a5fc34;
assign v3a6fbdd = hbusreq6_p & v3a6600c | !hbusreq6_p & v8455ab;
assign v3a66ab2 = hmaster2_p & v376b397 | !hmaster2_p & v3a6eaff;
assign v3a68d0e = hgrant4_p & v8455c2 | !hgrant4_p & v376fca4;
assign v3a70635 = hlock2_p & v3746b6e | !hlock2_p & v8455b7;
assign v3a7082c = hlock4 & v3758a9c | !hlock4 & v3a70791;
assign v8455ed = hgrant2_p & v8455ab | !hgrant2_p & !v8455ab;
assign v374721d = hlock1_p & v3a70edc | !hlock1_p & v372a837;
assign v3757f0d = hlock4_p & v3a6cf6a | !hlock4_p & v8455ab;
assign v3a68170 = hbusreq7_p & v372d691 | !hbusreq7_p & v376ae9f;
assign v37266d9 = hbusreq7_p & v3a6f74f | !hbusreq7_p & !v3a69df3;
assign v376062f = hlock4 & v3a7026f | !hlock4 & v3778787;
assign v374893c = hmaster0_p & v1e3778d | !hmaster0_p & v8455ab;
assign v374b074 = hbusreq5_p & cb09e1 | !hbusreq5_p & v3a5c196;
assign v3a57829 = hbusreq2_p & v3756716 | !hbusreq2_p & v8455ab;
assign v86d727 = hbusreq7 & v374bd7d | !hbusreq7 & v376e9ed;
assign v3a70244 = hlock4 & v3a71615 | !hlock4 & v3a6fd8f;
assign v3a6f81c = hbusreq5 & v376f51c | !hbusreq5 & v3a706c9;
assign v375c3eb = hlock4 & v37671b7 | !hlock4 & v373f4fb;
assign v376c5d3 = hmaster0_p & v3a61a7f | !hmaster0_p & v375f69e;
assign v3a60f22 = hbusreq6 & v373cd16 | !hbusreq6 & v8455ab;
assign v3a5e817 = hbusreq1_p & v37728d0 | !hbusreq1_p & !v8455ab;
assign v3756809 = hmaster0_p & v376ba62 | !hmaster0_p & v3778c61;
assign v3a66ea0 = hbusreq7 & v376a06c | !hbusreq7 & v373168f;
assign v37362fd = hlock7_p & v376848c | !hlock7_p & v3736320;
assign v377910a = hlock4 & v3770d22 | !hlock4 & v3a6774e;
assign v3a70532 = hlock4 & v377eaa3 | !hlock4 & v3a70791;
assign v37398f3 = hbusreq1_p & v3a6db4b | !hbusreq1_p & !v374e4c9;
assign v376957a = hbusreq8 & v3a60134 | !hbusreq8 & v3a5e611;
assign v377499f = hbusreq3_p & v37625a8 | !hbusreq3_p & !v2092faa;
assign v3a5b4ca = hbusreq5_p & v3a7126e | !hbusreq5_p & v3a5a1ef;
assign v3a61a76 = hbusreq0 & v3a70336 | !hbusreq0 & v3a70d44;
assign v37346be = hbusreq3_p & v8455ab | !hbusreq3_p & !v3a637dd;
assign v2093234 = hbusreq6 & v3744f0d | !hbusreq6 & v3a6f61f;
assign v373d68a = hmaster0_p & v374287d | !hmaster0_p & v3a70574;
assign v37578d4 = hbusreq6_p & v373997b | !hbusreq6_p & v37738fc;
assign v3745b07 = hbusreq3 & v3a5600a | !hbusreq3 & v373b3fb;
assign v374e8f7 = hbusreq8 & v376c6b3 | !hbusreq8 & v372d5e5;
assign v3a700b7 = hlock0 & v3748797 | !hlock0 & v3750c12;
assign v3a61336 = hmaster0_p & v377e784 | !hmaster0_p & v3a6b27e;
assign v377aae4 = hbusreq5_p & v377a8c3 | !hbusreq5_p & v3779470;
assign v3a605d3 = hgrant5_p & v3a67af1 | !hgrant5_p & v375be11;
assign v3a5784f = hlock0 & v3a58038 | !hlock0 & v375c52f;
assign v3a5a25a = hmaster3_p & v375d512 | !hmaster3_p & v3777d70;
assign v3a70b77 = hmaster0_p & v3747b2b | !hmaster0_p & v37412f3;
assign v3a592f7 = hready & v3a539ee | !hready & !v8455ab;
assign v3a6fcdc = hlock5 & v37548a5 | !hlock5 & v37318e3;
assign v3a701d3 = hgrant3_p & v3a68aa8 | !hgrant3_p & v3255a31;
assign v3a6f22b = hbusreq3_p & v3762700 | !hbusreq3_p & v8455b3;
assign v3a5538a = hlock6_p & v2aca977 | !hlock6_p & v8455ab;
assign v3a7101a = hlock8_p & v2acafeb | !hlock8_p & v3a6a03c;
assign v3775928 = hmaster2_p & v375058e | !hmaster2_p & v376a6f1;
assign v3a64718 = hbusreq5_p & v3a66f8d | !hbusreq5_p & v3769740;
assign v373ac15 = hmaster2_p & v8455ab | !hmaster2_p & !v376cf62;
assign v375119e = hmaster2_p & v37771a8 | !hmaster2_p & v37764c0;
assign v3763f05 = jx2_p & v3a6b368 | !jx2_p & v37432e1;
assign v3a70274 = hlock0_p & v375356f | !hlock0_p & v3a5e3d0;
assign v23fdbe6 = hmaster3_p & v373083d | !hmaster3_p & v374a528;
assign v3a60358 = hmaster2_p & d1e3dd | !hmaster2_p & v37674f6;
assign v375ec0b = hbusreq4 & v3a5f07a | !hbusreq4 & v3756018;
assign v3a70f74 = hlock2 & v3a700b5 | !hlock2 & v376f768;
assign v372da0b = hbusreq5_p & v3a63f9a | !hbusreq5_p & v3a59c5e;
assign v372379e = hmaster2_p & v37793a4 | !hmaster2_p & v375a697;
assign v37541ff = hbusreq0 & v372f02f | !hbusreq0 & v8455ab;
assign v3a5a8bf = hlock6_p & v3724a4b | !hlock6_p & adf78a;
assign v374813d = hgrant4_p & v376c1f7 | !hgrant4_p & v3a6eec9;
assign v375a2b5 = hgrant6_p & v3725fe1 | !hgrant6_p & v3722a0a;
assign v3743f54 = hlock0 & v37651c2 | !hlock0 & v373029d;
assign v2619ac3 = hgrant3_p & v3a6c2b6 | !hgrant3_p & v374c23c;
assign v372bcb0 = hgrant2_p & v3a70645 | !hgrant2_p & v3728d2a;
assign v3a5f458 = hgrant5_p & v37426ea | !hgrant5_p & v3a70ce8;
assign v3a7141c = hgrant4_p & v3774c1b | !hgrant4_p & v3736d03;
assign v375b0e4 = hmaster2_p & v3a6d21e | !hmaster2_p & v2ff8cae;
assign v3741906 = hgrant4_p & v8455ab | !hgrant4_p & v3a61d77;
assign v375d417 = hmaster0_p & v3a689bb | !hmaster0_p & v375842f;
assign v3758cc6 = hgrant7_p & v3a70c83 | !hgrant7_p & v376114f;
assign v374c98c = hgrant5_p & v3740a8a | !hgrant5_p & v3733d66;
assign v3723f2a = hbusreq4 & v3765e6a | !hbusreq4 & v3a6fba6;
assign v3a6ebdb = hgrant3_p & v374383b | !hgrant3_p & v3a62ed6;
assign v3a6fb6f = hmaster1_p & v377030a | !hmaster1_p & v3a65155;
assign v35b7168 = hbusreq5_p & v373014d | !hbusreq5_p & v377d107;
assign v3a6ff88 = hbusreq8 & v3a5f622 | !hbusreq8 & v375455d;
assign v3766f13 = hlock8_p & v37347cd | !hlock8_p & v3779e38;
assign v377aefe = hmaster2_p & v37728a5 | !hmaster2_p & v3775537;
assign v3a706d9 = hbusreq5 & v374fefc | !hbusreq5 & v376ab39;
assign v3729360 = hmaster2_p & v8455b0 | !hmaster2_p & !v8455ab;
assign v372d9a1 = hbusreq5_p & v1e379b9 | !hbusreq5_p & v8455ab;
assign v37522e4 = hbusreq0 & v3a6fefc | !hbusreq0 & v3731230;
assign v3a28da6 = decide_p & v37293c2 | !decide_p & v8455f9;
assign v3a70051 = hmaster2_p & v35b774b | !hmaster2_p & v37598ab;
assign v375521a = hbusreq8 & v3744824 | !hbusreq8 & v3a6f45d;
assign v3777efb = hbusreq5_p & v37360c0 | !hbusreq5_p & !v3749a4c;
assign v376f7a0 = hgrant6_p & v8455ca | !hgrant6_p & v375bc08;
assign v3758435 = hmaster1_p & v3a7069a | !hmaster1_p & v375b1a0;
assign v373d223 = hmaster1_p & v374502e | !hmaster1_p & v3a66645;
assign v37585e6 = hbusreq1 & v376b4e1 | !hbusreq1 & !v8455ab;
assign v3a70cc8 = hmaster0_p & v3756bd8 | !hmaster0_p & v3a5f992;
assign v3758f1b = hbusreq6 & v3756c25 | !hbusreq6 & v374f35a;
assign v3a6fe90 = hlock0_p & v3745f76 | !hlock0_p & !v8455ab;
assign v3777070 = hbusreq8 & v3a70d6b | !hbusreq8 & v8455ab;
assign v3744dca = hbusreq0 & v3a7104d | !hbusreq0 & v8455ab;
assign v3739386 = hbusreq6 & v3753e00 | !hbusreq6 & v376ef7a;
assign v373bb0f = hgrant3_p & v3758c35 | !hgrant3_p & v374b5d9;
assign v3741890 = hmaster3_p & v3a6f83f | !hmaster3_p & v377a5d4;
assign v3a7163c = hlock6_p & v37685bb | !hlock6_p & v373f503;
assign v3770d6d = hbusreq2 & v3777311 | !hbusreq2 & v3a56642;
assign v37354c1 = hmaster2_p & v376fcc3 | !hmaster2_p & !v3735b3e;
assign hgrant3 = !v3377c79;
assign v3a70480 = hbusreq6_p & v37504a9 | !hbusreq6_p & v372348c;
assign v375b40c = hbusreq6_p & v37232c0 | !hbusreq6_p & !v372df2a;
assign v374d273 = hlock2 & d9a7db | !hlock2 & v37415b2;
assign v3746e47 = hgrant2_p & v8455ab | !hgrant2_p & v3a57829;
assign v375c946 = hbusreq2 & v3754877 | !hbusreq2 & v3735525;
assign v3a6bee8 = hlock5_p & v8455ab | !hlock5_p & v374edba;
assign v3777d37 = hbusreq5 & v3766792 | !hbusreq5 & v3728f6d;
assign v3736113 = hmaster0_p & v3a6f4bd | !hmaster0_p & v373d9b3;
assign v3773ab1 = hbusreq5_p & v3a5395c | !hbusreq5_p & v3773838;
assign v3a70544 = hbusreq3_p & v3a635ea | !hbusreq3_p & v37577d8;
assign v3747b4e = hmaster1_p & v3a65b0a | !hmaster1_p & v376a411;
assign v3a6fe5c = hmaster2_p & v377d232 | !hmaster2_p & v374ccb3;
assign v377adbd = hmaster1_p & v3a709c3 | !hmaster1_p & !v373adb9;
assign v373e475 = hlock5_p & v3a6ff25 | !hlock5_p & v37717d0;
assign v376278c = hgrant3_p & v8455ab | !hgrant3_p & v3724121;
assign v372def3 = hmaster2_p & v375d9b1 | !hmaster2_p & !v3a6eb6e;
assign v375d1d0 = hmaster1_p & v8455ab | !hmaster1_p & d7cff8;
assign v23fe343 = hmaster1_p & v3a578af | !hmaster1_p & v8455ab;
assign v3a6aaea = hmaster2_p & v372433d | !hmaster2_p & !v8455ab;
assign v3808e6b = hmaster0_p & v3a6efc7 | !hmaster0_p & v3a7026a;
assign v3751807 = hburst0 & v37295fe | !hburst0 & v377d126;
assign v376a383 = hlock7 & v375c924 | !hlock7 & v3a70cd7;
assign v37772bf = hlock0_p & v3a68426 | !hlock0_p & v3a6f972;
assign v3a56f66 = hgrant3_p & ae7027 | !hgrant3_p & v376b33c;
assign v375d9ad = hmaster0_p & v3736610 | !hmaster0_p & v373f5ab;
assign v3a6ff8c = hbusreq5_p & v374a11d | !hbusreq5_p & !v8455ab;
assign v3a713c5 = hmaster0_p & v3a5f02e | !hmaster0_p & v3807a23;
assign v3a6f9e4 = hmaster2_p & v8455ab | !hmaster2_p & v37728c2;
assign v3742657 = hgrant2_p & v3a70115 | !hgrant2_p & v3a6dd65;
assign v375f742 = hbusreq5 & v3a6ffd9 | !hbusreq5 & v38070ea;
assign a5c257 = hmaster1_p & v3a6c4e4 | !hmaster1_p & v373e72e;
assign v3743e29 = hlock2_p & v3750aea | !hlock2_p & v3a5f991;
assign v3a2a348 = hbusreq2_p & v3a5c945 | !hbusreq2_p & !v3a619c0;
assign v3739166 = stateG10_1_p & v3774b25 | !stateG10_1_p & v376e00a;
assign v3a6079f = hbusreq2_p & v3a583dc | !hbusreq2_p & v37773c1;
assign v372ec1c = hbusreq0_p & v3723430 | !hbusreq0_p & v8455ab;
assign v374b13e = hmaster2_p & v3a5a510 | !hmaster2_p & v3759032;
assign v2092b2c = hmaster0_p & v3769ae2 | !hmaster0_p & v3742121;
assign v2092bae = hgrant3_p & v3a6505b | !hgrant3_p & v3a5b6ca;
assign v3a704ca = hmaster0_p & v3a71350 | !hmaster0_p & v3a5ef76;
assign v374b9f9 = hbusreq4 & v3a711e0 | !hbusreq4 & v3777666;
assign v3a6f0bd = hbusreq4 & v8455b0 | !hbusreq4 & v3a708a2;
assign v3a592bb = hbusreq8_p & v3a70578 | !hbusreq8_p & v3a5d62d;
assign v373706e = hmaster1_p & v372673d | !hmaster1_p & v37691d1;
assign v3725bd2 = hbusreq7_p & v3753aa5 | !hbusreq7_p & v3a6f2f8;
assign v39ea0c5 = hlock4_p & v3a70cdb | !hlock4_p & v8455b0;
assign v375c705 = hbusreq2 & v3a5d469 | !hbusreq2 & v3a69487;
assign v3a668da = hmaster2_p & v3a635ea | !hmaster2_p & v373ee52;
assign v3a7133d = hbusreq4_p & v3722f65 | !hbusreq4_p & v1e378da;
assign v3a70bff = hbusreq6 & v373081f | !hbusreq6 & v3a635ea;
assign v3a704ff = hlock7 & v3777c9b | !hlock7 & v375b56c;
assign v377222b = hbusreq3 & v3a63805 | !hbusreq3 & v8455b0;
assign v3776492 = hbusreq4 & v3750d4c | !hbusreq4 & v380988c;
assign v3a5db7f = hmaster0_p & v3733c51 | !hmaster0_p & v3a71420;
assign v3a6fc7b = hbusreq2_p & v3a6f22f | !hbusreq2_p & v3773856;
assign v3742725 = hmaster2_p & v3a635ea | !hmaster2_p & v37320ff;
assign v3a63f29 = hmaster2_p & v8455ab | !hmaster2_p & v3a6a8ee;
assign v3728f87 = hgrant2_p & d35b26 | !hgrant2_p & v37512a0;
assign v3737bff = hbusreq0_p & v38072fd | !hbusreq0_p & v3a66e91;
assign v37609e3 = hbusreq5 & v3725d18 | !hbusreq5 & v8455ab;
assign cae8ef = hbusreq7 & v3a67f12 | !hbusreq7 & !v8455b5;
assign v3748059 = hbusreq8 & v39eaae9 | !hbusreq8 & v3723d79;
assign v376b86f = hmaster2_p & v3a70641 | !hmaster2_p & v8455ab;
assign v3a707f1 = hgrant0_p & v8455ab | !hgrant0_p & v374710b;
assign v3a6f1ee = hbusreq6_p & v3a70788 | !hbusreq6_p & v209324e;
assign v3a70ce3 = stateG3_2_p & v8455ab | !stateG3_2_p & v3a712be;
assign v37362b5 = hlock0 & v3a6a934 | !hlock0 & v3a58a1b;
assign v3731383 = hbusreq6 & v3746265 | !hbusreq6 & !v8455ab;
assign v375f0d4 = hmaster1_p & v3a6ff36 | !hmaster1_p & !v3a6e0cc;
assign v373a876 = hmaster0_p & v3a61a7f | !hmaster0_p & v3741039;
assign v3a708ef = hgrant0_p & v8455ab | !hgrant0_p & !v3a6e7a7;
assign v3a7051a = hbusreq2 & v3775303 | !hbusreq2 & v8455ab;
assign v3768eb1 = hgrant3_p & v37c1a6f | !hgrant3_p & v3757746;
assign v3a5bb4e = hbusreq5 & c52384 | !hbusreq5 & v37554cd;
assign v3a6f5e4 = hmaster1_p & v3748266 | !hmaster1_p & !v3a69fcf;
assign v37605c1 = hbusreq2_p & v37261df | !hbusreq2_p & !v3a5ae7d;
assign v3a70bf4 = hgrant4_p & v37728a5 | !hgrant4_p & v37707d5;
assign v376ce06 = hmaster0_p & v375a023 | !hmaster0_p & v3a6fdea;
assign v3a7085c = hbusreq5 & v3a58687 | !hbusreq5 & v3742c68;
assign v3808ceb = hbusreq8_p & v372a027 | !hbusreq8_p & v372a48e;
assign v374544d = hlock8 & v376ae9f | !hlock8 & v3a6f3c2;
assign v37354f8 = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3a6617b;
assign v3745dae = hmaster1_p & v87be38 | !hmaster1_p & v3a5cfb0;
assign v3a5637b = hmaster0_p & v3a67dab | !hmaster0_p & v376db34;
assign v374b024 = hbusreq7_p & v3766260 | !hbusreq7_p & bfa92a;
assign bf29af = hlock0 & v37696b6 | !hlock0 & v3778430;
assign v3a5a2e4 = hlock6_p & v372a00b | !hlock6_p & v3a6fb2b;
assign v376a220 = hgrant2_p & b95be3 | !hgrant2_p & v3738766;
assign v3730343 = hbusreq0_p & v3809adf | !hbusreq0_p & !v3a70c07;
assign v3a57484 = hbusreq2_p & v376441d | !hbusreq2_p & v3737ad2;
assign v3a5b850 = hburst0 & v3a6ac2a | !hburst0 & v3a6fad0;
assign v375652a = hbusreq5_p & v375c3b6 | !hbusreq5_p & v1e37c60;
assign v372463a = hgrant4_p & v8455ab | !hgrant4_p & v3a5bff1;
assign v3a6eede = hbusreq5 & v3755b5c | !hbusreq5 & v373ca3d;
assign v373f91b = hbusreq2 & v3a6a939 | !hbusreq2 & v8455ab;
assign v3a708aa = hmastlock_p & v374592e | !hmastlock_p & v8455ab;
assign v373308b = hmaster2_p & v373b288 | !hmaster2_p & v376bb26;
assign v3a6de06 = hbusreq5 & bdb538 | !hbusreq5 & v373d5f4;
assign v3a6f433 = hbusreq5_p & v374a8e2 | !hbusreq5_p & v3a5a24d;
assign v375b736 = hbusreq2 & v372da4f | !hbusreq2 & v373c480;
assign v373c8ff = hlock6_p & v372d630 | !hlock6_p & v3a6f5d1;
assign v377e3ce = hbusreq4 & v3729852 | !hbusreq4 & v8455ab;
assign v3a71251 = hmaster2_p & v373cddc | !hmaster2_p & v8455ab;
assign v3a5ce35 = hmaster2_p & v3379037 | !hmaster2_p & v3765e46;
assign v37487f5 = hbusreq3 & v372eaaf | !hbusreq3 & v377395f;
assign v3775107 = hbusreq0_p & v8455ab | !hbusreq0_p & v374fb58;
assign v37484e7 = hbusreq7_p & v37249fe | !hbusreq7_p & v37774b6;
assign v3726605 = hgrant4_p & v3a6a213 | !hgrant4_p & d27e8c;
assign v3a6f046 = jx1_p & v8455ab | !jx1_p & v377f0dc;
assign v3a6fe99 = hmaster0_p & v3a6eff4 | !hmaster0_p & v8455e7;
assign v376a946 = hlock7 & v374bdac | !hlock7 & v3727a6d;
assign v3a6e005 = hlock5_p & v3a6b285 | !hlock5_p & !v377c49c;
assign v3a715fa = hmaster1_p & v374502e | !hmaster1_p & v374ddc7;
assign v37299fa = hgrant6_p & v3a6c7fe | !hgrant6_p & v37265f6;
assign v374b8c5 = hbusreq0 & v3a5a051 | !hbusreq0 & v3a6efb2;
assign v374e21e = hbusreq5_p & v3778138 | !hbusreq5_p & v374d969;
assign v3734db5 = hbusreq2_p & v37574d2 | !hbusreq2_p & v373b288;
assign v3773e41 = hbusreq2_p & v3a63f30 | !hbusreq2_p & !v3a672c9;
assign v3a5e2ee = hbusreq2 & v3740171 | !hbusreq2 & v8455e7;
assign v3765cd5 = hlock5_p & v8455ab | !hlock5_p & v1e3737d;
assign v374820d = hbusreq4_p & v37588c4 | !hbusreq4_p & !v3a7107a;
assign v373ac39 = hgrant2_p & v8455e7 | !hgrant2_p & v372efbe;
assign v3a6fe8e = hgrant2_p & v3758472 | !hgrant2_p & !v3a6f0b2;
assign v375e23b = hbusreq8_p & v3737103 | !hbusreq8_p & v3a6f786;
assign v376df3c = hmaster0_p & v3a5e24e | !hmaster0_p & v3770093;
assign v8c890d = hbusreq2_p & v372a711 | !hbusreq2_p & v3a5affd;
assign v372a958 = hbusreq3 & v373fe5e | !hbusreq3 & v8455ab;
assign v3a5fe00 = hmaster2_p & v37678fc | !hmaster2_p & v3760f4e;
assign v3752aa3 = hgrant5_p & v8455ab | !hgrant5_p & v3770b26;
assign v374e7fa = hbusreq5_p & v37711f0 | !hbusreq5_p & v37724fc;
assign v375a5b6 = hbusreq0 & v3774fa6 | !hbusreq0 & v376d566;
assign v37455cd = hmaster2_p & v3a707b5 | !hmaster2_p & v3a70272;
assign v3a683c1 = hmaster2_p & v3753dab | !hmaster2_p & v3a6f993;
assign v3735055 = hbusreq7 & v3765d9e | !hbusreq7 & v3a5fc34;
assign v3a5c350 = hbusreq6_p & v37288db | !hbusreq6_p & v3a70397;
assign v375dbe0 = hgrant3_p & v8455ab | !hgrant3_p & !v3a6fa9f;
assign v3a5a854 = hmaster0_p & v3a5e665 | !hmaster0_p & b2ea29;
assign v3733c9e = hbusreq0 & v372dde7 | !hbusreq0 & v3a6af0b;
assign v3738ed2 = hmaster0_p & v375b429 | !hmaster0_p & v3760be5;
assign v3a6f6cb = hbusreq5 & d3a479 | !hbusreq5 & v8455ab;
assign v3a70adb = hmaster0_p & v3a70557 | !hmaster0_p & v373296d;
assign v3a70232 = hbusreq2_p & v2092eaf | !hbusreq2_p & v8455ab;
assign v375c41e = hbusreq4 & v3733e0a | !hbusreq4 & v8455ab;
assign v3a66673 = hbusreq0_p & v375de18 | !hbusreq0_p & !v374cab9;
assign v3a5e611 = hlock7 & v3a6cd4f | !hlock7 & v37305e6;
assign v3a70ed0 = hbusreq7_p & v3a63b69 | !hbusreq7_p & v37542b2;
assign v3a70dfd = hmaster1_p & v3757568 | !hmaster1_p & v3a6f9a7;
assign v372e0b0 = hgrant4_p & v3733d6e | !hgrant4_p & v373d72e;
assign v3a63e68 = hmaster0_p & v3725198 | !hmaster0_p & v373f394;
assign v373b717 = hmaster0_p & v8455ca | !hmaster0_p & !v2ff8e8b;
assign v37555b4 = hmaster0_p & v3a566eb | !hmaster0_p & v3a71207;
assign v360d048 = hbusreq4 & v8455b0 | !hbusreq4 & v3a63805;
assign v3777cb9 = hlock6 & v3a6767d | !hlock6 & v373b759;
assign v3a708c2 = hlock0_p & v3747302 | !hlock0_p & v37538e1;
assign v3a6f3a2 = hmaster2_p & v3768b46 | !hmaster2_p & v377a434;
assign v37690fe = hmaster1_p & v3724e64 | !hmaster1_p & v3a557a1;
assign v3a6fbfc = hgrant0_p & v3a71452 | !hgrant0_p & v3a5a585;
assign v3768685 = hbusreq2_p & v37626d4 | !hbusreq2_p & v8455ab;
assign v3a6f01d = hbusreq7_p & v3a6f769 | !hbusreq7_p & cae8ef;
assign v374b340 = hlock0 & v374a637 | !hlock0 & v37507dd;
assign v3a606b0 = hmaster2_p & v3a702ee | !hmaster2_p & v8455ab;
assign v3740f94 = hmaster2_p & v375e854 | !hmaster2_p & v23fd83f;
assign v3766445 = hlock5 & v3744838 | !hlock5 & v3773cda;
assign v3a59c72 = hmaster1_p & v3a70d99 | !hmaster1_p & v375b4cb;
assign v373133d = hbusreq4_p & v377097a | !hbusreq4_p & v3a62a6d;
assign v3a6bab2 = hlock2 & v37458dc | !hlock2 & v3a623dc;
assign v3736b55 = hmaster0_p & v37429cc | !hmaster0_p & v8455b5;
assign v37399d0 = hmaster2_p & v377bd5c | !hmaster2_p & v37395a4;
assign v376610a = hmaster1_p & v8455e7 | !hmaster1_p & v375818b;
assign v3725f3b = stateG3_1_p & v845601 | !stateG3_1_p & !v845601;
assign v3a62d7d = hbusreq6 & v3760f4e | !hbusreq6 & v8455b3;
assign a54211 = hbusreq2_p & v3774c1b | !hbusreq2_p & !v38099c1;
assign v372809b = hlock7 & v3a6a208 | !hlock7 & v373ac84;
assign v2acaecc = hlock4_p & v3a56642 | !hlock4_p & v3730ffe;
assign v372e4cf = hbusreq4_p & v3a65bad | !hbusreq4_p & v8455ab;
assign v37523ea = hmaster0_p & v376aa57 | !hmaster0_p & v3a64147;
assign v372c007 = hbusreq6_p & v39a537f | !hbusreq6_p & !v1e38224;
assign v375cda1 = hmaster1_p & v3a6c6b1 | !hmaster1_p & v3a6f50c;
assign v375efa1 = hbusreq6_p & v374c33a | !hbusreq6_p & v8455ab;
assign v375ac48 = hbusreq3_p & v8455ab | !hbusreq3_p & v3a71682;
assign v37340b4 = hmaster0_p & v375b429 | !hmaster0_p & v3a6ff98;
assign v3a5e19b = hgrant5_p & v8455ab | !hgrant5_p & v373dff6;
assign v377b015 = hmaster2_p & v8455ab | !hmaster2_p & v3761d38;
assign v3a59c0b = jx1_p & v3a629a9 | !jx1_p & v37751ae;
assign v37505e1 = hmaster1_p & v373a27c | !hmaster1_p & v3764437;
assign v375f653 = hbusreq6_p & v373642c | !hbusreq6_p & !v8455ca;
assign v3a5ba5b = jx3_p & v3779955 | !jx3_p & v376c0dc;
assign v37445e5 = hlock0 & v3a6f044 | !hlock0 & v377a8e0;
assign v374465a = hbusreq4_p & v372ccc4 | !hbusreq4_p & v8455b0;
assign v37255a7 = hbusreq6_p & v372ff3a | !hbusreq6_p & v3a68d2e;
assign v3766f1c = hlock6_p & v3724a6e | !hlock6_p & v3760bd6;
assign v3a66d47 = hmaster0_p & v3a6f926 | !hmaster0_p & v3745b9c;
assign v3a58a8e = hgrant2_p & v3a70dc4 | !hgrant2_p & v3a70cea;
assign v3a70bb2 = hbusreq0_p & v3776670 | !hbusreq0_p & v374288a;
assign v374c4e9 = hbusreq2_p & v37790ef | !hbusreq2_p & v372c0f4;
assign v3a6f746 = hgrant6_p & v3a6fbe4 | !hgrant6_p & v37708e7;
assign v3761c68 = hlock2_p & v37237be | !hlock2_p & bd3d3d;
assign v3730383 = stateG3_2_p & v8455ab | !stateG3_2_p & !v37603af;
assign v376ed2b = hbusreq5_p & v3745181 | !hbusreq5_p & v3a5a04c;
assign c04cff = hmaster2_p & v3a70049 | !hmaster2_p & !v2092eb7;
assign v3750e0b = hmaster0_p & v375cbe2 | !hmaster0_p & !v3764b6e;
assign v3747929 = hbusreq5_p & v373e625 | !hbusreq5_p & v3a6ef5a;
assign v3742cd4 = hbusreq4_p & v8455bf | !hbusreq4_p & v2092abe;
assign v3a6f481 = hbusreq2 & v3743698 | !hbusreq2 & v8455ab;
assign v373cc5c = hbusreq6_p & v377803a | !hbusreq6_p & v374d749;
assign v3751460 = hgrant0_p & v8455ab | !hgrant0_p & v3a70274;
assign v3a6accb = hgrant5_p & v377d496 | !hgrant5_p & v37712e5;
assign v3a6eb98 = hmaster2_p & v380974c | !hmaster2_p & v8455b3;
assign v3736320 = hbusreq7 & v3766048 | !hbusreq7 & v3778901;
assign v3a70296 = hbusreq5_p & v37410bd | !hbusreq5_p & v2acae99;
assign v376604f = hbusreq4 & v3a6fd2d | !hbusreq4 & v3751100;
assign v376f504 = hmaster2_p & v3a69b74 | !hmaster2_p & v372de3b;
assign v3a6a4cf = hbusreq2 & v373d0af | !hbusreq2 & v37731c3;
assign v3a5d45c = hlock5_p & v37237a8 | !hlock5_p & v3a652b6;
assign v3a7155b = hmaster2_p & v372f309 | !hmaster2_p & v375b2e2;
assign v374853c = hbusreq0 & v3a70a03 | !hbusreq0 & v3a709ec;
assign v3760309 = hbusreq0 & v373a47e | !hbusreq0 & v1e37cd6;
assign v3a6f07b = hmaster1_p & v3736ef2 | !hmaster1_p & v37377d2;
assign v376b504 = hbusreq7 & v3a6177b | !hbusreq7 & v372f520;
assign v37368d3 = hlock0_p & v8455e7 | !hlock0_p & !v3744710;
assign v374648b = stateG10_1_p & v3a70c07 | !stateG10_1_p & v1e37d3f;
assign v37391ac = hmaster2_p & v1e377ba | !hmaster2_p & v3728e58;
assign v3a70be4 = hmaster1_p & v3a6826d | !hmaster1_p & v3748d55;
assign v3a707a7 = hmaster0_p & v374650c | !hmaster0_p & v376d312;
assign v3a6b49a = hgrant7_p & v8455ab | !hgrant7_p & v3a65a2e;
assign v372f8af = hgrant5_p & v3a710bf | !hgrant5_p & v3a6e37f;
assign v3731aac = hmaster0_p & v3a57046 | !hmaster0_p & v3a6fe9a;
assign v376c4c5 = hgrant2_p & v8455ab | !hgrant2_p & v37507da;
assign v3741240 = hbusreq4_p & v3a6fa86 | !hbusreq4_p & v3809240;
assign v37609d7 = hbusreq4_p & v374e7c5 | !hbusreq4_p & v3a58732;
assign v375f3f0 = hlock0_p & v376f73c | !hlock0_p & !v3732e1b;
assign v3a6471a = hbusreq8 & v377800b | !hbusreq8 & v3a70555;
assign v3a71685 = hbusreq6_p & v3a709a4 | !hbusreq6_p & !v8455ab;
assign v3743dc4 = hmaster1_p & v3807f45 | !hmaster1_p & v3a71405;
assign v3755ad0 = hmaster1_p & v377aae4 | !hmaster1_p & v373cada;
assign v3767fa5 = hgrant3_p & v8455ab | !hgrant3_p & v3779fbd;
assign v3a708a9 = hgrant4_p & v37758ad | !hgrant4_p & v377bc9c;
assign v3755289 = hmaster2_p & v373b02e | !hmaster2_p & v377d1dc;
assign v3764005 = hmaster1_p & v373bee7 | !hmaster1_p & v37630ff;
assign v3727d4c = hbusreq5_p & v372c6c4 | !hbusreq5_p & !v8455ab;
assign v3730d77 = hlock7_p & v3734f60 | !hlock7_p & v375ed19;
assign v3a5c983 = hmaster2_p & v3779680 | !hmaster2_p & v3767cc9;
assign v3a68a30 = hgrant0_p & v37773a9 | !hgrant0_p & v3a5979e;
assign v3766487 = hbusreq0 & v37507dd | !hbusreq0 & v374b340;
assign v372ed93 = hmaster0_p & v37443e0 | !hmaster0_p & v8455ab;
assign v374262d = hgrant3_p & v377b6ce | !hgrant3_p & v373a1f2;
assign v375c7f8 = hbusreq3 & v37738fc | !hbusreq3 & v35b774b;
assign v3a710b7 = hbusreq2 & v3760ab8 | !hbusreq2 & v8455bf;
assign v3a5f5f5 = hlock5_p & v3723ac4 | !hlock5_p & !v373b717;
assign v374fef0 = jx0_p & v3777bf4 | !jx0_p & v3a6fa10;
assign v3775a9f = hbusreq5 & d0e017 | !hbusreq5 & v3769740;
assign v3a70b3b = hmaster0_p & baec07 | !hmaster0_p & v3a706e1;
assign v375eb9c = stateG2_p & v8455ab | !stateG2_p & v37386f2;
assign v376a254 = hmaster2_p & v3a6f541 | !hmaster2_p & v3731fd8;
assign v3a5cb9d = hmaster1_p & v374948b | !hmaster1_p & v373e055;
assign v3a53709 = hbusreq7_p & v3a716a4 | !hbusreq7_p & v37756f8;
assign v377e60e = hlock6_p & v3732415 | !hlock6_p & v3a5e7fe;
assign v3741069 = hbusreq4 & v374f307 | !hbusreq4 & v8455b0;
assign v3a662fe = hbusreq6_p & v375156a | !hbusreq6_p & v3a6eeff;
assign v3745ece = hmaster2_p & v3723430 | !hmaster2_p & v376f2f8;
assign v3a65d01 = hbusreq2_p & v3747302 | !hbusreq2_p & v3a70a88;
assign v3a6ecd9 = hbusreq6_p & v3a5e95a | !hbusreq6_p & v3a6c066;
assign v377e9aa = hgrant2_p & v3752a0d | !hgrant2_p & v374e3c2;
assign v3a6ddd4 = hbusreq2 & v375d689 | !hbusreq2 & v3762502;
assign v3a6f83c = hgrant2_p & v8455ab | !hgrant2_p & v3a598b7;
assign v374fa21 = hgrant6_p & v372a20f | !hgrant6_p & v3a6f8f9;
assign v3a6db1a = hgrant6_p & v8455ab | !hgrant6_p & v373a349;
assign v3a71133 = hbusreq4_p & v8455cb | !hbusreq4_p & v3a6c2a9;
assign v3a689d1 = hbusreq7 & v374e74c | !hbusreq7 & v8455ab;
assign v375b801 = hmaster1_p & v376784b | !hmaster1_p & v23fd89c;
assign v3778aa6 = hmaster0_p & v37504f9 | !hmaster0_p & v377926d;
assign v372aacf = hmaster2_p & v3a68084 | !hmaster2_p & v375bb92;
assign v3a6f105 = hbusreq4 & v3a64056 | !hbusreq4 & v37771ca;
assign v3734788 = hbusreq4_p & v3726d1f | !hbusreq4_p & v377f401;
assign v3747994 = hlock0_p & v3a660f2 | !hlock0_p & v3775557;
assign v3726a8d = jx0_p & v8455ab | !jx0_p & v37571d0;
assign v37239ed = hlock4 & v3736cb8 | !hlock4 & v3753bb2;
assign v3743879 = hlock6_p & v3a617b4 | !hlock6_p & v3767437;
assign v374d781 = hlock5_p & v3a6fcb2 | !hlock5_p & v3a55aa3;
assign v375b7b5 = hbusreq2_p & v377eaf2 | !hbusreq2_p & v3a6006a;
assign c7658c = hbusreq5 & v3a580ca | !hbusreq5 & !v8455b9;
assign v3774314 = hbusreq7 & v3725a39 | !hbusreq7 & v3a67fd0;
assign v3757da6 = hbusreq4_p & v37386da | !hbusreq4_p & v3a63d55;
assign v39ebb74 = hgrant6_p & v3a69ae7 | !hgrant6_p & v373e6f1;
assign v37609a6 = hgrant2_p & v3a6f43e | !hgrant2_p & v3756ca5;
assign v374b70d = hlock0_p & v3a299d4 | !hlock0_p & v8455b0;
assign v374ad44 = hbusreq4_p & v3a70c9b | !hbusreq4_p & v37740ec;
assign v3770dcb = hgrant2_p & v3a646f5 | !hgrant2_p & v3772117;
assign v3745b52 = start_p & v8455ab | !start_p & v3730383;
assign v37783d2 = hbusreq8 & v3a701f7 | !hbusreq8 & v377386a;
assign v3a6ebee = hbusreq8 & v37751b4 | !hbusreq8 & v3734e70;
assign v376e587 = hbusreq8_p & v3763c1f | !hbusreq8_p & v3a6f8cf;
assign v37699c9 = hgrant3_p & v360d1cb | !hgrant3_p & v3a66e5d;
assign v3a6fa9a = hmaster2_p & v377234d | !hmaster2_p & v3730a3d;
assign v3a5bd48 = hbusreq1_p & v3a70316 | !hbusreq1_p & v8455b0;
assign v373c4c2 = hbusreq6_p & v3755dcd | !hbusreq6_p & !v3729421;
assign v3742623 = hmaster0_p & v37403ef | !hmaster0_p & v375c76b;
assign v377a345 = hgrant3_p & v35b7299 | !hgrant3_p & !v3a70524;
assign v3a63f0c = hbusreq4_p & v3a656b6 | !hbusreq4_p & v3726b10;
assign v374f76a = hlock0_p & v3747302 | !hlock0_p & v3748481;
assign v372bd06 = hmaster2_p & v3a56b60 | !hmaster2_p & v37427e9;
assign v377a308 = hmaster3_p & v360d099 | !hmaster3_p & v3a660a5;
assign v377619b = hmaster1_p & v3a635ea | !hmaster1_p & v3a5b109;
assign v3a7067d = hgrant5_p & v8455ab | !hgrant5_p & v373195f;
assign v3a6eaef = hmaster0_p & v3a71561 | !hmaster0_p & !v3a5f4b8;
assign v375b0d5 = hbusreq4_p & v3a62826 | !hbusreq4_p & v35b774b;
assign v376b164 = stateG2_p & v8455ab | !stateG2_p & v3759020;
assign v3a60cbd = hbusreq6 & v92acd8 | !hbusreq6 & v8455ab;
assign v3a63621 = stateA1_p & v3a635ea | !stateA1_p & !v35772a5;
assign v3a55c2f = hmaster0_p & v3a70d99 | !hmaster0_p & v9af5fc;
assign v375c9f0 = hbusreq4_p & v3752536 | !hbusreq4_p & !v8455ab;
assign v377b096 = hmaster2_p & v376489b | !hmaster2_p & v376d1bb;
assign v3a68276 = hbusreq2 & v3a5600a | !hbusreq2 & v8455ab;
assign v3747fa9 = hbusreq0 & v3a6d500 | !hbusreq0 & v3a5d2bc;
assign v3a6f000 = hmaster2_p & v3732dc6 | !hmaster2_p & v8455ab;
assign v37665e2 = hbusreq4_p & v372b24d | !hbusreq4_p & v3a709ea;
assign v3760eb3 = hbusreq4_p & v3a667b8 | !hbusreq4_p & v8455ab;
assign v3a65526 = hbusreq4 & v3a6b916 | !hbusreq4 & v3768c3e;
assign v372a823 = hbusreq0 & v3a65368 | !hbusreq0 & v372ba45;
assign v3752913 = hbusreq5_p & v3736ea9 | !hbusreq5_p & v8455ab;
assign v373f2fe = hbusreq8 & v3a70fea | !hbusreq8 & v3a71146;
assign v3a70ef8 = hmaster2_p & v3a635ea | !hmaster2_p & v37450b8;
assign v3a7074c = hgrant5_p & v3807587 | !hgrant5_p & v3a70be4;
assign v3a7012f = hlock4_p & v37604e9 | !hlock4_p & v35772a6;
assign v3a68834 = hbusreq6_p & v3a67983 | !hbusreq6_p & v377eb9d;
assign v373aa3d = hgrant4_p & v8455ab | !hgrant4_p & v357733c;
assign v37355ea = hmaster2_p & v375139d | !hmaster2_p & v3766ff7;
assign v37273b1 = hmaster2_p & v376501e | !hmaster2_p & v377234d;
assign v3a6ff35 = hmaster2_p & v377d7dc | !hmaster2_p & v3a6f0f9;
assign v377eac3 = hmaster1_p & v3a70209 | !hmaster1_p & v376a755;
assign v3a5ef2e = hbusreq7_p & v3a7042c | !hbusreq7_p & v3723d1a;
assign v3a6ef5f = hbusreq3_p & v376e040 | !hbusreq3_p & v3a6051a;
assign v3a621e6 = hmaster3_p & v376dae8 | !hmaster3_p & v3734a96;
assign v37727be = hgrant1_p & v374721d | !hgrant1_p & v8455ab;
assign v376bae4 = hmaster2_p & v3755e23 | !hmaster2_p & !v3a6ffe1;
assign v37267a5 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3809487;
assign v8455be = hbusreq3 & v8455ab | !hbusreq3 & !v8455ab;
assign v372bb35 = hbusreq7 & v3a70e80 | !hbusreq7 & v8455ab;
assign v37415ea = jx0_p & v3a70a44 | !jx0_p & v8455ab;
assign v37709bb = hgrant2_p & v376004c | !hgrant2_p & v374c718;
assign v3a607bd = hmaster1_p & v376a84d | !hmaster1_p & v3a573c2;
assign v377b2e1 = hmaster2_p & v3a5af28 | !hmaster2_p & v3748d67;
assign v3a6e986 = hmaster0_p & v3a54e41 | !hmaster0_p & !v3752b8f;
assign v3768502 = hbusreq8 & v3a56197 | !hbusreq8 & v3a6fb21;
assign v3a5e1e4 = hmaster0_p & v373a27c | !hmaster0_p & v3a61c51;
assign v373ac65 = hmaster1_p & v3a6fa11 | !hmaster1_p & v37435e9;
assign v372c492 = hlock7 & v35b7033 | !hlock7 & v373edf3;
assign v3755539 = hmaster2_p & v374da61 | !hmaster2_p & v3a5d5a4;
assign v3a65e1e = hgrant6_p & v374a664 | !hgrant6_p & v375e9a7;
assign v37476f7 = hgrant6_p & v3741b28 | !hgrant6_p & v3741cda;
assign v3a68356 = hmaster0_p & v3766746 | !hmaster0_p & v8455ab;
assign v3a569c8 = hbusreq5_p & v3a6b090 | !hbusreq5_p & v3a708fb;
assign v376d5a7 = hbusreq4_p & v8455b0 | !hbusreq4_p & v3753dab;
assign v3a6fb8f = hmaster1_p & v37682ce | !hmaster1_p & !v3a6fd84;
assign v374c0e4 = hgrant6_p & v8455ab | !hgrant6_p & v3766218;
assign v3a5c9d7 = hmaster2_p & v3753418 | !hmaster2_p & v3767b70;
assign v3a6aa9e = hgrant5_p & v8455ab | !hgrant5_p & v37536bf;
assign v865472 = stateG3_2_p & v8455ab | !stateG3_2_p & v37603af;
assign v3729115 = hbusreq3_p & v3732b81 | !hbusreq3_p & v3759947;
assign v3779071 = hmaster0_p & v3a6fb65 | !hmaster0_p & v374e6b1;
assign ce3eb4 = jx2_p & v3741b5a | !jx2_p & v3739c9a;
assign v375bf96 = hgrant4_p & v3a708d3 | !hgrant4_p & v3a68c0e;
assign v374bb02 = hbusreq2 & v372efbe | !hbusreq2 & v8455ab;
assign v3743f11 = hbusreq3_p & v377eaf2 | !hbusreq3_p & v3735512;
assign v373abcf = hmaster1_p & v3a635ea | !hmaster1_p & v3760bda;
assign v3a6eb83 = hbusreq3 & v8455b0 | !hbusreq3 & v37406d2;
assign v3733228 = hmaster0_p & v374743d | !hmaster0_p & v37599eb;
assign v3a6c3ae = hmaster1_p & v3a6810b | !hmaster1_p & v8455e7;
assign v3809b31 = hbusreq3_p & v3766877 | !hbusreq3_p & v3a68d2e;
assign v3a59613 = jx0_p & v8455ab | !jx0_p & v3a6f863;
assign v3a70f7c = hmaster3_p & v3a54484 | !hmaster3_p & v8455ab;
assign v3a6f53d = hbusreq3_p & v373d025 | !hbusreq3_p & !v3725f77;
assign v37472ea = hgrant5_p & v3733886 | !hgrant5_p & v37585bd;
assign v376956a = hbusreq8 & v3a5f205 | !hbusreq8 & v3745d1e;
assign v374494b = jx1_p & v3a70471 | !jx1_p & v3a70dc3;
assign cc2c2e = hbusreq2 & v3729d1a | !hbusreq2 & !v8455ab;
assign v23fdf1a = hmaster2_p & v3731b41 | !hmaster2_p & v3a700d8;
assign v3750857 = hlock7 & v372c20d | !hlock7 & v3a706ea;
assign v374845f = hmaster1_p & v375766c | !hmaster1_p & v377195f;
assign v3a71098 = hbusreq2_p & v3a66668 | !hbusreq2_p & v373a984;
assign v3723477 = hmaster2_p & v3740161 | !hmaster2_p & v3a5c30f;
assign v3747cdb = hgrant0_p & v3577306 | !hgrant0_p & v3740152;
assign v37551ac = hmaster0_p & v3778a5a | !hmaster0_p & v377a985;
assign v3756954 = hmaster2_p & v8455e7 | !hmaster2_p & v3a676d6;
assign v372b715 = hmaster3_p & v3a712a6 | !hmaster3_p & v375041a;
assign v3a6f1fd = hbusreq0_p & v3a635ea | !hbusreq0_p & v376bade;
assign v375eaea = hbusreq5 & v3806575 | !hbusreq5 & v3a5aad8;
assign v3a70394 = hbusreq2_p & v37403e5 | !hbusreq2_p & v8455ab;
assign v376a40d = hmaster2_p & v377d142 | !hmaster2_p & v3741f4b;
assign v377e9d7 = hlock0 & v37285eb | !hlock0 & v37264c9;
assign v3a70e4c = hlock5 & v3a6a02a | !hlock5 & v3730778;
assign v376c5f5 = hgrant6_p & v3a2a8f2 | !hgrant6_p & v374bec6;
assign v3a6f212 = hmaster3_p & v3a635ea | !hmaster3_p & v3751141;
assign v373d9e5 = stateA1_p & v8455ab | !stateA1_p & !v37481c3;
assign v373f262 = hbusreq7_p & c08050 | !hbusreq7_p & v374f645;
assign afa7f5 = hbusreq4 & v3a6dc08 | !hbusreq4 & v37406d2;
assign v3777daa = hbusreq4 & cff2df | !hbusreq4 & v3a70a7f;
assign v8455c1 = hbusreq4_p & v8455ab | !hbusreq4_p & !v8455ab;
assign v374cd51 = hgrant4_p & v8455ab | !hgrant4_p & v376455c;
assign v37458a3 = hgrant2_p & v375c7b9 | !hgrant2_p & v377022e;
assign v374d255 = hmaster0_p & v3a635ea | !hmaster0_p & v374d2d5;
assign v375b22c = hbusreq8 & v3771a24 | !hbusreq8 & v8455ab;
assign v3a71399 = hmaster0_p & v375b429 | !hmaster0_p & v377d142;
assign v3a703fc = hbusreq2_p & v39a5265 | !hbusreq2_p & v8455e1;
assign v372529a = hmaster2_p & cea55f | !hmaster2_p & v375c351;
assign v3744314 = hmaster2_p & v3a5e24e | !hmaster2_p & v1e38275;
assign v3a6f8c5 = hmaster3_p & v376b1aa | !hmaster3_p & v3a713c0;
assign v373f7a5 = hmaster2_p & v3a69c98 | !hmaster2_p & v375a3dc;
assign v3a65562 = hbusreq6 & v3a6bc65 | !hbusreq6 & v8455b9;
assign v373270f = hbusreq4_p & v377349f | !hbusreq4_p & v375f1ee;
assign v3759fca = hlock4_p & v3a637dd | !hlock4_p & !v8455ab;
assign v373e60c = hlock5 & v3747c20 | !hlock5 & v374b42b;
assign v3a70a00 = hbusreq5 & v3776150 | !hbusreq5 & v8455ab;
assign v377ea72 = hbusreq4_p & v372493b | !hbusreq4_p & !v3a6febd;
assign v373520f = hmaster0_p & v376285a | !hmaster0_p & v3a659eb;
assign v374748f = hbusreq4 & v3a6f04c | !hbusreq4 & v3a5f9e6;
assign v3a602c3 = hbusreq4_p & v37293d5 | !hbusreq4_p & v3a715ca;
assign v3379035 = hlock2_p & v3a6eb39 | !hlock2_p & v35772a6;
assign v3772e85 = hmaster0_p & v3a635ea | !hmaster0_p & v3a54580;
assign v3729b48 = hlock0 & v373bd6c | !hlock0 & v377419a;
assign v376ef42 = locked_p & v8455ab | !locked_p & v3a70c07;
assign v372630c = hmaster0_p & v377ecf0 | !hmaster0_p & v3a57e58;
assign v376a2e7 = hmaster3_p & v3a67fb5 | !hmaster3_p & v376b1ee;
assign v3765590 = hmaster1_p & v373ce86 | !hmaster1_p & v3a58139;
assign v3732c24 = hbusreq2 & v37379bb | !hbusreq2 & !v3736ebd;
assign v3729531 = hbusreq6 & v3733727 | !hbusreq6 & v3748797;
assign v3a5f43a = hmaster2_p & v374297b | !hmaster2_p & v3a6ce39;
assign v37485ec = hgrant2_p & v8455e7 | !hgrant2_p & !v3a70394;
assign v37316f3 = hmaster1_p & v8455b9 | !hmaster1_p & v3757301;
assign v3726ed7 = hmaster1_p & v3751e0a | !hmaster1_p & v3a6fbaf;
assign v3772f26 = hgrant6_p & v377938d | !hgrant6_p & v3a6ff5c;
assign v3771502 = hgrant5_p & v37431ac | !hgrant5_p & ad187c;
assign v377a60f = hbusreq5 & v374d59d | !hbusreq5 & v3774bad;
assign v37526e0 = hgrant1_p & v376e139 | !hgrant1_p & v3735ed0;
assign v375f60e = hbusreq7_p & v3766b23 | !hbusreq7_p & v372de8f;
assign v3a6f2dc = hmaster0_p & v375159d | !hmaster0_p & v3777817;
assign v3a6ddb3 = hbusreq8 & v3735ad0 | !hbusreq8 & v8455ab;
assign v3779f6b = hbusreq6_p & v3a586f1 | !hbusreq6_p & v8455ab;
assign v373c6b6 = hmaster2_p & v3a6be44 | !hmaster2_p & !v8455ab;
assign v3765734 = hbusreq7_p & v3757e32 | !hbusreq7_p & v3746444;
assign v39a4ef6 = hmaster2_p & v3750746 | !hmaster2_p & !v8455ab;
assign v372d811 = hmaster1_p & v8455ab | !hmaster1_p & v377077a;
assign v3752002 = hlock4 & v3758a9c | !hlock4 & v372e4de;
assign v3a68ebe = hmaster1_p & v37587a4 | !hmaster1_p & v3a64718;
assign v3a701de = hbusreq5_p & v3a5f066 | !hbusreq5_p & v3a5ec68;
assign v3751383 = hbusreq5 & v3755e61 | !hbusreq5 & v37493b4;
assign v3770bca = hmaster1_p & bb70de | !hmaster1_p & v3769b3f;
assign d5f283 = hbusreq4_p & v3776e9c | !hbusreq4_p & v8455ab;
assign v3a70e3d = hbusreq4 & v375a4fa | !hbusreq4 & v8455ab;
assign v1e38224 = stateA1_p & v8455ab | !stateA1_p & v39a5381;
assign v3a705dd = hbusreq6 & v39eb3bd | !hbusreq6 & v3738df9;
assign v3a70a85 = jx1_p & v376dee4 | !jx1_p & v3a532f2;
assign v3a66c9a = hmaster0_p & v377b015 | !hmaster0_p & v377f6ae;
assign v3a6392b = hlock4_p & v377989c | !hlock4_p & v8455e7;
assign v372cdec = hgrant5_p & v8455ab | !hgrant5_p & !v3a6fd10;
assign v38092e6 = hgrant4_p & v3a656d0 | !hgrant4_p & v3756883;
assign v3774913 = hbusreq3_p & b4444b | !hbusreq3_p & v8455ab;
assign v8ce84c = hbusreq8_p & v3a704b3 | !hbusreq8_p & v3a6f376;
assign v3a7011b = hbusreq7_p & v372543f | !hbusreq7_p & v377d9b2;
assign v374fa56 = hgrant3_p & v8455bd | !hgrant3_p & v3a6fa30;
assign v3756e39 = hmaster0_p & v374a668 | !hmaster0_p & v3770db3;
assign v3809f73 = hbusreq5_p & v3746d31 | !hbusreq5_p & !v377adf5;
assign v3773ba2 = hbusreq0_p & v375e309 | !hbusreq0_p & v8455ab;
assign v3773b7b = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a6e91d;
assign v3a6caa5 = hbusreq4_p & v3750d37 | !hbusreq4_p & !v3732dc6;
assign b6a7cc = hmaster0_p & v3769101 | !hmaster0_p & v8455ab;
assign v3a70f9c = hmaster2_p & v374cb9e | !hmaster2_p & v3a5d134;
assign v37720ca = hgrant3_p & v377057a | !hgrant3_p & v37455ec;
assign v38087e5 = hmaster0_p & v3723185 | !hmaster0_p & v37270b9;
assign v3725a6e = hgrant5_p & v3a578ef | !hgrant5_p & v376a556;
assign v374831d = jx0_p & v37470a5 | !jx0_p & !v3a594e8;
assign v3a7016b = hmaster0_p & v377ca40 | !hmaster0_p & v3a71609;
assign v3a672e5 = hbusreq4_p & v3a5faba | !hbusreq4_p & v3a6e089;
assign v373ec8e = hgrant6_p & v8455ab | !hgrant6_p & v1e379e9;
assign v37455ff = hmaster2_p & v377ca49 | !hmaster2_p & v373df13;
assign v372e031 = hmaster0_p & v8455b0 | !hmaster0_p & v377c71d;
assign v376cfae = hmaster0_p & v3770a82 | !hmaster0_p & v375449f;
assign v376265d = hmaster0_p & v375b429 | !hmaster0_p & v376a40d;
assign v3730b1c = hgrant5_p & v3a7159f | !hgrant5_p & v375822b;
assign v37345e9 = hlock0_p & v3a70b0d | !hlock0_p & v3765798;
assign v3a6e37f = hmaster1_p & v3a6ffa1 | !hmaster1_p & v3a69ad9;
assign v372fd12 = hbusreq2_p & v372310a | !hbusreq2_p & v3743b9e;
assign v3736dfd = hmaster1_p & v3a5c945 | !hmaster1_p & v374055c;
assign v373da1b = hmaster1_p & v3a696a7 | !hmaster1_p & v37695c7;
assign v376a74a = hbusreq8 & v3765e47 | !hbusreq8 & v8455ab;
assign v3a6cb62 = hbusreq4 & v3a5b4de | !hbusreq4 & v38072fd;
assign v3725d7b = hgrant6_p & v8455ab | !hgrant6_p & v3a6fa49;
assign v3a56e7a = hbusreq6 & v3a6fcc8 | !hbusreq6 & v8455ab;
assign v3a64a83 = hbusreq5 & v3a56eeb | !hbusreq5 & v8455ab;
assign v37770ed = hbusreq6 & v38094fb | !hbusreq6 & !v8455ab;
assign d78807 = hgrant2_p & v3a59bb4 | !hgrant2_p & v37693a9;
assign v3724908 = hbusreq8 & v374d121 | !hbusreq8 & v376673b;
assign v374a3db = hbusreq6_p & v3a6fd47 | !hbusreq6_p & v3a70142;
assign v3746b6e = hbusreq2 & v3730627 | !hbusreq2 & v3a5980d;
assign v38064d5 = hlock5 & v3a70c69 | !hlock5 & v3742303;
assign v3759fda = hlock7_p & v372bda4 | !hlock7_p & !v8455ab;
assign v3a69df1 = hgrant2_p & v3a60787 | !hgrant2_p & v3749380;
assign v375d861 = hbusreq6_p & v375e261 | !hbusreq6_p & v376096f;
assign v3754f2e = hlock4 & v3756c83 | !hlock4 & v373fe6f;
assign v373bbc1 = hmaster0_p & v3a661fe | !hmaster0_p & v99b6f5;
assign v375a86a = hmaster2_p & v37270bc | !hmaster2_p & v373bd76;
assign v37761ae = hbusreq3_p & v3774c1b | !hbusreq3_p & !v38099c1;
assign v3a65368 = hbusreq4 & v3a71319 | !hbusreq4 & v37235f9;
assign v37591ac = hlock0_p & v3a7153a | !hlock0_p & v373cc68;
assign v372ba93 = hmaster2_p & v3753eb2 | !hmaster2_p & v3a65dcf;
assign v3747fbf = hlock7 & v3a69677 | !hlock7 & v3a6f38b;
assign v3725dce = hgrant6_p & v3775b81 | !hgrant6_p & v8455ab;
assign v3a70114 = hbusreq0 & v3a6443d | !hbusreq0 & v3738ff9;
assign v3774b89 = hbusreq2_p & v375641f | !hbusreq2_p & !v3a6b0c7;
assign v373127e = hbusreq6_p & v8455bf | !hbusreq6_p & v3763a20;
assign v3777b2e = hbusreq4_p & v37536ae | !hbusreq4_p & v3a7103a;
assign v37793e4 = hgrant4_p & v3a635ea | !hgrant4_p & v3775f4f;
assign v3a70374 = hgrant4_p & v3747302 | !hgrant4_p & v3726d1f;
assign v377bc8e = hmaster0_p & a9e394 | !hmaster0_p & v3742cd4;
assign v3808c5f = hmaster1_p & v37c073f | !hmaster1_p & v374d7dc;
assign v3a70f29 = hbusreq6_p & v2acb5a2 | !hbusreq6_p & !v8455ab;
assign v3a5ad12 = hbusreq4 & v377b8ee | !hbusreq4 & v8455ab;
assign v3742dac = hmaster2_p & v3a6f6a4 | !hmaster2_p & v3750a9c;
assign v3a6eef8 = hlock8 & v374159f | !hlock8 & v3a710ff;
assign v3a61fd3 = hbusreq2_p & v3729ffd | !hbusreq2_p & v372f72b;
assign v3a62ad8 = hbusreq5_p & v374b362 | !hbusreq5_p & v3756045;
assign v3a6ff27 = hmaster0_p & v39ea76e | !hmaster0_p & v3a714d8;
assign v377b3a8 = hbusreq3 & v37583be | !hbusreq3 & v376b4e1;
assign v3779678 = hbusreq5_p & v372a55a | !hbusreq5_p & !v372d75a;
assign v3735cfb = hmaster0_p & v372d8e8 | !hmaster0_p & v3743113;
assign v373c2d7 = hgrant6_p & v8455ab | !hgrant6_p & v3a62d56;
assign v372ef39 = hmaster0_p & v37762cd | !hmaster0_p & v3a68cec;
assign v373ae22 = hgrant3_p & v3a64643 | !hgrant3_p & !v372f7c6;
assign v3a709aa = hgrant3_p & v3770f46 | !hgrant3_p & d08a74;
assign v3a6750f = hmaster2_p & v3a66110 | !hmaster2_p & !v1e38224;
assign v372b1e6 = hbusreq4_p & v37618ef | !hbusreq4_p & v3a6fc03;
assign v3a65827 = hlock2 & v3a700b0 | !hlock2 & v3747e8e;
assign v3a6f0fd = hlock2 & v375e577 | !hlock2 & b3d3ad;
assign v3a5c064 = hbusreq5_p & v37499a9 | !hbusreq5_p & v377adf7;
assign v3742676 = hbusreq7 & v3a5d8e0 | !hbusreq7 & v3a65afd;
assign v3a5575e = hmaster1_p & v37570f8 | !hmaster1_p & v3a65e6a;
assign v377dc99 = hmaster1_p & v3a5fc34 | !hmaster1_p & v3770ff9;
assign v3a574fc = hbusreq5_p & v3a70478 | !hbusreq5_p & v377a62e;
assign v3a70e8d = hgrant2_p & v3a70645 | !hgrant2_p & v377b086;
assign v377c47c = jx0_p & v37795a3 | !jx0_p & v375ae8d;
assign v3a705a6 = hgrant4_p & v3749b09 | !hgrant4_p & v37652eb;
assign v3a69b93 = hlock4 & v3a5f83c | !hlock4 & v3763d77;
assign v37662dc = hbusreq3_p & v3809adf | !hbusreq3_p & !v3a70c07;
assign v3a70c92 = hlock5 & v3762e54 | !hlock5 & v3755113;
assign v3a70d41 = hbusreq7_p & v3777f6f | !hbusreq7_p & v3a6f410;
assign v3a70948 = hbusreq0 & v37793c8 | !hbusreq0 & v373d41a;
assign v374d6dd = hlock4_p & v3a68426 | !hlock4_p & v8455b7;
assign v37379d7 = hbusreq2 & v372600f | !hbusreq2 & bf3e2b;
assign v3a712c8 = hmaster2_p & v373be25 | !hmaster2_p & v3a6b0c7;
assign v3746dd5 = hbusreq2_p & v3a57f59 | !hbusreq2_p & !v3a66110;
assign v375bb06 = hmaster1_p & v3a6ebd2 | !hmaster1_p & v374ec57;
assign v3a6f994 = hgrant6_p & v8455ab | !hgrant6_p & v1e37413;
assign v3a7047d = hmaster1_p & v3a703b0 | !hmaster1_p & v3a67555;
assign v9e6ddd = hbusreq5_p & v372b5bc | !hbusreq5_p & v3a6fe91;
assign v374c556 = jx0_p & v861ce0 | !jx0_p & v375c2d0;
assign v374760a = hbusreq6 & v3a6dc08 | !hbusreq6 & v8455b0;
assign v373a4cd = hbusreq5 & v37373bb | !hbusreq5 & v374e4fa;
assign v3a709a3 = hbusreq6_p & c61b3c | !hbusreq6_p & !v8455ab;
assign v37263bf = hbusreq5_p & v3736421 | !hbusreq5_p & v3767638;
assign v3a705bd = hbusreq8 & v373a59e | !hbusreq8 & v37285cd;
assign v3a6513d = hmaster0_p & v3736e19 | !hmaster0_p & v3a7094f;
assign v3a7121e = hmaster1_p & v3a5e24e | !hmaster1_p & v3758c5c;
assign d58c24 = hmaster2_p & v35b774b | !hmaster2_p & v8455ab;
assign v3a5d930 = hmaster3_p & v3a6f7eb | !hmaster3_p & v3a66988;
assign v37593c6 = hmaster1_p & v3763f95 | !hmaster1_p & v3728d1d;
assign v3a6e0ab = hgrant5_p & v3741566 | !hgrant5_p & v376277f;
assign v39eaa60 = hmaster0_p & v37bfc35 | !hmaster0_p & v37799ca;
assign v3a704a7 = hgrant5_p & v3744f6f | !hgrant5_p & v37482da;
assign v377e2f1 = stateG10_1_p & v3740171 | !stateG10_1_p & v3768c21;
assign v3a6f6ec = hmaster2_p & v3a6f995 | !hmaster2_p & v373a629;
assign v3a5aa3a = hbusreq4_p & v3739892 | !hbusreq4_p & v3a714e4;
assign v3a6f35b = hmaster2_p & v3a6f97b | !hmaster2_p & v3760513;
assign v376a4ec = hlock5 & v37581cf | !hlock5 & v372c3c7;
assign v3736679 = hbusreq0_p & v3a676d6 | !hbusreq0_p & v8455ab;
assign v37511c0 = hbusreq2_p & v372ff2c | !hbusreq2_p & v3a699d3;
assign v3a5b7e7 = hbusreq4_p & v3a701a0 | !hbusreq4_p & v3808c66;
assign v3749dc1 = hmaster0_p & v3759007 | !hmaster0_p & v3770fef;
assign v3768d1d = hbusreq8_p & v375d3e2 | !hbusreq8_p & v376cf03;
assign v3a7149e = hbusreq4 & v3736a23 | !hbusreq4 & v8455ab;
assign v375c7cd = hbusreq5_p & v3752e29 | !hbusreq5_p & v8455ab;
assign v3a6f794 = hgrant5_p & v1e37b48 | !hgrant5_p & v3735bef;
assign v375fc79 = jx0_p & v3766dfb | !jx0_p & v3a6fee5;
assign v373d5d6 = hlock3 & v375899b | !hlock3 & v374ec84;
assign v3766035 = hgrant1_p & v3a5dbb7 | !hgrant1_p & v3735ed0;
assign v3774d12 = hbusreq4_p & v3a66999 | !hbusreq4_p & cbb40b;
assign v376d4cb = hlock5_p & v3a68426 | !hlock5_p & v8455b7;
assign v37479ef = hbusreq4_p & v37427f8 | !hbusreq4_p & !v8455c2;
assign v3771724 = hlock7_p & v3a707e8 | !hlock7_p & v3771319;
assign v376d640 = hmaster0_p & v373f911 | !hmaster0_p & v373665b;
assign v3767feb = hgrant3_p & v8455be | !hgrant3_p & v3a70c11;
assign v37c007b = hbusreq4 & v37482f8 | !hbusreq4 & v8455ab;
assign v375b12b = hbusreq5_p & v3762873 | !hbusreq5_p & v3a71105;
assign v374e6c7 = hmaster2_p & v375cf36 | !hmaster2_p & v372e83f;
assign v37767fa = hmaster2_p & v2ff8c74 | !hmaster2_p & v3a70147;
assign v376021d = hmaster0_p & v372ff0a | !hmaster0_p & v374ebb6;
assign v372f38e = hmaster2_p & v374be5d | !hmaster2_p & v3728d9c;
assign v377d59e = hmaster1_p & v37475d9 | !hmaster1_p & v37695f7;
assign v3a5f717 = hgrant5_p & v3a56130 | !hgrant5_p & !v8455ab;
assign v3a7104e = hmaster0_p & v3a702d9 | !hmaster0_p & v3748179;
assign v3a65e9a = hgrant4_p & v3752a0d | !hgrant4_p & v3751719;
assign v3745a81 = hbusreq4 & v3a67b48 | !hbusreq4 & v3a685c7;
assign v3a6fd6a = hlock6 & v3a70bf1 | !hlock6 & v376e04c;
assign v37565a0 = hgrant2_p & v3764276 | !hgrant2_p & v3a713dc;
assign v372ae6f = hmaster2_p & v3a6f59d | !hmaster2_p & !v3744f62;
assign v3755914 = hmaster2_p & v374820d | !hmaster2_p & v23fdeaf;
assign v3a67261 = hlock2_p & v3735eb8 | !hlock2_p & v8455b3;
assign v376f051 = hbusreq5_p & v374a8bb | !hbusreq5_p & v37533f6;
assign v377c236 = hmaster1_p & v375c791 | !hmaster1_p & v3754d28;
assign v3766c68 = hmaster0_p & v8455ab | !hmaster0_p & !v377278b;
assign v372b304 = hbusreq2 & v372e305 | !hbusreq2 & v3379037;
assign v375b98c = hbusreq6_p & b66740 | !hbusreq6_p & !v2092faa;
assign v3753ff9 = hgrant3_p & v37579a9 | !hgrant3_p & v3765b08;
assign v372d5bb = hgrant2_p & v375d38f | !hgrant2_p & !v3a6feb9;
assign v3747238 = hmaster2_p & v8455ab | !hmaster2_p & v3a6f9d7;
assign v3768e79 = hgrant4_p & v3a7133d | !hgrant4_p & v372cd91;
assign v372f765 = hbusreq8 & v375aea8 | !hbusreq8 & v8455ab;
assign v376f271 = hmaster1_p & v3a6d874 | !hmaster1_p & !v377f640;
assign v373d7fe = hgrant0_p & v37773a9 | !hgrant0_p & v3723ac5;
assign v3a635ff = hbusreq1_p & v3763cf5 | !hbusreq1_p & !v37519ed;
assign v3a5e95a = hbusreq6 & v3749435 | !hbusreq6 & v8455ab;
assign v374b116 = hmaster2_p & v376b88d | !hmaster2_p & v3752e63;
assign v23fd970 = stateA1_p & v8455ab | !stateA1_p & !v3a6fa4f;
assign v3745b4f = hlock3_p & v372abd8 | !hlock3_p & v35772a6;
assign v3735cb2 = hmaster1_p & v3a6f556 | !hmaster1_p & !v3738826;
assign v3773bc6 = hbusreq6_p & v3a71558 | !hbusreq6_p & v3764bca;
assign v3a5ad94 = hgrant3_p & v377536e | !hgrant3_p & v8455ab;
assign v37658f5 = hgrant2_p & v8455ab | !hgrant2_p & v3770be3;
assign v3a6f310 = hbusreq0 & v3744f86 | !hbusreq0 & v8455ab;
assign v3741833 = hbusreq2_p & v372673b | !hbusreq2_p & v3742d37;
assign v372e6ad = hbusreq1 & v37583be | !hbusreq1 & v376b4e1;
assign v37419ca = hmaster2_p & v3a70147 | !hmaster2_p & v3775e81;
assign v3754229 = hgrant6_p & v3a57fff | !hgrant6_p & v37461e1;
assign v3728906 = hmaster0_p & v8455e7 | !hmaster0_p & v3a6fae3;
assign v37618bf = hmaster2_p & v3a57384 | !hmaster2_p & v3a641d5;
assign v373917f = jx1_p & v374b237 | !jx1_p & !v373cc0c;
assign v3a684bb = hgrant4_p & v8455ab | !hgrant4_p & v3a66123;
assign v3779008 = hlock4 & v3a71197 | !hlock4 & v3742b84;
assign v3a5cd0e = hmaster3_p & v8455ab | !hmaster3_p & v3a6f7db;
assign v372ce29 = hbusreq5_p & v3a707e0 | !hbusreq5_p & v3a61a2d;
assign v37621e0 = hmaster2_p & v373ad95 | !hmaster2_p & !v3a6b873;
assign v375f862 = jx1_p & v3769a2a | !jx1_p & v3a6fc1a;
assign v374122a = hbusreq5_p & v3a6eec4 | !hbusreq5_p & v3a70f1d;
assign v3752862 = hgrant6_p & v3a7156d | !hgrant6_p & v3a6fe3e;
assign v372bccc = jx1_p & v372de49 | !jx1_p & v37751ae;
assign v3748ba9 = hmaster0_p & v37793e4 | !hmaster0_p & v3a705d5;
assign v375ac09 = hmaster0_p & v37240a4 | !hmaster0_p & v377e51b;
assign v377709a = hmaster0_p & v375d76b | !hmaster0_p & !v37470e2;
assign v37699ec = jx1_p & v9d97fe | !jx1_p & v3771da0;
assign v3743b79 = hgrant2_p & v3a632f4 | !hgrant2_p & v3743f47;
assign v3748e09 = hlock5 & v37553f5 | !hlock5 & v3a6087b;
assign v374fc3b = hbusreq5 & bb0568 | !hbusreq5 & v8455ab;
assign v3723542 = hbusreq2_p & v372c60a | !hbusreq2_p & v3773982;
assign v3a5d8f6 = hmaster3_p & v3a70ae5 | !hmaster3_p & v3a715f8;
assign v372b12d = hmaster0_p & v375eee3 | !hmaster0_p & v3a71374;
assign v3a7126a = hbusreq1_p & v376dc2e | !hbusreq1_p & v3774494;
assign v3744f52 = hbusreq3 & v37479b4 | !hbusreq3 & v372b5b0;
assign v372e8ff = hmaster2_p & v3754fb0 | !hmaster2_p & v373ae1e;
assign v3751238 = hbusreq4 & v3379037 | !hbusreq4 & v8455ab;
assign v3a6f426 = hmaster0_p & v3a67d66 | !hmaster0_p & v374430e;
assign v3a71614 = hmaster2_p & a26159 | !hmaster2_p & v3a65e9a;
assign v377d232 = hgrant4_p & v1e37b99 | !hgrant4_p & !v3a7106d;
assign v372be5d = hbusreq5_p & v376e5b6 | !hbusreq5_p & v3808d7d;
assign v3740663 = hmaster1_p & v3a6870f | !hmaster1_p & v375ecab;
assign v3a70ad5 = jx0_p & v37531ca | !jx0_p & v37423c1;
assign v374b07c = hbusreq4 & v37566b2 | !hbusreq4 & !v8455ab;
assign v373afd5 = hbusreq5_p & v3756beb | !hbusreq5_p & v373274f;
assign v373c830 = hbusreq2 & v37583be | !hbusreq2 & !v8455ab;
assign v3748f17 = hgrant6_p & v8455c9 | !hgrant6_p & v33790e4;
assign v3a71019 = hlock6_p & v3730e98 | !hlock6_p & v3a63805;
assign v37502ca = hlock0 & v3731230 | !hlock0 & v3a6d4bf;
assign v3a70656 = hmaster1_p & v3743ff2 | !hmaster1_p & v3736f36;
assign v3a296d3 = hbusreq7 & v372f23a | !hbusreq7 & v8455bb;
assign v3a702cb = hlock0 & v3a60a68 | !hlock0 & v3a5f4b1;
assign v3a5bccf = hbusreq4_p & v3a70326 | !hbusreq4_p & v3766bc8;
assign v3776066 = hgrant5_p & a740cc | !hgrant5_p & v37630a8;
assign v376ff46 = hmaster0_p & v3a6c4e4 | !hmaster0_p & v37581a6;
assign v375d42d = hmaster2_p & v376b908 | !hmaster2_p & v3731737;
assign v3751fde = jx1_p & v866387 | !jx1_p & !v375e147;
assign v377dfec = hbusreq4 & v3760f4e | !hbusreq4 & v8455b3;
assign v3a5d469 = hbusreq0_p & v3a6f7bf | !hbusreq0_p & v8455ab;
assign v374cf44 = jx0_p & v374c885 | !jx0_p & v372ff79;
assign v375f2ba = hgrant4_p & v3a70b17 | !hgrant4_p & v3746ffa;
assign v3772c9f = hmaster0_p & v375cb5e | !hmaster0_p & !v3725496;
assign v3734916 = hgrant4_p & v3807afa | !hgrant4_p & v374fe39;
assign v3730878 = hmaster2_p & v37386f5 | !hmaster2_p & v3a71416;
assign v373c428 = hbusreq1_p & v37663a2 | !hbusreq1_p & v376cf85;
assign v3742f76 = hlock5 & v37410dc | !hlock5 & v3a63306;
assign v37533d5 = hgrant1_p & v377b159 | !hgrant1_p & v8455ab;
assign v3731508 = hmaster0_p & v3745cc6 | !hmaster0_p & v3a70f68;
assign v3a6ae54 = jx0_p & v3a29844 | !jx0_p & v23fd9fe;
assign v3a70d36 = hgrant5_p & v377cb3d | !hgrant5_p & v3750087;
assign v374f0f5 = hbusreq0 & v376f56d | !hbusreq0 & v8455be;
assign v3725252 = hbusreq2 & aab2b0 | !hbusreq2 & v8455e7;
assign v377f0dc = hmaster3_p & v3a59613 | !hmaster3_p & v3760e13;
assign v3a597d8 = hmaster3_p & v3779d09 | !hmaster3_p & !v3a6fee4;
assign v373df7f = hbusreq6_p & v376f56d | !hbusreq6_p & v3775653;
assign v377bd76 = hbusreq8 & v3751e7c | !hbusreq8 & v376ae9f;
assign v3a658a9 = hbusreq6_p & v3752fe6 | !hbusreq6_p & !v37234c3;
assign v3a701a6 = hbusreq2 & v8455b3 | !hbusreq2 & !v3768202;
assign v3808f75 = hmaster1_p & v375ba6d | !hmaster1_p & v376600a;
assign v3769d79 = hbusreq5_p & v3a6f4c9 | !hbusreq5_p & v8455ab;
assign v3a70ae8 = hmaster0_p & v377dacb | !hmaster0_p & v3a6edbe;
assign v3a5741c = hgrant6_p & v3748797 | !hgrant6_p & v8455ab;
assign v374c6aa = hbusreq7_p & v37612d0 | !hbusreq7_p & v373fdce;
assign v3a58fa7 = hmaster0_p & v3a6f781 | !hmaster0_p & v373c8c5;
assign v3a683c6 = hbusreq5_p & v3772f32 | !hbusreq5_p & v3a707b2;
assign v37250b5 = hmaster1_p & v8455ab | !hmaster1_p & v37290ab;
assign v375f83b = hmaster1_p & v3a55b39 | !hmaster1_p & v3746d57;
assign v3757f07 = hbusreq7 & v3757e15 | !hbusreq7 & v8455bf;
assign v373ad95 = locked_p & v8455fd | !locked_p & !v8455ab;
assign v3a70fd1 = hlock6 & v375c439 | !hlock6 & v3738df9;
assign v23fdf14 = hbusreq7 & v3a6f750 | !hbusreq7 & v3741b61;
assign v376c6a8 = hlock0 & v3a64af7 | !hlock0 & v376062f;
assign v372f87f = hgrant2_p & v3a6c580 | !hgrant2_p & v8d428b;
assign v3757c7f = hbusreq6_p & v3725d73 | !hbusreq6_p & v8455ab;
assign v3a5e015 = hbusreq5_p & v3761719 | !hbusreq5_p & v3777da6;
assign v373855c = hbusreq0 & v373ac12 | !hbusreq0 & v372e661;
assign v3a651b8 = hbusreq1 & v35b7808 | !hbusreq1 & v377eb9d;
assign v37655d6 = hgrant0_p & v3753e6a | !hgrant0_p & v37397c3;
assign v37754e6 = hmaster2_p & v376e72d | !hmaster2_p & v372b231;
assign v3769061 = stateG10_1_p & v8455ab | !stateG10_1_p & v39a5382;
assign v372a965 = hgrant5_p & v376bd96 | !hgrant5_p & v375e9ef;
assign v372c334 = hmaster1_p & v8455ab | !hmaster1_p & v3779da3;
assign v3a6375b = hmaster1_p & v3a70987 | !hmaster1_p & v373e944;
assign v3a67b3c = hgrant5_p & v3740a8a | !hgrant5_p & v372f6f9;
assign v3750f49 = hlock0 & v3a5741c | !hlock0 & v37724db;
assign be0e1a = hmaster2_p & v3735e84 | !hmaster2_p & v375a397;
assign v3736411 = hmaster0_p & v3a6fc3b | !hmaster0_p & !v37bfc8b;
assign v374ed57 = hlock0 & v373031f | !hlock0 & v3748ba4;
assign v3806fc0 = hmaster0_p & v373b4aa | !hmaster0_p & v373cde7;
assign v372f16b = hgrant2_p & v8455ab | !hgrant2_p & v38079d7;
assign v373c1e4 = hbusreq7_p & v37434eb | !hbusreq7_p & v373478e;
assign v3740232 = hbusreq6 & v3a5e881 | !hbusreq6 & v3765e79;
assign v3a70dc4 = hbusreq2_p & v3769cff | !hbusreq2_p & v37735a0;
assign v3a6fdb4 = hbusreq1_p & v376887c | !hbusreq1_p & !v8455ab;
assign v3a708d7 = hbusreq5 & v3a6f40f | !hbusreq5 & v3a64ff4;
assign v376513f = jx1_p & b539d9 | !jx1_p & v3a6f0f7;
assign v3736ab1 = hlock0_p & v37270d9 | !hlock0_p & !v1e38224;
assign v3747e73 = hmaster0_p & v8455ab | !hmaster0_p & v3766b05;
assign v376d432 = hmaster1_p & v372cdde | !hmaster1_p & v376644e;
assign v3a705d5 = hmaster2_p & v37793e4 | !hmaster2_p & v3a70374;
assign v3a71287 = hbusreq1_p & v3764834 | !hbusreq1_p & v3739d4a;
assign v3a6f831 = hbusreq5 & v374ab22 | !hbusreq5 & v3771c85;
assign v3a647e0 = hmaster1_p & v372673d | !hmaster1_p & v375ee2e;
assign v375ebdd = hbusreq2_p & v3a29706 | !hbusreq2_p & v372869e;
assign v37348f8 = hbusreq8_p & v3726d60 | !hbusreq8_p & v3778e2d;
assign af0958 = jx0_p & ac69a2 | !jx0_p & v3747133;
assign v39ea273 = hgrant3_p & v3a70272 | !hgrant3_p & !v373c703;
assign v372cb2c = hmaster1_p & bb49f9 | !hmaster1_p & v3a6fef5;
assign v373eea8 = hbusreq7_p & v374d1ed | !hbusreq7_p & !v372d07b;
assign v3a7072d = hmaster1_p & v3a5a6e6 | !hmaster1_p & v3761954;
assign v3771137 = hbusreq2_p & v3761cd3 | !hbusreq2_p & v3766485;
assign v3750eb8 = hgrant6_p & v3772362 | !hgrant6_p & v376614b;
assign v3724a65 = hbusreq5 & v3a6184c | !hbusreq5 & !v3743f4d;
assign v3a58803 = hbusreq5_p & v3772080 | !hbusreq5_p & v360d140;
assign v35772a6 = stateA1_p & v8455e1 | !stateA1_p & v35772a5;
assign v3a6a442 = hgrant6_p & v3759b2f | !hgrant6_p & v3743d58;
assign v377057a = hbusreq3_p & v3a6f43e | !hbusreq3_p & v372935c;
assign v373ea8d = hmaster0_p & v373b11a | !hmaster0_p & v3a53986;
assign v3728604 = hbusreq2_p & v3a6e327 | !hbusreq2_p & v8455ab;
assign v374047d = hbusreq0_p & v23fe285 | !hbusreq0_p & v8455b5;
assign v3a70297 = hbusreq6 & v3775303 | !hbusreq6 & v8455ab;
assign v377f5f2 = hmaster2_p & v3a641d5 | !hmaster2_p & v37450b8;
assign v377f45d = hmaster0_p & v3733a1e | !hmaster0_p & v3a6f291;
assign v377cbb6 = jx0_p & v3a66ca4 | !jx0_p & v37582e6;
assign d438fc = hmaster2_p & v3a635ea | !hmaster2_p & v37267d6;
assign v37658b1 = hbusreq3 & v8455b3 | !hbusreq3 & !v3768202;
assign v3a623ca = hbusreq4_p & v3a6ff08 | !hbusreq4_p & v376e772;
assign v374b20c = hbusreq6 & v377228d | !hbusreq6 & v3a6687c;
assign v3a70bf1 = hbusreq6 & v376e04c | !hbusreq6 & v1e378b4;
assign v3735f31 = hbusreq8_p & v3a6fe92 | !hbusreq8_p & v3a701af;
assign v377ba59 = hgrant4_p & v374f9c6 | !hgrant4_p & v3a58200;
assign v37449fc = hgrant4_p & v374bd09 | !hgrant4_p & v3a6f1fb;
assign v3a715d2 = hlock0_p & v3a70641 | !hlock0_p & v3a646f8;
assign v3a6c892 = hmaster2_p & v375646d | !hmaster2_p & !v8455ab;
assign v1e37dfd = hlock6 & v373ce84 | !hlock6 & v37436a8;
assign v375a579 = hbusreq6_p & v3a637ca | !hbusreq6_p & v374e29a;
assign v373ecd8 = hbusreq0 & v375ccc3 | !hbusreq0 & v3749cf7;
assign v374c13e = hlock4_p & v3378ef7 | !hlock4_p & v8455ab;
assign v380a1f3 = hmaster2_p & v3a29850 | !hmaster2_p & v37641ad;
assign v377d2bc = hbusreq4 & v3a5f0cf | !hbusreq4 & v8455ab;
assign v3731ab1 = hbusreq8_p & v3a6f01d | !hbusreq8_p & v373cf73;
assign v3724fdb = hbusreq0 & v3a6efe2 | !hbusreq0 & v3a70168;
assign v3740110 = hbusreq2_p & v3759032 | !hbusreq2_p & !v39a537f;
assign v3a69bbf = hgrant6_p & v3a69ae7 | !hgrant6_p & v376f505;
assign v8af425 = hmaster2_p & v377234d | !hmaster2_p & v3a6d590;
assign v3a5be6d = hgrant4_p & v3a643a0 | !hgrant4_p & v37545ea;
assign v3a6fc68 = hbusreq5_p & v3a6ef01 | !hbusreq5_p & v373b30b;
assign v373025a = hmaster2_p & v3769740 | !hmaster2_p & v375a397;
assign v375ad91 = hgrant0_p & v37773a9 | !hgrant0_p & v8455e7;
assign v1e378ea = hbusreq4_p & v3a6dbaa | !hbusreq4_p & v3747f81;
assign v3a6d525 = hgrant0_p & v3762cff | !hgrant0_p & !v3753cc4;
assign v38067b3 = hbusreq5_p & v37403b1 | !hbusreq5_p & v37512c1;
assign d7f9ec = hmaster3_p & v3a67d0d | !hmaster3_p & !v3759d9c;
assign v1e37972 = hlock6 & v3a6e105 | !hlock6 & v37686f6;
assign v376daa7 = hbusreq7 & v9d70f0 | !hbusreq7 & v3734d20;
assign v35b708f = hbusreq2 & v3a6f02e | !hbusreq2 & v374cba0;
assign v372309d = hmaster2_p & v360d136 | !hmaster2_p & v3a71133;
assign v3754ce8 = hbusreq5 & v372ab06 | !hbusreq5 & v3a6fa04;
assign v3a70c77 = hlock8_p & v3807a7d | !hlock8_p & v8455c7;
assign v3a56aa0 = hmaster1_p & v372dc8e | !hmaster1_p & v8455ab;
assign v23fe06e = hbusreq2_p & v374f871 | !hbusreq2_p & v8455b0;
assign v3a6c31f = hmaster0_p & v3730060 | !hmaster0_p & v375820e;
assign v3766799 = hlock5 & v3748972 | !hlock5 & v3a6efa1;
assign v3a6fd1c = jx0_p & v37253a5 | !jx0_p & v3a5b3f9;
assign db20f4 = hmastlock_p & v375eb9c | !hmastlock_p & v8455ab;
assign v3a60fa3 = hmaster2_p & v376c902 | !hmaster2_p & v8455ab;
assign b0ac65 = hbusreq7_p & v37585c9 | !hbusreq7_p & v373287a;
assign v3a695c9 = hbusreq4_p & b66740 | !hbusreq4_p & !v2092faa;
assign v372c30a = hbusreq8_p & v3752aa3 | !hbusreq8_p & v3763832;
assign v3a7066d = hlock8 & v372b7e6 | !hlock8 & v373055b;
assign v3733f37 = hbusreq6 & v3a6eb8b | !hbusreq6 & v380730d;
assign v37413d8 = hbusreq6_p & v3747302 | !hbusreq6_p & v37fc910;
assign v374a63c = stateG10_1_p & v373df21 | !stateG10_1_p & v375c956;
assign v3a6f65c = hbusreq0 & v3756430 | !hbusreq0 & v3a6fbd7;
assign v3a65dcf = hgrant4_p & v3a62826 | !hgrant4_p & v3743de1;
assign v3a70220 = hmaster1_p & v1e37405 | !hmaster1_p & v37750e4;
assign v3a6f052 = hbusreq3 & v3a6ab5f | !hbusreq3 & !v3776fa4;
assign v37548f4 = hmaster2_p & v3a5bf04 | !hmaster2_p & !v3728e09;
assign v3a60a84 = hmaster2_p & v3a62968 | !hmaster2_p & v3765740;
assign v3a70933 = hbusreq5 & v375a6be | !hbusreq5 & v3a6811a;
assign v3747917 = hlock7 & v376ea88 | !hlock7 & v3a5bc4f;
assign v373cee7 = hlock4_p & v3743da0 | !hlock4_p & v37406d2;
assign v3a65660 = hbusreq3_p & v376db8a | !hbusreq3_p & v3a708ef;
assign v94e9e0 = hmaster2_p & v3a56df7 | !hmaster2_p & v8455ab;
assign v374066d = hmaster0_p & v8455b3 | !hmaster0_p & !v8455ab;
assign v374d52a = hgrant4_p & v23fdf76 | !hgrant4_p & v3756506;
assign v3731eca = hbusreq5_p & v3a64a83 | !hbusreq5_p & v3722d5a;
assign v3a5897a = hmaster1_p & v8455e7 | !hmaster1_p & v3a5f60c;
assign v37418db = hbusreq5_p & v373f940 | !hbusreq5_p & v3a5d590;
assign v3a64c10 = hlock0_p & v35b774b | !hlock0_p & !v8455b5;
assign v374131b = hlock5_p & v37437c1 | !hlock5_p & v3a6d3f2;
assign v377a3ec = hlock0 & v375cf36 | !hlock0 & v374a67d;
assign v3a5b912 = hmaster2_p & v3a635ea | !hmaster2_p & v37651c2;
assign v373fc30 = hbusreq1_p & v360d1ca | !hbusreq1_p & v3a5c559;
assign v3a70a89 = hbusreq5 & v376d172 | !hbusreq5 & v23fd9e1;
assign v37694a0 = hmaster0_p & v37721cb | !hmaster0_p & v3a71251;
assign v376eb3c = hbusreq7 & v375a8a7 | !hbusreq7 & v3a647ce;
assign v37697ca = hbusreq5 & v3a6f65e | !hbusreq5 & v3747926;
assign v3a6ff16 = hmaster0_p & v3a70b63 | !hmaster0_p & v3a712d4;
assign v3a6fc5a = hmaster0_p & v3a6931f | !hmaster0_p & v8455e7;
assign v3a6557d = hbusreq1_p & v37568c8 | !hbusreq1_p & !v8455ab;
assign v3a6e81e = hgrant6_p & v3759032 | !hgrant6_p & v3a64d23;
assign v3a7143c = hbusreq2 & v37482f8 | !hbusreq2 & !v372b24d;
assign v3a70c17 = hmaster1_p & v376cd0d | !hmaster1_p & v3a60247;
assign v1e37c0d = hbusreq0 & v3a6f17b | !hbusreq0 & v37573a3;
assign v377d254 = hbusreq2 & v375309f | !hbusreq2 & !v8455ab;
assign v375d7bc = hmaster1_p & v375fb00 | !hmaster1_p & !v3a715d1;
assign v373e0ad = hgrant3_p & v8455be | !hgrant3_p & v37749fd;
assign v373a66d = hbusreq1 & v3740171 | !hbusreq1 & v8455e7;
assign v373ca53 = hgrant6_p & v377f09a | !hgrant6_p & v377b49d;
assign v37252d0 = hgrant2_p & v8455ba | !hgrant2_p & v3a68d3f;
assign v373e04e = hbusreq5_p & v376b4a2 | !hbusreq5_p & v3a6a4b0;
assign v3a70b51 = hgrant6_p & v373c81c | !hgrant6_p & v3a6599b;
assign v3722fc5 = hmaster0_p & v3a701a1 | !hmaster0_p & v372adb6;
assign v376bc8c = hmaster0_p & v3a66110 | !hmaster0_p & v3a6750f;
assign v3a705f1 = hbusreq5_p & v37525c8 | !hbusreq5_p & v377cef3;
assign v374953c = hmaster2_p & v8455ab | !hmaster2_p & v374c840;
assign v376ef47 = hmaster1_p & v376c2e6 | !hmaster1_p & v373adb9;
assign v3751ffd = hbusreq5 & v37572af | !hbusreq5 & v3755731;
assign v373700d = hbusreq5 & v38093a8 | !hbusreq5 & !v8455ab;
assign v3a6f77c = hgrant0_p & v8455ab | !hgrant0_p & d9767c;
assign v376410a = hgrant6_p & v37780cd | !hgrant6_p & v372d0de;
assign v3a609da = hmaster0_p & v374e855 | !hmaster0_p & v3777e7d;
assign v374b8fa = hgrant4_p & v3a53eeb | !hgrant4_p & v375c845;
assign v3a6efa1 = hmaster0_p & v3a5f7b8 | !hmaster0_p & v3a6ddea;
assign v375f3e2 = hbusreq6_p & v372d397 | !hbusreq6_p & !v8455ca;
assign v3a5f4b2 = hlock3_p & v377ea73 | !hlock3_p & !v8455ab;
assign v3749f9d = hbusreq7_p & v377118b | !hbusreq7_p & v3724f05;
assign v3a57d9e = hlock0 & v3757009 | !hlock0 & v3a5e3be;
assign v3759bf4 = hlock5 & v3756305 | !hlock5 & v375138c;
assign v377e124 = hgrant1_p & v3778528 | !hgrant1_p & v8455ab;
assign v3a6e8d9 = hmaster2_p & v37408e1 | !hmaster2_p & v374d6b2;
assign v376beea = hbusreq8_p & v3760da6 | !hbusreq8_p & v376b6ba;
assign v3770f48 = hbusreq5 & v3a59746 | !hbusreq5 & v3a7122f;
assign v3742ef6 = hbusreq3 & v3731258 | !hbusreq3 & v8455ab;
assign v3741cb9 = hbusreq3 & v3a6f7bf | !hbusreq3 & v8455e7;
assign v375c07c = hmaster1_p & v375f071 | !hmaster1_p & v376abd3;
assign v376ce55 = hbusreq5_p & v3a5c066 | !hbusreq5_p & v372e2cd;
assign v3755bbf = hlock5_p & v3a7083c | !hlock5_p & v3a6826d;
assign v376282b = stateG2_p & v3a5a496 | !stateG2_p & !v373180e;
assign v3a6eb4f = hbusreq8_p & v3a70ff2 | !hbusreq8_p & !v8455ab;
assign v3a5d04e = hbusreq3_p & v8455ab | !hbusreq3_p & v377c185;
assign v376e5d2 = hlock0 & v38072fd | !hlock0 & v37522ea;
assign v3760a58 = hbusreq4_p & v3727eda | !hbusreq4_p & v8455ab;
assign v375aa9b = hmaster1_p & v375db64 | !hmaster1_p & v37253dc;
assign v3a6446a = start_p & v3a59da9 | !start_p & v376de0b;
assign v3809f5f = hbusreq2_p & v377773f | !hbusreq2_p & v373125c;
assign v37558b4 = hgrant2_p & v8455ab | !hgrant2_p & v3a683a4;
assign v3a7012d = hgrant6_p & v8455ab | !hgrant6_p & v374c1a9;
assign v37349b9 = hmaster2_p & v37583be | !hmaster2_p & !v3a5f83e;
assign v3a6bf63 = hbusreq4 & v377fc4b | !hbusreq4 & v3727084;
assign v3a6f4f9 = hbusreq5_p & v3733e30 | !hbusreq5_p & v3a69b77;
assign v3809e3c = hmaster1_p & v374c0d0 | !hmaster1_p & v3730b8c;
assign v380880f = hbusreq8 & v8455b0 | !hbusreq8 & v3a69973;
assign v3746ea0 = hmaster2_p & v374fe8e | !hmaster2_p & v3a70118;
assign v372f04d = hlock5_p & v2acafaa | !hlock5_p & v3a60594;
assign v3732853 = hbusreq8 & v1e37af7 | !hbusreq8 & v372a2e4;
assign v375aea6 = hgrant6_p & v374d0e3 | !hgrant6_p & v380956e;
assign v9014db = hbusreq5_p & v3809561 | !hbusreq5_p & v374fb30;
assign v37569ec = hgrant2_p & v372d1a4 | !hgrant2_p & v3255a07;
assign v372f721 = hbusreq7_p & v3a55290 | !hbusreq7_p & v374bb16;
assign v3768c21 = hgrant1_p & v3a53877 | !hgrant1_p & v3740171;
assign v3766746 = hmaster2_p & v3730695 | !hmaster2_p & v8455ab;
assign v375134f = hbusreq5_p & v373e70e | !hbusreq5_p & !v3764c0d;
assign v372b75b = hbusreq2 & v37482f8 | !hbusreq2 & !v3a709ea;
assign v372923a = hbusreq2_p & v37273c2 | !hbusreq2_p & v37565ae;
assign v37647d8 = hgrant4_p & v8455ab | !hgrant4_p & v3a7115a;
assign v3a6581b = hmaster2_p & v373d27f | !hmaster2_p & v372988e;
assign v377cb0b = hbusreq5_p & v38076cf | !hbusreq5_p & v375f888;
assign v377dbd3 = hlock5 & v372787e | !hlock5 & v372f235;
assign v3a700c6 = hmaster0_p & v37245f8 | !hmaster0_p & v377609f;
assign v35ba1cf = hmaster0_p & v377c2d9 | !hmaster0_p & v3777817;
assign v9a641e = hmaster3_p & v3a71292 | !hmaster3_p & v37625d5;
assign b95be3 = hbusreq2_p & v3a70f3e | !hbusreq2_p & v374d479;
assign v3a57e56 = hmaster0_p & v3a6a678 | !hmaster0_p & !v3a58b9f;
assign v3a6f7b7 = jx3_p & v3724dfb | !jx3_p & v37348c9;
assign v3a6b4a6 = hgrant2_p & v37443ab | !hgrant2_p & v37607e8;
assign v3a65388 = hbusreq5_p & v3747d82 | !hbusreq5_p & v3a703a3;
assign v3a711df = hmaster2_p & v3a6ab5f | !hmaster2_p & v3773fdc;
assign v37665c9 = hmaster1_p & v37526ca | !hmaster1_p & !v372e1b6;
assign v37523c6 = hbusreq5 & v3a62cb7 | !hbusreq5 & v3a6f2ee;
assign v3770e77 = hgrant5_p & v88b8eb | !hgrant5_p & v3a6f72f;
assign v375446f = hmaster1_p & v3723ef8 | !hmaster1_p & v3736041;
assign v3763fdc = hbusreq0 & v8455b0 | !hbusreq0 & v8455ab;
assign v3759605 = hgrant2_p & v3751d98 | !hgrant2_p & v37441e0;
assign v377094b = hbusreq1_p & v3778ef8 | !hbusreq1_p & !v3a5bbed;
assign v3a707aa = hbusreq4 & v3a5af1e | !hbusreq4 & v375b9c1;
assign v37293ea = hgrant6_p & v8455ab | !hgrant6_p & v3754903;
assign v375c65a = hmaster2_p & v3772ee4 | !hmaster2_p & v3775ad3;
assign v374d85e = hlock0_p & v3732d4b | !hlock0_p & v8455ab;
assign v3a5ff76 = hbusreq2_p & v376c017 | !hbusreq2_p & !v3778a89;
assign v377b673 = hbusreq1_p & v3766452 | !hbusreq1_p & !v39a537f;
assign v3a6f2d5 = jx1_p & v375f069 | !jx1_p & v9bba04;
assign v3a6f6dd = jx1_p & v3762817 | !jx1_p & v3a6fa56;
assign v3751e62 = hbusreq5 & v3768e0e | !hbusreq5 & v3a63f9a;
assign v37796c5 = hgrant4_p & v377b94f | !hgrant4_p & v377e8ca;
assign v3a5e80e = hbusreq3_p & v373afb4 | !hbusreq3_p & v3776a6e;
assign v3768ec4 = hbusreq6_p & v3a6fc11 | !hbusreq6_p & v3a5ee3a;
assign v375cd4c = hbusreq0 & v3a6f618 | !hbusreq0 & v372bfd3;
assign v3a5e0cc = stateA1_p & v8455ab | !stateA1_p & !v3a6b059;
assign v3a71425 = hlock4 & v374c61d | !hlock4 & v3771ab9;
assign v3a5c816 = hbusreq5_p & v3775a9f | !hbusreq5_p & v3731aac;
assign v3751d7d = hbusreq4_p & v3a70641 | !hbusreq4_p & v8455e7;
assign v374771c = hmaster1_p & v3a634fd | !hmaster1_p & v8a7af6;
assign v3741418 = hlock7 & v3735a7f | !hlock7 & v3742676;
assign v3773aa0 = hbusreq2 & v3763a20 | !hbusreq2 & v8455bf;
assign d193f7 = hmaster1_p & v37776f0 | !hmaster1_p & v375652a;
assign v3a5b4d6 = hlock8 & v373bd70 | !hlock8 & v3377adc;
assign v3766b81 = hlock2 & v377c6e8 | !hlock2 & v37660d2;
assign v3a57012 = hbusreq6_p & v3a6f050 | !hbusreq6_p & v372cc25;
assign v372a264 = hmaster1_p & v3a6ff31 | !hmaster1_p & !v3755096;
assign v372f72b = hgrant3_p & v35b7299 | !hgrant3_p & !v8455ab;
assign v37732c0 = hlock1_p & v37502b7 | !hlock1_p & v376f9a8;
assign v37713fe = hlock0 & v3a6c5ee | !hlock0 & v3a6e7d8;
assign v37627f9 = hgrant2_p & v8455ba | !hgrant2_p & v375b4a7;
assign v373f3e4 = hlock7 & v3a54222 | !hlock7 & v3a64e75;
assign v374717a = hbusreq8_p & v37614fa | !hbusreq8_p & v39ebad8;
assign v374328c = hmaster2_p & v374502e | !hmaster2_p & !v8455ab;
assign v3752183 = hmaster0_p & v37469c4 | !hmaster0_p & v373ff5c;
assign v3a5e9b8 = hmaster0_p & v375c791 | !hmaster0_p & v3a60b90;
assign v3745236 = hbusreq3_p & v37261df | !hbusreq3_p & !v3a5ae7d;
assign v3723f0c = hmaster1_p & v377c5f8 | !hmaster1_p & v3a6570f;
assign v3767830 = hbusreq8_p & v3762802 | !hbusreq8_p & v3a5b03b;
assign v3760d74 = hgrant6_p & v372672f | !hgrant6_p & v3a712d6;
assign v373df14 = hgrant1_p & v3a637dc | !hgrant1_p & v3763961;
assign v376d9f8 = hmaster0_p & v3a6ff46 | !hmaster0_p & v8455ab;
assign v3736806 = hgrant4_p & v3a6fdde | !hgrant4_p & v3757aa1;
assign v3a5eeb4 = hgrant3_p & v3a62826 | !hgrant3_p & v3a70cc5;
assign v3a70013 = jx0_p & v377a6e2 | !jx0_p & v37548e7;
assign v3769639 = hlock5 & v3771c38 | !hlock5 & b8f5a8;
assign v3777cfc = hgrant4_p & v3a59505 | !hgrant4_p & v374bf59;
assign v372cc69 = hmaster0_p & v377df7d | !hmaster0_p & !v3a7163a;
assign v376bad7 = hmaster2_p & v2092bdc | !hmaster2_p & v3771dda;
assign v3744a9c = hbusreq5 & v3770425 | !hbusreq5 & v373497f;
assign v3a64977 = hmaster2_p & v3a6a289 | !hmaster2_p & v3a6da3b;
assign v3a6febe = hbusreq5 & v3a5e9b8 | !hbusreq5 & v3a55eda;
assign v3a6fa84 = hlock4_p & v3a710c6 | !hlock4_p & v8455bb;
assign v372e3db = hbusreq8_p & v37434eb | !hbusreq8_p & v373c1e4;
assign v3776b09 = hmaster2_p & v8455ca | !hmaster2_p & v37770ed;
assign v3734502 = hmaster0_p & v374314f | !hmaster0_p & v3a5f281;
assign v3a6effd = hlock7_p & d973ae | !hlock7_p & v375055f;
assign v3743a77 = hbusreq5 & v376a6f1 | !hbusreq5 & v377ac1e;
assign v377b3be = hmaster0_p & v3a5ce35 | !hmaster0_p & v3a69606;
assign v3a5e3c0 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a6e868;
assign v37392e0 = hbusreq5 & v3773633 | !hbusreq5 & v375e037;
assign v37c00f6 = hbusreq5 & v3769245 | !hbusreq5 & v3a7122f;
assign v3a655c3 = hbusreq1 & v376a8d5 | !hbusreq1 & v3a57309;
assign v3772b42 = hbusreq8_p & v3a6f76d | !hbusreq8_p & v3a6fc97;
assign v375be12 = hbusreq6_p & v3727ce4 | !hbusreq6_p & v372f5bd;
assign v3a6e516 = hgrant3_p & v37579a9 | !hgrant3_p & v3770bd9;
assign v375830c = hmaster1_p & v3744399 | !hmaster1_p & v3a6e675;
assign db1dc4 = hmaster0_p & v3768358 | !hmaster0_p & v372a674;
assign v3a6f0e7 = hbusreq6_p & v374ab1e | !hbusreq6_p & v3773d82;
assign v376e056 = hmaster2_p & v376029a | !hmaster2_p & v3a70e03;
assign v3756cf2 = hbusreq5_p & v3a700d9 | !hbusreq5_p & v8455ab;
assign v3a69ec5 = hmaster1_p & v360d0c7 | !hmaster1_p & v376a3f5;
assign v3755786 = hbusreq5_p & v37392e2 | !hbusreq5_p & !v8455ab;
assign v3a70ad1 = hbusreq7_p & v3759e04 | !hbusreq7_p & v3725bdd;
assign v372bfa1 = hbusreq6_p & v3731fc6 | !hbusreq6_p & v3a699a1;
assign v3a70a12 = locked_p & v3a635ea | !locked_p & !v373bce7;
assign v3772ab1 = hbusreq3_p & v372cd45 | !hbusreq3_p & v8455ab;
assign v377fbd5 = hbusreq5_p & v3749e8a | !hbusreq5_p & v37790c8;
assign v3a7044a = hgrant6_p & v8455ab | !hgrant6_p & v374d3b3;
assign v372b2ba = hgrant2_p & v374c523 | !hgrant2_p & v3a707c7;
assign v37240e8 = hgrant3_p & v37712f6 | !hgrant3_p & !v376c2e2;
assign v3a6f8e6 = hgrant4_p & v8455ab | !hgrant4_p & v377c4b8;
assign v2092f5e = hbusreq2 & v3a6b560 | !hbusreq2 & v3748797;
assign v3758e9e = hlock6_p & v376653d | !hlock6_p & v8455ab;
assign v373f691 = hmaster0_p & d58c24 | !hmaster0_p & v35b774b;
assign v3a5565d = hmaster0_p & v3a635ea | !hmaster0_p & v372d98c;
assign v3759fe8 = hlock2_p & v3772ae7 | !hlock2_p & v3728e25;
assign v3a70676 = hbusreq7 & v3730252 | !hbusreq7 & v376fdd4;
assign v3a54d04 = hbusreq8_p & v3731376 | !hbusreq8_p & !v8455ab;
assign v3a5a29e = hbusreq2_p & v3a713be | !hbusreq2_p & v3a635ea;
assign v3735fca = hgrant4_p & v3a70460 | !hgrant4_p & v3a714ad;
assign aac430 = hgrant2_p & v3a635ea | !hgrant2_p & b08e51;
assign v1e37556 = hbusreq4 & v31c369c | !hbusreq4 & v3a5f9e6;
assign v3730de2 = hgrant6_p & v3739884 | !hgrant6_p & v2ff9268;
assign v3728581 = hmaster3_p & v373fe61 | !hmaster3_p & v3739a9f;
assign v3a606b9 = hbusreq7 & bdc0a1 | !hbusreq7 & v39a5359;
assign v377f694 = hbusreq8 & v3777602 | !hbusreq8 & v3737808;
assign v33781df = hgrant4_p & v37622f5 | !hgrant4_p & v373f488;
assign v38064e5 = hmaster0_p & v376f111 | !hmaster0_p & v376a6f1;
assign v3a6fddd = hgrant2_p & v8455ab | !hgrant2_p & v3731906;
assign v3a5f239 = hbusreq4 & v3723430 | !hbusreq4 & v8455ab;
assign v3a5d153 = jx0_p & v375ece3 | !jx0_p & v3733249;
assign v377cdf1 = hmaster1_p & v3759611 | !hmaster1_p & v376f2fc;
assign v3a57dbb = hbusreq8_p & v3a5eb63 | !hbusreq8_p & v38097c4;
assign v372998c = hbusreq1_p & v3a635ea | !hbusreq1_p & !v377ed71;
assign v3a7045e = hmaster2_p & v377ba09 | !hmaster2_p & v3a70fdb;
assign v374bec6 = hgrant2_p & v3a59bb4 | !hgrant2_p & v39a4e8f;
assign v3777460 = hlock4_p & v3724a4b | !hlock4_p & v3730ffe;
assign v3a57108 = hbusreq5 & v3779797 | !hbusreq5 & v3771c85;
assign v3728a12 = hbusreq6_p & v376655b | !hbusreq6_p & v3740374;
assign v377564a = hgrant4_p & v377b6ce | !hgrant4_p & v3a53ffa;
assign v374cd2c = hmaster2_p & v3753dab | !hmaster2_p & v37386cb;
assign v373b0f5 = jx3_p & v3751fde | !jx3_p & v376f261;
assign v3761553 = hgrant4_p & v8455ab | !hgrant4_p & v3a70e79;
assign v3a5f6a8 = hbusreq7 & v37745e9 | !hbusreq7 & v3770edc;
assign v372981e = stateG10_1_p & v37328bf | !stateG10_1_p & v373178e;
assign v3a67ffd = hbusreq5_p & v3774e33 | !hbusreq5_p & v377a10f;
assign v3735554 = hgrant6_p & v375c7b9 | !hgrant6_p & !v3765722;
assign v3a6f9b3 = hgrant4_p & v8455ab | !hgrant4_p & v3a6ec1f;
assign v3a6f963 = hbusreq4_p & v3a5fc59 | !hbusreq4_p & !v8455ab;
assign v3a6f95a = hmaster2_p & v3778528 | !hmaster2_p & v8455ab;
assign v372f346 = hbusreq4_p & v375da82 | !hbusreq4_p & v3725717;
assign v3a6a918 = hbusreq7_p & v3a71675 | !hbusreq7_p & v35b708c;
assign v373fb22 = hbusreq5_p & v3a6ffee | !hbusreq5_p & v3a702f6;
assign v3a5fcf0 = hlock8_p & v372eb0f | !hlock8_p & v3a70333;
assign v3756eca = hgrant6_p & v8455ab | !hgrant6_p & v3a59391;
assign v373f349 = hmaster0_p & v8455c3 | !hmaster0_p & v377230a;
assign v23fda6c = hbusreq8 & v375b24f | !hbusreq8 & v3a71448;
assign v373f4a9 = hmaster0_p & v374cd2c | !hmaster0_p & v373ef01;
assign v3a5f451 = hmaster0_p & v3a5d678 | !hmaster0_p & v3770174;
assign v377d651 = hbusreq0 & v3a539af | !hbusreq0 & v3a64af7;
assign v3a6df62 = hgrant7_p & v8455ce | !hgrant7_p & v376e860;
assign v37617de = hgrant6_p & v37379fc | !hgrant6_p & v3a70832;
assign v3a70695 = hmaster1_p & v3a6f1c1 | !hmaster1_p & v3764805;
assign v3752d31 = hbusreq7 & v374e82c | !hbusreq7 & v37728cd;
assign v373335b = hbusreq5_p & v3a60b56 | !hbusreq5_p & !v8455ab;
assign v3726da1 = hbusreq5_p & v37752af | !hbusreq5_p & v37657be;
assign v3745e72 = hbusreq4_p & v3a5a2a7 | !hbusreq4_p & v3a7048d;
assign v3a706c5 = hmaster0_p & v3a58cfc | !hmaster0_p & v377bcf5;
assign v376cf62 = hbusreq2_p & v37332dd | !hbusreq2_p & v377957e;
assign v3737053 = hlock2_p & v3a5ec2d | !hlock2_p & v3a5a4a0;
assign v3a6f253 = hmaster1_p & v375f071 | !hmaster1_p & v373e30f;
assign v3748929 = hbusreq5_p & v3a70382 | !hbusreq5_p & v372815e;
assign v375dc43 = hmaster1_p & v372f11d | !hmaster1_p & v374c7e6;
assign v3a66cee = hbusreq8_p & v3757dea | !hbusreq8_p & v374a2b5;
assign v3809583 = hbusreq2 & v3770578 | !hbusreq2 & v8455ab;
assign v37736ad = hbusreq3_p & v3806912 | !hbusreq3_p & v3a5b9ea;
assign v3754685 = hmaster2_p & v3a6fe4e | !hmaster2_p & v375624e;
assign v375a2a7 = hmaster3_p & v3a65521 | !hmaster3_p & v3768ec3;
assign v376025f = hbusreq4_p & v376f56d | !hbusreq4_p & v3767f58;
assign v3a6af93 = hmaster2_p & v8455ab | !hmaster2_p & v3739c68;
assign v3739018 = hbusreq3_p & v375c8e8 | !hbusreq3_p & v3732aca;
assign v3a712da = hbusreq2 & v3752831 | !hbusreq2 & v376bade;
assign v372ffd3 = hbusreq5_p & v3a61a2d | !hbusreq5_p & v3a715d9;
assign v373a9a9 = hmaster0_p & v3a6e6a7 | !hmaster0_p & v373d4a6;
assign v372fb53 = hgrant5_p & v3a6f6af | !hgrant5_p & v3a6d2eb;
assign v377af98 = hgrant0_p & v8455ab | !hgrant0_p & v374ab5b;
assign v3755665 = hlock2 & v9c4c8d | !hlock2 & v374732a;
assign v3a5ebbf = hmaster0_p & v37464e4 | !hmaster0_p & v3764a7d;
assign v376f449 = hbusreq4_p & v3a70bf7 | !hbusreq4_p & v3761ed2;
assign v3a5dff7 = hbusreq7 & v3a64200 | !hbusreq7 & v3a6f1e8;
assign v3a6687c = hgrant2_p & v3748797 | !hgrant2_p & v8455ab;
assign v39eb3d2 = hbusreq5 & v37645bc | !hbusreq5 & v8455ab;
assign v37563cf = hlock5_p & v8455ab | !hlock5_p & v37514c2;
assign v3a6f356 = hbusreq7 & v3a715fa | !hbusreq7 & !v375e64d;
assign v3755b55 = hbusreq8_p & v3a7156c | !hbusreq8_p & v3a708f8;
assign v3a6fc73 = hbusreq5 & v377dfa2 | !hbusreq5 & v3378fc3;
assign v3763c04 = hbusreq2 & v373fe5e | !hbusreq2 & v8455ab;
assign v3a6b083 = hbusreq1_p & v3a6f7de | !hbusreq1_p & !v3754c0e;
assign v374a79e = hmaster1_p & v3a635ea | !hmaster1_p & v377eab7;
assign v3a710d0 = hmaster2_p & v377564a | !hmaster2_p & v2925c5b;
assign v374d121 = hmaster1_p & v3724394 | !hmaster1_p & v377e2e3;
assign v3765436 = hbusreq0_p & v8455ab | !hbusreq0_p & v37665bf;
assign v373b17e = hlock7 & v376ad04 | !hlock7 & v3a6209f;
assign v3a6f6a8 = hmaster0_p & v3a66110 | !hmaster0_p & v3a6f82c;
assign v3a7110e = hbusreq5 & v3a6870f | !hbusreq5 & !v8455c2;
assign v37376f9 = hgrant6_p & v1e37cd6 | !hgrant6_p & v372d238;
assign v3a70499 = hbusreq5_p & v37568c9 | !hbusreq5_p & v3778f46;
assign v360d166 = hmaster2_p & v3a635ea | !hmaster2_p & v377ad76;
assign v375351d = hmaster2_p & v3a64f7e | !hmaster2_p & v3769374;
assign v3a63a66 = hlock4_p & v3736ded | !hlock4_p & v8455bb;
assign v372b5af = hgrant3_p & v8455ab | !hgrant3_p & v3a70895;
assign v373ae91 = hgrant2_p & v8455b9 | !hgrant2_p & v375b713;
assign v38078e5 = hlock4 & v3769e4c | !hlock4 & v3a6fd6a;
assign v3a5a2d0 = hmaster3_p & v37594ae | !hmaster3_p & v3754bb9;
assign v3733e77 = hmaster2_p & v373ce86 | !hmaster2_p & v3750edc;
assign v3774b66 = hmaster1_p & v3a70f0c | !hmaster1_p & v3a6fd9b;
assign v3a702b5 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a68f4d;
assign v3742fbf = jx0_p & v3741286 | !jx0_p & v3768e31;
assign v3a53c87 = hbusreq5 & v377e283 | !hbusreq5 & v3778ab3;
assign v374df45 = hbusreq4 & v3a68e71 | !hbusreq4 & v3a62a6d;
assign v3a713be = hgrant3_p & v3a635ea | !hgrant3_p & v337830d;
assign v377f505 = hmaster2_p & v3a66110 | !hmaster2_p & !v3a5bf04;
assign v374d140 = hlock0_p & v376d9ad | !hlock0_p & v3a619c0;
assign v376c8ea = hlock0_p & v3a635ea | !hlock0_p & !v3a6fd2a;
assign v3a7029e = hmaster2_p & v377d107 | !hmaster2_p & v3a68084;
assign v37447e2 = hbusreq6_p & v3377b1b | !hbusreq6_p & v3727db9;
assign v377bde3 = hmaster1_p & v3758cec | !hmaster1_p & v372ed79;
assign v3a6d627 = hbusreq0 & v37678fc | !hbusreq0 & v8455ab;
assign v37523e9 = hbusreq6 & v374944b | !hbusreq6 & v3756c25;
assign v3767463 = hbusreq6_p & v3a6770f | !hbusreq6_p & v37526cd;
assign v375e0cb = hlock5_p & v3a5a510 | !hlock5_p & !v373e163;
assign v374dc99 = hmaster1_p & v374e4c5 | !hmaster1_p & v3779613;
assign v377e6fc = hmaster2_p & v3a70987 | !hmaster2_p & v373f6ee;
assign v3a5495d = hbusreq3 & v374362e | !hbusreq3 & v8455ab;
assign v3755a05 = hbusreq2_p & v373f0ee | !hbusreq2_p & v3a69946;
assign v37525c7 = hbusreq0 & v3a6af67 | !hbusreq0 & v37294db;
assign v374a7f0 = hgrant2_p & v3768486 | !hgrant2_p & v3732bc0;
assign v37764ee = hgrant3_p & v8455be | !hgrant3_p & !v3a65660;
assign v3a702f7 = hbusreq6_p & v372599c | !hbusreq6_p & v3737084;
assign v3729bf3 = hgrant6_p & v8455ab | !hgrant6_p & v35ba2dd;
assign v374e246 = hgrant6_p & v3730926 | !hgrant6_p & v374421d;
assign v3726ee7 = hlock5_p & v37644ff | !hlock5_p & v3a6fdcb;
assign v3a6efc8 = hbusreq6_p & v37367f1 | !hbusreq6_p & v3760b3d;
assign v3a6ca54 = hbusreq5 & v3a58c07 | !hbusreq5 & v8455ab;
assign v3762700 = hlock3_p & v3773ee6 | !hlock3_p & v8455b3;
assign v3a71299 = hmaster2_p & v37386f5 | !hmaster2_p & !v3a6bc65;
assign v3a671a2 = hgrant3_p & v3a6b873 | !hgrant3_p & v3a7003e;
assign v374b43d = hgrant2_p & v3739ca8 | !hgrant2_p & v37675f4;
assign v3a5bb6a = hbusreq4_p & v3740c8e | !hbusreq4_p & v8455ab;
assign v3a54a24 = hgrant7_p & v3a70008 | !hgrant7_p & v37393e8;
assign v3773f85 = hmaster1_p & v8455ab | !hmaster1_p & !v3a705a2;
assign v1e37cba = hmaster0_p & v3756a05 | !hmaster0_p & v3726262;
assign v37274a1 = hmaster3_p & v3755640 | !hmaster3_p & v374d14a;
assign v37497ce = hmaster0_p & v3752333 | !hmaster0_p & v3731bb5;
assign v37301d8 = hmaster2_p & v3775dbc | !hmaster2_p & v374eab4;
assign v3760513 = hbusreq4_p & v8455bb | !hbusreq4_p & v3727084;
assign v3a71202 = hmaster2_p & v3a61734 | !hmaster2_p & v3a6eb47;
assign v3a6c40d = jx1_p & v3a53f1c | !jx1_p & v3749b2e;
assign v3768ab0 = hgrant0_p & v3a5e24e | !hgrant0_p & c99197;
assign v3a5968c = hbusreq1 & v3740f3d | !hbusreq1 & !v8455ab;
assign v3a67cd1 = hlock0 & v373031f | !hlock0 & v376a149;
assign v3a6f8b5 = hmaster1_p & v3809cc0 | !hmaster1_p & v3a53fb5;
assign v3748932 = hlock3_p & v3a548b2 | !hlock3_p & v8455b0;
assign v3a5f41d = hgrant2_p & v3a70403 | !hgrant2_p & v3756ebb;
assign v3a7084c = hbusreq4 & v3a713cc | !hbusreq4 & v3771536;
assign v3a6de8c = hlock3_p & aefb3e | !hlock3_p & v3755381;
assign v3a5f894 = hmaster1_p & v376c248 | !hmaster1_p & v3a57721;
assign v375af99 = hmaster2_p & v3779736 | !hmaster2_p & !v380951e;
assign v3a681ed = hgrant4_p & v8455ab | !hgrant4_p & v3727b18;
assign v3a70ca4 = hmaster2_p & v8455ab | !hmaster2_p & v3a6a973;
assign v373f8fb = hbusreq1_p & v374270d | !hbusreq1_p & v3a56396;
assign v3a5a219 = hmaster0_p & v3a7149d | !hmaster0_p & v3771160;
assign v376572c = hlock6 & v376999e | !hlock6 & v39a5293;
assign v3745e0e = hmaster1_p & v3807183 | !hmaster1_p & v377f640;
assign v3727342 = hbusreq5 & v376babf | !hbusreq5 & v8455c7;
assign v375b82d = hbusreq4_p & v3a59158 | !hbusreq4_p & v8455ab;
assign v3a59264 = hgrant6_p & v37325cf | !hgrant6_p & v3a555d1;
assign v3769c6d = hmaster0_p & v3756dd8 | !hmaster0_p & v374e6b1;
assign v3a67996 = hlock5_p & v8455ab | !hlock5_p & v3758bfe;
assign v372bb82 = hgrant5_p & v8455ab | !hgrant5_p & v3a5a307;
assign v3a70554 = hbusreq0 & v3a5def2 | !hbusreq0 & v377c31d;
assign v3a63e9e = hlock2 & v37477dd | !hlock2 & v3725f24;
assign v375bd37 = hbusreq4 & v373a47e | !hbusreq4 & !v8455ab;
assign v37790bd = hbusreq8 & v3765f8e | !hbusreq8 & v8455ab;
assign v375946b = hgrant4_p & v3751968 | !hgrant4_p & !v375e3d1;
assign v3777342 = hbusreq4 & v373a588 | !hbusreq4 & v8455ab;
assign v3766222 = hbusreq5 & v372f151 | !hbusreq5 & v3730c3c;
assign v3a62ee2 = hmaster1_p & v37710c7 | !hmaster1_p & v3a545a7;
assign v3a6ffce = hmaster1_p & v3a6f469 | !hmaster1_p & v3776bc7;
assign v3a5e755 = jx0_p & v3a6f4cc | !jx0_p & v375b84e;
assign v376d287 = hbusreq5_p & v37363ae | !hbusreq5_p & v3a6c7e8;
assign v37485e0 = hlock3 & v3a70486 | !hlock3 & v3723247;
assign v3a6fe4d = hmaster2_p & v3751004 | !hmaster2_p & v373bb90;
assign v3a66170 = hlock5_p & v3a66161 | !hlock5_p & v3a6faae;
assign v3764d82 = hmaster2_p & v3739ab4 | !hmaster2_p & !v8455ab;
assign v37249f1 = hgrant3_p & v8455ab | !hgrant3_p & v3731688;
assign v373cada = hbusreq5_p & v375d15c | !hbusreq5_p & v3a6f08d;
assign v3a622f5 = hgrant6_p & v3a59b9e | !hgrant6_p & v3740e7d;
assign v3743332 = hlock0 & v3a6bf41 | !hlock0 & v3a63002;
assign v3a5a1ef = hmaster0_p & v37606e1 | !hmaster0_p & v3a6567f;
assign v3a5f9d5 = hmaster0_p & v372c03b | !hmaster0_p & v376d07b;
assign v374e5fa = hmaster0_p & v373464d | !hmaster0_p & v3a6d407;
assign v377f26e = hmaster0_p & v372673d | !hmaster0_p & v3756109;
assign v3762545 = hbusreq6_p & v375b7fa | !hbusreq6_p & v374a7b2;
assign v374f9cc = hmaster0_p & v3a6c0ab | !hmaster0_p & v8455bd;
assign v376c712 = hbusreq7_p & v3a53dfc | !hbusreq7_p & v3767919;
assign v3a6eeba = hbusreq6_p & v3a70970 | !hbusreq6_p & v3723ee7;
assign v38064a3 = hmaster1_p & v3775902 | !hmaster1_p & v3a64641;
assign v3a6891e = hbusreq1 & v3a581bd | !hbusreq1 & v3a635ea;
assign v3738ca1 = hbusreq5_p & v3a60974 | !hbusreq5_p & v3748460;
assign v374e843 = hmaster0_p & v3743726 | !hmaster0_p & v3a5ae95;
assign v3a67aaa = hlock3 & v3a710c2 | !hlock3 & v37317a9;
assign v3757656 = hbusreq2_p & v377ef7c | !hbusreq2_p & v3757fcc;
assign v3a70a51 = hgrant4_p & v3a5b6de | !hgrant4_p & v38078ed;
assign v3745790 = hmaster0_p & v8455ab | !hmaster0_p & v375792f;
assign v377f180 = hgrant6_p & v3743cd6 | !hgrant6_p & v372300f;
assign v3a57e01 = hbusreq8_p & v373c275 | !hbusreq8_p & v3769c72;
assign v3a572ee = hmaster1_p & v3762e8d | !hmaster1_p & v374fc17;
assign v3732632 = hbusreq7 & v3a71338 | !hbusreq7 & !v3765e47;
assign v373125c = hgrant3_p & v8455bd | !hgrant3_p & v375018e;
assign v3a6eb4a = hgrant2_p & v3a5a510 | !hgrant2_p & v3a702c6;
assign v3a56918 = hgrant5_p & v373ad69 | !hgrant5_p & v3a6f730;
assign v3745b60 = hlock0 & v3809ec3 | !hlock0 & v377bbbd;
assign v372fb48 = hbusreq4_p & v3a6a934 | !hbusreq4_p & v3a6ffcc;
assign v3a6f4a4 = hmaster0_p & v374b522 | !hmaster0_p & v3757966;
assign v3758ea7 = hbusreq0 & v3726cc1 | !hbusreq0 & v3a5e5d0;
assign v3a5dde0 = hbusreq4 & v3a6bc65 | !hbusreq4 & v8455b9;
assign v3739bcd = hgrant6_p & v377f09a | !hgrant6_p & v373f785;
assign v3a712a3 = hbusreq1 & v3a6ebb7 | !hbusreq1 & v3a635ea;
assign v37711dd = hbusreq0 & v374f7ec | !hbusreq0 & v3727bcb;
assign v3a5a967 = hgrant6_p & v8455ab | !hgrant6_p & v3758a0c;
assign v373823d = hmaster0_p & v3a71066 | !hmaster0_p & v372a520;
assign v37471f0 = hmaster2_p & v372b1dc | !hmaster2_p & v37379bb;
assign v3768e70 = hgrant6_p & v372ffaa | !hgrant6_p & v3772e33;
assign v375b2d9 = hbusreq0 & v3776492 | !hbusreq0 & v3776faf;
assign v374d552 = hgrant3_p & v3770559 | !hgrant3_p & v3a70df1;
assign v3755e1f = hlock5_p & v3a6fde5 | !hlock5_p & !v8455ab;
assign v3744f0d = hgrant2_p & v3a70f74 | !hgrant2_p & v37259bc;
assign v2619ad0 = hgrant1_p & v3a6c0b3 | !hgrant1_p & v8455ab;
assign v375624e = hbusreq0 & v37796c6 | !hbusreq0 & v8455ab;
assign v8a9c95 = hgrant4_p & v37c023b | !hgrant4_p & v375b878;
assign v3776f7f = hgrant2_p & v3758fa7 | !hgrant2_p & v37400bc;
assign v3a70c07 = stateA1_p & v8455ab | !stateA1_p & v3a708aa;
assign v37406a7 = hbusreq2_p & v3766a98 | !hbusreq2_p & v374b4a4;
assign v37798b9 = hmaster0_p & db6de7 | !hmaster0_p & v37793b9;
assign v37570f8 = hbusreq0 & v373e877 | !hbusreq0 & v8455ab;
assign v3a6f43e = hbusreq1_p & v376ef42 | !hbusreq1_p & v3733e9e;
assign v3a62a13 = hbusreq0 & v3729852 | !hbusreq0 & !v1e37cd6;
assign v3a5f40e = hbusreq6_p & v3726efb | !hbusreq6_p & v8455ab;
assign v3a565a1 = hbusreq5_p & v37786f3 | !hbusreq5_p & v377de7f;
assign v3728e58 = hgrant4_p & v374d92c | !hgrant4_p & v3a71028;
assign v372f8c1 = hbusreq3 & v3a5f265 | !hbusreq3 & v3762502;
assign v373f022 = hmaster0_p & v3a70806 | !hmaster0_p & v3726434;
assign v3758f19 = hgrant4_p & v3758e05 | !hgrant4_p & v3a6fe74;
assign v3772aa4 = hlock7_p & v3726d60 | !hlock7_p & !v374a50a;
assign v372673b = hgrant3_p & v8455ab | !hgrant3_p & v37311d6;
assign v3807b27 = hmaster1_p & v3a6906e | !hmaster1_p & v3a70b8f;
assign v3741172 = hgrant8_p & v3760860 | !hgrant8_p & v3a7138f;
assign v3736ecc = hbusreq8 & v3a66ad2 | !hbusreq8 & v8455ab;
assign v3779c09 = hlock7 & v3a6b58f | !hlock7 & v3729d06;
assign v35b70fa = hbusreq8 & v32558c4 | !hbusreq8 & !v8455ab;
assign v3778c7f = hbusreq5 & v9204d4 | !hbusreq5 & v3a5aad8;
assign v3a6a3e5 = hbusreq6_p & v3a6f87f | !hbusreq6_p & v3a6f804;
assign v373f6f0 = hbusreq5_p & v3a6eaba | !hbusreq5_p & v3a6f54e;
assign v377894f = hmaster1_p & v3757966 | !hmaster1_p & v3727e56;
assign v376c747 = hgrant3_p & v8455bd | !hgrant3_p & v3a6f884;
assign v3a6e118 = hmaster2_p & v3724394 | !hmaster2_p & v37326a0;
assign v37793a4 = hgrant4_p & v3722e5c | !hgrant4_p & v37259c7;
assign v375463e = hbusreq4_p & v3734b34 | !hbusreq4_p & v8455ab;
assign v3730e8f = jx1_p & v373e419 | !jx1_p & v8455d1;
assign v374cb97 = hbusreq4_p & v3a7136e | !hbusreq4_p & d2dc90;
assign v3756925 = hbusreq2_p & v3a6e3d1 | !hbusreq2_p & v372cc25;
assign v3743798 = hmaster1_p & v3a635ea | !hmaster1_p & v377638d;
assign v373a222 = hmaster2_p & v3735e39 | !hmaster2_p & !v37432c6;
assign v377c929 = hgrant3_p & v3a67eec | !hgrant3_p & v3a6eb0b;
assign v3a60d50 = hmaster0_p & v3a6f95a | !hmaster0_p & v8455ab;
assign v376e139 = hbusreq1 & v3a6dc08 | !hbusreq1 & v8455b0;
assign v374eb2d = hmaster1_p & v376bb43 | !hmaster1_p & v3a704d6;
assign v3a70d9e = hgrant5_p & v3a6f31d | !hgrant5_p & v3a70c17;
assign v3745b0f = hbusreq4 & v3775a92 | !hbusreq4 & v3a5741c;
assign v3a67603 = hgrant3_p & v376f768 | !hgrant3_p & v3a67698;
assign v3a5b517 = hmaster1_p & v3757169 | !hmaster1_p & v8455ab;
assign v1e37a34 = stateA1_p & v3a6efc9 | !stateA1_p & v3757c6f;
assign v377839d = hgrant2_p & v374a6fc | !hgrant2_p & v3772c89;
assign v3757047 = hgrant8_p & v8455ab | !hgrant8_p & v2093069;
assign v3a6b80e = hgrant2_p & v373dbb0 | !hgrant2_p & !v37275cf;
assign v375a159 = hbusreq7_p & v3a6cf15 | !hbusreq7_p & v3a70490;
assign v373bfd8 = hlock8_p & v375583c | !hlock8_p & v3a691fb;
assign v374cef4 = hbusreq5 & v1e37397 | !hbusreq5 & v374c5fc;
assign v38074ed = hbusreq8_p & v3759569 | !hbusreq8_p & v3807a93;
assign v3752407 = locked_p & v8455ab | !locked_p & v37563eb;
assign v3a6fafa = hbusreq3 & v3a6f7f0 | !hbusreq3 & v8455ab;
assign v3a7168a = hbusreq1_p & v37727be | !hbusreq1_p & v372de52;
assign v23fe20d = hmaster2_p & v3a710c6 | !hmaster2_p & v3736ded;
assign v3756943 = hgrant0_p & v37773a9 | !hgrant0_p & v23fe285;
assign v3727fcb = hmaster2_p & v37457fb | !hmaster2_p & v3a6f7bf;
assign v3759f8b = hbusreq3 & v3a5600a | !hbusreq3 & v375444e;
assign v374821f = hgrant4_p & v8455ab | !hgrant4_p & v3a6a66f;
assign v3a6ff43 = hbusreq0_p & v3757082 | !hbusreq0_p & bbbe50;
assign v3a701f2 = hmaster0_p & v376285a | !hmaster0_p & v373dd36;
assign v376ddb6 = hmaster2_p & v3733da4 | !hmaster2_p & v3a687a7;
assign v3a60974 = hmaster0_p & v376374b | !hmaster0_p & v3a7060a;
assign v3a707f5 = hmaster2_p & v376e3fb | !hmaster2_p & v3a5e8a0;
assign v3743677 = hmaster0_p & v3a6ebf7 | !hmaster0_p & !v3a6f31f;
assign v3755002 = hready & v376147f | !hready & !v8455ab;
assign v3766285 = hbusreq0 & v37701fd | !hbusreq0 & v372d967;
assign v3a6a40b = hbusreq7_p & v372ea2d | !hbusreq7_p & v372cfc2;
assign v3a7008a = hbusreq7_p & v3a69063 | !hbusreq7_p & v372e479;
assign v3a70c33 = hbusreq5 & v3a642c5 | !hbusreq5 & v376256c;
assign v372b396 = hgrant5_p & v8455ab | !hgrant5_p & v37257cf;
assign v3a692da = hmaster0_p & v375d65c | !hmaster0_p & v3a7074e;
assign v3743b49 = hbusreq8_p & v3a6f15d | !hbusreq8_p & v373f780;
assign v3a6eeb0 = hmaster2_p & v380881d | !hmaster2_p & v3769374;
assign v3a7106d = hbusreq4_p & v3a65fa5 | !hbusreq4_p & v8455ab;
assign v23fe379 = hbusreq3 & c511c2 | !hbusreq3 & v374f609;
assign v3a64879 = hbusreq5_p & v3a70134 | !hbusreq5_p & v372cdef;
assign v372a711 = hlock2_p & v3756416 | !hlock2_p & v3766b11;
assign v3a6ae2f = hmaster0_p & v3750eb9 | !hmaster0_p & v376b540;
assign v3a6daed = hmaster0_p & v372a1b5 | !hmaster0_p & v3775100;
assign v3773089 = hmaster0_p & v3770957 | !hmaster0_p & v3a296d8;
assign v37480f1 = hgrant4_p & v8455ab | !hgrant4_p & v372d10e;
assign v3a6406d = hbusreq6_p & v376ef7a | !hbusreq6_p & v8455b3;
assign v3a641c0 = hmaster0_p & v375139a | !hmaster0_p & !v3a702ce;
assign v3a6046d = hmaster1_p & v3755786 | !hmaster1_p & v3729bd1;
assign v38071a9 = hbusreq6 & v37566b2 | !hbusreq6 & !v8455ab;
assign v3a70577 = hgrant5_p & v3a69fe0 | !hgrant5_p & v375fac2;
assign v375cd0c = hbusreq1 & v3a70641 | !hbusreq1 & v8455ab;
assign cda4f0 = hmaster1_p & v3759031 | !hmaster1_p & v3744da3;
assign v3a5a52a = hgrant2_p & v3739ca8 | !hgrant2_p & v3a6fa5e;
assign v3a6961d = hmaster0_p & v37626ab | !hmaster0_p & v37665e1;
assign v377293c = hgrant6_p & v3a64045 | !hgrant6_p & v37558b4;
assign v37493ed = hbusreq8_p & v37431c0 | !hbusreq8_p & v37681ec;
assign a9f810 = hgrant1_p & v37599b1 | !hgrant1_p & v374e06f;
assign v375c845 = hgrant6_p & v377f09a | !hgrant6_p & v3a70a05;
assign v3a69910 = hmaster1_p & v3807aa1 | !hmaster1_p & v3a70943;
assign v372feb2 = hready & v3a705f6 | !hready & !v8455ab;
assign v3776323 = hgrant4_p & v37692c1 | !hgrant4_p & v3a5ab33;
assign v376147f = hmastlock_p & v3a6ac94 | !hmastlock_p & v8455ab;
assign v3a58bae = hbusreq5 & v376c5d3 | !hbusreq5 & v3730c96;
assign v375242f = hmaster1_p & v3757bac | !hmaster1_p & v3761019;
assign v37728b1 = hbusreq6 & v8455b0 | !hbusreq6 & v3730ffe;
assign a568f8 = hgrant4_p & v3a5e24e | !hgrant4_p & v37584c7;
assign v375a635 = hlock0 & v3a6efea | !hlock0 & v3a56cca;
assign v3762817 = hmaster3_p & v3a551bd | !hmaster3_p & v35b7d97;
assign v3729f3c = hmaster3_p & v8455ab | !hmaster3_p & !v3770891;
assign v37421c0 = hgrant5_p & v8455ab | !hgrant5_p & v3761e59;
assign v3a700ad = hbusreq2 & v3a6106c | !hbusreq2 & v3a713e3;
assign v3753f85 = jx0_p & v3779239 | !jx0_p & v3742358;
assign v3757ae7 = hbusreq3_p & a36a2a | !hbusreq3_p & v3778528;
assign v3a562b7 = hbusreq5 & v3776917 | !hbusreq5 & v37411ab;
assign v373a349 = hlock6 & v377c551 | !hlock6 & v377123e;
assign v374b2f7 = hbusreq6_p & v37349d3 | !hbusreq6_p & v3a5b41c;
assign v3a7028d = hgrant3_p & v3754227 | !hgrant3_p & v3a693af;
assign v3a6eb3e = hmaster0_p & v372be56 | !hmaster0_p & v3726983;
assign v3752b6d = hbusreq7 & v374b867 | !hbusreq7 & v376e66e;
assign v375c883 = hgrant6_p & v374306c | !hgrant6_p & v3a57496;
assign v373b571 = hgrant5_p & v3729720 | !hgrant5_p & v37411c1;
assign v3739311 = hgrant3_p & v8455ab | !hgrant3_p & v37596c8;
assign v37662e2 = hgrant6_p & v3766924 | !hgrant6_p & v375b143;
assign cb0c12 = hmaster1_p & v8455ab | !hmaster1_p & v3762f6e;
assign v2acaed7 = hlock5_p & v3a705cc | !hlock5_p & !v8455ab;
assign v3728373 = hmaster1_p & v3807f45 | !hmaster1_p & v3a60dd5;
assign v37636e3 = hmaster2_p & v377234d | !hmaster2_p & v3a7153c;
assign v372a465 = hmaster0_p & v37402d8 | !hmaster0_p & v377291b;
assign v3768e7e = hbusreq0 & v373ace1 | !hbusreq0 & v375e356;
assign v3745aae = hmaster0_p & v37329ec | !hmaster0_p & v37789ca;
assign v3a5b7e3 = hlock7 & v360d105 | !hlock7 & v3751fbe;
assign v3a704e6 = hbusreq8_p & v3a592bc | !hbusreq8_p & v3a636d2;
assign v3a6e5f0 = hlock4_p & v3755002 | !hlock4_p & !v8455ab;
assign v3766e55 = hbusreq4_p & v357731b | !hbusreq4_p & v3a5bb64;
assign v37302f1 = hbusreq2_p & v3755dcd | !hbusreq2_p & !v3729421;
assign v377a812 = hmaster1_p & v375121b | !hmaster1_p & v3772080;
assign v3a65762 = hbusreq0 & v3a63299 | !hbusreq0 & v373ad16;
assign v37602e0 = hbusreq5 & v377f26e | !hbusreq5 & v375ee2e;
assign bddd83 = hmaster2_p & v37245f8 | !hmaster2_p & !v374e28f;
assign v376c6ba = hmaster2_p & v37600c0 | !hmaster2_p & v3777c59;
assign v1e37ec1 = hlock8 & v373ef28 | !hlock8 & v3a6ccc6;
assign v372b790 = hlock2_p & v9c492b | !hlock2_p & v372c503;
assign v3a66dc0 = hgrant4_p & v3a6f0c9 | !hgrant4_p & v3a579a3;
assign v3731555 = hmaster1_p & v37386f5 | !hmaster1_p & v377c0ad;
assign v3764270 = hlock4 & v3745a81 | !hlock4 & v3a67b48;
assign v3726448 = hmaster1_p & v3a697b9 | !hmaster1_p & v375cfe0;
assign v3a58dac = hbusreq2_p & v3746e4e | !hbusreq2_p & v8455ab;
assign v37280a0 = hbusreq5 & v374cb24 | !hbusreq5 & !v8455ab;
assign v3758972 = hlock2 & v3757271 | !hlock2 & v3a6fd48;
assign v37725e7 = hbusreq6_p & v3a67729 | !hbusreq6_p & v3a5507a;
assign v3a6d499 = hmaster2_p & v3a635ea | !hmaster2_p & v3a641d5;
assign v37376c8 = hbusreq1_p & v3a6fd71 | !hbusreq1_p & v377e2f1;
assign v3731945 = hbusreq2 & v3a6fe46 | !hbusreq2 & v8455ab;
assign v3a61de8 = hlock5_p & v8455ab | !hlock5_p & v3776ada;
assign v377600d = hbusreq5 & v3725b77 | !hbusreq5 & v3a60bfb;
assign v3739239 = hmaster1_p & v376f979 | !hmaster1_p & !v3738eb0;
assign v3a5e537 = hbusreq5 & v3a6fc04 | !hbusreq5 & v8455ab;
assign v376d81a = hbusreq7_p & v380921b | !hbusreq7_p & v376fb37;
assign v3777eed = hlock6 & v3774df9 | !hlock6 & v3770075;
assign v3a69028 = hmaster0_p & v3a5a510 | !hmaster0_p & v375f95f;
assign v3754bc9 = hlock5_p & v3724249 | !hlock5_p & v8f7302;
assign v3a6d809 = hbusreq4_p & v3a557ea | !hbusreq4_p & v3a7131c;
assign v3764ca8 = hbusreq6_p & v38095b2 | !hbusreq6_p & v3769cd6;
assign v372f07d = hmaster2_p & v3759d41 | !hmaster2_p & v372348c;
assign v3a71652 = hlock2_p & v3a70526 | !hlock2_p & !v8455ab;
assign v377bf2b = hbusreq7_p & v374b7ea | !hbusreq7_p & v373e284;
assign v375045d = hbusreq2_p & v3756d07 | !hbusreq2_p & !v8455ab;
assign v3776cbb = hmaster2_p & v3a6fe96 | !hmaster2_p & v37627c3;
assign v374c5e2 = hmaster2_p & v8455ab | !hmaster2_p & v3774a77;
assign v360d07a = hgrant6_p & v3750d06 | !hgrant6_p & v3738419;
assign v3a572bd = hmaster1_p & v3a7069a | !hmaster1_p & v376e2fb;
assign v3a5d21b = hlock5 & v372d773 | !hlock5 & v37690da;
assign da4c01 = hbusreq6_p & v3737c86 | !hbusreq6_p & v3a6b4a6;
assign v3776e23 = hmaster3_p & v376b18f | !hmaster3_p & v37444ae;
assign v3a6f8a7 = hmaster2_p & v373325f | !hmaster2_p & !v3764978;
assign v3a70135 = hmaster0_p & v3a61f4c | !hmaster0_p & v3751925;
assign v3733b4e = hlock4 & v9762fd | !hlock4 & v37615aa;
assign v37673d6 = hbusreq6 & v37705de | !hbusreq6 & v8455ab;
assign v377122d = hbusreq1 & v37482f8 | !hbusreq1 & !v3a703df;
assign v375a8db = hbusreq7 & v3736b93 | !hbusreq7 & v3a56918;
assign v376111d = hburst1 & v372fe05 | !hburst1 & v377903c;
assign v375d4e5 = hgrant6_p & v3a68834 | !hgrant6_p & v3a67983;
assign v373cfd0 = hmaster0_p & v374d4e6 | !hmaster0_p & v3a707f9;
assign v3775100 = hmaster2_p & v3779cd7 | !hmaster2_p & v37290af;
assign v3a551d6 = hlock3_p & v3774710 | !hlock3_p & v372faf1;
assign v3a7056e = hmaster2_p & v8455e7 | !hmaster2_p & v3a54c77;
assign v375f147 = hbusreq0 & v377d1cd | !hbusreq0 & v376604f;
assign v372a696 = hmaster2_p & v3737860 | !hmaster2_p & v3a68b49;
assign v3a5e748 = hbusreq2_p & v376b21a | !hbusreq2_p & v3729d1a;
assign v3a6ff12 = hmaster0_p & v3a7113c | !hmaster0_p & v3755b4e;
assign v3726983 = hmaster2_p & v376ce4d | !hmaster2_p & v3a70bf7;
assign v3725799 = hgrant6_p & v3762502 | !hgrant6_p & v375b2fe;
assign v37748f0 = hbusreq0 & v3a71600 | !hbusreq0 & v3a7045f;
assign v377b4f7 = hbusreq3 & v37675e2 | !hbusreq3 & v8455ab;
assign v377596e = hmaster3_p & v3a6f8b2 | !hmaster3_p & !v376b1ee;
assign v37673e8 = hbusreq7 & v3a6fd36 | !hbusreq7 & !v8455bd;
assign a89e0c = hbusreq6_p & v372d1bf | !hbusreq6_p & v3a5cf22;
assign v380713a = hbusreq3 & v373fe5e | !hbusreq3 & v3a7136f;
assign v374b035 = hbusreq5 & v37295ce | !hbusreq5 & v8455ab;
assign v3778fab = hmaster0_p & a568f8 | !hmaster0_p & v375649a;
assign v376fe68 = hbusreq8_p & v376ae9f | !hbusreq8_p & v374544d;
assign v3771820 = hbusreq8 & v3a645c2 | !hbusreq8 & v3722f60;
assign v37477ca = hgrant6_p & v374530a | !hgrant6_p & !v3a6dddb;
assign v376b3a9 = hready_p & v374094a | !hready_p & v3a70a7b;
assign v376e358 = hbusreq5_p & v374326f | !hbusreq5_p & v3a71133;
assign v3a5971e = hgrant4_p & v3735cb3 | !hgrant4_p & v3a5ec7a;
assign v37409f6 = hmaster2_p & v373b288 | !hmaster2_p & v3748d67;
assign v3a70333 = hmaster1_p & v375345f | !hmaster1_p & !v376a3f5;
assign v3749f51 = hbusreq4 & v373a27c | !hbusreq4 & v8455e7;
assign v37414ed = hlock6_p & v8455ab | !hlock6_p & v373fe5e;
assign b0f188 = hbusreq2_p & v3a635ea | !hbusreq2_p & v377cc27;
assign v3760658 = hbusreq6 & v37386f5 | !hbusreq6 & !v8455b9;
assign v3a70124 = hmaster2_p & v3a5a6e6 | !hmaster2_p & v374e1c3;
assign v375542d = hbusreq4 & v3a6ffca | !hbusreq4 & v8455ab;
assign v373da8d = hlock6_p & v2925c39 | !hlock6_p & !v8455ab;
assign v3a2ae01 = hbusreq2 & v37482f8 | !hbusreq2 & v8455ab;
assign v3a5f7b8 = hmaster2_p & v3a70374 | !hmaster2_p & v3a5b51a;
assign v374b0a8 = hlock3_p & v373ecae | !hlock3_p & v37598c6;
assign v3a6f012 = hmaster0_p & v3776633 | !hmaster0_p & v376730a;
assign v376afdf = hgrant4_p & v8455ab | !hgrant4_p & v39ebb64;
assign v374a369 = hmaster0_p & v3a58bb0 | !hmaster0_p & v3739b7a;
assign v3a71386 = hmaster1_p & v3a5a510 | !hmaster1_p & v3a69028;
assign v373ee19 = hmaster2_p & v3a653e4 | !hmaster2_p & !v37648af;
assign v3a614df = jx1_p & v3a5aef2 | !jx1_p & v375b0f9;
assign v3a57b11 = hgrant8_p & v8455b9 | !hgrant8_p & v3a644d3;
assign v3769758 = hbusreq2 & v3751faf | !hbusreq2 & v8455ab;
assign v3757f96 = hbusreq8 & v372f7b4 | !hbusreq8 & v3775723;
assign v374a2cc = hbusreq6_p & v376c62d | !hbusreq6_p & v8455ab;
assign v1e37579 = hmaster0_p & v377839c | !hmaster0_p & v3a66292;
assign v3a2a13a = hbusreq4_p & v376a96b | !hbusreq4_p & v374cab5;
assign v375725f = hmaster2_p & v8455ab | !hmaster2_p & v8455b6;
assign v380879c = hgrant6_p & v3763fb5 | !hgrant6_p & v3a68255;
assign v3760237 = hbusreq8_p & v3763952 | !hbusreq8_p & v372d525;
assign v3a660e9 = hbusreq2_p & v374f1c3 | !hbusreq2_p & v37720ca;
assign v373d10f = hgrant6_p & v3735dae | !hgrant6_p & v3a6d4f9;
assign v93144b = hbusreq0 & ad3125 | !hbusreq0 & v3722e7a;
assign v3a68315 = hlock5 & v3730722 | !hlock5 & v3a5ed86;
assign v3779014 = hlock7 & v37758de | !hlock7 & v3a6e8db;
assign v3777628 = hmaster2_p & v3a5a807 | !hmaster2_p & v3739ddf;
assign v3747ec9 = hbusreq5 & v3745ab5 | !hbusreq5 & !v8455ab;
assign v3760452 = hmaster2_p & v3a5a6e6 | !hmaster2_p & v376e35e;
assign v37bfcae = hlock3_p & v37502d9 | !hlock3_p & a6f8c7;
assign v373c6a2 = hbusreq3_p & v3775a84 | !hbusreq3_p & v374b383;
assign v3737421 = hbusreq5_p & v3762873 | !hbusreq5_p & v3a5e541;
assign v3a705ac = hbusreq3_p & v37390ff | !hbusreq3_p & !v377b3a8;
assign v37695b1 = hlock0 & v376498f | !hlock0 & v3a6261b;
assign v376bd2f = hgrant5_p & v3a71020 | !hgrant5_p & v37451b6;
assign v376053f = hmaster2_p & v373b166 | !hmaster2_p & v3a65762;
assign v3a62348 = hbusreq6_p & v8455ab | !hbusreq6_p & v3a704c9;
assign v3763f38 = hmaster2_p & v373389a | !hmaster2_p & v377b774;
assign v3a7150d = hlock3_p & v37502b7 | !hlock3_p & v376f9a8;
assign v37728a5 = hbusreq2_p & v3725f4a | !hbusreq2_p & v8455ab;
assign v3744bac = hgrant1_p & v8455ab | !hgrant1_p & v38072fd;
assign v37615aa = hlock6 & v3a66773 | !hlock6 & v3a7025f;
assign v3808eaa = hgrant2_p & v3725475 | !hgrant2_p & v37780f6;
assign v3a70dab = hmaster0_p & v3a70198 | !hmaster0_p & !v373e15b;
assign v3758133 = hgrant4_p & v3a7156d | !hgrant4_p & v3752862;
assign v3a552d2 = hbusreq0 & v3a5bbeb | !hbusreq0 & v3a6bf41;
assign v377a0be = jx0_p & v3a6eb4f | !jx0_p & v37334c2;
assign v3a6eb11 = hmaster0_p & v3a712e2 | !hmaster0_p & v3a6c631;
assign v3760e2e = hbusreq6_p & d3068c | !hbusreq6_p & v377479e;
assign v3753a28 = hburst0 & v3749a12 | !hburst0 & v8455ab;
assign v377add5 = hbusreq2_p & v3a6f5da | !hbusreq2_p & v374d7ce;
assign v3a704f5 = hgrant5_p & v372e537 | !hgrant5_p & v3a5c9d3;
assign v373bb2c = hbusreq4 & v3766117 | !hbusreq4 & v3a70d64;
assign v3a57106 = hmaster2_p & v375946b | !hmaster2_p & v3a6ef5c;
assign v3a7132c = hmaster3_p & v3739d9b | !hmaster3_p & v3734a96;
assign v375ab8e = hlock8 & v3723f45 | !hlock8 & v3a69761;
assign v3755f2d = hmaster1_p & v376e3a0 | !hmaster1_p & v3809390;
assign v375168a = hbusreq0_p & ad2d05 | !hbusreq0_p & v8455b5;
assign v372f1d4 = hmaster2_p & v3a65e3c | !hmaster2_p & v3743de6;
assign v3743d30 = hmaster0_p & v377a121 | !hmaster0_p & v3751004;
assign v3a709e2 = hbusreq3_p & v373dcad | !hbusreq3_p & !v377b3a8;
assign v374fa66 = hmaster1_p & v1e379b9 | !hmaster1_p & !v8455ab;
assign v3a61ff9 = hbusreq5_p & v37647e3 | !hbusreq5_p & v3768551;
assign v3754295 = hlock7 & v3a6bb47 | !hlock7 & v377d428;
assign v37355d6 = hmaster2_p & v372c3d4 | !hmaster2_p & v3730e2a;
assign v3728876 = hmaster1_p & v37245f8 | !hmaster1_p & v373bd3d;
assign v3747467 = hgrant3_p & v374306c | !hgrant3_p & v376e76f;
assign v3a7045c = hgrant0_p & v3a69ac0 | !hgrant0_p & v375803a;
assign v3a5ad83 = hbusreq5_p & v37567ef | !hbusreq5_p & v377c690;
assign v3a6f3f0 = hmaster0_p & v375c432 | !hmaster0_p & v948ef2;
assign v3a571d1 = hmaster0_p & v3a70538 | !hmaster0_p & v37455cd;
assign v3779582 = hgrant2_p & v3a5f50e | !hgrant2_p & v3734465;
assign v377ccbf = hmaster1_p & v376c30b | !hmaster1_p & v8455ab;
assign v3a70b47 = stateG2_p & v8455ab | !stateG2_p & !v3a5cf0b;
assign v3a69c64 = hmaster1_p & v3a6fdd1 | !hmaster1_p & v3771be6;
assign v372a20c = hbusreq3_p & v3809da1 | !hbusreq3_p & v8455ab;
assign v3a70e23 = hgrant0_p & v375c7b9 | !hgrant0_p & !v8455e1;
assign v3776db6 = hgrant2_p & v8455ab | !hgrant2_p & v3737101;
assign v37434d6 = hbusreq3_p & v3759032 | !hbusreq3_p & !v39a537f;
assign v372b445 = hgrant0_p & v377b6ce | !hgrant0_p & !c1a4f5;
assign v23fda2f = stateG2_p & v8455ab | !stateG2_p & v3744037;
assign v373e5fb = hgrant0_p & v8455ab | !hgrant0_p & v377d5d7;
assign v37548e6 = hbusreq6_p & v374d2b3 | !hbusreq6_p & v3a6fd65;
assign v375925f = hbusreq0_p & v3740171 | !hbusreq0_p & v37270d9;
assign v91f9a4 = hbusreq5_p & v375cd8b | !hbusreq5_p & !v8455ab;
assign v374668c = hbusreq6 & v372dd89 | !hbusreq6 & v375b2fe;
assign v3a714b4 = hmaster2_p & v3724394 | !hmaster2_p & v3774bad;
assign v3a70149 = hlock5_p & v3728906 | !hlock5_p & v38072f0;
assign v3a7049e = hmaster0_p & v8455ab | !hmaster0_p & !v37577a4;
assign v3750b9d = hmaster2_p & v373d9e0 | !hmaster2_p & v3727472;
assign v373a8a1 = hmaster1_p & v3a635ea | !hmaster1_p & v3730b15;
assign v375987b = hbusreq3_p & v377b24b | !hbusreq3_p & v3746a04;
assign v3a626a1 = hlock1_p & v374306c | !hlock1_p & v3a6ffae;
assign v373cf8f = hbusreq2 & aa3e48 | !hbusreq2 & v3771e60;
assign v3806bc8 = hlock3 & v337907e | !hlock3 & v3728fb5;
assign v3a6f377 = hlock6 & v3a648d0 | !hlock6 & v3a625f8;
assign v374b9bb = hbusreq8_p & v3777c4e | !hbusreq8_p & v3a701d2;
assign v380911e = hmaster2_p & v3753eb2 | !hmaster2_p & v373891b;
assign v3a69d13 = hgrant6_p & v8455ca | !hgrant6_p & v375b7fa;
assign v3a703b0 = hbusreq5_p & v3733d3f | !hbusreq5_p & v3a6f6c0;
assign v3728916 = hbusreq5_p & v373373d | !hbusreq5_p & !v3729ddd;
assign v374de3d = hbusreq5 & v3a6aea3 | !hbusreq5 & beb41d;
assign v375f354 = hmaster0_p & v8455ab | !hmaster0_p & v375c8c4;
assign v3726699 = hmaster2_p & v3a67a41 | !hmaster2_p & v3a6912a;
assign v377c0ad = hmaster0_p & v37386f5 | !hmaster0_p & v3730878;
assign v3727acb = hmaster2_p & v375a10d | !hmaster2_p & v3a6dc08;
assign v37307a7 = hmaster0_p & v373014d | !hmaster0_p & v3761df7;
assign v3a60bfb = hmaster0_p & v3a71679 | !hmaster0_p & v3a7074e;
assign v3a6fe21 = hgrant6_p & v37604e9 | !hgrant6_p & !v3a70e2a;
assign v3a712d3 = hgrant6_p & v1e37cd6 | !hgrant6_p & v37255de;
assign v3a6ff59 = hbusreq2 & v375af3c | !hbusreq2 & v37c0077;
assign v3745941 = hbusreq8 & v3a60134 | !hbusreq8 & v375075b;
assign v375e444 = hmaster0_p & v3a63198 | !hmaster0_p & v372700a;
assign v3a5e291 = hgrant4_p & v3a6caa5 | !hgrant4_p & !v8455ab;
assign v3a6ffd2 = hlock5_p & v3a71602 | !hlock5_p & v3731d2d;
assign v3776914 = hmaster2_p & v377d107 | !hmaster2_p & v375a94a;
assign v374c9d1 = hbusreq7 & v3a6062e | !hbusreq7 & v3a60276;
assign v373cddc = hgrant4_p & v8455ab | !hgrant4_p & v3a68728;
assign v377dc82 = hmaster0_p & v3730dc4 | !hmaster0_p & v8455ab;
assign v376cbbe = hmaster2_p & v3727976 | !hmaster2_p & !v3a5cfac;
assign v3773f4e = hbusreq6_p & v377aede | !hbusreq6_p & v377eb7a;
assign v3a70b4f = hmaster1_p & v1e382e7 | !hmaster1_p & v3a70e25;
assign v3a680eb = hbusreq5_p & v3739b37 | !hbusreq5_p & v3771171;
assign v3754bb1 = hbusreq0 & v3778572 | !hbusreq0 & v377cf7f;
assign v375c735 = hlock7 & v3a65bb1 | !hlock7 & v377661b;
assign v374fd45 = hbusreq2_p & v37312e2 | !hbusreq2_p & v8455ab;
assign v3a5c9d3 = hmaster1_p & v3759be3 | !hmaster1_p & v3729988;
assign v373d293 = hgrant2_p & v8455ab | !hgrant2_p & v3a558f6;
assign v375f145 = hmaster2_p & v372d299 | !hmaster2_p & v3806ef3;
assign v373ef30 = hbusreq2 & v3755dcd | !hbusreq2 & !v8455bd;
assign v37335e0 = hmaster1_p & v376b7e1 | !hmaster1_p & v3744b87;
assign v376aedb = hgrant6_p & v377ab1f | !hgrant6_p & v377aede;
assign v3a6b90f = hbusreq6 & v3a5bca4 | !hbusreq6 & v3745f9b;
assign v3754a41 = hmaster2_p & v37392ad | !hmaster2_p & !v3a5e544;
assign v3725e96 = hgrant4_p & v8455ab | !hgrant4_p & v3a552d2;
assign v375fe7a = hmaster2_p & v3a70e4f | !hmaster2_p & !v8455bb;
assign v3a641d5 = hbusreq3_p & v3a635ea | !hbusreq3_p & v3a63621;
assign v373fde6 = hbusreq4 & v373a6c8 | !hbusreq4 & v3a6efad;
assign v37316bb = hbusreq4 & v377a35c | !hbusreq4 & v8455ab;
assign v3723555 = hbusreq6_p & v37709bb | !hbusreq6_p & v374a95d;
assign v3a70dbe = hlock6 & v37606ba | !hlock6 & v37672a5;
assign v373c22e = hmaster0_p & v37433f5 | !hmaster0_p & v35b71da;
assign v3731fab = hbusreq5 & v37534da | !hbusreq5 & v37c1a73;
assign v39eb56c = hlock4 & v375a92b | !hlock4 & v373eecc;
assign v375e752 = hbusreq4_p & v3a708ad | !hbusreq4_p & v3a6f310;
assign v3a5b121 = hbusreq6 & v372c60a | !hbusreq6 & v377caa3;
assign v8d4314 = hmaster2_p & v373b0d2 | !hmaster2_p & v372b8fd;
assign v3903ee2 = hmaster2_p & v8455ab | !hmaster2_p & !v8455c9;
assign v3a608fe = hbusreq4 & v35772c9 | !hbusreq4 & v8455ab;
assign v3765b9b = hgrant5_p & v375d98c | !hgrant5_p & v377a9b8;
assign v374e402 = hmaster0_p & v8455b0 | !hmaster0_p & v3a5a01b;
assign v3729e65 = hlock3_p & v3a63e82 | !hlock3_p & !v35772a6;
assign v3a6f113 = locked_p & v377e976 | !locked_p & v3727345;
assign v3729e38 = hbusreq4_p & v37661db | !hbusreq4_p & v375f1ee;
assign v3742c64 = hlock8_p & v37605db | !hlock8_p & v3a54059;
assign v3731115 = hgrant3_p & v37289d4 | !hgrant3_p & v8455ab;
assign v3768a11 = hbusreq5_p & v3724b20 | !hbusreq5_p & !v8455ab;
assign ba83e3 = hmaster2_p & v3738253 | !hmaster2_p & v373ad68;
assign v3766d24 = hmaster2_p & v3740187 | !hmaster2_p & v2ff8cae;
assign v375ca80 = hbusreq8_p & v3a6f794 | !hbusreq8_p & v373f057;
assign v377d1dc = hgrant4_p & v3a53eeb | !hgrant4_p & !v8455ab;
assign v3a55a75 = hmaster0_p & v3737d90 | !hmaster0_p & !v37c0294;
assign v3734b34 = hbusreq4 & v3740171 | !hbusreq4 & v8455ab;
assign v3777ad7 = hmaster2_p & v3a70c39 | !hmaster2_p & v8455ab;
assign v3734ed6 = hmaster1_p & v374306c | !hmaster1_p & v377975f;
assign v3a6eab2 = hmaster1_p & v3725a21 | !hmaster1_p & v373823e;
assign v37777ad = hbusreq4_p & v3a7092a | !hbusreq4_p & v3a6f48b;
assign v3a6fba2 = hbusreq8 & v373e88f | !hbusreq8 & v3a6ae12;
assign v375b282 = hmaster2_p & v3a637dd | !hmaster2_p & !v37326a1;
assign v374b424 = hbusreq3 & v3a6c0b3 | !hbusreq3 & v374cc2a;
assign v3a68787 = hmaster0_p & v376301d | !hmaster0_p & v3a64c71;
assign v3a54271 = jx1_p & v3738d54 | !jx1_p & v3a5c0f8;
assign v3761d7d = hmaster2_p & v3a5b7c2 | !hmaster2_p & !v3a60f71;
assign v3a70c87 = hbusreq5 & v372c6c4 | !hbusreq5 & v3765c08;
assign v37269de = hlock4 & v372f83b | !hlock4 & v376aba9;
assign v3a7005b = hmaster0_p & v3a6c628 | !hmaster0_p & v376ff64;
assign v374a4c2 = hmaster1_p & v376f56d | !hmaster1_p & v37384a9;
assign v3a714c6 = hlock0_p & v3a6c23b | !hlock0_p & v3745075;
assign v372b268 = hbusreq4_p & v3a71467 | !hbusreq4_p & !v376079f;
assign v373a832 = hbusreq7 & v3a6a413 | !hbusreq7 & v3a6cfa1;
assign v376b4e1 = hburst1 & v8455ab | !hburst1 & v373ef4b;
assign v3a70b12 = jx0_p & v3a5fc9c | !jx0_p & v8455ab;
assign v3a7010a = hbusreq7 & v3a5ae9f | !hbusreq7 & v37429c5;
assign v372f23a = hmaster1_p & v3a5b289 | !hmaster1_p & v3a6f674;
assign v3735826 = hgrant1_p & v3a6f2ef | !hgrant1_p & v37764a5;
assign v3750403 = hmaster2_p & v377855f | !hmaster2_p & v3a565ef;
assign v39a4e84 = hgrant6_p & v8455b5 | !hgrant6_p & v3a6f717;
assign v376e31a = hmaster2_p & v3a7151d | !hmaster2_p & !v3723b00;
assign v3779eea = hbusreq0 & v372c3a4 | !hbusreq0 & !v3a6fa19;
assign v37265b8 = hgrant6_p & v3a6ebe6 | !hgrant6_p & v3a6212b;
assign v377817b = hmaster2_p & v3a6fc7f | !hmaster2_p & v3764a2d;
assign v3742584 = hgrant8_p & v376079e | !hgrant8_p & v37673a3;
assign ac9d0d = hlock6 & v373698b | !hlock6 & v3a6199d;
assign b516f2 = hbusreq2 & v377a43e | !hbusreq2 & v37366b5;
assign v3a711fc = hbusreq4 & v3756057 | !hbusreq4 & v3a708c2;
assign v374f8b5 = jx0_p & v3779e21 | !jx0_p & v373ca17;
assign v3a63260 = hbusreq0_p & v375e459 | !hbusreq0_p & v8455ab;
assign v3765c1f = hmaster0_p & v373899b | !hmaster0_p & v3a711e5;
assign v3a6a9cf = stateG10_1_p & v95d97e | !stateG10_1_p & v373a391;
assign v3a71467 = hbusreq0 & v3a53e5b | !hbusreq0 & v8455ab;
assign v3767d4a = hlock7_p & v3a70e87 | !hlock7_p & v8455cb;
assign v373580d = hmaster2_p & v3742cd4 | !hmaster2_p & v3735afb;
assign v3732938 = hmaster2_p & v3a7059b | !hmaster2_p & v38076ec;
assign v3a70bdf = hbusreq8_p & v3a676f1 | !hbusreq8_p & v3a7023d;
assign v377149d = hgrant2_p & v37523f4 | !hgrant2_p & v3733da3;
assign v375d635 = hbusreq1 & v373cca3 | !hbusreq1 & v8455ab;
assign v3a6f73f = hmaster1_p & v3756c2e | !hmaster1_p & v37266a0;
assign v373d107 = hmaster2_p & v3a6b924 | !hmaster2_p & v3a69444;
assign v37464e4 = hmaster2_p & v3a567ec | !hmaster2_p & v3748d67;
assign v3745f9b = hbusreq2_p & v376e041 | !hbusreq2_p & v3748d67;
assign v3775179 = hbusreq6 & v3a58a39 | !hbusreq6 & v8455ab;
assign v377c798 = hlock7 & v3a6332f | !hlock7 & v3776779;
assign v3a60594 = hmaster0_p & v3a60147 | !hmaster0_p & v8455ab;
assign v3a5a6db = hlock3_p & v3778ed4 | !hlock3_p & v8455e7;
assign v37734f8 = hgrant6_p & v373cc5c | !hgrant6_p & v37735cb;
assign v37282cf = locked_p & v3a662f7 | !locked_p & v1e38224;
assign v3722bca = hgrant4_p & v376bb26 | !hgrant4_p & v3735c9d;
assign v3a65212 = hbusreq4 & v376a4d3 | !hbusreq4 & v3a6f07e;
assign v3a6f633 = hmaster2_p & v376eb1d | !hmaster2_p & v3a5bd83;
assign v3757c6f = hmastlock_p & v3a5cf0b | !hmastlock_p & v8455ab;
assign v3a6f5da = hgrant3_p & v8f30ee | !hgrant3_p & v3773aa9;
assign v377d047 = hbusreq2_p & v3a6ffe5 | !hbusreq2_p & v8455ab;
assign v3a62d36 = hgrant3_p & v8455ab | !hgrant3_p & v3a6fb78;
assign v3a6fb64 = hbusreq0_p & v374ab5b | !hbusreq0_p & v3723ac5;
assign v37728d3 = hgrant2_p & v3733d6e | !hgrant2_p & v3a71646;
assign v373f8f8 = hbusreq2_p & v3a69487 | !hbusreq2_p & v375d288;
assign aa6771 = hmastlock_p & v372c42d | !hmastlock_p & !v8455ab;
assign v37756e8 = hlock4_p & v373343b | !hlock4_p & v3741f69;
assign v374f1ae = hgrant6_p & v3a658a9 | !hgrant6_p & v3769c95;
assign v374127d = hbusreq8 & v37596a6 | !hbusreq8 & v37775c7;
assign v3736c97 = hgrant6_p & v8455e7 | !hgrant6_p & v374611e;
assign v373dd9b = hgrant3_p & v3a61a7f | !hgrant3_p & v3a66f81;
assign v3a71073 = hmaster2_p & v8455ab | !hmaster2_p & !v8455b3;
assign v3a67fd9 = hbusreq6 & v3729700 | !hbusreq6 & v37443ab;
assign v3a55aea = hbusreq7_p & v3746877 | !hbusreq7_p & v3777d70;
assign v3769f4e = hmaster0_p & v37435eb | !hmaster0_p & v3769923;
assign v3a60280 = hgrant4_p & v8455ab | !hgrant4_p & v3778754;
assign v374518c = hlock0 & v3a635ea | !hlock0 & v1e37339;
assign v377e3fe = hmaster1_p & v3a6f56b | !hmaster1_p & v377cf71;
assign v372ea2d = hgrant5_p & v375fcab | !hgrant5_p & v37424b8;
assign v3a6b78f = hbusreq5_p & v3a67dd5 | !hbusreq5_p & v3722ac4;
assign v3a5b00a = hlock6_p & v2acb5a2 | !hlock6_p & v3a6ac26;
assign v373adb9 = hbusreq5_p & v3744d2b | !hbusreq5_p & v3a6ca0b;
assign v3739da7 = hgrant2_p & v3735525 | !hgrant2_p & v3a70688;
assign v3756595 = hbusreq8 & v374efad | !hbusreq8 & v3a6f6e0;
assign v3752e29 = hbusreq5 & v374d781 | !hbusreq5 & v8455ab;
assign v3744f48 = hbusreq5 & v3766160 | !hbusreq5 & v3a635ea;
assign v3763d3a = hgrant0_p & d3b3b2 | !hgrant0_p & v374794f;
assign v372c3c0 = hbusreq7 & v3a69329 | !hbusreq7 & v3734ba4;
assign v3a5fe3c = hgrant4_p & v3a5e46d | !hgrant4_p & v3726f38;
assign v3a70791 = hgrant6_p & v372ea4b | !hgrant6_p & v3a57b70;
assign v3731a29 = hbusreq6_p & v372a5c8 | !hbusreq6_p & v372f192;
assign v37650c4 = hbusreq8_p & v37781fe | !hbusreq8_p & v372e47b;
assign v3a6ef56 = hgrant5_p & v3a5d11d | !hgrant5_p & v3a6fa58;
assign v3a70cd6 = hmaster0_p & v3a70209 | !hmaster0_p & v3a6fbad;
assign v377a18b = hlock5 & v3747084 | !hlock5 & v3a6fd98;
assign aab2b0 = hlock0_p & v3740171 | !hlock0_p & v375925f;
assign v3775303 = hbusreq1_p & v3770517 | !hbusreq1_p & v8455ab;
assign v3753eb2 = hgrant4_p & v35b774b | !hgrant4_p & v3735c92;
assign v373497f = hmaster0_p & v373e896 | !hmaster0_p & v3a6108b;
assign v37c0077 = hgrant3_p & v8455ab | !hgrant3_p & v374253f;
assign v37533c8 = hmaster0_p & v3a711ea | !hmaster0_p & !v3a6ff47;
assign v37631bf = hbusreq7_p & v3a704c4 | !hbusreq7_p & v3807472;
assign v373dff9 = hmaster1_p & v372b9c5 | !hmaster1_p & v37485e2;
assign v3a643a0 = hbusreq4_p & v3749cdf | !hbusreq4_p & v3a63938;
assign v37272df = hbusreq4_p & v376d41b | !hbusreq4_p & v3763b0a;
assign v3a7118e = hgrant5_p & v3747454 | !hgrant5_p & v3764678;
assign v373f661 = hgrant1_p & v375d635 | !hgrant1_p & v37764a5;
assign v3775622 = hbusreq7_p & v37761dd | !hbusreq7_p & v376597e;
assign v3767010 = hgrant8_p & v374f535 | !hgrant8_p & v373b0f5;
assign v376babf = hlock5_p & v8455e7 | !hlock5_p & !v3a6ff75;
assign v3743eed = hbusreq8_p & v3a6be07 | !hbusreq8_p & v375b0f9;
assign v3759ce2 = hmaster0_p & v3a70853 | !hmaster0_p & v373d55f;
assign v37438ca = hmaster0_p & v3a71469 | !hmaster0_p & v3a6a1b7;
assign v376dab5 = hgrant2_p & v3a5bb64 | !hgrant2_p & v3724f7b;
assign v375eaac = hbusreq4_p & v3755312 | !hbusreq4_p & v3a611b0;
assign v3a713e2 = hbusreq5 & v3a70987 | !hbusreq5 & v3a64624;
assign v3a7166f = hbusreq5 & v37583f0 | !hbusreq5 & v374c6b8;
assign v376f5e1 = hbusreq3_p & v374af0d | !hbusreq3_p & v3a6255b;
assign v23fde41 = hbusreq7_p & v374ce2a | !hbusreq7_p & v3a67beb;
assign v37416c8 = hbusreq0 & v3770c4c | !hbusreq0 & v39a53a4;
assign v3a68c27 = hlock7 & v3a60443 | !hlock7 & v377b8f9;
assign v3a7140b = hmaster1_p & v3a6f318 | !hmaster1_p & v3a598da;
assign v3a700d9 = hbusreq5 & v3a6f929 | !hbusreq5 & v8455ab;
assign v3a298b6 = hbusreq5_p & v3a614a0 | !hbusreq5_p & v373af26;
assign v3751d98 = hbusreq2_p & v3744983 | !hbusreq2_p & v3a6f386;
assign v374bbaf = hmaster1_p & v3730e7d | !hmaster1_p & v372c483;
assign v37739f4 = hlock4_p & v373fe5e | !hlock4_p & !v8455ab;
assign v373a9ac = hlock5_p & v375eac3 | !hlock5_p & v373cd5d;
assign v37644b7 = hgrant5_p & v8455ab | !hgrant5_p & v37360df;
assign v3a6ebc7 = hbusreq5 & v3258dc5 | !hbusreq5 & v376502e;
assign v3755423 = hmaster1_p & v37640e9 | !hmaster1_p & v37477d3;
assign v37285cd = hmaster1_p & v3767b70 | !hmaster1_p & v8b1055;
assign v377b0f8 = hmaster2_p & v376641b | !hmaster2_p & !v3775bd3;
assign v37247b2 = hbusreq5 & v3a66bc6 | !hbusreq5 & v373cae8;
assign v9d4353 = hmaster1_p & v3a55b39 | !hmaster1_p & v3765cf3;
assign v3a6dd5a = hbusreq0 & v3a645df | !hbusreq0 & v3a6487f;
assign v3a6f292 = hmaster1_p & v3a63fd2 | !hmaster1_p & v3a563c1;
assign v3733173 = hgrant5_p & v37300d3 | !hgrant5_p & v3a6df6c;
assign v37520d9 = hlock5_p & v37638fe | !hlock5_p & v3a59c91;
assign v3378302 = hlock4 & v3725bab | !hlock4 & v3a68601;
assign v375a6d8 = hbusreq7 & v372f99a | !hbusreq7 & v373c5b5;
assign v3a6fcb6 = hmaster2_p & v374729b | !hmaster2_p & v377cfd9;
assign v37453f0 = hbusreq0 & v3a5f0cf | !hbusreq0 & v3a58134;
assign v372cc25 = hbusreq1_p & v37721e6 | !hbusreq1_p & !v8455ab;
assign v3761847 = hmaster1_p & v3a6811a | !hmaster1_p & a52d64;
assign v3753ccf = hbusreq4_p & v8455ab | !hbusreq4_p & v3a6f817;
assign v375f985 = hlock7 & a0a219 | !hlock7 & v37425a8;
assign v375b046 = hmaster0_p & v3769b1d | !hmaster0_p & v3a6ff47;
assign v3722fc0 = hmaster2_p & v372b1dc | !hmaster2_p & !v3a703de;
assign v3a5d923 = hbusreq1_p & v374961f | !hbusreq1_p & !v8455ab;
assign v3a6cd35 = hbusreq4 & v3772c7a | !hbusreq4 & v3a712b1;
assign v3a69487 = hbusreq0_p & v8455e7 | !hbusreq0_p & v8455ab;
assign v37524cf = hmaster0_p & v3735486 | !hmaster0_p & v372c14d;
assign v3754aa8 = hmaster3_p & v3a704cd | !hmaster3_p & v8455ab;
assign v37605a5 = hlock8_p & v372bf1d | !hlock8_p & v35b776e;
assign v37761d1 = hmaster1_p & v3768da7 | !hmaster1_p & v8455ab;
assign v3751069 = hmaster2_p & v3724e8e | !hmaster2_p & v3a5f0b2;
assign v3776abb = hmaster0_p & v3a6ffae | !hmaster0_p & v376c047;
assign v3a704d9 = hgrant0_p & v8455ab | !hgrant0_p & !v374710b;
assign v3742f28 = hlock6_p & v3a56642 | !hlock6_p & adf78a;
assign v373530a = hbusreq6_p & v376c635 | !hbusreq6_p & v372d5bb;
assign v3a70ba7 = hbusreq6 & v3a70ee1 | !hbusreq6 & v373fc8a;
assign v3a6f8af = hgrant6_p & v3806cd2 | !hgrant6_p & v35b9d52;
assign v3a58b5a = hbusreq4 & v376dbdf | !hbusreq4 & v8455ab;
assign v3723e62 = hgrant5_p & v3809eb1 | !hgrant5_p & v3a6cf75;
assign v372d561 = hmaster1_p & v37296a5 | !hmaster1_p & v372dfba;
assign v3807074 = hbusreq5_p & v3a6ca54 | !hbusreq5_p & v8455ab;
assign v3727eca = hbusreq3_p & v3a5d923 | !hbusreq3_p & v3768931;
assign v377b6de = hmaster0_p & v3740893 | !hmaster0_p & v23fe28c;
assign v374b0cb = hgrant4_p & v3770719 | !hgrant4_p & v375e647;
assign v3777647 = hmaster0_p & v376f56d | !hmaster0_p & v37233e4;
assign v3732f03 = hlock4_p & v37474da | !hlock4_p & v377ea59;
assign v3760ab8 = hlock3_p & v3a6d4c2 | !hlock3_p & !v8455ab;
assign d383e7 = hmaster1_p & v3723211 | !hmaster1_p & v3a5bc5f;
assign v377c6b0 = hmaster3_p & v8455ab | !hmaster3_p & !v3a70485;
assign v3736079 = hgrant5_p & v8455ab | !hgrant5_p & !v373f880;
assign v3a5cc3c = hgrant3_p & v337948a | !hgrant3_p & v377c4bd;
assign v374cfee = hgrant4_p & v3a6b19d | !hgrant4_p & v8455ab;
assign v3a5f4ff = hgrant3_p & v8455ab | !hgrant3_p & v373da5b;
assign c60fa0 = hmaster2_p & v3a5c945 | !hmaster2_p & v3759032;
assign v3725058 = hmaster0_p & v376ea64 | !hmaster0_p & v3a5cdc1;
assign v3377c79 = decide_p & v37537cc | !decide_p & v3731f07;
assign v3747a5b = hmaster0_p & v376111d | !hmaster0_p & v37317ec;
assign v3a57959 = hbusreq3_p & v3747302 | !hbusreq3_p & v3a6c5ee;
assign v38072fe = hbusreq5 & v3770367 | !hbusreq5 & v372dd98;
assign v38076ec = hgrant4_p & v3a67403 | !hgrant4_p & v3778d07;
assign v3771607 = hlock4_p & v37453d8 | !hlock4_p & v380974c;
assign v3a59fbc = hbusreq5_p & v2ff87d2 | !hbusreq5_p & v3a60767;
assign v3a6f957 = hmaster2_p & v3a6f7dd | !hmaster2_p & v3a6f4ba;
assign v37646dc = jx3_p & v37311da | !jx3_p & v377c271;
assign v3a708e3 = hmaster2_p & v3a66387 | !hmaster2_p & v3a596c4;
assign v37244f4 = hmaster0_p & v375058e | !hmaster0_p & v3809f27;
assign v3a66651 = hburst1 & v3a6ff41 | !hburst1 & v3755a9f;
assign v3764bee = hlock8_p & v377f883 | !hlock8_p & v35b773b;
assign v3a65fa5 = hbusreq0 & v376a943 | !hbusreq0 & v377ad9c;
assign v3753b7d = hgrant3_p & v3739018 | !hgrant3_p & v3774a8f;
assign v3772d9a = hbusreq3_p & v2619ae8 | !hbusreq3_p & v2acaff4;
assign v3747514 = hbusreq5 & v3a6f6c7 | !hbusreq5 & v373e34e;
assign v3751012 = hmaster1_p & v377caa8 | !hmaster1_p & v376314e;
assign v375cbdf = hbusreq6_p & v3a6ac60 | !hbusreq6_p & v372d851;
assign v374214d = hmaster1_p & v8455b3 | !hmaster1_p & v3724926;
assign v3a679fd = hbusreq7 & v374d612 | !hbusreq7 & v35b71fc;
assign v3740e9c = hbusreq7_p & v3a713a9 | !hbusreq7_p & v3a57b00;
assign v375a166 = hgrant6_p & v8455ab | !hgrant6_p & v1e37dfd;
assign v3a6eb62 = hbusreq3_p & v3a6f7f0 | !hbusreq3_p & v3a618b7;
assign v3a6fa78 = hgrant4_p & v8455ab | !hgrant4_p & v3a6aee6;
assign v3724715 = hlock4 & v8e6c5f | !hlock4 & v3a70480;
assign v3740415 = locked_p & v374aa73 | !locked_p & v8455ab;
assign v377d377 = hbusreq0 & v3a6f616 | !hbusreq0 & v3735293;
assign v3766853 = hmaster1_p & v376bd2c | !hmaster1_p & v37733d9;
assign v3a70318 = hmaster2_p & v375fbf2 | !hmaster2_p & !v3a71330;
assign v3a5afe8 = hbusreq2 & v3733471 | !hbusreq2 & v8455ab;
assign v3a6e463 = hbusreq3_p & v377af98 | !hbusreq3_p & v3a693af;
assign v3809a58 = hlock0 & v37496fa | !hlock0 & v3753f0d;
assign v3a6f7d4 = jx3_p & v374ee76 | !jx3_p & v372bccc;
assign v376ed1f = hgrant2_p & v8455ab | !hgrant2_p & v3a6fed2;
assign v373109c = hbusreq0 & v377293c | !hbusreq0 & v3a70566;
assign v3776b9a = hbusreq6 & v3a5b289 | !hbusreq6 & v8455bb;
assign v37784ad = hbusreq4_p & v376085a | !hbusreq4_p & v3743b9e;
assign v373e873 = hmaster0_p & v37409f6 | !hmaster0_p & v37458ca;
assign v3a5d2a6 = hmaster0_p & v3a606b7 | !hmaster0_p & v373d4a6;
assign v3a5a39f = hmaster2_p & v3777b2e | !hmaster2_p & !v373d2bd;
assign v3a63df6 = hbusreq6_p & v3737c86 | !hbusreq6_p & v3808870;
assign v29256ae = hbusreq2 & v3762cc4 | !hbusreq2 & v38072fd;
assign v3a5b819 = hgrant5_p & v3727626 | !hgrant5_p & v3a6fc33;
assign v376d876 = hbusreq5_p & v3a556ab | !hbusreq5_p & v373cde5;
assign v374b08d = hmaster1_p & v375b48b | !hmaster1_p & v8455e7;
assign v374c2b4 = hbusreq3 & v3755002 | !hbusreq3 & v8455ab;
assign v3a66ad2 = hbusreq7 & v3a6b1b9 | !hbusreq7 & v969d5b;
assign v375a32c = hbusreq4 & bbab81 | !hbusreq4 & v8455ab;
assign v372cc3d = hbusreq8_p & v377444e | !hbusreq8_p & v373fb40;
assign v3728ee0 = hbusreq4 & v372fd0a | !hbusreq4 & !v8455ab;
assign v3728eeb = hbusreq2 & v39a5381 | !hbusreq2 & v8455ab;
assign v3774253 = hmaster3_p & v8455ab | !hmaster3_p & v3a6fee3;
assign v3743522 = hmaster2_p & v35772a5 | !hmaster2_p & !v3a70410;
assign v3746676 = hbusreq7_p & v3a5ccab | !hbusreq7_p & v3a6f684;
assign v37654e7 = hbusreq5 & v39eb413 | !hbusreq5 & v8455ab;
assign v3764703 = hgrant6_p & v3729f14 | !hgrant6_p & v3a70074;
assign v3a6db2d = hmaster2_p & v374306c | !hmaster2_p & v3722e5c;
assign v3752e13 = hbusreq2_p & v375bfd5 | !hbusreq2_p & v3a64d60;
assign v375b320 = hlock5 & v37349f9 | !hlock5 & v37560ef;
assign v376bbe8 = hbusreq1_p & v3764ba8 | !hbusreq1_p & !v8455ab;
assign v37658d9 = hbusreq5_p & v3a62b13 | !hbusreq5_p & v3a70650;
assign v3754c0e = stateG10_1_p & v35772a6 | !stateG10_1_p & v372d593;
assign v3a5f6d5 = hgrant4_p & v3727b03 | !hgrant4_p & v3a5794d;
assign v3750f8f = hlock6 & v3729531 | !hlock6 & v3733727;
assign v3760f87 = hbusreq1_p & v375984e | !hbusreq1_p & v8455ab;
assign v3a6911d = hgrant4_p & v8455ab | !hgrant4_p & v3a70850;
assign v3754d3a = hgrant4_p & v1e37d8b | !hgrant4_p & v3758187;
assign v375bde1 = hbusreq4_p & v3a6233b | !hbusreq4_p & v3a5907a;
assign v373fc07 = hbusreq4 & v374e64f | !hbusreq4 & !v8455b9;
assign v374fe9d = hmaster2_p & v3733da4 | !hmaster2_p & v3a6f4c7;
assign v89a228 = hmaster0_p & v372d842 | !hmaster0_p & v3a5cf5e;
assign v3a615c7 = hbusreq7 & v3a5bed2 | !hbusreq7 & v3a59ddc;
assign v3a62da7 = hlock8_p & v374183f | !hlock8_p & v3a6eee2;
assign v375cdd7 = hlock6_p & v37757e0 | !hlock6_p & v3a57309;
assign v3a64612 = hbusreq5 & v3779680 | !hbusreq5 & v380760a;
assign v37362ea = hgrant1_p & v373a66d | !hgrant1_p & v8455e7;
assign v3a6ca15 = hbusreq4_p & v374df64 | !hbusreq4_p & v2092abe;
assign v3730926 = hbusreq6_p & v3748e0b | !hbusreq6_p & v377a901;
assign v3a62846 = hmaster2_p & v372af77 | !hmaster2_p & v377e889;
assign c51df8 = hlock0_p & v374362e | !hlock0_p & v360bb9f;
assign v3a5e000 = hmaster0_p & v376f5d9 | !hmaster0_p & !v377e004;
assign v3742a8e = hbusreq7 & v3a70d36 | !hbusreq7 & v374a4cc;
assign v376ef09 = hgrant6_p & v377eaf2 | !hgrant6_p & v8455ab;
assign v377db1f = hlock4 & v377723a | !hlock4 & v3769a1e;
assign v3773fdc = hbusreq1_p & v337793f | !hbusreq1_p & !v8455ab;
assign v373227a = hgrant4_p & v3a70929 | !hgrant4_p & b6ae10;
assign v3a5cd53 = hbusreq4_p & v3a56c6d | !hbusreq4_p & v3770163;
assign v3767fd7 = hmaster1_p & v37475d9 | !hmaster1_p & v376f051;
assign v3a71609 = hmaster2_p & v376d5a7 | !hmaster2_p & v377b8ee;
assign v3776f07 = hmaster2_p & v3762034 | !hmaster2_p & v37283ff;
assign v3a6d665 = hlock8 & v376d4d9 | !hlock8 & v3a6ccfe;
assign v3a6eca6 = hmaster1_p & v3750ff0 | !hmaster1_p & v3726da1;
assign v3a70912 = hbusreq4_p & v3a59b8a | !hbusreq4_p & v377aa7a;
assign v375dcf8 = hgrant7_p & v377f5c9 | !hgrant7_p & v3a709ce;
assign v3a68fd3 = hbusreq4_p & v372e669 | !hbusreq4_p & v3a67588;
assign v3727f68 = hbusreq5 & v3a61714 | !hbusreq5 & v3a5f5f5;
assign v376373e = hgrant5_p & v3a6e8b1 | !hgrant5_p & !v8455ab;
assign v3a6f67e = hbusreq2_p & v372e61a | !hbusreq2_p & v37749bf;
assign v3a67ee6 = hbusreq0 & c3d672 | !hbusreq0 & v375cb83;
assign v3763aec = hbusreq0 & v3a713ae | !hbusreq0 & v3a6817a;
assign v37617b9 = hbusreq5_p & v37460de | !hbusreq5_p & !v8455ab;
assign v3a663c3 = hgrant4_p & v8455e7 | !hgrant4_p & v372ed34;
assign v3774cc2 = hbusreq5_p & v3a67bbd | !hbusreq5_p & v3732688;
assign v3a63fe2 = hbusreq5_p & v3762cd8 | !hbusreq5_p & !v8455ab;
assign v3742ecd = hbusreq7_p & v375ae53 | !hbusreq7_p & !v8455ab;
assign v37350c3 = hmaster0_p & v3a58218 | !hmaster0_p & v3730fc4;
assign v3741714 = hbusreq8_p & v375595c | !hbusreq8_p & v372b2b4;
assign v337901e = hbusreq2 & v3748f48 | !hbusreq2 & v8455ab;
assign v3763fb5 = hlock6 & v376f47f | !hlock6 & v37639c6;
assign v38073be = hgrant4_p & v37283bb | !hgrant4_p & v3778f6c;
assign v292556b = hmaster0_p & v3756f8a | !hmaster0_p & v3742851;
assign v3a6ff1a = hgrant6_p & v3743cd6 | !hgrant6_p & v376bb27;
assign v3743fee = jx0_p & v375961b | !jx0_p & v3772d8b;
assign v3735051 = hlock4 & v3a71054 | !hlock4 & v3763fb5;
assign v3a70188 = hlock6 & v3744adf | !hlock6 & v374401a;
assign v3a702e3 = hmaster1_p & v3a635ea | !hmaster1_p & v3750b29;
assign v372eeee = hbusreq6 & v37638ee | !hbusreq6 & v3a70c74;
assign v375c8e8 = hlock3_p & v3a6b9e8 | !hlock3_p & v3732aca;
assign a0cf3e = hbusreq4_p & v3a70a7d | !hbusreq4_p & v377422b;
assign v3765dda = hgrant6_p & v3a59c87 | !hgrant6_p & v377c32f;
assign v376be2c = hbusreq3 & v3a66b2b | !hbusreq3 & v373f0ee;
assign v37451f8 = hbusreq6_p & v375bc08 | !hbusreq6_p & v3a2981e;
assign v37670dd = hmaster1_p & v3762153 | !hmaster1_p & v3a6d2d3;
assign v377b8f9 = hgrant5_p & v373e07e | !hgrant5_p & v3a5f05e;
assign v37639fa = hmaster1_p & v3a670fb | !hmaster1_p & v3779ac0;
assign v377b0a0 = hgrant6_p & v8455ab | !hgrant6_p & v37640fd;
assign v3a62c0a = hmaster2_p & v3724e8e | !hmaster2_p & v8455ab;
assign v3761e19 = hbusreq4_p & v3a53f42 | !hbusreq4_p & v374df4b;
assign v374c251 = hmaster2_p & v3759c1f | !hmaster2_p & v3755b56;
assign v3a62628 = hlock2_p & v3a5b5d3 | !hlock2_p & v3a658bf;
assign v376342f = hmaster2_p & v37728a5 | !hmaster2_p & v3729f14;
assign v3a70dfc = hbusreq5 & v3a70540 | !hbusreq5 & v373b7b5;
assign v374cbe3 = hbusreq6_p & v376f56d | !hbusreq6_p & v37697fc;
assign v3a6e327 = hlock2_p & v377e586 | !hlock2_p & v37c0297;
assign v3777bf4 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3757e40;
assign v3754fb0 = hgrant4_p & v8455ab | !hgrant4_p & v377ec1c;
assign v373574c = hgrant4_p & v2ff87b0 | !hgrant4_p & v375b2d9;
assign v3a5c3eb = hlock5 & v3744f48 | !hlock5 & v3725bba;
assign v3a6f54f = hmaster1_p & v375fb00 | !hmaster1_p & !v374554d;
assign v3a701c6 = hmaster2_p & v3a5ef5c | !hmaster2_p & !v3730e2a;
assign v37781a8 = hlock0 & v38072fd | !hlock0 & v3a6512b;
assign v3a65565 = hbusreq5 & v37735b8 | !hbusreq5 & !v3745bbe;
assign v3a71523 = hbusreq8_p & v372c470 | !hbusreq8_p & v377371c;
assign v3757fcc = hgrant3_p & v8455ab | !hgrant3_p & v3a640c5;
assign v3a70f10 = hbusreq5_p & v37377cf | !hbusreq5_p & v3766e31;
assign v3a7006c = locked_p & v373eef7 | !locked_p & v3a5e24e;
assign v3750b03 = hgrant6_p & v377b6ce | !hgrant6_p & v3733234;
assign v3775aa7 = hmaster2_p & v377834b | !hmaster2_p & v3a5a158;
assign v372ca44 = hbusreq3_p & v376f768 | !hbusreq3_p & v376bb26;
assign v3a6651d = hlock0 & v3a7162d | !hlock0 & v3a56d86;
assign v3a6b70e = hbusreq4 & v37659e2 | !hbusreq4 & v376c76d;
assign v3a5dab7 = hgrant5_p & v37518c9 | !hgrant5_p & v374366a;
assign v3a6108b = hmaster2_p & v3a6fc78 | !hmaster2_p & v3a5bd99;
assign v376fc36 = hlock3 & v3a6f0cc | !hlock3 & v377d705;
assign v37482bb = hbusreq5 & v373a822 | !hbusreq5 & b5da28;
assign v3a6a720 = jx0_p & a0a219 | !jx0_p & v3808e56;
assign v376b600 = hlock6_p & v3735e39 | !hlock6_p & v376d856;
assign v3a5b7c2 = hbusreq6 & v376b4e1 | !hbusreq6 & !v8455ab;
assign v374b0e3 = hbusreq7_p & v3a6cd48 | !hbusreq7_p & v3a5a884;
assign v23fdf85 = hgrant3_p & v3747e8e | !hgrant3_p & v37251f6;
assign v372a79f = hlock4 & v3a679e7 | !hlock4 & v37775f9;
assign v37693af = hbusreq6_p & v3a5beb6 | !hbusreq6_p & v8455b0;
assign v375af43 = hbusreq0 & v3a617b4 | !hbusreq0 & v8455ab;
assign v3742101 = hlock0_p & v372dadb | !hlock0_p & v3a6ebf0;
assign v3758824 = hbusreq6_p & v3a6b710 | !hbusreq6_p & v3a5c210;
assign v3a585f5 = hgrant7_p & v3758fae | !hgrant7_p & v374d6b5;
assign v3a6fa11 = hbusreq5_p & v3a709ee | !hbusreq5_p & v377c7ae;
assign v3a6eace = hgrant5_p & v3a6ffce | !hgrant5_p & v3728ae9;
assign v372ffaa = hbusreq6_p & v8c8903 | !hbusreq6_p & v3a6ffae;
assign v3775a4a = hbusreq4 & v375b02a | !hbusreq4 & v3763104;
assign d27e8c = hgrant6_p & v3a6a213 | !hgrant6_p & v3775311;
assign v372d9ae = hmaster2_p & v3a63408 | !hmaster2_p & v374bb9c;
assign v37469ba = hbusreq5_p & v3a702d8 | !hbusreq5_p & v8455ab;
assign v3764049 = hbusreq4_p & v37639b1 | !hbusreq4_p & v3a682f0;
assign v3a62cff = hbusreq4_p & v37bfc8c | !hbusreq4_p & v37770c9;
assign v375a901 = hbusreq3_p & v3776615 | !hbusreq3_p & v3a6f483;
assign v3774a1b = jx0_p & v3737ca2 | !jx0_p & v37639a1;
assign v3a54d25 = hbusreq7 & v3a70129 | !hbusreq7 & v3737808;
assign v37c36bf = hmaster0_p & v3a635ea | !hmaster0_p & v3736eff;
assign v3a5414c = hbusreq5 & v3a6fda1 | !hbusreq5 & v372a465;
assign v37624a9 = hmaster3_p & v3a6ec29 | !hmaster3_p & v3726b63;
assign a69e17 = hgrant2_p & v3a5f50e | !hgrant2_p & v3a6ef74;
assign v377eed2 = hbusreq8_p & v373eeed | !hbusreq8_p & v3a6f227;
assign v3a5fc3c = hlock2_p & v3745993 | !hlock2_p & v3a669ae;
assign v3a6dc33 = hlock6_p & v3742122 | !hlock6_p & v373f058;
assign v3a61c80 = hlock5 & v3a626fe | !hlock5 & v377b0d8;
assign v376f2a7 = hlock6 & v3776125 | !hlock6 & v3755a0f;
assign v3769c95 = hbusreq6_p & v3a70988 | !hbusreq6_p & v1e37a04;
assign v37470c6 = hbusreq5_p & v3740d32 | !hbusreq5_p & v8455ab;
assign v3a70e7a = hbusreq8 & v374a0c4 | !hbusreq8 & v375295a;
assign v3a669ac = hbusreq3_p & v374f0c1 | !hbusreq3_p & v374e248;
assign v376c4fd = hbusreq7_p & v377bcfc | !hbusreq7_p & !v3a5e74c;
assign v3a70f6b = hgrant6_p & v8455ab | !hgrant6_p & v3a5be6a;
assign v37726d9 = hbusreq8 & v8455e7 | !hbusreq8 & v38076b7;
assign v3a5cfd9 = hbusreq0_p & v373be25 | !hbusreq0_p & !v372935c;
assign v3a7092b = jx3_p & v2ff8ee1 | !jx3_p & v3a6ec1b;
assign v3770eeb = hbusreq5_p & v3a70f9a | !hbusreq5_p & v3a6f235;
assign v3a61462 = hlock5_p & v37597c4 | !hlock5_p & v3725a73;
assign v3777474 = hmaster1_p & v3a57f59 | !hmaster1_p & v3766d53;
assign v3a6fe52 = hbusreq0 & v37420e2 | !hbusreq0 & v3741218;
assign v3753a8a = jx2_p & v377e7f8 | !jx2_p & !v372b2cb;
assign v3a5faf0 = hlock7 & v3737a8b | !hlock7 & v377bf7b;
assign v3a6c016 = hmaster0_p & v377bb3a | !hmaster0_p & v3a70222;
assign v3736e06 = hlock0 & v3a67cff | !hlock0 & v37239ed;
assign v3761932 = hlock3_p & v3a584bf | !hlock3_p & v37331b5;
assign v373cf3a = hbusreq2 & v325c976 | !hbusreq2 & v3a5b614;
assign v3a712de = hgrant2_p & v3a70dc4 | !hgrant2_p & v377e14d;
assign v375fac6 = hbusreq6_p & v3a7063c | !hbusreq6_p & !v3a56cdb;
assign v372c046 = hgrant7_p & v8455ab | !hgrant7_p & v8455cd;
assign v373f0ee = hlock0_p & v3a635ea | !hlock0_p & !v3807a92;
assign v3a6de03 = hbusreq4_p & v376d509 | !hbusreq4_p & v3723ace;
assign v3a707cc = hbusreq5_p & v3745d14 | !hbusreq5_p & !v37787ce;
assign v3a6fa44 = hmaster0_p & v374838d | !hmaster0_p & v3a583b0;
assign v3741bd8 = hbusreq5 & v33789ef | !hbusreq5 & bb70de;
assign v37419f2 = jx0_p & v3a6ec0e | !jx0_p & ade6f1;
assign v3755abd = hgrant6_p & v8455ab | !hgrant6_p & v374dc53;
assign b7df2b = hgrant6_p & v8455ab | !hgrant6_p & v3774add;
assign v3765c35 = hmaster2_p & v3a6f7b0 | !hmaster2_p & a34d2b;
assign v3a71674 = hmaster0_p & v374089d | !hmaster0_p & !v3770fa1;
assign v3806db7 = hready & v3a690ec | !hready & v373fe5e;
assign v3a70657 = jx0_p & v3a64eb3 | !jx0_p & v37247c8;
assign v3734c3a = hbusreq5_p & v3737bfb | !hbusreq5_p & v374fb02;
assign v3a60223 = hlock7 & v3a555a9 | !hlock7 & v3a6f474;
assign v3a6fb81 = hmaster2_p & v3725b27 | !hmaster2_p & v37778a2;
assign v375e21d = hlock7_p & v3a6f470 | !hlock7_p & v3739f49;
assign v37411df = hbusreq6_p & v374c1a9 | !hbusreq6_p & v3a593bb;
assign v3a6bb56 = hbusreq7 & v376f71a | !hbusreq7 & !v3a6f916;
assign v3a6eb5b = jx1_p & v3a71286 | !jx1_p & v8455ab;
assign v374b60b = hgrant6_p & v3738be9 | !hgrant6_p & v3a70bfa;
assign v373285a = hmaster1_p & v377b456 | !hmaster1_p & v372bd2b;
assign v3756531 = hbusreq8_p & v372760c | !hbusreq8_p & v3743b11;
assign v3a64dc2 = hbusreq4 & v3a6a129 | !hbusreq4 & v8455ab;
assign v375df5e = hlock5 & v3740d9a | !hlock5 & v3740975;
assign v3a6b710 = hgrant2_p & v3768b99 | !hgrant2_p & !v3a6fdf8;
assign v37522d3 = hbusreq2_p & v3a71417 | !hbusreq2_p & v8455ab;
assign v3a64058 = hbusreq7 & v377ab6b | !hbusreq7 & v375ccf3;
assign v376d509 = hbusreq4 & v37639c3 | !hbusreq4 & v37770c9;
assign v37403e5 = hbusreq2 & v37273c2 | !hbusreq2 & v8455ab;
assign v373a58c = hmaster1_p & v37293c3 | !hmaster1_p & !v8455ab;
assign v372825b = hbusreq6_p & b1ca9b | !hbusreq6_p & v3743256;
assign v3725589 = hmaster2_p & v8455ab | !hmaster2_p & v3746cc5;
assign v3775610 = hmaster0_p & v3a5b8b9 | !hmaster0_p & v377918a;
assign v375705a = hmaster0_p & v3779183 | !hmaster0_p & v377dbd7;
assign v3a61b9c = hbusreq4_p & v3778572 | !hbusreq4_p & v360d048;
assign v3a70fbb = hbusreq1 & v3a6f018 | !hbusreq1 & !v3a5db8a;
assign v372ee20 = hbusreq5 & v377a337 | !hbusreq5 & v8455ab;
assign v3774e9d = hmaster3_p & v3a702fd | !hmaster3_p & v377168f;
assign v3a5b615 = hbusreq5 & v3a65c31 | !hbusreq5 & !v8455bd;
assign v3a71097 = hbusreq5 & v372a22d | !hbusreq5 & v8455ab;
assign stateG10_2 = !v31461d5;
assign v3736eee = hmaster2_p & v377d1a3 | !hmaster2_p & !v374a2cc;
assign v375961b = hgrant5_p & v8455c6 | !hgrant5_p & v3a6fc5e;
assign v3770517 = hlock1_p & v375cd0c | !hlock1_p & v8455ab;
assign v3a68707 = hmaster1_p & v8455ab | !hmaster1_p & v373d661;
assign v37725ea = hbusreq4 & v376f56d | !hbusreq4 & !v8455ab;
assign v3a6b860 = hbusreq0 & v3a6fdc3 | !hbusreq0 & v8455ab;
assign v3727a10 = hbusreq5_p & v3755cf7 | !hbusreq5_p & v377a8dc;
assign v3762712 = hlock7 & v3731be2 | !hlock7 & v3731bd7;
assign v3a61f85 = hmaster0_p & v3a5f02e | !hmaster0_p & v37793b9;
assign v3807740 = hbusreq2_p & v3727703 | !hbusreq2_p & v3a6a82a;
assign v3741c91 = hmaster2_p & v3741384 | !hmaster2_p & v37350f9;
assign v3a6fc65 = hbusreq1 & v377ba55 | !hbusreq1 & v3724940;
assign v3731f35 = hmaster1_p & ca2eb2 | !hmaster1_p & v8455ab;
assign v3a5f9e6 = hgrant6_p & v8455ab | !hgrant6_p & v377728d;
assign v8455f3 = hgrant5_p & v8455ab | !hgrant5_p & !v8455ab;
assign v372984e = hmaster2_p & v377bfc0 | !hmaster2_p & v3745f9b;
assign v37645bc = hmaster0_p & v38097ee | !hmaster0_p & v8455b0;
assign v3a65e52 = hgrant2_p & v3a632f4 | !hgrant2_p & v37331ef;
assign v373bf79 = hbusreq4 & v37356f0 | !hbusreq4 & v8455ab;
assign v3775b30 = hgrant6_p & v8455ca | !hgrant6_p & v3762545;
assign v3a626ea = hgrant3_p & v8455ab | !hgrant3_p & v3775ee8;
assign v3a552f7 = hbusreq4 & v3a59dab | !hbusreq4 & v375cf36;
assign v3769d07 = hbusreq5 & v3738365 | !hbusreq5 & !v3a6f2c2;
assign v372c1bb = hlock7 & v3a66ea0 | !hlock7 & v376a06c;
assign v3a704ee = hgrant2_p & v372d3e8 | !hgrant2_p & v3a6f22f;
assign v3a5f147 = hbusreq0_p & v3750d37 | !hbusreq0_p & !v3732dc6;
assign v3a6cf6a = hbusreq2_p & v3753f1a | !hbusreq2_p & !v8455ab;
assign v374a4ca = hbusreq4 & v3756483 | !hbusreq4 & v38073c9;
assign v3a7119d = hmaster0_p & v377c9b1 | !hmaster0_p & v376bae4;
assign v3729a69 = hmaster2_p & v377c7c0 | !hmaster2_p & v377b774;
assign v3765ded = hgrant8_p & v3a56804 | !hgrant8_p & v3a68e41;
assign v376a8ee = hbusreq4 & v8455b0 | !hbusreq4 & v3a6fd81;
assign v373dfb5 = hbusreq4_p & v3a5aacb | !hbusreq4_p & v3735c9d;
assign v3a702c1 = hbusreq4_p & v35b6a6b | !hbusreq4_p & v375eb56;
assign v3a6fbd8 = hlock6_p & d99853 | !hlock6_p & !v8455ab;
assign v3a6074d = hbusreq4_p & v3723430 | !hbusreq4_p & v8455e7;
assign v3730e7d = hbusreq3_p & v3761c4e | !hbusreq3_p & v8455ab;
assign v3a65521 = jx0_p & v3739d69 | !jx0_p & v377da08;
assign v3a6f742 = hbusreq2_p & v3754272 | !hbusreq2_p & !v8455ab;
assign v3a59eab = hbusreq7 & v3a587a1 | !hbusreq7 & v372d811;
assign v3771102 = hgrant4_p & v376f449 | !hgrant4_p & v3a70bf7;
assign v374700b = hbusreq4_p & v374b15d | !hbusreq4_p & v3728957;
assign v3778e46 = hmaster1_p & v374f44c | !hmaster1_p & v8455ab;
assign v37493b4 = hmaster0_p & v3a64421 | !hmaster0_p & v37297ce;
assign v375baed = hgrant3_p & v8455ab | !hgrant3_p & v3a6df5a;
assign v3740627 = hmaster2_p & v3a6fcb0 | !hmaster2_p & v8455ab;
assign v37458ca = hmaster2_p & v373b7c5 | !hmaster2_p & v3725717;
assign v37528d5 = hgrant4_p & v3a53eeb | !hgrant4_p & v3742db5;
assign v37403cf = busreq_p & v377f4bb | !busreq_p & !v3749e1c;
assign v37385d2 = hgrant4_p & v372bf24 | !hgrant4_p & v8455ab;
assign v3724aa4 = hmaster1_p & v37641b8 | !hmaster1_p & v3a704d6;
assign v3a610da = hmaster0_p & v37729bf | !hmaster0_p & !v373197c;
assign v3a6f874 = hbusreq4_p & v372ac3b | !hbusreq4_p & v3a5fc8d;
assign v3a65a0f = hmaster0_p & v377700a | !hmaster0_p & v2ff8e8b;
assign v374a2b5 = hbusreq7_p & v37343d1 | !hbusreq7_p & v3743df6;
assign v37451ad = hbusreq4 & v8455b0 | !hbusreq4 & adf78a;
assign v375636e = hbusreq5 & aed6c7 | !hbusreq5 & !v374f9cc;
assign v3a7165c = hbusreq4 & v376beb4 | !hbusreq4 & v3a70a7f;
assign v3a70e5f = jx1_p & v3728bd6 | !jx1_p & v8455ab;
assign v376fd05 = hlock0_p & v3776aa8 | !hlock0_p & v8455ab;
assign v3732b3a = hmaster1_p & v3a70221 | !hmaster1_p & v376ce55;
assign v380775e = stateA1_p & v8455ab | !stateA1_p & !v3a5a225;
assign v37273f6 = hmaster0_p & v375e944 | !hmaster0_p & !v37280f3;
assign v37678bd = hmaster0_p & v3a700ce | !hmaster0_p & !v3a6607f;
assign b68bf2 = hgrant4_p & v8455ab | !hgrant4_p & v377fabb;
assign v374a289 = hmaster1_p & v3a6793d | !hmaster1_p & v37402ee;
assign b8ed55 = hbusreq7_p & v3a70b43 | !hbusreq7_p & v37572b6;
assign v372b163 = hbusreq2_p & v3750d37 | !hbusreq2_p & !v3732dc6;
assign v374c73d = hmaster0_p & v3757343 | !hmaster0_p & v8455ab;
assign v373cde7 = hmaster2_p & v3a6f2e1 | !hmaster2_p & v3a5c5f4;
assign v375b812 = hbusreq5_p & v3a6f790 | !hbusreq5_p & v3a5db06;
assign v3a6e29d = hlock8 & v3774a4b | !hlock8 & v37515a1;
assign v374c74f = hgrant4_p & v3a5b5d3 | !hgrant4_p & v3a5ef3e;
assign v3a7097f = hbusreq5_p & v37299dc | !hbusreq5_p & v3a6e08c;
assign v3759aca = hmaster0_p & v3747931 | !hmaster0_p & v375119e;
assign v3741aca = hbusreq4 & v37626d5 | !hbusreq4 & v8455ab;
assign v3740187 = hgrant4_p & v3a6425d | !hgrant4_p & !v8fc6a0;
assign v372599c = hgrant2_p & v8455e7 | !hgrant2_p & !v376064b;
assign v3a5be57 = hbusreq6_p & v37522d3 | !hbusreq6_p & v372ff72;
assign v372689b = hbusreq4_p & v37c006d | !hbusreq4_p & v8455b7;
assign v3735512 = hbusreq1_p & v3a7162d | !hbusreq1_p & v3778528;
assign v377e52e = hbusreq1 & v37282cf | !hbusreq1 & v37674c1;
assign v3a5949f = hbusreq5 & v377f579 | !hbusreq5 & v3a58c07;
assign v3a6ed14 = hmaster1_p & v3a6f1bf | !hmaster1_p & v3a5744d;
assign v3a70be7 = hmaster2_p & v3770754 | !hmaster2_p & v3a5db97;
assign v39ea663 = hmaster0_p & v376a2c0 | !hmaster0_p & v1e3773a;
assign v3728eef = hbusreq2_p & v3759b2f | !hbusreq2_p & !v373be25;
assign v3a7024b = hbusreq4 & v325b5fd | !hbusreq4 & v375556d;
assign v372580c = hmaster1_p & v377cc6d | !hmaster1_p & v374bc63;
assign v3a5a615 = hlock5 & v3a6add2 | !hlock5 & v3a6225d;
assign v3a579e2 = hlock7 & v3747598 | !hlock7 & v3a557d2;
assign v3379070 = hgrant6_p & v8455e1 | !hgrant6_p & !v3a6b23f;
assign v3a57c48 = hbusreq2 & v3809a76 | !hbusreq2 & v8455ab;
assign v3776bc7 = hbusreq5_p & v3736e12 | !hbusreq5_p & v374723b;
assign v3766218 = hgrant2_p & v8455ab | !hgrant2_p & v3747d3c;
assign v3a6ff26 = hbusreq0 & v3724fe8 | !hbusreq0 & v3a711b9;
assign v3a672a8 = hmaster2_p & v374b5b6 | !hmaster2_p & v375bf93;
assign v377e4d8 = hmaster0_p & v3a6c6ad | !hmaster0_p & v3729793;
assign v3735ed2 = hmaster2_p & v37593a1 | !hmaster2_p & v3723501;
assign v3a6fdef = hlock0_p & v3a635ea | !hlock0_p & v373ead8;
assign v373502e = hgrant2_p & v8455e7 | !hgrant2_p & !v3a6d364;
assign v3726a86 = hlock4_p & v3747c3e | !hlock4_p & v8455ab;
assign aef136 = hgrant0_p & v3734967 | !hgrant0_p & v375b21c;
assign v377ed6c = hgrant4_p & v3761cd5 | !hgrant4_p & v3a68d70;
assign v372d7ed = hgrant2_p & v8455ab | !hgrant2_p & v3a5754b;
assign v3a5b40f = jx0_p & v3755f22 | !jx0_p & v3757519;
assign a6f8c7 = hbusreq3 & v3a63805 | !hbusreq3 & v3755791;
assign v374fe8e = hbusreq4_p & v3755dcd | !hbusreq4_p & !v3729421;
assign v3a70581 = hbusreq7 & v3a5d7f7 | !hbusreq7 & v3a6f3df;
assign v377249b = hmaster0_p & v374b824 | !hmaster0_p & !v377624b;
assign v3a61c45 = hbusreq4 & v3764141 | !hbusreq4 & v37696b6;
assign v37566f4 = hgrant0_p & v3756899 | !hgrant0_p & v8455ab;
assign v375b16e = hbusreq6 & v37379bb | !hbusreq6 & !v3a703de;
assign v3767483 = hgrant5_p & v2acaee4 | !hgrant5_p & v375cd7b;
assign v8455e9 = hgrant0_p & v8455ab | !hgrant0_p & !v8455ab;
assign v375df97 = hbusreq8_p & v3735bf3 | !hbusreq8_p & v3a6fb44;
assign v37796bf = hmaster1_p & v374ec35 | !hmaster1_p & v3728d9c;
assign v3807729 = hmaster0_p & v3a70853 | !hmaster0_p & v3761178;
assign v3a6eb97 = hgrant5_p & v377807f | !hgrant5_p & v3a58d5f;
assign v376e3d3 = hbusreq2_p & v3725ba8 | !hbusreq2_p & v3a6f0d1;
assign v3a6edab = hbusreq1_p & v37567c7 | !hbusreq1_p & v373b288;
assign v373428e = hbusreq4_p & v37596d5 | !hbusreq4_p & v372cbfc;
assign v376a91d = hmaster2_p & v37793a4 | !hmaster2_p & v37580b3;
assign v3773a06 = hgrant5_p & v3759cad | !hgrant5_p & v375a4f6;
assign v3a6dd80 = hmaster2_p & v3767e7e | !hmaster2_p & v3a70c39;
assign v3a63d5f = hbusreq7_p & v3a63f49 | !hbusreq7_p & v3a71546;
assign v3a5d2c5 = hmaster0_p & v376c898 | !hmaster0_p & c536d5;
assign v3a713a3 = hmaster0_p & v3a57d1f | !hmaster0_p & !v3771e23;
assign v376b662 = hbusreq5_p & v376afff | !hbusreq5_p & v8455ab;
assign v3a705a5 = hgrant2_p & v3a70e21 | !hgrant2_p & v3a6fde9;
assign v3a6f4fc = hbusreq1_p & v3770b89 | !hbusreq1_p & v3a6f32a;
assign v374e2a0 = hbusreq8_p & v3a66c49 | !hbusreq8_p & v3766bbb;
assign v3a5a2a4 = hbusreq8_p & v375f3cf | !hbusreq8_p & v375c999;
assign v3732b15 = hbusreq5_p & v3a5e2a9 | !hbusreq5_p & v8455ab;
assign v3769bf7 = hburst1_p & v8455ab | !hburst1_p & !v845605;
assign v37749bf = hgrant3_p & v8455be | !hgrant3_p & v37447bf;
assign v3a6ec17 = hlock6 & v3733103 | !hlock6 & v3809259;
assign b56d1b = hbusreq1 & v3a5600a | !hbusreq1 & v37757e0;
assign v3a7066e = hgrant0_p & v8455ab | !hgrant0_p & v37682c6;
assign v3a7017a = jx0_p & v3a70a22 | !jx0_p & v3a66cee;
assign v35772a5 = hmastlock_p & v845605 | !hmastlock_p & !v8455ab;
assign v2092eac = hbusreq3 & v37757e0 | !hbusreq3 & v8455ab;
assign v23fd96e = hbusreq0 & v376d3d1 | !hbusreq0 & v3a70d8a;
assign v3777009 = hbusreq2_p & v3750dd3 | !hbusreq2_p & !v8455ab;
assign v3a6895d = hmaster1_p & v377e4b4 | !hmaster1_p & v376e441;
assign v3a58cfc = hbusreq4_p & v3a619c0 | !hbusreq4_p & v3a66110;
assign v3a6669b = hmaster2_p & v3a70893 | !hmaster2_p & v377961f;
assign v376055d = hbusreq5_p & v374e4fd | !hbusreq5_p & v372f0c7;
assign v37710ad = hmaster1_p & v3737b63 | !hmaster1_p & v37377fd;
assign v3758a7c = hmaster0_p & v374e855 | !hmaster0_p & v882147;
assign v93ca8c = hmaster0_p & v3747a0d | !hmaster0_p & !v376bae4;
assign v3a55672 = hmaster0_p & v3732b63 | !hmaster0_p & v8455ab;
assign v377144d = hlock2_p & v3a600b8 | !hlock2_p & v3a6a0b0;
assign v3726d00 = hbusreq0_p & v3766e3a | !hbusreq0_p & v8455ab;
assign v37627f6 = hbusreq5 & v373576f | !hbusreq5 & v3755220;
assign v3755670 = hmaster2_p & v3a582c5 | !hmaster2_p & v35772a6;
assign a8fef2 = hmaster2_p & v380881d | !hmaster2_p & v375624e;
assign v37581cf = hbusreq5 & v372c3c7 | !hbusreq5 & v3a703d7;
assign v376723e = hlock8 & v374127d | !hlock8 & v3776e45;
assign v376d5a4 = hlock3_p & v3770559 | !hlock3_p & v35772a6;
assign v3a70fb1 = hmaster3_p & v3a707b4 | !hmaster3_p & v376959b;
assign v3734046 = hgrant0_p & v3733090 | !hgrant0_p & v3752e8e;
assign v375f020 = hlock6_p & v3723af9 | !hlock6_p & v8455bf;
assign v3731d66 = hlock7_p & v3a5b9c3 | !hlock7_p & !v8455ce;
assign v3728d2a = hbusreq2_p & v8455ab | !hbusreq2_p & d22727;
assign v3736b3b = hmaster1_p & v3a65287 | !hmaster1_p & !v376a3f5;
assign v3a5db5f = hmaster0_p & v372b1dc | !hmaster0_p & v3722fc0;
assign v3a59cce = hgrant5_p & v3731780 | !hgrant5_p & v3a553bc;
assign v3a70a96 = hmaster2_p & v3a6b6ef | !hmaster2_p & v8455ab;
assign v374e380 = hbusreq4_p & v3763668 | !hbusreq4_p & v377167e;
assign v37485bd = hbusreq0_p & v8455b0 | !hbusreq0_p & v3753dab;
assign v3747d3d = hmaster2_p & v3763175 | !hmaster2_p & v3753dab;
assign v3738a63 = hbusreq5_p & v3726e48 | !hbusreq5_p & v37523ea;
assign v3723de9 = hbusreq7_p & v3a71442 | !hbusreq7_p & v8455b7;
assign v3a7051d = hbusreq5_p & v38088b6 | !hbusreq5_p & v3a58c07;
assign v3777790 = hbusreq6_p & v3a6d2ae | !hbusreq6_p & !v8455ab;
assign v3a6ffd7 = hmaster1_p & v375c92f | !hmaster1_p & !v37350b2;
assign v376ec9b = hlock5 & v3a703cb | !hlock5 & v3a700a3;
assign v3742dcb = hmaster1_p & v376bd2c | !hmaster1_p & v372348f;
assign v3727615 = hgrant2_p & ae0781 | !hgrant2_p & v3a6d3f3;
assign v3a6f83f = jx0_p & v8455ab | !jx0_p & v3735f31;
assign v37430f0 = hbusreq5_p & v3a633c5 | !hbusreq5_p & v3a5fc48;
assign db9e30 = hgrant6_p & v8455ab | !hgrant6_p & v3a709af;
assign v372acd3 = hmaster1_p & v8455ab | !hmaster1_p & v3a61d1f;
assign v3808884 = hbusreq8 & v373f4cf | !hbusreq8 & v38076b7;
assign v374975c = hbusreq5_p & v3730402 | !hbusreq5_p & v373ba2e;
assign v3a710c3 = hmaster2_p & v37578d4 | !hmaster2_p & v3775750;
assign v3a5e24e = busreq_p & v1e38275 | !busreq_p & !v39ebac7;
assign v3a577f2 = hlock2_p & v376ce37 | !hlock2_p & v3a71689;
assign v3a6e94b = hbusreq2 & v360cdfe | !hbusreq2 & v8455bf;
assign v377077a = hmaster0_p & v8455ab | !hmaster0_p & v375e133;
assign v3a70d64 = hbusreq3_p & v373f0ee | !hbusreq3_p & v3a69946;
assign v373a2f4 = hmaster0_p & v3725392 | !hmaster0_p & v3a61c70;
assign v3a6167d = hlock7_p & v37758e6 | !hlock7_p & v3a5e3d1;
assign v3760617 = hgrant5_p & v99b721 | !hgrant5_p & v3762617;
assign v373bb50 = hbusreq0 & v372de43 | !hbusreq0 & v377b68e;
assign v376beb3 = hgrant5_p & v374b873 | !hgrant5_p & v3a702ef;
assign v37312f4 = hbusreq7_p & v3755967 | !hbusreq7_p & v3a6199f;
assign v3738c5f = hmaster2_p & v3a70b92 | !hmaster2_p & v3748d67;
assign v37282f7 = hmaster2_p & v375f619 | !hmaster2_p & v3a621e7;
assign v2ff9348 = hbusreq6_p & v38072fd | !hbusreq6_p & v3a5df87;
assign v3a63c47 = hmaster2_p & v8455ab | !hmaster2_p & v3736739;
assign v372fe28 = hlock7_p & v374f3a9 | !hlock7_p & v3a643d6;
assign v3a65f7a = hbusreq6_p & v37244a0 | !hbusreq6_p & v3778323;
assign v377f61e = hgrant4_p & v377d78b | !hgrant4_p & v373e5a7;
assign v372ff72 = hbusreq2_p & v3a71417 | !hbusreq2_p & v3731300;
assign v377adf0 = hbusreq6_p & v375c505 | !hbusreq6_p & v8455b0;
assign v3773d39 = hbusreq6 & v3a7084e | !hbusreq6 & v8455bb;
assign v3a6fc27 = hbusreq4 & v3a70248 | !hbusreq4 & v8455ab;
assign v374a2be = hbusreq6_p & v3a66ef6 | !hbusreq6_p & v3a5b583;
assign v374153d = hlock5_p & v3a6fb8d | !hlock5_p & v3a645ac;
assign v377a01a = hmaster1_p & v3a70209 | !hmaster1_p & v3a712ed;
assign v3a6f8bb = hgrant3_p & v3774416 | !hgrant3_p & v373c331;
assign v374c05b = hbusreq7_p & v3758559 | !hbusreq7_p & v3744e62;
assign v3778637 = hgrant6_p & v3a67ffe | !hgrant6_p & v3a5ee7d;
assign v360d0fd = hgrant4_p & v3a5d2d3 | !hgrant4_p & v325b59f;
assign v2acaf4f = hlock5_p & v376a14f | !hlock5_p & v3a7151b;
assign v3742950 = hmaster0_p & v375a28e | !hmaster0_p & v3767e71;
assign v375f172 = hmaster0_p & v377c9cb | !hmaster0_p & v3808e2e;
assign v37509af = hbusreq0_p & v3a66140 | !hbusreq0_p & v37717f4;
assign v3a6f6b4 = hbusreq6_p & v3752c04 | !hbusreq6_p & v376e794;
assign v37c011c = hlock1_p & v37749b7 | !hlock1_p & !v8455ab;
assign v3737e57 = hmaster1_p & v3a7161a | !hmaster1_p & v3a6c573;
assign v3a708a6 = hlock7 & v3a5b448 | !hlock7 & v377b4b0;
assign v377cd41 = hbusreq7 & v377a422 | !hbusreq7 & v376fc7f;
assign v374c69c = hmaster0_p & v372580e | !hmaster0_p & v3a70b98;
assign v3a65096 = hmaster1_p & v376c652 | !hmaster1_p & v37266df;
assign v3765962 = jx0_p & v37470a5 | !jx0_p & v8455ab;
assign v373226c = hgrant1_p & v3742d60 | !hgrant1_p & v8455ab;
assign v373dd40 = hbusreq7 & v3a63688 | !hbusreq7 & v374d617;
assign v3748d3b = hbusreq3_p & v3a6fcf9 | !hbusreq3_p & v374f609;
assign v90829e = hbusreq2_p & v23fde92 | !hbusreq2_p & v3a704f8;
assign v3a70468 = hlock4_p & v3a713df | !hlock4_p & v8455b0;
assign v372715f = hlock5_p & v3733168 | !hlock5_p & !v8455ab;
assign v3a6faae = hmaster0_p & v3a59f7d | !hmaster0_p & v37527dc;
assign v373adae = hgrant0_p & v373bd24 | !hgrant0_p & v3777e08;
assign v3a62ef1 = jx1_p & v3768adf | !jx1_p & v3755898;
assign v372e6d0 = hbusreq8 & v374f26c | !hbusreq8 & v3a70a90;
assign v37654f4 = hbusreq0 & v377c842 | !hbusreq0 & v3735a71;
assign v3a701bc = hbusreq5_p & v377b0a3 | !hbusreq5_p & v3760927;
assign v3a5cc27 = hmaster0_p & v8455c1 | !hmaster0_p & v376a6f1;
assign v3776864 = hmaster0_p & v377cc52 | !hmaster0_p & v374677a;
assign v3a69bfd = hbusreq4_p & v2aca264 | !hbusreq4_p & v373422b;
assign v37457d1 = hlock0_p & v8455e7 | !hlock0_p & v373a07f;
assign v372d98c = hmaster2_p & v3a635ea | !hmaster2_p & v3a663b9;
assign v377002f = hgrant3_p & v3a70a7f | !hgrant3_p & v37756ac;
assign v3a5aacb = hgrant6_p & v375da10 | !hgrant6_p & v3a6f61f;
assign v3737209 = hlock2 & b516f2 | !hlock2 & v377a43e;
assign v375a8a7 = hmaster1_p & v3a5fa4c | !hmaster1_p & v8455ab;
assign v3a5cf57 = hbusreq8 & v373a0f8 | !hbusreq8 & v3756200;
assign v375c4ef = hmaster1_p & v373e376 | !hmaster1_p & v3a566c0;
assign v3a55773 = hbusreq0 & v3a703cd | !hbusreq0 & v372c3b9;
assign v3769a36 = hgrant2_p & v377d4a0 | !hgrant2_p & v3778345;
assign v37285c9 = hmaster2_p & v374a637 | !hmaster2_p & v8455ab;
assign v372dc39 = hbusreq5 & v3a6f455 | !hbusreq5 & v3a70135;
assign v3a6fac4 = hlock3 & v377b515 | !hlock3 & v39a5350;
assign v375fbba = hmaster2_p & v3736ded | !hmaster2_p & v3732415;
assign v374fd0b = hbusreq8 & v377a0cb | !hbusreq8 & v372e02c;
assign v375b8b9 = hgrant6_p & v3727d95 | !hgrant6_p & v3775aef;
assign v372640f = hlock4_p & v374caab | !hlock4_p & v8455e7;
assign v375f0af = hbusreq2_p & v3a6ffe5 | !hbusreq2_p & v373125c;
assign v373e0b5 = hlock7 & v373d25a | !hlock7 & v3a53392;
assign v37265c1 = hbusreq5 & v375671a | !hbusreq5 & v376cd02;
assign v373c642 = hmaster0_p & v3734967 | !hmaster0_p & v3751861;
assign v3a6ff98 = hmaster2_p & v375b429 | !hmaster2_p & v8455b0;
assign v3577388 = hbusreq7 & v8e4471 | !hbusreq7 & v373dafe;
assign v377015c = hbusreq4_p & v32562a3 | !hbusreq4_p & v3748146;
assign v3751db5 = hlock4 & b04260 | !hlock4 & v373c7a5;
assign v374514e = hmaster0_p & v28896b4 | !hmaster0_p & v377d4de;
assign v3a6ec0b = hmaster0_p & v373195f | !hmaster0_p & v3a5f000;
assign v3733bed = jx1_p & v377b61e | !jx1_p & v3a6b372;
assign v3724f6b = hgrant5_p & v3745428 | !hgrant5_p & v377586d;
assign v3a60aca = hgrant6_p & v3726bff | !hgrant6_p & v3a5b41c;
assign v3a5759a = hgrant3_p & v3a56aeb | !hgrant3_p & v1e3825d;
assign v372542e = hmaster2_p & v3a5e24e | !hmaster2_p & !v3733e9e;
assign dc57c8 = jx1_p & v8455ab | !jx1_p & v3a695ec;
assign v3a61f33 = jx0_p & v373e225 | !jx0_p & v377f6a5;
assign v3a6f562 = hlock0_p & v37376c8 | !hlock0_p & v3736d51;
assign v372abac = hgrant4_p & v8455ab | !hgrant4_p & v3745241;
assign v3a6d622 = hgrant4_p & v374d92c | !hgrant4_p & v37507f4;
assign v373ba25 = hmaster1_p & v3a61280 | !hmaster1_p & v373d32e;
assign v3a624da = hbusreq6_p & v3722e5c | !hbusreq6_p & v35772a6;
assign v3a67dd8 = hmaster1_p & v3a547ff | !hmaster1_p & v3a640fd;
assign v3a5ba8a = hmaster1_p & v3735f67 | !hmaster1_p & v3a70143;
assign v3a58589 = hmaster1_p & v37263bf | !hmaster1_p & v3a6776f;
assign v3730fc0 = hlock6 & v3a6e6e1 | !hlock6 & v37626a4;
assign v3748489 = hmaster2_p & v3a6fdef | !hmaster2_p & v374acbe;
assign v3758d2a = hmaster2_p & v3754dd0 | !hmaster2_p & v3a7153c;
assign v37414cd = hbusreq8_p & v3a70195 | !hbusreq8_p & v3739768;
assign v3774061 = hgrant0_p & v376e914 | !hgrant0_p & !v3a2a2fa;
assign v377f640 = hbusreq5_p & v3a65402 | !hbusreq5_p & !v376af1a;
assign v376fa76 = hgrant3_p & v8455ab | !hgrant3_p & v37664ab;
assign v375a251 = hbusreq7_p & v3a5dd8a | !hbusreq7_p & v3a5aa93;
assign v3727215 = hbusreq3 & v37674c1 | !hbusreq3 & !v8455ab;
assign v374874a = hbusreq6_p & v3741d99 | !hbusreq6_p & v3736f3b;
assign v3723abc = hbusreq6 & v374362e | !hbusreq6 & !v3a5e922;
assign v375efa4 = hgrant4_p & v375648e | !hgrant4_p & v3754aa3;
assign v3722b21 = hlock5 & v3a7008f | !hlock5 & v3727363;
assign v37433ef = hbusreq0 & v37232a6 | !hbusreq0 & v3a7156a;
assign v374c3f2 = hbusreq4_p & v39a537f | !hbusreq4_p & !v39a5381;
assign v37682ce = hmaster0_p & v3a6ebf7 | !hmaster0_p & !v8455ab;
assign v377f200 = hlock0_p & v376f56d | !hlock0_p & v3728826;
assign v3a6f17f = hbusreq4_p & v37446b5 | !hbusreq4_p & !v3a7107a;
assign v373dd5a = hmaster0_p & v3779680 | !hmaster0_p & v37297e8;
assign v374ce2a = hlock7_p & v3a67fc6 | !hlock7_p & v37743c6;
assign v376c1d6 = hmaster0_p & v375095a | !hmaster0_p & v3753a65;
assign v37591f2 = hbusreq7 & v375a543 | !hbusreq7 & v3a6f068;
assign v3a613da = hbusreq5_p & v375b6c3 | !hbusreq5_p & !v376eed1;
assign v3a6556a = hbusreq4 & v8455b0 | !hbusreq4 & v3722e7a;
assign v376ec4f = hlock8 & v3a70ab3 | !hlock8 & v3a6fb4f;
assign v375400b = hbusreq3 & v3737d44 | !hbusreq3 & v8455ab;
assign v3733b0c = hbusreq6_p & v3725ba8 | !hbusreq6_p & v376e3d3;
assign v3a70b94 = hburst0 & v3757c6f | !hburst0 & v3773092;
assign v374b697 = hlock0_p & v3a67983 | !hlock0_p & v8455b0;
assign v3769e8c = hgrant2_p & v8df61b | !hgrant2_p & v3a63ff3;
assign v360d00f = hlock5 & v3777517 | !hlock5 & v3a6bf3c;
assign v3779717 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3747314;
assign v3a6fde8 = hlock1_p & v8455ab | !hlock1_p & !v3a6ac26;
assign v3a70dc3 = hmaster3_p & v375be25 | !hmaster3_p & v3755db9;
assign v3a6fd31 = hmaster0_p & v3730a8b | !hmaster0_p & !v372362a;
assign v374705f = hmaster1_p & v3a6b8e8 | !hmaster1_p & v3a70cc7;
assign v3a61734 = hbusreq4_p & v3747302 | !hbusreq4_p & v377b946;
assign v92e5bb = hmaster2_p & v375139d | !hmaster2_p & v374a2cc;
assign v3a70edb = hlock3_p & v3a71263 | !hlock3_p & v3761181;
assign v3736610 = hgrant4_p & v39ea76e | !hgrant4_p & v3378d8f;
assign v3a615f7 = hbusreq3_p & v3773e2a | !hbusreq3_p & v3a6f986;
assign v3748858 = hbusreq0 & v3a707ae | !hbusreq0 & v37591ae;
assign v3a5f60c = hmaster0_p & v8455e7 | !hmaster0_p & v3a5ff26;
assign v37263bc = hlock0_p & v3760e7b | !hlock0_p & v3a63260;
assign v3737a29 = hbusreq6 & v37678fc | !hbusreq6 & v8455b3;
assign v373f408 = hbusreq8_p & v3737808 | !hbusreq8_p & v377577b;
assign v375b9b2 = hbusreq4 & v3a660f2 | !hbusreq4 & v8455ab;
assign v3a706f8 = hmaster2_p & v3779060 | !hmaster2_p & !v372391f;
assign v3a6eee8 = hmaster0_p & v3723c3f | !hmaster0_p & v37643e6;
assign v3a6fae9 = hgrant4_p & v8455ab | !hgrant4_p & v3754565;
assign v37465d7 = hbusreq8_p & v373dee7 | !hbusreq8_p & v3764c4a;
assign v374490b = hmaster0_p & v3a5d365 | !hmaster0_p & v373a822;
assign v375e813 = hbusreq5_p & v3725c13 | !hbusreq5_p & !v8455ab;
assign v3759a21 = hbusreq6 & v3a6f32f | !hbusreq6 & !v3a7101b;
assign v3741022 = hlock4_p & v377ba55 | !hlock4_p & !v8455ab;
assign v3770af1 = hbusreq1_p & v3730da3 | !hbusreq1_p & v3a63621;
assign v3777ee9 = hbusreq6 & v3a6fbd8 | !hbusreq6 & v373261f;
assign b412f3 = hlock7_p & v372b627 | !hlock7_p & !v8455ab;
assign v372bfbb = hbusreq6_p & v374faa9 | !hbusreq6_p & v37621ff;
assign v3769712 = hmaster1_p & v3a6e31f | !hmaster1_p & v3753927;
assign v37261df = hbusreq0_p & v1e37e66 | !hbusreq0_p & v8455ab;
assign cea42b = hbusreq7_p & v3731fe4 | !hbusreq7_p & v3777d70;
assign v3a57801 = hlock5 & v3727960 | !hlock5 & v292554f;
assign v3a6af0b = hlock0 & v373eaee | !hlock0 & v372dde7;
assign v377a9b8 = hmaster1_p & v37469c4 | !hmaster1_p & v3752183;
assign v39e9c97 = hbusreq2_p & v3a2981b | !hbusreq2_p & v372949c;
assign v3a55c0c = hgrant4_p & v3a6ef98 | !hgrant4_p & v1e37ebb;
assign v3760f4e = hbusreq3_p & v8455b3 | !hbusreq3_p & v3767437;
assign v3a641ea = hmaster2_p & v372b1dc | !hmaster2_p & !d1bf3b;
assign v376a9de = hgrant6_p & v3766924 | !hgrant6_p & v3730217;
assign v3a70cc5 = hbusreq1_p & v3a6f5c0 | !hbusreq1_p & v8455ab;
assign v3772db0 = stateG10_1_p & v8455ab | !stateG10_1_p & v3746f37;
assign v3739ab6 = hbusreq0 & v3751734 | !hbusreq0 & v8455ab;
assign v372d1b1 = jx0_p & v37430db | !jx0_p & v8455ab;
assign v3740174 = hbusreq4_p & v3a55dc3 | !hbusreq4_p & v3758c32;
assign v3378594 = hbusreq6 & v37440a8 | !hbusreq6 & v37372c9;
assign v3746312 = hbusreq8 & v3749544 | !hbusreq8 & v3776859;
assign v374d92c = hbusreq4_p & v3a6d5e9 | !hbusreq4_p & v37766f3;
assign v8455f5 = hgrant6_p & v8455ab | !hgrant6_p & !v8455ab;
assign v3a66856 = hmaster0_p & v373308b | !hmaster0_p & v3770cb8;
assign v3723495 = hgrant2_p & v3778fec | !hgrant2_p & v375abcd;
assign v3a6984f = hbusreq6_p & v3a635ea | !hbusreq6_p & v3a70b9a;
assign v374ac24 = hmaster2_p & v3733aa5 | !hmaster2_p & v3767f7f;
assign v375d337 = hgrant4_p & v375a268 | !hgrant4_p & v3a70f48;
assign v3724392 = hbusreq2_p & v3a6ffe5 | !hbusreq2_p & v3757fcc;
assign v372cfdf = hbusreq6 & b41a29 | !hbusreq6 & v3755c8b;
assign v3757735 = hmaster2_p & v3a6f7dd | !hmaster2_p & v3a5a6e6;
assign v3a2a41f = hbusreq5_p & v373a693 | !hbusreq5_p & v3769215;
assign v3a5b469 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a62caa;
assign v3a55466 = hbusreq5_p & v3734fba | !hbusreq5_p & v3a63f9a;
assign v3a6f6df = hgrant1_p & v3a653e4 | !hgrant1_p & !v8455ab;
assign v376e9e1 = hbusreq7 & v8f9a63 | !hbusreq7 & v8455ab;
assign v376daec = hbusreq4 & v3731991 | !hbusreq4 & v3a62a6d;
assign v3a62753 = hbusreq5 & v3a6f59e | !hbusreq5 & v376fbb5;
assign v8686c3 = jx1_p & v375e9c0 | !jx1_p & v3757fdd;
assign v3a5ba28 = hbusreq4_p & v37541a7 | !hbusreq4_p & v8455bb;
assign v377f6ae = hmaster2_p & v377d045 | !hmaster2_p & v3755a83;
assign v3a5aa64 = hbusreq8_p & v3a70cb4 | !hbusreq8_p & v3757e71;
assign v3723d73 = hbusreq5 & v3a704be | !hbusreq5 & v8455c7;
assign v375a500 = hmaster2_p & v375e721 | !hmaster2_p & v374e1c3;
assign v377a422 = hmaster1_p & v372bd46 | !hmaster1_p & v3757a04;
assign v375c482 = hlock2_p & v37336f0 | !hlock2_p & v376773b;
assign v37458d2 = hbusreq4 & v3a6dbf0 | !hbusreq4 & v3a6fba6;
assign v3a6fd9b = hbusreq5_p & v3765c49 | !hbusreq5_p & v373e891;
assign v3a7075b = hmaster0_p & v3a6f255 | !hmaster0_p & v3a70304;
assign v3765013 = hbusreq2 & v3a6b77d | !hbusreq2 & v8455ab;
assign v372cc0a = hgrant6_p & v35b774b | !hgrant6_p & v37542af;
assign v3726f6c = hbusreq3 & v37457fb | !hbusreq3 & v8455e7;
assign v375c7b9 = locked_p & v8455ab | !locked_p & !v8455e1;
assign v376d091 = hlock5_p & v3a555ae | !hlock5_p & v3a69ead;
assign v3759532 = hbusreq7 & v3a63f7b | !hbusreq7 & v3745d1e;
assign v375fcbf = hmaster2_p & v3a6f018 | !hmaster2_p & v375efa4;
assign v374ba61 = hlock4 & v3772567 | !hlock4 & v3754b98;
assign v3a54677 = hbusreq5 & v374ac2e | !hbusreq5 & v3771c85;
assign v35b7092 = hbusreq0 & v37266c2 | !hbusreq0 & v373a9ee;
assign v376da28 = hbusreq0_p & v374f1a1 | !hbusreq0_p & v8455ab;
assign v3a7010c = hmaster0_p & v374b25d | !hmaster0_p & !v8455bf;
assign v3a57721 = hmaster0_p & v376c248 | !hmaster0_p & v3a70ba9;
assign v37421bd = hbusreq5_p & v37385ee | !hbusreq5_p & !v3a678de;
assign v376a6d7 = hgrant0_p & v8455ab | !hgrant0_p & !v375c5a1;
assign v375693b = hgrant4_p & v3759b71 | !hgrant4_p & v3758ea7;
assign v373f14d = hmaster0_p & v3a6279b | !hmaster0_p & v3741e56;
assign v3767d1b = hgrant6_p & v3a6406d | !hgrant6_p & v3a594a5;
assign v3a59f7d = hmaster2_p & v373cc68 | !hmaster2_p & v8455ab;
assign v37329e1 = hbusreq6 & v376f542 | !hbusreq6 & !v8455ab;
assign v372e33d = hmaster2_p & v373e474 | !hmaster2_p & v37745c3;
assign v3a63bb0 = hbusreq1 & v3a64ee3 | !hbusreq1 & !v3a70131;
assign v375e431 = hmaster0_p & v8455ab | !hmaster0_p & !v3a6a5e6;
assign v3754777 = hbusreq6 & v3723e1f | !hbusreq6 & v3a635ea;
assign v376d143 = hgrant4_p & v8455ab | !hgrant4_p & v3a54560;
assign v37503bd = hmaster0_p & v374306c | !hmaster0_p & v3724398;
assign v3a71611 = hmaster2_p & v35ba1a5 | !hmaster2_p & v376a96b;
assign v3a71016 = hbusreq6_p & v372b59d | !hbusreq6_p & v8455ab;
assign v37474c1 = hmaster3_p & v373fe61 | !hmaster3_p & v3a6d0ae;
assign v375b389 = hbusreq5_p & v3a707f0 | !hbusreq5_p & v3a6fe50;
assign v372cd37 = hlock5_p & v3a5fd58 | !hlock5_p & !v3763c97;
assign v3a5fdfc = hgrant4_p & v37375ee | !hgrant4_p & v375444e;
assign v374ec84 = hgrant0_p & v372df47 | !hgrant0_p & v8455ab;
assign v375609e = hlock5_p & v372ef56 | !hlock5_p & v3a70ba1;
assign v1e3791d = hlock0_p & v373a841 | !hlock0_p & v3765e46;
assign v3a68dcb = hbusreq5 & v3736012 | !hbusreq5 & v8455ab;
assign v3a713d7 = hmaster3_p & v3a71312 | !hmaster3_p & v377740c;
assign v377772d = hmaster0_p & v376984d | !hmaster0_p & v337902c;
assign v3756d53 = hmaster0_p & v8455ca | !hmaster0_p & v3776b09;
assign v376596e = hmaster1_p & v376a31b | !hmaster1_p & v3753389;
assign v37525b0 = hmaster2_p & v377fb43 | !hmaster2_p & !v8455ab;
assign v3a6f04f = jx1_p & v3763a1e | !jx1_p & v3a70d5c;
assign v373afd0 = hmaster2_p & v3a5e24e | !hmaster2_p & !v3a70ee7;
assign v3a70515 = hlock5_p & v3773089 | !hlock5_p & v374949f;
assign v372bce5 = hbusreq7_p & v3a715d0 | !hbusreq7_p & v375d2ff;
assign v3728213 = hlock0 & v375da10 | !hlock0 & v3759f66;
assign v375a38e = hlock4 & v3745c75 | !hlock4 & v3743c51;
assign v37328f1 = hmaster2_p & v3741fc9 | !hmaster2_p & v372f553;
assign v3745803 = hmaster2_p & v37646e1 | !hmaster2_p & v3809a6a;
assign v3a6f2cf = hgrant6_p & v3a70240 | !hgrant6_p & v3a64417;
assign v372f216 = hbusreq4_p & v3a70ca3 | !hbusreq4_p & !v3a65526;
assign v37438ab = hlock4 & v374217a | !hlock4 & v3a6dfc9;
assign v3a5a17f = hmaster2_p & v3a68426 | !hmaster2_p & v372ab21;
assign v3a63f55 = hmaster1_p & v37261b3 | !hmaster1_p & c7ba89;
assign v375c691 = hlock8_p & v8455ab | !hlock8_p & b412f3;
assign v372ac1d = hbusreq5_p & v3a70943 | !hbusreq5_p & v3a6fb88;
assign v37485cb = hbusreq5 & v376eb68 | !hbusreq5 & v3760765;
assign v375ab6d = hbusreq2 & v372b5f5 | !hbusreq2 & v8455ab;
assign v3a6efd9 = hmaster0_p & v3a63ea7 | !hmaster0_p & v3759031;
assign v3771697 = hbusreq4_p & v3a7120c | !hbusreq4_p & v373fc07;
assign v3746d89 = hmaster2_p & v375de18 | !hmaster2_p & v37521ed;
assign v3a715b8 = hbusreq7 & v377e071 | !hbusreq7 & v3a6ec01;
assign v3a639e7 = hmaster0_p & v3a701c6 | !hmaster0_p & !v374677a;
assign v373f834 = hmaster0_p & v3772229 | !hmaster0_p & v390071e;
assign v360cd91 = jx1_p & v3a70f7c | !jx1_p & v3744dda;
assign v3a71580 = hmaster0_p & v373a3b9 | !hmaster0_p & v373c545;
assign v3808914 = hmaster1_p & v3a668e4 | !hmaster1_p & v3a714ab;
assign v37462e7 = hgrant4_p & v372f3e0 | !hgrant4_p & v376f1c0;
assign v374db48 = hbusreq5_p & v3a62d1c | !hbusreq5_p & !v952f44;
assign v3768172 = hbusreq5 & v374fde8 | !hbusreq5 & !v377a886;
assign v377167c = hmaster2_p & v33789b9 | !hmaster2_p & v3753258;
assign v372e096 = hbusreq4 & v37738fc | !hbusreq4 & v35b774b;
assign v373632b = hgrant0_p & v376ea4a | !hgrant0_p & !v3a70913;
assign v3a603b6 = hbusreq5 & v37524b2 | !hbusreq5 & v8bc0e2;
assign v3778857 = hbusreq5 & v376fbe3 | !hbusreq5 & v3755691;
assign v374464b = hgrant5_p & v3729808 | !hgrant5_p & v3a70df6;
assign v376a34d = hgrant3_p & v375d689 | !hgrant3_p & v3732b81;
assign v375859a = hmaster0_p & v3725b9b | !hmaster0_p & v3733767;
assign v372b6db = hbusreq6_p & v3767018 | !hbusreq6_p & !v8455ab;
assign v3a7156e = hbusreq5 & v3751d41 | !hbusreq5 & v37438fc;
assign v3753f0d = hlock4 & v3735ad2 | !hlock4 & v376f2a7;
assign v372a93f = hmaster0_p & v3744039 | !hmaster0_p & v375d507;
assign v3a6f4b9 = hmaster1_p & v373cb89 | !hmaster1_p & v374975c;
assign v1e37cec = hburst0 & v3a6ac2a | !hburst0 & v3750371;
assign v38076cf = hlock5_p & v8455ab | !hlock5_p & !v8455d9;
assign v3a6ffe5 = hlock2_p & v3a6bc47 | !hlock2_p & v35b70e6;
assign v3738a2b = hmaster2_p & v37718fb | !hmaster2_p & v374ebb0;
assign v3779b12 = hlock8 & v3a648a6 | !hlock8 & v3a6f194;
assign v37540d9 = hmaster2_p & v377b429 | !hmaster2_p & v8455ab;
assign v3a6f0d5 = hmaster0_p & v377f734 | !hmaster0_p & v376d0ff;
assign v23fdebb = hmaster2_p & v3768495 | !hmaster2_p & v376300a;
assign v3749629 = hbusreq3_p & v37427d3 | !hbusreq3_p & v3759947;
assign v3a5f587 = hmaster0_p & v377f85a | !hmaster0_p & v3a59caa;
assign v3a70bb7 = hgrant6_p & v372f87b | !hgrant6_p & v3a6837d;
assign v3a6c322 = hmaster1_p & v376c4ef | !hmaster1_p & v3728d9c;
assign v377ce5e = hmaster2_p & v3a6f501 | !hmaster2_p & v3a685c7;
assign v3760fb0 = hbusreq0 & v3a65384 | !hbusreq0 & v8455ab;
assign v3775e2e = hgrant4_p & v3747ed4 | !hgrant4_p & v374d153;
assign v3a70ebb = hbusreq7_p & v3752edb | !hbusreq7_p & v376ed36;
assign v373180e = start_p & v845605 | !start_p & v372c42d;
assign v3761d4c = hmaster2_p & v3763fdc | !hmaster2_p & v377988b;
assign v3a708c3 = hgrant4_p & v3a5690d | !hgrant4_p & v373109c;
assign v3725c68 = hlock3 & v377ac8a | !hlock3 & v3a6f757;
assign b3d3ad = hbusreq3_p & v373502a | !hbusreq3_p & v3a69946;
assign v377b0a3 = hmaster0_p & v3745181 | !hmaster0_p & v3a6fe5e;
assign v3767d4b = hbusreq0 & v3a71429 | !hbusreq0 & v3733be1;
assign v3a6df9a = hlock4_p & v377de7b | !hlock4_p & v373f058;
assign v37626ab = hmaster2_p & v2092faa | !hmaster2_p & v3a6f312;
assign v3a712b5 = hgrant5_p & v8455ab | !hgrant5_p & v3a67eb2;
assign v3a5e0f7 = hgrant2_p & v8455ba | !hgrant2_p & v3a55e7f;
assign v374c7e6 = hbusreq5_p & v376de5c | !hbusreq5_p & v3738ea9;
assign afa913 = hmaster2_p & v375af43 | !hmaster2_p & v375981e;
assign v3776dcd = hgrant4_p & v3a6f1ad | !hgrant4_p & v3a6ac26;
assign v3765bf4 = hmaster0_p & v3a6f9bd | !hmaster0_p & v3762dcf;
assign v3a683e2 = hlock6_p & v373c978 | !hlock6_p & v8455ab;
assign v3a6049f = hbusreq5 & v35b779e | !hbusreq5 & v3a2a107;
assign v376978e = hbusreq7_p & v35ba2cb | !hbusreq7_p & v3a715eb;
assign v3a598da = hbusreq5_p & v39ebb31 | !hbusreq5_p & v39ea0c2;
assign v377f486 = hbusreq4 & v3a705ad | !hbusreq4 & v964c47;
assign v3a5f946 = hbusreq5 & v3735e69 | !hbusreq5 & v374ffc1;
assign v375047c = hlock5 & v373d78f | !hlock5 & v3a61724;
assign v3766cd5 = hbusreq6_p & v3745069 | !hbusreq6_p & v3754940;
assign v3755a9f = hburst0 & v3a6ff41 | !hburst0 & v8455e1;
assign v374baac = hgrant6_p & v8455ab | !hgrant6_p & v377efd0;
assign v375de73 = hbusreq7 & v3a665ca | !hbusreq7 & v3a6b32d;
assign v377c31a = hgrant0_p & v3724057 | !hgrant0_p & v8455ab;
assign v3a55ecf = hlock6_p & v372f192 | !hlock6_p & v3a6f5d1;
assign v372c41f = hmaster2_p & v3a6e6fa | !hmaster2_p & v3750adf;
assign v37264c9 = hbusreq4 & v375a166 | !hbusreq4 & v37285eb;
assign v375ecd4 = hbusreq5 & v377d04f | !hbusreq5 & v3a6857b;
assign v376402f = stateA1_p & v3a70a83 | !stateA1_p & v8455ab;
assign v3745993 = hbusreq2 & v3a6d74f | !hbusreq2 & v8455ab;
assign v3776ca8 = hbusreq2_p & v372bf93 | !hbusreq2_p & v8455ab;
assign v3775f1f = hgrant4_p & v372d3ea | !hgrant4_p & v373f488;
assign v3a5af94 = hbusreq6_p & v3a619c0 | !hbusreq6_p & v3a66110;
assign v3779b9c = hmaster0_p & v3723c99 | !hmaster0_p & v3a5ef76;
assign v3724ab6 = hmaster2_p & v374a08a | !hmaster2_p & v37427e9;
assign v3a556ab = hmaster0_p & v3a6f90f | !hmaster0_p & v8455ab;
assign v3a6212a = hbusreq0_p & v3748797 | !hbusreq0_p & v372e169;
assign v209306f = hmaster1_p & v37793e4 | !hmaster1_p & v3763db6;
assign v37349cc = hmaster2_p & v376b88d | !hmaster2_p & v3768685;
assign v37637d5 = hbusreq6 & v377caa3 | !hbusreq6 & v8455bf;
assign v372495f = hbusreq6 & v3754b61 | !hbusreq6 & v372c500;
assign v375fb03 = hmaster2_p & v3a6fafd | !hmaster2_p & v3a71164;
assign v3a710e1 = hbusreq2_p & v372be4a | !hbusreq2_p & v8455b0;
assign v377d78b = hbusreq4_p & v3740672 | !hbusreq4_p & v32559c3;
assign v37620b4 = hlock5 & v3a70398 | !hlock5 & v3a6ef6f;
assign v37557a0 = hmaster0_p & v3756a6f | !hmaster0_p & v373af66;
assign v3773708 = hmaster2_p & v8455b0 | !hmaster2_p & v3752dd0;
assign v3753f35 = hmaster1_p & v8455ab | !hmaster1_p & v3a6eec5;
assign v3a70919 = hgrant5_p & v8455c6 | !hgrant5_p & v3731b53;
assign v3a5f4e0 = hmaster0_p & v3808d47 | !hmaster0_p & v3a59905;
assign v3a7046f = hbusreq7_p & v23fe1ca | !hbusreq7_p & !v373d0a2;
assign v3a6f772 = hmaster0_p & v376501e | !hmaster0_p & v372dcaa;
assign v3763bc4 = hbusreq5_p & v37680de | !hbusreq5_p & v3a6eb36;
assign v374e06d = hmaster3_p & v376c88f | !hmaster3_p & v3777d70;
assign v372c79f = hbusreq7_p & v376822d | !hbusreq7_p & !v8455ab;
assign v37273c2 = hgrant3_p & v3a6251b | !hgrant3_p & v3759b9a;
assign v3a71232 = hbusreq4_p & v8455ab | !hbusreq4_p & !v3a637dd;
assign v3a6f7fd = hbusreq2_p & v372ce8b | !hbusreq2_p & !v3a68591;
assign v376e093 = hbusreq2 & v3a6ff3f | !hbusreq2 & v8455ab;
assign v3739904 = hmaster0_p & v37526a5 | !hmaster0_p & v377ea20;
assign v3751887 = hbusreq5 & v3a6bf05 | !hbusreq5 & v3759aec;
assign v3722ad4 = hbusreq5 & v3a60dfb | !hbusreq5 & v3a5f5f5;
assign v377a9e7 = hbusreq2_p & v3a71528 | !hbusreq2_p & v3a70272;
assign v37c0170 = hbusreq8 & v37762ec | !hbusreq8 & v3737808;
assign v37267d6 = hbusreq0 & v3735e89 | !hbusreq0 & v37787da;
assign v377929d = hmaster1_p & v3a661fe | !hmaster1_p & v373bbc1;
assign v375f619 = hgrant4_p & v3a70a88 | !hgrant4_p & v38073c9;
assign v37403b1 = hlock5 & v3751383 | !hlock5 & v3755e61;
assign v37576b1 = hmaster0_p & v3a6e5f0 | !hmaster0_p & v95a0a1;
assign v3779924 = hbusreq4 & v3a697f1 | !hbusreq4 & !v372d924;
assign c511c2 = hgrant0_p & v8455ab | !hgrant0_p & !v372b351;
assign v373375c = hmaster0_p & v3a5d678 | !hmaster0_p & v3736a75;
assign v3743851 = hgrant4_p & v374d47d | !hgrant4_p & v3747800;
assign v3a711ec = hmaster2_p & v8455ab | !hmaster2_p & !v372cc25;
assign v37405a7 = stateG2_p & v8455ab | !stateG2_p & v3778565;
assign v374a0b1 = hbusreq5_p & v3779403 | !hbusreq5_p & v37342e7;
assign v375b737 = hbusreq1 & v3a7057b | !hbusreq1 & !v8455ab;
assign v3a6d88e = hgrant5_p & v372f55a | !hgrant5_p & v3764005;
assign v3a7162f = hmaster2_p & v3749437 | !hmaster2_p & v37786a6;
assign v374d258 = hlock8 & v3a70f61 | !hlock8 & v3a63b26;
assign v375e262 = hbusreq4_p & v37654f4 | !hbusreq4_p & v8455ab;
assign v23fd8c6 = hmaster2_p & v37343bc | !hmaster2_p & v3764d0b;
assign v3a59431 = hmaster0_p & v3a57584 | !hmaster0_p & v3730e75;
assign dc6ded = hlock6 & v372495f | !hlock6 & v3754b61;
assign v39a4c67 = hgrant4_p & v37796ce | !hgrant4_p & v373facf;
assign v375e12d = hlock6 & v373601e | !hlock6 & v3734db5;
assign v3a706e6 = hbusreq7_p & v1e378a8 | !hbusreq7_p & v3a57f7d;
assign v372a246 = hmaster2_p & v3748451 | !hmaster2_p & v37784b9;
assign v37718fb = hready & v3765f9e | !hready & !v3a5cf0b;
assign v3a70fca = hmaster1_p & v3a6ba08 | !hmaster1_p & v3757a04;
assign v372b6ec = hbusreq0 & v35b71af | !hbusreq0 & v3747d58;
assign v375352f = hgrant4_p & v8455ab | !hgrant4_p & v3a6a934;
assign v377ed24 = hbusreq0 & v3755928 | !hbusreq0 & v3a701ab;
assign v37290ab = hmaster0_p & v8455ab | !hmaster0_p & v375b019;
assign v3a7008f = hbusreq5 & v3727363 | !hbusreq5 & v37316cb;
assign v3736d03 = hgrant6_p & v3774c1b | !hgrant6_p & v377e545;
assign v3a70895 = hgrant0_p & v8455ab | !hgrant0_p & v3744bac;
assign v3729186 = hbusreq4 & v37bfc8c | !hbusreq4 & v8455ab;
assign v3a5a8f6 = hlock7_p & v3a66a8e | !hlock7_p & v37795eb;
assign v377e5ac = hmaster2_p & v3a6fa93 | !hmaster2_p & v37380c4;
assign v377c7c0 = hbusreq3_p & v375d304 | !hbusreq3_p & v8455ab;
assign v3a67a02 = hlock7_p & v3a6f317 | !hlock7_p & v377632d;
assign v3743da3 = hlock6_p & v3774a7e | !hlock6_p & v375e9a7;
assign v373f5d3 = hgrant3_p & v37645ec | !hgrant3_p & v3a6eb62;
assign v3a55d66 = hbusreq1_p & v3778176 | !hbusreq1_p & v8455ab;
assign v3747892 = hmaster2_p & v3a55d66 | !hmaster2_p & v3a6a261;
assign v3a60077 = hbusreq4_p & v377cfd9 | !hbusreq4_p & !v372ee7e;
assign v3807386 = hmaster1_p & v375dd87 | !hmaster1_p & v3724b5a;
assign v3a60103 = hbusreq4 & v3a5ba1a | !hbusreq4 & v3a6f994;
assign v3a55076 = hbusreq8 & v3735d01 | !hbusreq8 & v3a60276;
assign v3a6f345 = hmaster1_p & v374e033 | !hmaster1_p & v373ec60;
assign v377a8c3 = hbusreq5 & v3a66aa4 | !hbusreq5 & v3a71530;
assign v3a66014 = hbusreq6 & v3767f33 | !hbusreq6 & v8455e7;
assign v376fafe = hbusreq6_p & v3767420 | !hbusreq6_p & v35772a6;
assign v3a6eba9 = hbusreq0 & v3a6f07e | !hbusreq0 & v3733542;
assign v3728034 = hbusreq4 & v373f9db | !hbusreq4 & v373484e;
assign v374dae3 = hmaster3_p & v3727477 | !hmaster3_p & v8455ab;
assign v3a58792 = hmaster3_p & v8455ab | !hmaster3_p & !v3a6fb41;
assign v372c2bf = hgrant4_p & v3759d08 | !hgrant4_p & v3753eb3;
assign v37308a9 = hbusreq0 & v3748ba4 | !hbusreq0 & v374ed57;
assign v3740fef = hbusreq2 & v3a6f9c3 | !hbusreq2 & v8455bf;
assign v376d258 = hbusreq8 & v37644ee | !hbusreq8 & v373a005;
assign v3751d87 = hgrant0_p & v3a713fb | !hgrant0_p & v360d0a7;
assign v377fc15 = hgrant6_p & v3770c9d | !hgrant6_p & v3a56338;
assign v3732759 = hgrant2_p & v3758472 | !hgrant2_p & !v3a63329;
assign v3a69923 = hbusreq5_p & v3a635ea | !hbusreq5_p & v3a5ba93;
assign v372c60a = hbusreq2 & v3760ab8 | !hbusreq2 & v377caa3;
assign v37399b4 = hbusreq2 & v377c7c0 | !hbusreq2 & v377b774;
assign v3723fec = hmaster2_p & v8455ab | !hmaster2_p & v3a5b978;
assign v375722a = hbusreq8 & v8455e7 | !hbusreq8 & v3a702f0;
assign v3752d24 = hlock5_p & v3a5cc79 | !hlock5_p & !v8455ab;
assign v372c6b3 = hbusreq8_p & v3a6f684 | !hbusreq8_p & v8455ab;
assign v3732d82 = hlock6 & v3744877 | !hlock6 & v37688df;
assign v3a6f8c0 = hmaster1_p & v372a24d | !hmaster1_p & v377535e;
assign v3a69eb7 = hbusreq6 & v37414ed | !hbusreq6 & v8455ab;
assign v39eb590 = hbusreq6_p & v3729801 | !hbusreq6_p & v8455ab;
assign v3a6fdc5 = hgrant3_p & v8455ab | !hgrant3_p & v373a3dd;
assign v374cfd8 = hbusreq5_p & v376e0f5 | !hbusreq5_p & !v8455ab;
assign v377a180 = hlock4 & v3a60103 | !hlock4 & v3a5ba1a;
assign v3726f10 = hbusreq6_p & v373e877 | !hbusreq6_p & v3736fc4;
assign v3a6f9d1 = hbusreq4 & v373dd66 | !hbusreq4 & v8455ab;
assign v3a6c42b = jx1_p & v3753f59 | !jx1_p & v3a7109b;
assign v377ba41 = hmaster2_p & v376a6f1 | !hmaster2_p & v375e53a;
assign v376ef3d = hmaster1_p & v3754a39 | !hmaster1_p & v8455ab;
assign v3a5965e = hmaster1_p & v3726357 | !hmaster1_p & v3a64641;
assign v375021b = hbusreq2 & v37383f6 | !hbusreq2 & v37366b5;
assign v3740152 = hbusreq1_p & v37393f0 | !hbusreq1_p & v373217b;
assign v372766c = jx1_p & v372b715 | !jx1_p & v37676e0;
assign v3a70448 = hmaster0_p & v37790c6 | !hmaster0_p & v8455ab;
assign v3808fc8 = hmaster0_p & v377d1dc | !hmaster0_p & a7394c;
assign v3a5e3d0 = hbusreq0_p & v375356f | !hbusreq0_p & v3a551a4;
assign v37447bf = hgrant0_p & v8455ab | !hgrant0_p & v8455b6;
assign v372f4ea = hmaster2_p & v3a70fb2 | !hmaster2_p & v3768685;
assign v39eb1dc = hmaster3_p & v37415e4 | !hmaster3_p & v374a516;
assign v3a6fc33 = hmaster1_p & v372ef39 | !hmaster1_p & b52e7d;
assign v375b142 = hbusreq6_p & v3726c67 | !hbusreq6_p & v3731383;
assign v373b6ca = hbusreq2_p & v374bf71 | !hbusreq2_p & v1e3755f;
assign v37735b8 = hmaster0_p & v3a710e3 | !hmaster0_p & v375f847;
assign v3a712e2 = hgrant4_p & v3a5fc34 | !hgrant4_p & v3807604;
assign v3757009 = hgrant6_p & v8455ab | !hgrant6_p & v373f492;
assign v3a6ac26 = stateA1_p & v2aca977 | !stateA1_p & v2acb5a2;
assign v3773a6b = hgrant2_p & v37598ab | !hgrant2_p & v3a709c4;
assign v375f95f = hmaster2_p & v3a5a510 | !hmaster2_p & !v3735e39;
assign v3747a0e = hlock6 & v3774df9 | !hlock6 & v3a646fb;
assign v3a5ab05 = hmaster2_p & v3a6f880 | !hmaster2_p & v8455ab;
assign v3771a62 = hbusreq5_p & v372a9a5 | !hbusreq5_p & v37390d5;
assign v3740404 = hmaster2_p & v8455ab | !hmaster2_p & v360bc71;
assign v3737462 = hbusreq1_p & v3a6fd6f | !hbusreq1_p & v35772a6;
assign v3a6f622 = hbusreq7 & v3a713d2 | !hbusreq7 & v3a70d99;
assign v3778528 = locked_p & v372a023 | !locked_p & v8455ab;
assign v375d078 = hmaster0_p & v374b35e | !hmaster0_p & v372c14d;
assign v3a6f90c = hmaster2_p & v3a70c19 | !hmaster2_p & v3758ab0;
assign v3771e6d = hbusreq5 & v3a2976f | !hbusreq5 & v1e37407;
assign v3a62f13 = hlock6 & v375b90a | !hlock6 & v374f351;
assign v3a6fc63 = hbusreq2 & v3a689eb | !hbusreq2 & v8455ab;
assign v3765b09 = hbusreq3_p & v3a6ebf1 | !hbusreq3_p & !v8455ab;
assign v3a69c7b = hlock7_p & v377beee | !hlock7_p & v372fade;
assign v373cb82 = jx0_p & v375b0f9 | !jx0_p & v3a5d51a;
assign v3a71682 = hgrant0_p & v374c01f | !hgrant0_p & v373905f;
assign v37623f5 = hmaster0_p & v3756ef1 | !hmaster0_p & v3728813;
assign v376c047 = hmaster2_p & v3a6ffae | !hmaster2_p & v35772a6;
assign v373a2fc = stateG10_1_p & v8455ab | !stateG10_1_p & v373d4e8;
assign v37691fa = hbusreq2_p & v3a5d555 | !hbusreq2_p & !v380a1a6;
assign v3a5b070 = hmaster1_p & v3742c62 | !hmaster1_p & v3808fc8;
assign v3a6f25b = hbusreq7 & v3a7159f | !hbusreq7 & v3a671f2;
assign v3a70006 = hbusreq6_p & v376b21a | !hbusreq6_p & v3a5e748;
assign v376bf97 = hmaster2_p & v8455ab | !hmaster2_p & !v2678c40;
assign v373899b = hgrant4_p & v3739896 | !hgrant4_p & v3764381;
assign v37410d9 = hbusreq3 & v37566b2 | !hbusreq3 & !v8455ab;
assign v37751bb = hmaster1_p & v3a5a510 | !hmaster1_p & v374cceb;
assign v374355f = hbusreq4_p & v373127e | !hbusreq4_p & v3a6fc2f;
assign v376e513 = hlock4_p & v37315da | !hlock4_p & v8455b0;
assign v37507d6 = hmaster2_p & v375d4e5 | !hmaster2_p & v373bf45;
assign v3a561aa = hlock5_p & v376f9ca | !hlock5_p & !v8455ab;
assign v377adaa = hgrant5_p & v377a522 | !hgrant5_p & v376596e;
assign v372efee = hmaster2_p & v37651c2 | !hmaster2_p & v374af22;
assign v3763150 = hlock0 & v3a64af7 | !hlock0 & v3725cc8;
assign v3a65384 = hgrant6_p & v8455ab | !hgrant6_p & v3a6eec2;
assign v376ab5d = hbusreq4_p & v3a6851f | !hbusreq4_p & v3a5e5f3;
assign v37334c2 = hbusreq8_p & v3a6f41f | !hbusreq8_p & !v8455ab;
assign v373ce4e = hmaster0_p & v3a5a807 | !hmaster0_p & v3a6d9ac;
assign v3728a6a = hbusreq4 & v376eeea | !hbusreq4 & v8455ab;
assign v33789b9 = hbusreq0 & v375add0 | !hbusreq0 & v3744452;
assign v3777825 = hbusreq5 & v3a5cc14 | !hbusreq5 & v377c174;
assign v375b506 = hgrant3_p & v377dd3b | !hgrant3_p & v37361aa;
assign v3776e5b = hbusreq4_p & v376e033 | !hbusreq4_p & v376ab51;
assign v3a54350 = hgrant4_p & v37510a5 | !hgrant4_p & v3806b78;
assign v37776c8 = hgrant5_p & v8455ab | !hgrant5_p & v3a6faaa;
assign v377bd79 = hbusreq6_p & v376ca93 | !hbusreq6_p & v373a542;
assign v3738061 = hgrant4_p & v3a70230 | !hgrant4_p & v375f88a;
assign v376ce4d = hbusreq4_p & v373f52e | !hbusreq4_p & v8455b0;
assign v37331e1 = hbusreq7 & v37581f6 | !hbusreq7 & v374dfe3;
assign v3a6b714 = hbusreq2 & v3a6bd87 | !hbusreq2 & !v8455ab;
assign v377eab5 = hbusreq5_p & v3745871 | !hbusreq5_p & v376af8d;
assign v3736b93 = hgrant5_p & v377cdf1 | !hgrant5_p & v3a680eb;
assign v374abee = hmaster2_p & v376025f | !hmaster2_p & v8455ab;
assign v3725149 = hbusreq4_p & v3778921 | !hbusreq4_p & v3a6ebf2;
assign v3a6fc01 = hbusreq0 & v3a636a7 | !hbusreq0 & v3755ed8;
assign v37614a9 = hbusreq7_p & a0a219 | !hbusreq7_p & v377ccb7;
assign v3a7152a = hbusreq5 & v376a2de | !hbusreq5 & v373a6d9;
assign v3732bf9 = hmaster2_p & v3a635ea | !hmaster2_p & v376c7d1;
assign v3a701ab = hgrant6_p & v3a6ffb6 | !hgrant6_p & v375602e;
assign v372cdde = hbusreq5_p & v8455ab | !hbusreq5_p & v375058e;
assign v3a6fd65 = hgrant2_p & v375975b | !hgrant2_p & v3a68b74;
assign v3a6467a = hbusreq2 & v3768ecc | !hbusreq2 & v8455e7;
assign v3a5cb2c = hmaster0_p & v37285c9 | !hmaster0_p & v8455ab;
assign v3a70a65 = hmaster0_p & v375fc83 | !hmaster0_p & v3a5c026;
assign v3738602 = hbusreq6_p & v374faa9 | !hbusreq6_p & v377661c;
assign v3a71076 = hmaster1_p & v3a69de7 | !hmaster1_p & v373a57d;
assign v380985a = jx0_p & v3743e3c | !jx0_p & v3a6a25c;
assign v375646d = hready & v3a66651 | !hready & v8455ab;
assign v3a6cce9 = hlock8 & v37741d7 | !hlock8 & v3743b2f;
assign v37315d0 = hmaster2_p & v3a707f2 | !hmaster2_p & v3a6eaff;
assign v3749d74 = hgrant2_p & v3734967 | !hgrant2_p & v3763c82;
assign v37738fc = hbusreq1_p & v3752a45 | !hbusreq1_p & v8455ab;
assign v373a158 = hbusreq4_p & v373c3ba | !hbusreq4_p & v3742b54;
assign v376d68d = hmaster0_p & v3a6c4e4 | !hmaster0_p & v3767dc8;
assign v3a66316 = hbusreq0 & v3a70f28 | !hbusreq0 & v3743fe3;
assign v3a709a4 = hbusreq6 & v376dcd0 | !hbusreq6 & !v3a57aad;
assign v3728fb5 = hgrant0_p & v8455ab | !hgrant0_p & v3a6a7a1;
assign v3751d9c = hbusreq5_p & v373899b | !hbusreq5_p & v3756ef1;
assign v3a6f2dd = hgrant0_p & v3727517 | !hgrant0_p & v3776670;
assign v375f0de = hbusreq7 & v3a6f873 | !hbusreq7 & v37775c7;
assign v376b23a = hgrant0_p & v376dfed | !hgrant0_p & v3731b88;
assign v3a67092 = hmaster0_p & v3a54b31 | !hmaster0_p & d26e1e;
assign v3a683d9 = hmaster0_p & v3a6ffb6 | !hmaster0_p & v377ba78;
assign v3a5a496 = hburst0_p & v8455ab | !hburst0_p & v8455d7;
assign v3736a9a = hgrant2_p & v8455ab | !hgrant2_p & v377ab2c;
assign v3749001 = hbusreq4 & v373997b | !hbusreq4 & v35b774b;
assign v3740f7e = hlock5_p & v3a6f443 | !hlock5_p & !v377a92d;
assign v37302b7 = hmaster1_p & v376e72d | !hmaster1_p & v3743f3b;
assign v372eeda = hbusreq0 & afa7f5 | !hbusreq0 & v8455ab;
assign v3769010 = hgrant2_p & v3a702a0 | !hgrant2_p & v3741a9b;
assign v375a750 = hlock6_p & v3a68838 | !hlock6_p & v8455b0;
assign v3755113 = hmaster0_p & v3a70bcb | !hmaster0_p & v8455ab;
assign v3a5ffdd = hmaster2_p & v8455ab | !hmaster2_p & v373f72a;
assign v3a70db3 = hmaster0_p & v373014d | !hmaster0_p & v3a67462;
assign v372ab46 = hbusreq2_p & v8455b3 | !hbusreq2_p & v3767437;
assign v3a67a6f = hbusreq4_p & v3a5d94a | !hbusreq4_p & !v8455ab;
assign v3778a91 = jx0_p & v37231e5 | !jx0_p & !v373327e;
assign v3731c4b = hlock4_p & v2aca977 | !hlock4_p & v8455ab;
assign v3779288 = hmaster0_p & v3a5af94 | !hmaster0_p & v37489a0;
assign v3751c68 = hbusreq6_p & v2aca977 | !hbusreq6_p & v3a6ee22;
assign v373b647 = hbusreq8_p & v3737808 | !hbusreq8_p & v37628f3;
assign v374fe73 = hgrant2_p & v37320bb | !hgrant2_p & v374e753;
assign v23fd9e1 = hmaster0_p & v3760a52 | !hmaster0_p & v373a759;
assign v372e0fc = hgrant5_p & v8455ab | !hgrant5_p & v3724936;
assign v3a56dd5 = hgrant2_p & v8455b0 | !hgrant2_p & v375e5d4;
assign v3a6e221 = hbusreq8_p & v3738c33 | !hbusreq8_p & v3a6ed49;
assign v372de1e = hbusreq0 & v377598f | !hbusreq0 & v374baea;
assign v3a705bc = hbusreq4_p & v373e814 | !hbusreq4_p & v372d967;
assign v3a6dbec = hbusreq8 & v3a620f2 | !hbusreq8 & v373c3ac;
assign v39eb44a = hmaster0_p & v37354c1 | !hmaster0_p & !v3771e23;
assign v377bf9f = hgrant6_p & v3772362 | !hgrant6_p & a89e0c;
assign v376adaf = hlock6 & v37352a5 | !hlock6 & v372e6f4;
assign v37c101a = hlock1_p & v375b265 | !hlock1_p & v3729bd7;
assign v373924d = hmaster2_p & v375ced2 | !hmaster2_p & v375444a;
assign v3760d8d = hbusreq6 & v376cad6 | !hbusreq6 & v376bade;
assign v37373bb = hmaster0_p & v3750f4c | !hmaster0_p & v3769923;
assign v3a7135e = hmaster1_p & v3a5fe3c | !hmaster1_p & v3a7005d;
assign v376ab0f = hgrant5_p & v372dd77 | !hgrant5_p & v3a71309;
assign v3a551e4 = hbusreq2_p & v3a6f949 | !hbusreq2_p & v374abc9;
assign v3a6f138 = hbusreq4_p & v3751081 | !hbusreq4_p & v3a5bb64;
assign v37744a3 = hmaster0_p & v372fd00 | !hmaster0_p & v37665c5;
assign v3775e46 = jx0_p & v37370f1 | !jx0_p & v3a706ba;
assign v3736d5e = hmaster2_p & v3779060 | !hmaster2_p & v3a6f43e;
assign ab4f60 = hmaster1_p & v375d078 | !hmaster1_p & v3a60e4c;
assign v23fdc4f = hbusreq5 & v377dc65 | !hbusreq5 & v372d92b;
assign v3a70906 = hgrant6_p & v3753bac | !hgrant6_p & v3a6fc11;
assign v3a6ff9f = hlock4_p & v3759c5d | !hlock4_p & v3a6fe46;
assign v3a7080c = hbusreq5_p & v3778998 | !hbusreq5_p & v3a65607;
assign v3a612af = hlock4 & v37570db | !hlock4 & v377b67d;
assign v37722c4 = hbusreq2_p & v3a6fc17 | !hbusreq2_p & v3a6f032;
assign v372b96c = hbusreq4_p & v3a65a19 | !hbusreq4_p & v3744f86;
assign v3a64082 = hmaster0_p & v37430c6 | !hmaster0_p & v375d8a6;
assign v376a87f = hbusreq5 & v3a70c8c | !hbusreq5 & v3777f05;
assign v373b31d = hbusreq1_p & v3758ef5 | !hbusreq1_p & !v8455ab;
assign ab15ca = hmaster2_p & v3a6ffd3 | !hmaster2_p & v37745a0;
assign v3a2a0f9 = hmaster2_p & v3a61a7f | !hmaster2_p & v3747302;
assign v376d780 = hmaster2_p & v3764881 | !hmaster2_p & !v3752fbc;
assign v3a70415 = hlock1_p & v2ff9190 | !hlock1_p & v8455ab;
assign v3a6e52e = hmaster0_p & v37640e9 | !hmaster0_p & v375f94a;
assign v3775fa5 = hmaster0_p & v37418dc | !hmaster0_p & v37662e7;
assign v337907e = hbusreq3 & v3728fb5 | !hbusreq3 & v3a68523;
assign v3a6af83 = hmaster2_p & v3735417 | !hmaster2_p & v3752a0d;
assign v3a70e09 = hbusreq7_p & v8455c7 | !hbusreq7_p & v375e813;
assign v3a6f62b = hmaster2_p & v3a5c640 | !hmaster2_p & v374e855;
assign v3771360 = hgrant6_p & v377b6ce | !hgrant6_p & v377754d;
assign v3a70e97 = hbusreq4 & v3a614cb | !hbusreq4 & v3a635ea;
assign v3a6fdf4 = hgrant3_p & v8455be | !hgrant3_p & v374005b;
assign v3776c95 = hmaster2_p & v3738855 | !hmaster2_p & v3746caf;
assign v3a703cd = hlock4 & v37355ce | !hlock4 & v3a6c1ec;
assign v37579f7 = hlock5 & v3751261 | !hlock5 & v3764910;
assign v3a70c12 = hmaster0_p & v37430c6 | !hmaster0_p & v37787d1;
assign v3a701ee = hbusreq7 & v37276a0 | !hbusreq7 & v380735e;
assign v3a704be = hlock5_p & v8455e7 | !hlock5_p & !v375792c;
assign v3746df7 = hbusreq8 & v3a55fe8 | !hbusreq8 & v3a6f1e8;
assign v372a406 = hgrant3_p & v8455ab | !hgrant3_p & v2093127;
assign v3a6f0a9 = hgrant3_p & v35b7299 | !hgrant3_p & !v3768933;
assign v37427cf = hbusreq3_p & v3a6fc29 | !hbusreq3_p & !v374d654;
assign v375b64b = hgrant6_p & v3737223 | !hgrant6_p & v374b0a9;
assign v37684a8 = hgrant6_p & v8455ab | !hgrant6_p & v3a703d3;
assign v37440c0 = hmaster2_p & v3a6e6fa | !hmaster2_p & v377ad76;
assign v3a5600a = hready & v3726dfa | !hready & v37295fe;
assign v3757568 = locked_p & v37403cf | !locked_p & v3a6e7b3;
assign v3779aa8 = hmaster0_p & v3a58e93 | !hmaster0_p & v3771e23;
assign d35b26 = hbusreq2_p & v376021f | !hbusreq2_p & v3a6ee06;
assign v37425c6 = hbusreq0 & v3a702c2 | !hbusreq0 & v3a6fd81;
assign v3a6ff2e = hmaster1_p & v3726ba5 | !hmaster1_p & v3a5fe51;
assign v3758a7b = hbusreq0 & v3a706e2 | !hbusreq0 & v1e37cd6;
assign v376cfd9 = hmaster2_p & v8455ab | !hmaster2_p & v375d616;
assign v3772318 = hbusreq5 & v3a56ba2 | !hbusreq5 & v3742c68;
assign v3a630b7 = hbusreq4_p & v3a635ea | !hbusreq4_p & v376bade;
assign v360d0a9 = hmaster0_p & v3a6fa3a | !hmaster0_p & v3a6cf46;
assign v3764a16 = hgrant3_p & v3754e5a | !hgrant3_p & v375d7b6;
assign v3748016 = hgrant4_p & v8e4f94 | !hgrant4_p & v3765758;
assign v375243f = hmaster0_p & v37283c0 | !hmaster0_p & v3a68426;
assign v3a70377 = hmaster0_p & v3728d9c | !hmaster0_p & v375899a;
assign v3a6fb30 = hbusreq6_p & v376fbd0 | !hbusreq6_p & !v8455ab;
assign v373301a = hbusreq5 & a19873 | !hbusreq5 & v376502e;
assign v37591e8 = hmaster0_p & v3a5a868 | !hmaster0_p & !v3746ea0;
assign v3778657 = hbusreq5_p & v3a706b3 | !hbusreq5_p & v377a9e2;
assign v3748db2 = hmaster2_p & v3a65dcf | !hmaster2_p & v8455ab;
assign v3764869 = hbusreq5_p & v3742649 | !hbusreq5_p & v37366d5;
assign v3a58a34 = hmaster2_p & v3a70e2e | !hmaster2_p & v372a0b0;
assign v373561e = hgrant4_p & v8455ab | !hgrant4_p & v3a6f9d9;
assign v3a6aa8d = jx0_p & v3756531 | !jx0_p & v372b34d;
assign v3773262 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3a70674;
assign v375b203 = hgrant0_p & v3759c2e | !hgrant0_p & !v360d0a7;
assign v373121b = hlock8 & v377d9fa | !hlock8 & v3a5ee7a;
assign v3736d0d = hmaster0_p & v374f307 | !hmaster0_p & v376af20;
assign v372c37f = hbusreq6 & v376b21a | !hbusreq6 & !v8455ab;
assign v3762a37 = hmaster2_p & v37583be | !hmaster2_p & !v377df2e;
assign v3a6f790 = hmaster0_p & v3a58ddb | !hmaster0_p & v3775c6e;
assign v372a837 = hbusreq1 & v3a6a939 | !hbusreq1 & v8455ab;
assign v3735fee = hlock0_p & v372b351 | !hlock0_p & v37266e1;
assign v3a65f0f = hlock3_p & v3a69d06 | !hlock3_p & !v8455ab;
assign v37574c0 = hmaster2_p & v375b429 | !hmaster2_p & v37624a2;
assign v37787ac = hbusreq5_p & v3728a3d | !hbusreq5_p & v372587b;
assign v373a0dc = hbusreq5_p & v3a68525 | !hbusreq5_p & v3a570ee;
assign v3758b3f = hlock0_p & v3767f33 | !hlock0_p & v3728e09;
assign v374f749 = hbusreq7_p & v376ef47 | !hbusreq7_p & v373c38b;
assign v376eaf1 = hmaster2_p & v3807f45 | !hmaster2_p & v3809ebc;
assign v377e59a = hmaster0_p & v377817b | !hmaster0_p & v372f59c;
assign v374ab4c = hbusreq7_p & v35b7734 | !hbusreq7_p & v372c09e;
assign v3742825 = jx0_p & v3734c16 | !jx0_p & v3a6f7a7;
assign v3a712bb = hmaster1_p & v3a702be | !hmaster1_p & v38064e3;
assign v3a70bcb = hmaster2_p & v3764825 | !hmaster2_p & v8455ab;
assign v373afb4 = hlock3_p & v8455ab | !hlock3_p & v3771ce2;
assign c8e1cc = jx0_p & v376e587 | !jx0_p & v375ce2d;
assign v372a53e = hmaster2_p & v3742cd4 | !hmaster2_p & v3a70ba8;
assign v376739f = hmaster2_p & v372673d | !hmaster2_p & v377d74c;
assign ae4185 = hbusreq5_p & v3a70cf4 | !hbusreq5_p & v3a61b59;
assign v3a70bd6 = hbusreq2_p & v35b774b | !hbusreq2_p & v9ed516;
assign v373432d = hlock8 & v374d31a | !hlock8 & v374c576;
assign v3a642ab = hmaster1_p & v3763571 | !hmaster1_p & v3a298b6;
assign d4de60 = hgrant2_p & v37283fc | !hgrant2_p & c58ea1;
assign v377233c = hbusreq5_p & v374c9ab | !hbusreq5_p & v8455ab;
assign v3a6d0ef = hbusreq1_p & v39e9c6f | !hbusreq1_p & v376cf85;
assign v376bf83 = hmaster0_p & v37230ec | !hmaster0_p & v3a5cdc1;
assign v3a6f7ee = hmaster2_p & v377d232 | !hmaster2_p & v3807686;
assign v3808899 = hmaster0_p & v3a70853 | !hmaster0_p & v375f94a;
assign v3a7129d = hmaster1_p & v375585e | !hmaster1_p & v374b36f;
assign v372c6cb = hbusreq2_p & v2aca978 | !hbusreq2_p & v8455ab;
assign v376b67d = hmaster0_p & v37430c6 | !hmaster0_p & v3751004;
assign v37516cc = hbusreq2_p & v37625a8 | !hbusreq2_p & !v2092faa;
assign v376cff4 = hmaster1_p & v373bbd0 | !hmaster1_p & v377b8fb;
assign v375e051 = hmaster2_p & v375a10d | !hmaster2_p & v3753dab;
assign v376afff = hbusreq5 & v3a6fb9f | !hbusreq5 & v8455ab;
assign v3a5c4c6 = hmaster0_p & v376053f | !hmaster0_p & v3a6fb52;
assign v373dd66 = hlock4_p & v376b11a | !hlock4_p & v373dd77;
assign v372e499 = hmaster0_p & v375a03b | !hmaster0_p & v372529a;
assign v3a704e7 = hlock4 & v377870b | !hlock4 & v377d9bb;
assign v373e0d3 = hbusreq0 & v372baaf | !hbusreq0 & v372818d;
assign v3a58762 = hbusreq2_p & v375c705 | !hbusreq2_p & v377e39f;
assign v373eff1 = hmaster2_p & v37737aa | !hmaster2_p & v9f823e;
assign v3755aca = hmaster0_p & v37369d7 | !hmaster0_p & v377cccb;
assign v3a70ff7 = hlock5_p & v8455ab | !hlock5_p & v375a12e;
assign v374e20c = hlock3_p & v3747c3e | !hlock3_p & v8455ab;
assign v376c777 = hbusreq0_p & v3a635ea | !hbusreq0_p & v3a6f757;
assign v3a6fb5a = hmaster0_p & v3749d86 | !hmaster0_p & v375cdf8;
assign v374faf5 = hmaster2_p & v3747302 | !hmaster2_p & v376d1bb;
assign v37514c7 = hbusreq0 & v375911a | !hbusreq0 & v8455ab;
assign v374edd8 = hmaster0_p & v3759ad6 | !hmaster0_p & v94e9e0;
assign v3a6f55a = hmaster1_p & v3a6eecb | !hmaster1_p & !v376acd9;
assign v3a70609 = hmaster2_p & v3731210 | !hmaster2_p & v373a415;
assign v373e1d0 = hgrant4_p & v8455ab | !hgrant4_p & v3a64af7;
assign v2acb095 = hbusreq4_p & v373d262 | !hbusreq4_p & v8455ab;
assign v92aebd = hbusreq7_p & v3a53dfc | !hbusreq7_p & v372e479;
assign v37351ff = hbusreq7_p & v3763c1f | !hbusreq7_p & v375b5d6;
assign v3a713b2 = hburst0 & v3a5815e | !hburst0 & v3a70a2e;
assign v3a7041c = hbusreq7_p & v372fe28 | !hbusreq7_p & v3a715f8;
assign v3766485 = hbusreq2 & v3a6fe0d | !hbusreq2 & !v8455b5;
assign v374a11d = hmaster0_p & v3738b8a | !hmaster0_p & v8455ab;
assign v3a65ca8 = hbusreq2_p & v3764caf | !hbusreq2_p & v37677ee;
assign v37762ec = hlock7 & v37339b7 | !hlock7 & v37730b3;
assign v3a7083b = hbusreq6_p & v376944c | !hbusreq6_p & v3a5b581;
assign v37690af = hbusreq2_p & v3779227 | !hbusreq2_p & v3a6fcef;
assign v376a35c = hmastlock_p & v3a6ffe0 | !hmastlock_p & v8455ab;
assign v372773c = hmaster1_p & v375f071 | !hmaster1_p & v374c000;
assign v373cde8 = hgrant2_p & v3a6cfe0 | !hgrant2_p & v3765d2a;
assign v375cc8b = hbusreq5 & v376581d | !hbusreq5 & v3738726;
assign v3a6b46d = hlock4 & v37263b9 | !hlock4 & v3a5e10c;
assign v3a65acb = hbusreq8 & v373ddfc | !hbusreq8 & v374214d;
assign v372c8d0 = hmaster0_p & v372c00b | !hmaster0_p & v372d9ae;
assign v37270bc = hbusreq0 & v376ffbf | !hbusreq0 & v3a64e2a;
assign v3a5d9e7 = hbusreq4_p & v37728a5 | !hbusreq4_p & v3a70d99;
assign v373a3fa = hgrant4_p & v3735cb3 | !hgrant4_p & v377dae8;
assign v37574b0 = hbusreq6_p & v3a6e6c9 | !hbusreq6_p & v8455ab;
assign v3a71535 = hmaster1_p & v376640a | !hmaster1_p & v8455ab;
assign v3a68822 = hgrant6_p & v374510e | !hgrant6_p & v3a714e9;
assign v374743d = hgrant4_p & v3763b9b | !hgrant4_p & v3a701a0;
assign v3a6fb57 = hmaster2_p & v3a635ea | !hmaster2_p & v372e711;
assign v372fe5f = hbusreq0_p & v3a6bddd | !hbusreq0_p & v373b288;
assign v37294db = hlock0 & v373abde | !hlock0 & v3a6af67;
assign b02944 = hmaster1_p & v372a93f | !hmaster1_p & v3728040;
assign v3a70cb2 = hmaster0_p & v37498bd | !hmaster0_p & v3a6ff47;
assign v376ba4d = hbusreq2 & v3806db7 | !hbusreq2 & v372fba5;
assign v377a369 = hmaster2_p & v3a6c5ee | !hmaster2_p & v3a57959;
assign v373f6ee = hbusreq6_p & v3a6fb71 | !hbusreq6_p & v8455ab;
assign v3746f4c = hbusreq8 & v3a6f5e4 | !hbusreq8 & v375f27b;
assign v3a66279 = hgrant6_p & v3a59b9e | !hgrant6_p & v37578a2;
assign v3726dfa = hmastlock_p & v37405a7 | !hmastlock_p & v8455ab;
assign v3729beb = hbusreq8_p & v3a6f511 | !hbusreq8_p & v23fdbce;
assign v3733726 = hgrant6_p & v8455ab | !hgrant6_p & v3a66c2f;
assign v3779544 = hbusreq6 & v3a70200 | !hbusreq6 & !v3a70caf;
assign v373506a = hbusreq0 & v3a6cc67 | !hbusreq0 & v3a6fd89;
assign v373fb42 = hbusreq7 & v376592c | !hbusreq7 & v3a712b5;
assign v374f432 = hbusreq5_p & v377a3bd | !hbusreq5_p & v372ff0a;
assign v3762fc3 = hbusreq3 & v3723b00 | !hbusreq3 & v8455ab;
assign v3a5db66 = hgrant1_p & v3743745 | !hgrant1_p & v37665bf;
assign v3a61123 = jx0_p & v377a0e7 | !jx0_p & v377a883;
assign v377e0a4 = hmaster3_p & v8455ab | !hmaster3_p & v3761340;
assign v3727363 = hmaster0_p & v372f2ed | !hmaster0_p & !v37328f1;
assign v3a70304 = hmaster2_p & v377eac7 | !hmaster2_p & v3a708a9;
assign v375ebe9 = hbusreq0 & v373de8a | !hbusreq0 & v37649a0;
assign v3771b20 = hbusreq0_p & v376a8cf | !hbusreq0_p & v3734312;
assign v375556d = hlock4_p & v3742122 | !hlock4_p & v373f058;
assign v373adaa = hmaster0_p & v375fbba | !hmaster0_p & v3741320;
assign v377882e = hgrant6_p & v8455b9 | !hgrant6_p & v3146177;
assign v3741748 = hmaster2_p & v8455c3 | !hmaster2_p & v3729f25;
assign v360d080 = hgrant2_p & v3a5f50e | !hgrant2_p & v375c771;
assign v37482f5 = hbusreq7_p & v376bfe6 | !hbusreq7_p & v373461a;
assign v3a578ef = hmaster1_p & v3775dbc | !hmaster1_p & v3762a26;
assign v375408d = hbusreq8 & v37751cb | !hbusreq8 & v3a5c733;
assign aa783c = hmaster0_p & v377108d | !hmaster0_p & v3a6aa59;
assign v3737a6e = hmaster2_p & v3a70557 | !hmaster2_p & v37745a0;
assign v3a65afa = hlock6_p & v3770116 | !hlock6_p & v3a71350;
assign v3741197 = hmaster0_p & v3a7000f | !hmaster0_p & v377e0d2;
assign v374a6fc = hbusreq2_p & v3a6467a | !hbusreq2_p & v377b4ad;
assign v38078ea = hbusreq8 & v37507a8 | !hbusreq8 & v3778211;
assign v3775d56 = hbusreq2 & v3a6fdc5 | !hbusreq2 & v3a558f6;
assign v3776ea4 = hgrant6_p & v3a70272 | !hgrant6_p & v3766345;
assign v3756d6e = hmaster1_p & v3a635ea | !hmaster1_p & v3772f74;
assign v372ea9a = hbusreq3_p & v3752c04 | !hbusreq3_p & v37467a3;
assign v3a6ab8c = hbusreq6_p & v3a6fdd8 | !hbusreq6_p & v3a710ba;
assign v35b6c3a = hbusreq5_p & v372402f | !hbusreq5_p & v8455ab;
assign v3770032 = hbusreq4_p & v3a6e31f | !hbusreq4_p & !v3a5af94;
assign v3807601 = hmaster0_p & v3a70609 | !hmaster0_p & v94e9e0;
assign v3a6367f = hmaster1_p & v3a700e2 | !hmaster1_p & v3a70bbd;
assign v2acafb4 = hmaster0_p & v3a7002c | !hmaster0_p & v377a8ea;
assign v3a5b8a2 = hmaster2_p & v374e51a | !hmaster2_p & v3a70e9e;
assign v37510e5 = hbusreq5_p & v3a6b60d | !hbusreq5_p & v3762929;
assign v377baeb = hgrant2_p & v3a5f50e | !hgrant2_p & v3a6bf86;
assign v375865a = hbusreq2_p & v3769d3e | !hbusreq2_p & v3a70f03;
assign v376894a = hmaster2_p & v377e904 | !hmaster2_p & v3a684bb;
assign v372946a = hbusreq8 & v376a383 | !hbusreq8 & v373c26c;
assign v3a6aee6 = hbusreq0 & v3729b48 | !hbusreq0 & v373bd6c;
assign v2092bcb = hlock4 & v374e3a9 | !hlock4 & v3773575;
assign v3a6cf19 = hlock2 & v3a70a4c | !hlock2 & v377881b;
assign v375a187 = hbusreq5 & v3a652b6 | !hbusreq5 & v3731d2d;
assign v372c18e = hlock6 & v38072fd | !hlock6 & v3a640ab;
assign v3737e8c = hbusreq2_p & v3747346 | !hbusreq2_p & v3a6f22f;
assign v3a54c9b = hgrant4_p & v8455c1 | !hgrant4_p & v375a637;
assign v3a69583 = hbusreq5 & v3a5b86c | !hbusreq5 & v3a5e783;
assign b46885 = hbusreq5_p & v3a67e25 | !hbusreq5_p & v8455ab;
assign v3a6f7a7 = hbusreq8_p & v3759569 | !hbusreq8_p & v3778676;
assign v3809e71 = hbusreq8_p & v3a616f0 | !hbusreq8_p & v376d191;
assign v37653d1 = hmaster2_p & v375a9d0 | !hmaster2_p & v3a6c8b4;
assign v372a5fc = hgrant6_p & v8455ab | !hgrant6_p & v374a23a;
assign v3a573c2 = hbusreq5_p & v375a16a | !hbusreq5_p & !v377a808;
assign v3743f3c = hbusreq4_p & v3a635ea | !hbusreq4_p & v37715d9;
assign v3a70eac = hmaster0_p & v377adf5 | !hmaster0_p & v37635f0;
assign ca9b68 = hmaster2_p & v23fdd06 | !hmaster2_p & v373a629;
assign v37404da = hlock6 & v373af5d | !hlock6 & v37650bd;
assign v3764ecd = hbusreq8 & v3a6c96a | !hbusreq8 & v376f51a;
assign v37606b1 = hmaster2_p & v37392ad | !hmaster2_p & !v8455ab;
assign v35b77ae = hbusreq5 & v374544c | !hbusreq5 & v3731aaf;
assign v3779cf6 = hlock5 & v3a538b3 | !hlock5 & v39372d9;
assign v376646f = hgrant4_p & v8455ab | !hgrant4_p & aa52b8;
assign v376c06f = hlock3 & v37560c7 | !hlock3 & v3730946;
assign v3739b40 = hlock2_p & v3778ed4 | !hlock2_p & v8455e7;
assign v377e976 = busreq_p & v3a6fa4f | !busreq_p & !v23fd970;
assign v3753e6a = hlock0_p & v374306c | !hlock0_p & v3a6ffae;
assign v3a63f49 = hlock7_p & v3774d2a | !hlock7_p & v377ae0c;
assign v372d59e = hgrant3_p & v8455ab | !hgrant3_p & v3727293;
assign v33790da = hgrant0_p & v8455ab | !hgrant0_p & v37241fd;
assign v2093127 = hgrant0_p & v8455ab | !hgrant0_p & !v374b4d6;
assign v37366df = jx3_p & v372e0b7 | !jx3_p & v374f048;
assign v376114f = jx1_p & v374e304 | !jx1_p & v3756bd1;
assign v3a6b5ba = hmaster0_p & v3a6e31f | !hmaster0_p & v3a6ef21;
assign v3a70bbd = hmaster0_p & v3a700e2 | !hmaster0_p & v374182b;
assign v3a55d3b = hlock0 & v377c6b3 | !hlock0 & v3a70261;
assign v3a6799a = hlock7_p & v380651a | !hlock7_p & !v3742360;
assign v3764218 = hbusreq6_p & v3a70e6f | !hbusreq6_p & v35772a6;
assign v375aa18 = hbusreq5 & v374518e | !hbusreq5 & v3758661;
assign v376f583 = hbusreq7_p & v3763c1f | !hbusreq7_p & v3a70be1;
assign v3744c88 = hbusreq5_p & v8455c6 | !hbusreq5_p & !v8455ab;
assign v3738641 = hmaster1_p & v372d8ff | !hmaster1_p & v3a5c064;
assign v3a70ed5 = hmaster1_p & v374ff15 | !hmaster1_p & v3a5b4ca;
assign v3a5ae1b = hbusreq6_p & v38072fd | !hbusreq6_p & v372c18e;
assign v3766597 = hbusreq8_p & v375a338 | !hbusreq8_p & v376550d;
assign v3a665ab = hbusreq2_p & v37c0190 | !hbusreq2_p & v3a62986;
assign v845605 = stateG3_2_p & v8455ab | !stateG3_2_p & !v8455ab;
assign v37419b4 = hmaster0_p & v375c769 | !hmaster0_p & v3a64977;
assign v3a701fa = hmaster0_p & v377b59e | !hmaster0_p & v3753b80;
assign v3727c91 = hbusreq5 & v3a5e2eb | !hbusreq5 & v3727b10;
assign v2aca81d = hbusreq5 & v3749dc1 | !hbusreq5 & v376af8d;
assign v3a71131 = hlock6 & v3748797 | !hlock6 & v3a6fa7e;
assign v3a6f61f = hgrant2_p & v375da10 | !hgrant2_p & v3a6f949;
assign v3753ee8 = hmaster1_p & v2ff9371 | !hmaster1_p & v3a557a1;
assign v374ec37 = hbusreq5_p & v37480c6 | !hbusreq5_p & v377af0b;
assign v373da33 = hmaster0_p & v3763175 | !hmaster0_p & v3747d3d;
assign v376ac74 = hbusreq4 & v3725230 | !hbusreq4 & v8455ab;
assign v3a70d6b = hgrant5_p & v3a66e3d | !hgrant5_p & v3a6f8e1;
assign v3a53f43 = hbusreq2_p & v376c02d | !hbusreq2_p & v3a699d3;
assign v3724731 = hbusreq0 & v3746d4a | !hbusreq0 & v3808fce;
assign v375cde6 = hbusreq4_p & v373583d | !hbusreq4_p & !v8455ab;
assign v8c0e15 = hbusreq1 & v3a593ee | !hbusreq1 & v37496fa;
assign v372f326 = hmaster2_p & v3762f51 | !hmaster2_p & v37229c2;
assign v3a5f8d0 = hbusreq1_p & v375cd0c | !hbusreq1_p & v8455ab;
assign v3a6fc9c = hbusreq0 & v8455b0 | !hbusreq0 & v3a708a2;
assign v3a707f6 = hbusreq6 & v3768685 | !hbusreq6 & v3a70d99;
assign v3a6fd3e = hbusreq0 & v3726f10 | !hbusreq0 & v375564e;
assign v37739c6 = hgrant6_p & v3765fcf | !hgrant6_p & !v3764218;
assign v38073bb = hmaster2_p & v3747302 | !hmaster2_p & v374db6a;
assign v3746d07 = hlock2 & v360d18d | !hlock2 & v3a6ffa0;
assign v372706f = hlock8_p & v3750b9b | !hlock8_p & v3a6f049;
assign v3a70615 = hmaster1_p & v8455ab | !hmaster1_p & v37519d9;
assign v373c9c1 = hmaster0_p & v373e74b | !hmaster0_p & v3a60195;
assign v3808943 = hbusreq7_p & v3772aa4 | !hbusreq7_p & !v374a50a;
assign v3a7067e = hlock5 & v3777b5f | !hlock5 & v375b96f;
assign v3754d28 = hlock5 & v3a6febe | !hlock5 & v3a5e9b8;
assign v3a56346 = stateA1_p & v8455ab | !stateA1_p & v375b258;
assign v3778b73 = hbusreq7_p & v373ab3d | !hbusreq7_p & v8455d3;
assign v3a66fb3 = hbusreq6_p & v3749674 | !hbusreq6_p & v3770735;
assign v376537c = hmaster0_p & v3a6e7b3 | !hmaster0_p & v3741365;
assign v3a70d30 = hbusreq5_p & v3a7070c | !hbusreq5_p & v8455ab;
assign v3a701d2 = hmaster1_p & v3a29814 | !hmaster1_p & v3a70021;
assign v3a6fd2d = hlock4_p & v3a6c23b | !hlock4_p & v3a63805;
assign v3a6f724 = hbusreq5_p & v3736421 | !hbusreq5_p & v3758532;
assign v372b0b0 = hmaster1_p & v37447b9 | !hmaster1_p & v3760c32;
assign v3756dd6 = hbusreq5 & v3a5dec3 | !hbusreq5 & !v8455b5;
assign v376ca07 = hlock0_p & v2aca784 | !hlock0_p & v3a6fcc5;
assign v3757c5c = hmaster2_p & v376a6f1 | !hmaster2_p & !v373a158;
assign v3a66988 = hbusreq7_p & v3a6f5f9 | !hbusreq7_p & v3734de2;
assign v372320e = hgrant6_p & v8455ab | !hgrant6_p & v3762fcb;
assign v3a5c2f4 = hgrant3_p & v3a5b5d3 | !hgrant3_p & !v3769157;
assign v3748194 = hbusreq6_p & v3735e39 | !hbusreq6_p & !v3a6d684;
assign v3729caa = jx0_p & v3743407 | !jx0_p & v3742cce;
assign v37487a4 = hgrant2_p & v8455ab | !hgrant2_p & v3764b3f;
assign v3a58d22 = hbusreq6 & v39a537f | !hbusreq6 & v8455ab;
assign v376053b = hmaster1_p & v3754a25 | !hmaster1_p & v372b006;
assign v3724b72 = stateA1_p & v3752b8c | !stateA1_p & !v3a54427;
assign v373f780 = hbusreq7_p & v3a60030 | !hbusreq7_p & v3766645;
assign v37284b7 = hbusreq7_p & v3a70042 | !hbusreq7_p & v3a62da7;
assign v376ee03 = hbusreq6 & v3a644e6 | !hbusreq6 & v3a59391;
assign v3730eae = hbusreq4_p & v375cd4c | !hbusreq4_p & v3808f44;
assign v3a62c49 = hgrant6_p & v8455ab | !hgrant6_p & v3725f3e;
assign v375e6b2 = hbusreq4_p & v3a6439a | !hbusreq4_p & v3746ffa;
assign v3744f6f = hmaster1_p & v374d6de | !hmaster1_p & v1e379fa;
assign v372ebbf = hbusreq4 & v377e089 | !hbusreq4 & !v8455bd;
assign v3a6e4b8 = hbusreq8 & v3747587 | !hbusreq8 & v3766472;
assign v8e4749 = hgrant6_p & v8455ab | !hgrant6_p & v376a4dd;
assign v375e1a1 = hbusreq6_p & v3a6efac | !hbusreq6_p & v37728b1;
assign v3729801 = hbusreq6 & v373ee17 | !hbusreq6 & v8455ab;
assign v3745012 = hbusreq0 & v3a70a8f | !hbusreq0 & v3755090;
assign v374188e = hbusreq6 & v3a6c82f | !hbusreq6 & v8455ab;
assign v373e679 = hbusreq8_p & v377225c | !hbusreq8_p & v3a59e1b;
assign v373765a = hbusreq8_p & v3a6f394 | !hbusreq8_p & v3a65100;
assign v3723686 = hbusreq7_p & v37661e4 | !hbusreq7_p & v8455ab;
assign v377960b = hgrant4_p & v374e849 | !hgrant4_p & v3756f17;
assign v376fb60 = hgrant4_p & v376de99 | !hgrant4_p & v3731a1f;
assign v3726bdb = hgrant5_p & v372642b | !hgrant5_p & v3737e57;
assign v373a891 = hbusreq4 & d039bc | !hbusreq4 & v8455ab;
assign v3a6ebfc = hmaster1_p & v3779071 | !hmaster1_p & v37735aa;
assign v374288a = hbusreq1_p & v1e37d3f | !hbusreq1_p & v1e38224;
assign v3747dd0 = hbusreq1_p & v373226c | !hbusreq1_p & v8455ab;
assign v374bb76 = hbusreq4_p & v3733da4 | !hbusreq4_p & v3743b9e;
assign v3a648f2 = stateG2_p & v3a5a496 | !stateG2_p & v374592e;
assign be181b = hmaster2_p & v376fb60 | !hmaster2_p & v372f853;
assign v3a6fa1c = hmaster0_p & v3a7018b | !hmaster0_p & v373a246;
assign v377ad63 = hlock5_p & v3a6fc5a | !hlock5_p & !v8455ab;
assign v3a5fcbc = hlock3 & v37560c7 | !hlock3 & v374a266;
assign v372e3d8 = hgrant6_p & v8455ab | !hgrant6_p & v37369eb;
assign v3752df5 = hmaster0_p & v377cc69 | !hmaster0_p & v3741b5e;
assign v3a70a3e = hmaster2_p & v375f2ba | !hmaster2_p & v3a711f9;
assign v3754586 = stateG10_1_p & v3a57330 | !stateG10_1_p & v3773091;
assign v372e250 = hmaster2_p & v8455b0 | !hmaster2_p & v3a6f0f6;
assign v3a655e9 = hgrant4_p & v8455c2 | !hgrant4_p & v3a6a209;
assign v3a6f1b7 = hmaster2_p & v377c931 | !hmaster2_p & v376bb26;
assign v372fd00 = hgrant4_p & v8455ab | !hgrant4_p & v3a6aabc;
assign v3a6cfe0 = hbusreq2_p & v3a70e02 | !hbusreq2_p & v376d6f9;
assign v3a6fcf3 = hbusreq4 & v3a7015f | !hbusreq4 & !v8455b9;
assign v3736cdb = hbusreq6 & v37790df | !hbusreq6 & v3a6f408;
assign v374d847 = hmaster2_p & v376773f | !hmaster2_p & v3a6f09f;
assign v372989d = hbusreq2_p & v37796c6 | !hbusreq2_p & cee4af;
assign v3a70f23 = hmaster1_p & v8455ab | !hmaster1_p & v377e310;
assign v37415b2 = hgrant3_p & v3731ffc | !hgrant3_p & v3a6f48f;
assign v35b7096 = hmaster3_p & v3a70ae5 | !hmaster3_p & v3750a17;
assign v3a55039 = hbusreq3 & v372ade8 | !hbusreq3 & v372cc25;
assign v3779613 = hbusreq5_p & v3770c99 | !hbusreq5_p & !v377300f;
assign v958697 = hgrant7_p & v8455ab | !hgrant7_p & v3a6d198;
assign v374ba88 = hmaster2_p & v37430c6 | !hmaster2_p & v373f058;
assign v3748bb7 = hgrant1_p & v8455ab | !hgrant1_p & v3748797;
assign v37289b0 = hbusreq8 & v3a6ec28 | !hbusreq8 & v3a6f847;
assign v3a6f64e = hbusreq4_p & v3a6f365 | !hbusreq4_p & v373f82c;
assign v376243f = hmaster1_p & v373ff97 | !hmaster1_p & !v3a5cf3c;
assign v39ebac7 = stateA1_p & v8455ab | !stateA1_p & v373c3bd;
assign v3a6f09f = hbusreq0 & v8455ab | !hbusreq0 & v375feba;
assign a50cea = hmaster0_p & v3a63777 | !hmaster0_p & v3723740;
assign v3a2a105 = hmaster1_p & v3725bdc | !hmaster1_p & v3763dd4;
assign v37604e9 = hbusreq2_p & v3722e5c | !hbusreq2_p & v35772a6;
assign v3a55cf3 = hbusreq8_p & v3740a1e | !hbusreq8_p & v3a6fc93;
assign v372e49a = hmaster3_p & v3a68183 | !hmaster3_p & v37518f0;
assign v373280e = hbusreq7 & v3a58673 | !hbusreq7 & v1e37943;
assign v3771394 = hbusreq4 & v3a6f0f9 | !hbusreq4 & !v8455ab;
assign v374fe54 = hgrant4_p & v8455e7 | !hgrant4_p & !v372d744;
assign v3a71528 = hlock0_p & v3a5891c | !hlock0_p & v3a66d1b;
assign v375649e = hbusreq4_p & v377d7dc | !hbusreq4_p & !v8455ab;
assign v3808f6f = hbusreq0 & v37255d9 | !hbusreq0 & !v1e37cd6;
assign v3753923 = hbusreq6 & v38090f6 | !hbusreq6 & v375de7f;
assign v37413fc = hlock6_p & v3a6ac2a | !hlock6_p & v8455ab;
assign v374a37e = hmaster1_p & v377adf5 | !hmaster1_p & v37443a2;
assign v3a622a9 = jx0_p & a61746 | !jx0_p & v3a656bd;
assign v377521b = hmaster0_p & v374f307 | !hmaster0_p & v3739f75;
assign v374f543 = hbusreq4 & v3752862 | !hbusreq4 & v8455ab;
assign v3775a4f = hlock6 & v3a6e02d | !hlock6 & v37429b9;
assign v377f37e = hgrant5_p & v375446f | !hgrant5_p & v3723df0;
assign v3a6eead = hlock2 & v3a6ddd4 | !hlock2 & v375d689;
assign v3764898 = hbusreq4 & v3734af2 | !hbusreq4 & v8455ab;
assign v372e9b1 = hbusreq8_p & v3a67eb4 | !hbusreq8_p & v376723e;
assign v3a71037 = hbusreq4 & v37285ad | !hbusreq4 & v3762502;
assign v3a29dbd = hgrant6_p & v375c7b9 | !hgrant6_p & v3a6356b;
assign v3a6f807 = hgrant3_p & v3733e9e | !hgrant3_p & v376049c;
assign v3759d41 = hbusreq0 & v37333bb | !hbusreq0 & v37393ed;
assign v374765b = hgrant2_p & v377cbad | !hgrant2_p & v377e1e8;
assign v3a705b2 = hmaster0_p & v375e183 | !hmaster0_p & !v3a6e4cd;
assign v3a5cc1a = hbusreq4 & v37482f8 | !hbusreq4 & !v37661b2;
assign v3735c5a = hlock4 & v3729ae9 | !hlock4 & v3a6eddd;
assign v37790c6 = hmaster2_p & v373bb90 | !hmaster2_p & v8455ab;
assign v376a015 = hbusreq6 & v3a7156d | !hbusreq6 & v8455ab;
assign v376f70a = hmaster2_p & v39a537f | !hmaster2_p & v37521ed;
assign v37598ab = hbusreq3_p & v3a62826 | !hbusreq3_p & v35b774b;
assign v3746a67 = hmaster0_p & v3739ab4 | !hmaster0_p & v3a65612;
assign v3746b0c = hlock7 & v373d89b | !hlock7 & v3a54769;
assign d692cc = hgrant5_p & v3759611 | !hgrant5_p & v3a680eb;
assign v3a6b090 = hbusreq5 & v9ed0ba | !hbusreq5 & v376f920;
assign v377e8da = hgrant6_p & v3a57959 | !hgrant6_p & v3a702a7;
assign v3a6faff = hmaster0_p & v37691e6 | !hmaster0_p & v3a7004b;
assign v3a5ff5a = hgrant2_p & v3807f45 | !hgrant2_p & v373568c;
assign v372eabb = hlock4_p & v2925c39 | !hlock4_p & !v8455ab;
assign v3a70fe6 = hmaster0_p & v373c828 | !hmaster0_p & v372f9cf;
assign v3a610a4 = hmaster2_p & d68a4d | !hmaster2_p & v37274c2;
assign v37347d9 = hbusreq8_p & v3a68977 | !hbusreq8_p & v374bce5;
assign v373a493 = hbusreq6 & cf45c3 | !hbusreq6 & v3a6efad;
assign acbf77 = hmaster0_p & v37731ce | !hmaster0_p & v3a66cd7;
assign v3745eab = hbusreq2 & v376495e | !hbusreq2 & v8455ab;
assign jx2 = v35d37b1;
assign v377d6fc = hmaster0_p & v3a6f6e2 | !hmaster0_p & v372e58c;
assign v374fb58 = locked_p & v8455ab | !locked_p & !v3a637dd;
assign v373e9a5 = hlock6_p & v3743da0 | !hlock6_p & v37406d2;
assign v3a714a6 = hbusreq5_p & v3742649 | !hbusreq5_p & v3a68356;
assign v3a7127e = hbusreq6_p & v3a6e6c9 | !hbusreq6_p & v374e26d;
assign v375b247 = hmaster1_p & v3753418 | !hmaster1_p & v374d042;
assign v3a707ad = hbusreq2 & v374362e | !hbusreq2 & v8455ab;
assign v373343b = hgrant6_p & v377938d | !hgrant6_p & v3769f88;
assign v372ea48 = hlock4_p & v23fe06e | !hlock4_p & v377c57a;
assign v96f7ab = hmaster0_p & v3a7097c | !hmaster0_p & !v3733cd1;
assign v3a614a1 = hmaster2_p & v3a70374 | !hmaster2_p & v375f9e9;
assign v3772590 = hbusreq8 & v3a7024a | !hbusreq8 & v3a6feab;
assign v23fe061 = hbusreq4_p & v374f0c1 | !hbusreq4_p & v377cbc9;
assign v3a7135a = hbusreq8_p & v3756202 | !hbusreq8_p & v3738f1b;
assign v373240c = hmaster0_p & v373e6d2 | !hmaster0_p & v3a705e2;
assign v375f4c8 = hlock3_p & v3a6fcfe | !hlock3_p & v376430b;
assign v375bd53 = hgrant2_p & v8455ab | !hgrant2_p & v3a5f4ff;
assign v374ec57 = hbusreq5_p & v375471b | !hbusreq5_p & v3731999;
assign v376374b = hmaster2_p & v3a70f68 | !hmaster2_p & v3770b26;
assign v3728196 = hlock4_p & v3a56642 | !hlock4_p & adf78a;
assign v3734632 = hbusreq8_p & v37429d9 | !hbusreq8_p & v3a6e614;
assign v3761470 = hbusreq6 & v3a64ee3 | !hbusreq6 & v8455ab;
assign v3a66335 = hbusreq5_p & v3741d83 | !hbusreq5_p & v373d8d8;
assign v375b429 = hlock1_p & v3755002 | !hlock1_p & !v8455ab;
assign v3a6297f = hgrant4_p & v3a65053 | !hgrant4_p & v37592a3;
assign v3a53877 = hbusreq1 & v39a537f | !hbusreq1 & !v8455ab;
assign v379318b = hmaster2_p & v3377c6c | !hmaster2_p & v3751cd1;
assign v3a5dcd4 = hbusreq7_p & v3a70d4e | !hbusreq7_p & v991591;
assign v3a6d1b9 = hbusreq0 & v3a70ff1 | !hbusreq0 & v373d7ea;
assign v3769e3a = hgrant6_p & v8455ab | !hgrant6_p & v3807341;
assign v3a65b3e = hgrant5_p & v9d4353 | !hgrant5_p & v37533e5;
assign v3764586 = hmaster2_p & v3734827 | !hmaster2_p & v374fc82;
assign v3748d2f = hmaster0_p & v3766462 | !hmaster0_p & v3a5f992;
assign v37463ae = hgrant2_p & v8455ba | !hgrant2_p & v3a70aa4;
assign v376a399 = hbusreq6_p & v372d630 | !hbusreq6_p & v3769e8c;
assign c858c6 = hbusreq0_p & v3a60bc8 | !hbusreq0_p & v8455b5;
assign v37523de = hgrant5_p & v3726d60 | !hgrant5_p & v3a700e6;
assign v377f85a = hmaster2_p & v8455ab | !hmaster2_p & v3a6ffc7;
assign v372fe3c = hbusreq5 & v377c0ad | !hbusreq5 & !v8455b9;
assign v37677e2 = hmaster1_p & v3a70236 | !hmaster1_p & v3a6f072;
assign v3a6f8a2 = hmaster3_p & v37474fc | !hmaster3_p & v375e7bb;
assign v37556ae = hmaster2_p & v376ace2 | !hmaster2_p & !v8455ab;
assign v3a63ef6 = hbusreq8 & v3a6f6d1 | !hbusreq8 & v3779c26;
assign v3751a0b = hbusreq1 & v374f307 | !hbusreq1 & v8455b0;
assign v375d5ac = hbusreq2_p & v3a6a895 | !hbusreq2_p & !v8455ab;
assign c8a454 = hbusreq4_p & v3a5d80f | !hbusreq4_p & v8455ab;
assign v37611c1 = hbusreq2_p & v3a6d621 | !hbusreq2_p & v3736319;
assign v3a7031a = hmaster2_p & v3a619c0 | !hmaster2_p & v8455ab;
assign v3769cd3 = hbusreq6_p & v3a58218 | !hbusreq6_p & v3a6f778;
assign v373861f = hmaster0_p & v374bfd2 | !hmaster0_p & v373fdae;
assign v3a6ff7c = hbusreq2_p & v3a6fda4 | !hbusreq2_p & v37749bf;
assign v374dfd5 = hmaster2_p & v373e52d | !hmaster2_p & v37606dc;
assign v375c196 = hbusreq1 & v3769cad | !hbusreq1 & v380662a;
assign v3725f4a = hbusreq2 & v3723430 | !hbusreq2 & v8455ab;
assign v372db12 = hbusreq7_p & v3a63c8e | !hbusreq7_p & v3761026;
assign v3a575d6 = hgrant2_p & v3750269 | !hgrant2_p & v375fbc0;
assign v37237e8 = hmaster2_p & v374c7f4 | !hmaster2_p & v3732569;
assign v3777f01 = hbusreq5 & v3a6f541 | !hbusreq5 & v37613bf;
assign v3a616ad = hgrant4_p & v3724fdb | !hgrant4_p & v374b8c5;
assign v3a60b56 = hbusreq5 & v374fde8 | !hbusreq5 & !v375aa0d;
assign v37773a9 = hlock0_p & v8455e7 | !hlock0_p & !v8455ab;
assign v3772c92 = hbusreq2_p & v376021f | !hbusreq2_p & v3a586d0;
assign v372952d = hbusreq4 & v3774acc | !hbusreq4 & v375aea6;
assign v373bb6c = hmaster2_p & v3a5f8a2 | !hmaster2_p & v3753258;
assign v3765396 = hbusreq0 & v3a5b39d | !hbusreq0 & v372ddfa;
assign v3a58bb0 = hgrant4_p & v376a6f1 | !hgrant4_p & v37706dd;
assign v373ca0e = hbusreq3_p & cb89d9 | !hbusreq3_p & v8455ab;
assign v376445f = hmaster2_p & v3a635ea | !hmaster2_p & v374acbe;
assign v375c06a = hbusreq6 & v3766f1c | !hbusreq6 & !v8455ab;
assign v377ce47 = hmaster2_p & v209312a | !hmaster2_p & v3a5971e;
assign v3a68931 = hgrant5_p & v3a5b01c | !hgrant5_p & v373d071;
assign v376f23f = hlock6 & v37649d3 | !hlock6 & v3a646fb;
assign v3a60859 = hmaster1_p & v2925d03 | !hmaster1_p & v3a713da;
assign v3a70da8 = hbusreq7_p & v37240c0 | !hbusreq7_p & v3a56918;
assign v3a70f03 = hgrant3_p & v8455be | !hgrant3_p & v375a901;
assign v884deb = hlock2 & aebd68 | !hlock2 & v373e296;
assign v37296db = hlock0_p & v3a5ad13 | !hlock0_p & v37737f9;
assign v3a67715 = hbusreq7 & v3a593b0 | !hbusreq7 & v3734279;
assign v375cd7b = hmaster1_p & v373ed5c | !hmaster1_p & v372f9b4;
assign v3a700e6 = hmaster1_p & v3a54aa0 | !hmaster1_p & v37229ba;
assign v3730d16 = hmaster0_p & v380952f | !hmaster0_p & !v372a520;
assign v3a70405 = hlock4 & v3772edc | !hlock4 & v372a94e;
assign v3a5a16b = hbusreq2 & v3a5617a | !hbusreq2 & v3748797;
assign v3a6e50e = hlock4 & v3a5d6c6 | !hlock4 & v3a70cb1;
assign v376a348 = hbusreq4 & v3a6dc08 | !hbusreq4 & v373f058;
assign v3a565a8 = hbusreq4_p & v3a55dc3 | !hbusreq4_p & v380919d;
assign v3a6fbaa = hmaster2_p & v3735324 | !hmaster2_p & v8455ab;
assign v3a626fe = hbusreq5 & v377b0d8 | !hbusreq5 & v3a5584b;
assign v3744ff3 = hbusreq0 & v3a6c6f6 | !hbusreq0 & v3767d14;
assign v3a6ebb0 = hbusreq2 & v37624a2 | !hbusreq2 & v3a7153a;
assign v372a7c9 = hgrant1_p & v8455b0 | !hgrant1_p & v8455ab;
assign v37728c2 = hgrant4_p & v8455ab | !hgrant4_p & v37442e1;
assign v3a61a1d = jx3_p & v3a70f3f | !jx3_p & !v8455ab;
assign v3a669c2 = hbusreq6_p & v3757aa1 | !hbusreq6_p & v377b576;
assign v37507dc = hmaster0_p & v3a712ca | !hmaster0_p & v3a5b071;
assign v3a6471e = hbusreq7_p & v3a57759 | !hbusreq7_p & !v374e590;
assign v3377c6c = hbusreq4_p & v380922b | !hbusreq4_p & v3a5b079;
assign v3a6f4ea = hbusreq7 & v3a62229 | !hbusreq7 & a0a219;
assign v377cbad = hbusreq2_p & v3a68c1f | !hbusreq2_p & !v3a66110;
assign v35b779f = hgrant2_p & v8455ab | !hgrant2_p & v3a6fb14;
assign v3a5d76d = hbusreq5_p & v375f159 | !hbusreq5_p & v3a6a693;
assign v377fc87 = hbusreq2_p & v375c379 | !hbusreq2_p & v376d817;
assign v3741a83 = hmaster2_p & v8455ab | !hmaster2_p & v3730ffe;
assign v3769628 = hlock2_p & v3775b81 | !hlock2_p & v8455ab;
assign v3a6e4cd = hmaster2_p & v3a613f4 | !hmaster2_p & v3a70d66;
assign v3761c72 = hmaster2_p & v3a6b60d | !hmaster2_p & v37745c3;
assign v37261ad = hbusreq5 & v3a65e55 | !hbusreq5 & v3a6eaf8;
assign v376d1bb = hbusreq0 & v3729fa0 | !hbusreq0 & v3a71166;
assign v37247f2 = hbusreq4 & v3753dab | !hbusreq4 & v8455ab;
assign v37488fe = hgrant6_p & v3a6f61e | !hgrant6_p & !v3770ab9;
assign v377871a = hbusreq4 & v3752f2e | !hbusreq4 & v8455ab;
assign v3734ba4 = hmaster1_p & v375e037 | !hmaster1_p & v3a6f4da;
assign v3a636c0 = hbusreq7_p & v377456d | !hbusreq7_p & v3768734;
assign v37495ed = hmaster2_p & v3a635ea | !hmaster2_p & v3a6eb7b;
assign v3750d4c = hgrant6_p & v3a6f3aa | !hgrant6_p & v372ea14;
assign v3744280 = hmaster0_p & v37705f3 | !hmaster0_p & v372f1d4;
assign v377fb09 = hbusreq4_p & v3a6fc9c | !hbusreq4_p & v8455b0;
assign v377c487 = hbusreq7 & v375439c | !hbusreq7 & v8455ab;
assign v3745186 = hmaster2_p & v37245f8 | !hmaster2_p & v3a70d99;
assign v3a7161c = hmaster0_p & v8455ab | !hmaster0_p & v37520fc;
assign v3730f21 = hbusreq5_p & v3a6e916 | !hbusreq5_p & !v8455ab;
assign v372b6d0 = hmaster2_p & v376a6f1 | !hmaster2_p & v372cacb;
assign v3a68016 = hgrant3_p & v8455ab | !hgrant3_p & v3a2a770;
assign v3a5fb37 = hbusreq6_p & v37558b4 | !hbusreq6_p & v3a6be6d;
assign v3a62eaa = hbusreq7_p & v3a6f622 | !hbusreq7_p & v3a714ed;
assign v9644fd = hgrant2_p & v372f09a | !hgrant2_p & v3a701e7;
assign v377aad8 = hbusreq1_p & v376b97b | !hbusreq1_p & v3754c0e;
assign v3755f9b = hbusreq0 & v372cdf6 | !hbusreq0 & v8455ab;
assign v3a682f9 = hbusreq5_p & v3761671 | !hbusreq5_p & !v3a6fb9b;
assign v3a62082 = hgrant6_p & v3a7083b | !hgrant6_p & v3a6f6b8;
assign v3a6bf89 = hgrant6_p & v8455ab | !hgrant6_p & v375d6ba;
assign v3775902 = hmaster0_p & v3a628d4 | !hmaster0_p & v373197c;
assign v3a5fd58 = hmaster0_p & v37370f0 | !hmaster0_p & v3a63f29;
assign v377bbd1 = hgrant0_p & v3a6faac | !hgrant0_p & v23fe03a;
assign v3a70c37 = hmaster1_p & v377e36c | !hmaster1_p & v373db68;
assign v3a6f860 = hbusreq8_p & v373afa4 | !hbusreq8_p & v3a71041;
assign v373cbf9 = hbusreq4_p & v3a7162d | !hbusreq4_p & v3778528;
assign v3770919 = hbusreq2_p & v3729ffd | !hbusreq2_p & v37797ef;
assign v3a70369 = hmaster2_p & v3a6a8ee | !hmaster2_p & v3a70ff5;
assign v3739ec6 = hmaster0_p & v2acb0a5 | !hmaster0_p & v375d2b3;
assign v377ba37 = hbusreq4 & v377d8d6 | !hbusreq4 & !v3a5aca8;
assign b27f78 = hbusreq1_p & v3770b89 | !hbusreq1_p & v1e38224;
assign v3774641 = hmaster1_p & v3743b12 | !hmaster1_p & v374b747;
assign v3a61eea = hbusreq6 & v3a5b7b5 | !hbusreq6 & v8455ab;
assign v374550d = hbusreq0 & v3a70906 | !hbusreq0 & v377c31d;
assign v3736011 = hmaster1_p & v376ec9b | !hmaster1_p & v376a40c;
assign v3a707ec = hmaster0_p & v375df8e | !hmaster0_p & v3a5e371;
assign v3a6ca24 = hbusreq2 & v3737d44 | !hbusreq2 & v8455ab;
assign v3a64709 = hmaster2_p & v3a635ea | !hmaster2_p & v3a70a7f;
assign v3a7089e = hgrant5_p & d5e2c2 | !hgrant5_p & v373ebd2;
assign v3733d6e = hlock0_p & v376ef42 | !hlock0_p & v37736a6;
assign v37573b9 = hgrant3_p & v35b7299 | !hgrant3_p & !v3738b0c;
assign v3a58f56 = hmaster2_p & v3a6fc7f | !hmaster2_p & v375f9e9;
assign v3769605 = hbusreq3 & v3a559f0 | !hbusreq3 & v3733c39;
assign v373d4e8 = hgrant1_p & v3a7151d | !hgrant1_p & v8455ab;
assign v374d95f = hmaster1_p & v3a5a807 | !hmaster1_p & v37621d5;
assign v373b733 = hbusreq7 & v37668b8 | !hbusreq7 & v3737808;
assign v3a6f569 = hgrant5_p & v3a70578 | !hgrant5_p & v373fb1a;
assign v37523f8 = hmaster1_p & v3a635ea | !hmaster1_p & v3a5f4c6;
assign v3a672b6 = hlock8 & v38079db | !hlock8 & v375c3c5;
assign v3a57e21 = hgrant1_p & v3a619c0 | !hgrant1_p & v3744a2f;
assign v372ffd2 = hbusreq3_p & v3a6efdd | !hbusreq3_p & v3740655;
assign v3745458 = hmaster0_p & v3a6380f | !hmaster0_p & !v374b68a;
assign v376beaa = hbusreq0 & v372339a | !hbusreq0 & v3a6f447;
assign v374f29f = hbusreq3_p & v374fbca | !hbusreq3_p & !v8455ab;
assign v3a5d6f3 = hlock7 & v37679f0 | !hlock7 & v37402b8;
assign v3a6f3aa = hbusreq6_p & v3764ac0 | !hbusreq6_p & v374c0c9;
assign v3a70570 = hmaster1_p & v8455c6 | !hmaster1_p & v373700d;
assign v3a615a2 = hgrant3_p & v373b4ce | !hgrant3_p & v2aca977;
assign v3760881 = hbusreq0 & v3a5f4b1 | !hbusreq0 & v3a702cb;
assign v3a701b7 = hbusreq5 & v373eadd | !hbusreq5 & v8455ab;
assign v3a6b90e = hbusreq5_p & v374e968 | !hbusreq5_p & v3769b7e;
assign v3747ef9 = hlock5 & v3a6ae23 | !hlock5 & v373fa48;
assign v37549e1 = hbusreq3 & v3725230 | !hbusreq3 & v8455ab;
assign v3779d6b = hmaster1_p & v3a63556 | !hmaster1_p & v3a6f3f2;
assign v372dab0 = hgrant2_p & v3a70c0b | !hgrant2_p & !v209310e;
assign v3772b14 = hmaster2_p & v3759b2f | !hmaster2_p & v376ea4a;
assign v3a6c467 = hbusreq3 & v3a5600a | !hbusreq3 & v3773b23;
assign v38094fb = hlock6_p & v373c755 | !hlock6_p & v8455ab;
assign v3a70aae = hmaster2_p & v3a661fe | !hmaster2_p & v3a702c2;
assign v37474da = hgrant6_p & v3a5cb5f | !hgrant6_p & v375c463;
assign v2ff8f77 = hmaster1_p & v8455b0 | !hmaster1_p & v3a6f87e;
assign v3a6fd8f = hbusreq4 & v3748de3 | !hbusreq4 & v377b67d;
assign v3726381 = hlock0 & v3757009 | !hlock0 & v3a6f8fd;
assign v374a0ab = hmaster1_p & v3763571 | !hmaster1_p & v3747271;
assign v3752ebb = hbusreq5_p & v3777da6 | !hbusreq5_p & v3731b41;
assign v376156f = hbusreq5 & v377282c | !hbusreq5 & v3a5e859;
assign v374fef7 = hbusreq2 & v3a5f0cf | !hbusreq2 & v8455ab;
assign v3737bc8 = hgrant2_p & v375c55a | !hgrant2_p & v3768eb1;
assign v3a5b9c3 = hbusreq8 & v3a714e0 | !hbusreq8 & v3a6dcbf;
assign v3a6f827 = hmaster3_p & v3a29835 | !hmaster3_p & v3a5bd12;
assign v3a62d1c = hbusreq5 & v37360c8 | !hbusreq5 & v38076cf;
assign v3a6f9b6 = hmaster1_p & v3751e0a | !hmaster1_p & v3734c3a;
assign v3770b33 = hmaster1_p & v3764530 | !hmaster1_p & !v37420de;
assign v377855f = hbusreq4_p & v3759fca | !hbusreq4_p & v3a637dd;
assign v372bd5f = hmaster2_p & v377e089 | !hmaster2_p & !v3729421;
assign v8455eb = hgrant1_p & v8455ab | !hgrant1_p & !v8455ab;
assign v3764d1f = hbusreq2 & v377094b | !hbusreq2 & v8455ab;
assign v3a6fb9e = hbusreq7 & v97b684 | !hbusreq7 & v3a70265;
assign v3a64994 = hlock1 & v3a70378 | !hlock1 & v372ab85;
assign v3773a25 = hmaster2_p & v3a58218 | !hmaster2_p & v3753dab;
assign v3742eaf = hbusreq6 & v372422d | !hbusreq6 & v3762223;
assign v377e5fd = hgrant0_p & v875999 | !hgrant0_p & v23fe285;
assign v3a70432 = hgrant6_p & v921bc8 | !hgrant6_p & v8455ab;
assign v375439c = hmaster1_p & v37356f0 | !hmaster1_p & v39a53eb;
assign v3a70400 = jx2_p & v3a56e15 | !jx2_p & v3769524;
assign v3732208 = hmaster2_p & v3753c73 | !hmaster2_p & v373f24b;
assign v3a68240 = hbusreq2_p & v3a6eeca | !hbusreq2_p & v2092bae;
assign c99197 = hlock0_p & v3740d36 | !hlock0_p & v3a5e24e;
assign v37474fc = jx0_p & v3755b55 | !jx0_p & v37301f9;
assign v37c025b = hmaster1_p & v3a29814 | !hmaster1_p & v37560b0;
assign v3746f58 = hgrant5_p & v373c1a2 | !hgrant5_p & v3a6602d;
assign v37397ba = hbusreq5 & v3738e3c | !hbusreq5 & v3a6eece;
assign v376f8ea = hbusreq5_p & v3749bc0 | !hbusreq5_p & !v3757cd1;
assign v360cdfe = hbusreq3_p & v3755806 | !hbusreq3_p & v8455ab;
assign v373c56f = hgrant5_p & v3a5a807 | !hgrant5_p & v3a7072d;
assign v3a6d198 = jx1_p & v373fc52 | !jx1_p & adaeff;
assign v375c7cf = hmaster0_p & v375fe58 | !hmaster0_p & v373a822;
assign v37383d3 = hbusreq5_p & v3a584fd | !hbusreq5_p & v3a70736;
assign v3a712a6 = hbusreq8_p & v374ba3c | !hbusreq8_p & v8455ab;
assign v377d4de = hmaster2_p & v3777844 | !hmaster2_p & v3a5eaaf;
assign v3a6eec2 = hgrant2_p & v8455ab | !hgrant2_p & v376eeac;
assign v3809964 = hlock5 & v3733294 | !hlock5 & v3a70dcb;
assign v3a5b7b5 = hgrant2_p & v3723430 | !hgrant2_p & v374bf71;
assign v3a71061 = hgrant3_p & v3a615f7 | !hgrant3_p & v377c185;
assign v376ef20 = hgrant5_p & v373ad69 | !hgrant5_p & v3a5c349;
assign v3777a6c = hlock6_p & v3a54c77 | !hlock6_p & !v8455ab;
assign v3778281 = hbusreq0 & v37282f3 | !hbusreq0 & v374a7ab;
assign v3766014 = hmaster0_p & v8455ab | !hmaster0_p & v3a7128e;
assign v3767415 = hmaster1_p & v3a70b77 | !hmaster1_p & v374b747;
assign v37330d3 = hbusreq5_p & v3727f68 | !hbusreq5_p & !v3a6333a;
assign v373acc2 = hgrant6_p & v3a69146 | !hgrant6_p & v3743285;
assign v3a7017f = hmaster3_p & v3a712b5 | !hmaster3_p & v3766f30;
assign v374247d = hbusreq8_p & v3a6e40f | !hbusreq8_p & v3a6f411;
assign v3a710ba = hbusreq6 & v3737d44 | !hbusreq6 & !v8455ab;
assign v3779470 = hbusreq5 & v3a6fe0d | !hbusreq5 & !v8455b5;
assign v37763d1 = hgrant4_p & v8455e7 | !hgrant4_p & !v8455ab;
assign v375aacf = hbusreq5 & v3a6fdee | !hbusreq5 & v374949f;
assign v376a39c = hgrant6_p & v372ffaa | !hgrant6_p & v374fe73;
assign v3a6efaa = hbusreq1_p & v376b0e6 | !hbusreq1_p & !v8455ab;
assign v3a70cd9 = hgrant2_p & v8455ab | !hgrant2_p & v375ea72;
assign v3752ac9 = hgrant6_p & v8455c9 | !hgrant6_p & v3729620;
assign v377defb = hgrant6_p & v3743ded | !hgrant6_p & v3a6f91a;
assign v3744b3d = hmaster0_p & v3760799 | !hmaster0_p & v374974e;
assign v3a6650e = hbusreq6 & v3767ea6 | !hbusreq6 & !v8455ab;
assign v3775508 = hlock5 & v3a6f28a | !hlock5 & v3a6934e;
assign v3755ae2 = hbusreq7 & v375e9ca | !hbusreq7 & v3a6f1d8;
assign v377dc8f = hbusreq7 & v3757afc | !hbusreq7 & v3a71551;
assign v3770ecc = hbusreq5_p & v8455bb | !hbusreq5_p & v3760513;
assign v3741ae7 = hgrant6_p & v3724475 | !hgrant6_p & v377149d;
assign v3770be6 = hbusreq7_p & v37343bd | !hbusreq7_p & v3760066;
assign v3a6f6c8 = hbusreq7_p & v3a70655 | !hbusreq7_p & v3749520;
assign v3743d8b = hgrant6_p & v8455ab | !hgrant6_p & v3a5688f;
assign v374cbc0 = hgrant4_p & v8455ab | !hgrant4_p & v3a59eb3;
assign v3806579 = hmaster1_p & v3a6f7dd | !hmaster1_p & v3a58dfc;
assign v3772ac1 = hbusreq7 & v3a648c8 | !hbusreq7 & v3766472;
assign v374a430 = hlock2 & v37551e3 | !hlock2 & v3378a34;
assign v376b7a8 = jx0_p & v374ea7e | !jx0_p & v374717a;
assign v3770f6e = hgrant2_p & v9ed516 | !hgrant2_p & v374dfea;
assign v3a6fb45 = hgrant2_p & v372b163 | !hgrant2_p & !v8455ab;
assign v1e37413 = hbusreq6_p & v3a5ee6e | !hbusreq6_p & v3770735;
assign v376dee4 = hmaster3_p & v8455ab | !hmaster3_p & v2092bfc;
assign v37445ff = hmaster2_p & v372be16 | !hmaster2_p & v3a706a4;
assign v3753298 = hmaster2_p & v37297cb | !hmaster2_p & v3a5b7db;
assign v3732e48 = hmaster1_p & v372ba1c | !hmaster1_p & v3a61038;
assign v3755e35 = hbusreq2 & v3a5689e | !hbusreq2 & v375c1d1;
assign v3743adf = hlock0 & v3a7162d | !hlock0 & v374021a;
assign v374a3b8 = hlock0 & v38072fd | !hlock0 & v3728f3a;
assign v37293f6 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3a5b47c;
assign v372317f = hbusreq5_p & v374c6b8 | !hbusreq5_p & v375ede6;
assign v3753e28 = hbusreq7_p & v3779b12 | !hbusreq7_p & v3728e91;
assign v37611a9 = hbusreq4 & v377d9bb | !hbusreq4 & v37434ce;
assign v3737e97 = hgrant5_p & v373d10a | !hgrant5_p & v376eb57;
assign v372615f = hgrant4_p & v3768c78 | !hgrant4_p & v3a70393;
assign v3a6e927 = hmaster1_p & v3a70f0c | !hmaster1_p & v3726da1;
assign v3a70219 = hbusreq3 & v3a5eac0 | !hbusreq3 & v8455ab;
assign v3738eb0 = hbusreq5_p & v3a5f449 | !hbusreq5_p & !v3a571d1;
assign v3a6261c = hmaster1_p & v372f2fe | !hmaster1_p & v3a6ed27;
assign v375833e = hlock3_p & v3a6f668 | !hlock3_p & v8455ab;
assign v3756aea = hbusreq0 & v3a6becb | !hbusreq0 & v3770d93;
assign v3749a17 = hmaster0_p & v3736610 | !hmaster0_p & v3749846;
assign v3a6ea66 = hgrant4_p & v3a7137c | !hgrant4_p & v3a712af;
assign v3740dcc = hbusreq7 & v3740489 | !hbusreq7 & !v8455bd;
assign v373db8f = hlock6_p & v3742122 | !hlock6_p & v375d616;
assign v377a801 = hgrant4_p & v8455ab | !hgrant4_p & v3a5d830;
assign v3742905 = hlock2 & v374172f | !hlock2 & v373502a;
assign v37678eb = hmaster0_p & v3a70124 | !hmaster0_p & v377402f;
assign v3774f07 = hmaster1_p & v3a5373e | !hmaster1_p & v372af40;
assign b62443 = hmaster2_p & v37793a4 | !hmaster2_p & v377bb6d;
assign v3a68523 = hgrant0_p & v8455ab | !hgrant0_p & v3a5ae6d;
assign v3a709d0 = hgrant2_p & v376e04c | !hgrant2_p & v3a5574a;
assign v3741e12 = hready & v3a54d59 | !hready & v8455ab;
assign v3a661fe = hlock6_p & v3755002 | !hlock6_p & !v8455ab;
assign v3a70154 = hmaster0_p & v39a4d8a | !hmaster0_p & v3761c61;
assign v3739983 = hmaster3_p & v374139a | !hmaster3_p & v3a6d8f4;
assign v3a5e8f6 = stateG10_1_p & v8455e7 | !stateG10_1_p & !v3a70056;
assign v3a70106 = hbusreq5_p & v3a5b7ad | !hbusreq5_p & v3a5ba93;
assign v23fde9c = hbusreq7 & v3a70c67 | !hbusreq7 & v373b837;
assign v377d7a4 = hbusreq6_p & v37757e0 | !hbusreq6_p & v3773b23;
assign v3746a78 = stateG10_1_p & v8455ab | !stateG10_1_p & !v3723430;
assign v376a4ba = hmaster0_p & v37519cb | !hmaster0_p & !v3731bb5;
assign v373013d = hbusreq5 & v3752115 | !hbusreq5 & v37567f5;
assign v373cf96 = hbusreq0 & v3a6fadb | !hbusreq0 & v3726c8d;
assign v3737c86 = hbusreq6 & v3a705f4 | !hbusreq6 & v8455ab;
assign v375ad7d = hlock8_p & v374cd37 | !hlock8_p & v8455ab;
assign v2619b04 = hgrant4_p & v3a53eeb | !hgrant4_p & v373b8e2;
assign v3a6ebe7 = hbusreq1 & v3737554 | !hbusreq1 & v8455ab;
assign v3a69adb = hgrant0_p & v3779060 | !hgrant0_p & v3a70ab7;
assign v3725410 = hbusreq1_p & v3a71014 | !hbusreq1_p & v8455ab;
assign v376600a = hbusreq5 & v376265d | !hbusreq5 & v373fcbf;
assign v8455d5 = hburst0_p & v8455ab | !hburst0_p & !v8455ab;
assign v3746696 = hlock6 & v38072fd | !hlock6 & v3a6fa76;
assign v37506fb = hbusreq3_p & v376d5a4 | !hbusreq3_p & v35772a6;
assign v374b3e1 = hbusreq0_p & a38ed7 | !hbusreq0_p & v37775c4;
assign v374ae4a = hgrant6_p & v377edba | !hgrant6_p & !v3a5d373;
assign v3764257 = hgrant5_p & v8455ab | !hgrant5_p & !v3765222;
assign v3a57118 = hgrant4_p & v3a602c3 | !hgrant4_p & v3772a3f;
assign v3a62250 = hmaster0_p & v3a635ea | !hmaster0_p & v3a70e7d;
assign v3727345 = busreq_p & v8455ab | !busreq_p & v373cdb4;
assign v3a62508 = hbusreq4_p & v37558eb | !hbusreq4_p & v3759d3c;
assign v374cab9 = locked_p & v3a70a29 | !locked_p & v39a5381;
assign v3a6c6c3 = jx0_p & v3a66b6e | !jx0_p & v3a71342;
assign v374a65c = hmaster2_p & v374571d | !hmaster2_p & v376d374;
assign v3774a7e = hgrant2_p & v3751931 | !hgrant2_p & v375f4fd;
assign v3a6c905 = hbusreq5 & v3a66c9a | !hbusreq5 & v3a6ff12;
assign v377ebc9 = jx0_p & v3a29856 | !jx0_p & v3756471;
assign v37452d5 = hgrant3_p & v8455ab | !hgrant3_p & v3a5ef37;
assign v3a62f70 = hbusreq5_p & v3778c64 | !hbusreq5_p & v3771994;
assign v3740d4a = hmaster2_p & v375b7b0 | !hmaster2_p & v3a70b80;
assign v3a5bfbd = hmaster1_p & v37438ba | !hmaster1_p & v3764daf;
assign v37733c0 = hbusreq4_p & v3731549 | !hbusreq4_p & v377d256;
assign v3728040 = hbusreq5_p & v376c2d6 | !hbusreq5_p & v1e37dcd;
assign v37334ff = hbusreq7_p & v376c17d | !hbusreq7_p & v3733b84;
assign v3a6f8f5 = hlock3_p & v3765e46 | !hlock3_p & !v8455ab;
assign v3a69761 = hlock7 & v375f6e3 | !hlock7 & v3a69961;
assign v3753fc9 = hmaster1_p & v377ef09 | !hmaster1_p & v375e30f;
assign v37718d5 = hbusreq8_p & c5b5f4 | !hbusreq8_p & v3a6fd90;
assign v3a684af = hgrant0_p & v374fb58 | !hgrant0_p & v3a6f656;
assign v3737edc = hmaster3_p & v3a5ed64 | !hmaster3_p & v3a6a635;
assign v3a53f2b = hbusreq6 & v375f98a | !hbusreq6 & v8455ab;
assign v3a6ec6d = hlock2 & v3750547 | !hlock2 & v37415b2;
assign v374949d = hmaster0_p & v375d7df | !hmaster0_p & !v374b1a4;
assign v397d85e = hgrant6_p & v377f09a | !hgrant6_p & v3a70c54;
assign v3a5bfe6 = hbusreq4_p & v377f46d | !hbusreq4_p & v3776f8c;
assign v3a7059e = hmaster1_p & v3a62cac | !hmaster1_p & v3a6f601;
assign v37684c0 = hbusreq8_p & v376ae9f | !hbusreq8_p & v3a5f586;
assign v373abe2 = hbusreq2 & v376430b | !hbusreq2 & v376653d;
assign v8d428b = hbusreq2_p & v3777749 | !hbusreq2_p & v3a6fe5d;
assign v3726979 = hlock0 & v3a70a88 | !hlock0 & v3a6d03c;
assign v37488ed = hbusreq3 & v375ed5a | !hbusreq3 & v376a6d7;
assign v374b30b = hbusreq4 & v3a6dc08 | !hbusreq4 & v375d616;
assign v3730f35 = hbusreq4 & v23fe101 | !hbusreq4 & v3a635ea;
assign v37380d5 = hbusreq7_p & v377c56c | !hbusreq7_p & v37652d7;
assign v373e845 = hbusreq5 & v3762eeb | !hbusreq5 & v3777c0c;
assign v377d320 = locked_p & v374f0c1 | !locked_p & v3577306;
assign v375562a = hbusreq4_p & v3a6f42e | !hbusreq4_p & !v3755252;
assign v3a68004 = hbusreq4 & v372c3d4 | !hbusreq4 & v3760f87;
assign v37360c1 = jx0_p & v3731211 | !jx0_p & v3a61ceb;
assign v3725bdc = hready & v3a703dd | !hready & v8455ab;
assign v3767f58 = hbusreq6_p & v8d9a96 | !hbusreq6_p & !v8455ab;
assign v3757d5b = hbusreq5 & v3a5b4bd | !hbusreq5 & v373a693;
assign v3729b37 = hgrant3_p & v8455be | !hgrant3_p & !v376db8a;
assign v3769753 = hlock5 & v3727bc1 | !hlock5 & v3a70572;
assign v377312b = hmaster1_p & v3a702c5 | !hmaster1_p & v372ee5a;
assign v3a6ca4e = hbusreq6_p & v373e933 | !hbusreq6_p & v3756b48;
assign v374c9c7 = busreq_p & v377adc8 | !busreq_p & !v3a6fc6e;
assign v377f829 = hmaster1_p & v3a70f8b | !hmaster1_p & v3738826;
assign v3a6fce1 = hbusreq4 & v3a5b037 | !hbusreq4 & v8455ab;
assign v372bee9 = hbusreq7_p & v9ac541 | !hbusreq7_p & !v39a4dc7;
assign v374c9e1 = hmaster3_p & v3733cf4 | !hmaster3_p & af0958;
assign v3a6368a = stateG10_1_p & v3809adf | !stateG10_1_p & !v3a5c5ae;
assign v3a70a23 = hlock6_p & v37624a2 | !hlock6_p & v8455b0;
assign v2092ef2 = hmaster2_p & v37315e2 | !hmaster2_p & v377d1dc;
assign v3a71604 = hbusreq5 & v3778bb4 | !hbusreq5 & v8455ab;
assign v3729880 = hbusreq0_p & v375e60f | !hbusreq0_p & !v3a672c9;
assign v3766afa = hmaster1_p & v8455ab | !hmaster1_p & v3775a8e;
assign v373a1d0 = hbusreq5_p & v377984a | !hbusreq5_p & aa9893;
assign v3742a57 = hmaster0_p & v374dd8f | !hmaster0_p & v376189d;
assign v374ad7d = hbusreq0 & v377bb3a | !hbusreq0 & v3a61f4c;
assign v372fba5 = hready & v3a690ec | !hready & !v3a5f308;
assign v3766b5a = hbusreq5 & v3727981 | !hbusreq5 & v3a6542a;
assign v3753bac = hbusreq6_p & v380a2f5 | !hbusreq6_p & v3725a56;
assign v3a5b359 = hlock6_p & v373e209 | !hlock6_p & v377af44;
assign jx3 = !v39af33c;
assign v3378a03 = hlock2 & v360c6b6 | !hlock2 & v3a55ba9;
assign v3768b07 = hbusreq2_p & v3a6f5f6 | !hbusreq2_p & v375dcdb;
assign v3806b0a = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3a7162d;
assign v3a6d531 = hmaster2_p & v37666f6 | !hmaster2_p & v8455ab;
assign v3772827 = hbusreq4 & v3a5952d | !hbusreq4 & v3a707c4;
assign v372ce88 = hbusreq6 & v3a7096e | !hbusreq6 & v376ef7a;
assign v2619aa5 = hmaster2_p & v3a5fe9e | !hmaster2_p & v3775688;
assign v8455f9 = hgrant8_p & v8455ab | !hgrant8_p & !v8455ab;
assign v375e944 = hmaster2_p & v3a6f23a | !hmaster2_p & v374e0f6;
assign v377021d = hgrant6_p & v37369b2 | !hgrant6_p & v3a70cd9;
assign v372647c = hgrant5_p & v3740f78 | !hgrant5_p & v3a62e77;
assign v37315af = hmaster0_p & v3a712c2 | !hmaster0_p & v376b1a1;
assign v377d7dc = hlock4_p & v3a6a939 | !hlock4_p & !v8455ab;
assign v372e88a = hgrant3_p & v8455e7 | !hgrant3_p & !v3768933;
assign v3a6f11b = hbusreq5 & v377e089 | !hbusreq5 & !v8455bd;
assign v374bfcf = hgrant4_p & v376a6f1 | !hgrant4_p & c35240;
assign v372e03f = hlock6_p & v374b8ad | !hlock6_p & v3a5be6a;
assign v376f56d = hready & v3749a12 | !hready & v8455ab;
assign v3779863 = hlock8 & v374a0f0 | !hlock8 & v3765224;
assign v3754c99 = hmaster1_p & v37383da | !hmaster1_p & v3724ced;
assign v3737dee = hlock5_p & v37640e2 | !hlock5_p & v3739646;
assign v37785f8 = hbusreq5 & v3a65e55 | !hbusreq5 & v374d255;
assign v97e702 = hmaster1_p & v3723923 | !hmaster1_p & v3729830;
assign v376b5bc = hbusreq2_p & v3759fe8 | !hbusreq2_p & v8455ab;
assign v3a70a44 = hbusreq8_p & v3723c25 | !hbusreq8_p & v3a299ba;
assign v374fcf6 = hbusreq2_p & v37316b7 | !hbusreq2_p & v374fa56;
assign v3753bb4 = hmaster0_p & v3a5fc34 | !hmaster0_p & v8e06bc;
assign v3757e32 = hlock8 & v375ad79 | !hlock8 & v3a60f1a;
assign v3730289 = hbusreq7_p & v373d64d | !hbusreq7_p & !v377dc8f;
assign v37443e0 = hmaster2_p & v8455ab | !hmaster2_p & !v3a6f48b;
assign v3768c76 = hmaster1_p & v377a18b | !hmaster1_p & v374e7fa;
assign v377844d = hlock3 & v3736cc7 | !hlock3 & v3776b61;
assign v1e3737d = hmaster0_p & v8455ab | !hmaster0_p & v3776ada;
assign v377e142 = hlock0_p & v372ac5c | !hlock0_p & v3a6f2a2;
assign v37325ad = hgrant3_p & v8455ab | !hgrant3_p & !v3a703a4;
assign v3a5ae95 = hmaster2_p & v375166c | !hmaster2_p & v375d059;
assign v3a704b7 = hmaster3_p & v3738aef | !hmaster3_p & v3728085;
assign v376b83d = hlock6_p & v377169f | !hlock6_p & v3a65da7;
assign v35b7768 = hmaster3_p & v3a649da | !hmaster3_p & !v3746f18;
assign v37773a0 = hbusreq4_p & v3758636 | !hbusreq4_p & v3a667a7;
assign v37712f6 = hbusreq3_p & v3a70272 | !hbusreq3_p & !v3a5b68a;
assign v376c08d = hlock7_p & v374e855 | !hlock7_p & v8455cb;
assign v3809240 = hbusreq4 & v8455b0 | !hbusreq4 & v3a702c2;
assign v3a5998b = hmaster2_p & v9f823e | !hmaster2_p & v3a5b978;
assign v3a704d6 = hbusreq5_p & v3a63628 | !hbusreq5_p & v3a63e9b;
assign v3722ae9 = hmaster2_p & v37419bc | !hmaster2_p & v372a9c7;
assign v374cffd = hlock7 & v3753e3b | !hlock7 & v37798bb;
assign v3777a66 = hlock6 & v3a55aa8 | !hlock6 & v3a60ba3;
assign v373f03e = hbusreq6_p & v377eaf2 | !hbusreq6_p & v3762b55;
assign v3a6ed55 = hmaster1_p & v3738e62 | !hmaster1_p & !v3a2abf4;
assign v376070d = hbusreq6_p & v3778962 | !hbusreq6_p & v374500f;
assign v3a61279 = hbusreq2_p & cd348d | !hbusreq2_p & !v8455ab;
assign v373395b = hmaster0_p & v3733940 | !hmaster0_p & v373fc36;
assign v3746746 = hmaster1_p & v3a57b57 | !hmaster1_p & v37558f2;
assign v3a588ef = hgrant6_p & v1e37cd6 | !hgrant6_p & v37411df;
assign v3735f0b = hbusreq6 & v3773d82 | !hbusreq6 & b6390c;
assign v3a6a1f4 = hgrant3_p & v3a59ffa | !hgrant3_p & v3741dce;
assign v376046c = hbusreq5_p & v3a7077a | !hbusreq5_p & !v3749fd0;
assign v374215e = hbusreq8 & v3744cf1 | !hbusreq8 & v8455ab;
assign v37317f2 = hmaster2_p & v3a5bf5f | !hmaster2_p & v3a5fe9e;
assign v3a53cc2 = hbusreq8_p & v3755f80 | !hbusreq8_p & v3779863;
assign v372514f = hlock2 & v372a960 | !hlock2 & v377b4f2;
assign v3770359 = hgrant8_p & v8455ab | !hgrant8_p & v3a702dd;
assign v3a5d28b = hlock2_p & v3a703ac | !hlock2_p & !v8455ab;
assign v3739460 = hbusreq6_p & v3a5b91d | !hbusreq6_p & v3a632e8;
assign v375c0e8 = hlock5 & v3740bee | !hlock5 & v377e9a5;
assign v3728bff = hbusreq7_p & v3a655d2 | !hbusreq7_p & v37271ad;
assign v374378e = hbusreq4_p & v3a6f6bd | !hbusreq4_p & v3725b75;
assign v3a6c088 = hburst1 & v376c211 | !hburst1 & v376d387;
assign v3758561 = hmaster0_p & v3758524 | !hmaster0_p & v375d2b3;
assign v37638ee = hlock2 & v37711e1 | !hlock2 & v37699f2;
assign v3750c12 = hlock4 & v3748797 | !hlock4 & v3736b57;
assign v372ff3a = hlock6 & v3a6ffab | !hlock6 & v37523e9;
assign v3777b5f = hbusreq5 & v375b96f | !hbusreq5 & v377de7f;
assign v372fe1b = hbusreq6 & v3a5a8c3 | !hbusreq6 & v3766e4a;
assign v3761671 = hlock5_p & v3a5a1e8 | !hlock5_p & !v373c379;
assign v374f559 = hbusreq4 & v37796c6 | !hbusreq4 & v8455ab;
assign v372791c = hmaster1_p & v3a7152b | !hmaster1_p & v372794f;
assign v376dc58 = hbusreq3_p & v374f609 | !hbusreq3_p & v3a71644;
assign v3728e89 = hmaster2_p & v3a5b289 | !hmaster2_p & v8455bb;
assign v3a70dea = hgrant6_p & v8455ab | !hgrant6_p & v375c0cd;
assign v3743e7b = hmaster0_p & v8455bb | !hmaster0_p & v377ed5e;
assign v3a66274 = hbusreq7 & v377b3a2 | !hbusreq7 & v3730c0b;
assign v3745498 = hgrant5_p & v375f0f0 | !hgrant5_p & v3768690;
assign v3a55aa8 = hbusreq6 & v3a60ba3 | !hbusreq6 & v3766e4a;
assign v3a6eb65 = hmaster2_p & v374502e | !hmaster2_p & !v37583be;
assign v3739e39 = hlock2 & v2acaffd | !hlock2 & v374b310;
assign v3725506 = hlock2 & v375ddb7 | !hlock2 & v3731ffc;
assign v374b37d = hlock4 & v3a713ec | !hlock4 & v3a70dbe;
assign v3755cc3 = hmaster1_p & v8455ab | !hmaster1_p & v375a412;
assign v3a6f8ef = hmaster1_p & v8455ab | !hmaster1_p & v3746efa;
assign v3768c16 = hbusreq6_p & v3726229 | !hbusreq6_p & v37798ad;
assign v376fbb5 = hmaster0_p & v37288bc | !hmaster0_p & v3a6e318;
assign v374f95d = hbusreq4_p & v37578f3 | !hbusreq4_p & v3763cfa;
assign v373cdd5 = hlock0 & v376bade | !hlock0 & v375c3eb;
assign v376187f = hbusreq2_p & v376ba53 | !hbusreq2_p & v8455ab;
assign v3a71484 = hbusreq0 & v372d772 | !hbusreq0 & v3379037;
assign cc9d04 = hlock1_p & v3a5b5d3 | !hlock1_p & v3a658bf;
assign v3a68f16 = hbusreq4 & v3a6f586 | !hbusreq4 & !v3a6f3cf;
assign v3a6fe46 = hbusreq1_p & v3737d55 | !hbusreq1_p & !v8455ab;
assign v3a6fb07 = jx0_p & v37378a3 | !jx0_p & v374247d;
assign v3a70943 = hmaster0_p & v3807aa1 | !hmaster0_p & v372b686;
assign v372f6ec = hmaster1_p & be54b2 | !hmaster1_p & v372bc0c;
assign v3729620 = hbusreq6_p & v37439b2 | !hbusreq6_p & v3a6f7a0;
assign v377ef09 = hgrant4_p & v3a53eeb | !hgrant4_p & v373ca53;
assign v374a297 = hlock4 & v3a7168b | !hlock4 & v3577354;
assign v3a6a6eb = hbusreq0 & v373b548 | !hbusreq0 & !v8455ab;
assign v3a5e96b = hbusreq0 & v3a59e74 | !hbusreq0 & v3a6000d;
assign v3765e79 = hbusreq2_p & v3a635ea | !hbusreq2_p & v373b288;
assign v3727084 = hbusreq6_p & v8455bb | !hbusreq6_p & v37443ab;
assign v377ef58 = hbusreq5 & v3771be6 | !hbusreq5 & v8455b3;
assign v375409b = hbusreq4_p & v3a56b19 | !hbusreq4_p & v3756f42;
assign v3742efb = hmaster2_p & v8455ab | !hmaster2_p & v380881d;
assign v3a703d0 = hgrant2_p & v3a70f74 | !hgrant2_p & v372afd2;
assign v373720a = hlock1_p & v3762414 | !hlock1_p & v8455b0;
assign v37535e7 = hbusreq6 & v37bfd10 | !hbusreq6 & v8455ab;
assign v3730d6a = hgrant6_p & v1e37cd6 | !hgrant6_p & v375a83f;
assign v377703d = hmaster0_p & v3735ac3 | !hmaster0_p & v8455e7;
assign v374d40b = hbusreq2 & v23fdf85 | !hbusreq2 & v37730bf;
assign v377b576 = hbusreq1_p & v3a70fbb | !hbusreq1_p & !v8455ab;
assign v3a6fcad = hgrant4_p & v374195f | !hgrant4_p & v3771fd8;
assign v3752f15 = hmaster1_p & v8455ab | !hmaster1_p & v37302fa;
assign v3808db6 = hmaster0_p & v3769090 | !hmaster0_p & v374974e;
assign v37797c2 = hmaster0_p & v374b160 | !hmaster0_p & b05db7;
assign v3754f72 = hbusreq8 & v3a70461 | !hbusreq8 & v3a62bc6;
assign v374a48c = hlock2 & v3a70752 | !hlock2 & v3747527;
assign v3a713c7 = hbusreq2 & v3a6f8f5 | !hbusreq2 & v8455bf;
assign v3a5dd70 = hmaster1_p & v3751d9c | !hmaster1_p & v37519bf;
assign v3a702ed = hbusreq0_p & v374e0ba | !hbusreq0_p & v3a6ea51;
assign v374fc57 = hlock4 & v3764a07 | !hlock4 & v376e5fe;
assign v3779d24 = hgrant5_p & v8455c6 | !hgrant5_p & v3a68ebe;
assign v376b89f = hmaster1_p & v3a6a8c0 | !hmaster1_p & v3a69a9f;
assign v374c0c9 = hbusreq6 & v3a6fb2b | !hbusreq6 & v8455bf;
assign v3809093 = hbusreq1_p & v3a64994 | !hbusreq1_p & v373b288;
assign v375589b = hbusreq0_p & v37682c6 | !hbusreq0_p & v8455b6;
assign v3a7026c = hmaster2_p & v3a70374 | !hmaster2_p & v3727472;
assign v3725e9a = hlock7 & v374e650 | !hlock7 & v3a70301;
assign v3a7015b = hgrant5_p & v3a70a1f | !hgrant5_p & v372981a;
assign v377ceea = hbusreq0 & v375b8b9 | !hbusreq0 & v8455ab;
assign v3a68757 = hbusreq8_p & v3a70578 | !hbusreq8_p & v377d4dd;
assign v3a5e46d = hbusreq4_p & d7f8bb | !hbusreq4_p & v373bf79;
assign v3a5fdd3 = hbusreq2_p & v3a707cd | !hbusreq2_p & v37432c6;
assign v3775293 = hbusreq6_p & v3a635ea | !hbusreq6_p & v373c219;
assign v37330b1 = hmaster2_p & v2ff8cfd | !hmaster2_p & v3a6d175;
assign v3a60b0f = hmaster1_p & v37784b3 | !hmaster1_p & v3750113;
assign v377c5f8 = hbusreq5_p & v1e37d35 | !hbusreq5_p & v3a6f8a8;
assign v374657b = hmaster0_p & v3768953 | !hmaster0_p & !v3a70d93;
assign v3770733 = hlock5 & v3a6fb43 | !hlock5 & v3773078;
assign v3a68cb5 = hbusreq5_p & v373dd3c | !hbusreq5_p & v375345f;
assign v373f883 = hbusreq6 & v3a544de | !hbusreq6 & v8455ab;
assign v372421d = hmaster2_p & v3a5a6e6 | !hmaster2_p & v374158d;
assign v3a69248 = hlock6_p & v3753f1a | !hlock6_p & v8455ab;
assign v37c014e = hbusreq0_p & v373da69 | !hbusreq0_p & v3a6f4fc;
assign v3746063 = hbusreq0_p & v3a5600a | !hbusreq0_p & v8455ab;
assign v3a6f701 = jx0_p & v375178a | !jx0_p & v8455ab;
assign v375331e = hbusreq6_p & v3a667e7 | !hbusreq6_p & v8455ab;
assign v3a71453 = hbusreq2_p & v3a55e8e | !hbusreq2_p & v8455ab;
assign v2093018 = hmaster2_p & v377bfc0 | !hmaster2_p & v3a6f71a;
assign v3770bb9 = hgrant3_p & v376f0c1 | !hgrant3_p & v3a5c4d5;
assign v3a715ab = hgrant6_p & v375f653 | !hgrant6_p & v374a95d;
assign v37750e0 = jx0_p & v37510d7 | !jx0_p & v3741714;
assign v3a6437e = hmaster1_p & v377b6ce | !hmaster1_p & !v3a7159b;
assign v3a6efc1 = hmaster2_p & v3766487 | !hmaster2_p & v8455ab;
assign v3735e69 = hmaster0_p & v3a6e5f0 | !hmaster0_p & v376c85c;
assign v3a554b9 = hbusreq2 & v3a6f586 | !hbusreq2 & !v3a6f3cf;
assign v3734c75 = jx3_p & v3a61ad3 | !jx3_p & v37499c4;
assign v3a6fe33 = hbusreq4_p & v372e790 | !hbusreq4_p & v3a6ef22;
assign v3740f25 = hmaster1_p & v376d9ad | !hmaster1_p & v375874f;
assign v375d1fa = hbusreq2_p & v3745a47 | !hbusreq2_p & v37501fd;
assign v3752d10 = hbusreq3_p & v375f4c8 | !hbusreq3_p & !v8455ab;
assign v37572d0 = hmaster2_p & v3762ea7 | !hmaster2_p & v37386da;
assign v376489a = hlock4_p & v3778e71 | !hlock4_p & v3760854;
assign v376e06b = hbusreq3 & v373d8e5 | !hbusreq3 & v3736fdd;
assign v372da7e = hmaster1_p & v377845d | !hmaster1_p & v3759602;
assign v3a65716 = hbusreq4 & v37521ed | !hbusreq4 & !v8455ab;
assign v3a70ef4 = hbusreq4 & v3743a66 | !hbusreq4 & v2acaecc;
assign v3a5ee6e = hgrant2_p & v3a62e1b | !hgrant2_p & v8455ab;
assign v377a312 = hmaster2_p & b66740 | !hmaster2_p & !v372493b;
assign v3a578c3 = hbusreq8 & v3806b0b | !hbusreq8 & v373216d;
assign v376de0b = hburst0_p & v3730383 | !hburst0_p & v3a6f453;
assign v37794e5 = hmaster2_p & v3a64f5e | !hmaster2_p & !v8455ab;
assign v3a6a56e = hmaster2_p & v8455b0 | !hmaster2_p & v8455ab;
assign bfae74 = hbusreq5_p & v3a63831 | !hbusreq5_p & v3a5bb4e;
assign v374cb0f = hmaster0_p & v372abac | !hmaster0_p & v374b24a;
assign v3738253 = hgrant4_p & v372410a | !hgrant4_p & v3763b9e;
assign v3757388 = hlock3_p & v3a7081b | !hlock3_p & v3731ed2;
assign v377c49c = hmaster0_p & v3a58cfc | !hmaster0_p & !v3a6ad0b;
assign v3a5db97 = hgrant4_p & v8455ab | !hgrant4_p & v3a6e8a6;
assign v3740d4e = hmaster0_p & v37349b9 | !hmaster0_p & !v376ef9f;
assign v37568c9 = hmaster0_p & v3a6ef01 | !hmaster0_p & v373aa96;
assign v37661e4 = hbusreq7 & v376f549 | !hbusreq7 & v8455ab;
assign v3a70d48 = jx0_p & v380946e | !jx0_p & v3753fe6;
assign v3a62a71 = hgrant2_p & v8455e7 | !hgrant2_p & !v3a5cf3d;
assign v377261b = hlock0 & v3a70ad6 | !hlock0 & v3378302;
assign v3742290 = hbusreq6 & v3a70cc2 | !hbusreq6 & v3a6687c;
assign v3a712d8 = hmaster0_p & v3750883 | !hmaster0_p & v3763fec;
assign v3730f97 = hbusreq8_p & v376ae9f | !hbusreq8_p & v376e7c1;
assign v377f73c = hgrant6_p & v8455ab | !hgrant6_p & v1e37972;
assign v3a6fed3 = hbusreq3 & v376c8ea | !hbusreq3 & v373f0ee;
assign v3a6eb37 = hbusreq7_p & v3758526 | !hbusreq7_p & !v3771252;
assign v377ce30 = hgrant2_p & v372f09a | !hgrant2_p & v3a6f42c;
assign v377b4ad = hbusreq2 & v3737d44 | !hbusreq2 & !v8455ab;
assign v377c77a = hbusreq6 & v374f307 | !hbusreq6 & v8455b0;
assign v374c790 = hmaster1_p & v3731720 | !hmaster1_p & v3759cb9;
assign v37451db = hmaster3_p & v3759569 | !hmaster3_p & v8455ab;
assign v8bc0e2 = hmaster0_p & v3a6fb95 | !hmaster0_p & v375fb03;
assign v375f46d = hbusreq5_p & v3a704e3 | !hbusreq5_p & v373ae4a;
assign v37753dc = hlock5 & v3a70933 | !hlock5 & v375a6be;
assign v3a70c4d = hbusreq3 & v37482f8 | !hbusreq3 & v8455ab;
assign v37395e8 = hbusreq2_p & v3a6f3b1 | !hbusreq2_p & v8455ab;
assign v380921b = hgrant5_p & v8455ab | !hgrant5_p & v3a6fd87;
assign v3757921 = hlock0 & v3a70b92 | !hlock0 & v37438ab;
assign v3a7103d = hlock6 & v373e789 | !hlock6 & v39eb3bd;
assign v23fe0ff = hgrant5_p & v3769384 | !hgrant5_p & v3725403;
assign v2acaf2d = hmaster2_p & v376081b | !hmaster2_p & v3a6c549;
assign v37232c0 = hbusreq6 & v37482f8 | !hbusreq6 & !v377c3a1;
assign v376b56b = hbusreq8_p & v3a70578 | !hbusreq8_p & v3a5e0e5;
assign v3a61254 = busreq_p & v3a6f04a | !busreq_p & !v374c234;
assign v3a6f93b = hlock5_p & v372a599 | !hlock5_p & v37586e4;
assign v3a66ea9 = hbusreq0 & v3a6f37f | !hbusreq0 & v8455ab;
assign v3730cce = stateA1_p & v8455ab | !stateA1_p & !v3a5cf0b;
assign v3764383 = hmaster1_p & v3a60d50 | !hmaster1_p & v8455ab;
assign v3a70c51 = hbusreq5 & v3a6e1ed | !hbusreq5 & v3743efa;
assign v3765c08 = hlock5_p & v3738a87 | !hlock5_p & !v8455ab;
assign v3a6f8ae = hmaster2_p & v8455ab | !hmaster2_p & v377e9bb;
assign v3a675bc = hbusreq6_p & v376572c | !hbusreq6_p & v3727db9;
assign v376485c = hbusreq3 & v37567c7 | !hbusreq3 & v3a635ea;
assign v3a6ffd3 = hgrant4_p & v3a6f443 | !hgrant4_p & v3733027;
assign v373e2db = hgrant2_p & v8455b9 | !hgrant2_p & v3a6fe58;
assign v3a71093 = hmaster1_p & v38087c5 | !hmaster1_p & v3a6fd52;
assign v3a65287 = hmaster0_p & v3a70ca1 | !hmaster0_p & !v3a56512;
assign v37472f4 = hmaster1_p & v376c0c8 | !hmaster1_p & v3a6ffec;
assign v376a58a = hbusreq7 & v37520b7 | !hbusreq7 & v374d643;
assign v3a700c7 = hbusreq6_p & v3a563d3 | !hbusreq6_p & v8455ab;
assign v377da37 = hlock4_p & v87cef3 | !hlock4_p & v37395f5;
assign v375398e = hmaster0_p & v8455bf | !hmaster0_p & v3756820;
assign v374bdfe = hbusreq6_p & v3762333 | !hbusreq6_p & v8455ab;
assign v3a61f4c = hbusreq3_p & v3a6f539 | !hbusreq3_p & v8455ab;
assign v3a70eb8 = jx0_p & v3a6ef60 | !jx0_p & v374dd11;
assign v3770cf6 = hlock6 & v3759ca7 | !hlock6 & v37537ef;
assign v3a6ef21 = hmaster2_p & v3a6e31f | !hmaster2_p & v3759032;
assign v3731edf = hmaster3_p & v3806624 | !hmaster3_p & v374a795;
assign v37691ab = hbusreq5 & v3730e7d | !hbusreq5 & v3a62a6d;
assign v3779ba9 = hbusreq8 & v374148a | !hbusreq8 & v3a5666f;
assign v9c9e05 = hbusreq8_p & v3725bd2 | !hbusreq8_p & v3759dc9;
assign v375dc46 = hgrant2_p & v8455ba | !hgrant2_p & v377ac7e;
assign v375aceb = hbusreq5 & v3732775 | !hbusreq5 & v37c014f;
assign v3a70a92 = hgrant2_p & v3a637dc | !hgrant2_p & d27546;
assign v3a65db0 = start_p & v3a54fb2 | !start_p & !v37603af;
assign v372e44d = hmaster0_p & v375a3dd | !hmaster0_p & !v373e267;
assign v37363f8 = hmaster2_p & v373ad95 | !hmaster2_p & !v37346be;
assign v3a6e548 = hgrant4_p & v377d78b | !hgrant4_p & v3a5cd5c;
assign v3a6f329 = hgrant4_p & v3751081 | !hgrant4_p & v3777d39;
assign v3744a91 = hmaster0_p & v3759172 | !hmaster0_p & v3a5e371;
assign v375a68d = jx2_p & v372d0db | !jx2_p & v375c7b0;
assign v3a5f4a8 = hgrant8_p & v3767651 | !hgrant8_p & v3a65383;
assign hmaster2 = !v329f8b7;
assign v23fe217 = hmaster2_p & v3757b16 | !hmaster2_p & v3a655e9;
assign v3749760 = hgrant6_p & v3a6f8f6 | !hgrant6_p & v3a5a2be;
assign v3a626da = hmaster1_p & v3a6e124 | !hmaster1_p & v37386c0;
assign v377e9c9 = hmaster1_p & v3a66aa4 | !hmaster1_p & v37313e4;
assign v3726d7a = hbusreq1 & v3a64ee3 | !hbusreq1 & v8455ab;
assign v3a6757a = decide_p & d1331f | !decide_p & v8455e7;
assign v3a70e28 = hgrant4_p & v374db6a | !hgrant4_p & v3750d61;
assign v3753c73 = hgrant4_p & v8455ab | !hgrant4_p & v373031f;
assign v3779d06 = hgrant5_p & v8455ab | !hgrant5_p & v374d5fa;
assign v3a709b2 = hmaster2_p & v3730ffe | !hmaster2_p & v3a6f0f6;
assign v3a70e2e = hbusreq2_p & v3a2ae01 | !hbusreq2_p & v8455ab;
assign v3a709ea = hburst1 & v3a6ac2a | !hburst1 & v3a6f456;
assign cf45c3 = hbusreq2_p & v3751f72 | !hbusreq2_p & v3a641d5;
assign v376faab = hbusreq4_p & v38072fd | !hbusreq4_p & v3a6fc01;
assign v3731099 = hbusreq6_p & v377149d | !hbusreq6_p & v3768573;
assign v374bee4 = hbusreq3_p & v3759b9a | !hbusreq3_p & v3a63197;
assign v3a55526 = hbusreq6 & v3a70a23 | !hbusreq6 & v3a71019;
assign v375a268 = locked_p & v374b394 | !locked_p & v3577306;
assign v3778a55 = hbusreq8_p & v375a4a9 | !hbusreq8_p & v3730dc1;
assign v373828a = hbusreq4_p & v377ef6e | !hbusreq4_p & v3a53f53;
assign v3a707b2 = hmaster0_p & v3a7097d | !hmaster0_p & v3770cb8;
assign v3a61886 = hbusreq6_p & v3768383 | !hbusreq6_p & v372f16b;
assign v377f61c = hmaster0_p & v37380e2 | !hmaster0_p & !v37411c6;
assign v37660d9 = hmaster1_p & v2619ad7 | !hmaster1_p & v3759a08;
assign v37430c2 = hbusreq2 & v37300c9 | !hbusreq2 & v3778cdd;
assign v3a62aa3 = hmaster1_p & v1e37e29 | !hmaster1_p & v377f887;
assign v3a6ff6e = hmaster1_p & v2aca977 | !hmaster1_p & v3744151;
assign v3727e59 = hlock6_p & v375ecd5 | !hlock6_p & v8455ab;
assign v3a70130 = hbusreq0 & v3a6fab9 | !hbusreq0 & v3a56b4e;
assign v37345de = hmaster0_p & v3730398 | !hmaster0_p & v8455ab;
assign v3776454 = hmaster0_p & v37615a2 | !hmaster0_p & v3a5f43a;
assign v377efac = hbusreq2 & v3743da0 | !hbusreq2 & v3a6f5ea;
assign v3a705ad = hbusreq0_p & d44200 | !hbusreq0_p & v8455ab;
assign v3a55bf6 = hbusreq2 & v3a66051 | !hbusreq2 & v373f0ee;
assign v3a7004b = hmaster2_p & a0cf3e | !hmaster2_p & v8455ab;
assign v3a53c9d = hgrant2_p & v377097a | !hgrant2_p & v3723f24;
assign v3724a6d = hmaster1_p & v3757966 | !hmaster1_p & v374c9e9;
assign v3a659f5 = hbusreq5 & v375afe9 | !hbusreq5 & v372294a;
assign v3a70fae = hmaster2_p & v377b5f6 | !hmaster2_p & v3a6ff9e;
assign v3a64a7b = hbusreq8_p & v3756ebf | !hbusreq8_p & v372b6a1;
assign v3a59283 = hbusreq7_p & v3a575e5 | !hbusreq7_p & !v3778023;
assign v374801c = hmaster0_p & v3a5b289 | !hmaster0_p & v3a70bec;
assign be2682 = hbusreq6_p & v3a55755 | !hbusreq6_p & v8455ab;
assign v3739c94 = hbusreq4_p & v3a69cd8 | !hbusreq4_p & v3a7012e;
assign v375a92d = hmaster0_p & v3a70622 | !hmaster0_p & v3a5fd4a;
assign v3737a8b = hbusreq7 & v377bf7b | !hbusreq7 & v373c52e;
assign v3a6df32 = hgrant4_p & v8455ab | !hgrant4_p & !v373b76d;
assign v3a5dbd1 = hbusreq4_p & v37601a1 | !hbusreq4_p & v8455ab;
assign v37730bf = hgrant3_p & v3a70b92 | !hgrant3_p & v3724f24;
assign v373e8de = jx3_p & v3a5f375 | !jx3_p & !v37726b0;
assign v3768349 = hbusreq6_p & v3747302 | !hbusreq6_p & v3a5dc35;
assign v3760276 = hlock5 & v3a66c12 | !hlock5 & v3a6f610;
assign v372cfc2 = hgrant5_p & v373f0d2 | !hgrant5_p & v3a61ff4;
assign v377f78c = hlock5_p & v376f979 | !hlock5_p & !v372e44d;
assign v3731b33 = hbusreq2_p & v376f73c | !hbusreq2_p & !v3728e09;
assign v2acb06f = hbusreq5_p & v3777b5b | !hbusreq5_p & v3776fc5;
assign v372ce1e = hbusreq7 & v377c0c3 | !hbusreq7 & v376ae9f;
assign v372a027 = hbusreq7_p & v372e374 | !hbusreq7_p & v3a6f569;
assign v375ea89 = hbusreq0 & v373cf60 | !hbusreq0 & v37397f0;
assign v3258dc5 = hmaster0_p & v3a635ea | !hmaster0_p & v3a5f78a;
assign v3725b77 = hmaster0_p & v37646a9 | !hmaster0_p & v376b540;
assign v3a696ed = hbusreq1_p & v3723430 | !hbusreq1_p & v8455e7;
assign v3775687 = hmaster0_p & v3a70ef8 | !hmaster0_p & v377b2f3;
assign v3a6f5ff = hmaster1_p & v3a6e31f | !hmaster1_p & v3a6b5ba;
assign v3a65206 = hmastlock_p & v3751860 | !hmastlock_p & !v8455ab;
assign v3a7048a = locked_p & v3749dad | !locked_p & v3a637dc;
assign v3731202 = hbusreq7_p & v3a5b819 | !hbusreq7_p & v3741abd;
assign v3a6f650 = hmaster1_p & v8455ab | !hmaster1_p & v3742649;
assign v372de43 = hgrant6_p & v377938d | !hgrant6_p & v372ae4c;
assign v3752781 = hmaster1_p & v3762c7c | !hmaster1_p & v3a5cfbb;
assign v3a7079c = hmaster1_p & v3a70474 | !hmaster1_p & v8455ab;
assign v37676e0 = hmaster3_p & v375a025 | !hmaster3_p & v8455ab;
assign v3a6b1b9 = hmaster1_p & v3a60c82 | !hmaster1_p & v3777efb;
assign v3a5fc59 = hbusreq4 & v3a697f1 | !hbusreq4 & !v39ebbae;
assign v3a70cab = hmaster2_p & v3a53d1e | !hmaster2_p & !v377d2a0;
assign v3769820 = hmaster2_p & v373785d | !hmaster2_p & v3760ff4;
assign v376cfaa = hlock0_p & v2925c39 | !hlock0_p & !v8455ab;
assign v373e13a = hmaster2_p & v8455e7 | !hmaster2_p & !v3753f1a;
assign v3a6431f = hbusreq4 & v3a6f32f | !hbusreq4 & !v3a706ce;
assign v3a6f99c = hbusreq4_p & v3a5e7fe | !hbusreq4_p & v377af09;
assign v3809788 = hlock2 & v374809d | !hlock2 & v372ca44;
assign v37780cc = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3a603a1;
assign v3a5cb14 = hbusreq4 & v3723903 | !hbusreq4 & v23fe101;
assign v3a673d3 = hmaster0_p & v3a5902f | !hmaster0_p & v3a583b0;
assign v37408e4 = hmaster1_p & v3766d4b | !hmaster1_p & v373a26b;
assign v376e150 = hmaster0_p & v376f8ba | !hmaster0_p & !v3a713a7;
assign v3a57eae = hmaster1_p & v37702f3 | !hmaster1_p & v377b8fb;
assign v3764ee3 = hmaster0_p & v376d9c6 | !hmaster0_p & v3760513;
assign v3774524 = hmaster2_p & v377b774 | !hmaster2_p & v373389a;
assign v3a6497b = hmaster2_p & v373e474 | !hmaster2_p & v375a1ab;
assign v3770c9d = hbusreq6_p & v1e374cc | !hbusreq6_p & v3725a56;
assign v37507da = hlock2 & v3a5cef4 | !hlock2 & v372777c;
assign v377f46e = hmaster1_p & v3a5642f | !hmaster1_p & !v376f051;
assign v9342d1 = jx1_p & v3a6f9bb | !jx1_p & v375d366;
assign v376a4c0 = hbusreq3 & v8455ab | !hbusreq3 & !v373aecf;
assign v375f106 = jx0_p & v8455ab | !jx0_p & v37586e2;
assign v37594ae = jx0_p & v3756234 | !jx0_p & !v3776cda;
assign v373511d = hgrant4_p & v3a57959 | !hgrant4_p & v377e8da;
assign v3a54222 = hbusreq7 & v3a64e75 | !hbusreq7 & v376195b;
assign v3a70ac0 = hbusreq6_p & v375208a | !hbusreq6_p & v374a8df;
assign v3a61c49 = hlock4_p & v28896da | !hlock4_p & v3750dd3;
assign v3a63028 = hbusreq2_p & v372ec1c | !hbusreq2_p & v3a69487;
assign v3724112 = hbusreq0_p & ad2d05 | !hbusreq0_p & v8455ab;
assign v3762806 = hbusreq5 & v372d538 | !hbusreq5 & v2acaed7;
assign v2acaf9d = hbusreq8_p & v3a712b9 | !hbusreq8_p & v8455ab;
assign v3a6f728 = hbusreq5_p & v374e0b8 | !hbusreq5_p & v3255a0c;
assign v3a5d8a9 = hmaster0_p & v8455ab | !hmaster0_p & !v372809d;
assign v3735d6f = hmaster2_p & v37770ed | !hmaster2_p & v8455ca;
assign v3a5aaf9 = hmaster2_p & v3a59e1c | !hmaster2_p & v8455b0;
assign v374eec1 = hmaster3_p & v3774cf5 | !hmaster3_p & v3763e92;
assign v3a710ea = hmaster1_p & v372685c | !hmaster1_p & v3747271;
assign v377e851 = hbusreq7 & v955d7b | !hbusreq7 & v8455ab;
assign v3a706c0 = hready & v373b288 | !hready & v3a635ea;
assign v373132b = hgrant0_p & v8455b3 | !hgrant0_p & v3749207;
assign v3a7094d = hbusreq2_p & v3a658be | !hbusreq2_p & v8455b0;
assign v3775d1d = hbusreq6 & v37274c2 | !hbusreq6 & !v8455b5;
assign v3768a41 = hbusreq6_p & v3a6fce5 | !hbusreq6_p & v8455ab;
assign v3738dc0 = hmaster0_p & v3a5bf5f | !hmaster0_p & v3a70097;
assign v37674a5 = hbusreq6_p & v3754543 | !hbusreq6_p & v372f87f;
assign v3a6fc60 = hgrant2_p & v8455b9 | !hgrant2_p & v3a6f7fb;
assign v3a6324b = hbusreq6 & v3779f67 | !hbusreq6 & v8455ab;
assign v3a64d23 = hgrant2_p & v3768c3c | !hgrant2_p & v376a7e8;
assign v3723118 = stateA1_p & v3a6efc9 | !stateA1_p & a81487;
assign v3a6ef18 = hlock2_p & v372a98e | !hlock2_p & !v8455ab;
assign v3a5cfac = hbusreq3_p & v3762fc3 | !hbusreq3_p & v8455ab;
assign v3751e09 = hgrant3_p & v37645ec | !hgrant3_p & v3a6e463;
assign v3a70f48 = hgrant6_p & v375a268 | !hgrant6_p & v3764df7;
assign v37232bd = hlock0_p & v3730627 | !hlock0_p & v3770187;
assign v3a7122f = hmaster0_p & v8455ab | !hmaster0_p & v8455dd;
assign v3737298 = hmaster1_p & v3730e01 | !hmaster1_p & v376055d;
assign v375af5d = hbusreq6 & v3a5f0cf | !hbusreq6 & v8455ab;
assign v37730ff = hlock5_p & v3754018 | !hlock5_p & v3a53904;
assign v3a71656 = hbusreq5_p & v377bd9b | !hbusreq5_p & v3766445;
assign v3731eff = hbusreq6_p & v3a635ea | !hbusreq6_p & v3743c51;
assign v376daf2 = hbusreq5 & v35b987f | !hbusreq5 & !v374e0f6;
assign v3a6fabf = hmaster0_p & v3772c5a | !hmaster0_p & v3774878;
assign v375d134 = hgrant6_p & v374352b | !hgrant6_p & v3731a29;
assign v3a59d59 = hgrant6_p & v3767463 | !hgrant6_p & v373ffa0;
assign v3a2975f = hbusreq0 & v3a6f5ea | !hbusreq0 & v8455ab;
assign v3a6f65e = hmaster0_p & v375945f | !hmaster0_p & v37429c2;
assign v3734374 = hmaster2_p & v8f695f | !hmaster2_p & v37261b3;
assign v3a577ed = hgrant7_p & v8455ab | !hgrant7_p & v3a5bc70;
assign v3a70bd0 = hlock3_p & v3742ef6 | !hlock3_p & v37509c7;
assign v374d1ed = hmaster1_p & v375a4a0 | !hmaster1_p & v372bd2b;
assign v3a6a6c1 = hbusreq4 & a25d5b | !hbusreq4 & v8455ab;
assign v3a6885a = hburst1 & v3a5f308 | !hburst1 & v3a671f4;
assign v374fa2a = hmaster3_p & v3a7003d | !hmaster3_p & v3745c20;
assign v3765224 = hlock7 & v374ef3e | !hlock7 & v377b647;
assign v373f694 = hmaster2_p & v3763f95 | !hmaster2_p & v3a6dc08;
assign v3751831 = hbusreq3 & v3763d3a | !hbusreq3 & v37427d3;
assign v3a54f8a = hmaster2_p & v3734967 | !hmaster2_p & v3a60787;
assign v374571d = hbusreq6_p & v3a6a6b4 | !hbusreq6_p & v8455ab;
assign v3760d46 = hbusreq4_p & v375ed63 | !hbusreq4_p & v3a6f29c;
assign v377d408 = hlock1_p & v3763f8b | !hlock1_p & !v8455ab;
assign v3771be4 = hmaster2_p & v3764276 | !hmaster2_p & !v8455ab;
assign v37325e0 = hmaster1_p & v377989c | !hmaster1_p & v377098c;
assign v3731159 = hmaster1_p & v377984a | !hmaster1_p & v3735bbc;
assign v375b61a = hmaster3_p & v3724579 | !hmaster3_p & v3a6b161;
assign v373b0be = hgrant6_p & v375f653 | !hgrant6_p & v3a70b55;
assign v3a64102 = hbusreq8 & v3a5ec6b | !hbusreq8 & v376f51a;
assign v377933b = hbusreq8 & v377281c | !hbusreq8 & v3a6f369;
assign v3809b0a = hmaster1_p & v8455ab | !hmaster1_p & v377133f;
assign v3a70a99 = hmaster0_p & v372ded7 | !hmaster0_p & v3773ca3;
assign v3a710de = hbusreq5_p & v3a63f9a | !hbusreq5_p & v37725c6;
assign v374a46d = hmaster2_p & v8455ab | !hmaster2_p & v3755791;
assign v3768828 = hmaster0_p & v3a54c2e | !hmaster0_p & v377c71d;
assign v3745de0 = hlock8 & v374b0d9 | !hlock8 & v3a5cf6f;
assign v3731487 = hbusreq3_p & v3a6f8f5 | !hbusreq3_p & !v8455ab;
assign v3769b7e = hmaster0_p & v3a70a3e | !hmaster0_p & v3764d26;
assign v39a53b3 = hbusreq2_p & v377327b | !hbusreq2_p & v377c7b2;
assign v372a77f = hlock5 & v3a6ae0f | !hlock5 & v3744a9c;
assign v3a6eb44 = hbusreq6 & v3756e01 | !hbusreq6 & v375bfa6;
assign v377ea86 = hbusreq3_p & v39a5265 | !hbusreq3_p & v8455e1;
assign v37616e0 = hgrant2_p & v3809ee9 | !hgrant2_p & v3a55b93;
assign v3a6fd62 = hbusreq5 & v376a6f1 | !hbusreq5 & v3728392;
assign v3761340 = hbusreq8_p & v376a59f | !hbusreq8_p & a0a219;
assign v3733aa5 = hgrant4_p & v3a5ed4b | !hgrant4_p & v3775654;
assign v3a7093a = hbusreq6 & v3a6fce6 | !hbusreq6 & v8455cb;
assign v372c614 = hbusreq6 & v3a61604 | !hbusreq6 & v8455ab;
assign v869938 = hmaster0_p & v3a6d499 | !hmaster0_p & v37710a1;
assign v3724af9 = hbusreq0 & v37652a5 | !hbusreq0 & v8455ab;
assign v376b363 = hbusreq3_p & v3a60787 | !hbusreq3_p & !v377cfd9;
assign v37532ee = hmaster0_p & v372c638 | !hmaster0_p & v37281fb;
assign v375580b = hgrant5_p & v8455ab | !hgrant5_p & v3a6bc32;
assign v37596f3 = hlock7_p & v3a704fe | !hlock7_p & v8455c7;
assign v3a59df2 = hbusreq6_p & v376bb27 | !hbusreq6_p & v377bfb6;
assign v3776917 = hmaster0_p & v3723477 | !hmaster0_p & v3a66615;
assign v3a694bb = hbusreq6_p & v3734dd8 | !hbusreq6_p & v8455ab;
assign v3760690 = hbusreq5_p & v37744a3 | !hbusreq5_p & v3a713c5;
assign v3a713ab = hlock5_p & v3a6a2d7 | !hlock5_p & v8455ab;
assign v3a6f72a = hgrant2_p & v3742033 | !hgrant2_p & v372a4c4;
assign v3a6f925 = hgrant5_p & v3a6ff1f | !hgrant5_p & v3735749;
assign v3772bff = hmaster0_p & v3747fbc | !hmaster0_p & !v373f2a6;
assign v3a713a7 = hmaster2_p & v8455ab | !hmaster2_p & v3731bc8;
assign v3a709b9 = hmaster2_p & v8455ab | !hmaster2_p & !v373006f;
assign v3a705ec = hmaster2_p & v37481e4 | !hmaster2_p & v375884e;
assign v190eb62 = hready_p & v37255d6 | !hready_p & !v3722e5a;
assign v3a603bb = hbusreq3_p & v3747302 | !hbusreq3_p & v373e521;
assign v37322ca = hbusreq4 & v3730ae3 | !hbusreq4 & !v8455ab;
assign v3727187 = hbusreq5_p & v3a6fdb7 | !hbusreq5_p & v375d94c;
assign v3a5cf5e = hmaster2_p & c8a454 | !hmaster2_p & v3a5ba28;
assign v3a712c0 = hmaster0_p & v8455ab | !hmaster0_p & v3a71282;
assign v3a5a05d = hbusreq5_p & v375eeb9 | !hbusreq5_p & v37244f4;
assign v377d39f = hbusreq2_p & v3a6b4d7 | !hbusreq2_p & v3a6fdf4;
assign v3744b16 = jx3_p & v3775630 | !jx3_p & v8455ab;
assign v373fc77 = hready_p & v3a70772 | !hready_p & v3985138;
assign v3a6f7f9 = hbusreq3 & v37441b5 | !hbusreq3 & v37775d9;
assign v3a6f122 = hlock5_p & v376d979 | !hlock5_p & v3a6f387;
assign v3758b25 = hbusreq8_p & b0b0c6 | !hbusreq8_p & v3770be6;
assign v375bdaf = hlock0 & v373031f | !hlock0 & v376d7c6;
assign v3a6fe92 = hbusreq8 & v3a69fe5 | !hbusreq8 & v37613b3;
assign v375ed43 = hmaster1_p & v3a6f352 | !hmaster1_p & v3a6c573;
assign v3a6f318 = hbusreq5_p & v3772083 | !hbusreq5_p & v3766222;
assign v3a70b61 = hmaster1_p & v3a6ffca | !hmaster1_p & v372efc8;
assign v376ef36 = hbusreq2_p & v3a70dd6 | !hbusreq2_p & v3a6a7b4;
assign v1e373d9 = hgrant5_p & v374b330 | !hgrant5_p & v380705b;
assign v377018e = hbusreq2 & v376111d | !hbusreq2 & v8455ab;
assign v3a63556 = hmaster0_p & v3779069 | !hmaster0_p & v376db34;
assign v377b5f4 = hbusreq7_p & v3742395 | !hbusreq7_p & v3769870;
assign v3a5af86 = hbusreq3 & v3a5b68a | !hbusreq3 & !v8455ab;
assign v3762414 = hbusreq1 & v3a5600a | !hbusreq1 & v3773b23;
assign v3771fe5 = hready_p & v3a5f5d0 | !hready_p & !v375a68d;
assign v37705de = hgrant2_p & v376f2f8 | !hgrant2_p & v37251cc;
assign v3757ad8 = hmaster0_p & v3a641d5 | !hmaster0_p & v37710a1;
assign v3768fb7 = hmaster2_p & v3a706fe | !hmaster2_p & v3730986;
assign v3737647 = hbusreq0 & v3a7073b | !hbusreq0 & v3764601;
assign v3a5fcfc = start_p & v3730a0f | !start_p & v3a7111f;
assign v3745dc7 = hgrant3_p & v3734bc3 | !hgrant3_p & v8455ab;
assign v3741572 = hlock7 & v37494a7 | !hlock7 & v372f56c;
assign v374ad1e = hgrant3_p & v374f307 | !hgrant3_p & v23fd7d9;
assign v3a628ef = jx0_p & v380958f | !jx0_p & v3a6eb37;
assign v3a6fe0d = hbusreq1_p & v373b80b | !hbusreq1_p & v8455ab;
assign v373c856 = hlock0 & v37285eb | !hlock0 & v1e374ce;
assign v3a6eb0a = hlock0 & v377b946 | !hlock0 & v3753526;
assign v374bce0 = hbusreq0 & v3750c12 | !hbusreq0 & v3a700b7;
assign v2925d19 = hgrant6_p & v376f2a7 | !hgrant6_p & v37404da;
assign v375a367 = hmaster0_p & v3a68d0e | !hmaster0_p & v3a7152d;
assign v3747d33 = hmaster0_p & v3a706d5 | !hmaster0_p & v372dcf7;
assign v3762858 = hmaster2_p & v35772a6 | !hmaster2_p & v3a6eb39;
assign v3a70a60 = stateG10_1_p & v8455ab | !stateG10_1_p & v372df69;
assign v376a2df = hmaster2_p & v8455c3 | !hmaster2_p & v372e4cf;
assign v375c24b = hbusreq7_p & v3a5a4c0 | !hbusreq7_p & v376faf0;
assign v3743c40 = hbusreq4_p & v37430e7 | !hbusreq4_p & v3a6f240;
assign v374c288 = hbusreq5 & v372f478 | !hbusreq5 & v3742cd5;
assign v372cbac = hmaster1_p & v375c7b9 | !hmaster1_p & !v38074a8;
assign v3739f22 = hbusreq2_p & v37765e1 | !hbusreq2_p & v3a62e1e;
assign v377db21 = hbusreq2_p & v376c569 | !hbusreq2_p & v3809583;
assign v3772612 = hmaster1_p & v3743ff2 | !hmaster1_p & v374546c;
assign v3747b97 = hbusreq5 & v377e59a | !hbusreq5 & v3743fc1;
assign v8455c9 = hbusreq6_p & v8455ab | !hbusreq6_p & !v8455ab;
assign v376938e = hbusreq4 & v37606e5 | !hbusreq4 & v8455ab;
assign v3757f9b = hgrant0_p & v3a5be72 | !hgrant0_p & v8455ab;
assign v3a6f593 = hmaster1_p & v375c65f | !hmaster1_p & v3734658;
assign v921bc8 = hbusreq6_p & v377eaf2 | !hbusreq6_p & v3735512;
assign v3a692c3 = hmaster2_p & v3734967 | !hmaster2_p & v3733d6e;
assign v3a6f114 = hmaster2_p & v373ab12 | !hmaster2_p & !v8455c3;
assign v376d6ef = hmaster2_p & v377bf71 | !hmaster2_p & v37514c7;
assign v3a7050d = jx0_p & v3734279 | !jx0_p & v3729c9a;
assign v3726ea3 = hmaster0_p & v3728c5b | !hmaster0_p & v3a70666;
assign v37390f9 = hgrant4_p & v37484e0 | !hgrant4_p & v37282c1;
assign v377c039 = hbusreq2_p & v3761efb | !hbusreq2_p & c0d46a;
assign v3a5c700 = hlock2 & v375ddb7 | !hlock2 & v3a5fcbc;
assign v375d434 = hbusreq5_p & v3a6b27d | !hbusreq5_p & v377e056;
assign v2acaf23 = hgrant0_p & v3a5d822 | !hgrant0_p & v3a5ca02;
assign v37554b1 = hbusreq4_p & v3a679ae | !hbusreq4_p & v3a6f896;
assign v3a66c84 = hbusreq5_p & v372cafb | !hbusreq5_p & !v376bc8c;
assign v3767852 = hmaster1_p & v3757261 | !hmaster1_p & v3737f8b;
assign v37350e9 = jx0_p & v3739077 | !jx0_p & v8455ab;
assign v3774a1e = hbusreq0 & v3730afc | !hbusreq0 & v3a6bdd1;
assign v3768082 = hmaster1_p & v374e5ad | !hmaster1_p & v8455ab;
assign v3a70c63 = hgrant6_p & v373cc5c | !hgrant6_p & v3767b98;
assign v375d715 = hgrant2_p & v376b5f8 | !hgrant2_p & d1f2e2;
assign v2acb088 = hbusreq3_p & v373588a | !hbusreq3_p & !v376d9d4;
assign v3731999 = hmaster0_p & v3a711e4 | !hmaster0_p & !v37712b7;
assign v373785d = hbusreq6_p & v3a635ea | !hbusreq6_p & v377c6b3;
assign v373c2ec = hbusreq2_p & v3747302 | !hbusreq2_p & v3778b8d;
assign v377af47 = hbusreq4 & v37366d0 | !hbusreq4 & v8455ab;
assign v373d142 = hbusreq8 & v3a71101 | !hbusreq8 & v3807414;
assign v3a677ce = hmaster2_p & v3a70641 | !hmaster2_p & v3806db7;
assign v3749ece = hgrant1_p & v8455ab | !hgrant1_p & !v374e78f;
assign v375c525 = hbusreq8_p & v3a5cae1 | !hbusreq8_p & !v8455ab;
assign v374c73c = hmaster0_p & v3746d52 | !hmaster0_p & !v37bfc8b;
assign v38079d7 = hgrant3_p & v8455ab | !hgrant3_p & v3770f51;
assign v3776022 = hbusreq4 & v373cd16 | !hbusreq4 & v8455ab;
assign v3a573e3 = hbusreq1_p & v3a635ea | !hbusreq1_p & !v3a709a0;
assign v3a643ef = hbusreq7_p & v3a6f590 | !hbusreq7_p & v3a674c9;
assign v3a70f7a = hbusreq4_p & v38072fd | !hbusreq4_p & v375ae91;
assign v373fee1 = hgrant2_p & v8455ba | !hgrant2_p & v3a5797b;
assign v375b7e1 = hbusreq6 & v3a5dcfc | !hbusreq6 & v3a635ea;
assign v3a70ae5 = hgrant5_p & v8455ab | !hgrant5_p & v3728d9c;
assign v3a6f98e = hbusreq7 & v375c009 | !hbusreq7 & !v376fa50;
assign v3a6eb1e = hlock6 & v3a6a322 | !hlock6 & v374d8bb;
assign v3755045 = hlock5_p & v37510b9 | !hlock5_p & !v8455ab;
assign v3a6c6f6 = hlock4 & v372e618 | !hlock4 & v3778390;
assign v3a703b1 = hmaster2_p & v372c546 | !hmaster2_p & v3a6f1e4;
assign v37790c8 = hmaster0_p & v377e298 | !hmaster0_p & v37458ca;
assign v3749e1c = hmastlock_p & v37690db | !hmastlock_p & v8455ab;
assign v3a603a1 = hbusreq0 & v3a56d86 | !hbusreq0 & v3a6651d;
assign v3734c7e = hgrant6_p & v3a5cc17 | !hgrant6_p & v3a62539;
assign v3745754 = hmaster0_p & v3a7117c | !hmaster0_p & v3776cbb;
assign v374e5e9 = hbusreq8_p & v3a635ea | !hbusreq8_p & v3753e28;
assign v373374d = hgrant2_p & v3a6c33a | !hgrant2_p & !v377005e;
assign v3a6cd1b = start_p & v845605 | !start_p & v3a7111f;
assign v3726204 = hbusreq6_p & v37414d1 | !hbusreq6_p & !v372df2a;
assign v3753389 = hmaster0_p & v376a31b | !hmaster0_p & v376e7f5;
assign v372f9c3 = hbusreq2 & v3a70e03 | !hbusreq2 & v8455ab;
assign v3a6ff93 = hmaster2_p & v374513e | !hmaster2_p & v8455ab;
assign v3a71389 = hbusreq6_p & v3734918 | !hbusreq6_p & v3a657bf;
assign v375b7fa = hgrant2_p & v8455ba | !hgrant2_p & v3729b37;
assign v3758c0d = hbusreq0_p & v3a5891c | !hbusreq0_p & v3759032;
assign v3a56d2e = hbusreq7_p & v3779e38 | !hbusreq7_p & v3738641;
assign v3a713d5 = hbusreq5 & v373e219 | !hbusreq5 & v374c6b8;
assign v374f838 = hgrant5_p & v3a70578 | !hgrant5_p & v372c016;
assign v37263c1 = hmaster0_p & v377c7c0 | !hmaster0_p & v3729a69;
assign v3751c65 = jx0_p & v376f39f | !jx0_p & v3776ff3;
assign v3747302 = locked_p & v8455ab | !locked_p & !v35772a5;
assign v3809892 = hmaster0_p & v8a94c2 | !hmaster0_p & !v374514c;
assign v3a6fb84 = hgrant0_p & v8455ab | !hgrant0_p & v3a6e7a7;
assign c7d478 = hbusreq4_p & v37337b3 | !hbusreq4_p & v3778528;
assign v3a6f3ef = hlock5_p & v377e5e1 | !hlock5_p & !v8455ab;
assign v37bfca2 = hbusreq3 & v3a676d6 | !hbusreq3 & v8455ab;
assign v376fb18 = hgrant3_p & v3a67ab9 | !hgrant3_p & v8455ab;
assign v3a601a0 = hbusreq2_p & v3a6ef18 | !hbusreq2_p & !v8455ab;
assign v3a6c2a9 = hbusreq6_p & v3726838 | !hbusreq6_p & !v8455ab;
assign v3a6f4ba = hgrant4_p & v3a5a807 | !hgrant4_p & v377b2d0;
assign v374e8b4 = hmaster2_p & v3731857 | !hmaster2_p & !v3777b2e;
assign v3766986 = hlock5 & v376bfb9 | !hlock5 & v3a65ce7;
assign v375b019 = hmaster2_p & v8455ab | !hmaster2_p & !v373c3ba;
assign v376bb81 = hlock8_p & v20d166d | !hlock8_p & v3754afa;
assign v373e484 = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v372adaa;
assign v37358f3 = hgrant5_p & v377af89 | !hgrant5_p & v3a6f526;
assign v3a6620b = hlock0 & v373bd6c | !hlock0 & v377d6d3;
assign v37681ec = hgrant5_p & v3a63cf5 | !hgrant5_p & v3a60bc1;
assign v37500ac = hbusreq2 & v3a6672b | !hbusreq2 & v8455ab;
assign v3767399 = stateG10_1_p & v3a6f252 | !stateG10_1_p & v376eb2b;
assign cd743d = hmaster0_p & v3728962 | !hmaster0_p & v3a296dc;
assign v3a60888 = hmaster0_p & v374e985 | !hmaster0_p & v3723be4;
assign v372fecf = hbusreq4 & v3741338 | !hbusreq4 & v3a5741c;
assign v372d643 = hbusreq5 & v3759aca | !hbusreq5 & v1e37cba;
assign v3777d6c = hmaster0_p & v8455ab | !hmaster0_p & v3a6dc60;
assign v3a70a6d = hbusreq0_p & v3a67e64 | !hbusreq0_p & !v3a5952d;
assign v37656cd = hbusreq8 & v3a7092f | !hbusreq8 & v8455ab;
assign v3a6fb2b = hbusreq2_p & v8455bf | !hbusreq2_p & v3763a20;
assign v3777536 = hmaster2_p & v373b7c5 | !hmaster2_p & v3a6f43a;
assign v39a5350 = hgrant0_p & v3a705f7 | !hgrant0_p & v37777bf;
assign v3a711c6 = hlock5_p & v3743b12 | !hlock5_p & cfaa3a;
assign v3a5dd8a = hlock8 & v2aca987 | !hlock8 & v3779014;
assign v3a63a18 = hmaster2_p & v3a635ea | !hmaster2_p & v376358f;
assign v376209f = hbusreq7_p & v37341ff | !hbusreq7_p & !v375c28e;
assign v3744037 = start_p & v845605 | !start_p & v3730383;
assign v3776cb6 = hlock5_p & v372bd5e | !hlock5_p & !v37419b2;
assign v37799f4 = hgrant4_p & v8455ab | !hgrant4_p & v3733d71;
assign v3747dfc = hgrant3_p & v37506fb | !hgrant3_p & v374d4c1;
assign v3747c90 = hlock4 & v3759ef7 | !hlock4 & v3755abd;
assign v3730b5a = hmaster3_p & v37266bd | !hmaster3_p & v3734a96;
assign v3735c5f = hmaster2_p & v3763175 | !hmaster2_p & v8455b0;
assign v375b2e2 = hbusreq0 & v376d1e2 | !hbusreq0 & v8455ab;
assign v3a6fba3 = hgrant5_p & v373ad69 | !hgrant5_p & v37262ab;
assign v3723220 = hmaster1_p & cd0aed | !hmaster1_p & v3a6db7f;
assign v377e934 = hbusreq4 & v37270d9 | !hbusreq4 & v8455e7;
assign v3a6f29a = hbusreq0 & v375ca93 | !hbusreq0 & v8455ab;
assign v3a66559 = hbusreq1_p & b4fa3c | !hbusreq1_p & v3a69d9b;
assign v3761da2 = hbusreq7 & v375ad90 | !hbusreq7 & v3750fa9;
assign v3a63cf5 = hmaster1_p & v3a5c945 | !hmaster1_p & v3730a73;
assign v3733174 = hmaster0_p & v8455ab | !hmaster0_p & !v3a5c3ba;
assign v374b36f = hbusreq5_p & v37480ad | !hbusreq5_p & !v375f708;
assign v3a7042a = hbusreq6_p & v374aca8 | !hbusreq6_p & v372d48d;
assign v3769bec = hbusreq4_p & v3741e5c | !hbusreq4_p & v374a23b;
assign v3739681 = hmaster1_p & v372b1dc | !hmaster1_p & v37430f5;
assign v3737695 = hlock8_p & v3778baf | !hlock8_p & v374fe51;
assign v3736b71 = hgrant4_p & v373f17f | !hgrant4_p & v376e17a;
assign v3a7046e = hlock5_p & v3a71159 | !hlock5_p & v375fbef;
assign v3a70bce = hbusreq1_p & v1e37d3f | !hbusreq1_p & v3a6f32a;
assign v3736d43 = hlock0 & v374f35a | !hlock0 & v23fdf30;
assign v37317c4 = hbusreq4_p & v3a68407 | !hbusreq4_p & v8455ab;
assign v3a6fa4f = stateG2_p & v8455ab | !stateG2_p & v2092f0a;
assign v3770dbf = hgrant7_p & v3a6f7a9 | !hgrant7_p & v37689aa;
assign v372fd45 = hgrant2_p & v377b6ce | !hgrant2_p & v3747035;
assign v3742122 = hbusreq2_p & v3754eb1 | !hbusreq2_p & v8455ab;
assign v3a712b6 = hgrant3_p & v3a7029b | !hgrant3_p & v3a5c366;
assign v3a5dc35 = hlock6 & v3a71582 | !hlock6 & v372310a;
assign v376bbbe = hmaster2_p & v3a676ce | !hmaster2_p & v3a6fb68;
assign v3a58d67 = hlock0 & v3a64af7 | !hlock0 & v3a6f160;
assign v372ab63 = hmaster1_p & v3a6fc99 | !hmaster1_p & v374f5a1;
assign v375022e = hbusreq6 & v3743040 | !hbusreq6 & v8455ab;
assign v372d19a = hbusreq0 & v3a6784d | !hbusreq0 & v372a1b4;
assign v3a562a9 = locked_p & v37624b2 | !locked_p & v8455ab;
assign v3a70a68 = hbusreq1_p & v360d1ca | !hbusreq1_p & v3730bb7;
assign v3807071 = hmastlock_p & v3738cfc | !hmastlock_p & !v8455ab;
assign v3a70a2c = hmaster1_p & v3a64ebb | !hmaster1_p & v3a6b90e;
assign v3727e33 = hmaster2_p & v3807f45 | !hmaster2_p & v3a70b17;
assign v3a665b4 = hgrant5_p & v3742146 | !hgrant5_p & v3743e4a;
assign v375f5c1 = hmaster1_p & v374f307 | !hmaster1_p & v373f3dd;
assign v374a528 = jx0_p & v3a55ec0 | !jx0_p & v3728bff;
assign v3a5fc48 = hmaster0_p & v3a70c3e | !hmaster0_p & v374b887;
assign v375d4d9 = hbusreq6 & v37526d6 | !hbusreq6 & v377c6b3;
assign v37253a5 = hbusreq8_p & v3a7042c | !hbusreq8_p & v3a5ef2e;
assign v3724bf3 = hlock5 & v37337e7 | !hlock5 & v3a5ebbf;
assign v372838e = hmaster2_p & a96343 | !hmaster2_p & v3765740;
assign v375524c = hmaster1_p & v3734914 | !hmaster1_p & v3a6fd9b;
assign v3a66835 = hmaster2_p & v3a5e817 | !hmaster2_p & !v8455ab;
assign v360bc71 = hgrant4_p & v8455ab | !hgrant4_p & v3a71684;
assign v37317f1 = hbusreq6_p & v37617a9 | !hbusreq6_p & v373dc73;
assign v3755785 = hbusreq6_p & v376648e | !hbusreq6_p & !v37433ff;
assign v3748332 = hgrant2_p & v8455ab | !hgrant2_p & v3a71006;
assign v3759ef7 = hbusreq4 & v3755abd | !hbusreq4 & v3a6a934;
assign v376a8be = hmaster0_p & v3a6e065 | !hmaster0_p & v37455cd;
assign v375fa71 = hbusreq6_p & v3a714ff | !hbusreq6_p & v3a6e305;
assign v3757253 = hbusreq3_p & v373e296 | !hbusreq3_p & v373b288;
assign v3a67af1 = hmaster1_p & v3a6c793 | !hmaster1_p & v376f9ac;
assign v375c10c = hlock7 & v372c00a | !hlock7 & v3779b5b;
assign v3a54c8d = hbusreq3_p & v376f56d | !hbusreq3_p & !v8455ab;
assign v3733993 = hbusreq5 & v360d0c7 | !hbusreq5 & !v8455ab;
assign v3a62b35 = hbusreq7 & v373402f | !hbusreq7 & v3768734;
assign v3a70e75 = hlock6 & v37366fc | !hlock6 & v3809788;
assign v3a70d32 = hgrant6_p & v8455ca | !hgrant6_p & v3776e85;
assign v372ec9f = hbusreq5_p & v3777d7c | !hbusreq5_p & v37273f6;
assign v374f857 = hmaster2_p & v375e60f | !hmaster2_p & v3a6b0c7;
assign v3a6f585 = hbusreq4_p & v3775a4a | !hbusreq4_p & v375c05f;
assign v3a6f30f = hgrant2_p & v37639c6 | !hgrant2_p & v374cb05;
assign v3a5a051 = hlock0 & v37790fb | !hlock0 & v3a70704;
assign v377e002 = hgrant4_p & v1e37b99 | !hgrant4_p & !v3775269;
assign v3a69057 = hmaster1_p & v39a53e9 | !hmaster1_p & v3a557a1;
assign v3739884 = hbusreq6_p & v3a68b34 | !hbusreq6_p & v3762886;
assign v372a421 = hmaster1_p & v3a635ea | !hmaster1_p & v37497d6;
assign v372dcd4 = hbusreq3_p & v376ea4a | !hbusreq3_p & !v3728e09;
assign v37341b2 = hbusreq6_p & v373a29c | !hbusreq6_p & v372d1bf;
assign v3a64e05 = hbusreq6_p & v37401f0 | !hbusreq6_p & v374ea45;
assign v3a6f7d0 = hbusreq5 & v3a697d2 | !hbusreq5 & v374b549;
assign v3756883 = hbusreq0 & v37297b2 | !hbusreq0 & v374638c;
assign v374d6bd = hmaster2_p & v8455ab | !hmaster2_p & v3768091;
assign v3a58cb2 = hgrant8_p & v374e7f2 | !hgrant8_p & v374d802;
assign v37430fb = hmaster2_p & v3769740 | !hmaster2_p & v3750edc;
assign v3778138 = hlock5 & v3a6708d | !hlock5 & v3740762;
assign v37445f1 = hlock6 & v3733dd8 | !hlock6 & v3a5ef89;
assign v3a583cd = hmaster1_p & v8455ab | !hmaster1_p & d9e2a4;
assign v3766dcc = hmaster2_p & v3767b70 | !hmaster2_p & v3a67de3;
assign v3769923 = hmaster2_p & v3a703bf | !hmaster2_p & v372b4cb;
assign v3a6ac94 = stateG2_p & v8455ab | !stateG2_p & v3a71137;
assign v372c28d = hbusreq5_p & v373b9ab | !hbusreq5_p & v3a6fa04;
assign v3a58134 = hgrant6_p & v3727b41 | !hgrant6_p & v3a7037c;
assign v3752bcc = hgrant0_p & v8455ab | !hgrant0_p & v37296db;
assign v3a6fdf7 = hgrant3_p & v375c1d1 | !hgrant3_p & v374a97f;
assign v372d86d = hmaster3_p & c76b50 | !hmaster3_p & v375b6fe;
assign v3731e91 = hbusreq6_p & v3a6f8f9 | !hbusreq6_p & v3766c97;
assign v37337b3 = hbusreq0 & v37269de | !hbusreq0 & v3a58c2f;
assign v3a6f342 = hbusreq3_p & v37390ed | !hbusreq3_p & v3a6f95f;
assign v3729949 = hbusreq5_p & v3725371 | !hbusreq5_p & v3726dfd;
assign v3a5880b = hlock0_p & v376ea4a | !hlock0_p & !v3728e09;
assign v3a56df7 = hbusreq4_p & v3732dac | !hbusreq4_p & v3731210;
assign v3764ddc = hmaster0_p & v3a70513 | !hmaster0_p & v372c46e;
assign v38097ee = hmaster2_p & v3a702c2 | !hmaster2_p & v8455b0;
assign v3a7115a = hbusreq0 & v3a70362 | !hbusreq0 & v372e3d8;
assign v3a5f580 = hlock0 & v3733b4e | !hlock0 & v376fc77;
assign v375fbe1 = hbusreq8_p & v372bb25 | !hbusreq8_p & v37494da;
assign v3a6a516 = hmaster2_p & v35772a6 | !hmaster2_p & v375518f;
assign v3a5978c = hbusreq3_p & v3748797 | !hbusreq3_p & v3a6fad9;
assign v37307de = hbusreq0_p & v3a70c07 | !hbusreq0_p & v1e38224;
assign v3a60332 = hmaster0_p & v372cdb8 | !hmaster0_p & v375d4aa;
assign v372d96e = hgrant2_p & v8455ab | !hgrant2_p & v37782ff;
assign v3807969 = hmaster1_p & v3779b9c | !hmaster1_p & v3a70bee;
assign v3769e10 = hmaster1_p & v3748d63 | !hmaster1_p & v8455ab;
assign v375a116 = hgrant6_p & v3771fb3 | !hgrant6_p & v377de92;
assign v3737352 = hbusreq4_p & v3a6f56c | !hbusreq4_p & v3a6ffcc;
assign v375f963 = hmaster0_p & v37559c4 | !hmaster0_p & v374d4d3;
assign v377870b = hbusreq4 & v377d9bb | !hbusreq4 & v3725799;
assign v372ac3b = hbusreq0 & v3a6fb8c | !hbusreq0 & v3754229;
assign v3809f1c = hbusreq3_p & v375a250 | !hbusreq3_p & v376b23a;
assign v3a6b059 = hmastlock_p & v373cb9c | !hmastlock_p & !v8455ab;
assign v37237a8 = hmaster0_p & v8a21c4 | !hmaster0_p & v374e758;
assign v3770362 = hmaster3_p & v3a70dfd | !hmaster3_p & v3a6fb41;
assign v3a6f627 = hbusreq3_p & v3748932 | !hbusreq3_p & v3739417;
assign v3a6162f = hgrant4_p & v3a663b9 | !hgrant4_p & v3733c9e;
assign v3749ec0 = hlock0 & v3765e79 | !hlock0 & v374d80f;
assign v3759032 = locked_p & v8455ab | !locked_p & !v39a537f;
assign v375795d = hmaster0_p & v377e6f5 | !hmaster0_p & v373b59f;
assign v8455cf = hlock7_p & v8455ab | !hlock7_p & !v8455ab;
assign v377b3ff = hmaster0_p & v3725bdc | !hmaster0_p & v37744e0;
assign v376c2d6 = hmaster0_p & v3761769 | !hmaster0_p & !v3a70cab;
assign v374184c = hmaster2_p & v3a70374 | !hmaster2_p & v37431ec;
assign v373d5af = hmaster1_p & v372a0ed | !hmaster1_p & v377cb41;
assign v3749008 = hlock4 & v377d1ab | !hlock4 & v37302c5;
assign v373f64f = hbusreq5 & v374490b | !hbusreq5 & v375c7cf;
assign a374cd = hlock5 & v3a6080b | !hlock5 & v3a68904;
assign v3a70913 = hbusreq1_p & v37469db | !hbusreq1_p & !v3a645f6;
assign v374d7dd = hbusreq6_p & v377915c | !hbusreq6_p & c98f7c;
assign v3a586d0 = hbusreq2 & v3a6dc08 | !hbusreq2 & v376648d;
assign v3a5f609 = hlock8 & v373766f | !hlock8 & v3a6fa99;
assign v3741039 = hmaster2_p & v3a61a7f | !hmaster2_p & v3a635ea;
assign v3a7079b = hmaster0_p & v3750746 | !hmaster0_p & v39a4ef6;
assign v376e6ac = hmaster0_p & v377a312 | !hmaster0_p & !v3722caa;
assign v3a57759 = hmaster1_p & v37582a2 | !hmaster1_p & v3a70f10;
assign v374e03d = hgrant0_p & v37487ca | !hgrant0_p & b27f78;
assign v3a6edbe = hmaster2_p & v377dacb | !hmaster2_p & v8455ab;
assign v377435d = jx0_p & v3a6514f | !jx0_p & v373c268;
assign v37501e6 = hbusreq8_p & v3737aee | !hbusreq8_p & v372de63;
assign v3767091 = hmaster1_p & v8455c5 | !hmaster1_p & !v372d9a1;
assign db6de7 = hmaster2_p & v3807a23 | !hmaster2_p & v3a7047c;
assign v3727ce4 = hlock0_p & v3378ef7 | !hlock0_p & v8455ab;
assign v3a70ea1 = hmaster0_p & v3a57bd7 | !hmaster0_p & !v374b68a;
assign v3757684 = hbusreq2_p & v375a08b | !hbusreq2_p & !v3a68591;
assign v374beee = hbusreq5_p & v3723923 | !hbusreq5_p & v3729308;
assign v3a56ffa = hbusreq5_p & v377de7f | !hbusreq5_p & v3735e52;
assign v3a53d1e = hgrant4_p & v3a6faeb | !hgrant4_p & !v374a580;
assign v3752933 = hlock6 & v3733dd8 | !hlock6 & v3a70466;
assign v3a59ff7 = hgrant6_p & v3744142 | !hgrant6_p & v3a70bf5;
assign v376e4da = hgrant2_p & v3730e2e | !hgrant2_p & d22727;
assign v372dc34 = hbusreq8_p & v374e455 | !hbusreq8_p & v3a70485;
assign v3a6c1ec = hlock6 & v3a715ae | !hlock6 & v372c903;
assign v3a6ebc3 = hbusreq4_p & v3a7115a | !hbusreq4_p & v3a5b57a;
assign v37649e9 = hmaster1_p & v8455ab | !hmaster1_p & v37637d4;
assign v3758395 = hmaster2_p & v374446c | !hmaster2_p & v376acd5;
assign v375ed19 = hbusreq7 & v37500db | !hbusreq7 & v8455ab;
assign v37441e0 = hbusreq2_p & v37325ad | !hbusreq2_p & v3a70c01;
assign v3a714f6 = hbusreq5_p & cfaa3a | !hbusreq5_p & v375977c;
assign v3a5ee62 = hbusreq4_p & v3773f83 | !hbusreq4_p & v37767cd;
assign v3723296 = hlock4_p & v376e914 | !hlock4_p & !v3a658bf;
assign v377cdf0 = hgrant6_p & v8455ab | !hgrant6_p & v373fbc9;
assign v3a6fa8b = hbusreq5_p & v3809505 | !hbusreq5_p & v3a6727a;
assign v2619ae8 = hlock0_p & v95d97e | !hlock0_p & v8455ab;
assign v376ed63 = hmaster0_p & v3806a78 | !hmaster0_p & v8455ab;
assign v3731476 = hmaster1_p & v3a6fb28 | !hmaster1_p & v2ff87d3;
assign v3a5be3f = hbusreq8 & v3a70819 | !hbusreq8 & v373bfdd;
assign v377970b = hbusreq0 & v3a6f09a | !hbusreq0 & v3723e77;
assign v3a6d37f = hgrant3_p & v3759512 | !hgrant3_p & v3a70654;
assign v3749c2f = hmaster2_p & v3a703de | !hmaster2_p & !v373b5f0;
assign v3a70e02 = hlock2_p & v373fcf4 | !hlock2_p & v3a713c7;
assign v377f0fb = hlock8_p & v3771820 | !hlock8_p & v8455b7;
assign v374d4c1 = hgrant0_p & v3779ea0 | !hgrant0_p & v377aad8;
assign v375d6e8 = hlock0 & v3770234 | !hlock0 & v3748d1f;
assign v3733641 = hbusreq5_p & v3a6eede | !hbusreq5_p & !v3a6196d;
assign v3745871 = hmaster0_p & v372de68 | !hmaster0_p & v374e1dc;
assign v37539cd = hmaster2_p & v376d856 | !hmaster2_p & v3728e09;
assign v373547f = hlock5 & v376a052 | !hlock5 & v972988;
assign v374f658 = hgrant4_p & v375cdee | !hgrant4_p & v376e65d;
assign v37315d5 = hgrant2_p & v372919a | !hgrant2_p & v3a70976;
assign v35b724d = hbusreq0 & v3a6f2cf | !hbusreq0 & v3758418;
assign v37534da = hmaster0_p & v3a66835 | !hmaster0_p & !v3a610a4;
assign v373d737 = hbusreq4_p & v380919d | !hbusreq4_p & v3758c32;
assign v3a70809 = hgrant4_p & v372b77b | !hgrant4_p & v3765758;
assign v374ed0a = hlock6 & v3748797 | !hlock6 & v37391a1;
assign v1e37d8b = hbusreq4_p & v3733fad | !hbusreq4_p & v3806f70;
assign v373c04a = hmaster0_p & v3a71243 | !hmaster0_p & v37286e9;
assign v374fa4d = hgrant6_p & v8455ca | !hgrant6_p & v37316fd;
assign v3a6f6c6 = hbusreq2_p & v3a6a4d4 | !hbusreq2_p & v3731906;
assign v3a6a259 = hgrant0_p & v3757568 | !hgrant0_p & v3a66151;
assign v8c5d6a = hbusreq8 & v3a57be6 | !hbusreq8 & v375adcd;
assign cbfab3 = hbusreq5_p & v377e355 | !hbusreq5_p & v37c36bf;
assign v375492b = hbusreq6 & v3749149 | !hbusreq6 & v3a6da8a;
assign v3a29803 = hbusreq1 & v3a54c77 | !hbusreq1 & v377ba55;
assign v871244 = hbusreq0 & v3753fea | !hbusreq0 & v8455ab;
assign v8d2bbf = hbusreq5 & v374fad8 | !hbusreq5 & !v3755a96;
assign v372f09a = hbusreq2_p & v3743dfc | !hbusreq2_p & v373ab4a;
assign v3779a3c = hbusreq5_p & v3752ab6 | !hbusreq5_p & v3756f9b;
assign v3a6f1e2 = hmaster2_p & v3a7127f | !hmaster2_p & !v3a5f83e;
assign v3a6f3e7 = hgrant4_p & v3745f9b | !hgrant4_p & v3770234;
assign v373f42a = hbusreq3_p & v3a6dc32 | !hbusreq3_p & v373421c;
assign v377cbcb = hgrant2_p & v375d12e | !hgrant2_p & v37629e2;
assign v37353d9 = stateA1_p & v8455ab | !stateA1_p & v3a635ea;
assign v37471e0 = hgrant2_p & v3a6c33a | !hgrant2_p & !v3a6b908;
assign v3731c7b = hmaster2_p & v377097a | !hmaster2_p & v3a5e544;
assign v3725f02 = hbusreq2_p & v377773f | !hbusreq2_p & v3763acf;
assign v37579a9 = hbusreq3_p & v3740140 | !hbusreq3_p & !v37761b6;
assign bc7f17 = hgrant0_p & v3a6f43e | !hgrant0_p & v3a70bce;
assign v3a68601 = hbusreq4 & v3a6a493 | !hbusreq4 & v3757f45;
assign v375b2fe = hgrant2_p & v3762502 | !hgrant2_p & v3a5b2fd;
assign v23fde7c = hbusreq4_p & v3749fd7 | !hbusreq4_p & v3a5c2d7;
assign v377022e = hgrant3_p & v375c7b9 | !hgrant3_p & v3a70e23;
assign v376a8cf = hbusreq1_p & v38071c1 | !hbusreq1_p & !v373dc2f;
assign v375bd8c = hmaster2_p & v374449e | !hmaster2_p & v3a57118;
assign v37509a3 = hgrant6_p & v8455c9 | !hgrant6_p & v3a60c05;
assign v3757a04 = hbusreq5_p & v37711f0 | !hbusreq5_p & v3a707b2;
assign v37605db = hbusreq8 & v3a708f9 | !hbusreq8 & v3a5d33e;
assign v3a65c81 = hmaster1_p & v377a968 | !hmaster1_p & v8455ab;
assign v39ebad8 = hbusreq7_p & v990999 | !hbusreq7_p & v3a5b6a3;
assign v3779fd2 = hbusreq5_p & v360d10b | !hbusreq5_p & v3a5dbd7;
assign v3767b98 = hbusreq6_p & v37461e1 | !hbusreq6_p & v3757fde;
assign v376502e = hmaster0_p & v3a635ea | !hmaster0_p & v374bfa6;
assign v38095ed = hbusreq2_p & v3a6fb2a | !hbusreq2_p & v35772a6;
assign v374e314 = hgrant6_p & v374fb58 | !hgrant6_p & v375fd38;
assign v3a70528 = hmaster0_p & v3a683c1 | !hmaster0_p & v3736184;
assign v375c861 = hmaster1_p & v374c73d | !hmaster1_p & v8455ab;
assign v3a68c19 = hgrant2_p & v8455ba | !hgrant2_p & v3a6f98c;
assign v3730b62 = hgrant3_p & v8455bd | !hgrant3_p & v3a56866;
assign v3a6fb6a = hbusreq8 & v3763105 | !hbusreq8 & v373abcf;
assign v3730ba6 = hbusreq6_p & v3a70209 | !hbusreq6_p & v8455ab;
assign v3770a83 = hgrant5_p & v372e47b | !hgrant5_p & v3751a0d;
assign v3745181 = hgrant4_p & v37733c0 | !hgrant4_p & !v3a6f6d3;
assign v37496c6 = hbusreq7_p & v3a704eb | !hbusreq7_p & !v8455ab;
assign v3762a9f = hgrant4_p & v372642c | !hgrant4_p & v375c845;
assign v3a5f991 = hbusreq2 & v3a63805 | !hbusreq2 & v8455b0;
assign v3752552 = hbusreq7_p & v37471c2 | !hbusreq7_p & v3a5e998;
assign v3a7110f = hbusreq8 & v374f8a5 | !hbusreq8 & !v8455ab;
assign v3a5c93e = hmaster0_p & v3a6fa7a | !hmaster0_p & v3a61cb5;
assign v3739635 = hgrant6_p & v8455ab | !hgrant6_p & v3a6bada;
assign v3762db6 = hmaster1_p & v3751a94 | !hmaster1_p & v3a6f54b;
assign v373453a = hbusreq0_p & v3769ae2 | !hbusreq0_p & v375a135;
assign v37391e5 = hgrant5_p & v8455ab | !hgrant5_p & v375acae;
assign v3a6ca53 = hbusreq2_p & v3737c2f | !hbusreq2_p & v2acae91;
assign v3a648c8 = hmaster1_p & v37359cb | !hmaster1_p & v3a6fd9b;
assign v3743425 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3a704d0;
assign v37450aa = hlock5_p & v3a667ba | !hlock5_p & v373f940;
assign v377b3bd = hlock5 & v376e979 | !hlock5 & v3a6ed2b;
assign v37739c7 = hburst0 & v3a6ffa9 | !hburst0 & v8455ab;
assign v376f250 = hbusreq8_p & v3764257 | !hbusreq8_p & v3a636d2;
assign v3733343 = hgrant4_p & v3809400 | !hgrant4_p & !v3a7146f;
assign v3770b24 = hbusreq7_p & v374e00b | !hbusreq7_p & v3726654;
assign v3a6c2d2 = hmaster1_p & v380974c | !hmaster1_p & v37640ff;
assign v375a234 = hgrant6_p & v3728d84 | !hgrant6_p & v3769c2e;
assign v3a6ac33 = hmaster0_p & v2093083 | !hmaster0_p & v373d43a;
assign v23fd8cb = hbusreq0 & v373dd4a | !hbusreq0 & v376a0fc;
assign v3727740 = hbusreq0_p & v3756bc9 | !hbusreq0_p & v3a6d684;
assign v3a70980 = hmaster0_p & v374571a | !hmaster0_p & v376e056;
assign v3a6fdce = hbusreq7_p & v372a1bd | !hbusreq7_p & !v23fd8b7;
assign v35b71da = hmaster2_p & v8455ab | !hmaster2_p & v377db81;
assign v3a6f48b = hbusreq1_p & v39eb57c | !hbusreq1_p & !v8455ab;
assign v376f980 = hbusreq5 & v3a5c511 | !hbusreq5 & v8455ab;
assign v373bff4 = hgrant3_p & v35b774b | !hgrant3_p & v376ed91;
assign v3a6fc98 = hmaster1_p & v8455ab | !hmaster1_p & v3a71329;
assign v374b7e8 = hmaster0_p & v37469c4 | !hmaster0_p & v3771160;
assign v3a710c5 = hbusreq5_p & v375c7cf | !hbusreq5_p & v376a04d;
assign v377c9b3 = hmaster1_p & v8455c1 | !hmaster1_p & v3a6903e;
assign v3a5b23c = hmaster0_p & v373de18 | !hmaster0_p & !v377f34a;
assign v3a7018d = hbusreq7 & v37776eb | !hbusreq7 & v3a6cf44;
assign v375135a = hgrant2_p & v8455e7 | !hgrant2_p & !v3a5eaa1;
assign v372b5f5 = hlock3_p & v3a6fa39 | !hlock3_p & !v8455ab;
assign v377722d = hgrant6_p & v372a51d | !hgrant6_p & v374a7f0;
assign v37363ae = hmaster0_p & v372e959 | !hmaster0_p & v372d51c;
assign a29a96 = hgrant3_p & v8455ab | !hgrant3_p & v37533ac;
assign v372b2aa = hbusreq0 & v3760f4e | !hbusreq0 & v373e814;
assign v37764f7 = hmaster2_p & v8455ab | !hmaster2_p & !v373c991;
assign v37494a7 = hbusreq7 & v372f56c | !hbusreq7 & v374d617;
assign v37297d0 = hgrant4_p & v8455e7 | !hgrant4_p & !v3a7106d;
assign v3770cb8 = hmaster2_p & v3a5f1d4 | !hmaster2_p & v3a5bb64;
assign v3760a1c = hgrant4_p & v8455ab | !hgrant4_p & v37522e4;
assign v3756ca5 = hgrant3_p & v3a6f43e | !hgrant3_p & bc7f17;
assign v374cc43 = hbusreq7 & v3a6f945 | !hbusreq7 & v3a29814;
assign v3773076 = hbusreq7 & v8455b0 | !hbusreq7 & v3724488;
assign v3a7047b = hmaster1_p & v3a6f1a6 | !hmaster1_p & v3a299f8;
assign v3a70498 = hlock8_p & v3a6ec83 | !hlock8_p & v35772a6;
assign v3a65680 = hlock5 & v3761e45 | !hlock5 & v3a71196;
assign v3a6c8b4 = hgrant4_p & v3a6c97d | !hgrant4_p & v375581b;
assign v3a7050f = hbusreq7_p & v37336b4 | !hbusreq7_p & v37523f8;
assign v3a5b78f = hmaster3_p & v3809e77 | !hmaster3_p & v3a6fd1c;
assign v3a53b76 = hlock5_p & v3775303 | !hlock5_p & v3776135;
assign v37275ef = hgrant3_p & v375b3af | !hgrant3_p & v372b9c6;
assign v3a6854c = hbusreq4_p & v3a585d1 | !hbusreq4_p & !v8455ab;
assign v3a702dd = jx3_p & v376726e | !jx3_p & v3809e41;
assign v3737c1c = hbusreq7 & v3a65160 | !hbusreq7 & v3762396;
assign v377d1a3 = hbusreq4_p & v3739b80 | !hbusreq4_p & v3765627;
assign v3734397 = hbusreq7_p & v3767902 | !hbusreq7_p & !v8455ab;
assign v3a6fb38 = hlock8_p & v372a352 | !hlock8_p & v374fcac;
assign v372c5e4 = hbusreq0 & v3a55fc6 | !hbusreq0 & v373f647;
assign v3a5d994 = hmaster2_p & v37566b2 | !hmaster2_p & !v374cab9;
assign v3a6f4af = hlock4 & v3a6e793 | !hlock4 & v3754b2c;
assign v37690da = hmaster0_p & v3a635ea | !hmaster0_p & v372a683;
assign v377d414 = hmaster3_p & v374cf44 | !hmaster3_p & v37422af;
assign v3a5f0cf = hlock0_p & v3a5600a | !hlock0_p & v8455b0;
assign v376aa62 = hbusreq7 & v3772c08 | !hbusreq7 & v3765e47;
assign v3a60691 = hmaster0_p & v3a70a79 | !hmaster0_p & v3a6f53a;
assign v3a60e78 = hbusreq7 & v373d5af | !hbusreq7 & !v3767baa;
assign v377997f = hmaster0_p & v3a5e784 | !hmaster0_p & v373ef01;
assign v3a67403 = hlock0_p & v3a62826 | !hlock0_p & v372d65f;
assign v3744887 = hbusreq5 & v374b3b5 | !hbusreq5 & v8455ab;
assign v376d62b = hbusreq6 & v3a703d0 | !hbusreq6 & v3744f0d;
assign v37706a7 = hbusreq0 & v3a6f323 | !hbusreq0 & v3777e0e;
assign v3750547 = hbusreq2 & v37415b2 | !hbusreq2 & v3a6a393;
assign v3a5e9e9 = hbusreq5 & v1e37a06 | !hbusreq5 & v8455bf;
assign a2e8c8 = hbusreq6_p & v3a7033b | !hbusreq6_p & v8455ab;
assign v3723a94 = hmaster1_p & v375add1 | !hmaster1_p & v3a6f2ce;
assign v3a63624 = hmaster0_p & v3a61bac | !hmaster0_p & !v3755914;
assign v3776311 = jx0_p & v3a67251 | !jx0_p & v3a6f144;
assign v3a7159a = hbusreq4_p & v377e2a4 | !hbusreq4_p & v8455ab;
assign v3743fc1 = hmaster0_p & v3747fda | !hmaster0_p & v3a6f90c;
assign v37705d1 = hgrant3_p & v3770f46 | !hgrant3_p & v375825a;
assign v37389d5 = hbusreq4_p & v3764978 | !hbusreq4_p & v376ecc8;
assign v376ce15 = hbusreq4 & v3a6f2e7 | !hbusreq4 & !v8455ab;
assign v377bc9f = hbusreq8 & v372a965 | !hbusreq8 & v37476d9;
assign v376e0b5 = hmaster2_p & v3755791 | !hmaster2_p & v8455ab;
assign v372f99a = hmaster1_p & v3739c66 | !hmaster1_p & v3a6fef5;
assign v3a647b8 = hbusreq5_p & v376f980 | !hbusreq5_p & v8455ab;
assign v3a64320 = hmaster2_p & v3757966 | !hmaster2_p & v376fbfe;
assign v3765798 = hbusreq0_p & v373b31d | !hbusreq0_p & v376bbe8;
assign v3a6fc74 = hgrant4_p & v8455c1 | !hgrant4_p & v3731511;
assign v39ebb49 = stateA1_p & v8455ab | !stateA1_p & !v3777191;
assign v375faac = hgrant5_p & v3a674e2 | !hgrant5_p & v3a7132e;
assign v3a5aa93 = hgrant5_p & v3a71264 | !hgrant5_p & v3806c70;
assign v3a6eba0 = hlock0 & v3a635ea | !hlock0 & v374733b;
assign v3a6c7ab = hbusreq0 & v37678fc | !hbusreq0 & v373e814;
assign v3a70e80 = hmaster1_p & v3775303 | !hmaster1_p & v372a599;
assign v3a66e3d = hmaster1_p & v3727d4c | !hmaster1_p & v373e30f;
assign v3742dae = hbusreq6_p & v37369eb | !hbusreq6_p & v375d0cf;
assign v3a5fdc8 = hmaster1_p & v377e5e1 | !hmaster1_p & !v8455ab;
assign v3a6a831 = hlock2_p & v375eb97 | !hlock2_p & v3725092;
assign v3a6fac1 = hlock5 & v3a6c1f1 | !hlock5 & v3756fbd;
assign v372d9ad = hbusreq4 & acc1e3 | !hbusreq4 & v3a5a807;
assign v375e147 = hmaster3_p & v373b287 | !hmaster3_p & !v375ff1e;
assign v37603f4 = hgrant1_p & v3733e9e | !hgrant1_p & v3a70c07;
assign v376d45e = hbusreq6_p & v376dcd0 | !hbusreq6_p & !v8455ab;
assign a72315 = hbusreq6_p & v374faa9 | !hbusreq6_p & v3727db9;
assign v37617dd = hmaster2_p & v3757966 | !hmaster2_p & v37480f1;
assign v3a6f7c0 = hlock0_p & v3a5b563 | !hlock0_p & v377af64;
assign v3a5b9ba = hlock1_p & v35772b3 | !hlock1_p & v35772a6;
assign v3a6fc2e = hlock0_p & b254e2 | !hlock0_p & v3739c05;
assign v37390ca = jx0_p & v3773341 | !jx0_p & v3773796;
assign v3a55b39 = hbusreq5_p & v3730055 | !hbusreq5_p & v3a6f831;
assign v37525c8 = hbusreq5 & v3a6f5cb | !hbusreq5 & v377234d;
assign v372f0bb = hbusreq5 & v377a6fe | !hbusreq5 & v8455ab;
assign v374ee47 = stateA1_p & v3a5b585 | !stateA1_p & v3a65206;
assign v373b589 = hbusreq6_p & v3740171 | !hbusreq6_p & v37270d9;
assign v3768a88 = hbusreq2_p & v3a645d7 | !hbusreq2_p & v8455b0;
assign v2aca396 = decide_p & v376b8e1 | !decide_p & v374f0bb;
assign v3a70fb2 = hbusreq2_p & v3a707ad | !hbusreq2_p & v8455ab;
assign v372794f = hbusreq5_p & c17a4a | !hbusreq5_p & v8455ab;
assign v374d643 = hgrant5_p & v373f6b1 | !hgrant5_p & v373419f;
assign v3760d54 = hmaster2_p & v8455ab | !hmaster2_p & v374cd51;
assign v3a65174 = hmaster2_p & v3760a58 | !hmaster2_p & v377234d;
assign v3a6bbeb = hbusreq6_p & v372f1a0 | !hbusreq6_p & v3a5d5cc;
assign v3a64147 = hmaster2_p & v376a6f1 | !hmaster2_p & !v3755793;
assign v3749435 = hlock0_p & v3a7042b | !hlock0_p & v3a69487;
assign v3a5d32a = hmaster2_p & v376b11e | !hmaster2_p & v376bb26;
assign v37729c7 = hbusreq6_p & v374d2b3 | !hbusreq6_p & v3a703d3;
assign v3749b09 = hbusreq4_p & v37536c3 | !hbusreq4_p & v3a6708c;
assign v37701a0 = hmaster2_p & v3744ada | !hmaster2_p & v373f2b6;
assign v3750e9a = hgrant0_p & v373aa23 | !hgrant0_p & v375024d;
assign v3724e61 = hbusreq3 & v3a6ab5f | !hbusreq3 & !v3a6ee22;
assign v373a9db = hmaster3_p & v8455ab | !hmaster3_p & v375a59f;
assign v377aaba = hbusreq5_p & v374b393 | !hbusreq5_p & v375058e;
assign v375a7cd = hbusreq3 & v39a537f | !hbusreq3 & v8455ab;
assign v3a7169d = hbusreq5_p & v3749ab1 | !hbusreq5_p & !v8455ab;
assign d6eddf = hlock0 & v3a5f9e6 | !hlock0 & v3a715a8;
assign v37418bf = hmaster0_p & v375121b | !hmaster0_p & v373a54d;
assign v373e5ad = hlock0_p & v377b673 | !hlock0_p & v376a6d6;
assign v376c484 = hbusreq4_p & v3728d5a | !hbusreq4_p & v37247f2;
assign v3a562a7 = hmaster2_p & v3a7142f | !hmaster2_p & v376f903;
assign v375af00 = hbusreq1 & v3a6f018 | !hbusreq1 & !v3740f3d;
assign v375ea58 = hbusreq3 & v8455e7 | !hbusreq3 & v8455ab;
assign v3a70afd = hbusreq8_p & v376e954 | !hbusreq8_p & v372919e;
assign v37455c2 = hbusreq2 & v3731991 | !hbusreq2 & v3a62a6d;
assign v3a61d1f = hmaster0_p & v8455ab | !hmaster0_p & v377e81a;
assign v3a55ea1 = hlock5 & v3731fb9 | !hlock5 & v3747d33;
assign v377a965 = hgrant6_p & v3725fe1 | !hgrant6_p & v3a6f485;
assign v377b4b0 = hgrant5_p & v372a421 | !hgrant5_p & v3730038;
assign v372cab6 = hbusreq4_p & v380956d | !hbusreq4_p & v3a709f8;
assign v380947a = hbusreq0 & v373f924 | !hbusreq0 & v373c65b;
assign v3745d8c = hmaster2_p & v3773262 | !hmaster2_p & v3768aa4;
assign v3a71557 = hbusreq5 & v3755bbf | !hbusreq5 & v8455ab;
assign v3a5d555 = hbusreq2 & v3a58429 | !hbusreq2 & v3736679;
assign v3a5b333 = hbusreq8_p & v375e516 | !hbusreq8_p & v3a6eee3;
assign v3255b27 = hmaster1_p & v37430c6 | !hmaster1_p & v3a6fa5d;
assign v3772b8a = hlock5 & v3a704f0 | !hlock5 & v3771c5f;
assign v3a70df5 = hbusreq8_p & v3a560d9 | !hbusreq8_p & v3763562;
assign v3a5fbb0 = hbusreq6 & v3759c6c | !hbusreq6 & v380730d;
assign v3759d3c = hbusreq0 & v374f559 | !hbusreq0 & v8455ab;
assign v3a6f446 = hbusreq5_p & v37255f6 | !hbusreq5_p & !v374cb21;
assign v3a5a2e2 = hbusreq2 & v3a6d810 | !hbusreq2 & v3a635ea;
assign v3a5fefa = hbusreq0 & v3738937 | !hbusreq0 & v3a6fb83;
assign v377eb00 = hbusreq4 & v3a63ea7 | !hbusreq4 & v8455ab;
assign v3a5a76d = hbusreq2 & v375fa8b | !hbusreq2 & v375c1d1;
assign v3759d9c = hbusreq7_p & v3761702 | !hbusreq7_p & !v3736b3b;
assign v3756a20 = hmaster1_p & v3777c0c | !hmaster1_p & v3a70d99;
assign v37251e7 = hlock6_p & v37453d8 | !hlock6_p & v380974c;
assign v372580e = hgrant4_p & v1e37b99 | !hgrant4_p & v3a594f1;
assign v376575c = hbusreq0 & v3758f94 | !hbusreq0 & v8455ab;
assign v3a5408e = hmaster2_p & v1e38224 | !hmaster2_p & !v3728e09;
assign v375cb14 = hlock4 & v373e6cf | !hlock4 & v3728d72;
assign v372dcc2 = hgrant2_p & v3a5e24e | !hgrant2_p & v3577416;
assign v3750037 = hgrant0_p & v3723b00 | !hgrant0_p & v3730f98;
assign v3755b07 = hmaster2_p & v3a65da7 | !hmaster2_p & v3a7084e;
assign v3a6edf6 = hmaster1_p & v3a70b5b | !hmaster1_p & v37418db;
assign v3a65cfb = hbusreq3 & v376fe30 | !hbusreq3 & v8455ab;
assign v3754a8e = hlock5_p & v376111d | !hlock5_p & v376285a;
assign v3809127 = hbusreq4 & v3a70e03 | !hbusreq4 & v8455ab;
assign v374ea7d = hbusreq5_p & v3a63f9a | !hbusreq5_p & v375f5f0;
assign v3745249 = hmaster1_p & v372be5d | !hmaster1_p & v8455ab;
assign v37741d7 = hbusreq8 & v3743b2f | !hbusreq8 & v3723025;
assign v3735758 = hmaster1_p & v8455ab | !hmaster1_p & v373e04e;
assign v3a61e6a = hmaster1_p & v372f309 | !hmaster1_p & v374f5d6;
assign v377d0e6 = hmaster0_p & v3a54e42 | !hmaster0_p & !v376bae4;
assign v3a70dd3 = hmaster0_p & v372ff54 | !hmaster0_p & v3764a7d;
assign v376be60 = hlock0 & v3a6a934 | !hlock0 & v376d6b2;
assign v3a70f93 = hbusreq5 & v3a6bee8 | !hbusreq5 & v8455ab;
assign v3739849 = hgrant6_p & v8455c9 | !hgrant6_p & v3a714f2;
assign v374183f = hbusreq8 & v3a612fa | !hbusreq8 & v8455ab;
assign v3a6f888 = hmaster2_p & v375b429 | !hmaster2_p & v3a63805;
assign v37734ba = hlock3_p & v3a6ac81 | !hlock3_p & !v8455ab;
assign v3a62a08 = hgrant4_p & v3754b58 | !hgrant4_p & v3a625d8;
assign v373647a = hbusreq5_p & v376ab39 | !hbusreq5_p & v3a705c7;
assign v3725f9b = hbusreq2 & v3a67603 | !hbusreq2 & v3a6741a;
assign v373d0a2 = hmaster1_p & v3724aa0 | !hmaster1_p & !v37629b0;
assign v3a5bffe = hbusreq4_p & v3735e39 | !hbusreq4_p & !v3a6d684;
assign v37714e6 = hgrant0_p & v8455ab | !hgrant0_p & v3a6f316;
assign v3a6f2d2 = hbusreq5_p & v3723ec6 | !hbusreq5_p & v37332fa;
assign v3762dc3 = hmaster0_p & v3768589 | !hmaster0_p & v372abac;
assign v3a702f1 = hbusreq5 & v377b3be | !hbusreq5 & v8455ab;
assign v3a6f964 = hmaster1_p & v3a62a6d | !hmaster1_p & v3759144;
assign v372a786 = hgrant3_p & v3a5f9f2 | !hgrant3_p & v1e3780f;
assign v3744cd7 = hmaster2_p & v375dc01 | !hmaster2_p & v372c029;
assign v3778251 = hlock3 & v3a61668 | !hlock3 & v3736e1d;
assign v3a618b7 = hgrant0_p & v37773a9 | !hgrant0_p & v3760af0;
assign v3731fe4 = hbusreq7 & v3a6f820 | !hbusreq7 & v3777d70;
assign v3a58be6 = hbusreq5 & v3734fc3 | !hbusreq5 & v3a54466;
assign v3a6307d = hgrant8_p & v376f032 | !hgrant8_p & v325c93a;
assign v37581f6 = hgrant5_p & v3a6f37d | !hgrant5_p & v3a6eb4b;
assign v39a4e1f = hmaster0_p & v3a6c922 | !hmaster0_p & v37662e7;
assign v3744c29 = hgrant3_p & v8455ab | !hgrant3_p & v37378ca;
assign v3743d21 = hgrant2_p & v377d4a0 | !hgrant2_p & v3758adb;
assign v376f111 = hmaster2_p & v376a6f1 | !hmaster2_p & v8455c1;
assign v373b719 = hbusreq3 & v37583be | !hbusreq3 & !v8455ab;
assign v3741922 = hmaster2_p & v372650c | !hmaster2_p & !v37634d8;
assign v3a669c6 = hbusreq5 & v374b025 | !hbusreq5 & v374e92a;
assign v3a61901 = hlock6 & v373e3d5 | !hlock6 & v372d7a4;
assign v37705c0 = hbusreq4_p & v3754bb1 | !hbusreq4_p & v373276f;
assign v8455df = hmaster3_p & v8455ab | !hmaster3_p & !v8455ab;
assign v3756ebf = hlock8_p & v3736107 | !hlock8_p & v37695c1;
assign v3734247 = hgrant6_p & v3726bff | !hgrant6_p & v2092b01;
assign v23fdaf1 = jx0_p & v3a5c40b | !jx0_p & v3a5b517;
assign v3736048 = hmaster2_p & v374fb58 | !hmaster2_p & v3726139;
assign v375ff99 = hgrant5_p & v3740052 | !hgrant5_p & v374294c;
assign v3a71518 = hmaster2_p & v375afe9 | !hmaster2_p & v3770bcd;
assign v3a6fb56 = hmaster0_p & v37710fb | !hmaster0_p & !v3764b6e;
assign v3a5d96d = hbusreq5 & v373e475 | !hbusreq5 & v8455ab;
assign v373a373 = hlock8 & v373c617 | !hlock8 & v380909f;
assign v376cebe = hmaster2_p & v3a6f32f | !hmaster2_p & !v372cc25;
assign v3764306 = hmaster0_p & v3774247 | !hmaster0_p & v3a7090f;
assign v3a54580 = hmaster2_p & v3a635ea | !hmaster2_p & v372348c;
assign v3757271 = hbusreq2 & v3a6fd48 | !hbusreq2 & v3a6f6e7;
assign v3a71319 = hgrant6_p & v37725e7 | !hgrant6_p & v38072fb;
assign v3806818 = hlock3_p & v373aea0 | !hlock3_p & v1e37bab;
assign b755d3 = hgrant3_p & v8455ab | !hgrant3_p & v3743eb5;
assign v3806f19 = hbusreq6_p & v23fd967 | !hbusreq6_p & v3a629a6;
assign v377215c = hbusreq5 & v374f7cb | !hbusreq5 & v3a5f587;
assign v3741cd7 = hbusreq2 & v3a6c2d4 | !hbusreq2 & v37731c3;
assign v3745614 = hmaster1_p & v3a5c42c | !hmaster1_p & v3a70e76;
assign v376ef2d = hmaster0_p & v3747b2b | !hmaster0_p & v377b774;
assign v3a708a1 = hbusreq8 & v3751c54 | !hbusreq8 & v377b951;
assign v3725bfb = hbusreq4_p & v3a6a1b4 | !hbusreq4_p & v374b05b;
assign v3a63512 = hmaster0_p & v3a703e4 | !hmaster0_p & !v375f847;
assign v3a6d684 = locked_p & v39ebac7 | !locked_p & v1e38224;
assign v3a6209f = hmaster1_p & v3750ff0 | !hmaster1_p & v3a6fd9b;
assign v3774cd5 = hgrant3_p & v3a67403 | !hgrant3_p & v37256c4;
assign v3740469 = hlock4 & v377564e | !hlock4 & v3a58674;
assign v3a6dddb = hbusreq6_p & v373502e | !hbusreq6_p & v376f345;
assign v1e3778c = hmaster1_p & v3a6b266 | !hmaster1_p & v3729798;
assign v3a71395 = hbusreq6 & v8455b0 | !hbusreq6 & v373f058;
assign a14297 = hmaster0_p & v3748acd | !hmaster0_p & v37614c1;
assign v3a67118 = hlock6_p & v8455ab | !hlock6_p & v3773fdc;
assign v3a6fe48 = hbusreq6_p & v3a6f0a2 | !hbusreq6_p & v3743b9e;
assign v3725804 = hbusreq5 & v3a70c4c | !hbusreq5 & !v3762847;
assign v3a71505 = hmaster2_p & v3752446 | !hmaster2_p & v377167e;
assign v3a709c6 = hburst0 & v39ebac7 | !hburst0 & !v8455e1;
assign v3a61e33 = hmaster2_p & v3a6f942 | !hmaster2_p & v8455ab;
assign v3740c75 = hgrant4_p & v3a702b3 | !hgrant4_p & v3734788;
assign v2ff87d7 = hbusreq8_p & v3759569 | !hbusreq8_p & v3779810;
assign v376652f = hmaster2_p & v374502e | !hmaster2_p & !v372a4c1;
assign v3740890 = hbusreq3_p & v3a70a48 | !hbusreq3_p & v8455ab;
assign v3a713e8 = jx0_p & v37642fa | !jx0_p & v373e5e7;
assign v374d07a = hmaster1_p & v87be38 | !hmaster1_p & v375dc75;
assign v3a5ed4b = hbusreq4_p & v3a68f04 | !hbusreq4_p & v3a6a6eb;
assign v37436e6 = hmaster1_p & v3774937 | !hmaster1_p & v377e406;
assign v3730f6f = hgrant5_p & v3a6b288 | !hgrant5_p & v372cd1f;
assign c39398 = hbusreq0 & v3733df1 | !hbusreq0 & v37721df;
assign v3a6fc18 = hmaster0_p & v8455ab | !hmaster0_p & !v3a57d41;
assign v3a66fd9 = hmaster2_p & v3747302 | !hmaster2_p & v3a6f3c6;
assign v3a6a546 = hgrant4_p & v37617ad | !hgrant4_p & v8455ab;
assign v3724c77 = hbusreq6_p & v3a68bb1 | !hbusreq6_p & v37774e4;
assign v375d800 = hbusreq4_p & v3a708a4 | !hbusreq4_p & v3a63621;
assign v3a711b7 = hbusreq1 & v3740171 | !hbusreq1 & v8455ab;
assign v3a6f36f = hmaster1_p & v2acb06f | !hmaster1_p & v3778628;
assign a740cc = hmaster1_p & v3a6eb67 | !hmaster1_p & v3728435;
assign v3a707ae = hgrant6_p & v377c147 | !hgrant6_p & v3749586;
assign v3a6f6f2 = hlock7 & v375c144 | !hlock7 & v3a6ddc7;
assign v376241e = hbusreq7_p & v3771724 | !hbusreq7_p & v3771319;
assign v37456d2 = hgrant6_p & v8455ab | !hgrant6_p & v3722da3;
assign v3737bb4 = hmaster2_p & v374b8fa | !hmaster2_p & v3a603fc;
assign v375c728 = hlock0 & v3a635ea | !hlock0 & v39eb56c;
assign v3a703e4 = hmaster2_p & v3723da9 | !hmaster2_p & !v376e854;
assign v3778627 = hlock7_p & v37611f5 | !hlock7_p & v3a5e998;
assign v3731906 = hgrant3_p & v3731d69 | !hgrant3_p & v8455ab;
assign v375c439 = hbusreq6 & v3738df9 | !hbusreq6 & v3731004;
assign v3770bd9 = hbusreq3_p & v374a891 | !hbusreq3_p & v3726f97;
assign v3747f46 = hmaster1_p & v3a7101d | !hmaster1_p & v377f640;
assign a85c8e = hbusreq5 & v372c6c4 | !hbusreq5 & v3a550c2;
assign v372bae3 = hmaster2_p & v37476bd | !hmaster2_p & v376bb26;
assign v3745014 = hbusreq2 & v3a6f018 | !hbusreq2 & !v3740f3d;
assign v28896dc = hmaster2_p & v37330dc | !hmaster2_p & v37320ff;
assign v377cb05 = hgrant5_p & v8455ab | !hgrant5_p & v3a6ef7d;
assign v374d1d7 = hlock8_p & v3736958 | !hlock8_p & v3a2a0e9;
assign v377338f = hbusreq4 & v3a6eb1e | !hbusreq4 & v377c6b3;
assign v374aabf = hmaster2_p & v3730ffe | !hmaster2_p & v8455ab;
assign v3a6db03 = hbusreq5_p & v3a70fed | !hbusreq5_p & v3a5b567;
assign v3769bb0 = hlock7 & v374e828 | !hlock7 & v376f7d1;
assign v376be50 = hbusreq0 & v3a7148e | !hbusreq0 & v3a65aba;
assign v377cccb = hmaster2_p & v376f0fb | !hmaster2_p & v3a6a295;
assign v375ac26 = hbusreq5_p & v3a5ec50 | !hbusreq5_p & v376e5de;
assign v3a6f49b = jx1_p & v374c9e1 | !jx1_p & v3745e63;
assign v37617d8 = hbusreq7_p & v3808d2f | !hbusreq7_p & !v8455ab;
assign v3768e0e = hmaster0_p & v375b5ca | !hmaster0_p & v8455ab;
assign v37707db = hbusreq5 & v3a703aa | !hbusreq5 & v1e379c4;
assign v3a5ab24 = hbusreq8 & v375c009 | !hbusreq8 & v8455c3;
assign v3748eaa = hmaster1_p & v3a71678 | !hmaster1_p & v3a5a381;
assign v3a59178 = hgrant4_p & v3731bc8 | !hgrant4_p & v3733734;
assign v3a5bda4 = hbusreq5 & v37356ec | !hbusreq5 & v8455ab;
assign v372c3b9 = hlock0 & v38072fd | !hlock0 & v3a703cd;
assign v8a21c4 = hmaster2_p & v372d203 | !hmaster2_p & v3a6f0f6;
assign v375d9f8 = hlock0_p & v8455ab | !hlock0_p & v373fe5e;
assign v3a6f76a = hlock5_p & v8455ab | !hlock5_p & v3a6fce0;
assign v3762656 = hbusreq4 & v376f23f | !hbusreq4 & v372348c;
assign v377286e = hlock2_p & v3773ee6 | !hlock2_p & v8455b3;
assign v3776cce = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3a635f8;
assign v3a70b00 = hlock0 & v3775999 | !hlock0 & v3751db5;
assign v3769101 = hmaster2_p & v375ecd5 | !hmaster2_p & v8455ab;
assign v377915c = hgrant2_p & v3a5f50e | !hgrant2_p & d0b9d7;
assign v375a688 = hbusreq5 & v3743792 | !hbusreq5 & v8455ab;
assign v37375ee = hbusreq4_p & v375444e | !hbusreq4_p & v373b3fb;
assign v375d455 = hmaster0_p & v3a5998b | !hmaster0_p & v3744cd7;
assign v2acafdf = hgrant6_p & v375f2ec | !hgrant6_p & v23fe10f;
assign v3a67bce = hmaster0_p & v37247cf | !hmaster0_p & v3729793;
assign v374362e = locked_p & v3755019 | !locked_p & v39a537f;
assign v3770ffb = hbusreq8 & v3a5a48f | !hbusreq8 & v373340f;
assign v37549cd = hmaster0_p & v3773fdc | !hmaster0_p & bbba6b;
assign v3761fd7 = hbusreq5 & v375818b | !hbusreq5 & v8455ab;
assign v377904f = hmaster2_p & v372ee06 | !hmaster2_p & v3776b2a;
assign v37612d4 = hlock0 & v3752767 | !hlock0 & b95629;
assign v375ecc7 = hbusreq0_p & v3a70131 | !hbusreq0_p & v376b4e1;
assign v37681ed = hbusreq4 & v375e0e3 | !hbusreq4 & v3a6f3c6;
assign v3763398 = hgrant6_p & v3a57b60 | !hgrant6_p & v39eb4d4;
assign v3742b31 = hlock3 & v376485c | !hlock3 & v3a5a3be;
assign v3728f6d = hmaster0_p & v3763550 | !hmaster0_p & v3807a26;
assign v375df25 = hbusreq2 & v374fd4a | !hbusreq2 & v3a6e3bb;
assign v3728ac4 = hmaster1_p & v3a70b19 | !hmaster1_p & !v8455ab;
assign v3a70488 = hbusreq0 & v3a6f35f | !hbusreq0 & v3a64af7;
assign v3752a43 = hmaster0_p & v3a5c473 | !hmaster0_p & v3774878;
assign v3a6ec0d = hlock1_p & v3759e9d | !hlock1_p & !v8455ab;
assign v3a6fe83 = hbusreq5_p & v3a6f45c | !hbusreq5_p & v3738844;
assign v3a70f1e = hbusreq5_p & v3769d07 | !hbusreq5_p & !v3765e5b;
assign v373c23c = hbusreq5_p & v372a80a | !hbusreq5_p & v37753b4;
assign v3a6fc1c = hmaster0_p & v8455ab | !hmaster0_p & v376cfd9;
assign v3a70e36 = hgrant3_p & v3774550 | !hgrant3_p & v3725f48;
assign v376cc8d = hbusreq2 & v3728cfe | !hbusreq2 & v3a5f5bb;
assign v3a6fb24 = hmaster1_p & v376e72d | !hmaster1_p & v373f012;
assign v37670ac = hmaster2_p & v377a876 | !hmaster2_p & v3757684;
assign v3a573d2 = hlock5 & v3a63f9a | !hlock5 & v3724547;
assign v3725ccb = hbusreq3_p & v3a551d6 | !hbusreq3_p & v3a5cd20;
assign jx1 = v357748a;
assign v3a5aaed = hbusreq4_p & v3756de3 | !hbusreq4_p & v3a6c2a9;
assign v3a565ef = hlock0_p & v3a637dd | !hlock0_p & !v374b962;
assign v3a71526 = hgrant4_p & v377d58d | !hgrant4_p & v373d12a;
assign v3a70b63 = hmaster2_p & v375cf36 | !hmaster2_p & v3a70c74;
assign v374132e = hbusreq8 & v37751b4 | !hbusreq8 & v3779749;
assign v3a6ef23 = hgrant2_p & v3a70ee7 | !hgrant2_p & v3758dfe;
assign v3a6edb9 = hlock2 & v3742cfe | !hlock2 & v23fdf85;
assign v372ce8b = hbusreq2 & v37482f8 | !hbusreq2 & !v377c3a1;
assign v3a6fd15 = hgrant2_p & v8455ab | !hgrant2_p & v37722c6;
assign v3739d88 = hbusreq6_p & v3255a16 | !hbusreq6_p & v8455ab;
assign v3a69544 = hbusreq2_p & v3a6eead | !hbusreq2_p & v3a5bb64;
assign v372391f = hbusreq1_p & v37502b7 | !hbusreq1_p & v3735e39;
assign v3a5b41c = hgrant2_p & v8df61b | !hgrant2_p & v374c4bc;
assign v372f55a = hmaster1_p & v99797a | !hmaster1_p & v3a596df;
assign v3a6f871 = hmaster2_p & v375e2bc | !hmaster2_p & v35b71cf;
assign v374ee8d = hlock0 & v3a6fdef | !hlock0 & v376d902;
assign v377456d = hlock8 & v3771c6a | !hlock8 & v3a6f92d;
assign v1e37e29 = hmaster0_p & v1e37d3a | !hmaster0_p & v3a5fc34;
assign v372953c = hbusreq7_p & v373501a | !hbusreq7_p & !v3a6efb7;
assign v37673fe = hmaster2_p & v3759c1f | !hmaster2_p & v3739b4c;
assign v3a6aba6 = hbusreq7_p & v3a6cc28 | !hbusreq7_p & v37441dc;
assign v3778395 = hmaster2_p & v372eaaf | !hmaster2_p & v8455e7;
assign v3757264 = hbusreq3_p & v3a7037c | !hbusreq3_p & v3746f84;
assign v376af81 = hlock8_p & v3a581fb | !hlock8_p & v3a6d8a9;
assign v3a6fd27 = hbusreq2_p & v37647aa | !hbusreq2_p & v37673dd;
assign v375c7d3 = hlock0_p & v377eb9d | !hlock0_p & v8455b0;
assign v372b7fb = hmastlock_p & v3a6e431 | !hmastlock_p & v8455ab;
assign v3a62d54 = hbusreq2 & v3a6ab8d | !hbusreq2 & v3769de7;
assign v3a5907a = hbusreq4 & v3763175 | !hbusreq4 & v8455ab;
assign v3735c84 = hlock5 & v3a6fbdb | !hlock5 & v3740681;
assign v3a6de60 = hmaster1_p & v377316f | !hmaster1_p & v3a62424;
assign v3a6f7a0 = hgrant2_p & v8455b9 | !hgrant2_p & v37677d8;
assign v3774e7b = hmaster1_p & v3a61a7f | !hmaster1_p & v3a65680;
assign v2678bee = hbusreq1_p & v8455ab | !hbusreq1_p & v8455eb;
assign v3767a21 = hmaster0_p & v372edf8 | !hmaster0_p & v3774492;
assign v3741e5c = hbusreq4 & v3a5f8d0 | !hbusreq4 & v8455ab;
assign v1e38241 = hgrant6_p & v376d45e | !hgrant6_p & !v8455ab;
assign v3757e40 = hlock8 & v3768737 | !hlock8 & v372586f;
assign v37643e5 = hbusreq0 & v37235f9 | !hbusreq0 & v372ba45;
assign v373c828 = hmaster2_p & v3a5f8d0 | !hmaster2_p & v3749907;
assign v376faad = hgrant0_p & v8455ab | !hgrant0_p & v3a70a68;
assign v3725b27 = hgrant4_p & v8455ab | !hgrant4_p & v3737647;
assign v3a58a0d = hgrant5_p & v372cbac | !hgrant5_p & v373a66b;
assign v372d060 = hmaster0_p & v376c644 | !hmaster0_p & v373f911;
assign v3753576 = hlock5_p & v376f9ca | !hlock5_p & !v3731f3c;
assign v3a710e0 = hgrant5_p & v8455ab | !hgrant5_p & v3a6c322;
assign v377d04f = hmaster0_p & v3a6e5f0 | !hmaster0_p & v3759586;
assign v3733294 = hbusreq5 & v3a70dcb | !hbusreq5 & v3a635ea;
assign v3a71375 = hmaster0_p & v3a635ea | !hmaster0_p & v37c03ad;
assign v3731cf0 = hgrant4_p & v8455ab | !hgrant4_p & v376ae9c;
assign v37480b3 = hmaster0_p & v373bac2 | !hmaster0_p & v3a5fd4a;
assign v3a5842b = hmaster3_p & v373e6d8 | !hmaster3_p & v3a715e8;
assign v3776a6e = hlock0_p & v8455ab | !hlock0_p & v3744710;
assign v3763bb8 = hmaster2_p & v377ed6c | !hmaster2_p & v3a5fbd6;
assign v3753f82 = hlock5_p & v374b9e6 | !hlock5_p & !v3764818;
assign v9e78af = hbusreq5_p & v3a6cc93 | !hbusreq5_p & v375f989;
assign v3a6086a = hready_p & v3760ce0 | !hready_p & v373e02a;
assign v3742c87 = hmaster2_p & v8455ab | !hmaster2_p & v3a58eed;
assign v3777844 = hgrant4_p & v8455ab | !hgrant4_p & v372b5a3;
assign v373b130 = hbusreq5_p & v377de07 | !hbusreq5_p & v3729435;
assign v3a58b04 = hgrant5_p & v3731780 | !hgrant5_p & v3a71057;
assign v3776d3e = hlock8 & v3740ff7 | !hlock8 & v3a6a367;
assign v3a58527 = hmaster0_p & v3a635ea | !hmaster0_p & v372c53a;
assign v3a7099b = hbusreq6_p & v38072fd | !hbusreq6_p & a16ae7;
assign v3a59caa = hmaster2_p & v37385d2 | !hmaster2_p & v3722d9b;
assign v373823e = hbusreq5_p & v3a70134 | !hbusreq5_p & v3a6f387;
assign v3a5706c = hgrant2_p & v8455ab | !hgrant2_p & v3a66668;
assign v3740614 = hbusreq5 & v374f307 | !hbusreq5 & v3a58c07;
assign v377308e = hbusreq4_p & v374e4c0 | !hbusreq4_p & !v8455ab;
assign v37755d5 = hbusreq4_p & v3a6aaaa | !hbusreq4_p & v3a588ec;
assign v3a6f2fd = hmaster1_p & v372ec32 | !hmaster1_p & !v3779003;
assign v3734c20 = hlock6 & v3a54f85 | !hlock6 & v37328fc;
assign v375dcdb = hgrant3_p & v37427cf | !hgrant3_p & !v3a6f36e;
assign v37770ae = hmaster2_p & v3a687be | !hmaster2_p & v3a67967;
assign v3a70ff9 = hgrant3_p & v376e914 | !hgrant3_p & !v37345f3;
assign v377d3b9 = hbusreq4 & v3a55efa | !hbusreq4 & v3735525;
assign v3769950 = hbusreq4_p & v37519e3 | !hbusreq4_p & v8455ab;
assign v375f7d1 = hgrant4_p & v8455ab | !hgrant4_p & v3741ef3;
assign v3a62550 = hgrant6_p & v377f09a | !hgrant6_p & v3a57ad0;
assign v3a5d836 = hgrant2_p & v8455ab | !hgrant2_p & v3a6fe0a;
assign v375aff6 = hmaster0_p & v3763f20 | !hmaster0_p & v373185b;
assign v373c433 = hbusreq7 & v3a70b40 | !hbusreq7 & v8455ab;
assign v3750b61 = hgrant4_p & v3750d06 | !hgrant4_p & v360d07a;
assign d435c2 = hgrant0_p & v37416b5 | !hgrant0_p & v3775bf6;
assign v3731376 = hlock8_p & v3762199 | !hlock8_p & !v8455ab;
assign v3a58fef = stateG10_1_p & v37764a5 | !stateG10_1_p & v373f661;
assign v3a7097c = hmaster2_p & v3a70464 | !hmaster2_p & v374b5c5;
assign v37323a5 = hlock6_p & v3747c3e | !hlock6_p & v8455ab;
assign v3a6e404 = hmaster1_p & v8455ab | !hmaster1_p & v3766014;
assign v3771088 = hmaster1_p & v3a56069 | !hmaster1_p & v375c70a;
assign v3a69f8e = hbusreq5 & v3776ada | !hbusreq5 & v1e3737d;
assign v3762389 = hlock3 & v3a6b8a2 | !hlock3 & v3768062;
assign v3a55584 = hbusreq0 & v372c480 | !hbusreq0 & v3735112;
assign v3726eb4 = hgrant5_p & v37346fe | !hgrant5_p & d383e7;
assign v376993b = hbusreq6_p & v372300f | !hbusreq6_p & v376baef;
assign v3a70ec9 = hbusreq6_p & v3a701d9 | !hbusreq6_p & v8455ab;
assign v374158d = hgrant4_p & v376ac08 | !hgrant4_p & v3a7157e;
assign v3a70351 = hbusreq3_p & v377d393 | !hbusreq3_p & v3a6fee8;
assign v3737a06 = hmaster0_p & v8455ab | !hmaster0_p & v3a6f441;
assign v3a6fa2d = hmaster0_p & v3771076 | !hmaster0_p & v375bf61;
assign v3a5ccab = hlock8_p & v3a5b0ea | !hlock8_p & v8455ab;
assign v3a704e5 = hlock2_p & v3a6fa39 | !hlock2_p & !v8455ab;
assign v3731003 = hmaster1_p & v377d202 | !hmaster1_p & !v3779a66;
assign v373f418 = hbusreq7_p & v3a71442 | !hbusreq7_p & v23fe156;
assign v3379430 = hmaster2_p & v37470c7 | !hmaster2_p & v372ea9b;
assign v3732bc1 = hbusreq2 & v9181c9 | !hbusreq2 & v8455ab;
assign v3a68c1f = locked_p & v8455ab | !locked_p & !v3807bf8;
assign v375d65c = hmaster2_p & v3a6fdef | !hmaster2_p & v3735525;
assign v3a5b213 = hlock0_p & v3a57309 | !hlock0_p & !v8455ab;
assign v3731c2f = hmaster2_p & v3755000 | !hmaster2_p & v377d232;
assign v3a5ef0d = hmaster3_p & v3753f36 | !hmaster3_p & !v3a66e7f;
assign v372fade = hmaster1_p & v374502e | !hmaster1_p & v3748b2c;
assign v3a6c179 = hmaster0_p & v376c198 | !hmaster0_p & v375c621;
assign v374d011 = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3735512;
assign v3a5923e = hmaster0_p & v3a568e8 | !hmaster0_p & v3a6f379;
assign v3727e80 = hmastlock_p & v3732fec | !hmastlock_p & v8455ab;
assign v376c4e8 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3760d46;
assign v377065f = hbusreq8_p & v3773165 | !hbusreq8_p & !v8455ab;
assign v3a7096e = hlock6_p & v37269f4 | !hlock6_p & v374b3cf;
assign v3743bde = hmaster0_p & v37712aa | !hmaster0_p & v3a700db;
assign v3728723 = hmaster3_p & v8455ab | !hmaster3_p & v377e539;
assign v37771cc = hmaster3_p & v374ebac | !hmaster3_p & v374dd5f;
assign v376f858 = hmaster2_p & v380760a | !hmaster2_p & v3a6ca15;
assign v3739ddf = hbusreq6_p & v373691d | !hbusreq6_p & v8455ab;
assign v373cc0c = hmaster3_p & v373539e | !hmaster3_p & v373ea50;
assign v3762a68 = hbusreq8 & v373a832 | !hbusreq8 & v373c183;
assign v3a5463b = hbusreq5_p & v3770690 | !hbusreq5_p & v3a6f4ca;
assign v3759c8c = hbusreq5_p & v372b6bf | !hbusreq5_p & v3a6f360;
assign v3746ae3 = hmaster0_p & v375fe7a | !hmaster0_p & !v8455bb;
assign v3771d70 = hbusreq8 & v3a58e15 | !hbusreq8 & !v3a6eb28;
assign v3a710f1 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3a6fdef;
assign v8455d7 = hburst1_p & v8455ab | !hburst1_p & !v8455ab;
assign v3a6fd81 = hbusreq6 & v3a702c2 | !hbusreq6 & v8455ab;
assign v37396eb = hbusreq3 & v3a54c77 | !hbusreq3 & v377ba55;
assign v2acb0ef = hmaster1_p & v3a69f0e | !hmaster1_p & v377cb41;
assign v377de72 = hbusreq8_p & v3771214 | !hbusreq8_p & v8455ab;
assign v37500e0 = hmaster2_p & v3779060 | !hmaster2_p & v3759b2f;
assign v3723e23 = hbusreq5_p & v3a6fa7c | !hbusreq5_p & v3a66856;
assign v3a5b583 = hgrant2_p & v8455b9 | !hgrant2_p & v3732b12;
assign v3a67f58 = hbusreq5 & v37540dd | !hbusreq5 & v3a5eae2;
assign v3a6a9d3 = hgrant5_p & v3765e47 | !hgrant5_p & v374c2e2;
assign v3a55d41 = hbusreq3_p & v3741cb9 | !hbusreq3_p & v3757663;
assign v376062b = hmaster3_p & v8455ab | !hmaster3_p & v3753445;
assign v3a66aa6 = hmaster0_p & v3a5ad26 | !hmaster0_p & v8d4314;
assign v3a58182 = hmaster0_p & v3734967 | !hmaster0_p & v3a54f8a;
assign v374af6a = hbusreq3 & v373a27c | !hbusreq3 & v8455e7;
assign v3743b2f = hlock7 & v374e873 | !hlock7 & v372fcfc;
assign v3a631f7 = hbusreq8 & v3a705d2 | !hbusreq8 & v3777d70;
assign v3a711d8 = hgrant6_p & v3770c9d | !hgrant6_p & v372a5c8;
assign v377f579 = hmaster0_p & v374f307 | !hmaster0_p & v372b679;
assign v376f3c8 = hlock3 & v3a6ffcf | !hlock3 & v3a6772f;
assign v3756a6f = hmaster2_p & v376158d | !hmaster2_p & v372a1d6;
assign v3736b0e = hmaster1_p & v35b774b | !hmaster1_p & v372b607;
assign v3a704ae = hmaster2_p & v8455ab | !hmaster2_p & !v374be32;
assign v3763a1e = hmaster3_p & v8455ab | !hmaster3_p & v3765f61;
assign v3a70e5a = hbusreq6_p & v3a5b121 | !hbusreq6_p & v2acb056;
assign v37231c2 = hmaster0_p & v8455ab | !hmaster0_p & v3a71635;
assign v98083e = hmaster2_p & v37763d1 | !hmaster2_p & v377d1dc;
assign v337830d = hgrant0_p & v3a635ea | !hgrant0_p & v3772c19;
assign v3a60ac5 = jx1_p & v37298b2 | !jx1_p & v3739983;
assign v3a5878e = hlock5 & v3779a80 | !hlock5 & v3a70dd3;
assign v376ce1a = hbusreq7_p & v375a1fd | !hbusreq7_p & v376323b;
assign v3731549 = hbusreq4 & v3a70987 | !hbusreq4 & v3a5a807;
assign v37682d5 = hmaster0_p & v3774161 | !hmaster0_p & !v3762e85;
assign v3a6f17e = hbusreq6_p & v3739386 | !hbusreq6_p & v3a70ad4;
assign v376dd80 = hmaster3_p & v3a70b12 | !hmaster3_p & v3a6582d;
assign v373bded = hmaster2_p & v3a6f442 | !hmaster2_p & v3a5b51a;
assign bda6d5 = hgrant1_p & v3a68c1f | !hgrant1_p & !v3a700a5;
assign v3766216 = hmaster0_p & v3a6f1e2 | !hmaster0_p & !v376ef9f;
assign v3a6fde5 = hmaster0_p & v3a619c0 | !hmaster0_p & v377224f;
assign v3778e98 = hmaster1_p & v377e7ac | !hmaster1_p & v372fbb1;
assign v3a681f5 = hbusreq7_p & v374237b | !hbusreq7_p & !v3a6ed14;
assign v3725d14 = hbusreq8 & v3a6eb29 | !hbusreq8 & v3775790;
assign v37621eb = hlock4 & v3a64b83 | !hlock4 & v3760a55;
assign v374179c = hlock4_p & v3a58261 | !hlock4_p & !v8455ab;
assign v374602f = hlock5_p & v3731839 | !hlock5_p & v3724733;
assign v3a57cc8 = hmaster0_p & v375cb51 | !hmaster0_p & v3a71202;
assign bd1306 = hbusreq8 & v375f28d | !hbusreq8 & v376fdd4;
assign v3a6f373 = hbusreq0_p & v377d5d7 | !hbusreq0_p & v375cea7;
assign v3a6f548 = jx1_p & v377115c | !jx1_p & v3752986;
assign v37720f9 = hmaster0_p & v3741748 | !hmaster0_p & v372fd0a;
assign v3a7024c = hlock6 & v37233e7 | !hlock6 & v375da9c;
assign v372fdd0 = hmaster1_p & v3a635ea | !hmaster1_p & v3772e85;
assign v3a7026e = jx0_p & v375fe15 | !jx0_p & v37277ab;
assign v3a6a352 = hlock5_p & v8455ab | !hlock5_p & v3a6f8f0;
assign v3a7149d = hgrant4_p & v3772d6e | !hgrant4_p & v375460c;
assign v39ea259 = hgrant5_p & v372450e | !hgrant5_p & v376e2a4;
assign v3a57210 = hgrant7_p & v9bba04 | !hgrant7_p & v37572eb;
assign v3a5874e = hbusreq7 & v3a5def7 | !hbusreq7 & a0a219;
assign v3725036 = hmaster0_p & v8455ab | !hmaster0_p & v3a704ae;
assign v3a7158e = hmaster0_p & v3a6a56e | !hmaster0_p & v3776c95;
assign v3a6ce39 = hgrant4_p & v8455ab | !hgrant4_p & ac1a2c;
assign v3a6a54d = hmaster2_p & v37c048c | !hmaster2_p & v377b038;
assign v372cdd5 = hmaster2_p & v375c4e6 | !hmaster2_p & v3a70e3d;
assign v3a5ada9 = hmaster0_p & v3a5a510 | !hmaster0_p & v373d593;
assign v3733090 = hlock0_p & v8455ab | !hlock0_p & v3a5f20c;
assign v3a7165a = hmaster0_p & v8455b0 | !hmaster0_p & v375ea85;
assign v3a661c2 = hmaster0_p & v3a708ce | !hmaster0_p & !v375449f;
assign v376abd9 = hbusreq5_p & v37536bf | !hbusreq5_p & v3a620f1;
assign v37407b3 = hgrant0_p & v375039e | !hgrant0_p & v3a573e3;
assign v3a70417 = hlock0 & v373b687 | !hlock0 & v3775831;
assign v376b6c9 = hgrant3_p & v8455ab | !hgrant3_p & v3a7078a;
assign v3a698b7 = hbusreq7 & v3765f8e | !hbusreq7 & v8455ab;
assign v373d848 = hgrant2_p & v8455ba | !hgrant2_p & v377d39f;
assign v38073c9 = hgrant6_p & v3a70a88 | !hgrant6_p & v37372c9;
assign v37650bd = hgrant2_p & v3755a0f | !hgrant2_p & v3764994;
assign v374a45c = hbusreq1_p & b4fa3c | !hbusreq1_p & v372b4ba;
assign v92a03a = hlock0 & v3a5741c | !hlock0 & v3723e5d;
assign v372ba0f = hbusreq4 & v377af44 | !hbusreq4 & v8455ab;
assign v3a70710 = hbusreq3_p & v372fbf4 | !hbusreq3_p & !v3727fd0;
assign v37569b8 = hbusreq8_p & d18baa | !hbusreq8_p & v3a6f670;
assign v9edb6a = hlock6_p & v3754e5e | !hlock6_p & v8455ab;
assign v3a6fcc1 = hgrant1_p & v1e37e66 | !hgrant1_p & !v8455ab;
assign v3778f19 = hlock5 & v3a6f3a9 | !hlock5 & v3745790;
assign v37288c3 = jx0_p & v37457a8 | !jx0_p & v3733cf4;
assign v37512f3 = hgrant6_p & v373557c | !hgrant6_p & v3a6dae5;
assign v3759ad8 = hgrant4_p & v3778ed4 | !hgrant4_p & !v8455ab;
assign v377374f = hbusreq0_p & v3a6fe46 | !hbusreq0_p & v8455ab;
assign v3a704c7 = hbusreq6_p & v3a60787 | !hbusreq6_p & v3733d6e;
assign v3a57422 = hmaster2_p & v377e419 | !hmaster2_p & v37747f8;
assign v376015e = hbusreq3_p & v38072fd | !hbusreq3_p & v376efcf;
assign v3773837 = hbusreq3_p & v3a2a770 | !hbusreq3_p & v3751460;
assign v38079db = hbusreq8 & v375c3c5 | !hbusreq8 & v3a6b303;
assign v3762dd5 = hmaster1_p & v375e512 | !hmaster1_p & v372e741;
assign v3a56794 = hlock5 & v3a714c8 | !hlock5 & v372b794;
assign v3a70287 = hbusreq8_p & v3a6cc28 | !hbusreq8_p & v3a6aba6;
assign v372da95 = jx0_p & v3a6fe15 | !jx0_p & v8455ab;
assign v37789da = hlock6 & v373af5d | !hlock6 & v39a5293;
assign v3744abe = hlock5_p & v373449d | !hlock5_p & v3776da7;
assign v3a6a0a6 = hmaster2_p & v374b8fa | !hmaster2_p & v3771a0d;
assign v3a547ff = hbusreq5_p & v375e0cb | !hbusreq5_p & !v1e382e7;
assign v3a60c82 = hmaster0_p & v3769c70 | !hmaster0_p & v37733e3;
assign v375aa44 = hlock7_p & v377d3bf | !hlock7_p & v3a6fec5;
assign v374ea27 = hgrant2_p & v3a5f50e | !hgrant2_p & v377d67a;
assign v372d07b = hmaster1_p & v3a63fe2 | !hmaster1_p & !v372bd2b;
assign v373340d = hbusreq6_p & v3a5dd17 | !hbusreq6_p & v3778528;
assign v375c551 = hbusreq8_p & v377adaa | !hbusreq8_p & v3a7089e;
assign v3a6ef27 = hbusreq8 & v8455b0 | !hbusreq8 & v3a71504;
assign v372f744 = jx0_p & v3a573ec | !jx0_p & v3a6eff6;
assign v3778e28 = hbusreq4_p & v3723da9 | !hbusreq4_p & v3a62a13;
assign v37742f4 = hbusreq8 & v3739681 | !hbusreq8 & v3763ca1;
assign v8455b5 = hbusreq1_p & v8455ab | !hbusreq1_p & !v8455ab;
assign v376cd91 = hbusreq3_p & v2aca977 | !hbusreq3_p & v3748900;
assign v3775725 = hlock0 & v3a5e2e1 | !hlock0 & v37652f1;
assign v3765466 = hmaster2_p & v3a70ee7 | !hmaster2_p & v3a6f312;
assign v35b86d1 = hmaster1_p & v375cf11 | !hmaster1_p & !v377f640;
assign v380700c = hbusreq4 & v3a6fcd3 | !hbusreq4 & !v374c13e;
assign v3a53cf1 = hmaster1_p & v373e474 | !hmaster1_p & v3778333;
assign v3a5c0de = hbusreq2_p & b66740 | !hbusreq2_p & !v2092faa;
assign v3739f1d = hmaster1_p & v373b6ee | !hmaster1_p & v37558f2;
assign bba7f1 = hlock3 & v3a5a985 | !hlock3 & v3a6ca99;
assign v373e5f1 = stateG2_p & v8455ab | !stateG2_p & v3a65db0;
assign v3a533ae = hbusreq2_p & v377ba5a | !hbusreq2_p & v38079d7;
assign v2acaf6f = hbusreq2_p & d0b9d7 | !hbusreq2_p & ae13ec;
assign v37692e3 = hbusreq7 & v3a6f697 | !hbusreq7 & v3a5666f;
assign v372cbfc = hbusreq4 & v375a4fa | !hbusreq4 & !v8455ab;
assign v37229e6 = hbusreq5_p & v373e0d8 | !hbusreq5_p & v373dcdd;
assign v372e91a = hbusreq5_p & v3764219 | !hbusreq5_p & v3740490;
assign v3767cb7 = hbusreq6 & v3a5be20 | !hbusreq6 & v374fc8e;
assign v3a54e42 = hmaster2_p & v376fcc3 | !hmaster2_p & !v372a0b0;
assign v3722e5a = hmaster3_p & v37723fb | !hmaster3_p & v8455db;
assign v376cdf3 = hbusreq0 & v37612dd | !hbusreq0 & v3a6fd9d;
assign v3772dc6 = hbusreq3_p & v3a65546 | !hbusreq3_p & v3728b05;
assign v372bf24 = hbusreq4_p & v377eaf2 | !hbusreq4_p & v3730695;
assign v3a70cb6 = hbusreq6 & v8455b0 | !hbusreq6 & b6390c;
assign v373f07d = hmaster0_p & v37793e4 | !hmaster0_p & v3a70890;
assign v3a70c81 = hlock7_p & v2acb015 | !hlock7_p & v3a69631;
assign v37466d4 = hbusreq4_p & v35772a2 | !hbusreq4_p & v3a70cc3;
assign v3a67eb4 = hgrant5_p & v3a70638 | !hgrant5_p & v373fb1a;
assign v3a6af67 = hlock4 & v3a70728 | !hlock4 & v376dc16;
assign v37449d1 = hbusreq7_p & v3778362 | !hbusreq7_p & v37556c0;
assign v3a6c717 = hgrant6_p & v3739d45 | !hgrant6_p & v3741f3c;
assign v3a6ff1f = hmaster1_p & v3808cf7 | !hmaster1_p & !v373a11f;
assign v3a56518 = hgrant2_p & v3a6cfe0 | !hgrant2_p & v373a101;
assign v380886b = hmaster2_p & v3577306 | !hmaster2_p & v3a5b5d3;
assign v377bb38 = hbusreq5 & v3738e3c | !hbusreq5 & v3a6fa7c;
assign v3a71182 = hmaster2_p & v3a66910 | !hmaster2_p & !v376d86c;
assign v3a6eae6 = hbusreq6 & v375a750 | !hbusreq6 & v3a58dc1;
assign v377faa6 = hbusreq5_p & v3a5b571 | !hbusreq5_p & !v8455ab;
assign c5fc63 = hgrant4_p & v3779717 | !hgrant4_p & v373187a;
assign v3749dc2 = hbusreq7_p & v37249fe | !hbusreq7_p & v3732899;
assign bb611d = hbusreq2 & cee4af | !hbusreq2 & v8455ab;
assign v3775c6e = hmaster2_p & v3a58ddb | !hmaster2_p & v8455ab;
assign v3a6bba5 = hbusreq7 & v3a58b04 | !hbusreq7 & v3a59cce;
assign v37385c6 = hbusreq5 & v374b23d | !hbusreq5 & v3a67b76;
assign v3a6c437 = hlock4_p & v37534a4 | !hlock4_p & v3a62550;
assign v3a703a3 = hbusreq5 & v3a5d2a6 | !hbusreq5 & v373a9a9;
assign v3a5c3d7 = hmaster2_p & v374729b | !hmaster2_p & !v3725f77;
assign aef673 = hgrant2_p & v8455ab | !hgrant2_p & v3a6c2ad;
assign v3729440 = jx0_p & v8455ab | !jx0_p & v376e66e;
assign v375fbe8 = hbusreq2 & v380930a | !hbusreq2 & v3778cdd;
assign v3725dbb = hbusreq8 & v374407c | !hbusreq8 & v3778211;
assign v374e3a9 = hbusreq4 & v3773575 | !hbusreq4 & v3a6f044;
assign b66740 = hlock0_p & v37502b7 | !hlock0_p & v3735e39;
assign v37519e3 = hbusreq4 & v3746b4f | !hbusreq4 & v8455ab;
assign v3a5fdab = hbusreq0_p & v375e657 | !hbusreq0_p & !v3a69591;
assign v3767f7f = hgrant4_p & v8455c1 | !hgrant4_p & v3a705bc;
assign v376bc75 = jx0_p & v3a6e221 | !jx0_p & v3a71150;
assign v37626d5 = hlock4_p & v3766ea9 | !hlock4_p & v3a57309;
assign v3a6fd11 = hgrant6_p & v376f175 | !hgrant6_p & v337897a;
assign v373c1ed = hmaster1_p & v37241db | !hmaster1_p & v374ec37;
assign v373a8d6 = hgrant1_p & v3a69de7 | !hgrant1_p & v3a635ea;
assign v3a6f0f6 = hgrant2_p & v3a5a6f4 | !hgrant2_p & v3778fb2;
assign v3774df9 = hbusreq6 & v3770075 | !hbusreq6 & v372348c;
assign v3a70f35 = hlock7 & v37626b9 | !hlock7 & v374ecf9;
assign v377c0c3 = hmaster1_p & v8455ab | !hmaster1_p & v3a55b5b;
assign v37710d4 = hgrant4_p & v8455ab | !hgrant4_p & v3749e96;
assign v3a6a4b0 = hmaster0_p & v8455ab | !hmaster0_p & v37731d8;
assign v3a712d5 = hbusreq8 & v3a59b6d | !hbusreq8 & v3a67beb;
assign v37789ca = hmaster2_p & v37329ec | !hmaster2_p & v374449e;
assign v377f5e0 = hmaster2_p & v3775b81 | !hmaster2_p & v8455ab;
assign v372b6bf = hmaster0_p & v37342ef | !hmaster0_p & v3a5c94c;
assign v3742938 = hmaster2_p & v3a5e2a3 | !hmaster2_p & !v8455ab;
assign v37279dc = hgrant5_p & v3a5d6e3 | !hgrant5_p & v3a70dfa;
assign v372870d = hlock6_p & v3a6ac26 | !hlock6_p & v8455ab;
assign v3a5cff8 = hmaster0_p & v3776a3e | !hmaster0_p & v372f9cf;
assign v3808eb8 = hgrant5_p & v373b0b2 | !hgrant5_p & v373940c;
assign v37635de = hmaster2_p & v376285a | !hmaster2_p & v8455ab;
assign v3773f83 = hbusreq4 & v373b589 | !hbusreq4 & v8455e7;
assign d0a27e = hbusreq2 & v373b317 | !hbusreq2 & v3737ad2;
assign v37429d9 = hbusreq7_p & v3a5bbc1 | !hbusreq7_p & v373c8bb;
assign v3a7015f = hbusreq6_p & v3a71416 | !hbusreq6_p & !v3a6bc65;
assign v3a5b3dc = hbusreq7 & v37645f6 | !hbusreq7 & v376e66e;
assign v3a621d5 = hbusreq8_p & v3728373 | !hbusreq8_p & v3a6ff04;
assign v3753f1a = locked_p & v3807071 | !locked_p & v8455ab;
assign v3771440 = hlock5 & v374a509 | !hlock5 & v3a70467;
assign v376cf85 = stateG10_1_p & v8455ab | !stateG10_1_p & v372a7c9;
assign v3a6f8ee = hbusreq0 & v3a5bd05 | !hbusreq0 & v3a635ea;
assign v377324f = hbusreq8_p & v376ae69 | !hbusreq8_p & v1e37c44;
assign v373185f = hlock0 & v3752cf6 | !hlock0 & v3a6f52c;
assign v373a588 = hlock4_p & v373580a | !hlock4_p & v3722a7e;
assign aa52b8 = hbusreq0 & v373a196 | !hbusreq0 & v373a305;
assign v3740328 = hmaster1_p & v3a6a478 | !hmaster1_p & !v37229e6;
assign v3a707d0 = hmaster2_p & v3730e98 | !hmaster2_p & v8455ab;
assign v3a5cb92 = hbusreq7 & v3a6ebd0 | !hbusreq7 & v3767b70;
assign v377bf71 = hbusreq0 & v37348ee | !hbusreq0 & v8455ab;
assign v3a59d5f = hgrant4_p & v374409a | !hgrant4_p & v3a706a6;
assign v3a7025c = hmaster3_p & v374fef0 | !hmaster3_p & v37525c5;
assign v3730ffe = hlock3_p & v3a60132 | !hlock3_p & !v8455ab;
assign v373e41c = hmaster0_p & v374502e | !hmaster0_p & v39eb1df;
assign v3765d74 = hgrant4_p & v3a56580 | !hgrant4_p & v3769ad7;
assign v3255a0c = hmaster0_p & v377d1dc | !hmaster0_p & v3a55377;
assign v3728435 = hbusreq5_p & v373e587 | !hbusreq5_p & v376158e;
assign v3759c90 = hlock1 & v3a6b381 | !hlock1 & v3a685cd;
assign v375de7f = hgrant2_p & v3a708c2 | !hgrant2_p & v3757955;
assign v37bfc8b = hmaster2_p & v3a70446 | !hmaster2_p & !v3747400;
assign v3378e07 = hgrant6_p & v8455ab | !hgrant6_p & v374f5e3;
assign v372aa55 = hlock6_p & v3a6f331 | !hlock6_p & v37765fb;
assign v3746acf = hmaster1_p & v376501e | !hmaster1_p & v3a6f772;
assign v3755e66 = hlock7_p & v374aa82 | !hlock7_p & !v8455ab;
assign v374d9fe = hmaster0_p & v374d926 | !hmaster0_p & v373a02b;
assign v3a67acf = hmaster1_p & v3a70484 | !hmaster1_p & v9e6ddd;
assign v3a6772f = hgrant0_p & v8455ab | !hgrant0_p & v3777787;
assign v3772e33 = hgrant2_p & v37320bb | !hgrant2_p & v3a5561b;
assign v3755bc2 = hgrant3_p & v3a68aa8 | !hgrant3_p & v37359d8;
assign v374672f = hbusreq4_p & v3749831 | !hbusreq4_p & d90332;
assign v377163d = hlock4_p & v3a6ac2a | !hlock4_p & v8455ab;
assign v37702dc = hbusreq5_p & v38064d5 | !hbusreq5_p & v3a6f573;
assign v3763863 = hmaster2_p & v372ee7e | !hmaster2_p & !v373e8ad;
assign v3753a2e = hmaster2_p & v3a6ff99 | !hmaster2_p & v37697a3;
assign v3a6e37c = hmaster2_p & v3a66910 | !hmaster2_p & !v375fbbb;
assign v372ee18 = hmaster1_p & v3808d7d | !hmaster1_p & v8455ab;
assign v37627c3 = hgrant4_p & v37436bc | !hgrant4_p & v3739aa6;
assign v373a755 = hbusreq6_p & v374e542 | !hbusreq6_p & v8455ab;
assign v375d3a2 = hgrant4_p & v8455ab | !hgrant4_p & v37285eb;
assign v374dfea = hgrant3_p & v9ed516 | !hgrant3_p & v37775d9;
assign v3a6e985 = hbusreq4_p & v3747302 | !hbusreq4_p & v3a70c35;
assign v372b390 = hmaster2_p & v3a5c85c | !hmaster2_p & v3747a41;
assign v375c099 = hmaster1_p & v37763d1 | !hmaster1_p & v3a68525;
assign v3779e38 = hmaster1_p & v3a6efe8 | !hmaster1_p & v37499a9;
assign v376acf0 = busreq_p & v3a2a766 | !busreq_p & v8455e1;
assign v37780cd = hbusreq6_p & v373142a | !hbusreq6_p & !v3a67221;
assign v3764568 = hgrant4_p & v3771042 | !hgrant4_p & v3767d4b;
assign v3a580a0 = busreq_p & v3a703cf | !busreq_p & v37562fd;
assign v372afda = hbusreq6_p & v3a5a2be | !hbusreq6_p & v3757fde;
assign v37735aa = hbusreq5_p & v373859f | !hbusreq5_p & v375f172;
assign v3a6fba9 = hbusreq4 & v37572f7 | !hbusreq4 & v377c6b3;
assign v8b397d = hlock0_p & v3750d37 | !hlock0_p & v3a5f147;
assign v3722fe6 = hlock5_p & v3a62481 | !hlock5_p & v3737fca;
assign v374bc20 = hbusreq7_p & v3a5fae4 | !hbusreq7_p & !v3a67d49;
assign v375c3a2 = hbusreq4 & v3a6f709 | !hbusreq4 & v375f9df;
assign v37671eb = hlock0 & v374f35a | !hlock0 & v37366ed;
assign v373ebcf = hmaster0_p & v3759a4a | !hmaster0_p & v3a705e6;
assign v374a115 = hbusreq4 & cb1cc0 | !hbusreq4 & v375cf36;
assign v373b6ba = hbusreq5 & v37678bd | !hbusreq5 & v373112c;
assign v37368ce = hgrant4_p & v372b77b | !hgrant4_p & v377a9cb;
assign v373faf3 = hmaster3_p & v377f037 | !hmaster3_p & v8455ab;
assign v3778fda = hgrant2_p & v373a568 | !hgrant2_p & v376c883;
assign v37770d2 = hgrant2_p & v376ea4a | !hgrant2_p & v3736da4;
assign v3768e1e = jx3_p & v372969d | !jx3_p & v374c4c0;
assign v37535d9 = hbusreq5_p & v37320f4 | !hbusreq5_p & v8455ab;
assign v374c70d = hbusreq6_p & v3726c67 | !hbusreq6_p & v3a657bf;
assign v37659e2 = hgrant6_p & v3a6dfc9 | !hgrant6_p & v8f559e;
assign v9f7a48 = hbusreq3_p & v3745b4f | !hbusreq3_p & v35772a6;
assign v3a6f70d = hbusreq3_p & v3a635ea | !hbusreq3_p & v376d98c;
assign v3773103 = hbusreq5_p & v37763d1 | !hbusreq5_p & v373b02e;
assign v3777e08 = hbusreq1_p & v3748bb1 | !hbusreq1_p & v3767399;
assign v374d6b2 = hbusreq2_p & v3a62a6d | !hbusreq2_p & v3a70b17;
assign v373dbbb = hbusreq7_p & v377cd7f | !hbusreq7_p & v375aeb3;
assign v375ad1d = hgrant4_p & v376e914 | !hgrant4_p & v3a5f3e3;
assign v3a6bb84 = hgrant6_p & v3743b9e | !hgrant6_p & v3727db9;
assign v3744f62 = hbusreq4 & v3751734 | !hbusreq4 & v8455ab;
assign v3a6f938 = hlock7_p & v377d91c | !hlock7_p & !v3a6eb09;
assign v372c467 = hlock5 & v37325ed | !hlock5 & afadd1;
assign v3747a0d = hmaster2_p & v374282f | !hmaster2_p & !v372a0b0;
assign v3809d45 = hbusreq0 & v372b858 | !hbusreq0 & v373e76a;
assign v3728a45 = hmaster0_p & v3a709ee | !hmaster0_p & v376b561;
assign v3a6fc5d = hmaster1_p & v374a0ac | !hmaster1_p & v3777527;
assign v3754877 = hlock3 & v373dfb8 | !hlock3 & v376f332;
assign v3774acc = hgrant6_p & v3a5836e | !hgrant6_p & v3729cbe;
assign v3a64d96 = hbusreq7_p & v3777988 | !hbusreq7_p & v3a6ef8f;
assign v373b956 = hmaster0_p & v374729b | !hmaster0_p & !v3a692c3;
assign v3a70a90 = hmaster1_p & v3807aa1 | !hmaster1_p & v37383d3;
assign v376bca9 = hgrant4_p & v375f486 | !hgrant4_p & !v8455ab;
assign v375dbda = hbusreq7 & v3a5baf5 | !hbusreq7 & v3a62f14;
assign v3a70caf = hlock6_p & v3a615a2 | !hlock6_p & v8455ab;
assign v3a710c1 = hbusreq6_p & v373014d | !hbusreq6_p & v3752000;
assign v3757440 = hgrant6_p & v8455c9 | !hgrant6_p & v1e3732b;
assign v376af64 = hmaster0_p & v375808f | !hmaster0_p & v37333a4;
assign v3747956 = hlock1_p & v37673f7 | !hlock1_p & v374668d;
assign v376a21e = hgrant6_p & v37796ee | !hgrant6_p & v3a63203;
assign v377adc8 = stateA1_p & v8455ab | !stateA1_p & !v3a5a496;
assign v374e590 = hmaster1_p & v374ab34 | !hmaster1_p & !v3a70f10;
assign v3a6fde9 = hbusreq2_p & v37291d1 | !hbusreq2_p & v373d4c6;
assign v3749d3f = hbusreq4 & v374852b | !hbusreq4 & v3a6eb47;
assign v3a70fed = hmaster0_p & v3a5950d | !hmaster0_p & v3a7045e;
assign v372863f = hmaster1_p & v3a635ea | !hmaster1_p & v375d9df;
assign v3a6fcfe = hbusreq3 & v373aecf | !hbusreq3 & !v8455ab;
assign v3778425 = hbusreq2 & v3733c46 | !hbusreq2 & v8455ab;
assign v3a69ed9 = hbusreq4_p & v3749001 | !hbusreq4_p & v3735f25;
assign v374ce92 = hgrant0_p & v8455ab | !hgrant0_p & v3753233;
assign v376ffb4 = hlock5_p & v3733e4f | !hlock5_p & v3a57b46;
assign v377f734 = hgrant4_p & v8455ab | !hgrant4_p & v37355d8;
assign v374e43d = hlock2 & v3747569 | !hlock2 & v373f622;
assign v37779ea = locked_p & v373414c | !locked_p & !v8455ab;
assign v3a70927 = hmaster0_p & v3a6c050 | !hmaster0_p & v3a55cc4;
assign v3809dfb = hbusreq5 & v3a7017d | !hbusreq5 & v3a7161b;
assign v3a6f70b = hmaster1_p & v37793e4 | !hmaster1_p & v3748ba9;
assign v3a6ac2a = stateA1_p & v37440c3 | !stateA1_p & v2acb5a2;
assign v377e869 = hmaster0_p & v3a5e60c | !hmaster0_p & v374b68a;
assign v23fe03a = hlock0_p & v374ab5b | !hlock0_p & v3769283;
assign v372ed55 = hbusreq4_p & v3739ea3 | !hbusreq4_p & v3757a57;
assign v376db8f = hbusreq4 & v37577e7 | !hbusreq4 & v8455ab;
assign v3a6373e = hbusreq5_p & v372c524 | !hbusreq5_p & v8455ab;
assign v3750c92 = hlock3_p & v3775b81 | !hlock3_p & v8455ab;
assign v3a6fa35 = hmaster2_p & v35772a6 | !hmaster2_p & v377bb6d;
assign v37610e5 = hmaster2_p & v3a701c4 | !hmaster2_p & v3a6152c;
assign v3807ddf = stateG10_1_p & v3767642 | !stateG10_1_p & v3a5db66;
assign v372e365 = hlock5_p & v3a66667 | !hlock5_p & v376dea1;
assign v3a29844 = hgrant5_p & v8455c6 | !hgrant5_p & bb41ad;
assign v3a64f05 = hlock2 & v3748797 | !hlock2 & v3a5a16b;
assign v3a66e9f = hmaster0_p & v37358ab | !hmaster0_p & !v3a70da2;
assign v3a6f0cc = hbusreq3 & v377d705 | !hbusreq3 & v377437a;
assign v377de7b = hbusreq2_p & v3a708d1 | !hbusreq2_p & v8455ab;
assign v3a7143d = hbusreq5 & v8455b0 | !hbusreq5 & v377edd6;
assign v3726c8e = hgrant5_p & v8455ab | !hgrant5_p & v3a71659;
assign v377f32e = hgrant4_p & v3758e05 | !hgrant4_p & v3731803;
assign v37756df = hbusreq7 & v37581f6 | !hbusreq7 & v3a6fdab;
assign v372b765 = hlock3_p & v37285a1 | !hlock3_p & v3a6f8dc;
assign v3768734 = hgrant5_p & v375478f | !hgrant5_p & v3a71693;
assign v37345a4 = hbusreq7_p & v3723698 | !hbusreq7_p & v3731800;
assign v3747931 = hmaster2_p & v8455ab | !hmaster2_p & v376646f;
assign v3a70210 = hbusreq4 & v3755820 | !hbusreq4 & v2092abe;
assign v3a716a4 = hgrant5_p & v8455ab | !hgrant5_p & v372a24d;
assign v3a6f48f = hlock3 & v376aa7a | !hlock3 & v372d880;
assign v373be9e = hgrant0_p & v8455ab | !hgrant0_p & v373fc30;
assign v373687f = hbusreq3_p & v3773871 | !hbusreq3_p & v3806912;
assign v3a6130e = hbusreq7 & v3a6fd76 | !hbusreq7 & v3736684;
assign v3a62e3c = hbusreq7_p & v3725948 | !hbusreq7_p & v3758bbf;
assign v3736fb4 = hbusreq5 & v376e74b | !hbusreq5 & v377ee7c;
assign v375de43 = hmaster2_p & v8455ab | !hmaster2_p & v377c44f;
assign v3a705d2 = hgrant5_p & v8455c6 | !hgrant5_p & v376b89f;
assign v3744117 = hbusreq4 & v3a6bf12 | !hbusreq4 & v3a6b53f;
assign v3a6fbfd = hmaster1_p & v37566b2 | !hmaster1_p & v376a752;
assign a65142 = hmaster0_p & v3a71654 | !hmaster0_p & be54b2;
assign v3a708fb = hbusreq5 & v3a7016b | !hbusreq5 & v373eadd;
assign v375b21c = hlock0_p & v374e0ba | !hlock0_p & v3a702ed;
assign v377a478 = hbusreq6_p & v3a69e8c | !hbusreq6_p & v373ae91;
assign v3756bc9 = locked_p & v39ebac7 | !locked_p & v3a70c07;
assign v3a714b9 = hlock5_p & v3a6e31f | !hlock5_p & !v3772e82;
assign v3a6faef = hgrant6_p & v3a70d99 | !hgrant6_p & v1e37a04;
assign v3a707b4 = jx0_p & v8b32e5 | !jx0_p & v2ff8e3d;
assign v3a708d8 = hgrant5_p & v3742dcb | !hgrant5_p & v37398a1;
assign v375d263 = hgrant4_p & v3a6ffb6 | !hgrant4_p & v377ed24;
assign v3a59900 = hbusreq7 & v376025c | !hbusreq7 & !v8455c2;
assign v3724a2c = hgrant6_p & v377938d | !hgrant6_p & v373f63e;
assign v3739443 = stateG10_1_p & v3a6fe6a | !stateG10_1_p & v3a703df;
assign v377a6c4 = hready_p & v372fddd | !hready_p & v3744f80;
assign a12203 = hlock0_p & v375803a | !hlock0_p & v3a6f849;
assign v3a5ae05 = hbusreq5 & v23fe1ad | !hbusreq5 & v3a6ff16;
assign v375d640 = hmaster0_p & v3728d9c | !hmaster0_p & v3738906;
assign v375956a = hmastlock_p & v8455e3 | !hmastlock_p & v8455ab;
assign v373a0d6 = hmaster2_p & v373d9e0 | !hmaster2_p & v3764a2d;
assign v376d3cb = hmaster1_p & v3a70a57 | !hmaster1_p & v373bbb4;
assign v37588c4 = hbusreq4 & v37482f8 | !hbusreq4 & !v377acae;
assign v372802c = hlock0_p & v3a635ea | !hlock0_p & v3a6f1fd;
assign v376980f = hmaster0_p & v3a6dfb2 | !hmaster0_p & v3a63989;
assign v3a705b9 = hbusreq4_p & v3a6f9c4 | !hbusreq4_p & v3766285;
assign v3a7015e = hmaster1_p & v372ba66 | !hmaster1_p & v373a7ab;
assign v3a6784d = hbusreq2_p & v3a67261 | !hbusreq2_p & v8455b3;
assign v3a6eec5 = hbusreq5_p & v3255a34 | !hbusreq5_p & v37741bd;
assign v3a70103 = hmaster2_p & v372adb5 | !hmaster2_p & v3a70ca8;
assign v372b32f = hmaster2_p & v8455ab | !hmaster2_p & v3a603fc;
assign v3a7116b = hbusreq1_p & v37684ed | !hbusreq1_p & v8455ab;
assign v377766c = hbusreq0 & v3737c2f | !hbusreq0 & v8455ab;
assign v3a71615 = hbusreq4 & v3748de3 | !hbusreq4 & v373f0ee;
assign v374ff84 = hbusreq5 & v3a70a01 | !hbusreq5 & v8455ab;
assign v374c1a9 = hgrant2_p & v8455ab | !hgrant2_p & v3a65a33;
assign v3768ba1 = hbusreq4_p & v3a6a261 | !hbusreq4_p & v372e6a1;
assign v3a6b8e8 = hlock5 & v3a6094b | !hlock5 & v3a6fec1;
assign v3a6eef7 = hmaster2_p & v3a71484 | !hmaster2_p & v3765e46;
assign v3a6fddb = hgrant5_p & v373ad69 | !hgrant5_p & v37435e1;
assign v3750002 = hgrant6_p & v374f7b7 | !hgrant6_p & v377f15c;
assign v3a5c40b = hmaster1_p & v3a6fc18 | !hmaster1_p & v8455ab;
assign v3a7072e = hmaster1_p & v374875f | !hmaster1_p & v3a70144;
assign v3a6f44e = hlock0 & v38072fd | !hlock0 & v3a6ef4d;
assign v3a5507a = hbusreq6 & v3723542 | !hbusreq6 & v3a6da8a;
assign v3778151 = hbusreq6_p & v3806e0e | !hbusreq6_p & v3758988;
assign v377dacb = hgrant4_p & v8455ab | !hgrant4_p & v3a55641;
assign v3a69606 = hmaster2_p & v374ecd5 | !hmaster2_p & v373aaa8;
assign v376b6fb = hbusreq8_p & cc8eeb | !hbusreq8_p & v8455ab;
assign v3a5c576 = hmaster0_p & v3747c23 | !hmaster0_p & d26e1e;
assign v376c8f2 = hlock7 & v376c313 | !hlock7 & v3771428;
assign v3739e36 = hmaster0_p & v376bd43 | !hmaster0_p & v37270a2;
assign v3729eb0 = hlock5_p & v8455ab | !hlock5_p & v372d727;
assign v3a61cbf = hlock3 & v3a6fb62 | !hlock3 & v375969d;
assign v3776018 = hbusreq7_p & v3746877 | !hbusreq7_p & v3762c4c;
assign v374a7b2 = hgrant2_p & v8455ba | !hgrant2_p & v9ccd8a;
assign v37476fd = hbusreq6_p & v8455b7 | !hbusreq6_p & v3a6dcdc;
assign v3a6fb40 = hmaster0_p & v376ea59 | !hmaster0_p & v3a58d68;
assign v3a5fe72 = hlock2_p & v3a564a8 | !hlock2_p & v373cb2d;
assign v3767f9a = hmaster0_p & v3a7002c | !hmaster0_p & bb4062;
assign v3a5e7e8 = hmaster3_p & v3a712b5 | !hmaster3_p & a7e544;
assign v37652ae = hbusreq7_p & v3809380 | !hbusreq7_p & v39a4ca6;
assign v377230a = hmaster2_p & v8455c3 | !hmaster2_p & !v373ab12;
assign v3739e70 = hgrant2_p & v374bf8a | !hgrant2_p & v3765968;
assign v37474b8 = hlock2 & v374dd61 | !hlock2 & v3773c69;
assign v3a60bae = hmaster1_p & v37509fc | !hmaster1_p & v3773ee7;
assign d18baa = hmaster1_p & v377234d | !hmaster1_p & v377bd63;
assign v3a6f8a1 = hmastlock_p & v374ca2d | !hmastlock_p & v8455ab;
assign v37586e2 = hbusreq8_p & v35b7174 | !hbusreq8_p & v372d2d2;
assign v374177f = hgrant2_p & v8455ab | !hgrant2_p & !v3a6eb3c;
assign v3a540f3 = hbusreq1 & v375de18 | !hbusreq1 & v8455ab;
assign v375da09 = hbusreq3 & v3747cf5 | !hbusreq3 & !v8455ab;
assign v376d979 = hmaster0_p & v377dfbf | !hmaster0_p & v374f6f9;
assign v373c076 = hmaster2_p & v2ff8bbc | !hmaster2_p & v37320ff;
assign v376c945 = hmaster2_p & v8455ab | !hmaster2_p & v375bf9a;
assign v375fe58 = hmaster2_p & v377e31b | !hmaster2_p & v3a6fd72;
assign v3a6f706 = hmaster1_p & v3a6b924 | !hmaster1_p & v37419df;
assign v372ea14 = hbusreq6 & v3770a77 | !hbusreq6 & v3763004;
assign v3754a74 = hmaster0_p & v372a161 | !hmaster0_p & v373e16b;
assign v3a709e8 = hbusreq8 & v3a61e6a | !hbusreq8 & v377dc99;
assign v3a5d33e = hmaster1_p & v8455ab | !hmaster1_p & v3744806;
assign v3a7107a = hbusreq4 & v37583be | !hbusreq4 & v376b4e1;
assign v37731ec = hbusreq5 & v3a6f7ef | !hbusreq5 & v3739b5c;
assign v3a6ff15 = hmaster2_p & v3a6f995 | !hmaster2_p & v3726605;
assign v3748a5d = hlock8 & v375d8f8 | !hlock8 & v3a5de59;
assign v3768076 = hbusreq4 & v3a70fb2 | !hbusreq4 & v3a705c5;
assign v3a5aef2 = hmaster3_p & v3a6fb07 | !hmaster3_p & v1e378ce;
assign v375107e = hgrant4_p & v373d4ff | !hgrant4_p & v3749d78;
assign v3a6fdc0 = hmaster0_p & v3a6f000 | !hmaster0_p & v8455ab;
assign v373fe74 = hgrant6_p & v8455ca | !hgrant6_p & v376a006;
assign v3770e0e = hbusreq5 & v375eef0 | !hbusreq5 & v37c0296;
assign v3a6b0eb = hbusreq7 & v3a6094e | !hbusreq7 & v3757ebc;
assign v3728fa6 = hbusreq5 & v37500ae | !hbusreq5 & v357742d;
assign v3a675eb = hbusreq7 & v3a5f80f | !hbusreq7 & v373a8a1;
assign v3739808 = hbusreq8_p & v3776d62 | !hbusreq8_p & v3778032;
assign v373c665 = hbusreq6_p & v3739bd5 | !hbusreq6_p & !v8455ab;
assign v3775adf = hlock5_p & v3736894 | !hlock5_p & !v375a9c1;
assign v3a558c5 = hgrant2_p & v3a5c823 | !hgrant2_p & v3770bb9;
assign v3a70874 = hmaster0_p & v374c251 | !hmaster0_p & v374e6b1;
assign v3777f6f = hbusreq8 & v372cbdf | !hbusreq8 & v8455b3;
assign v3a55d64 = hmaster0_p & v3a6ac17 | !hmaster0_p & v3a6af83;
assign v37433d5 = hmaster0_p & v8455ab | !hmaster0_p & v376c945;
assign v373e8e3 = hmaster1_p & v8455e7 | !hmaster1_p & v37772c0;
assign v3722ac4 = hmaster0_p & v3a71291 | !hmaster0_p & v3a296dc;
assign v3762aaf = jx0_p & v3a712ae | !jx0_p & v377bbfc;
assign v37338bb = hmaster2_p & v373b166 | !hmaster2_p & v377d58d;
assign v3a59299 = hmaster2_p & v3a5a807 | !hmaster2_p & v37466cb;
assign v375df71 = hlock5 & v3a62753 | !hlock5 & v3a6f59e;
assign v3736e8e = hbusreq0 & v37444b2 | !hbusreq0 & c7355c;
assign v376078d = hmaster1_p & v3806c9a | !hmaster1_p & v3743580;
assign v375d1d1 = hmaster0_p & v37793a6 | !hmaster0_p & v377a985;
assign v373ba4a = hbusreq6_p & v37434f6 | !hbusreq6_p & !v3747167;
assign v3777962 = hgrant0_p & v8455ab | !hgrant0_p & v37747fc;
assign v3a6113b = hlock6_p & v372ae4c | !hlock6_p & v3a5be6a;
assign v3a7031f = hbusreq3_p & v3a69de7 | !hbusreq3_p & v3a635ea;
assign d3a24d = hbusreq8 & v3a6a52c | !hbusreq8 & v3a57f04;
assign v375d7fc = hmaster2_p & v3766b95 | !hmaster2_p & v3a67d2f;
assign v372afd2 = hlock2 & v3752400 | !hlock2 & v3a67603;
assign v3761865 = hbusreq2 & v372e305 | !hbusreq2 & v8455ab;
assign v375d877 = hbusreq6_p & v39eb5ab | !hbusreq6_p & v37462e3;
assign v374b285 = hmaster2_p & v3a635ea | !hmaster2_p & v3a70374;
assign v3a588e5 = hbusreq5_p & v37702a1 | !hbusreq5_p & !v2092ac3;
assign v3739b18 = hbusreq7 & v377e9c9 | !hbusreq7 & v35b774b;
assign v3a71140 = hmaster0_p & v37770ae | !hmaster0_p & v3774878;
assign v3753964 = hlock0_p & v374c693 | !hlock0_p & v3738700;
assign v3762720 = hbusreq7_p & v37250b5 | !hbusreq7_p & v3a704d1;
assign v3a6a03c = hmaster1_p & v3a7152b | !hmaster1_p & v3751159;
assign v375c85c = hmaster1_p & v3a703d7 | !hmaster1_p & v3765dbe;
assign v2acafcc = hgrant4_p & v3759032 | !hgrant4_p & v3a6e81e;
assign v376fa86 = hlock7_p & v37385e9 | !hlock7_p & v3a296d3;
assign v3a6ccc4 = hlock5 & v3747ea2 | !hlock5 & v3a5e496;
assign v3749540 = hmaster0_p & v372e889 | !hmaster0_p & v3a66615;
assign v3740bb7 = hmaster0_p & v3a70e6a | !hmaster0_p & v373af66;
assign v372c0fd = hlock5 & v377142b | !hlock5 & v3a705d1;
assign v94b9e7 = hbusreq8 & v37667d3 | !hbusreq8 & v376fc7f;
assign v3a60229 = hmaster2_p & v3a635ea | !hmaster2_p & v374e9c0;
assign v2925cef = hbusreq7 & v37309ae | !hbusreq7 & v3762100;
assign v373058e = hmaster2_p & v3a6fcad | !hmaster2_p & v3a70cfc;
assign v3a697f1 = hlock4_p & v39a5265 | !hlock4_p & !v8455ab;
assign v377aa7a = hbusreq0 & v3726905 | !hbusreq0 & v8455ab;
assign v37675f1 = hmaster0_p & v8455c2 | !hmaster0_p & !v37470e2;
assign v3776cad = hmaster1_p & v3a5762d | !hmaster1_p & v372ef3e;
assign v3763295 = hbusreq6_p & v3a69eb7 | !hbusreq6_p & v8455ab;
assign v3a5bac7 = hlock0 & v3a6f43a | !hlock0 & v376a97b;
assign v3a6c835 = hgrant2_p & v377b6ce | !hgrant2_p & v373f4a5;
assign v372f9cf = hmaster2_p & v3a5cb57 | !hmaster2_p & v377c38c;
assign v3764312 = hlock2 & v3748797 | !hlock2 & v376144f;
assign v3a71581 = hmaster1_p & v3a6ff25 | !hmaster1_p & v3771555;
assign v3778f25 = hlock7 & v3a5f546 | !hlock7 & v3741736;
assign v3727807 = hbusreq6 & aef673 | !hbusreq6 & v3a7011e;
assign v3748de3 = hlock6 & v3744877 | !hlock6 & v3742905;
assign v3a6f3af = hgrant6_p & v8455ab | !hgrant6_p & v375adaa;
assign v37309cf = hlock2_p & v3a64f4f | !hlock2_p & !v8455ab;
assign v3724940 = hready & v3732eca | !hready & v3a5ca7b;
assign v377c258 = hbusreq6_p & v3a70d86 | !hbusreq6_p & v8455ab;
assign v3a70384 = hgrant4_p & v3a6f71a | !hgrant4_p & v37763c2;
assign v373aa76 = hlock8_p & v376faa6 | !hlock8_p & v374df88;
assign v3a6f731 = hbusreq8_p & v3779c8d | !hbusreq8_p & v3a6299c;
assign v375a0ad = hlock5 & v3735760 | !hlock5 & v373809d;
assign v3a6f139 = hbusreq4 & v376cf3f | !hbusreq4 & v373bd6c;
assign v3737193 = hbusreq6_p & v375e7aa | !hbusreq6_p & v8455ab;
assign v3752201 = hgrant3_p & v8455e7 | !hgrant3_p & !v3772ab1;
assign v375c432 = hmaster2_p & v3a70374 | !hmaster2_p & v3a63df4;
assign v37409c7 = hbusreq5 & v380971d | !hbusreq5 & v376d091;
assign v37438fc = hmaster0_p & v3a6f475 | !hmaster0_p & v374e0a9;
assign v3736c7e = hmaster1_p & v374d4e6 | !hmaster1_p & v37363da;
assign v376f9a8 = locked_p & v3a70cd5 | !locked_p & v3809adf;
assign v37716b0 = hbusreq8 & v37756df | !hbusreq8 & v37331e1;
assign v3768aaa = hbusreq1_p & v8455ab | !hbusreq1_p & !v8455b0;
assign v3771728 = hbusreq1_p & v3a6ebff | !hbusreq1_p & !v3760582;
assign v373ace1 = hlock4 & v372c1b0 | !hlock4 & v3728ea7;
assign v3a634eb = hmaster2_p & v3736be1 | !hmaster2_p & v8455ab;
assign v373397b = hbusreq2_p & v377eaf2 | !hbusreq2_p & v3a6f79e;
assign v3a5f5d0 = hgrant8_p & v376a129 | !hgrant8_p & v3a6f77b;
assign v3a5c7a2 = hmaster0_p & v372625f | !hmaster0_p & v3761300;
assign v3a70049 = hgrant4_p & v3a5b5d3 | !hgrant4_p & !v3a5f3e3;
assign v3737b63 = hlock5 & v23fdec8 | !hlock5 & v3a70927;
assign v3722d5a = hmaster0_p & v375058e | !hmaster0_p & v376ad77;
assign v372eff2 = hgrant4_p & v8455ab | !hgrant4_p & v373f200;
assign v3724798 = hbusreq5_p & v3a6f4f3 | !hbusreq5_p & v375cd50;
assign v3a66a8e = hbusreq8 & v3a6fc84 | !hbusreq8 & v8455ab;
assign v372b7a3 = hmaster2_p & v37423d1 | !hmaster2_p & v3a6eeef;
assign v3a2976f = hmaster0_p & v3807020 | !hmaster0_p & !v3a56b7c;
assign v373c228 = hbusreq7 & v3a66c94 | !hbusreq7 & v3744c5e;
assign v374b497 = hmaster0_p & v8455c2 | !hmaster0_p & v374da1a;
assign v3807765 = hmaster2_p & v8455ab | !hmaster2_p & !v3a71133;
assign v3772dd2 = hmaster0_p & v376999f | !hmaster0_p & v3a61dca;
assign v3a7009f = hmaster0_p & v8455ab | !hmaster0_p & v37493c7;
assign v3806e7b = hgrant6_p & v37c039c | !hgrant6_p & v3a7042a;
assign v3a6f164 = hmaster2_p & v375ac50 | !hmaster2_p & v3736b71;
assign v37342e7 = hmaster0_p & v376f858 | !hmaster0_p & v376bbbe;
assign v373ec34 = hmaster0_p & v3a6e846 | !hmaster0_p & v37766fb;
assign v3a5e485 = hbusreq3_p & v3735e39 | !hbusreq3_p & !v3a6d684;
assign v3726464 = hbusreq0_p & v3740171 | !hbusreq0_p & v37457fb;
assign v37658de = hlock8_p & v3a66da0 | !hlock8_p & v374af1f;
assign v92bc1e = jx0_p & v3770ee4 | !jx0_p & v374cb5e;
assign v3a6f6ba = hbusreq2_p & v374ba65 | !hbusreq2_p & v3a710d2;
assign v37702e6 = hbusreq7_p & v374fa66 | !hbusreq7_p & v8455ab;
assign v37560ef = hmaster0_p & v3a713b8 | !hmaster0_p & v373f7a5;
assign v372d880 = hgrant0_p & v3a714f5 | !hgrant0_p & v3758e5f;
assign v376a6d6 = hbusreq0_p & v377b673 | !hbusreq0_p & b27f78;
assign v3770187 = hbusreq0_p & v8455b7 | !hbusreq0_p & v374e61f;
assign v3a5aca8 = hlock4_p & v37507d0 | !hlock4_p & v8455ab;
assign v375d387 = hbusreq5_p & v3726594 | !hbusreq5_p & !v3a66110;
assign v377bdb2 = hbusreq5_p & v3762790 | !hbusreq5_p & v8455ab;
assign v3a6f3cd = hmaster2_p & v3a71267 | !hmaster2_p & v3725717;
assign v3a587a1 = hmaster1_p & v8455ab | !hmaster1_p & v3806b2d;
assign v3a6a289 = hgrant4_p & v3a6ef50 | !hgrant4_p & !v373554b;
assign v3a625f8 = hgrant2_p & v8455ab | !hgrant2_p & v374e43d;
assign v3761678 = hgrant3_p & v372abd8 | !hgrant3_p & v376d251;
assign v377118b = hlock8 & v3a6a1d9 | !hlock8 & v3748d6c;
assign v3736ad7 = hmaster0_p & v372625f | !hmaster0_p & v374d1dc;
assign v3a705f0 = hlock6_p & v3a709ea | !hlock6_p & v3a70131;
assign v3a7137d = hmaster1_p & v375fb00 | !hmaster1_p & v3a5cf3c;
assign v3776a27 = hgrant2_p & v375d12e | !hgrant2_p & v3806fa6;
assign v375d6ba = hgrant2_p & v8455ab | !hgrant2_p & v373fbc7;
assign v374b8cb = hgrant3_p & v3a70272 | !hgrant3_p & !v374db9d;
assign v377d34b = hgrant0_p & v3a70233 | !hgrant0_p & v376f30a;
assign v3809e97 = hmaster1_p & v3734f6d | !hmaster1_p & v3a68377;
assign v375ed52 = busreq_p & v3726dfa | !busreq_p & v377670f;
assign v3a70662 = hbusreq8 & b44720 | !hbusreq8 & v3a5666f;
assign v3758299 = hlock0 & v37450b8 | !hlock0 & v3a697e4;
assign v3754cb0 = hmaster2_p & v37270bc | !hmaster2_p & v3a6f2cb;
assign v372d24d = hbusreq8_p & v3760ac5 | !hbusreq8_p & v377a75f;
assign v3a5c5e1 = hmaster1_p & v8455ab | !hmaster1_p & v3734df5;
assign v375a1a7 = hbusreq5_p & v3730055 | !hbusreq5_p & v373cc82;
assign v375e551 = hgrant3_p & v376ace9 | !hgrant3_p & v3761af1;
assign v3a5dba4 = hmaster2_p & v3a70c39 | !hmaster2_p & v3752dd0;
assign v3758466 = hmaster0_p & v3a65d93 | !hmaster0_p & v37281fb;
assign v3a5915c = hgrant4_p & v8455ab | !hgrant4_p & v3809ec3;
assign v37649c2 = hmaster2_p & v8455b0 | !hmaster2_p & v3770116;
assign v3a5dcfc = hlock2 & v372dc5c | !hlock2 & v3a6f70d;
assign v373c583 = hmaster2_p & v373006f | !hmaster2_p & v373f503;
assign v3778cba = hmaster0_p & v3a6f463 | !hmaster0_p & v3a56512;
assign v3731a5a = hgrant6_p & v3764486 | !hgrant6_p & v3a5a5d1;
assign v375eb56 = hbusreq4 & v3a71453 | !hbusreq4 & !v8455b9;
assign v3752edb = hlock7_p & v377933b | !hlock7_p & v376ed36;
assign v3775de3 = hbusreq6 & v3729f6a | !hbusreq6 & v373867c;
assign v380678d = hbusreq0 & v3764a07 | !hbusreq0 & v3753903;
assign v376256f = hbusreq5_p & v3a6fd84 | !hbusreq5_p & !v3a7122f;
assign v373ef69 = hbusreq4_p & v3739fff | !hbusreq4_p & !v3a7151d;
assign v3761bee = hmaster2_p & v3752cc5 | !hmaster2_p & v3734634;
assign b9f306 = hmaster1_p & v3808865 | !hmaster1_p & v3750edc;
assign v3a694ec = hmaster2_p & v8455ab | !hmaster2_p & !v3a69cd8;
assign v376d240 = hgrant2_p & v377182c | !hgrant2_p & v37699c9;
assign v3a6dafc = hmaster2_p & v376ac08 | !hmaster2_p & v3739ddf;
assign v376a3c2 = hmaster2_p & v3a635ea | !hmaster2_p & v3743b9e;
assign v377e9c4 = hbusreq3_p & v3a7045c | !hbusreq3_p & v373dafc;
assign v3a6f434 = hgrant2_p & v3755c7c | !hgrant2_p & v372ccbb;
assign v3756483 = hgrant6_p & v3728d72 | !hgrant6_p & v3770cf6;
assign v374ad45 = hmaster0_p & v3a635ea | !hmaster0_p & v3732bf9;
assign v373809d = hmaster0_p & v3740f94 | !hmaster0_p & v375d2b3;
assign v3a6f485 = hgrant2_p & v372f09a | !hgrant2_p & v3a6fff7;
assign v376f0f6 = hmaster2_p & v3747302 | !hmaster2_p & v376e041;
assign v3a6f0bc = hgrant4_p & v3a6143f | !hgrant4_p & v3747c3d;
assign v37369f2 = hbusreq0 & v376791c | !hbusreq0 & v372ecd8;
assign v35b7169 = hbusreq5_p & v372b9c5 | !hbusreq5_p & v3a6f0d5;
assign v37722c6 = hgrant3_p & v37765fe | !hgrant3_p & v3774913;
assign bde868 = hmaster0_p & v3a696a7 | !hmaster0_p & v3a62efa;
assign v373165b = hmaster2_p & v8455ab | !hmaster2_p & v3a56642;
assign v376df9f = hmaster0_p & v3a606e6 | !hmaster0_p & !v3770a68;
assign v3a6ae0f = hbusreq5 & v3770425 | !hbusreq5 & v3a6eed9;
assign v3a585b7 = hmaster0_p & v37657e4 | !hmaster0_p & v8455bd;
assign v3a6f9ac = hlock0 & v3a635ea | !hlock0 & v376a272;
assign v376e2a4 = hmaster1_p & v375f2a3 | !hmaster1_p & v376d215;
assign v372ff70 = hbusreq4 & v376495e | !hbusreq4 & v8455ab;
assign v3753329 = hlock4_p & v3a6672b | !hlock4_p & !v8455ab;
assign v3748cbd = hlock0_p & v372dadb | !hlock0_p & cf4a8f;
assign v375610e = hbusreq8 & v377cd68 | !hbusreq8 & v372ad2c;
assign v37293e9 = hmaster1_p & v377bdb2 | !hmaster1_p & v3a70550;
assign v372428a = hmaster1_p & v3a619c0 | !hmaster1_p & v3a6eaba;
assign v3758539 = hbusreq2_p & v3a577f2 | !hbusreq2_p & !v3a687ea;
assign v3a65909 = hmaster2_p & v8455ab | !hmaster2_p & v3765e46;
assign v375a4f8 = hbusreq5_p & v376a915 | !hbusreq5_p & v3774449;
assign v375dbd4 = hbusreq2_p & v8455e1 | !hbusreq2_p & v3a6f549;
assign v373ac84 = hgrant5_p & v3728a53 | !hgrant5_p & v3a5d185;
assign v3738686 = hmaster2_p & v8455ab | !hmaster2_p & v37346be;
assign v3a6f63a = hmaster0_p & v3769ae2 | !hmaster0_p & v37311fa;
assign v375bf36 = hbusreq7 & v23fe343 | !hbusreq7 & a0a219;
assign v37740f9 = hgrant2_p & v3a6fa0d | !hgrant2_p & v374f29f;
assign v373de13 = hbusreq6_p & v3747302 | !hbusreq6_p & v3a6ff18;
assign v3726be0 = hbusreq6_p & v37261df | !hbusreq6_p & !v3a5ae7d;
assign v3730a6a = hgrant5_p & v8455bd | !hgrant5_p & v3776eff;
assign v2acafff = hbusreq3 & v373be9e | !hbusreq3 & v8455ab;
assign v3747623 = hbusreq2_p & v3a71065 | !hbusreq2_p & v3a5b68a;
assign v3a6fc91 = hbusreq5_p & v3a64abe | !hbusreq5_p & v3a70d5d;
assign b6390c = hgrant2_p & v8455b0 | !hgrant2_p & v37677ee;
assign v3a709c2 = jx0_p & v37565d3 | !jx0_p & v8455ab;
assign v374544c = hmaster0_p & v3806ff5 | !hmaster0_p & v3a5f992;
assign v3744a2f = locked_p & v374c9c7 | !locked_p & v3a619c0;
assign v37283fc = hbusreq2_p & a875ea | !hbusreq2_p & v3761d4e;
assign cb1cc0 = hlock6 & v37577db | !hlock6 & v377d41d;
assign v3a68c23 = hlock4_p & v3742122 | !hlock4_p & v375d616;
assign v375523e = hbusreq5_p & v3722a6f | !hbusreq5_p & v3a6ff16;
assign v3723e00 = hmaster1_p & v97ea11 | !hmaster1_p & v372d237;
assign v373bd70 = hbusreq8 & v3377adc | !hbusreq8 & v376775d;
assign v3733b9a = hbusreq7 & v3763a12 | !hbusreq7 & v3a6f9fa;
assign v37337d2 = hbusreq0 & v376b5ad | !hbusreq0 & v3a6f03e;
assign v3a714a3 = hmaster0_p & v8455b0 | !hmaster0_p & v3a715c5;
assign v3a70ac7 = hgrant6_p & v377f09a | !hgrant6_p & !v3a6fbdd;
assign v376ce90 = hbusreq8 & v3a6fda8 | !hbusreq8 & v374a262;
assign v3758a96 = hmaster2_p & v3a67d66 | !hmaster2_p & ca01e4;
assign v3a7103c = hbusreq1 & v39a5265 | !hbusreq1 & !v3a6ac26;
assign v3a6f50c = hbusreq5_p & v3736a50 | !hbusreq5_p & !v8455ab;
assign v373cf60 = hgrant6_p & v3a70bd6 | !hgrant6_p & v3a60130;
assign v38076b7 = hmaster1_p & v3a29814 | !hmaster1_p & v3a6acd3;
assign v3a70bcd = hmaster2_p & v377766c | !hmaster2_p & !v3767e76;
assign v373fd4c = hmaster2_p & v8455ab | !hmaster2_p & v3769e7f;
assign v38096d8 = jx1_p & v374b237 | !jx1_p & !v3a69feb;
assign v372d366 = hgrant6_p & v8455ab | !hgrant6_p & v3a63df6;
assign v3a6f415 = hlock0_p & v3779324 | !hlock0_p & v373da69;
assign v372e02d = hbusreq7 & v376cb10 | !hbusreq7 & v3a5f55e;
assign v3722f58 = hbusreq3 & v37566f4 | !hbusreq3 & v3a6c5fc;
assign v37664c5 = hbusreq5 & v372c6c4 | !hbusreq5 & v3a70041;
assign v3a70c3e = hgrant4_p & v8455c1 | !hgrant4_p & v373141b;
assign v3a695fc = hbusreq3_p & v376fa38 | !hbusreq3_p & !v1e38224;
assign v3a6fcba = hgrant6_p & v3772c51 | !hgrant6_p & v3740f3d;
assign v3a63559 = hbusreq0 & v8455e1 | !hbusreq0 & v8455ab;
assign v375f87b = hmaster2_p & v37386f5 | !hmaster2_p & !v376641b;
assign v376b27a = hmaster0_p & v377d1dc | !hmaster0_p & v375d06a;
assign v3a7002a = hlock4 & v3779a88 | !hlock4 & v375c976;
assign v3808fce = hlock0 & v3a5aacb | !hlock0 & v3746d4a;
assign v37285fa = hmaster0_p & v3746a81 | !hmaster0_p & v37628cd;
assign v8b51d2 = hgrant4_p & v3a6eaf3 | !hgrant4_p & v3730ad2;
assign v3a70f09 = hbusreq5 & v3a7161b | !hbusreq5 & v2925d03;
assign v3764276 = locked_p & v3a637dc | !locked_p & v3750746;
assign v374145d = hbusreq0 & v3768c16 | !hbusreq0 & !v3733278;
assign v3759536 = hbusreq6 & v3a7116e | !hbusreq6 & v3755a05;
assign v3a6e7ae = hgrant8_p & v3756f21 | !hgrant8_p & v374ea10;
assign v3774d9c = hbusreq7_p & v3a6f28b | !hbusreq7_p & v377e852;
assign v374b824 = hmaster2_p & v3777b2e | !hmaster2_p & !v374cb97;
assign v376bfa7 = hbusreq5 & v374657b | !hbusreq5 & !v3a614d1;
assign v374a266 = hlock0_p & v374d836 | !hlock0_p & v3746824;
assign v3767640 = hbusreq8_p & v37621c1 | !hbusreq8_p & v376bd96;
assign v374f9c6 = hbusreq4_p & v37496fa | !hbusreq4_p & v3743b9e;
assign v372af77 = hgrant4_p & v37784ad | !hgrant4_p & v3a70183;
assign v3761287 = hbusreq5_p & v374ea19 | !hbusreq5_p & v23fe353;
assign v3a54b77 = hmaster0_p & v37594d4 | !hmaster0_p & v3775f25;
assign v374fc95 = hmaster1_p & v3a5c3a0 | !hmaster1_p & v376824b;
assign v372bf35 = hbusreq6 & v3a6f8de | !hbusreq6 & v3a62a6d;
assign v3752fbe = hmaster0_p & v8455e1 | !hmaster0_p & v374e409;
assign v3753d51 = hgrant6_p & v3a5a591 | !hgrant6_p & v3a6837d;
assign v376b035 = hmaster1_p & v3757966 | !hmaster1_p & v3a6f4a4;
assign v3a5d08a = hgrant6_p & v3741f22 | !hgrant6_p & v3769d5c;
assign v374c007 = hbusreq5 & v372e426 | !hbusreq5 & v374602f;
assign v3745c84 = hmaster0_p & v3734982 | !hmaster0_p & v3a6e93d;
assign v3774662 = hlock8_p & v3771df4 | !hlock8_p & !v8455ab;
assign v3a6fee5 = hgrant5_p & v3754328 | !hgrant5_p & v37770af;
assign v3727651 = hbusreq7 & v374c2d6 | !hbusreq7 & v3a70d99;
assign v3a6eff8 = hlock5_p & v3764ddc | !hlock5_p & v8f7302;
assign v3a637a1 = hmaster0_p & v37719a1 | !hmaster0_p & v8455b9;
assign v3a6f22a = hmaster2_p & v3a6fe0d | !hmaster2_p & v3a6143b;
assign v3736041 = hbusreq5_p & v3a6d7cd | !hbusreq5_p & v37d8c61;
assign v376ad4e = hlock0_p & v3770cd8 | !hlock0_p & v3a5cfed;
assign v3775cca = hbusreq5_p & v3a6fc73 | !hbusreq5_p & v3a5e38d;
assign v3a6f274 = hmaster3_p & v3727b7f | !hmaster3_p & v372ce4b;
assign v376822d = hlock7_p & v3769ee7 | !hlock7_p & !v8455ab;
assign v3753e23 = hbusreq5 & v3767f9a | !hbusreq5 & v3a70d26;
assign v3a70a7f = hbusreq3_p & v3a635ea | !hbusreq3_p & v373b288;
assign v3778091 = hgrant4_p & v8455ab | !hgrant4_p & v8955d0;
assign v374a6a5 = hbusreq6_p & v3a70c34 | !hbusreq6_p & !v8455ab;
assign v372b172 = hbusreq8 & v3723749 | !hbusreq8 & !v3a70570;
assign v37764a5 = hready & v3a6de33 | !hready & !v8455ab;
assign v3a6f8c1 = hlock1_p & v373fe5e | !hlock1_p & !v8455ab;
assign v3a54769 = hmaster1_p & v3a635ea | !hmaster1_p & v376c028;
assign v37645f6 = hmaster1_p & v374f307 | !hmaster1_p & v377521b;
assign v3a70f3b = hmaster1_p & v3a6f7dd | !hmaster1_p & v37754f6;
assign v3a6f8be = hmaster2_p & v376e914 | !hmaster2_p & v377b6ce;
assign v3a6f72e = hbusreq8_p & v372589e | !hbusreq8_p & v3a6be9f;
assign v3a541ee = hgrant2_p & v3a5f50e | !hgrant2_p & v3a552d4;
assign v3767abc = hbusreq1 & v3733383 | !hbusreq1 & v8455ab;
assign v37300d7 = hmaster1_p & v3a5d015 | !hmaster1_p & v3728203;
assign v37441dc = hgrant5_p & v8455ab | !hgrant5_p & v37665f9;
assign b4fa3c = hgrant1_p & v3743252 | !hgrant1_p & v8455ab;
assign v3a6f402 = hbusreq6_p & v372797f | !hbusreq6_p & v3a62d7d;
assign v3a5e776 = jx1_p & v375fa66 | !jx1_p & v3a6bd5a;
assign v373d35f = hbusreq6_p & v372d83d | !hbusreq6_p & !v8455ab;
assign v3769a2a = hmaster3_p & v372f039 | !hmaster3_p & v3751539;
assign v3743ada = hgrant2_p & v3a62524 | !hgrant2_p & v373449a;
assign v3a6beff = hlock7_p & v3a5b0b3 | !hlock7_p & v3726156;
assign v375f6e3 = hbusreq7 & v3a69961 | !hbusreq7 & v3a71478;
assign v374daa9 = hmaster1_p & v3763224 | !hmaster1_p & !v3a56847;
assign v3a70e47 = hlock5 & v3a6f8a9 | !hlock5 & v3a5eae2;
assign v3a625b1 = hmaster2_p & v3742cd4 | !hmaster2_p & !v8455ab;
assign v37287bd = hbusreq4 & v39a5381 | !hbusreq4 & v8455ab;
assign v373c151 = hbusreq3 & v3a6ab5f | !hbusreq3 & !v3a6ac26;
assign v3a6fb14 = hbusreq2_p & v373cf3a | !hbusreq2_p & v3a5b614;
assign v3a7033a = hbusreq4 & v3733383 | !hbusreq4 & v8455ab;
assign v375be2d = hgrant5_p & v373ad69 | !hgrant5_p & v3a5ba8a;
assign v3a714e0 = hbusreq7 & v3a5bc27 | !hbusreq7 & v8455b0;
assign v3752fcb = hlock5 & v3a700d7 | !hlock5 & v3758561;
assign v374578a = hgrant0_p & v3a58964 | !hgrant0_p & v3a71542;
assign v373fa04 = hmaster2_p & v373a1b4 | !hmaster2_p & v8455ab;
assign v3a70622 = hmaster2_p & v374da61 | !hmaster2_p & v374d54c;
assign v3743b64 = hmaster2_p & v3a6f806 | !hmaster2_p & v8455ab;
assign v3a70cf5 = hbusreq8 & v374dc99 | !hbusreq8 & !v376cef0;
assign v376f9ca = hmaster0_p & v8455e7 | !hmaster0_p & v377d769;
assign v2092abd = hmaster1_p & v373e376 | !hmaster1_p & v374e1f6;
assign v37671d3 = hmaster1_p & v3a6d3f2 | !hmaster1_p & v3a70bee;
assign v374513e = hbusreq3_p & v3a6f7a5 | !hbusreq3_p & v8455ab;
assign v3734b5a = hbusreq8 & v3a7132d | !hbusreq8 & v3723ddc;
assign v3727830 = hbusreq5 & v376c6fb | !hbusreq5 & v374e5fa;
assign v375b902 = hbusreq3 & v95d97e | !hbusreq3 & v8455ab;
assign v3757a57 = hbusreq0 & v377aa06 | !hbusreq0 & v372d967;
assign v372904d = hbusreq3_p & v3759f4c | !hbusreq3_p & v3a6eb83;
assign v376f152 = hgrant1_p & v37467f3 | !hgrant1_p & v8455ab;
assign v3727026 = hlock5 & v374cf82 | !hlock5 & v372bfd0;
assign v3a6fc04 = hmaster0_p & v3723fec | !hmaster0_p & v3744cd7;
assign v377ae32 = hmaster2_p & v3a62b5f | !hmaster2_p & v3728d9c;
assign v3a5fe5e = hgrant4_p & v8455ab | !hgrant4_p & v374f89b;
assign v376924d = hmaster1_p & v3743094 | !hmaster1_p & v3773dc6;
assign v375bdd4 = hlock0_p & v39a5265 | !hlock0_p & !v8455ab;
assign v3743b66 = hbusreq5_p & v3756b5c | !hbusreq5_p & v3a67c8e;
assign v376c94b = hbusreq7 & v37739af | !hbusreq7 & v8455ab;
assign v360d2c6 = hmaster0_p & v3a6fc9f | !hmaster0_p & !v8455ab;
assign v373738e = hbusreq8_p & v377f66c | !hbusreq8_p & v3a59283;
assign b2eec3 = hbusreq4_p & v3a635ea | !hbusreq4_p & v376819e;
assign v37457a8 = hbusreq8_p & v37563bc | !hbusreq8_p & v37576af;
assign v3a70e45 = hmaster0_p & v3763424 | !hmaster0_p & v3a6fad5;
assign v3a6535f = hmaster1_p & v3a6f875 | !hmaster1_p & !v3725042;
assign v3771a24 = hmaster1_p & v3752cac | !hmaster1_p & v3764daf;
assign v3a67c9e = hbusreq8_p & v3726ec0 | !hbusreq8_p & v37730ab;
assign v23fd9fe = hgrant5_p & v8455c6 | !hgrant5_p & v3a55162;
assign v373af1f = hbusreq4 & v372dccf | !hbusreq4 & v3a69487;
assign v375cda2 = hgrant4_p & v8455ab | !hgrant4_p & v3a687e0;
assign v3a62a8c = hgrant2_p & v3a62524 | !hgrant2_p & v3a70dd6;
assign v3a6f4ed = hbusreq0 & v3765021 | !hbusreq0 & v3a6f78a;
assign v375c6c1 = hmaster0_p & v37372a1 | !hmaster0_p & v374e51a;
assign v376f9d3 = hmaster1_p & v37430f0 | !hmaster1_p & v376fdbe;
assign v377b416 = hmaster0_p & v3a68b7b | !hmaster0_p & v3a70304;
assign v37691b8 = hbusreq7_p & v377d497 | !hbusreq7_p & v3a70cfa;
assign v3a708c1 = hbusreq5_p & v37775ff | !hbusreq5_p & v3a5ae8d;
assign v35b6a6b = hbusreq4 & v3752e63 | !hbusreq4 & v3a70d99;
assign v3a6ebf0 = hbusreq0_p & v372dadb | !hbusreq0_p & v377d8dd;
assign v374fb93 = hgrant3_p & v372abd8 | !hgrant3_p & !v3774061;
assign v37696a2 = hbusreq0 & v3772f26 | !hbusreq0 & v3724a2c;
assign v3a299f8 = hbusreq5_p & v37697ca | !hbusreq5_p & v3a5fa82;
assign v376b044 = hmaster2_p & v37267d6 | !hmaster2_p & v377d58d;
assign v3a6fab4 = hbusreq5_p & v37419df | !hbusreq5_p & v377405e;
assign v3728840 = hbusreq8 & v376079d | !hbusreq8 & v3a6ec01;
assign v373b166 = hbusreq0 & v3a6f908 | !hbusreq0 & v3752131;
assign v3a57796 = hlock8_p & v377d999 | !hlock8_p & !v8455ab;
assign v37331a1 = hbusreq0 & v3a709f3 | !hbusreq0 & v8455ab;
assign v37717ed = hmaster1_p & v377050f | !hmaster1_p & v37658d9;
assign v373c437 = hbusreq5_p & v3a6f45c | !hbusreq5_p & v3733fd0;
assign v3a711b2 = hbusreq4 & a0d21b | !hbusreq4 & v3a70d32;
assign v3a6f9a2 = hbusreq2_p & v3a6ae3e | !hbusreq2_p & v3a69946;
assign v3a67142 = hbusreq0 & v377e3ce | !hbusreq0 & !v1e37cd6;
assign v1e379d2 = hbusreq4 & v3a6fb29 | !hbusreq4 & v8455ab;
assign v3a6764b = hbusreq8_p & v3722f8e | !hbusreq8_p & v8455ab;
assign v3a5a6e6 = hgrant4_p & v3a5a807 | !hgrant4_p & ade0d8;
assign v3a708f4 = hmaster0_p & v37289f0 | !hmaster0_p & v37409cd;
assign v3726c67 = hbusreq6 & v3a5d469 | !hbusreq6 & v3a69487;
assign v376d98c = hlock3 & v3a70e84 | !hlock3 & v3806507;
assign v3a70b9a = hlock6 & v3a5f75a | !hlock6 & v3a6fa2c;
assign v3779d09 = jx0_p & v3a5a2d4 | !jx0_p & v8455ab;
assign v3a6857b = hmaster0_p & v377ce1a | !hmaster0_p & v3759586;
assign v377f887 = hmaster0_p & v3a5fc34 | !hmaster0_p & v3a6f2de;
assign v3a6d8ce = hbusreq1_p & v3a6e66e | !hbusreq1_p & !v3a5e8f6;
assign v37781fe = hmaster1_p & v3764276 | !hmaster1_p & v3a710a3;
assign v374e788 = hgrant5_p & v3a6046d | !hgrant5_p & !v8455ab;
assign v377a673 = hmaster1_p & v3a54aa0 | !hmaster1_p & v3a61a15;
assign v37508c4 = hmaster1_p & v380974c | !hmaster1_p & v375f67d;
assign v375d577 = hbusreq5 & v3778484 | !hbusreq5 & v3a71530;
assign v376cd02 = hmaster0_p & v3a6fac9 | !hmaster0_p & v380760a;
assign v3a663b9 = hbusreq0 & v373e2d3 | !hbusreq0 & v3a70275;
assign v3a694a5 = hlock8_p & v3750f1e | !hlock8_p & v3a6d3bc;
assign v3765cf3 = hbusreq5_p & d09db6 | !hbusreq5_p & ab11fe;
assign v3771214 = hlock8_p & v3744af7 | !hlock8_p & v3a714f8;
assign v3739b7a = hmaster2_p & v3770bcd | !hmaster2_p & v3a6f541;
assign v373cedd = hmaster2_p & v3735e39 | !hmaster2_p & !v376ea4a;
assign v3760066 = hbusreq8 & v376a9f5 | !hbusreq8 & v8455ab;
assign v37793cd = hbusreq5_p & v3735302 | !hbusreq5_p & !v8455ab;
assign v37776b6 = hbusreq6 & v3749907 | !hbusreq6 & v8455ab;
assign v3a5b885 = hgrant6_p & v8455ab | !hgrant6_p & v376b795;
assign v373d703 = hmaster0_p & v3748234 | !hmaster0_p & v23fe0c9;
assign v37551b9 = hgrant4_p & v3a6eb95 | !hgrant4_p & v373ec98;
assign v375f989 = hmaster0_p & v374a4d2 | !hmaster0_p & v3a69e22;
assign v3747d51 = hgrant8_p & v3a5397f | !hgrant8_p & !v3744b16;
assign v376c2a1 = hbusreq0 & v3a6b51b | !hbusreq0 & v375aa6b;
assign v3a5bea0 = hbusreq4 & v3737d44 | !hbusreq4 & v8455ab;
assign v3a6ef75 = hbusreq6_p & v37611c3 | !hbusreq6_p & v8455ab;
assign v375138c = hmaster0_p & v3a60976 | !hmaster0_p & v337902c;
assign v37324e7 = hmaster1_p & v373b2ba | !hmaster1_p & v377faa6;
assign v373557c = hbusreq6_p & v3a635ea | !hbusreq6_p & v3765e79;
assign v3769b1d = hmaster2_p & v3a5b7c2 | !hmaster2_p & !v3752fbc;
assign v3a6f1f5 = hmaster0_p & v8455ab | !hmaster0_p & v3741a83;
assign v3a70a5e = hbusreq0 & v3a715a8 | !hbusreq0 & d6eddf;
assign v374569b = hgrant2_p & v3758fa7 | !hgrant2_p & !v8455ab;
assign v3a6b15d = hbusreq6 & v37565a5 | !hbusreq6 & v3a57959;
assign v3773b55 = hbusreq2_p & v3a5d1fb | !hbusreq2_p & v3736da4;
assign v374aab3 = hbusreq7 & v375682e | !hbusreq7 & v3757b0f;
assign v3755252 = hbusreq0 & v3a5ae7d | !hbusreq0 & !v8455ab;
assign v373894d = hgrant4_p & v8455ab | !hgrant4_p & v372e669;
assign b08e51 = hgrant3_p & v3a69de7 | !hgrant3_p & v3a635ea;
assign v3a70433 = hmaster1_p & v376072e | !hmaster1_p & v3a702fc;
assign v377d745 = hmaster2_p & v373cc68 | !hmaster2_p & v3a6a609;
assign v376af6a = hbusreq4_p & v3a675f7 | !hbusreq4_p & v376bb26;
assign v372af91 = hbusreq1 & v372eaaf | !hbusreq1 & v377395f;
assign v374aa0f = hgrant5_p & v373b2ba | !hgrant5_p & !v8455ab;
assign v325c93e = hmaster2_p & v3739b80 | !hmaster2_p & !v3a60f71;
assign v37512c1 = hmaster0_p & v3a635ea | !hmaster0_p & v3763da5;
assign v375b04f = hgrant2_p & v3a6fbe2 | !hgrant2_p & v3755296;
assign v3a5749e = hmaster0_p & v3742582 | !hmaster0_p & v37384a3;
assign v375d8a6 = hmaster2_p & v3751004 | !hmaster2_p & v377de7b;
assign v377fbb9 = stateA1_p & v8455e1 | !stateA1_p & !v3a70df9;
assign v3741e61 = hbusreq7 & v3767059 | !hbusreq7 & v3a627a1;
assign v3731ffc = hlock3 & v3a6f3ad | !hlock3 & v3730946;
assign v376b1ee = hbusreq7 & v3764fd7 | !hbusreq7 & !v377a468;
assign v1e37368 = hmaster1_p & v374e855 | !hmaster1_p & v3756a59;
assign v3a63884 = hlock4 & v375cc06 | !hlock4 & v372d95c;
assign v372490a = hmaster0_p & v3a710f4 | !hmaster0_p & v3a634eb;
assign v372e96f = hbusreq4 & v3733c46 | !hbusreq4 & v8455ab;
assign v3a6f40a = hlock5_p & v3725612 | !hlock5_p & v8455ab;
assign v2acaef3 = hbusreq1 & v3a5600a | !hbusreq1 & v8455ab;
assign v3a6fe22 = hmaster2_p & v8455bb | !hmaster2_p & v376a96b;
assign v3a6f898 = hbusreq6 & v3a58b4c | !hbusreq6 & v3a6dc33;
assign v373e4ca = hbusreq8 & v37355e3 | !hbusreq8 & v3768734;
assign v37511a1 = hbusreq4_p & v3a5e55e | !hbusreq4_p & v372ac3b;
assign v3a59d40 = hbusreq3 & v3737d44 | !hbusreq3 & !v8455ab;
assign v376d21d = hmaster2_p & v3777adb | !hmaster2_p & v37751d9;
assign v3748ac8 = hbusreq5_p & v375121b | !hbusreq5_p & v37480b7;
assign v3a5a223 = hmaster2_p & v376c7d1 | !hmaster2_p & v3a70e98;
assign v3772007 = hmaster2_p & v3a707c4 | !hmaster2_p & v372cc25;
assign v3747630 = hgrant5_p & v8455ab | !hgrant5_p & v37366eb;
assign v3727d4d = hmaster2_p & v8455ab | !hmaster2_p & v37484de;
assign v377386a = hmaster1_p & v3a635ea | !hmaster1_p & v375d417;
assign v35b71af = hbusreq4 & v3a711d8 | !hbusreq4 & v8455ab;
assign v37740fd = hbusreq0 & v3a5c80e | !hbusreq0 & v377497c;
assign v3767adc = hbusreq0 & v37307dd | !hbusreq0 & v373e814;
assign v377bdec = hbusreq5 & v373e944 | !hbusreq5 & v3a64624;
assign v3a7162d = locked_p & v3a6ac94 | !locked_p & v8455ab;
assign v375bacc = hmaster2_p & v35772a6 | !hmaster2_p & v375a697;
assign v373f1a5 = hbusreq3 & v3a6f32f | !hbusreq3 & !v3a5614c;
assign v373e7d9 = hbusreq2 & v3809516 | !hbusreq2 & v376bade;
assign v3772200 = hmaster0_p & v374e0f6 | !hmaster0_p & !v37280f3;
assign v3a5b6ac = hmaster2_p & v37674f6 | !hmaster2_p & v8455ab;
assign v377c068 = hlock6 & v3a7118a | !hlock6 & v376d62b;
assign v3a6ffc0 = hbusreq5_p & v376156f | !hbusreq5_p & v3a5ba58;
assign v3771d2d = hgrant6_p & v37781ac | !hgrant6_p & v372f4f1;
assign v376a9f5 = hmaster1_p & v3a705ba | !hmaster1_p & v376055d;
assign v337859c = hbusreq3 & v37246f1 | !hbusreq3 & v3a70c74;
assign v37366b7 = hbusreq8_p & v375f8b1 | !hbusreq8_p & v374b86c;
assign v3a69f2b = hlock7_p & v3740a8a | !hlock7_p & v3a70652;
assign v376bb04 = hlock6_p & v374c5b2 | !hlock6_p & v8455bf;
assign v373c52e = hmaster1_p & v376bc32 | !hmaster1_p & v3a6f4da;
assign v3a71041 = hmaster1_p & v3779060 | !hmaster1_p & v3a695b7;
assign v3a6826d = hmaster0_p & v3764586 | !hmaster0_p & v3741dea;
assign v3779c40 = hbusreq8_p & v375dea9 | !hbusreq8_p & v3a58541;
assign v37693e7 = hmaster2_p & v3a62826 | !hmaster2_p & v8455ab;
assign v3a706dc = hmaster2_p & v8455ab | !hmaster2_p & v3a696ed;
assign v35b987f = hmaster0_p & v375fbf2 | !hmaster0_p & v374fda1;
assign v37642f9 = hbusreq6 & v3a63805 | !hbusreq6 & v8455ab;
assign v3a6f3dc = hbusreq7 & v3a6f371 | !hbusreq7 & v3a6d34c;
assign v3772b34 = hbusreq6_p & v3734067 | !hbusreq6_p & !v3a68b49;
assign v37573f5 = hmaster0_p & v3a6a56e | !hmaster0_p & v37527dc;
assign v375820e = hmaster2_p & v3773506 | !hmaster2_p & v8455ab;
assign v3760954 = hbusreq4_p & v3a712f2 | !hbusreq4_p & v374e345;
assign v3a55e7d = hlock1_p & v1e377bd | !hlock1_p & !v8455ab;
assign v376ba33 = hbusreq3_p & v3749ea2 | !hbusreq3_p & v3a6255b;
assign v3726f89 = hbusreq0 & v377623c | !hbusreq0 & !v8455ab;
assign v372be56 = hmaster2_p & v37757e0 | !hmaster2_p & v376ddc6;
assign v372f76a = hlock3 & v3741694 | !hlock3 & v39a4e5f;
assign v3758418 = hgrant6_p & v3a70240 | !hgrant6_p & v3a603cf;
assign v376b651 = hbusreq6 & v375ff74 | !hbusreq6 & !v8455ab;
assign v3a6fc84 = hbusreq7 & v3740f25 | !hbusreq7 & v3a56bb5;
assign v2093069 = hgrant7_p & v8455ab | !hgrant7_p & v3726c8e;
assign v373e6eb = hbusreq5 & ab808e | !hbusreq5 & v3771739;
assign v37640dc = hbusreq5 & v373f834 | !hbusreq5 & v3755d19;
assign v373df71 = hbusreq3 & v3763191 | !hbusreq3 & v35b774b;
assign v37679f0 = hbusreq7 & v37402b8 | !hbusreq7 & v3773ccd;
assign v3742f38 = stateG10_1_p & v8455ab | !stateG10_1_p & v3378a0a;
assign v3a6fb4e = jx0_p & v37496c6 | !jx0_p & b3ccfa;
assign v39a5265 = stateA1_p & v37295fe | !stateA1_p & !v3757c6f;
assign v376d387 = hburst0 & v376c211 | !hburst0 & v8455ab;
assign v374e753 = hgrant3_p & v372f657 | !hgrant3_p & v3a5fa18;
assign v3a5c3a0 = hgrant4_p & v373ff91 | !hgrant4_p & v3764702;
assign v372f853 = hgrant4_p & v3a6e543 | !hgrant4_p & v372b2aa;
assign v3759ee4 = hlock4 & v37657ef | !hlock4 & v3757f45;
assign v377432b = hbusreq5_p & v375a2a3 | !hbusreq5_p & v375b9cc;
assign v374bc9c = hmaster0_p & v372ddde | !hmaster0_p & v3a57912;
assign v3a6f0ed = hgrant6_p & v372aacd | !hgrant6_p & v1e379f7;
assign v39a4df7 = hmaster0_p & v373c6b6 | !hmaster0_p & v8455bd;
assign v3a6e138 = hgrant3_p & v8455be | !hgrant3_p & v375463f;
assign v3777d51 = hgrant5_p & v3752def | !hgrant5_p & v3a6f733;
assign v3a6db4b = hgrant1_p & v3778ed4 | !hgrant1_p & !v8455ab;
assign v3a6ec2a = hlock4_p & v37665bf | !hlock4_p & v3a6a939;
assign v3750fee = hlock5 & v3a62e92 | !hlock5 & v376e1fd;
assign v3744d60 = hmaster2_p & v3a7006c | !hmaster2_p & !v3759032;
assign v3a650a7 = hbusreq5_p & v3a6e005 | !hbusreq5_p & !v3a706c5;
assign v372ae9d = hbusreq6 & v360c3d7 | !hbusreq6 & !v8455ab;
assign v3766202 = hbusreq6_p & v3a6fbd4 | !hbusreq6_p & v8455ab;
assign v3a6f7a9 = hmaster3_p & v373ca17 | !hmaster3_p & v37505cd;
assign v39eb431 = hmaster2_p & v3a6b60d | !hmaster2_p & v375a1ab;
assign v375f3f4 = hbusreq4 & v3a6fa39 | !hbusreq4 & v8455ab;
assign v8f30ee = hbusreq3_p & v37528b9 | !hbusreq3_p & v376f911;
assign v3750382 = hbusreq8_p & v376419b | !hbusreq8_p & v8455ab;
assign v376dc91 = hbusreq4 & v376b11a | !hbusreq4 & v8455ab;
assign v373c983 = hgrant2_p & v3a710e1 | !hgrant2_p & v3a65ca8;
assign v3a70321 = hlock0_p & v376d327 | !hlock0_p & v373593a;
assign v3738c33 = hlock8_p & v3735ad7 | !hlock8_p & v3a6ed49;
assign v372ced7 = hmaster2_p & v3a57f59 | !hmaster2_p & v3733e9e;
assign d9fd79 = hbusreq8_p & v3735f03 | !hbusreq8_p & !v8455ab;
assign v3a6ffca = busreq_p & v373deb5 | !busreq_p & v3730dea;
assign v3a64b41 = hgrant3_p & v8455e7 | !hgrant3_p & !v3a70f04;
assign v372a9bd = hbusreq1_p & v3a6f6df | !hbusreq1_p & !v3a5a374;
assign v3a6ad22 = hmaster2_p & v8455ab | !hmaster2_p & v375f7d1;
assign v373c3e4 = hbusreq3 & v3a6500c | !hbusreq3 & v3726006;
assign v3a6f04d = hmaster2_p & v292555a | !hmaster2_p & v8455ab;
assign v3a6c6cf = hbusreq6 & v374e64f | !hbusreq6 & !v8455b9;
assign v372e132 = hlock2 & v2889703 | !hlock2 & v3a70923;
assign v375d78f = hbusreq5_p & v9fc6a0 | !hbusreq5_p & v373285d;
assign v37328fc = hbusreq6 & v3766b81 | !hbusreq6 & v3a5dcfc;
assign v3747114 = hbusreq0 & v3a58cd4 | !hbusreq0 & v3a6218f;
assign v3a56f67 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f061;
assign v3730595 = hmaster1_p & v372b4b4 | !hmaster1_p & v372dc39;
assign v3749655 = hbusreq0 & v375eeb0 | !hbusreq0 & v3726460;
assign v372c14d = hmaster2_p & v3a71250 | !hmaster2_p & v8455ab;
assign v374a0eb = hmaster2_p & v376a6f1 | !hmaster2_p & !v373c111;
assign v3a570ee = hmaster0_p & v373b02e | !hmaster0_p & v3a65069;
assign v3759dc9 = hbusreq7_p & v3753aa5 | !hbusreq7_p & v3a704d2;
assign v374d654 = hbusreq3 & v376b509 | !hbusreq3 & v3a5c1a5;
assign v3a6fdf0 = hgrant2_p & v8455ba | !hgrant2_p & v376d4b7;
assign v374a601 = jx0_p & v3722ba9 | !jx0_p & v3723bf9;
assign v373342f = hgrant2_p & v3a5e221 | !hgrant2_p & v373d506;
assign v37477d3 = hmaster0_p & v37640e9 | !hmaster0_p & v3a6fec8;
assign v3a70ee6 = hbusreq5 & v3730057 | !hbusreq5 & v376de5c;
assign v3a5d5cc = hgrant2_p & v3758472 | !hgrant2_p & !v374fd45;
assign v373ac1c = hgrant4_p & v8455ab | !hgrant4_p & v3a5efb8;
assign v3a6fd9c = hmaster1_p & v373016b | !hmaster1_p & v376c505;
assign v377320c = hbusreq3_p & v37675e2 | !hbusreq3_p & v375c806;
assign v374ea45 = hbusreq1_p & v373720a | !hbusreq1_p & v8455b0;
assign v3a6c91f = hbusreq0 & v3a6f579 | !hbusreq0 & v97f405;
assign v374c840 = hgrant4_p & v8455ab | !hgrant4_p & v3a62415;
assign stateG10_4 = !v379318f;
assign d9e2a4 = hmaster0_p & v8455ab | !hmaster0_p & v3773804;
assign v3766ce0 = hbusreq0 & v374b3cf | !hbusreq0 & !v8455ab;
assign v3a6c20e = hgrant4_p & v8455ab | !hgrant4_p & v3778546;
assign v3a64d60 = hbusreq2 & v8455b0 | !hbusreq2 & v3730ffe;
assign v3a710d9 = hlock0 & v3a6fdef | !hlock0 & v373d8f2;
assign v3a57658 = hbusreq4 & v3747bea | !hbusreq4 & v3a5e2e1;
assign v3739b80 = hbusreq6 & v37583be | !hbusreq6 & !v8455ab;
assign v3a714bf = hgrant6_p & v8455ab | !hgrant6_p & v3763898;
assign v3a70f11 = hgrant6_p & v8455ab | !hgrant6_p & !v37466c1;
assign v372ac64 = hmaster1_p & v3a5af94 | !hmaster1_p & v37232a3;
assign v375969d = hlock0_p & v3747302 | !hlock0_p & v3a648c3;
assign v3a705a9 = hbusreq0 & v3731a5a | !hbusreq0 & v3735112;
assign v37703a5 = hbusreq4_p & v3a70315 | !hbusreq4_p & v3a60258;
assign v374ad23 = hmaster1_p & v3759031 | !hmaster1_p & v37503c2;
assign v3770f55 = hlock0 & v375da82 | !hlock0 & v376af98;
assign v3a64361 = hbusreq5_p & v3a70642 | !hbusreq5_p & v3a6f932;
assign v374f0bf = hmaster2_p & v3773b23 | !hmaster2_p & v37685bb;
assign v3731e0f = hbusreq3 & v37244e7 | !hbusreq3 & v8455ab;
assign v3752ed7 = jx0_p & v3766597 | !jx0_p & v3a70a5f;
assign v37566c9 = hbusreq5 & v3779071 | !hbusreq5 & v377234d;
assign v37676b6 = jx1_p & v3761f13 | !jx1_p & v3a70a3d;
assign v373e450 = hbusreq4 & v3809e93 | !hbusreq4 & v3745f9b;
assign v3742dc6 = hbusreq2_p & v3a6f764 | !hbusreq2_p & v8455ab;
assign v3a6ef90 = hgrant6_p & v8455ab | !hgrant6_p & v373fef5;
assign v3a5e24d = hbusreq3 & v372dccf | !hbusreq3 & v3a69487;
assign v3a6b18c = hlock0 & v373031f | !hlock0 & v3a5f154;
assign v3a58db9 = hgrant6_p & v37571ad | !hgrant6_p & v3a7089f;
assign v373222d = hgrant4_p & v8455ab | !hgrant4_p & v3769945;
assign v3766c97 = hbusreq3_p & v377f730 | !hbusreq3_p & !v8455ab;
assign v3744aca = hmaster3_p & v3747462 | !hmaster3_p & v3775544;
assign v3a6847c = hlock6_p & v374ebb0 | !hlock6_p & v3a71350;
assign v3740af7 = hmaster1_p & v37469c4 | !hmaster1_p & v372dcc0;
assign v375af91 = hmaster1_p & v3a5ebc2 | !hmaster1_p & v3a6fb0e;
assign v3751929 = hbusreq7 & v3749f2e | !hbusreq7 & v377cbf0;
assign v3a5d5a4 = hbusreq4_p & v3729f25 | !hbusreq4_p & !v8455ab;
assign v372c06f = hgrant3_p & v8455be | !hgrant3_p & !v3a7065a;
assign v3761be0 = hgrant3_p & v377dd3b | !hgrant3_p & v3767d7c;
assign v3a71342 = hbusreq8_p & v372aafa | !hbusreq8_p & !v8455ab;
assign c88c38 = hlock4_p & v3770415 | !hlock4_p & v8455bb;
assign v376704f = hbusreq5_p & v37567ef | !hbusreq5_p & v375c062;
assign v3a706c7 = hbusreq1_p & v3a7148d | !hbusreq1_p & v3732b98;
assign v3a6c044 = hbusreq5 & v374a157 | !hbusreq5 & v3a5e783;
assign v373481c = hbusreq6_p & v3a6a880 | !hbusreq6_p & v8455b3;
assign v3733cfb = hmaster0_p & v3a6f8be | !hmaster0_p & v377b6ce;
assign v3773b30 = hmaster2_p & v8455e7 | !hmaster2_p & v35772c9;
assign v3a69169 = hgrant4_p & v8455ab | !hgrant4_p & v373c2d7;
assign v3736739 = hgrant6_p & v3748a4f | !hgrant6_p & v3a70e86;
assign v3758cf5 = hbusreq4_p & v3739d88 | !hbusreq4_p & v373f6ee;
assign v3778834 = hlock3_p & v377f01a | !hlock3_p & v37373ea;
assign v37698ab = hbusreq7_p & v3760233 | !hbusreq7_p & v3764238;
assign v373f53e = hbusreq5_p & v3744aaa | !hbusreq5_p & !v8455ab;
assign v3741759 = hgrant5_p & v376139f | !hgrant5_p & v3747210;
assign v373cfbd = hmaster2_p & v372ba1c | !hmaster2_p & v3769740;
assign c7f8d6 = hlock0_p & v376f73c | !hlock0_p & !v373cff4;
assign v376d0bc = hmaster2_p & v375ed6f | !hmaster2_p & v3a6f99c;
assign v3735236 = hbusreq5_p & v3725a21 | !hbusreq5_p & v3736b43;
assign v3a672c8 = hmaster2_p & v377accc | !hmaster2_p & v3a6fa93;
assign v3727626 = hmaster1_p & v37358d5 | !hmaster1_p & v3a62424;
assign v3a6aac8 = hmaster0_p & v3a70ca4 | !hmaster0_p & v3806882;
assign v3727c6e = hmaster1_p & v377d1dc | !hmaster1_p & v3a6f728;
assign v377981b = hbusreq8 & v3762892 | !hbusreq8 & v375a510;
assign v37579b8 = hmaster2_p & v3a6fcba | !hmaster2_p & !v374044c;
assign v37538e1 = hbusreq0_p & v3747302 | !hbusreq0_p & v3a6c5ee;
assign v374d8bb = hlock2 & v375b261 | !hlock2 & v29256bb;
assign v373e76c = hmaster1_p & v3a6e8b1 | !hmaster1_p & v3a6f89b;
assign v3761e62 = hmaster2_p & v35772a6 | !hmaster2_p & v3728dc7;
assign v373af26 = hlock5 & v3a6799d | !hlock5 & v3761d9f;
assign v3a55954 = hgrant2_p & v8455ba | !hgrant2_p & v3726a2c;
assign v3a70a8f = hlock4 & v3768eac | !hlock4 & v3a7001d;
assign v3736948 = jx0_p & v3a7157f | !jx0_p & v372363e;
assign v380651a = hmaster1_p & v3a6f92f | !hmaster1_p & v3a5a1e8;
assign v3724b26 = hmaster1_p & v3a67ffd | !hmaster1_p & v37324da;
assign v3736df1 = hmaster1_p & v3749ba6 | !hmaster1_p & v375a311;
assign v3777bf9 = hbusreq0 & v375d1d9 | !hbusreq0 & v3a7129b;
assign v37297b2 = hgrant6_p & v37711cc | !hgrant6_p & v3776be1;
assign v3a71502 = hmaster2_p & v2ff9190 | !hmaster2_p & v8455ab;
assign v3a70e16 = hlock5 & v3748966 | !hlock5 & v3743ec6;
assign v3a5be20 = hbusreq2_p & v37583be | !hbusreq2_p & v373fda2;
assign v37629db = hgrant7_p & v8455ab | !hgrant7_p & v3a689b8;
assign v3761d2f = hbusreq5_p & v3758fa8 | !hbusreq5_p & v1e37b76;
assign v3a53a2d = hmaster2_p & v3a706fe | !hmaster2_p & v3722bca;
assign v2678c97 = hbusreq4_p & v3739ab6 | !hbusreq4_p & v3760309;
assign v3809a8b = hgrant2_p & v3a7031f | !hgrant2_p & v3a635ea;
assign v372e873 = hlock0 & v375da82 | !hlock0 & v3a6f4af;
assign v373ed9a = hlock2 & v375b736 | !hlock2 & v375767e;
assign v3a6ff04 = hmaster1_p & v3807f45 | !hmaster1_p & v3766803;
assign v376dfed = hlock0_p & v3a68c1f | !hlock0_p & !v3a5e357;
assign v37519ed = stateG10_1_p & v8455e1 | !stateG10_1_p & !v3763cf5;
assign v374e78a = hmaster0_p & v8455ab | !hmaster0_p & v3a5c538;
assign v3a5a93a = hlock0 & v373abde | !hlock0 & v3a627b3;
assign v377f06c = hmaster0_p & v8455ab | !hmaster0_p & v373ea29;
assign v3728fcd = hmaster2_p & v3a6c4e4 | !hmaster2_p & v375139d;
assign v3740d05 = hmaster0_p & v3760512 | !hmaster0_p & v3a710c3;
assign v3760d53 = hlock4_p & v377de7b | !hlock4_p & v375d616;
assign v3a6dd7e = hbusreq4 & v3a5b8e4 | !hbusreq4 & v3a70c74;
assign c86567 = hmaster2_p & v3a635ea | !hmaster2_p & v376e90a;
assign v3a70015 = hmaster1_p & v3777498 | !hmaster1_p & v3751606;
assign v3a648f6 = hbusreq7_p & v1e37ec1 | !hbusreq7_p & v3a60276;
assign v374fc8e = hbusreq2_p & v376b4e1 | !hbusreq2_p & v3723efc;
assign v913004 = hmaster0_p & v3a6a63c | !hmaster0_p & !v3a700a8;
assign v3a53cc3 = stateG10_1_p & v375bbe9 | !stateG10_1_p & v3a5fe1d;
assign v372d7a4 = hlock2 & v372d608 | !hlock2 & v37288b6;
assign v3a6f8e1 = hmaster1_p & v3758bfe | !hmaster1_p & v3740bf5;
assign v374d31a = hbusreq8 & v374c576 | !hbusreq8 & v3736684;
assign v377a883 = hbusreq8_p & v3a5bc5d | !hbusreq8_p & v3a70a97;
assign v37469c4 = hgrant4_p & v3772d6e | !hgrant4_p & v3748f09;
assign v3a70e53 = hbusreq7_p & v3a56c18 | !hbusreq7_p & v37673e8;
assign v3a6a084 = hlock7 & v377fbeb | !hlock7 & v3a64dbb;
assign ae0781 = hlock2 & v3a70715 | !hlock2 & v3a61cbf;
assign v376ab29 = hmaster0_p & v376bd43 | !hmaster0_p & v375cc17;
assign v3764c57 = hgrant6_p & v3743eae | !hgrant6_p & v3761bb6;
assign v3767e79 = hmaster0_p & v3a70950 | !hmaster0_p & v3a57912;
assign v3a6261f = hgrant8_p & v3a67131 | !hgrant8_p & !v374dddd;
assign v3a6512b = hlock4 & v3a6cb62 | !hlock4 & v3a5b4de;
assign v3a703f2 = hgrant4_p & v3a6ffb6 | !hgrant4_p & v3a701ab;
assign v3a70acb = hbusreq7_p & a0a219 | !hbusreq7_p & v376f92f;
assign v376142a = hgrant4_p & v8455ab | !hgrant4_p & v374a3b2;
assign v373f42f = hlock4_p & v373146d | !hlock4_p & v3a6f4ec;
assign v3775bca = hbusreq6 & v3a5cebe | !hbusreq6 & v8455ab;
assign v37278c2 = hbusreq2_p & v3a6ffe5 | !hbusreq2_p & v3763acf;
assign v3a66306 = hlock4 & v3a6fa55 | !hlock4 & v374b320;
assign v372cb44 = hgrant6_p & v8455ab | !hgrant6_p & v95151c;
assign v3775e78 = hlock4 & v3a62197 | !hlock4 & v3743c51;
assign v376766e = jx0_p & v3776ce3 | !jx0_p & v8455ab;
assign v37261a6 = hbusreq8_p & v376f0c2 | !hbusreq8_p & b412f3;
assign v3737438 = hbusreq8_p & dacf90 | !hbusreq8_p & v3a6eef0;
assign v3a62615 = hgrant8_p & v3773e52 | !hgrant8_p & v3729c71;
assign v3a6f249 = hmaster2_p & v3a58218 | !hmaster2_p & v3a6dc08;
assign v373046c = hbusreq8 & v3a6856a | !hbusreq8 & v373ba84;
assign v375b3be = hlock0 & v38072fd | !hlock0 & v3a704de;
assign v373f953 = hbusreq6 & v3a582d6 | !hbusreq6 & v376e041;
assign v377803f = hbusreq2_p & v8455ab | !hbusreq2_p & v8455bd;
assign v3a6fb68 = hbusreq4_p & v37541a7 | !hbusreq4_p & v3727084;
assign v3a711e5 = hmaster2_p & v373899b | !hmaster2_p & v3a6b6ef;
assign v39a536d = hbusreq3 & v3a6143b | !hbusreq3 & !v8455b5;
assign v3a6f8fd = hlock4 & v377f70a | !hlock4 & v3a6134b;
assign v3a69efa = hbusreq6 & v375b044 | !hbusreq6 & v373f0ee;
assign v374f511 = hbusreq6_p & v3a6f9bc | !hbusreq6_p & v35772a6;
assign v3a6fd0a = hmaster2_p & v20930c6 | !hmaster2_p & v3767f7f;
assign v3a6f5f6 = hgrant3_p & v3744ca2 | !hgrant3_p & !v3a64e91;
assign v3761781 = hgrant5_p & v8455ab | !hgrant5_p & v376b035;
assign v377c72c = hmaster3_p & v3746d92 | !hmaster3_p & v37419f2;
assign v373ead4 = hgrant1_p & v3767abc | !hgrant1_p & v3735ed0;
assign v3770f76 = hlock5_p & v3a6c179 | !hlock5_p & v373285d;
assign v373acce = hbusreq2 & v39a4ca8 | !hbusreq2 & v8455b5;
assign v3a6c849 = hbusreq8_p & v377e871 | !hbusreq8_p & v3756e63;
assign v3a6f723 = hgrant4_p & v8455ab | !hgrant4_p & v3768364;
assign v3a70e0e = hbusreq5_p & v3a70924 | !hbusreq5_p & !v8455ab;
assign b4ede7 = hmaster3_p & v3a6f53e | !hmaster3_p & v3a66a4f;
assign v3a6670c = hbusreq6 & v3733334 | !hbusreq6 & v391331d;
assign v3773107 = hmaster0_p & v8455ab | !hmaster0_p & !v37794e5;
assign v3a53dbb = hgrant4_p & v8455ab | !hgrant4_p & !v3a713dd;
assign v3a6a8b2 = hgrant5_p & v3a706ea | !hgrant5_p & v377c236;
assign v374bbca = jx1_p & v376964c | !jx1_p & v3a5d930;
assign v360d0a7 = hlock0_p & v3737462 | !hlock0_p & v3a5d34b;
assign v3a5b289 = hlock2_p & v3a6ffca | !hlock2_p & !v8455ab;
assign v3a682e5 = hbusreq7_p & v3778627 | !hbusreq7_p & v3a5e998;
assign v37483ff = hgrant4_p & v8455ab | !hgrant4_p & v3a572b4;
assign v3a7101b = hbusreq1_p & v372fca8 | !hbusreq1_p & !v8455ab;
assign v3a62542 = hgrant4_p & v3a5c945 | !hgrant4_p & v374c53a;
assign v3a7038d = jx3_p & v3a5f375 | !jx3_p & !v3a6de5e;
assign v3a6f32d = hbusreq4_p & be0bbd | !hbusreq4_p & v35772a6;
assign v3752428 = hbusreq5_p & v9af7ec | !hbusreq5_p & v3779680;
assign v3779cb5 = hbusreq7_p & v373aaf0 | !hbusreq7_p & v8455ab;
assign v3a714fd = hbusreq4_p & v3a70e0f | !hbusreq4_p & !v8455ab;
assign v3736f6d = hbusreq7 & v944e42 | !hbusreq7 & v3750bc4;
assign v3a64483 = hmaster0_p & v37771ed | !hmaster0_p & v375d77d;
assign v372a8d9 = jx0_p & v3736c86 | !jx0_p & v3743b49;
assign v3a704d5 = hlock6_p & v3a66750 | !hlock6_p & v3759daf;
assign v3a55bd0 = hbusreq6_p & v3763a20 | !hbusreq6_p & v374c163;
assign v375e682 = hbusreq6_p & v8455b0 | !hbusreq6_p & v3753dab;
assign v39ed7ea = decide_p & v3a71352 | !decide_p & v3742ed3;
assign v3764f60 = hmaster2_p & v23fdd06 | !hmaster2_p & v3726605;
assign v37600ad = jx0_p & v374c009 | !jx0_p & v3772616;
assign v3726bcc = hmaster2_p & v377c7c0 | !hmaster2_p & v3724e8e;
assign v3741b59 = hmaster2_p & v3a6f240 | !hmaster2_p & v3766ce0;
assign v3741b5e = hmaster2_p & v8455ab | !hmaster2_p & v376d306;
assign v3733e0a = hlock4_p & v3752577 | !hlock4_p & v377c34f;
assign v372865e = hgrant1_p & v3722e5c | !hgrant1_p & v35772a6;
assign v376513c = hgrant6_p & v8455ab | !hgrant6_p & v9a07a5;
assign v3743546 = hbusreq6 & v377af44 | !hbusreq6 & v8455ab;
assign v3a5551b = hmaster1_p & v3a6fc0f | !hmaster1_p & v372b3ca;
assign v376ddc6 = hbusreq1_p & v3a620e2 | !hbusreq1_p & v8455b0;
assign v3a59b6d = hmaster1_p & v3a6ebe2 | !hmaster1_p & v8455ab;
assign v3778d73 = hmaster2_p & v3771076 | !hmaster2_p & v3a6fc7f;
assign v3a65b64 = hbusreq7_p & v376a3cb | !hbusreq7_p & v37581d2;
assign v3771fec = hmaster0_p & v3755002 | !hmaster0_p & v3a70116;
assign v372cafb = hlock5_p & v3760e6e | !hlock5_p & !v374fad5;
assign v3a714da = hmaster1_p & v375a858 | !hmaster1_p & v374a9eb;
assign v3a6f3ee = hbusreq4_p & v37707d5 | !hbusreq4_p & v3a6faef;
assign v372a85f = hgrant4_p & v3725717 | !hgrant4_p & v3a69c57;
assign v374a849 = hmaster1_p & v377a6bf | !hmaster1_p & v3a60247;
assign v3a67fc6 = hbusreq7 & v3a62cb5 | !hbusreq7 & v3a5c3c4;
assign v3a70f45 = hmaster2_p & v3779680 | !hmaster2_p & v377308e;
assign v3a715b0 = hbusreq3_p & v3a70d67 | !hbusreq3_p & !v8455ab;
assign v3730b98 = hgrant4_p & v8455ab | !hgrant4_p & v3730e90;
assign v3a711d5 = hmaster1_p & v23fe20c | !hmaster1_p & v3a569c8;
assign v375a95b = hgrant4_p & v372b268 | !hgrant4_p & v3755a02;
assign v1e37a04 = hgrant2_p & v8455ab | !hgrant2_p & v3776c44;
assign v91ebb9 = hmaster0_p & v8455ab | !hmaster0_p & v3768a3c;
assign v3725bea = hgrant2_p & v3726139 | !hgrant2_p & v375bdf0;
assign v3a6ebc6 = hmaster1_p & v8455ab | !hmaster1_p & v3a7094b;
assign v373c8cb = hbusreq4 & v37302f1 | !hbusreq4 & !v8455bd;
assign v37598a3 = hbusreq2 & v3723b00 | !hbusreq2 & v8455ab;
assign v374e6a5 = hbusreq2_p & v3a635ea | !hbusreq2_p & v3739e39;
assign v3a6ab7f = hmaster2_p & v3751d7d | !hmaster2_p & v3a715d2;
assign v373f1db = hmaster2_p & v37666f6 | !hmaster2_p & !v8455ab;
assign v98381a = hbusreq4 & v3755a70 | !hbusreq4 & v3a7164a;
assign v375cd00 = hgrant6_p & v3743ded | !hgrant6_p & v3a70055;
assign v376beed = hgrant6_p & v8455ab | !hgrant6_p & v3a5d836;
assign v3a71164 = hbusreq3_p & v3760933 | !hbusreq3_p & v8455ab;
assign v37672ac = hbusreq3_p & v3730181 | !hbusreq3_p & v8455ab;
assign v3a58c07 = hmaster0_p & v8455b0 | !hmaster0_p & v3a6a56e;
assign v3a6a7b4 = hgrant3_p & v3777d79 | !hgrant3_p & v1e3825d;
assign v37375bc = hbusreq2_p & v3753f37 | !hbusreq2_p & !v8455ab;
assign v373a6c8 = hlock6 & v3a6872e | !hlock6 & v3725556;
assign v375c1c5 = hmaster2_p & v39a4dbb | !hmaster2_p & !v3748609;
assign v37582dc = hmaster2_p & v3722e5c | !hmaster2_p & v3a6eb39;
assign v3a5be6a = hgrant2_p & v8455ab | !hgrant2_p & bf6063;
assign v3a6c39b = hbusreq4 & v3a6f993 | !hbusreq4 & v8455ab;
assign v3768aa4 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3a5e2b9;
assign v3a682f0 = hbusreq0 & v8455b0 | !hbusreq0 & v3a6f0bd;
assign v3809e93 = hlock6 & v3a6b90f | !hlock6 & v3a5bca4;
assign v3a593cc = hbusreq8 & v3756546 | !hbusreq8 & v373496c;
assign v3a668a4 = hbusreq4 & v3a7156d | !hbusreq4 & v8455ab;
assign v3767d57 = hmaster2_p & v3a55198 | !hmaster2_p & v8455ab;
assign v3a58218 = hlock0_p & v373cca3 | !hlock0_p & !v8455ab;
assign v3a57156 = hbusreq0 & v3734c7e | !hbusreq0 & v8455ab;
assign v374ca02 = hmaster0_p & v3a71073 | !hmaster0_p & v8455ab;
assign v372d078 = hbusreq3_p & v3a635ea | !hbusreq3_p & v3a6ef1e;
assign v376d93b = hmaster2_p & v3a5c3a0 | !hmaster2_p & v375a1ab;
assign v3761c19 = hmaster0_p & v374729b | !hmaster0_p & v3a6f0c8;
assign v375f98a = hbusreq2_p & v37406d2 | !hbusreq2_p & v3753dab;
assign v3776a59 = hmaster0_p & v3751891 | !hmaster0_p & v3a58b9f;
assign v37582a2 = hmaster0_p & v3a6dfdb | !hmaster0_p & v3758c58;
assign v3757b0e = hgrant2_p & v3a57f59 | !hgrant2_p & v3766709;
assign v3760198 = hgrant7_p & v8455ab | !hgrant7_p & !v376a966;
assign v375bb15 = hgrant6_p & v8455ab | !hgrant6_p & v3a70178;
assign v3731d8f = hmaster0_p & v3a635ea | !hmaster0_p & v3743fba;
assign v3731e3c = stateG3_1_p & v845601 | !stateG3_1_p & v8455ab;
assign v37600da = hbusreq4_p & v3737dad | !hbusreq4_p & v3774a1e;
assign v373a341 = hbusreq6_p & v3a635ea | !hbusreq6_p & v3a641d5;
assign v337904e = hgrant1_p & v37470eb | !hgrant1_p & !v8455e7;
assign v38079c2 = hbusreq7_p & v3a6f680 | !hbusreq7_p & v3a6d89d;
assign v3732772 = hmaster2_p & v3a6ffca | !hmaster2_p & v3a71484;
assign v375e0e3 = hbusreq6_p & v3a68f98 | !hbusreq6_p & v3748d67;
assign v3808c39 = hlock0_p & v374f87c | !hlock0_p & v8455b0;
assign v377047a = hgrant4_p & v375058e | !hgrant4_p & v3a68fd3;
assign v3a70452 = hgrant0_p & v8455ab | !hgrant0_p & v375d8fb;
assign v373cd0a = hbusreq0 & v3753073 | !hbusreq0 & v3a706d2;
assign v37b64f8 = hlock5_p & v373d199 | !hlock5_p & !v3757ca4;
assign v373d0eb = hbusreq8_p & v894fb9 | !hbusreq8_p & v374071d;
assign v3775f56 = hmaster0_p & v3740b82 | !hmaster0_p & v374b1a4;
assign cf1ae7 = hbusreq3 & v37406d2 | !hbusreq3 & v8455ab;
assign v3748b0e = hmaster0_p & v3753883 | !hmaster0_p & !c04cff;
assign v3a6279b = hmaster2_p & v8455ab | !hmaster2_p & v3728c08;
assign v3744d2a = hbusreq5 & v3751d33 | !hbusreq5 & v3a6f5d4;
assign v3748984 = hmaster1_p & v3a619c0 | !hmaster1_p & v3a6fde5;
assign v3774ad3 = hburst0 & v3a563ad | !hburst0 & !v8455ab;
assign v37661dc = hbusreq5 & v3a6ef30 | !hbusreq5 & !v3769ca2;
assign v3a6efd1 = hgrant0_p & v8455e7 | !hgrant0_p & !v374063d;
assign v3733734 = hgrant6_p & v8455ab | !hgrant6_p & v3737193;
assign v3735c51 = hbusreq3_p & v3a712e7 | !hbusreq3_p & v8455b3;
assign v3a68904 = hmaster0_p & v3a6f4df | !hmaster0_p & v3770da3;
assign v375c69e = hburst0 & v39a537f | !hburst0 & v372dd8e;
assign v37482c8 = hbusreq3 & v3729ae4 | !hbusreq3 & v8455ab;
assign v374c47e = hbusreq2 & v374f307 | !hbusreq2 & v8455b0;
assign v3734a92 = hbusreq4_p & v374ab4f | !hbusreq4_p & v374fe0f;
assign v375cc28 = hbusreq3_p & v3a70910 | !hbusreq3_p & v3a70452;
assign v374d47d = hbusreq4_p & v3a708ad | !hbusreq4_p & v37307d7;
assign v37612dd = hgrant6_p & v372a51d | !hgrant6_p & v3808ee4;
assign v375e9ca = hmaster1_p & v3a635ea | !hmaster1_p & v372e571;
assign v3a6fdbd = hmaster2_p & v377f734 | !hmaster2_p & v3a71555;
assign v377d714 = hbusreq6 & v3a6dc08 | !hbusreq6 & v37406d2;
assign v3a55bd3 = hlock5_p & v3779477 | !hlock5_p & v37494ce;
assign v372e83a = jx0_p & v372bce5 | !jx0_p & v3773ad7;
assign v377601b = hmaster1_p & v39ea76e | !hmaster1_p & v377ea6c;
assign v37510fb = hmaster0_p & v3a6669b | !hmaster0_p & v375355a;
assign v3773ee6 = hlock0_p & v8455ab | !hlock0_p & v8455e7;
assign v372348f = hbusreq5_p & v374d525 | !hbusreq5_p & v3a60836;
assign v372a309 = hbusreq5 & v37345de | !hbusreq5 & v377de7f;
assign v373f4d3 = stateG2_p & v8455ab | !stateG2_p & v37464c8;
assign v3a6f549 = hbusreq3_p & v8455e1 | !hbusreq3_p & v3744f35;
assign v376d4f3 = hbusreq5_p & v377672d | !hbusreq5_p & v3a70556;
assign v372d86a = hgrant6_p & v3752a0d | !hgrant6_p & v376c13c;
assign v373d8e5 = hgrant0_p & v8455ab | !hgrant0_p & v3726d00;
assign v37266c6 = hgrant6_p & v3739761 | !hgrant6_p & v372ac03;
assign v3a667ba = hmaster0_p & v3a5fc61 | !hmaster0_p & v377a083;
assign v37267f3 = hmaster0_p & v3756a9e | !hmaster0_p & v374eaf4;
assign v3a6fad9 = hlock3 & v3748797 | !hlock3 & v376d34b;
assign v37520fc = hmaster2_p & v8455ab | !hmaster2_p & v3738d63;
assign v3a6eb1b = hbusreq4 & v3769112 | !hbusreq4 & v3748797;
assign v375e721 = hgrant4_p & v3728c23 | !hgrant4_p & v373d735;
assign v376faa6 = hlock7_p & v373c82f | !hlock7_p & v3743ab6;
assign v3725c41 = hmaster2_p & v3a635ea | !hmaster2_p & v3723fcc;
assign v3a70a18 = hlock4 & v3a6ead6 | !hlock4 & v3a70a4d;
assign v377fb50 = hmaster1_p & v374743d | !hmaster1_p & v3723e2f;
assign v3738ff9 = hgrant6_p & v3a71389 | !hgrant6_p & v3a5f41d;
assign b3a152 = hmaster0_p & v3765c70 | !hmaster0_p & !v37733e3;
assign v3a700eb = hmaster0_p & v374aabf | !hmaster0_p & v3a5bd69;
assign v374dcfb = hmaster0_p & v8455ab | !hmaster0_p & !v372eb00;
assign v375c381 = hbusreq5_p & v3a6ffc1 | !hbusreq5_p & v3a713ad;
assign v3a6c03d = hmaster2_p & v374c78e | !hmaster2_p & v3730b98;
assign v375058e = hbusreq4_p & v8455ab | !hbusreq4_p & v375564e;
assign v3a6f5a0 = hbusreq4 & v3a6fc2f | !hbusreq4 & v2092abe;
assign v3725580 = hgrant4_p & v377a036 | !hgrant4_p & v376e844;
assign v377a7f8 = hmaster2_p & v37234c3 | !hmaster2_p & !v3729f14;
assign v3a5bc70 = jx1_p & v3a6f274 | !jx1_p & v373cdef;
assign v376aa10 = hbusreq4 & v3a6f8f5 | !hbusreq4 & v8455bf;
assign v3769bcb = hbusreq2_p & v3747302 | !hbusreq2_p & v3725506;
assign v3722e49 = hbusreq8 & v3a6f578 | !hbusreq8 & v8455ab;
assign v3a6ec22 = hbusreq5_p & v3755d20 | !hbusreq5_p & v3750f27;
assign v372d299 = hbusreq4_p & v3a635ea | !hbusreq4_p & v3a63621;
assign v37502d9 = hbusreq3 & v3a6c23b | !hbusreq3 & v3a70cdb;
assign v3747b02 = hlock5_p & v3740f65 | !hlock5_p & v3a6826d;
assign v3a5b6ca = hbusreq3_p & v3758c62 | !hbusreq3_p & v37355db;
assign v3a715e2 = hbusreq2 & v3725410 | !hbusreq2 & v3a706d1;
assign v3a6b3df = hbusreq2_p & v3759cce | !hbusreq2_p & v8455b0;
assign v3774fa6 = hgrant6_p & v8455ca | !hgrant6_p & v3a64f97;
assign v3732128 = hbusreq3_p & v3752fe9 | !hbusreq3_p & !v8455ab;
assign v1e37c60 = hlock5 & v3747b97 | !hlock5 & v3a6e81d;
assign v3730b6d = hgrant3_p & v8455ab | !hgrant3_p & v3a5eb73;
assign v3a6be79 = hmaster2_p & v3724c55 | !hmaster2_p & v3a607af;
assign v3809e77 = hgrant5_p & v8455ab | !hgrant5_p & v3761719;
assign v3754a27 = hgrant3_p & v3a5c5ca | !hgrant3_p & v3761224;
assign c8ca6f = hmaster1_p & v3a57f59 | !hmaster1_p & v3760e6e;
assign v3a6eeef = hbusreq2_p & v3745eab | !hbusreq2_p & v8455ab;
assign v3a5b03b = hbusreq7_p & v3767a08 | !hbusreq7_p & v3a71333;
assign v37483f9 = hmaster2_p & v373ad2b | !hmaster2_p & v3a67869;
assign v3a6f173 = hmaster0_p & v37781b7 | !hmaster0_p & v3731079;
assign v37533e5 = hmaster1_p & v373d27f | !hmaster1_p & v39ebb7b;
assign v3743393 = hbusreq6_p & v3a6bf6d | !hbusreq6_p & v3756b48;
assign v375356f = hgrant1_p & v8455ab | !hgrant1_p & v3747c3e;
assign v3a70fd2 = hlock2 & v3a6f418 | !hlock2 & v3a5cf53;
assign v3725bab = hbusreq4 & v3a6a493 | !hbusreq4 & v3a70ad6;
assign v3743702 = hbusreq6_p & v3735134 | !hbusreq6_p & v89c52e;
assign v37295fe = hmastlock_p & v3a70b47 | !hmastlock_p & !v8455ab;
assign v377329c = hbusreq4_p & v3a53cf5 | !hbusreq4_p & !v8455ab;
assign v3a60c4f = hmaster2_p & v3a5c562 | !hmaster2_p & v3727e66;
assign v37317ec = hmaster2_p & v376111d | !hmaster2_p & !v23fe324;
assign v3a705ae = hbusreq5 & v3a70fc4 | !hbusreq5 & v3766cfb;
assign v3762312 = hgrant6_p & v3a654c1 | !hgrant6_p & v3a6ffff;
assign v337793f = hlock1_p & v372ef7c | !hlock1_p & !v8455ab;
assign v3730be2 = hbusreq4 & v3a6f7bf | !hbusreq4 & v8455ab;
assign v376d191 = hbusreq7_p & v374e7b5 | !hbusreq7_p & v3724b26;
assign v3751d30 = hlock4_p & v3a6f5ea | !hlock4_p & v37406d2;
assign v3772a15 = hmaster1_p & v9375a3 | !hmaster1_p & v374e21e;
assign v3a6eab3 = hgrant3_p & v37579a9 | !hgrant3_p & v372e92b;
assign v372c959 = hmaster3_p & v8455ab | !hmaster3_p & v374c556;
assign v3a6d6be = hbusreq0 & v3a6f9e5 | !hbusreq0 & v3761bb7;
assign v3a5e371 = hmaster2_p & v3a6898d | !hmaster2_p & v3a66316;
assign v3a706ed = hlock6 & v2093234 | !hlock6 & v3744f0d;
assign v3731994 = hlock5 & v3755207 | !hlock5 & v3a6329a;
assign v373be4d = jx1_p & v8a1014 | !jx1_p & v373eb05;
assign v3a706b3 = hbusreq5 & v3a5e1e4 | !hbusreq5 & v8455e7;
assign v3a6f3ab = hlock2_p & v9c492b | !hlock2_p & v8455e7;
assign v376de4e = hbusreq3_p & v3a6fac5 | !hbusreq3_p & v8455ab;
assign v3a5deb7 = locked_p & v8455ab | !locked_p & !v373c3bd;
assign v373c0b4 = hbusreq7 & v3a5fa29 | !hbusreq7 & v375a510;
assign v37536b2 = hbusreq5 & v373014d | !hbusreq5 & v8455bf;
assign v3a554d8 = hmaster2_p & v8455ab | !hmaster2_p & v3a6b873;
assign v376778a = hbusreq8_p & v377073f | !hbusreq8_p & v3a6c15d;
assign v3729b52 = hmaster0_p & v372b902 | !hmaster0_p & v3a59979;
assign v3a6f19d = hmaster1_p & v37586d3 | !hmaster1_p & v3a63812;
assign v3762fdb = hmaster0_p & v3735fe8 | !hmaster0_p & v8455ab;
assign v3743788 = hbusreq5_p & v3752798 | !hbusreq5_p & v39eaa60;
assign v376fe7d = hmaster1_p & v375a64f | !hmaster1_p & v8455ab;
assign v375b1a0 = hbusreq5 & v3a6f810 | !hbusreq5 & v37551b8;
assign v37361ad = hbusreq8_p & v3765e47 | !hbusreq8_p & !v8455ab;
assign v3778d7f = hmaster2_p & v3723b5b | !hmaster2_p & v37697a3;
assign v3a6f409 = hmaster3_p & v3a558dc | !hmaster3_p & v8455ab;
assign v372b22b = hgrant2_p & v375d38f | !hgrant2_p & !v3a5927f;
assign v3a7092a = hbusreq1_p & v3a5e9a3 | !hbusreq1_p & !v8455ab;
assign v376a2bf = hlock2 & v3a6fea8 | !hlock2 & v372b373;
assign v375f2a3 = hbusreq5_p & v37306c6 | !hbusreq5_p & v3773eeb;
assign v39a4ca8 = hbusreq1_p & v3a6254e | !hbusreq1_p & !v8455ab;
assign v372b9c6 = hbusreq3_p & v2092ffc | !hbusreq3_p & v3765ce2;
assign v375fec7 = hlock6_p & v8455ab | !hlock6_p & v3a70a05;
assign v372faf3 = hbusreq5_p & v38076cf | !hbusreq5_p & v376142a;
assign v38072f9 = hgrant6_p & v8455ab | !hgrant6_p & v376bf0a;
assign v372bd46 = hbusreq5_p & v3a6eb67 | !hbusreq5_p & v37790c8;
assign v3a6f37d = hmaster1_p & v37787ac | !hmaster1_p & v3a65388;
assign v3378f4c = hgrant2_p & v8455ba | !hgrant2_p & v373301d;
assign v37780f6 = hgrant3_p & v376e7bc | !hgrant3_p & v374e03d;
assign v3a70592 = hmaster0_p & v3750ea5 | !hmaster0_p & v3a708a7;
assign v3a5750b = hbusreq5 & v3a6caa7 | !hbusreq5 & v3731720;
assign v3a6eb0d = hmaster0_p & v372d905 | !hmaster0_p & v8455e7;
assign v377d521 = hgrant5_p & v8455c6 | !hgrant5_p & v3745614;
assign v3a71149 = hmaster0_p & v374f658 | !hmaster0_p & v3723988;
assign v376efb6 = hlock0 & v3730695 | !hlock0 & v3741ccb;
assign v37565b0 = hmaster2_p & v3a70f68 | !hmaster2_p & v3765511;
assign v3777a52 = hbusreq6 & v3a6f496 | !hbusreq6 & v3a69487;
assign v3a5f315 = hgrant2_p & v375d288 | !hgrant2_p & v3745484;
assign v3a5971d = hbusreq8_p & v37646ce | !hbusreq8_p & v3a6724f;
assign v3733278 = hbusreq2_p & v377d254 | !hbusreq2_p & !v8455ab;
assign v373e48c = hbusreq5_p & v372523e | !hbusreq5_p & v8455ab;
assign v3a563ad = stateA1_p & v8455ab | !stateA1_p & v3745b85;
assign v3a59979 = hmaster2_p & v372b902 | !hmaster2_p & v380760a;
assign v380663a = hlock6_p & v3a703fc | !hlock6_p & !v8455ab;
assign v37385ee = hlock5_p & v3a7124d | !hlock5_p & !v3a678de;
assign v37445a8 = hmaster2_p & v9f823e | !hmaster2_p & v37314fa;
assign v377cc52 = hmaster2_p & v9ed516 | !hmaster2_p & v3730e2a;
assign v372fc51 = locked_p & v377b24b | !locked_p & v3577306;
assign v3a684ef = hgrant0_p & v3a5880b | !hgrant0_p & !v3a6918e;
assign v3757559 = hbusreq6_p & v37674c1 | !hbusreq6_p & v372914b;
assign v3808d2e = hbusreq2 & v3a67c13 | !hbusreq2 & !v8455ab;
assign v3a70772 = hgrant8_p & v8455c9 | !hgrant8_p & v372debd;
assign v3a7138f = jx3_p & v3752d7a | !jx3_p & v373df5c;
assign v3a67312 = hmaster1_p & v8455ab | !hmaster1_p & v376b1ad;
assign v37580b3 = hgrant4_p & v3a6eb39 | !hgrant4_p & v3778fa0;
assign v3a6e2ec = hgrant5_p & v3773f85 | !hgrant5_p & v3a7087c;
assign v37258d6 = hmaster1_p & v372b8a5 | !hmaster1_p & !v3a56847;
assign v3a67698 = hlock3 & v3809b44 | !hlock3 & v37407b3;
assign v3a66e7f = jx0_p & v37702e6 | !jx0_p & v372fe3d;
assign v37453d8 = hlock0_p & v3a70d71 | !hlock0_p & v8455e7;
assign v373e02a = jx2_p & v3a6b368 | !jx2_p & v3765ded;
assign v3a6f8c6 = hgrant7_p & dc57c8 | !hgrant7_p & v3a6897b;
assign v37480ad = hbusreq5 & v375859a | !hbusreq5 & !v3a5fc05;
assign v3a5c27f = hlock3 & v3744f52 | !hlock3 & v37479b4;
assign v37512f6 = hmaster1_p & v376fd84 | !hmaster1_p & v8455ab;
assign v37306c6 = hlock5 & v3754ba1 | !hlock5 & v3a6f4a3;
assign v374fdeb = hmaster1_p & v375db64 | !hmaster1_p & d9e97c;
assign v3a69a00 = hbusreq7_p & v3724f6b | !hbusreq7_p & v377b5dc;
assign v375f52b = hgrant0_p & v37773a9 | !hgrant0_p & v374f1a1;
assign v3a70118 = hbusreq3_p & v375400b | !hbusreq3_p & v8455ab;
assign v37543d8 = hbusreq2_p & v3761c68 | !hbusreq2_p & v3a5a76d;
assign v3a623dc = hbusreq2 & v373e521 | !hbusreq2 & v3a67eec;
assign v3a6f058 = jx0_p & v3a66988 | !jx0_p & v3a2981d;
assign v3a70da3 = hbusreq0 & v3743da0 | !hbusreq0 & v8455ab;
assign v3763f1d = hgrant7_p & v3729139 | !hgrant7_p & c8bdc6;
assign v3a6fc95 = hgrant7_p & v3766ef7 | !hgrant7_p & v3740a9c;
assign v3a70b2d = hmaster1_p & v3a6e7b3 | !hmaster1_p & v377d789;
assign v3a706a2 = hgrant2_p & v8455ab | !hgrant2_p & v372b5af;
assign v374db21 = hbusreq4_p & v372febd | !hbusreq4_p & v3725717;
assign v37365f8 = hlock5 & cbc7dd | !hlock5 & v3809542;
assign v376ad73 = hlock8 & v376ae9f | !hlock8 & v3741b49;
assign v3731bd7 = hmaster1_p & v3a6f7b4 | !hmaster1_p & v3a66811;
assign v3772327 = hmaster2_p & v3767e76 | !hmaster2_p & !v3751510;
assign v3a57b3c = hbusreq4 & v380992b | !hbusreq4 & v8455ab;
assign v3a666a9 = hgrant5_p & v375d98c | !hgrant5_p & v3737b19;
assign v3764702 = hgrant6_p & v377618a | !hgrant6_p & v3806e0e;
assign v376a9ee = hbusreq0 & v372a13a | !hbusreq0 & v3741f08;
assign v374961f = hlock1_p & bad3a6 | !hlock1_p & !v8455ab;
assign v3763ce3 = hbusreq4_p & v8455ab | !hbusreq4_p & v374e314;
assign v37508b9 = hmaster2_p & v3a6f541 | !hmaster2_p & v3a711e8;
assign v3736c86 = hbusreq8_p & v37676a5 | !hbusreq8_p & v37445e6;
assign v3a6ef3f = hbusreq0 & v374648f | !hbusreq0 & v8455ab;
assign v3a6501d = hlock7_p & v3a64e18 | !hlock7_p & v3a55c44;
assign v3a60a9b = hmaster0_p & v377a0da | !hmaster0_p & v3a6fad5;
assign v3a6848c = hgrant4_p & v3767b6e | !hgrant4_p & v3a700ec;
assign v376edbb = hlock5 & v3735ac0 | !hlock5 & v3755691;
assign v3764418 = hbusreq0 & v376480c | !hbusreq0 & v372ce45;
assign v3a6f2d7 = hlock6_p & v3a6c60e | !hlock6_p & v3760f4e;
assign v3724273 = hgrant6_p & v3a71389 | !hgrant6_p & a8fc27;
assign v3a56b60 = hgrant4_p & v3a6f7a1 | !hgrant4_p & v3772541;
assign v3a70b5c = jx1_p & v374b237 | !jx1_p & !v3a597d8;
assign v3a640c5 = hgrant0_p & v8455b3 | !hgrant0_p & v8455ab;
assign v3734067 = hbusreq2_p & v3759b2f | !hbusreq2_p & v3a6f43e;
assign v3a6face = hbusreq4_p & v3a6e0f4 | !hbusreq4_p & v3a70349;
assign v3a66027 = hbusreq2 & v3730fd2 | !hbusreq2 & v8455ab;
assign v3735e18 = jx1_p & v3723df5 | !jx1_p & v3777243;
assign v377ace4 = hbusreq8 & v3767153 | !hbusreq8 & a0a219;
assign v373b58a = stateA1_p & v8455ab | !stateA1_p & v3a70df9;
assign v3771994 = hmaster0_p & v3a7074d | !hmaster0_p & v37329ec;
assign v3a651b5 = hgrant6_p & v3735906 | !hgrant6_p & v3a57cd0;
assign v3767266 = hgrant2_p & v377bfc0 | !hgrant2_p & v3a53bb3;
assign v3a6f0c8 = hmaster2_p & v374729b | !hmaster2_p & v3a5ace5;
assign v374f6a0 = hbusreq6 & v373f058 | !hbusreq6 & v8455ab;
assign v3a5b079 = hbusreq4 & v8455b0 | !hbusreq4 & v373f058;
assign v3a6e91e = hmaster2_p & v8455ab | !hmaster2_p & v377ba55;
assign v3747ed4 = hbusreq0 & v372ab46 | !hbusreq0 & v8455ab;
assign v376e605 = hbusreq5_p & v3a705fc | !hbusreq5_p & v377273d;
assign v374b7b2 = hlock7_p & v3a6dd8f | !hlock7_p & v377e031;
assign v3a656d0 = hbusreq4_p & v3771cf0 | !hbusreq4_p & v376157e;
assign v375db62 = hgrant2_p & v3a709df | !hgrant2_p & v37360b3;
assign v3756a8f = hlock7_p & v375d46e | !hlock7_p & !v374a37e;
assign v3754d8a = hgrant2_p & v3a6f312 | !hgrant2_p & !v3744161;
assign v377ef7c = hlock2_p & v373c97a | !hlock2_p & v375c771;
assign v3772c51 = hbusreq6_p & v3740f3d | !hbusreq6_p & v3a5db8a;
assign v3735fb2 = hbusreq7 & v3724600 | !hbusreq7 & v37782a8;
assign v3a67e64 = hbusreq1_p & v3726d7a | !hbusreq1_p & v8455ab;
assign v37266df = hmaster0_p & v8455ab | !hmaster0_p & v377ecac;
assign v37526ca = hbusreq5_p & v374ffd5 | !hbusreq5_p & v3739b38;
assign v376d856 = locked_p & v3a70cd5 | !locked_p & v39a537f;
assign v3a6deaa = hmaster1_p & v377b848 | !hmaster1_p & v3a6f601;
assign v375f41f = hmaster0_p & v3769093 | !hmaster0_p & v374d138;
assign v3a71452 = hlock1 & v380693e | !hlock1 & v3743b9e;
assign v3a70987 = hbusreq6_p & v9450a2 | !hbusreq6_p & v8455ab;
assign v3a6f03f = hlock2 & v2acaffd | !hlock2 & v3757253;
assign v375e91f = hbusreq6_p & v3775d59 | !hbusreq6_p & v374bfc8;
assign v3a6e3e0 = hbusreq4_p & v3739ea3 | !hbusreq4_p & v377aa06;
assign v372c546 = hbusreq4_p & v377a7e9 | !hbusreq4_p & v8455cb;
assign v3777c6f = hbusreq8_p & v3753ee5 | !hbusreq8_p & v377d607;
assign v3a55cf2 = hlock4_p & v37269f4 | !hlock4_p & v374b3cf;
assign v23fd9e7 = hmaster0_p & v3746a87 | !hmaster0_p & v37289f0;
assign v374edff = hgrant6_p & v3a62b8d | !hgrant6_p & v3743d21;
assign v377dae8 = hbusreq0 & v3a61120 | !hbusreq0 & v3a57d2f;
assign v3a6738f = hready_p & v374140e | !hready_p & v8455e1;
assign v376f319 = hmaster1_p & v8455ab | !hmaster1_p & v3762552;
assign v3767f52 = hlock4_p & v374c5b2 | !hlock4_p & v8455bf;
assign v374726f = hlock8_p & v3a593cc | !hlock8_p & v3a6fba2;
assign v3745a47 = hgrant3_p & v8455ab | !hgrant3_p & v375461f;
assign v325c93a = hgrant7_p & v374b83f | !hgrant7_p & v8ac028;
assign v375f888 = hmaster0_p & v376142a | !hmaster0_p & v3726b90;
assign v3a70233 = hlock0_p & v3a5c945 | !hlock0_p & !v3a619c0;
assign v3768522 = hmaster3_p & v8455ab | !hmaster3_p & v374cf68;
assign v3a70a29 = hburst1 & v3745b85 | !hburst1 & v375b990;
assign v374cb5e = hbusreq7_p & d23562 | !hbusreq7_p & v377f6af;
assign v3741acc = hbusreq6_p & v3a66014 | !hbusreq6_p & v3763011;
assign v3a630dc = hlock4 & v373bb2c | !hlock4 & v3766117;
assign v3a60a32 = hbusreq0 & v37311a4 | !hbusreq0 & !v3a61279;
assign v373bf7c = stateA1_p & v8455ab | !stateA1_p & !v373a7d4;
assign v3a6602e = hmaster0_p & v3a660c0 | !hmaster0_p & v3a57e58;
assign v3758079 = hburst0 & v8455ab | !hburst0 & !v3a563ad;
assign v373bb2d = hgrant3_p & v375c7b9 | !hgrant3_p & !v37477d2;
assign v3a6fcf9 = hbusreq3 & v373d9aa | !hbusreq3 & v374f609;
assign v2ff937f = hgrant4_p & v3769ed3 | !hgrant4_p & v37265b8;
assign v3a6ae12 = hbusreq7 & v3255b27 | !hbusreq7 & v3a61519;
assign v3a67de3 = hbusreq0 & v3a56eb1 | !hbusreq0 & v8455ab;
assign v37604d6 = hbusreq5_p & v3a715e5 | !hbusreq5_p & !v8455ab;
assign v3a6ff55 = hbusreq7_p & v3a6ffd8 | !hbusreq7_p & v3777d70;
assign v3a712c5 = hbusreq4 & v3769cd3 | !hbusreq4 & v8455ab;
assign v377b2ce = hgrant2_p & v3748792 | !hgrant2_p & v3a6bbed;
assign v372914b = hbusreq2_p & v37674c1 | !hbusreq2_p & v3761ad0;
assign v3766f7d = hlock2_p & v37266b1 | !hlock2_p & v8455e7;
assign v3777d63 = hlock5_p & v37263c1 | !hlock5_p & v3a656ca;
assign v3761915 = hbusreq5_p & v3a708a0 | !hbusreq5_p & v374c9ab;
assign v3a70c91 = hmaster2_p & v3a54c9b | !hmaster2_p & v3771715;
assign v3732d55 = hbusreq2_p & v3a6ac7e | !hbusreq2_p & !v8455ab;
assign v37563bc = hbusreq7_p & v3733cf4 | !hbusreq7_p & v3a592bc;
assign v3a62dec = hgrant7_p & v8455ce | !hgrant7_p & v3766809;
assign v3723ded = hgrant2_p & v8455ba | !hgrant2_p & v372c06f;
assign v3a70e87 = hmaster1_p & v3753921 | !hmaster1_p & v374e855;
assign v3a70c66 = stateG10_1_p & v372dab1 | !stateG10_1_p & v372e5d3;
assign v3743c7e = hmaster2_p & v8455ab | !hmaster2_p & v37258b7;
assign v3a6dea7 = jx1_p & v380a20c | !jx1_p & v3a713d7;
assign v3a71400 = hbusreq3_p & v373a374 | !hbusreq3_p & v37584fe;
assign v3761cec = hbusreq1_p & v3a6b4fb | !hbusreq1_p & v3732b98;
assign v3a6fea8 = hbusreq2 & v372b373 | !hbusreq2 & v3a6f6e7;
assign v3a60755 = hbusreq5 & v374c6ff | !hbusreq5 & v3a61323;
assign v3a71635 = hmaster2_p & v8455ab | !hmaster2_p & !v3778ed4;
assign v375f368 = hmaster0_p & v377a2f2 | !hmaster0_p & v3755914;
assign v3a6f6a4 = hbusreq4_p & v3a5d494 | !hbusreq4_p & v8455ab;
assign v3751406 = hlock8 & v37509c4 | !hlock8 & v372c1bb;
assign v987445 = hlock5_p & v3742b92 | !hlock5_p & v3722b6c;
assign v37364a3 = hmaster1_p & v3a64eba | !hmaster1_p & v3776bc7;
assign v377946d = hmaster1_p & v3733d3f | !hmaster1_p & v3729381;
assign v3767897 = hmaster2_p & v3a61081 | !hmaster2_p & !v374a2cc;
assign v23fe156 = hbusreq5_p & v8455b7 | !hbusreq5_p & v372433d;
assign v3a6dfa3 = hmaster0_p & v3746e8b | !hmaster0_p & v3a63033;
assign a7b390 = hmaster0_p & v3725198 | !hmaster0_p & v37659e4;
assign v3a2a8f2 = hbusreq6_p & v3a636d9 | !hbusreq6_p & v3a533d3;
assign v3a6e130 = hmaster2_p & v3772f85 | !hmaster2_p & v3808eed;
assign v3a58519 = hmaster2_p & v8455ab | !hmaster2_p & !v3a66af8;
assign v3748755 = hbusreq2 & v37251b9 | !hbusreq2 & v376f768;
assign v3a6ef22 = hgrant6_p & v3a60a68 | !hgrant6_p & a72315;
assign v373c5f5 = hbusreq2 & v3a6dc08 | !hbusreq2 & v3730ffe;
assign v3a706bd = hbusreq5 & v376f56d | !hbusreq5 & !v3768e52;
assign v3a5c4e8 = hgrant4_p & v8455ab | !hgrant4_p & v3a56da3;
assign v3766b05 = hmaster2_p & v8455ab | !hmaster2_p & v3760e75;
assign v3728d57 = hlock5 & v3a61302 | !hlock5 & v3a62819;
assign v3a70b46 = hmaster1_p & v3a5e24e | !hmaster1_p & v3a5dd60;
assign v376f6e4 = hmaster2_p & v3a6f92f | !hmaster2_p & v3768c3c;
assign v360d177 = hmaster1_p & v3a70efe | !hmaster1_p & !v8455b3;
assign v372f1a8 = hgrant5_p & v3766afa | !hgrant5_p & v3a5b01a;
assign v3a6eeff = hgrant2_p & v8455ba | !hgrant2_p & v3724002;
assign v37434e1 = hmaster2_p & v8455ab | !hmaster2_p & v3742f64;
assign v374c28e = hgrant5_p & v37250b1 | !hgrant5_p & v3743156;
assign v375b01a = hbusreq6_p & v372ce88 | !hbusreq6_p & v375deaa;
assign v3a700c8 = hmaster0_p & v375c044 | !hmaster0_p & v374e39c;
assign v374fda1 = hmaster2_p & v375fbf2 | !hmaster2_p & !v375d9b1;
assign v37565be = hbusreq6 & v3768130 | !hbusreq6 & v377728d;
assign v3736958 = hbusreq8 & v3a70081 | !hbusreq8 & v375aa9b;
assign c03a6a = hmaster0_p & v3a6d768 | !hmaster0_p & !v377e004;
assign v37514dd = hlock8 & v3a6fc58 | !hlock8 & v3734e23;
assign v3751389 = hbusreq4_p & v3a69584 | !hbusreq4_p & v3a6ffae;
assign v3a7163f = hbusreq0 & v3a6620b | !hbusreq0 & v373bd6c;
assign v3a7016e = hlock7 & v3a5ed98 | !hlock7 & v3a299f3;
assign v3a6ff33 = hmaster0_p & v3a7052e | !hmaster0_p & v376ff64;
assign v37686f6 = hgrant2_p & v8455ab | !hgrant2_p & v3a702fe;
assign v3767c92 = hbusreq8 & v3724600 | !hbusreq8 & v8455ab;
assign v37301f9 = hbusreq8_p & v374bdfb | !hbusreq8_p & v3756cea;
assign v3738aef = jx0_p & v375fbe1 | !jx0_p & v8455ab;
assign v373098e = hmaster0_p & v3753eb2 | !hmaster0_p & v380911e;
assign v3741566 = hmaster1_p & v37330d3 | !hmaster1_p & v3a70503;
assign v37308bf = hmaster2_p & v8455ab | !hmaster2_p & v3806f67;
assign v3a6f0f7 = hmaster3_p & v37600ad | !hmaster3_p & v3769c19;
assign v3750fea = stateG2_p & v8455ab | !stateG2_p & !v377f108;
assign v374b330 = hmaster1_p & v8455ab | !hmaster1_p & v377bd81;
assign v3a6eb6b = hgrant3_p & v8455ab | !hgrant3_p & !v3752ec0;
assign v3730587 = hmaster1_p & v3a66d47 | !hmaster1_p & v376046c;
assign v37510ae = hgrant3_p & v373e12e | !hgrant3_p & !v374fa0a;
assign a80fe2 = hmaster1_p & v3a635ea | !hmaster1_p & v3a6eaf8;
assign v3a62a9d = stateA1_p & v8455e1 | !stateA1_p & !v373513a;
assign v3755508 = hbusreq5_p & v3a5e859 | !hbusreq5_p & v3a71658;
assign v375967d = hlock8 & v373c126 | !hlock8 & v37597fa;
assign v3a538b3 = hbusreq5 & v3a62d5d | !hbusreq5 & v3a635ea;
assign v375e2ab = hlock2_p & v3763c04 | !hlock2_p & !v373abe2;
assign v373714f = hbusreq8_p & v37742c5 | !hbusreq8_p & v8455ab;
assign v37280b0 = hbusreq2_p & v377caa3 | !hbusreq2_p & v377efdc;
assign v3a70ce8 = hmaster1_p & v374caf9 | !hmaster1_p & v3a71656;
assign v372cd04 = hmaster2_p & v3754df4 | !hmaster2_p & v373ae83;
assign v3a6ff41 = busreq_p & v377fbb9 | !busreq_p & !v373b58a;
assign v3a53329 = hbusreq4 & v3750c9f | !hbusreq4 & v8455ab;
assign v3a6a8aa = hmaster1_p & v3777f05 | !hmaster1_p & v3745871;
assign v3a6ff6f = hbusreq5 & v372a22f | !hbusreq5 & v8455ab;
assign v3779177 = hmaster1_p & v3a6dc83 | !hmaster1_p & v374db73;
assign v37749b7 = hbusreq1 & v39a5265 | !hbusreq1 & !v2aca977;
assign v3747192 = hmaster0_p & v8455ab | !hmaster0_p & v3746211;
assign v3729bd7 = hbusreq1 & v3a6ac26 | !hbusreq1 & v2aca977;
assign v3725092 = hbusreq2 & v373aaa8 | !hbusreq2 & v8455ab;
assign v3a7100a = hbusreq8 & v375f985 | !hbusreq8 & a0a219;
assign v3a59ee0 = hbusreq6 & v3a7163c | !hbusreq6 & v8455ab;
assign v3a70696 = hmaster2_p & v3a710c6 | !hmaster2_p & v3732415;
assign v3a5ec68 = hbusreq5 & v94faa4 | !hbusreq5 & v8455ab;
assign v3744724 = hlock6_p & v375444e | !hlock6_p & v8455b0;
assign v37270b9 = hmaster2_p & v3752aa5 | !hmaster2_p & v8455ab;
assign v3764fad = hmaster1_p & v377316f | !hmaster1_p & v3751b9a;
assign v3724547 = hbusreq5 & v3769325 | !hbusreq5 & v3a63f9a;
assign v2092ac1 = hmaster1_p & v3765bf4 | !hmaster1_p & v3a6eed9;
assign v3775e7e = hmaster0_p & v374e079 | !hmaster0_p & v3777ee7;
assign v3a70dd6 = hgrant3_p & v37362fc | !hgrant3_p & v3740ee1;
assign v3740cb5 = hmaster1_p & v3a70557 | !hmaster1_p & v3a6d5e2;
assign v37293b1 = hbusreq3_p & v3a70c38 | !hbusreq3_p & v35772a6;
assign v3a6504e = hgrant6_p & v37332c8 | !hgrant6_p & v37487a4;
assign v37467a6 = hbusreq2 & v373fe5e | !hbusreq2 & !v376430b;
assign v374f7b7 = hbusreq6_p & v3a6f9df | !hbusreq6_p & !v377cd5b;
assign v940c77 = hmaster0_p & v375d6b4 | !hmaster0_p & v375c76b;
assign v3759470 = hbusreq3_p & v3a6f7f0 | !hbusreq3_p & v373d7fe;
assign v3771b8a = hbusreq5_p & v3776b93 | !hbusreq5_p & !v375818a;
assign v3a6e8db = hbusreq7 & v3776066 | !hbusreq7 & v37305e6;
assign v375e815 = hbusreq4 & v37413d8 | !hbusreq4 & v3763209;
assign v372fa3a = hmaster2_p & v377d1dc | !hmaster2_p & v373b02e;
assign v3256555 = hmaster1_p & v3a7066c | !hmaster1_p & v3a54dd4;
assign v375ac23 = hbusreq3_p & v3a63805 | !hbusreq3_p & v8455b0;
assign v380992b = hlock4_p & v37366d0 | !hlock4_p & v3a715d2;
assign v377bb21 = hgrant2_p & v3733d6e | !hgrant2_p & v3a6eee6;
assign v377395f = locked_p & v3773ca9 | !locked_p & !v8455ab;
assign v3a673d9 = hmaster1_p & v3a55672 | !hmaster1_p & v8455ab;
assign v3a63ee6 = hmaster2_p & v35b7808 | !hmaster2_p & v373bf45;
assign v376e966 = hmaster3_p & v3a7017a | !hmaster3_p & v3762aaf;
assign v374fd4a = hgrant3_p & v3771d77 | !hgrant3_p & v3756398;
assign v3775c24 = hlock5_p & v376fd84 | !hlock5_p & v8455ab;
assign v3767153 = hlock7 & a0a219 | !hlock7 & v3a6165b;
assign v375095a = hmaster2_p & v374362e | !hmaster2_p & v3767f33;
assign v3773c69 = hbusreq3_p & v37250a3 | !hbusreq3_p & v3a69946;
assign ac6831 = hbusreq7_p & v376d892 | !hbusreq7_p & v380702c;
assign v39a52e6 = hgrant6_p & v3a6fbe4 | !hgrant6_p & v3a7145f;
assign v374109e = hgrant4_p & v37346be | !hgrant4_p & v3777573;
assign v3a5c94c = hbusreq4_p & v8455b3 | !hbusreq4_p & v3767437;
assign v377a7e9 = hbusreq4 & v3a6fc48 | !hbusreq4 & v375a38b;
assign v373abdd = hgrant4_p & v372e7f8 | !hgrant4_p & v8455ab;
assign v3a6f61e = hbusreq6_p & v372a2f5 | !hbusreq6_p & !v3a6fb1f;
assign v37396f7 = hmaster2_p & v37782c9 | !hmaster2_p & v375c675;
assign v3751913 = hgrant4_p & v3744637 | !hgrant4_p & v3a7112a;
assign v376f182 = hmaster0_p & v373a4e4 | !hmaster0_p & v377da14;
assign v3a70618 = hbusreq8 & v372b386 | !hbusreq8 & v37727f9;
assign v3a6fa4c = hbusreq4_p & v37625ef | !hbusreq4_p & v373b288;
assign v3a702f6 = hlock5 & v3756ead | !hlock5 & v37606f4;
assign v3a69758 = hmaster0_p & v8455ab | !hmaster0_p & v3a6bc0e;
assign v3a6fb88 = hmaster0_p & v3807aa1 | !hmaster0_p & v3a6ef26;
assign v374908e = hmaster2_p & v374502e | !hmaster2_p & !v376b4e1;
assign v3a61992 = hbusreq7 & v3765121 | !hbusreq7 & v3a67f49;
assign v87be38 = hbusreq5_p & v3a5b289 | !hbusreq5_p & v3a701a1;
assign v1e379e9 = hgrant2_p & v8455ab | !hgrant2_p & v3741797;
assign v3740766 = hlock7_p & v37586cd | !hlock7_p & v37799a0;
assign v3758bfe = hmaster0_p & v3737bb4 | !hmaster0_p & v3761bee;
assign v375f3cf = hgrant5_p & v8455ab | !hgrant5_p & v3a6f8c0;
assign v3a707e3 = hmaster1_p & v3809561 | !hmaster1_p & v3724df8;
assign v3a6f744 = hlock0_p & v3740f3d | !hlock0_p & v8455ab;
assign v1e37bdd = hbusreq0_p & v3730f98 | !hbusreq0_p & v8455ab;
assign v3762886 = hbusreq6 & bbab81 | !hbusreq6 & v8455ab;
assign v3a6fafb = hbusreq5_p & v3a70a00 | !hbusreq5_p & v372ee20;
assign v37317a9 = hbusreq1_p & v3a635ea | !hbusreq1_p & !a4a7a5;
assign v3724e8e = hbusreq3_p & v37471cb | !hbusreq3_p & v8455ab;
assign v375c423 = hbusreq4 & v3a6fcb9 | !hbusreq4 & v8455ab;
assign v3a70159 = hbusreq3 & v23fd7d9 | !hbusreq3 & v3743e56;
assign v3a5eb73 = hgrant0_p & v8455ab | !hgrant0_p & v3746368;
assign v3a6eb94 = hgrant2_p & v377d4a0 | !hgrant2_p & v3a6ebdb;
assign v3770a6d = hbusreq5 & v3733e30 | !hbusreq5 & v8455c2;
assign v3a608c4 = hmaster1_p & v3a6f724 | !hmaster1_p & v3a5463b;
assign v376438f = hmaster2_p & v3a70f53 | !hmaster2_p & v3a53e66;
assign d27546 = hgrant3_p & v3a637dc | !hgrant3_p & v3a70208;
assign v3a702be = hmaster0_p & v376db9c | !hmaster0_p & v88d9b8;
assign v3a6cf46 = hmaster2_p & v8455ab | !hmaster2_p & v3a6911d;
assign v3a70ed6 = hbusreq6 & v3a5f8d0 | !hbusreq6 & v8455ab;
assign v374a9e7 = hgrant3_p & v376e914 | !hgrant3_p & v3769157;
assign v3a5d494 = hbusreq4 & v3a5600a | !hbusreq4 & v8455ab;
assign v372d3b2 = hbusreq5_p & v37267f3 | !hbusreq5_p & v374a41b;
assign v3756ef1 = hgrant4_p & v37300a5 | !hgrant4_p & v3723701;
assign v375d76b = hmaster2_p & v3a5d94a | !hmaster2_p & v8455c2;
assign v3754afa = hmaster1_p & v20d166d | !hmaster1_p & v3741d83;
assign v372e5a8 = hgrant5_p & v376530c | !hgrant5_p & v3a5c653;
assign v3a60d86 = hgrant6_p & v374ca88 | !hgrant6_p & v375b34f;
assign v37388a7 = hbusreq4_p & v3a71188 | !hbusreq4_p & v3a712d3;
assign v373a18b = hlock0 & v3a7162d | !hlock0 & v8827d7;
assign v3a5f0d0 = hbusreq5_p & v377eb8b | !hbusreq5_p & v3808d85;
assign v37306d8 = hbusreq2 & v375f8b0 | !hbusreq2 & v375fbc0;
assign v3a6324e = hgrant5_p & v3739940 | !hgrant5_p & a27bd0;
assign v372cd91 = hbusreq0 & v376311f | !hbusreq0 & v3760d74;
assign v3724d8b = hlock7 & v3a607ba | !hlock7 & v3741e9f;
assign v3a6c610 = hmaster0_p & v3770bc0 | !hmaster0_p & v3757966;
assign v3779cd7 = hbusreq4_p & v373f058 | !hbusreq4_p & v3753dab;
assign v375cd5d = hbusreq4_p & v373d7f9 | !hbusreq4_p & v377b0f7;
assign v375fbd7 = hbusreq1_p & v372dec8 | !hbusreq1_p & v3a71345;
assign v3a5881c = hmaster3_p & v8455ab | !hmaster3_p & v372ee18;
assign v37691e6 = hmaster2_p & v3763fdc | !hmaster2_p & v3769374;
assign v3738321 = hmaster2_p & v8455ab | !hmaster2_p & !v3729430;
assign v376e238 = hgrant3_p & v377dd3b | !hgrant3_p & v375ad91;
assign v3753e74 = hbusreq7 & v37593c6 | !hbusreq7 & v8455ab;
assign v3a6fda4 = hbusreq2 & v377ac7e | !hbusreq2 & v37749bf;
assign v3a7134d = hbusreq2_p & v3a635ea | !hbusreq2_p & v376bade;
assign v3a54952 = hgrant5_p & v37335e0 | !hgrant5_p & v37239a5;
assign v3a62dfa = hmaster2_p & v373feaa | !hmaster2_p & v3a6f4eb;
assign v375896e = hbusreq4 & v37379bb | !hbusreq4 & !v3a703de;
assign v3758fa7 = hbusreq2_p & v3a61a3d | !hbusreq2_p & !v8455ab;
assign v3a6f025 = hmaster2_p & v3a635ea | !hmaster2_p & v3759f09;
assign v3a66af8 = hbusreq4_p & v3755cb2 | !hbusreq4_p & v3a6ffe1;
assign v3a53f38 = hmaster0_p & v3a5e24e | !hmaster0_p & v3a6aada;
assign v3a603c1 = hlock5_p & v3a6581d | !hlock5_p & !v3a6f3b8;
assign v374c671 = hbusreq2 & v374ad1e | !hbusreq2 & v8455b0;
assign v374bdfb = hgrant5_p & v3a6f8e7 | !hgrant5_p & v3a5bcc4;
assign v374291b = hgrant6_p & v372952e | !hgrant6_p & v3a6d299;
assign v3a6cc93 = hmaster0_p & v374df63 | !hmaster0_p & v372f997;
assign v2acae4c = hlock4 & v3761466 | !hlock4 & v37255a7;
assign v3a70c5d = hbusreq0 & v3a65503 | !hbusreq0 & v37532ac;
assign v3778ef8 = hbusreq1 & v37482f8 | !hbusreq1 & !v3a6fe6a;
assign v3a5c484 = hbusreq8_p & v376ae9f | !hbusreq8_p & v3773bf5;
assign v3a6f031 = hlock8_p & v3a7131f | !hlock8_p & v3a7007c;
assign v3a70460 = hbusreq4_p & v3a635ea | !hbusreq4_p & v1e37c0d;
assign v3a6f4c9 = hbusreq5 & v3a5a81d | !hbusreq5 & v8455ab;
assign v3a6f81f = hbusreq1 & v374f87c | !hbusreq1 & v8455ab;
assign v377df9c = hgrant4_p & v3a7025d | !hgrant4_p & v3a6f3fb;
assign v375607f = hgrant4_p & v3a6fac2 | !hgrant4_p & v3746ab1;
assign v376e370 = hmaster2_p & v3a62a6d | !hmaster2_p & v374513e;
assign v37533e3 = hlock3_p & v35772b3 | !hlock3_p & v35772a6;
assign v3a70bc6 = hbusreq4 & v3723b00 | !hbusreq4 & v8455ab;
assign v3a6f487 = hmaster1_p & v372d8e8 | !hmaster1_p & v375a5f9;
assign v376e3a3 = hgrant5_p & v3a679b5 | !hgrant5_p & v3a706b8;
assign v3759590 = hgrant0_p & v3a6b873 | !hgrant0_p & !v372a9bd;
assign v37798ad = hbusreq2_p & v375bdd4 | !hbusreq2_p & v3a6f549;
assign v3a63f30 = hlock2_p & v372391f | !hlock2_p & v375e60f;
assign v3a5b6c5 = hgrant2_p & v8455ab | !hgrant2_p & !v3742d37;
assign v3763502 = hbusreq7_p & v3a6167d | !hbusreq7_p & v37649a5;
assign v376e77e = hbusreq5_p & v374d9c0 | !hbusreq5_p & v3767ee9;
assign v372a1b6 = hmaster2_p & v38087c5 | !hmaster2_p & v3772f85;
assign v37668b8 = hmaster1_p & v8455ab | !hmaster1_p & v3a59ce1;
assign v374d542 = hbusreq2_p & v3a5a01a | !hbusreq2_p & v3731be6;
assign v3a6f6af = hmaster1_p & v375c62d | !hmaster1_p & v3779678;
assign v372b1c8 = hgrant6_p & v37432c6 | !hgrant6_p & v374b36e;
assign v37387e6 = hgrant5_p & v8455ab | !hgrant5_p & !v97e702;
assign v3a54ba7 = hbusreq0 & v374262b | !hbusreq0 & v3750d44;
assign v373c377 = hbusreq6 & v910050 | !hbusreq6 & v3a7011e;
assign v3a6fb8c = hgrant6_p & v3a57fff | !hgrant6_p & v3747ec5;
assign v373a3e7 = hlock5_p & v3a70b19 | !hlock5_p & !v8455ab;
assign v3a624d7 = hbusreq5 & v3764334 | !hbusreq5 & v8455ab;
assign v3a71109 = hgrant1_p & v3762de1 | !hgrant1_p & !v37457fb;
assign v3a61603 = hbusreq4_p & v373d136 | !hbusreq4_p & v373f4ce;
assign v3a70042 = hlock8_p & v372c298 | !hlock8_p & v375b22c;
assign v3a702fc = hbusreq5_p & v3727b10 | !hbusreq5_p & v3728f6d;
assign v373b50e = hbusreq4 & v3768349 | !hbusreq4 & v3753bb2;
assign v3a6d81d = hgrant6_p & v374352b | !hgrant6_p & v3a5e1bc;
assign v375416d = hgrant3_p & v374306c | !hgrant3_p & v37614c8;
assign v3a6f769 = hlock7_p & v3739b18 | !hlock7_p & cae8ef;
assign v3a705e4 = hmaster0_p & v374ac8c | !hmaster0_p & v3a715c3;
assign v3778ed4 = locked_p & v8455e1 | !locked_p & !v8455ab;
assign v3a70821 = hlock0 & v375c70c | !hlock0 & v3a57ec9;
assign v374dabe = hmaster0_p & v8455ab | !hmaster0_p & v377d21c;
assign v372a2f5 = hbusreq6 & v3a70fb2 | !hbusreq6 & v3a705c5;
assign v376fd33 = hmaster0_p & v375c1c5 | !hmaster0_p & !v3747dd8;
assign v3a6f84c = hmaster2_p & v3a57584 | !hmaster2_p & !v3a707c4;
assign v377d2bb = hbusreq5 & v373c8ba | !hbusreq5 & v3a700af;
assign v3a569b7 = hbusreq0 & v39eb4ca | !hbusreq0 & v3a6499e;
assign v1e377ba = hgrant4_p & v3723299 | !hgrant4_p & v3a6f8a0;
assign v375d4aa = hmaster2_p & v3768bbc | !hmaster2_p & v3a6f0bc;
assign v3732202 = hbusreq6_p & v3a594a5 | !hbusreq6_p & v3750134;
assign v3a6efc3 = hmaster3_p & v37493ed | !hmaster3_p & v3a66988;
assign v377a8dc = hbusreq5 & v377109a | !hbusreq5 & !v8455bd;
assign v37383b1 = hbusreq7 & v3a65dce | !hbusreq7 & v8455ab;
assign v3767527 = hlock0_p & v3771728 | !hlock0_p & v3773069;
assign b736f4 = hbusreq5_p & v3731f6b | !hbusreq5_p & v3724696;
assign v3a57ed1 = hbusreq6 & v372b304 | !hbusreq6 & v8455ab;
assign v3a595fe = hmaster2_p & v3a62542 | !hmaster2_p & v37745a0;
assign v375928d = hbusreq3 & v3733383 | !hbusreq3 & v8455ab;
assign v37411bc = hbusreq4 & v3762385 | !hbusreq4 & v3a6f71a;
assign v37747c0 = hgrant4_p & v373ef69 | !hgrant4_p & v3a6de03;
assign v3764486 = hbusreq6_p & v375a0b3 | !hbusreq6_p & v37715af;
assign v3a6f89b = hbusreq5_p & v37655ff | !hbusreq5_p & !v8455ab;
assign v3730df7 = hmaster1_p & v3a712d8 | !hmaster1_p & v3729ed5;
assign v37386af = hbusreq7 & v3a6fa2a | !hbusreq7 & v3a62aa3;
assign v372a7e7 = hmaster3_p & v3736948 | !hmaster3_p & v3a6f850;
assign v3a6c631 = hmaster2_p & v3a712e2 | !hmaster2_p & v3736026;
assign v3762c73 = hbusreq6 & b4f73f | !hbusreq6 & v3767429;
assign v3a6f222 = hmaster0_p & v3a60d5e | !hmaster0_p & v376dd15;
assign v3a6ecf6 = hlock4_p & v35b7769 | !hlock4_p & v372d10e;
assign v3747400 = hgrant4_p & v3807a80 | !hgrant4_p & v373abbb;
assign v376fd84 = hmaster0_p & v376c224 | !hmaster0_p & v8455ab;
assign v3a6fd4b = hbusreq4 & v374ad67 | !hbusreq4 & v376c76d;
assign v373ee52 = hbusreq0 & v375a7d3 | !hbusreq0 & v376aa99;
assign v375685b = hbusreq6 & v3763191 | !hbusreq6 & v35b774b;
assign v374c234 = stateA1_p & v8455ab | !stateA1_p & v3a6f8a1;
assign v374b1bc = hbusreq4_p & v8455e7 | !hbusreq4_p & v374f307;
assign v3a714d2 = hbusreq6 & v3723495 | !hbusreq6 & v375b2fe;
assign v373afc3 = hgrant4_p & a8c5c5 | !hgrant4_p & v325c960;
assign v376a799 = hbusreq5 & v3761bd1 | !hbusreq5 & v375f906;
assign v3756149 = hbusreq2 & v3746c51 | !hbusreq2 & v8455ab;
assign v3733471 = hlock0_p & v3a63805 | !hlock0_p & v3745075;
assign v3a6f7ed = hbusreq4 & v374829e | !hbusreq4 & v3775999;
assign v376f584 = hbusreq6 & v3a70a50 | !hbusreq6 & v3a70b92;
assign v3761e97 = hbusreq5_p & v3777647 | !hbusreq5_p & v375ed5c;
assign v372c4bd = hgrant0_p & v374d140 | !hgrant0_p & v380853c;
assign v3748fe0 = hmaster2_p & v377d7dc | !hmaster2_p & v3729f25;
assign v325b5df = hlock4 & v3a70511 | !hlock4 & v3a5c462;
assign v3752a05 = hgrant8_p & v8455ab | !hgrant8_p & !v3739e0d;
assign v373b42b = hbusreq2 & v377dcbc | !hbusreq2 & v372c151;
assign v37361aa = hgrant0_p & v8455e7 | !hgrant0_p & ad2d05;
assign v37687ce = stateA1_p & v375956a | !stateA1_p & v3a6feed;
assign v3738df9 = hgrant2_p & v3a6f20d | !hgrant2_p & baf7ba;
assign v38063ce = hmaster0_p & v37229db | !hmaster0_p & v372f9cf;
assign v3772698 = hbusreq3_p & v3769ae2 | !hbusreq3_p & v37574f8;
assign v3742c62 = hmaster0_p & v98083e | !hmaster0_p & v377d1dc;
assign v375deaa = hbusreq6 & v374b3cf | !hbusreq6 & v8455b3;
assign v3725a21 = hmaster0_p & v372f326 | !hmaster0_p & v3767121;
assign v3a6830a = hbusreq4 & v1e38224 | !hbusreq4 & v8455ab;
assign v3a5e2a3 = hgrant4_p & v8455b0 | !hgrant4_p & v38090f4;
assign v3a70509 = hbusreq4 & v3759c49 | !hbusreq4 & v2092abe;
assign v3a6dcdc = hbusreq2_p & v8455b7 | !hbusreq2_p & v3753d60;
assign v3a660b5 = hlock4_p & v37581c2 | !hlock4_p & v3722a7e;
assign v377bae8 = hmaster0_p & v3a70235 | !hmaster0_p & v375f6c7;
assign v3a5d176 = jx0_p & v372ff37 | !jx0_p & v3752cc4;
assign v3a710ff = hlock7 & v3a707e1 | !hlock7 & v3724cce;
assign v373f2d1 = hgrant6_p & v3a6ab8c | !hgrant6_p & v377839d;
assign v3a7079f = hmaster0_p & v375058e | !hmaster0_p & v376a6f1;
assign v376bebb = hlock4 & v3728034 | !hlock4 & v373f9db;
assign v3779fdf = hbusreq8_p & v375d351 | !hbusreq8_p & v374a9fa;
assign v3748ca3 = hready & v375eb9c | !hready & v3a70b47;
assign v3a70f18 = hlock4 & v3a70753 | !hlock4 & v3a6582b;
assign v3739c9a = hgrant8_p & v3768e1e | !hgrant8_p & dc3a01;
assign v3a6ae99 = hbusreq1_p & v376e00a | !hbusreq1_p & !v375d651;
assign v3a6ef86 = hgrant2_p & v373744b | !hgrant2_p & v3722bcf;
assign v3a62fd2 = hmaster1_p & v3a6f382 | !hmaster1_p & !v3a5733c;
assign v3a713dc = hgrant3_p & v3764276 | !hgrant3_p & v376e9e2;
assign v376625e = hgrant5_p & v3765e47 | !hgrant5_p & v3724c46;
assign v3737084 = hgrant2_p & v3758472 | !hgrant2_p & !v376064b;
assign v37680a7 = hmaster0_p & v377576e | !hmaster0_p & v8455ab;
assign v3a5b6b0 = hmaster0_p & v376a11d | !hmaster0_p & v3a70fae;
assign v374794f = hlock0_p & v372dadb | !hlock0_p & v3a6fe5b;
assign v3730b67 = hmaster1_p & v373e625 | !hmaster1_p & v377eada;
assign v37592c9 = hbusreq8_p & v3a5b660 | !hbusreq8_p & v375982a;
assign v3767e66 = hmaster2_p & v375d337 | !hmaster2_p & !v2ff8cfd;
assign v3a6fc9b = hbusreq6_p & v3758a0c | !hbusreq6_p & v37571da;
assign v2925ca9 = hbusreq0 & v3753e49 | !hbusreq0 & v374eda5;
assign v3a62197 = hbusreq4 & v375b349 | !hbusreq4 & v3a635ea;
assign v3a6fd77 = hmaster1_p & v3a710c5 | !hmaster1_p & v373647a;
assign v373d2bd = hbusreq4_p & v3751510 | !hbusreq4_p & v3764eb2;
assign v377206b = hbusreq0 & v376bebb | !hbusreq0 & v3a7080b;
assign v3a5ad1d = hgrant6_p & v3a5cd51 | !hgrant6_p & v373e10f;
assign v37784b9 = hgrant4_p & v3a7133d | !hgrant4_p & v3767650;
assign v3a666e8 = hlock6_p & v37757e0 | !hlock6_p & v8455b0;
assign v375e093 = hbusreq8 & v39ebaee | !hbusreq8 & v3a6f1d8;
assign v374d28d = hgrant6_p & v8455ab | !hgrant6_p & v3a5b841;
assign v37467f3 = hlock1_p & v3774911 | !hlock1_p & v3a6f10f;
assign v3725901 = hmaster2_p & v3767b70 | !hmaster2_p & v3a67905;
assign v3a637e0 = hlock2 & v373cf3a | !hlock2 & v325c976;
assign v3a701ce = hmaster0_p & v3a5b8b9 | !hmaster0_p & v3a6f818;
assign v3a6ff08 = hbusreq0 & v37281e7 | !hbusreq0 & v3a714be;
assign v374caab = hbusreq3_p & v8455ab | !hbusreq3_p & v37665bf;
assign v376f45e = stateG10_1_p & v3a57330 | !stateG10_1_p & v3a6cf18;
assign v374f033 = stateG10_1_p & v3750746 | !stateG10_1_p & v3730de9;
assign v37631d9 = hgrant4_p & v8455ab | !hgrant4_p & v375026b;
assign v377c977 = hbusreq5_p & v3751887 | !hbusreq5_p & v3a70ed3;
assign v3a6fdcb = hmaster0_p & v3753825 | !hmaster0_p & v3a6230b;
assign v3a702ef = hmaster1_p & v3737c04 | !hmaster1_p & v3a63812;
assign v3a6f4cc = hgrant5_p & v8455ab | !hgrant5_p & d3482c;
assign v3a6f657 = hmaster3_p & v8455ab | !hmaster3_p & b1f79b;
assign v372ff2c = hbusreq2 & v3a6fcb9 | !hbusreq2 & v8455ab;
assign v3772c95 = hmaster0_p & v3747e1f | !hmaster0_p & v8455e7;
assign v3a656a4 = hmaster0_p & v374c8a8 | !hmaster0_p & v3a6d407;
assign v3a6eb77 = hgrant1_p & v3a66110 | !hgrant1_p & v3a70ecf;
assign v3a6f4d3 = hbusreq1 & v373a27c | !hbusreq1 & v8455e7;
assign v37428b3 = hmaster2_p & v376e89b | !hmaster2_p & v3752e63;
assign v3a70033 = hmaster0_p & v377e692 | !hmaster0_p & v3a70caa;
assign v37341d3 = hmaster2_p & v2acb095 | !hmaster2_p & b038e6;
assign v3779680 = hbusreq4_p & v3a6fbf8 | !hbusreq4_p & !v8455ab;
assign v37293f2 = hmaster2_p & v376d9ad | !hmaster2_p & v3740171;
assign v373d98d = hbusreq5_p & v37525c8 | !hbusreq5_p & v3754717;
assign v8f695f = hbusreq3_p & v3a705d7 | !hbusreq3_p & v8455ab;
assign v3757b58 = hbusreq4_p & v3a5dde7 | !hbusreq4_p & v3a70a3b;
assign v375eef0 = hlock5_p & v3a67a48 | !hlock5_p & v9a3ffa;
assign v3a63dbf = hlock6 & v3748797 | !hlock6 & v3768d29;
assign v372bcbc = hbusreq0_p & v374ab5b | !hbusreq0_p & v8455ab;
assign v377d0fc = hgrant4_p & v8455ab | !hgrant4_p & v375a677;
assign v3a5810a = hbusreq3 & v3759b9a | !hbusreq3 & v8455ab;
assign v3a70e9e = hbusreq0 & v376f56d | !hbusreq0 & v8455b6;
assign v37400d8 = hbusreq5_p & v372d060 | !hbusreq5_p & v37613bf;
assign v377e630 = hmaster2_p & v376e717 | !hmaster2_p & v8455ab;
assign c7f1d0 = hgrant6_p & v3a6f3d9 | !hgrant6_p & v37650e3;
assign v37797ef = hgrant3_p & v8455e7 | !hgrant3_p & !v8455ab;
assign v376665a = hbusreq5_p & v376f56d | !hbusreq5_p & v376025f;
assign v3a66d50 = hbusreq2 & v3809516 | !hbusreq2 & v3a55b2d;
assign v374d95a = hmaster2_p & v3a6ffae | !hmaster2_p & v3a658bf;
assign v377cd0d = hbusreq2_p & v3a6bab2 | !hbusreq2_p & v3743b9e;
assign v3a6fbda = hbusreq5 & v3a5b289 | !hbusreq5 & v8455bb;
assign v3770690 = hbusreq5 & v3a6f3fa | !hbusreq5 & v3a5fc34;
assign v3a67d49 = hmaster1_p & v3a6dfb2 | !hmaster1_p & v377ce5a;
assign v3747a5f = hbusreq4 & v3a608b9 | !hbusreq4 & !v377163d;
assign v376e822 = hgrant5_p & v375b03c | !hgrant5_p & v3723e00;
assign v37729fa = hbusreq5 & v373ae6a | !hbusreq5 & v373ae4a;
assign v37795d9 = hlock5_p & v8455ab | !hlock5_p & v3750f20;
assign v37293d5 = hbusreq4 & v3a62f60 | !hbusreq4 & v3a63a66;
assign v377accc = hgrant4_p & v3a57f59 | !hgrant4_p & v3778567;
assign v3a6a1df = hgrant6_p & v1e37cd6 | !hgrant6_p & v3a71686;
assign v3a572d0 = hmaster2_p & v3a6ffca | !hmaster2_p & v3379037;
assign v373bce1 = hbusreq7_p & v375e33e | !hbusreq7_p & v373b571;
assign v374d13d = hmaster0_p & v8455ab | !hmaster0_p & v3a5c11a;
assign v375e973 = hbusreq6_p & v37577d7 | !hbusreq6_p & v8455b3;
assign v3774542 = hmaster0_p & v3a5e24e | !hmaster0_p & v37287be;
assign v376b5c0 = hgrant5_p & v3a6b078 | !hgrant5_p & v37786f9;
assign v3734d9a = hbusreq5_p & v3a70105 | !hbusreq5_p & v3749628;
assign v3762db3 = hbusreq6 & v377d4dc | !hbusreq6 & v3a66a6c;
assign v377ea01 = hbusreq6 & v375a750 | !hbusreq6 & v372a3cb;
assign v3a5e55e = hbusreq0 & a90ef2 | !hbusreq0 & v3749760;
assign v2ff8e5c = hmaster2_p & v3a70374 | !hmaster2_p & v3725827;
assign v37640e2 = hmaster0_p & v3a6fa7a | !hmaster0_p & v37362e9;
assign v375959a = hmaster2_p & v3739d88 | !hmaster2_p & v3757c7f;
assign v377fb9d = hbusreq3 & v3a696ed | !hbusreq3 & v8455ab;
assign v3a593ee = locked_p & v8455ab | !locked_p & v37386a9;
assign v3755b4e = hmaster2_p & v37429a1 | !hmaster2_p & v3a691eb;
assign v3a610f7 = hgrant7_p & v3a6fbcc | !hgrant7_p & v3767c3e;
assign v3a5c6d8 = hgrant6_p & v37517d2 | !hgrant6_p & !v3728621;
assign v377caa8 = hlock5 & v3a6b643 | !hlock5 & v1e377f7;
assign v372ad83 = jx1_p & v37766b2 | !jx1_p & v3a70f2c;
assign v376f6d1 = stateG10_1_p & v3a592f7 | !stateG10_1_p & v37526e0;
assign v3752def = hmaster1_p & v3a65540 | !hmaster1_p & v3a613da;
assign v3766b94 = hmaster2_p & v377ea20 | !hmaster2_p & v375dbf3;
assign v3752bbd = hmaster1_p & v376a2c0 | !hmaster1_p & v39ea663;
assign v377c22b = hmaster1_p & v3746c51 | !hmaster1_p & v375eac3;
assign v376f98e = hmaster3_p & v8455ab | !hmaster3_p & v3734279;
assign v3737c3f = hmaster2_p & v8a9c95 | !hmaster2_p & v3722a9c;
assign v3a6f528 = hbusreq5 & v3776bdf | !hbusreq5 & d7669b;
assign v377a975 = hmaster0_p & v8455e7 | !hmaster0_p & v3751369;
assign v3750b29 = hlock5 & v3757e93 | !hlock5 & v372713b;
assign v37747fc = hbusreq1_p & v37637db | !hbusreq1_p & v3769061;
assign v3a630bc = hbusreq7 & v3a55ab6 | !hbusreq7 & v3741b61;
assign v3a6ffd9 = hmaster0_p & v3a661fe | !hmaster0_p & v3a6eae9;
assign v3a567ea = hmaster1_p & v376891a | !hmaster1_p & v3a70cc7;
assign v3a6f1e8 = hmaster1_p & v3a635ea | !hmaster1_p & v3770aee;
assign v372e38f = hlock2 & v374cd48 | !hlock2 & v3757ae7;
assign v3a6f435 = hmaster1_p & v3778b48 | !hmaster1_p & v376c505;
assign v3773ce0 = hmaster2_p & v373014d | !hmaster2_p & v3763a20;
assign v3a6218f = hlock0 & v3a6bf41 | !hlock0 & v3a58cd4;
assign v374f319 = hbusreq0 & v3752aa5 | !hbusreq0 & v3744713;
assign v3a63172 = hbusreq6_p & v3759a21 | !hbusreq6_p & !v3a66a6e;
assign v3777e7d = hmaster2_p & v8455ab | !hmaster2_p & v374e855;
assign v3a5f218 = hmaster1_p & v3a6542a | !hmaster1_p & v8f1dd1;
assign v373b7c5 = hbusreq6_p & v3747302 | !hbusreq6_p & v3743b9e;
assign v3a70b87 = hmaster2_p & v35b774b | !hmaster2_p & v3a62826;
assign v3a6f97b = hbusreq4_p & v3a67d66 | !hbusreq4_p & v380714c;
assign v3a6f3f2 = hbusreq5_p & v3a5c73c | !hbusreq5_p & v3742623;
assign v37278fd = hbusreq5 & v373f911 | !hbusreq5 & v372d060;
assign v3a6f4ac = hbusreq3_p & v3747302 | !hbusreq3_p & v376c06f;
assign v377997c = jx1_p & v377c06f | !jx1_p & v3a6d8af;
assign v3a5dffe = hbusreq5 & v377997f | !hbusreq5 & v372b72d;
assign v3773eeb = hmaster0_p & v373cd03 | !hmaster0_p & v375bdcc;
assign v3a55b6c = stateG10_1_p & v3a70ecf | !stateG10_1_p & !v3a64566;
assign v37368d0 = jx1_p & v3774e9d | !jx1_p & v3a703b8;
assign v37681cc = hmaster2_p & v37433ef | !hmaster2_p & v8455ab;
assign v3a714b3 = hgrant2_p & v8455ab | !hgrant2_p & v3a53356;
assign v3809dcb = hmaster3_p & v3724e60 | !hmaster3_p & v3756da3;
assign v37420bb = hmaster2_p & v373f410 | !hmaster2_p & v373222d;
assign v3a6c80b = hbusreq2_p & v3a5e2ee | !hbusreq2_p & v3a704f8;
assign v3a606e6 = hmaster2_p & v8455ab | !hmaster2_p & !v3a70cc0;
assign v3a6fc21 = hbusreq0 & v374f9c5 | !hbusreq0 & v3a5ec91;
assign v3a71335 = hbusreq2_p & v3a6613e | !hbusreq2_p & v37510ae;
assign v3749e8a = hlock5 & v3747ea2 | !hlock5 & v373d955;
assign v3745072 = hbusreq5 & v374efb3 | !hbusreq5 & v8455ab;
assign v3759a4a = hmaster2_p & v372af77 | !hmaster2_p & v3a5b7db;
assign v37737aa = hgrant4_p & v8455e7 | !hgrant4_p & v37639c3;
assign v3765c70 = hmaster2_p & v376b4e1 | !hmaster2_p & !v3a709e2;
assign v2ff8c74 = hgrant4_p & v3772d6e | !hgrant4_p & adf1da;
assign v37314f0 = hmaster0_p & v376a14f | !hmaster0_p & v3a6fdbf;
assign v3806575 = hmaster0_p & v3736d47 | !hmaster0_p & v3a6817f;
assign v3a632e8 = hgrant2_p & v8455ba | !hgrant2_p & v3757c91;
assign v3757fa5 = hmaster1_p & v375b429 | !hmaster1_p & v37340b4;
assign v3a57f6c = hmaster2_p & v3a635ea | !hmaster2_p & v3747302;
assign v3759512 = hbusreq3_p & v8455ab | !hbusreq3_p & v3776a6e;
assign v3a703e0 = hgrant3_p & v3a59ffa | !hgrant3_p & v3a706b5;
assign v3a70d3a = hmaster2_p & v3a619c0 | !hmaster2_p & !v1e38224;
assign v3725f98 = hbusreq2_p & v3a6ff9b | !hbusreq2_p & !v3732bc1;
assign v3a66e5d = hgrant0_p & v372fc9d | !hgrant0_p & v375803a;
assign v3a69f4e = hmaster1_p & v3a56130 | !hmaster1_p & v91f9a4;
assign v375ca93 = hbusreq4 & v372dd09 | !hbusreq4 & v8455ab;
assign v37475be = hbusreq7_p & v3a6fd8a | !hbusreq7_p & !v3a7068f;
assign v3a66ca0 = hmaster0_p & v8455ab | !hmaster0_p & ba7f1c;
assign v3a6eff4 = hmaster2_p & v3a6909a | !hmaster2_p & v8455e7;
assign v3a6937a = hgrant4_p & v376d285 | !hgrant4_p & !v23fe329;
assign v3a5c65e = hbusreq0 & v37544cb | !hbusreq0 & v3732086;
assign v3a61517 = hgrant4_p & v3a6c5ee | !hgrant4_p & v3752cf6;
assign v376a967 = stateA1_p & v2aca977 | !stateA1_p & v3a70e3a;
assign v377839c = hmaster2_p & v37674f6 | !hmaster2_p & v3a70096;
assign v373732f = hmaster0_p & v3a639a2 | !hmaster0_p & v374677a;
assign v3730fd2 = hgrant3_p & v37645ec | !hgrant3_p & v3759470;
assign v3a5c366 = hbusreq3_p & v3a6eb0b | !hbusreq3_p & v37366d2;
assign v3a6887f = hbusreq6_p & v3758fc7 | !hbusreq6_p & v3a68c19;
assign v3a700b6 = hlock0 & v3748797 | !hlock0 & v372539e;
assign v3722e7a = hgrant6_p & v8455b0 | !hgrant6_p & b6390c;
assign v3a5f7c5 = hgrant4_p & v8455ab | !hgrant4_p & v3a6f994;
assign v3a5903a = hgrant0_p & v3a5b71a | !hgrant0_p & !v3776a6e;
assign v3a6f394 = hbusreq7_p & v3a71039 | !hbusreq7_p & v3a71675;
assign v39eb418 = hbusreq8_p & v375ea88 | !hbusreq8_p & v3746976;
assign v3769283 = hbusreq0_p & v374ab5b | !hbusreq0_p & v3760af0;
assign v3a7148d = hgrant1_p & v3743b9e | !hgrant1_p & v3a63621;
assign v1e377f7 = hmaster0_p & v3a6f7e9 | !hmaster0_p & v23fe28c;
assign v3738636 = hbusreq4_p & v3748609 | !hbusreq4_p & !v3732569;
assign v375c4e0 = hbusreq5 & v372893a | !hbusreq5 & v8455ab;
assign v37270b5 = hmaster1_p & v3a709ee | !hmaster1_p & v3a71273;
assign v3746ed6 = hmaster1_p & v3a57baa | !hmaster1_p & v373c23c;
assign v3724779 = hmaster2_p & v8455ab | !hmaster2_p & v377d27a;
assign v3770aee = hmaster0_p & v3a635ea | !hmaster0_p & v3763548;
assign v373aef5 = hbusreq4 & v3a70e2e | !hbusreq4 & !v3a55033;
assign v3a5b58e = hmaster1_p & v376ed2b | !hmaster1_p & v3a701bc;
assign d09db6 = hbusreq5 & v377a470 | !hbusreq5 & v357742d;
assign v3a7070c = hbusreq5 & v374da93 | !hbusreq5 & v8455ab;
assign v3a6c44c = hgrant4_p & v8455ab | !hgrant4_p & v3a66f3e;
assign v372d967 = hgrant6_p & v8455c9 | !hgrant6_p & v376b57e;
assign v3807dc9 = hbusreq5 & v3a67092 | !hbusreq5 & v8455ab;
assign v3739934 = hmaster2_p & v3755002 | !hmaster2_p & v3a5600a;
assign v3744aa9 = hmaster0_p & v3a703f2 | !hmaster0_p & v3a701e0;
assign v3a7058c = jx0_p & v3a6ff55 | !jx0_p & v374da33;
assign v3a6eb02 = hmaster0_p & v37721fa | !hmaster0_p & v376a6f1;
assign v3a706f0 = hgrant5_p & v8455ab | !hgrant5_p & v372fb63;
assign v3a62cda = hgrant5_p & v3a53d98 | !hgrant5_p & v376eef5;
assign v37287e1 = hmaster2_p & v3763a86 | !hmaster2_p & v3730986;
assign v372ead5 = hbusreq2_p & v3a6d621 | !hbusreq2_p & v3a63597;
assign v3a6f7b9 = hbusreq5_p & v3756b5c | !hbusreq5_p & v3a5604a;
assign v3a6faf3 = hmaster2_p & v380974c | !hmaster2_p & v37678fc;
assign v373ff97 = hmaster0_p & v37363f8 | !hmaster0_p & !v937864;
assign v374a075 = hmaster2_p & v3746c51 | !hmaster2_p & v3a70893;
assign v376204f = hmaster0_p & v3a6d040 | !hmaster0_p & v374f6f9;
assign v38074bc = hbusreq6 & v376bfc3 | !hbusreq6 & v3766e4a;
assign v377bc9c = hbusreq0 & v375ee2a | !hbusreq0 & v373f2d1;
assign v37382eb = hmaster2_p & v8455b9 | !hmaster2_p & !v8455ab;
assign v3a6c527 = hmaster1_p & v376891a | !hmaster1_p & v375b389;
assign v3774f24 = hgrant4_p & v8455ab | !hgrant4_p & v37443b5;
assign v3a70f04 = hbusreq3_p & v377b4f7 | !hbusreq3_p & v8455ab;
assign v3a7044c = hbusreq1_p & v373ae2e | !hbusreq1_p & !v3733350;
assign v377609a = hbusreq8_p & v3750d4d | !hbusreq8_p & v37255e9;
assign v377988b = hbusreq4_p & v3769374 | !hbusreq4_p & v3755e97;
assign v3a60642 = hmaster1_p & v374b7d8 | !hmaster1_p & v3a56200;
assign v3727a04 = hmaster1_p & v374a9d0 | !hmaster1_p & v3a6f449;
assign v373927b = hbusreq5_p & v3a706bd | !hbusreq5_p & !v3768e52;
assign v373330f = hbusreq0 & v37748b2 | !hbusreq0 & v3a702e8;
assign v37765cf = hmaster2_p & v37624a2 | !hmaster2_p & v8455ab;
assign v3a58761 = hmaster0_p & v374f0c1 | !hmaster0_p & v3774c98;
assign v3778674 = hbusreq8 & v374244e | !hbusreq8 & v375da52;
assign v3770c0d = hbusreq8 & v373bbce | !hbusreq8 & v8455ab;
assign v377bf21 = hbusreq5_p & v3777f05 | !hbusreq5_p & v3a706f6;
assign v374eaeb = hbusreq0 & v3772513 | !hbusreq0 & v8455ab;
assign v375075b = hgrant5_p & v3a60509 | !hgrant5_p & v373ec83;
assign v3a6fe5f = hbusreq5_p & v3a70e45 | !hbusreq5_p & v3726a7e;
assign v377740c = jx0_p & v3730862 | !jx0_p & v37287fa;
assign v3a70a78 = hbusreq5 & v37280b2 | !hbusreq5 & v377cebd;
assign v3738f36 = jx0_p & v374f003 | !jx0_p & v3a6f6f0;
assign v3a6f9e5 = hlock4 & v3748797 | !hlock4 & v372fc07;
assign v3742472 = hmaster3_p & v37629ba | !hmaster3_p & !v374e02b;
assign v3a6f6d1 = hmaster1_p & v3a58218 | !hmaster1_p & v37350c3;
assign v3a7033d = hbusreq6_p & v3a6ebaf | !hbusreq6_p & !v8455ab;
assign v374220d = hgrant4_p & v1e37d8b | !hgrant4_p & v28896e3;
assign v23fdadd = hmaster0_p & v376a14f | !hmaster0_p & v3764ec5;
assign v3755b56 = hbusreq4_p & v3a5f974 | !hbusreq4_p & v8455ab;
assign v3750d4d = hbusreq7_p & v3756087 | !hbusreq7_p & v3751aab;
assign v3774e33 = hmaster0_p & v3a6fe22 | !hmaster0_p & v374fe44;
assign v374fe51 = hmaster1_p & v376e72d | !hmaster1_p & v3a6fc67;
assign v3725c13 = hbusreq5 & v8455c7 | !hbusreq5 & !v8455ab;
assign v374f5d6 = hmaster0_p & v372f309 | !hmaster0_p & v377b460;
assign v3a7007c = hbusreq8 & v3a5e388 | !hbusreq8 & v8455bb;
assign v3726991 = hmaster2_p & v3a6f1ab | !hmaster2_p & v8455ab;
assign v1e3732b = hbusreq6_p & v3808870 | !hbusreq6_p & v37474e8;
assign v3730118 = hgrant4_p & v3a624da | !hgrant4_p & !v372dfc1;
assign v3772362 = hbusreq6_p & v3a70cf0 | !hbusreq6_p & v1e37cab;
assign v3a53eeb = hbusreq4_p & v3a6f2a8 | !hbusreq4_p & !v8455ab;
assign v375ac12 = hbusreq5_p & v37290ab | !hbusreq5_p & v375210d;
assign v3726d60 = hmaster1_p & v3734967 | !hmaster1_p & v3a58182;
assign v2acb5c8 = hmaster1_p & v3755002 | !hmaster1_p & v3743327;
assign v3a5fd4a = hmaster2_p & v375d887 | !hmaster2_p & v3771758;
assign v3773015 = hbusreq5 & v3a711bd | !hbusreq5 & v37682d5;
assign v373cd5d = hmaster0_p & v37356f0 | !hmaster0_p & v3a7161f;
assign v3735417 = hbusreq4_p & v35b774b | !hbusreq4_p & v9ed516;
assign v3258db3 = hbusreq2 & v3750866 | !hbusreq2 & v375cf36;
assign v3748529 = stateA1_p & v2aca977 | !stateA1_p & v376a35c;
assign v376233b = hready_p & v374c144 | !hready_p & v3a64c73;
assign v3729382 = hmaster0_p & v3755539 | !hmaster0_p & v3a296dc;
assign v37304a2 = hready_p & v3737186 | !hready_p & v373da11;
assign v374d7dc = hbusreq5_p & v3a6b73b | !hbusreq5_p & v3a6f948;
assign v3a62415 = hbusreq4_p & v89a0d1 | !hbusreq4_p & v8455ab;
assign v374bba3 = hbusreq5_p & v3770b26 | !hbusreq5_p & v377f734;
assign v3728bd6 = hmaster3_p & v37670b6 | !hmaster3_p & v374e463;
assign v3a5a7fd = hbusreq2_p & v3747302 | !hbusreq2_p & v3806e34;
assign v3a66123 = hgrant6_p & v8455ab | !hgrant6_p & v3a6e9b8;
assign v3a6fb7a = hbusreq6 & v372f74f | !hbusreq6 & v8455ab;
assign v3774647 = hgrant4_p & v8455ab | !hgrant4_p & v375b626;
assign v3a70ba9 = hmaster2_p & v376c248 | !hmaster2_p & v3a61cd7;
assign v374f0ac = hlock5 & v3763e30 | !hlock5 & v3a66aa6;
assign v3a70ef2 = hbusreq0_p & v38072fd | !hbusreq0_p & v3a6430c;
assign v374978c = hlock2_p & v372eada | !hlock2_p & !v8455ab;
assign v37701fd = hgrant6_p & v3724475 | !hgrant6_p & v3731099;
assign v3728760 = hgrant1_p & v374721d | !hgrant1_p & v37665bf;
assign v3a70d79 = hlock6_p & v3a607af | !hlock6_p & v373aaa8;
assign v374c6ff = hmaster0_p & v3a5e846 | !hmaster0_p & v3731d67;
assign v3779925 = hlock0 & v3a6f994 | !hlock0 & v377a180;
assign v37778cf = hbusreq6 & v373e2c3 | !hbusreq6 & v8455e7;
assign c35240 = hbusreq4_p & v37684a8 | !hbusreq4_p & v3a6a1df;
assign v3a70c75 = hmaster2_p & v3a635ea | !hmaster2_p & v37476bd;
assign v377e85e = hlock1_p & v3741500 | !hlock1_p & !v8455b6;
assign v3a6f696 = hbusreq6 & v3746c51 | !hbusreq6 & v8455ab;
assign v375c505 = hbusreq6 & v3756e01 | !hbusreq6 & v3a666e8;
assign d8a786 = hgrant6_p & v377f21b | !hgrant6_p & v3736cdb;
assign v3a6a678 = hmaster2_p & v37234c3 | !hmaster2_p & !v3775537;
assign v3a6fc54 = hgrant2_p & v8455ab | !hgrant2_p & v3a7010f;
assign v3749d78 = hgrant6_p & v373d4ff | !hgrant6_p & v37452c7;
assign v37686c1 = hgrant3_p & v8455be | !hgrant3_p & v3a6fdd0;
assign v37390f0 = hbusreq5 & v372d1f0 | !hbusreq5 & v3a705c7;
assign v374262b = hgrant6_p & v8455ca | !hgrant6_p & v3773390;
assign v3730389 = hbusreq5 & v373a4e4 | !hbusreq5 & v3a70d99;
assign v3758e8d = hmaster1_p & v3a55d4c | !hmaster1_p & !v375ecab;
assign d2afa4 = hmaster0_p & v37469c4 | !hmaster0_p & v37767fa;
assign v3744940 = hbusreq8 & v38092a9 | !hbusreq8 & v3a70555;
assign v3774c55 = hmaster0_p & v3747b81 | !hmaster0_p & v3a6fc05;
assign v3738a45 = hmaster3_p & v37318cb | !hmaster3_p & v3a6ffc5;
assign v3a6152c = hgrant4_p & v3742241 | !hgrant4_p & v374d970;
assign v3a59746 = hmaster0_p & v3a67577 | !hmaster0_p & v3762ba2;
assign v3a6de93 = hmaster2_p & v3757765 | !hmaster2_p & v374f0f5;
assign v373cb2d = hbusreq2 & v3760f4e | !hbusreq2 & v8455b3;
assign v3777baa = hgrant0_p & v37773a9 | !hgrant0_p & v3777e08;
assign v37290fa = hbusreq7 & v37375ed | !hbusreq7 & v3767483;
assign v3728f0a = hbusreq7_p & v374fe51 | !hbusreq7_p & v372fd4a;
assign v374449e = hgrant4_p & v3a6fe35 | !hgrant4_p & v3a6f874;
assign baea86 = hgrant4_p & v8455ab | !hgrant4_p & v3747114;
assign v3a6fa62 = hmaster0_p & v3773950 | !hmaster0_p & v3a6af83;
assign v3759daf = hlock2_p & v375d25d | !hlock2_p & !v8455ab;
assign v3a6d4f8 = hmaster1_p & v8455ab | !hmaster1_p & v3a66cad;
assign v2acb0c1 = stateG10_1_p & v35b9d52 | !stateG10_1_p & v3733ea2;
assign v3a6f7b0 = hbusreq4_p & v3a6008f | !hbusreq4_p & v8455ab;
assign v3a6851f = hbusreq4 & v3a714b1 | !hbusreq4 & v8455ab;
assign v3a618b3 = hbusreq2 & v376a34d | !hbusreq2 & v3a5b2fd;
assign v3729c6b = hlock2_p & v3a704f3 | !hlock2_p & v8455e7;
assign v3763e55 = hmaster2_p & v3770b26 | !hmaster2_p & v372fd5d;
assign v3722b64 = hbusreq2 & v37660d2 | !hbusreq2 & v3a6f70d;
assign v377a3bd = hgrant4_p & v3a70aeb | !hgrant4_p & v3a64190;
assign v37775d9 = hgrant0_p & v9ed516 | !hgrant0_p & v373eedf;
assign v3724e4b = hmaster0_p & v375930e | !hmaster0_p & v3760f64;
assign v3a6eee2 = hbusreq8 & v3a5544e | !hbusreq8 & v8455ab;
assign v3a6f443 = hbusreq4_p & v3a5c945 | !hbusreq4_p & v3a57f59;
assign v3723ba5 = hbusreq4_p & v3a5585e | !hbusreq4_p & v8455ab;
assign v372b27e = hmaster0_p & v3a62c11 | !hmaster0_p & v37614c1;
assign v37485f0 = hgrant0_p & v3733e9e | !hgrant0_p & v375da3a;
assign v35772dd = hmaster3_p & v3739cdb | !hmaster3_p & v3763ca5;
assign v3723e5f = hmastlock_p & v376df43 | !hmastlock_p & v8455ab;
assign v380910e = hlock8 & v3745941 | !hlock8 & v376957a;
assign v9c0027 = hmaster2_p & v3a5ddc1 | !hmaster2_p & v3769740;
assign d1375e = hmaster0_p & v1e382e7 | !hmaster0_p & !v374b13e;
assign v3a67d8d = hgrant4_p & v3763209 | !hgrant4_p & v373d10f;
assign v376f017 = hmaster0_p & v3a6ff35 | !hmaster0_p & v3747666;
assign v3744fa5 = hbusreq3 & v1e38224 | !hbusreq3 & v8455ab;
assign v3739e31 = hbusreq5_p & v3745072 | !hbusreq5_p & v8455ab;
assign v3a71215 = hmaster0_p & v3739698 | !hmaster0_p & !v373e267;
assign v3a712d0 = hmaster2_p & v8455ab | !hmaster2_p & v375ecd5;
assign v374fe44 = hmaster2_p & v3745539 | !hmaster2_p & v8455bb;
assign v3760700 = hbusreq4_p & v3769dfe | !hbusreq4_p & v8455ab;
assign v37643eb = hgrant2_p & v3a6fd27 | !hgrant2_p & v3a67d59;
assign v3a6fe09 = hmaster2_p & v8455ab | !hmaster2_p & v376e9e9;
assign v3762a54 = hbusreq5_p & v3747453 | !hbusreq5_p & v3751285;
assign v37294f4 = hgrant7_p & v376faf9 | !hgrant7_p & !v8455ab;
assign v376e4c5 = hbusreq7_p & v374763e | !hbusreq7_p & v3778211;
assign v3746b91 = hlock7_p & v377e851 | !hlock7_p & v3a63cf3;
assign v374a97c = hbusreq6_p & v3766a28 | !hbusreq6_p & !v8455ab;
assign v374b4f8 = hbusreq5 & v373794a | !hbusreq5 & v3a6ff12;
assign v3737265 = hbusreq8 & v374ffb8 | !hbusreq8 & v3769a6c;
assign v3a632f4 = hbusreq2_p & v37666bd | !hbusreq2_p & v3a699d3;
assign v373f880 = hgrant4_p & v8455ab | !hgrant4_p & v375bd0e;
assign v376ab01 = hlock0 & v37285eb | !hlock0 & v372f759;
assign v375ec98 = hgrant6_p & v3a5a63c | !hgrant6_p & v3a5aee5;
assign v374b07b = hbusreq1 & v8455ab | !hbusreq1 & v8455b0;
assign v375add0 = hlock4 & v3a6fba9 | !hlock4 & v37572f7;
assign v3a6eec4 = hmaster0_p & v37453dd | !hmaster0_p & v3766573;
assign v3754e7b = hgrant0_p & v376bb26 | !hgrant0_p & v372998c;
assign v3a56e53 = hmaster0_p & v3a5b8b9 | !hmaster0_p & v3a6a197;
assign v372e3b4 = hmaster2_p & v374f138 | !hmaster2_p & !v8455ab;
assign v372cd45 = hbusreq3 & v3a6fd17 | !hbusreq3 & v8455ab;
assign v35772a2 = hbusreq2_p & v1e37932 | !hbusreq2_p & v8455ab;
assign v3a539bf = hmaster2_p & v8455ab | !hmaster2_p & v3a70b1e;
assign v3a6f4d7 = hmaster0_p & v3778083 | !hmaster0_p & v375eb99;
assign v373ac67 = hbusreq4 & v3a71314 | !hbusreq4 & v8455ab;
assign v3a70484 = hmaster0_p & v3773666 | !hmaster0_p & v3a6f3cd;
assign v373b2ce = hbusreq3_p & v37675e2 | !hbusreq3_p & v3a70d90;
assign v3a71379 = hbusreq2 & v3a5b68a | !hbusreq2 & !v8455ab;
assign v377152e = hbusreq4_p & v37c006d | !hbusreq4_p & v37759b6;
assign v3761d06 = hbusreq4 & v377cd6c | !hbusreq4 & v8455ab;
assign v3765b5a = hbusreq7 & v845765 | !hbusreq7 & v8455ab;
assign v3746e85 = hgrant4_p & v376495e | !hgrant4_p & v3a6995c;
assign v3743f47 = hgrant3_p & v37669b4 | !hgrant3_p & v37244e7;
assign v3a5bc77 = hbusreq6 & v374f351 | !hbusreq6 & v39a4e43;
assign v372f3f1 = hbusreq0 & v37299fa | !hbusreq0 & v37436cf;
assign v3a70877 = hmaster1_p & v376d287 | !hmaster1_p & v1e37561;
assign v3a6ef61 = hgrant5_p & v3a62c28 | !hgrant5_p & v3a70c37;
assign v37446e0 = hgrant5_p & v3a6f555 | !hgrant5_p & v37356aa;
assign v3735f9b = hlock6_p & v8455ab | !hlock6_p & a69e17;
assign v37640fd = hbusreq6_p & v37535e7 | !hbusreq6_p & v3736a9a;
assign v3a5e1ab = hlock4_p & v375d9f8 | !hlock4_p & v8455b3;
assign v3767080 = hmaster0_p & v374e0e9 | !hmaster0_p & v3751b35;
assign v3757044 = hbusreq5_p & v37531fd | !hbusreq5_p & v3a70dfc;
assign v3a64fce = hbusreq5_p & v2619aa7 | !hbusreq5_p & v3a5a37a;
assign v3761df7 = hmaster2_p & v373014d | !hmaster2_p & v377caa3;
assign v37457fb = locked_p & v8455ab | !locked_p & !v39a5381;
assign v3750c27 = hgrant4_p & v8455ab | !hgrant4_p & v376c2a1;
assign v3a6fb8d = hmaster0_p & v3759031 | !hmaster0_p & v372ef80;
assign v373dde1 = hmaster0_p & v8455ab | !hmaster0_p & v3a64987;
assign v3745dac = hgrant0_p & v3808553 | !hgrant0_p & v373eedf;
assign v377439e = hmaster0_p & v376d550 | !hmaster0_p & v377e004;
assign v3a6f96e = hmaster0_p & v37693ce | !hmaster0_p & !v373b59f;
assign v2acaf74 = hbusreq3 & v375f52b | !hbusreq3 & v8455ab;
assign v372cf41 = hlock8_p & v3746f89 | !hlock8_p & !v8455ab;
assign v373594b = hmaster2_p & v3a6fd7b | !hmaster2_p & v37453f0;
assign v37598c6 = hgrant0_p & v37773a9 | !hgrant0_p & ad2d05;
assign cbb40b = hbusreq0 & v3a7035f | !hbusreq0 & v3a69bbf;
assign v376e7e8 = hlock4_p & v8455ab | !hlock4_p & v375c845;
assign v929796 = hgrant2_p & v8455ab | !hgrant2_p & v375ef1e;
assign v3a701e0 = hmaster2_p & v375d263 | !hmaster2_p & v3a60b88;
assign v3a58429 = hbusreq0_p & v374362e | !hbusreq0_p & v8455ab;
assign v3a57db6 = hmaster0_p & v1e37d82 | !hmaster0_p & v8455ab;
assign v3a5a381 = hmaster0_p & v3a71678 | !hmaster0_p & v3756aaa;
assign v37603d4 = hbusreq5_p & v374b035 | !hbusreq5_p & v376b2a3;
assign v3a60509 = hmaster1_p & v374851a | !hmaster1_p & v3a6fa7c;
assign v3751d41 = hmaster0_p & v37770f5 | !hmaster0_p & v374e0a9;
assign v3a6ad38 = hbusreq0 & v3a7151e | !hbusreq0 & v3a7018a;
assign v375a00a = hbusreq2 & v376b6c9 | !hbusreq2 & b755d3;
assign v3750f60 = hmaster2_p & v1e38224 | !hmaster2_p & !v3a59e87;
assign v3a71031 = jx0_p & v372a64f | !jx0_p & v375b84e;
assign v3a56687 = hbusreq5_p & v377451f | !hbusreq5_p & v3a5ba93;
assign v3806b2d = hlock5 & v3770322 | !hlock5 & v3a7136b;
assign v3a5689e = hbusreq3_p & v373014d | !hbusreq3_p & !v8455ab;
assign v3736c8d = hlock6 & v37685ea | !hlock6 & v3a6f0fd;
assign v374c9e9 = hmaster0_p & v3775f0b | !hmaster0_p & v3757966;
assign v376f4c5 = hmaster0_p & v372da78 | !hmaster0_p & v375820e;
assign v3a5fd0a = hmaster0_p & v8455ab | !hmaster0_p & v377529a;
assign v376b374 = hmaster0_p & v3a6e6c2 | !hmaster0_p & v3777536;
assign v3a70894 = hmaster0_p & dafc4e | !hmaster0_p & v375d42d;
assign v372a652 = hgrant5_p & v3a5aef8 | !hgrant5_p & v374a9db;
assign v375dc9b = hmaster2_p & v3807aa1 | !hmaster2_p & !v375a67c;
assign v3772b7e = hbusreq4_p & v3a68f04 | !hbusreq4_p & v3a60f18;
assign v3765cfd = hbusreq0_p & v373e67e | !hbusreq0_p & v3a70e52;
assign v372dec3 = hbusreq4 & v376ba2e | !hbusreq4 & v3770234;
assign v377ce5a = hmaster0_p & v3a6dfb2 | !hmaster0_p & v372f006;
assign v3773c70 = hmaster0_p & v375e8aa | !hmaster0_p & !v3755914;
assign v375c5a1 = hbusreq1_p & v3a711f1 | !hbusreq1_p & !v8455ab;
assign v375e183 = hmaster2_p & v3a5952d | !hmaster2_p & v372cc25;
assign v3737c21 = jx1_p & v380a20c | !jx1_p & v372a9c2;
assign v377b3d5 = hgrant5_p & v8455ab | !hgrant5_p & v3738da4;
assign v3a7010b = hmaster0_p & v377d596 | !hmaster0_p & v377e004;
assign v375c4cb = hmaster2_p & v373d9e0 | !hmaster2_p & v374b526;
assign v37246f1 = hlock0_p & v37317a9 | !hlock0_p & v3a70dfb;
assign v3a7013a = hbusreq5 & v3a5f451 | !hbusreq5 & v3760bda;
assign v360d0c7 = hmaster0_p & v376f70a | !hmaster0_p & v3a56512;
assign v374de43 = hmaster0_p & v3736d47 | !hmaster0_p & v3a6f6a9;
assign v3759144 = hmaster0_p & v3a62a6d | !hmaster0_p & v372754b;
assign v374ebbf = hbusreq8 & v3749fc1 | !hbusreq8 & v3734d20;
assign v375bb92 = hbusreq4_p & v3a6f8f5 | !hbusreq4_p & v375c334;
assign v374deba = hbusreq8 & v376c69d | !hbusreq8 & v3a63ac4;
assign v3a6f77e = hlock2 & v377b27b | !hlock2 & v37599cb;
assign v376b220 = hmaster1_p & v3a69913 | !hmaster1_p & v376d215;
assign v374c052 = hgrant6_p & v3a5a510 | !hgrant6_p & v3a6eb4a;
assign v3a6022f = hlock7 & v37431ce | !hlock7 & v375df28;
assign v3a70478 = hmaster0_p & v377181f | !hmaster0_p & !v373a3c8;
assign v377c125 = hmaster2_p & v373891b | !hmaster2_p & v377b030;
assign v3a6fdb6 = hmaster0_p & v377234d | !hmaster0_p & b8f82c;
assign v377e1f6 = hbusreq6_p & v3a65da7 | !hbusreq6_p & v37338d8;
assign v3a63fd5 = hbusreq8 & v3a61661 | !hbusreq8 & v374f6c0;
assign v3a6fbcc = jx1_p & v3739a33 | !jx1_p & v8455ab;
assign v37532a8 = hmaster1_p & v8455ab | !hmaster1_p & v3a7009f;
assign v3a5d90a = hgrant2_p & v374f617 | !hgrant2_p & v3752511;
assign v372cede = hgrant2_p & v375e7cc | !hgrant2_p & v360d109;
assign v3a6a374 = hbusreq0 & v3a6f430 | !hbusreq0 & v3a6fa5c;
assign v374a9e4 = hbusreq5_p & v3a6f6c0 | !hbusreq5_p & v3a70786;
assign v373aca2 = hbusreq0 & v3768202 | !hbusreq0 & !v8455ab;
assign v3731d75 = hbusreq4_p & v3733e9e | !hbusreq4_p & v1e38224;
assign v3775144 = hbusreq4 & v3730bf9 | !hbusreq4 & v373b687;
assign v375a4a9 = hbusreq7_p & v3a6af87 | !hbusreq7_p & v8455ab;
assign v3a6ebd4 = jx0_p & v3a704e0 | !jx0_p & v375dfc6;
assign v377dfa2 = hlock5_p & a7b390 | !hlock5_p & v3a6f674;
assign v375c2b1 = hlock6_p & v3757684 | !hlock6_p & v377167e;
assign v375b597 = hmaster1_p & v3778c64 | !hmaster1_p & v3a70cf4;
assign v373ea00 = hbusreq7 & v3a6f5e9 | !hbusreq7 & v3a605d3;
assign v3774b2b = hmaster2_p & v3a705f2 | !hmaster2_p & v375981e;
assign v38065aa = hgrant3_p & v37655d3 | !hgrant3_p & v3730cda;
assign ca602f = hlock3 & v3769605 | !hlock3 & v3a559f0;
assign v3766025 = hlock4_p & v374f78c | !hlock4_p & v3748e81;
assign v373346a = hbusreq5 & v377ac0f | !hbusreq5 & !v8455ab;
assign v374572e = hbusreq0 & v372d86a | !hbusreq0 & v3a7035a;
assign v374a262 = hbusreq7 & v375269c | !hbusreq7 & v3725a6e;
assign v3730452 = hbusreq3 & v3734046 | !hbusreq3 & v3774a8f;
assign v3737700 = hmaster1_p & v372d905 | !hmaster1_p & v374a650;
assign v3730de9 = hgrant1_p & v3764276 | !hgrant1_p & v3750746;
assign v3a5c59f = hbusreq4 & v375331e | !hbusreq4 & !v3a640a0;
assign v3a70514 = hbusreq4 & v373c7a5 | !hbusreq4 & v374829e;
assign v374d2b3 = hgrant2_p & v8455ab | !hgrant2_p & v3a6eb6b;
assign v3a7098f = hmaster0_p & v372c221 | !hmaster0_p & d1e3dd;
assign v3a69ac0 = hlock0_p & v3a70641 | !hlock0_p & v8455b0;
assign v3a6fc89 = hmaster0_p & a012c1 | !hmaster0_p & v377eee2;
assign v3a6f773 = hbusreq8_p & v37271fd | !hbusreq8_p & v23fde66;
assign v3a6a893 = hbusreq8_p & v3a6cbfa | !hbusreq8_p & v375c67c;
assign v374077c = hmaster2_p & v37693af | !hmaster2_p & v37319d5;
assign v3a6f04e = hmaster2_p & v3733e9e | !hmaster2_p & v376ea4a;
assign v3a6b6f2 = hmaster0_p & v3a63111 | !hmaster0_p & !v372ee6a;
assign v3779c26 = hmaster1_p & v8455ab | !hmaster1_p & v37299dc;
assign v3a66f8d = hbusreq5 & a65142 | !hbusreq5 & v3769740;
assign v3a6ad04 = hbusreq6_p & v377550d | !hbusreq6_p & v3a58102;
assign v2ff8e9c = hbusreq4_p & v37652cb | !hbusreq4_p & v3a5f9e6;
assign v375e647 = hbusreq0 & v3751db5 | !hbusreq0 & v3a70b00;
assign v3751b6b = hbusreq8_p & v373f262 | !hbusreq8_p & v377f3ba;
assign v375a025 = jx0_p & v374c22d | !jx0_p & v9f56fd;
assign v372f320 = jx3_p & v3a5f375 | !jx3_p & !v377a9fc;
assign v3a6f365 = hbusreq0 & v375c7a9 | !hbusreq0 & v8455ab;
assign v3a6305e = hbusreq2_p & v3a5e7a5 | !hbusreq2_p & v3761865;
assign v372a55a = hbusreq5 & v3740bce | !hbusreq5 & v374ef20;
assign v3a6f674 = hmaster0_p & v3a5b289 | !hmaster0_p & v3728e89;
assign v375c6c7 = hgrant3_p & v377dd3b | !hgrant3_p & v3a55347;
assign v3761fda = hmaster2_p & v3a6c4e4 | !hmaster2_p & !v377d1a3;
assign v3776bb6 = hbusreq6_p & v3742370 | !hbusreq6_p & v3758e68;
assign v3738c45 = hbusreq6_p & v3a5457f | !hbusreq6_p & v3a632e8;
assign v3742f0b = hmaster2_p & v3733d6e | !hmaster2_p & v372493b;
assign v3728eca = hmaster0_p & v377b096 | !hmaster0_p & v3a7026a;
assign v3a5982a = hmaster0_p & v3a635ea | !hmaster0_p & v376ba2b;
assign v38087ee = hmaster2_p & v372ee7e | !hmaster2_p & !v3a6febd;
assign v3755296 = hgrant3_p & v37506fb | !hgrant3_p & v3a5ea7b;
assign v3a70cd1 = hbusreq6 & v376b88d | !hbusreq6 & v3a70d99;
assign v3729e32 = hgrant6_p & v3756057 | !hgrant6_p & v3a67dbc;
assign v376f0c2 = hbusreq7_p & v380929f | !hbusreq7_p & v375c691;
assign v3771431 = hbusreq8_p & v3a635ea | !hbusreq8_p & v373a36a;
assign v375b3af = hbusreq3_p & v3a635ea | !hbusreq3_p & v3734fa9;
assign v374151e = jx2_p & v37315ae | !jx2_p & v3741172;
assign v3773f88 = hmaster2_p & v8455e7 | !hmaster2_p & v3a696ed;
assign v37556c1 = hbusreq5 & v3771ddb | !hbusreq5 & v377011b;
assign v3a6dd22 = hbusreq5 & v376a6f1 | !hbusreq5 & v3761a8f;
assign v3a6667c = hbusreq8 & v23fde9c | !hbusreq8 & v376f37e;
assign v3726111 = hbusreq8_p & v375d36b | !hbusreq8_p & v375a55d;
assign v3a71554 = hlock4_p & v375444e | !hlock4_p & v8455b0;
assign v374b747 = hbusreq5_p & v372b60b | !hbusreq5_p & v3750b86;
assign v3a710b5 = hbusreq3 & v374f307 | !hbusreq3 & v8455ab;
assign v3724398 = hmaster2_p & v374306c | !hmaster2_p & !v376e914;
assign v377e582 = hgrant2_p & v3a5c823 | !hgrant2_p & v37526a0;
assign v37683f8 = hmaster3_p & v37701a5 | !hmaster3_p & v3760251;
assign v372f73c = hbusreq2 & v3a6773a | !hbusreq2 & v35b774b;
assign v3756918 = hgrant6_p & v8455ab | !hgrant6_p & v3a65f7a;
assign v3a55f2b = hbusreq4 & v37413b6 | !hbusreq4 & v3a6eb47;
assign v374ed99 = hlock6 & v376f9b5 | !hlock6 & v3a6f30f;
assign v37237f1 = hbusreq5_p & v373d943 | !hbusreq5_p & v377e056;
assign v3a617a6 = hmaster2_p & v3a7024f | !hmaster2_p & v3748d67;
assign v3a6225d = hbusreq5 & v3a712c0 | !hbusreq5 & v374b42b;
assign v375b0ad = hmaster0_p & v37350f0 | !hmaster0_p & v3a70388;
assign v374da36 = hgrant6_p & v3770559 | !hgrant6_p & v3757a13;
assign v372c134 = hbusreq3 & v3a66b2b | !hbusreq3 & v376c8ea;
assign v373e1fb = hlock5 & v3a650a6 | !hlock5 & v375a6e8;
assign v1e374ce = hlock4 & v37264c9 | !hlock4 & v375a166;
assign v377a9fc = jx1_p & v380a20c | !jx1_p & v3732be9;
assign v3768274 = hmaster1_p & v3779595 | !hmaster1_p & v3743017;
assign v3a5dec3 = hmaster0_p & v3a6fe0d | !hmaster0_p & v3a6f22a;
assign v3a6f427 = hmaster2_p & v376d9ad | !hmaster2_p & v37270d9;
assign v374e459 = hbusreq2 & v3745053 | !hbusreq2 & !v8455b3;
assign v3a70f8f = hbusreq4_p & v3a634db | !hbusreq4_p & v3809240;
assign v3a7076e = hmaster2_p & v37297cb | !hmaster2_p & v377e889;
assign v377c79a = hlock5_p & v3a5a854 | !hlock5_p & v377dc65;
assign v375620b = hmaster0_p & v373b48c | !hmaster0_p & v3a714d5;
assign v37c023b = hbusreq4_p & v3743b98 | !hbusreq4_p & v8455b7;
assign v360bedd = hbusreq5 & v3731d8f | !hbusreq5 & v37759a7;
assign v3a695a8 = hmaster0_p & v375fd99 | !hmaster0_p & v376b540;
assign v37717ac = hgrant6_p & v38075aa | !hgrant6_p & v8455ab;
assign v3771ea6 = hlock2_p & v3a6ebb0 | !hlock2_p & v373086c;
assign v37739ed = hmaster0_p & v3736539 | !hmaster0_p & !v8455ab;
assign v3a674d5 = hmaster3_p & v373ca17 | !hmaster3_p & v3a6fbc6;
assign v376d98d = hgrant4_p & v3743de6 | !hgrant4_p & v3a69ca2;
assign v373d2e0 = stateG2_p & v8455ab | !stateG2_p & v37643ee;
assign v3775dbc = hbusreq6_p & v377c77a | !hbusreq6_p & v8455b0;
assign v3a62d18 = hlock6_p & v372391f | !hlock6_p & v375e60f;
assign v3729030 = hlock4 & v1e37556 | !hlock4 & v31c369c;
assign v37711f0 = hlock5 & v35b85ad | !hlock5 & v3a6eb1c;
assign v37765d0 = hgrant6_p & v372abd8 | !hgrant6_p & v3764e95;
assign v3766ff3 = hmaster0_p & aa421e | !hmaster0_p & v376d060;
assign v3739d23 = hmaster2_p & v3736026 | !hmaster2_p & v374eedb;
assign v3732939 = hbusreq6_p & v3a5acca | !hbusreq6_p & v8455ab;
assign v3769dfe = hbusreq4 & v3734e58 | !hbusreq4 & v8455ab;
assign v3739b37 = hbusreq5 & v3735272 | !hbusreq5 & v1e37b76;
assign v3756de7 = hmaster2_p & v3a6fe0d | !hmaster2_p & v3754ec1;
assign v372a1bd = hlock7_p & v3a6f5ff | !hlock7_p & !v23fd8b7;
assign v3a67462 = hmaster2_p & v373014d | !hmaster2_p & v374b077;
assign v376456d = hmaster2_p & v3a635ea | !hmaster2_p & v37c3782;
assign v3a6f5d4 = hmaster0_p & v8455b9 | !hmaster0_p & v37382eb;
assign v3a63f77 = hbusreq8_p & v372dc20 | !hbusreq8_p & v3a67beb;
assign v376fe0c = hbusreq5_p & v376d4cb | !hbusreq5_p & v8455b7;
assign v3743f5b = hbusreq5_p & v3a67971 | !hbusreq5_p & !v3739acd;
assign v3a64dbd = hbusreq1_p & v3768095 | !hbusreq1_p & !v3752648;
assign v377a876 = hbusreq6_p & v3a6dcf0 | !hbusreq6_p & !v372df2a;
assign v374373c = hlock8 & v3a7100a | !hlock8 & v375f985;
assign v3735ee1 = hbusreq7_p & v377f829 | !hbusreq7_p & !v3735cb2;
assign v37393ed = hlock0 & v3a5fc82 | !hlock0 & v37333bb;
assign v372ef36 = hmaster2_p & v3a704cc | !hmaster2_p & v3752dd0;
assign v3a70d0f = hbusreq4 & v375f6ef | !hbusreq4 & v377e8da;
assign v3748472 = jx0_p & v377b5f4 | !jx0_p & v3770b24;
assign v3a6e39a = hmaster0_p & v374a277 | !hmaster0_p & v3737721;
assign v3a6fd1b = hmaster0_p & v8455bf | !hmaster0_p & v374d4ae;
assign v3766e29 = hgrant6_p & v3764276 | !hgrant6_p & v37565a0;
assign v3807474 = hmaster0_p & v372ad34 | !hmaster0_p & v3746ea0;
assign v372b1ed = hlock6_p & v375adaa | !hlock6_p & v2ff8e00;
assign v3770f96 = hgrant4_p & v3a7133d | !hgrant4_p & v3a569a9;
assign v3a571de = hbusreq5_p & v37505a2 | !hbusreq5_p & v3772dd2;
assign v372e213 = hmaster2_p & v3a66d94 | !hmaster2_p & v3a71377;
assign v3a6cae3 = hbusreq5_p & v3730d64 | !hbusreq5_p & v3a58c07;
assign v3a6f617 = hbusreq5_p & v376c248 | !hbusreq5_p & v3a68d0e;
assign v373e654 = hbusreq2 & v3a6ffca | !hbusreq2 & v8455ab;
assign v373ad69 = hbusreq5_p & v8455ab | !hbusreq5_p & v376a6f1;
assign v374a8df = hgrant2_p & v3768b99 | !hgrant2_p & !v37493b9;
assign v3771646 = hbusreq5_p & v3a6fd19 | !hbusreq5_p & v3a610da;
assign da0ed3 = hbusreq8 & v374f768 | !hbusreq8 & !v3a6f330;
assign v3741dac = hlock6 & v3a70125 | !hlock6 & v376c351;
assign v3a5a162 = hbusreq5_p & v3a638aa | !hbusreq5_p & v3a570ee;
assign v3a712e3 = hgrant3_p & v3725b4f | !hgrant3_p & !v3731b11;
assign v3a70373 = hbusreq4 & v375cbe3 | !hbusreq4 & v8455ab;
assign v372840a = hmaster2_p & v3a6ca1f | !hmaster2_p & v3a7044d;
assign v3741e2a = hgrant2_p & v3753f17 | !hgrant2_p & v3a53f45;
assign v376c203 = hlock0 & v3a6fba6 | !hlock0 & v3739391;
assign v3a5ee12 = hgrant2_p & v8455b9 | !hgrant2_p & v37655ac;
assign v37696c4 = hmaster2_p & v375607f | !hmaster2_p & v37745c3;
assign v37286e9 = hgrant4_p & v3765305 | !hgrant4_p & v3a6ff29;
assign v372bf72 = hbusreq7_p & v372d732 | !hbusreq7_p & v3738bdf;
assign v377a653 = hmaster1_p & v3761333 | !hmaster1_p & v3728d9c;
assign v3a705fb = hbusreq6_p & v372f475 | !hbusreq6_p & v3741dab;
assign v3a64b57 = hmaster0_p & v374729b | !hmaster0_p & v3a5c3d7;
assign v376ea80 = hgrant5_p & v8455ab | !hgrant5_p & v2ff9229;
assign v374326f = hbusreq5 & v375e94c | !hbusreq5 & v3a7130e;
assign v3762396 = hgrant5_p & v373ad69 | !hgrant5_p & v3a5ea57;
assign v3732926 = hmaster1_p & v375795d | !hmaster1_p & v374b36f;
assign hgrant2 = !v2aca396;
assign v39eb4a5 = hmaster0_p & v3a70d99 | !hmaster0_p & v373a8b4;
assign v373eef9 = hmaster1_p & v3a6fb85 | !hmaster1_p & v8455dd;
assign v37585a0 = hbusreq1 & v35b7808 | !hbusreq1 & v3a67983;
assign v3a6b4db = hlock7_p & v3733a0e | !hlock7_p & v3a6869f;
assign v3a5ae9f = hmaster1_p & v374e34f | !hmaster1_p & v372c9eb;
assign v3734f9f = hbusreq1 & v3a70131 | !hbusreq1 & !v8455ab;
assign v376589f = hmaster2_p & v3a5690e | !hmaster2_p & v3750a9c;
assign v375fbae = hmaster2_p & v3753418 | !hmaster2_p & v375af43;
assign v3a6422d = hbusreq0 & v3769cc2 | !hbusreq0 & !v8455ab;
assign v373a3b9 = hmaster2_p & v3a700c7 | !hmaster2_p & v3a5a01b;
assign v374c523 = hbusreq2_p & a875ea | !hbusreq2_p & v3808d2e;
assign v3a563c1 = hbusreq5_p & v374edd8 | !hbusreq5_p & v3807601;
assign v3722968 = hmaster1_p & v37447b9 | !hmaster1_p & v37229e6;
assign v3a5cb68 = hbusreq3 & v3809093 | !hbusreq3 & v376bade;
assign v3a5aad8 = hmaster0_p & v3736d47 | !hmaster0_p & v3754caa;
assign v3a5996e = hbusreq0_p & v3754ec1 | !hbusreq0_p & !v3a5e817;
assign v372586f = hbusreq8 & v3764461 | !hbusreq8 & v3754295;
assign v3a5c317 = jx1_p & v3737edc | !jx1_p & v3771dd8;
assign v3a6908b = hgrant4_p & v3744934 | !hgrant4_p & v3a5787a;
assign v3a5c645 = hmaster2_p & v3806c9a | !hmaster2_p & v374b8fa;
assign v3a5fd6a = hlock4_p & v3a6c60e | !hlock4_p & v3760f4e;
assign v373ec60 = hbusreq5_p & v3770f48 | !hbusreq5_p & v3a7122f;
assign v37711ec = hbusreq5 & v3a69758 | !hbusreq5 & v373790d;
assign v3a5727d = hgrant4_p & v3a63eaf | !hgrant4_p & v372936a;
assign v372d828 = hbusreq3_p & v3729b63 | !hbusreq3_p & !v8455ab;
assign v2ff8e00 = hgrant2_p & v8455ab | !hgrant2_p & v3770651;
assign v1e3746e = hburst0 & v3a299c1 | !hburst0 & v3772e90;
assign v3a715fd = stateA1_p & v8455e1 | !stateA1_p & !v376a35c;
assign v373ba84 = hbusreq7 & v3a6856a | !hbusreq7 & v374170e;
assign v3a7114b = hmaster2_p & v37248fd | !hmaster2_p & v3726c20;
assign v375b68b = hbusreq6 & v372dccf | !hbusreq6 & v3a69487;
assign v3a7157d = hmaster0_p & v377a121 | !hmaster0_p & v3a6fe4d;
assign v375912e = jx0_p & v3a70533 | !jx0_p & v3a6a893;
assign v3a6054b = hmaster1_p & v372ebc8 | !hmaster1_p & v8455ab;
assign v3a5f000 = hmaster2_p & v3770b26 | !hmaster2_p & v373195f;
assign v374b1a4 = hmaster2_p & c9bec3 | !hmaster2_p & v3a650bb;
assign v3739077 = hbusreq8_p & v373c590 | !hbusreq8_p & v375e3fd;
assign v1e37b52 = hgrant7_p & v37500d0 | !hgrant7_p & v3a6feb5;
assign v3a62f14 = hmaster1_p & v3a555ae | !hmaster1_p & v8455ab;
assign v3a66534 = hgrant4_p & v3a67cff | !hgrant4_p & v374165f;
assign v3a68b49 = hbusreq2_p & v373be25 | !hbusreq2_p & !v372935c;
assign v3a70b15 = hmaster0_p & v8455ab | !hmaster0_p & v3747a7b;
assign v3a661f1 = hmaster2_p & v3a6ffb6 | !hmaster2_p & v372c3d4;
assign v3745828 = hbusreq4_p & v3747302 | !hbusreq4_p & v3733b77;
assign v3a7094f = hmaster2_p & v3a6d569 | !hmaster2_p & v3a70fa6;
assign v3a711fb = hbusreq3 & v37774c7 | !hbusreq3 & v3a70c74;
assign v3a6acd3 = hbusreq5_p & v377e0c6 | !hbusreq5_p & v8455ab;
assign v3a6a939 = hmastlock_p & v3a70a83 | !hmastlock_p & v8455ab;
assign v372750b = hmaster0_p & v376111d | !hmaster0_p & v375dc5f;
assign v372bfd3 = hgrant6_p & v374530a | !hgrant6_p & !v373502e;
assign v377f342 = hbusreq3_p & v3726cf7 | !hbusreq3_p & !v3a658bf;
assign v377550d = hbusreq6 & v3a6ff2d | !hbusreq6 & v3a58102;
assign v375139a = hmaster2_p & v8455ab | !hmaster2_p & !v3a714aa;
assign v3a6b423 = hlock2_p & v8455ab | !hlock2_p & !v3753f1a;
assign v372b50b = hmaster0_p & v377e298 | !hmaster0_p & v3764a7d;
assign v3a661b5 = hbusreq6_p & v372cd3f | !hbusreq6_p & v8455ab;
assign v3729a07 = hbusreq8 & v3a68c27 | !hbusreq8 & v374a4cc;
assign v376beca = hbusreq7_p & v3a70d9e | !hbusreq7_p & v3764f39;
assign v3732f4d = hbusreq7 & v3a70e68 | !hbusreq7 & v373d40c;
assign v3751fbe = hbusreq7 & v3772b81 | !hbusreq7 & v3734868;
assign v376300a = hgrant4_p & v376a6f1 | !hgrant4_p & v37577b7;
assign v376067f = hbusreq0 & v3760854 | !hbusreq0 & v3a6f145;
assign v3a6fbad = hmaster2_p & v3a70209 | !hmaster2_p & !v373325f;
assign v373f8b1 = hgrant6_p & v3727cd0 | !hgrant6_p & v376c635;
assign v3723d16 = hmaster3_p & v3a6f900 | !hmaster3_p & !v3747d69;
assign v3a5a260 = hgrant5_p & v8455ab | !hgrant5_p & v3727e10;
assign v3378fc3 = hlock5_p & v3736ded | !hlock5_p & v8455bb;
assign v372993f = hbusreq5_p & v3a71470 | !hbusreq5_p & v376bc6b;
assign v3a6f02c = hburst0 & v3a6f8df | !hburst0 & v376acf0;
assign v3a6c6aa = hlock0_p & v373905f | !hlock0_p & v375168a;
assign v87762a = hmaster1_p & v377c7c0 | !hmaster1_p & v37263c1;
assign v3778b51 = hlock6_p & v372abd8 | !hlock6_p & v35772a6;
assign v372ee06 = hbusreq0 & v3a66606 | !hbusreq0 & v8455ab;
assign v3a702a2 = hbusreq4_p & v3747302 | !hbusreq4_p & v37496fa;
assign v3a65e9d = hmaster0_p & v376d6ef | !hmaster0_p & v3a6fd53;
assign v3a6f42c = hgrant3_p & v37331e7 | !hgrant3_p & v376faad;
assign v37735cb = hbusreq6_p & v377c003 | !hbusreq6_p & db3b98;
assign v372600f = hgrant3_p & v8455ab | !hgrant3_p & v375a28a;
assign v3735ba1 = hbusreq7 & v3a71556 | !hbusreq7 & v3a60276;
assign v3a6f968 = hlock6_p & v372ab21 | !hlock6_p & v8455b7;
assign v3a5fc33 = hmaster0_p & v373040b | !hmaster0_p & v35b774b;
assign v373666f = hmaster0_p & v372567a | !hmaster0_p & v23fe28c;
assign v3755312 = hbusreq0 & v3722e5e | !hbusreq0 & v8455ab;
assign v3a6f709 = hlock6 & v3a7144a | !hlock6 & v3770e35;
assign v3a70144 = hbusreq5_p & v3774628 | !hbusreq5_p & !v375f44a;
assign v3a70960 = hlock4 & v3a6eb1b | !hlock4 & v3769112;
assign v3a6a489 = hbusreq6 & v37235ee | !hbusreq6 & v8455ab;
assign v3a6feb5 = jx1_p & v38064a1 | !jx1_p & v3a7017f;
assign v376bd2a = start_p & v3726abd | !start_p & v8455ab;
assign v3a6f0d9 = hbusreq6 & v3a6dc08 | !hbusreq6 & v372d0ad;
assign v3a700ae = hbusreq6_p & v375641f | !hbusreq6_p & !v3a6b0c7;
assign v377eda6 = hbusreq4_p & v3a70554 | !hbusreq4_p & v3768b3d;
assign v3a70994 = hmaster2_p & v37782c9 | !hmaster2_p & v37416c6;
assign v3725ca4 = hlock7_p & v3a70fd9 | !hlock7_p & v3a66fb0;
assign v35b7734 = hbusreq8 & v377a812 | !hbusreq8 & !v3779f92;
assign b5a5ab = hmaster1_p & v377d0e6 | !hmaster1_p & !v37702c5;
assign v372757f = hmaster2_p & v37771e3 | !hmaster2_p & v3764978;
assign v3723089 = hbusreq7 & v3a6fa70 | !hbusreq7 & v3a70bf0;
assign v37546a4 = hbusreq7_p & v376c17d | !hbusreq7_p & v3776d32;
assign v374f691 = hmaster0_p & v377a51b | !hmaster0_p & v3753097;
assign v372628c = hgrant4_p & v372abd8 | !hgrant4_p & v3a6f31c;
assign v3a5f265 = hlock0_p & v3747302 | !hlock0_p & v3726c36;
assign v3736901 = hbusreq2 & v3757d20 | !hbusreq2 & v3a70a7f;
assign v376ba56 = hmaster0_p & v3a6f406 | !hmaster0_p & v3a6a1af;
assign v377cda9 = hbusreq5 & c81b97 | !hbusreq5 & v375b0ad;
assign v3a6eefa = hlock8_p & v3a62009 | !hlock8_p & v3a70892;
assign v3777142 = hlock5 & v374a806 | !hlock5 & v3a6f2d8;
assign v37550ac = hlock8_p & v3a618f6 | !hlock8_p & !v8455ab;
assign v3a70eb0 = hbusreq5_p & v3774b16 | !hbusreq5_p & v39eb520;
assign v3744b11 = hbusreq7 & v3725bb3 | !hbusreq7 & v376e8e3;
assign v373fecd = hmastlock_p & v372cf62 | !hmastlock_p & v8455ab;
assign v374febd = hbusreq0 & v3748d1f | !hbusreq0 & v375d6e8;
assign v3726bb7 = jx0_p & v3775ec8 | !jx0_p & v3a6df51;
assign v375dcac = hgrant4_p & v376983e | !hgrant4_p & v3753eb3;
assign v3a70739 = hmaster1_p & v3a6f467 | !hmaster1_p & v8455ab;
assign v3a70fce = hmaster0_p & v3a6f6a2 | !hmaster0_p & v3756d28;
assign v3a5d5d3 = hbusreq2 & v8455b0 | !hbusreq2 & v8455ab;
assign v3748e6a = hbusreq7 & v372f1a8 | !hbusreq7 & v3a6ec01;
assign v3a7162b = hbusreq7_p & v373a77b | !hbusreq7_p & v3a6f925;
assign v3757993 = hmaster2_p & v3744835 | !hmaster2_p & v3a6eb2f;
assign v3a698d8 = hbusreq8 & v3757f07 | !hbusreq8 & v3736e7c;
assign v3a713df = hbusreq6_p & aa5556 | !hbusreq6_p & v8455ab;
assign v3749658 = hlock5_p & v377c174 | !hlock5_p & v8455ab;
assign v3765583 = hgrant5_p & v3a70769 | !hgrant5_p & v37270b5;
assign v374a97f = hbusreq3_p & v3a640c5 | !hbusreq3_p & v3a5cd20;
assign v3766d29 = hmaster2_p & v3a6f998 | !hmaster2_p & v3730986;
assign v3a7137c = hbusreq4_p & v3a712af | !hbusreq4_p & v373fb71;
assign v373e6d8 = jx0_p & v3751983 | !jx0_p & v3a6f816;
assign v3731e3a = hbusreq6_p & v3a61eea | !hbusreq6_p & v8455ab;
assign v3a59085 = hbusreq5 & v3727c07 | !hbusreq5 & v3775687;
assign v3738cab = hgrant4_p & v8455ab | !hgrant4_p & v37456d2;
assign v3767638 = hbusreq5 & v3a70fd5 | !hbusreq5 & !v3745bbe;
assign v3a59c1d = hbusreq5_p & v3754392 | !hbusreq5_p & v8455ab;
assign v37748b7 = hbusreq4 & v3a5468d | !hbusreq4 & v8455ab;
assign v35b71fc = hmaster1_p & v3a635ea | !hmaster1_p & v3752616;
assign v3758166 = hbusreq2_p & v3759032 | !hbusreq2_p & v3733e9e;
assign v3759d78 = hbusreq6 & v3a6f4bc | !hbusreq6 & v372781d;
assign cc8eeb = hbusreq7_p & v372706f | !hbusreq7_p & v35b7070;
assign v377c8c8 = hmaster3_p & v8455ab | !hmaster3_p & v374e18a;
assign v37793d4 = hbusreq5_p & v3727342 | !hbusreq5_p & !v8455ab;
assign v3a5f0b2 = hbusreq3_p & v375fcfb | !hbusreq3_p & v8455ab;
assign v374ac8c = hmaster2_p & v372cac6 | !hmaster2_p & v373a3fa;
assign v3a71247 = hbusreq0 & v3730b63 | !hbusreq0 & v3a5e90f;
assign v37293e0 = hmaster2_p & v37793e4 | !hmaster2_p & v374aec2;
assign v3a6ebb8 = hbusreq4_p & v377349f | !hbusreq4_p & v3749a32;
assign v3a6870f = hmaster0_p & v375bb10 | !hmaster0_p & v372cdd5;
assign v3a5857e = jx0_p & v37632c6 | !jx0_p & v8455ab;
assign v377ef6e = hbusreq4 & v3739d88 | !hbusreq4 & v3a5a807;
assign v3729214 = hbusreq6_p & v3a6f09c | !hbusreq6_p & !v3a704c2;
assign v3806a7b = hbusreq5_p & v3a708b5 | !hbusreq5_p & !v3a6dfb2;
assign v3a6e5e1 = hbusreq4 & v375c263 | !hbusreq4 & v8455ab;
assign v3a7116e = hbusreq2_p & v3742905 | !hbusreq2_p & v3a69946;
assign v380a2f5 = hbusreq6 & v376d1e2 | !hbusreq6 & v3a69487;
assign v3a68467 = hgrant5_p & v8455ab | !hgrant5_p & v3a7017b;
assign v3a5a6fb = hmaster2_p & v376a6f1 | !hmaster2_p & !v374bbc7;
assign v3762d06 = hmaster2_p & v376e3fb | !hmaster2_p & v3733343;
assign v3a6edfb = hbusreq5_p & v3740fc3 | !hbusreq5_p & v8455ab;
assign v3778a5a = hmaster2_p & v3a70cc3 | !hmaster2_p & v377928c;
assign v37591ae = hgrant6_p & v377c147 | !hgrant6_p & v3724887;
assign v37452a4 = hmaster2_p & v373a4e4 | !hmaster2_p & v376e89b;
assign v3a5a211 = hbusreq6_p & v373a29c | !hbusreq6_p & v3a5cf22;
assign v3a6f48c = hgrant4_p & v3a653e4 | !hgrant4_p & !v3763ce3;
assign v3a6443d = hgrant6_p & v3a71389 | !hgrant6_p & v3737416;
assign v3a5be72 = hlock0_p & v3a70cdb | !hlock0_p & v8455b0;
assign v3753b5e = hbusreq2 & v3770ae6 | !hbusreq2 & v38072fd;
assign v37314cc = hbusreq4 & v376111d | !hbusreq4 & v8455ab;
assign v3a707a0 = hlock6 & v375a80c | !hlock6 & v377bb66;
assign v3761026 = hmaster1_p & v374457a | !hmaster1_p & v3774359;
assign v3a7026a = hmaster2_p & v375b42e | !hmaster2_p & v3759b71;
assign v3a71194 = hmaster0_p & v3808d48 | !hmaster0_p & v3a6cf7f;
assign bc9e23 = hbusreq0_p & v372dadb | !hbusreq0_p & v3a6123e;
assign v377a87d = hmaster1_p & v39ea76e | !hmaster1_p & v3a6ff27;
assign v3808d7d = hmaster0_p & v8455ab | !hmaster0_p & v3a5b404;
assign v375248f = hbusreq4_p & v8455ab | !hbusreq4_p & v37604b3;
assign v3a5f642 = hlock4_p & v373a841 | !hlock4_p & v3765e46;
assign v375058a = hbusreq5_p & v3736260 | !hbusreq5_p & v8455ab;
assign v374cd15 = hmaster1_p & v3751d33 | !hmaster1_p & !v3779613;
assign v374203a = hbusreq2_p & v373e782 | !hbusreq2_p & !v3725f77;
assign v3750519 = hbusreq5_p & v3a6f047 | !hbusreq5_p & !v8455ab;
assign v372818d = hbusreq4 & v3732f03 | !hbusreq4 & v8455ab;
assign v374e304 = hmaster3_p & v3779910 | !hmaster3_p & v3a6f47d;
assign v3a6f9ce = hmaster0_p & v3a6f9ed | !hmaster0_p & v3a7026a;
assign v375d445 = hlock4 & v38079dc | !hlock4 & v3a5966b;
assign v376a2ea = hlock0_p & v377989c | !hlock0_p & v3a6ffca;
assign v3a70922 = hmaster0_p & v3a70696 | !hmaster0_p & v3741320;
assign v372b388 = hgrant6_p & v37781ac | !hgrant6_p & v37643eb;
assign v374ad24 = hbusreq6_p & v375bdd4 | !hbusreq6_p & v8455e1;
assign v3a70c36 = hbusreq3_p & v372c3d4 | !hbusreq3_p & !v3a5ef5c;
assign v3752281 = hmaster2_p & v3a6ef95 | !hmaster2_p & v3a6848c;
assign v372e749 = hbusreq5_p & v375fdb5 | !hbusreq5_p & v37551ac;
assign v3745c8f = hgrant3_p & v8455ab | !hgrant3_p & v374a681;
assign v372adaa = hbusreq6_p & v3a6650e | !hbusreq6_p & !v8455ab;
assign v377e13b = hbusreq6_p & v3a707f6 | !hbusreq6_p & v377671e;
assign v3a6f314 = hlock3_p & v374b0c1 | !hlock3_p & v37720e5;
assign v3a7063e = hbusreq0 & v3734e69 | !hbusreq0 & v377a6dc;
assign v3a70647 = hmaster0_p & v374502e | !hmaster0_p & v376652f;
assign v3a5e3d1 = hbusreq7 & v3771a24 | !hbusreq7 & v3749ca6;
assign v3757746 = hgrant0_p & v3753edb | !hgrant0_p & v376e364;
assign v37615d0 = hbusreq5_p & v3775533 | !hbusreq5_p & v3752df5;
assign v3747084 = hbusreq5 & v3a6fd98 | !hbusreq5 & v2925d03;
assign v3a6dc32 = hlock3_p & v375b8b2 | !hlock3_p & v37406d2;
assign v3736539 = hmaster2_p & v3a70385 | !hmaster2_p & !v8455ab;
assign v3751022 = hmaster0_p & v3a6672b | !hmaster0_p & c536d5;
assign v3a6a116 = hgrant2_p & v372b17b | !hgrant2_p & v375f71d;
assign v375179a = hlock4_p & v3745131 | !hlock4_p & v372c706;
assign v3722d85 = hmaster1_p & v3a6f51e | !hmaster1_p & v3738826;
assign v3771622 = hlock8 & v3a6a76d | !hlock8 & v3758892;
assign v3a7026d = hbusreq5 & v3766acb | !hbusreq5 & v3772e85;
assign v376498a = hgrant1_p & v3a6e591 | !hgrant1_p & v3a6f436;
assign v3a67967 = hbusreq2_p & v372c502 | !hbusreq2_p & v8455ab;
assign v375624b = hbusreq4_p & v3a635ea | !hbusreq4_p & v372e8d8;
assign v3a6a1b4 = hbusreq0 & v3807a8d | !hbusreq0 & v373e858;
assign v3a59d07 = hbusreq0 & v375d1a6 | !hbusreq0 & v37513b7;
assign v3a71088 = hbusreq2_p & v37765e1 | !hbusreq2_p & v373c480;
assign v377613d = hgrant3_p & v3a6cdbc | !hgrant3_p & v37598c6;
assign v3a70d60 = hlock8_p & v3a68c63 | !hlock8_p & v3a6c127;
assign v3a67f0c = hmaster0_p & v8455ab | !hmaster0_p & v3747a3f;
assign v37544ab = hmaster3_p & v3779879 | !hmaster3_p & !v8455ab;
assign v374c163 = hbusreq2_p & v3763a20 | !hbusreq2_p & v377cd7a;
assign v3736e1d = hbusreq1_p & v3727507 | !hbusreq1_p & v3748797;
assign v3725be9 = hbusreq8 & v3a6f4dd | !hbusreq8 & cd5e35;
assign v3a5a220 = hburst0 & v3a6ffa9 | !hburst0 & v377ac6f;
assign v374797c = hmaster2_p & v3a635ea | !hmaster2_p & v377b946;
assign v375f847 = hmaster2_p & v3a6b8aa | !hmaster2_p & v3751acf;
assign v3a705f7 = hlock0_p & v3a635ea | !hlock0_p & v3775e66;
assign v3a58dfc = hmaster0_p & v3a6f7dd | !hmaster0_p & v3a6f957;
assign v3a6f8d5 = hbusreq4 & v3773575 | !hbusreq4 & v373b78b;
assign v372e4e3 = hbusreq4_p & v3751e80 | !hbusreq4_p & v3755420;
assign v375515c = hbusreq7_p & v3725e12 | !hbusreq7_p & v8455ab;
assign v3739c68 = hgrant4_p & v8455ab | !hgrant4_p & v3743d8b;
assign v3a69c05 = hlock6_p & v3a56642 | !hlock6_p & v3730ffe;
assign v373e962 = hbusreq2 & v3742d54 | !hbusreq2 & v3a6fdef;
assign v3768d29 = hbusreq6 & v3a56608 | !hbusreq6 & v3748797;
assign v3a6ff37 = hgrant6_p & v3730926 | !hgrant6_p & v37c038c;
assign v376ba96 = jx0_p & v3760237 | !jx0_p & v3a54242;
assign v374c3bf = hgrant5_p & v3a6eb8c | !hgrant5_p & v3758291;
assign v3750cfa = hbusreq5_p & v3a5c4e1 | !hbusreq5_p & v8455ab;
assign v377a617 = hbusreq4_p & v375641f | !hbusreq4_p & !v3a6b0c7;
assign v373763f = hmaster1_p & v373c15d | !hmaster1_p & v374b747;
assign v3a711d1 = hbusreq5 & v23fda7e | !hbusreq5 & v8455ab;
assign v37707b6 = hmaster2_p & v3727f14 | !hmaster2_p & v8455ab;
assign v3a70430 = hbusreq8_p & v3a6ebd8 | !hbusreq8_p & v376a74a;
assign v374aa4f = hmaster1_p & v375b046 | !hmaster1_p & !v372f9b4;
assign v3739ec9 = hmaster2_p & v374571d | !hmaster2_p & v3a5f40e;
assign v3a62245 = hmaster2_p & v3a635ea | !hmaster2_p & v9b03cc;
assign v3722dfe = hmaster2_p & v3735d9c | !hmaster2_p & v3a54b63;
assign v3a5b0dd = hbusreq0 & v3737028 | !hbusreq0 & v8455ab;
assign v2ff87c6 = hmaster0_p & v3a637dc | !hmaster0_p & v3a68b0a;
assign v360d1cb = hbusreq3_p & v924b19 | !hbusreq3_p & v3a60132;
assign v374401a = hlock2 & v3a712da | !hlock2 & v3752831;
assign v374b867 = hmaster1_p & v374f307 | !hmaster1_p & v3736d0d;
assign v8cb684 = hbusreq4 & v3723ace | !hbusreq4 & v8455b0;
assign v375d887 = hbusreq4_p & v37422b5 | !hbusreq4_p & !v8455ab;
assign v37707eb = hgrant0_p & v373cf42 | !hgrant0_p & v37775c4;
assign v3759abe = hbusreq2_p & v8455ab | !hbusreq2_p & v373125c;
assign v375ab35 = stateG3_2_p & v8455ab | !stateG3_2_p & v3731e3c;
assign v3a6adf2 = hmaster1_p & v375c7cf | !hmaster1_p & v376ab39;
assign v3a6fbb8 = jx3_p & v3743172 | !jx3_p & v3a6f233;
assign v3a643d7 = hbusreq6 & v3a714b3 | !hbusreq6 & v377728d;
assign v3745bee = hmaster0_p & v3a6fa35 | !hmaster0_p & v3a5f76b;
assign v3a6a045 = hmaster0_p & v3a6c4b3 | !hmaster0_p & v3729004;
assign v3a29810 = hbusreq0 & v3a702e1 | !hbusreq0 & v3a7062f;
assign v3a5fa22 = hgrant4_p & v3776cce | !hgrant4_p & v8455ab;
assign v376c630 = hbusreq6_p & v377fb00 | !hbusreq6_p & v3378f4c;
assign v3753976 = hmaster0_p & v3a703fa | !hmaster0_p & !v3a703be;
assign v3a6f5cb = hmaster0_p & v3a6dc83 | !hmaster0_p & v375bfe5;
assign v3756203 = hbusreq4_p & v3a5f8d0 | !hbusreq4_p & v3775303;
assign v3a57913 = hmaster1_p & v3a57db6 | !hmaster1_p & v8455ab;
assign v3a7152b = hbusreq5_p & v374067c | !hbusreq5_p & v8455ab;
assign v376f5d9 = hmaster2_p & v3766bc8 | !hmaster2_p & !v3a627cc;
assign v3741b92 = hbusreq4_p & v3a6fc8f | !hbusreq4_p & !v3a5bf04;
assign v3728d1d = hmaster0_p & v3763f95 | !hmaster0_p & v3a71560;
assign v3772bda = hbusreq5 & v3a7140f | !hbusreq5 & v37494c3;
assign v3a6f820 = hgrant5_p & v8455c6 | !hgrant5_p & be54b2;
assign v3a5be93 = hbusreq6_p & v374535e | !hbusreq6_p & v8455ab;
assign v3760b3d = hbusreq2_p & v8455ab | !hbusreq2_p & v3731300;
assign v3747527 = hgrant3_p & v8455ab | !hgrant3_p & v376f3c8;
assign v3a7062f = hbusreq4 & v3a702e1 | !hbusreq4 & v3a70088;
assign v374f617 = hbusreq2_p & v3a557b1 | !hbusreq2_p & v3744590;
assign v3a5af26 = hmaster0_p & v372f309 | !hmaster0_p & v3a7155b;
assign v377d7e1 = hgrant3_p & v3743f11 | !hgrant3_p & v8455ab;
assign v377ce91 = hbusreq8_p & v374fb2f | !hbusreq8_p & v37519e2;
assign v3762b55 = hlock6 & v375a41b | !hlock6 & v37642a0;
assign v374ec22 = hlock0_p & v3a6ee22 | !hlock0_p & v8455ab;
assign v3a70586 = hbusreq5 & v377a0d8 | !hbusreq5 & v360bc74;
assign v3778a4f = jx0_p & v3a6fb49 | !jx0_p & v3724579;
assign v360d01e = hgrant5_p & v3a6f650 | !hgrant5_p & v3739e05;
assign v37602cf = hbusreq6_p & v95151c | !hbusreq6_p & v375d6ba;
assign a5679d = hbusreq1 & v376dbdf | !hbusreq1 & v8455ab;
assign v3a60132 = hbusreq3 & v8455b0 | !hbusreq3 & v8455ab;
assign v377a511 = hgrant2_p & v37234e0 | !hgrant2_p & !v374c425;
assign v3737f16 = jx0_p & v3761781 | !jx0_p & v3730c49;
assign v3a64112 = hbusreq6 & v3a70cc3 | !hbusreq6 & v8455ab;
assign v377e547 = hbusreq8 & v3748299 | !hbusreq8 & v3730c0b;
assign v374d0ad = jx0_p & v37414be | !jx0_p & v3a6f665;
assign v3a5ebc2 = hbusreq5_p & v374c6b8 | !hbusreq5_p & v373e873;
assign v37313e4 = hmaster0_p & v3a66aa4 | !hmaster0_p & v373fe1f;
assign v375aeca = hgrant2_p & v8455ab | !hgrant2_p & v3746d07;
assign v375fae9 = hmaster1_p & v8455ab | !hmaster1_p & v375df5e;
assign v3a70f52 = hbusreq8 & v3a5a8e6 | !hbusreq8 & v8455ab;
assign v3730e43 = hmaster2_p & v3a5fc34 | !hmaster2_p & !v3755252;
assign v374db73 = hmaster0_p & v3a6dc83 | !hmaster0_p & v3a6c9aa;
assign v3750113 = hbusreq5_p & v3a70ee6 | !hbusreq5_p & v3a6f237;
assign v3738e45 = hbusreq8_p & v37385fc | !hbusreq8_p & v3740923;
assign v3a6e8a6 = hbusreq4_p & v37706a7 | !hbusreq4_p & v3a6bf89;
assign v372a1a9 = hmaster1_p & v3764d40 | !hmaster1_p & !v373e055;
assign v3a70295 = hbusreq0_p & v37397c3 | !hbusreq0_p & v37341bc;
assign v3a5e239 = hbusreq0 & v3735708 | !hbusreq0 & v37483c5;
assign v376ca86 = hgrant6_p & v3a635ea | !hgrant6_p & v3a6fc0b;
assign v372a201 = stateG10_1_p & v8455ab | !stateG10_1_p & v3a6bdd7;
assign v373f704 = hgrant2_p & v3a71121 | !hgrant2_p & v3777c39;
assign v3a6fa3f = hbusreq0 & v3a715ab | !hbusreq0 & v37473a3;
assign v3736ee0 = hgrant4_p & v3a6b7e9 | !hgrant4_p & v3761433;
assign v3763550 = hmaster2_p & v373a7a5 | !hmaster2_p & v375b880;
assign v3a7126c = hlock6 & v37565be | !hlock6 & v3768130;
assign v3762c7f = hbusreq5_p & v89fdcf | !hbusreq5_p & v372efcb;
assign v3a6a680 = hbusreq4_p & v3a66381 | !hbusreq4_p & v3774ee5;
assign v3724023 = hmaster0_p & d893c7 | !hmaster0_p & v8455ab;
assign v3753883 = hmaster2_p & v2ff8cfd | !hmaster2_p & v3754b35;
assign v37712fa = hbusreq5_p & v3809505 | !hbusreq5_p & v8455cb;
assign v37244f1 = hmaster1_p & v3a55542 | !hmaster1_p & v3762c7f;
assign v37674d1 = hbusreq5 & v37586bb | !hbusreq5 & v3769215;
assign v38090f6 = hgrant2_p & v3a710a2 | !hgrant2_p & v376aeae;
assign v3a6b8d8 = hgrant6_p & v8455ab | !hgrant6_p & v372a902;
assign v3a7081b = hbusreq3 & v3757746 | !hbusreq3 & v8455ab;
assign v373c96e = hbusreq6 & v373aaa8 | !hbusreq6 & v8455ab;
assign v3766a8d = hbusreq4_p & v3763a20 | !hbusreq4_p & v3a55bd0;
assign v3a6f3fa = hmaster0_p & v372f309 | !hmaster0_p & v377d8c8;
assign v3a6de33 = locked_p & v377e976 | !locked_p & v37563eb;
assign v374c107 = hgrant4_p & v3741b92 | !hgrant4_p & !v377d821;
assign v3a6f23a = hbusreq4_p & ae317f | !hbusreq4_p & v3768c3e;
assign v3732a41 = stateA1_p & v8455e1 | !stateA1_p & !v3a6feed;
assign v3a6f3d6 = hready_p & v3a627a8 | !hready_p & v3a70680;
assign bbcc5e = hgrant4_p & v3a6eb47 | !hgrant4_p & v3a6b53f;
assign v372618d = hgrant0_p & v8455ab | !hgrant0_p & v37241cc;
assign v3738373 = hlock7_p & v3a70956 | !hlock7_p & v3736dfe;
assign v3770a77 = hgrant2_p & v3a702b4 | !hgrant2_p & cd3a92;
assign v3a590fb = hbusreq2 & v3377af7 | !hbusreq2 & v377c6b3;
assign v3767b66 = hgrant6_p & v8455ca | !hgrant6_p & v376975e;
assign v3737ca3 = hbusreq2 & v3760740 | !hbusreq2 & v8455ab;
assign v3a702d8 = hbusreq5 & v3a70380 | !hbusreq5 & v8455ab;
assign v3739e7a = hlock4 & v3a6f0a5 | !hlock4 & v3762312;
assign v3a70a87 = hlock6 & v372c944 | !hlock6 & v376c4c5;
assign v3725ba5 = hbusreq5 & v373497f | !hbusreq5 & v3a6eed9;
assign v377c38c = hbusreq2_p & v3a5f8d0 | !hbusreq2_p & v3775303;
assign v39ebb8a = hbusreq5_p & v37384a9 | !hbusreq5_p & v3a70b3b;
assign v3723a30 = hmaster0_p & v3757568 | !hmaster0_p & v3a6a36d;
assign v2925d2c = hgrant6_p & v8455ab | !hgrant6_p & v3807026;
assign v3776ce0 = hbusreq1_p & v3806507 | !hbusreq1_p & v3a63621;
assign v3744796 = hgrant3_p & v377052f | !hgrant3_p & v8455ab;
assign v3742851 = hmaster2_p & v3760eeb | !hmaster2_p & v3768ecc;
assign v37449b3 = hbusreq4_p & v37316bb | !hbusreq4_p & v372ba0f;
assign v376cddf = hmaster1_p & v37667f8 | !hmaster1_p & v3757272;
assign v3725fe5 = hgrant2_p & v8455ba | !hgrant2_p & v3a6ff7c;
assign v37725c6 = hlock5 & v3a63f9a | !hlock5 & v375e5ed;
assign v3a70315 = hgrant6_p & v8455ab | !hgrant6_p & v3736a9a;
assign v3a708b5 = hlock5_p & v3779060 | !hlock5_p & !v3a6fbe8;
assign v3a5b037 = hbusreq3_p & v3a6cb50 | !hbusreq3_p & v8455ab;
assign v37605ab = hbusreq5_p & v3a602cd | !hbusreq5_p & v3a6e8bc;
assign v373df9c = hbusreq0_p & v372e169 | !hbusreq0_p & v3748797;
assign v3a713c0 = jx0_p & v373fd51 | !jx0_p & v3765298;
assign v37439ad = hlock0_p & v372b24d | !hlock0_p & v375ecc7;
assign v3735fdc = hlock0 & v3a635ea | !hlock0 & v372a79f;
assign v3a70c21 = hgrant8_p & v3745d3f | !hgrant8_p & v3a5fc64;
assign v375e737 = hlock8_p & v375d388 | !hlock8_p & v373d687;
assign v3a68377 = hbusreq5_p & v3755c0e | !hbusreq5_p & !v3779288;
assign v3779e9b = hmaster1_p & v373ea09 | !hmaster1_p & v374e7fa;
assign d23bf8 = hlock4_p & v1e38275 | !hlock4_p & v39a537f;
assign v37346e8 = hlock0 & v3765e79 | !hlock0 & v375ef49;
assign v374a9d0 = hbusreq5_p & v3a64421 | !hbusreq5_p & v3a635ea;
assign v3a5cfed = hbusreq0_p & v3770cd8 | !hbusreq0_p & v376b3b0;
assign v3763f8e = hbusreq5 & v37262ad | !hbusreq5 & v8455ab;
assign v3734914 = hlock5 & v3772bda | !hlock5 & v3a7140f;
assign v375c4ac = hlock4 & v375cdf4 | !hlock4 & v3736c8d;
assign v377e283 = hmaster0_p & v37710d4 | !hmaster0_p & v373cddc;
assign v374f533 = hmaster0_p & v3724e45 | !hmaster0_p & v3741320;
assign fc6f92 = hmaster0_p & v28896b4 | !hmaster0_p & v373d69f;
assign v3a6ff9a = hmaster1_p & v3a61a7f | !hmaster1_p & v375fe83;
assign v37262ec = hgrant5_p & v8455ab | !hgrant5_p & v3a6fc68;
assign v3a6a1fd = hgrant2_p & v3746dd5 | !hgrant2_p & v37705d1;
assign v3747eef = hgrant0_p & v3759032 | !hgrant0_p & v3770cd8;
assign v3764f06 = hmaster0_p & v3740ab8 | !hmaster0_p & !v375f847;
assign v377bc89 = hgrant3_p & v8455e7 | !hgrant3_p & !v35b7160;
assign v3722dba = hbusreq1 & v3724940 | !hbusreq1 & v8455ab;
assign v375c94e = hmaster0_p & v37538af | !hmaster0_p & b0e59c;
assign v372b59f = hmaster1_p & v3747d5a | !hmaster1_p & v377cf71;
assign v374db32 = hgrant6_p & v8455ab | !hgrant6_p & v3a70ec9;
assign v3a578af = hlock5 & v3a7038a | !hlock5 & v3753804;
assign v3758d56 = hgrant4_p & v8455ab | !hgrant4_p & v3a6bf41;
assign v3757169 = hmaster0_p & v8455ab | !hmaster0_p & !v375e624;
assign v3806636 = hmaster0_p & v3a635ea | !hmaster0_p & v372a417;
assign v3a6ebda = hbusreq8_p & v3a620fd | !hbusreq8_p & v3a6ebc6;
assign v374ad67 = hgrant6_p & v3a6f3da | !hgrant6_p & dc6ded;
assign v375d7df = hmaster2_p & d1bf3b | !hmaster2_p & !v373b5f0;
assign v3730fb0 = hbusreq6_p & v3776e85 | !hbusreq6_p & v3378f4c;
assign v3775252 = hlock0 & v374617d | !hlock0 & v373cd41;
assign v3a5f89e = hlock6_p & v35b9d52 | !hlock6_p & v8455ab;
assign v372e959 = hmaster2_p & v3806db0 | !hmaster2_p & v374f501;
assign v3a70af0 = hbusreq5 & v3a70a75 | !hbusreq5 & v3a6d6fb;
assign v372b3dd = hbusreq5_p & v374f8f6 | !hbusreq5_p & !v3768918;
assign v374f26c = hmaster1_p & v3807aa1 | !hmaster1_p & v372ac1d;
assign v3758ff4 = hgrant6_p & v3752304 | !hgrant6_p & v3a5ee3a;
assign v375e7d6 = hbusreq2_p & v373a181 | !hbusreq2_p & v35772a6;
assign v3730a2f = hlock0 & v38073c9 | !hlock0 & v3a7082c;
assign v376cb10 = hmaster1_p & v3a6fa77 | !hmaster1_p & v376e441;
assign v37533c3 = hgrant0_p & v8455ab | !hgrant0_p & v377fabc;
assign v3a6feab = hmaster1_p & v8455ab | !hmaster1_p & v37433d5;
assign v3a6fe44 = hlock6 & v374d9b3 | !hlock6 & v372fd12;
assign v3a70aef = hmaster2_p & v372d727 | !hmaster2_p & v3776ada;
assign v3761dda = hbusreq5 & v376fbe3 | !hbusreq5 & v37366d5;
assign v3a69b91 = hmaster1_p & v3a706c9 | !hmaster1_p & v372c23b;
assign v3a635b1 = hmaster1_p & v3a70225 | !hmaster1_p & !v37421bd;
assign v377d4a0 = hbusreq2_p & v3a7051a | !hbusreq2_p & v3a5d5d3;
assign v3a57496 = hgrant2_p & v374306c | !hgrant2_p & v3747467;
assign v3764261 = hbusreq3 & v35b7808 | !hbusreq3 & v3a67983;
assign v3a6f431 = hgrant2_p & v37709d2 | !hgrant2_p & v373b6ca;
assign v1e37784 = hmaster2_p & v3a5e24e | !hmaster2_p & b66740;
assign v374d057 = hbusreq6_p & v373bcea | !hbusreq6_p & v8455ab;
assign v3747454 = hmaster1_p & v377233c | !hmaster1_p & v3807074;
assign v3a7139c = hbusreq4 & v3760740 | !hbusreq4 & v8455ab;
assign v374cb4a = hbusreq3 & v3a6f149 | !hbusreq3 & v3748797;
assign v37767d7 = hmaster0_p & v376f53e | !hmaster0_p & !v3747dd8;
assign v3764870 = hbusreq4_p & v3a5f26f | !hbusreq4_p & v375ebe9;
assign v372cacb = hbusreq4_p & v8455ab | !hbusreq4_p & v372a1b4;
assign v3a627a4 = hgrant4_p & v37408e1 | !hgrant4_p & v372f236;
assign v3a54e41 = hmaster2_p & v376da22 | !hmaster2_p & v373698e;
assign v3776f25 = hmaster1_p & v372cc69 | !hmaster1_p & !v374610d;
assign v3a5c349 = hbusreq5_p & b5da28 | !hbusreq5_p & v3a55cda;
assign v3752987 = hmaster2_p & v8455ab | !hmaster2_p & v3a708a2;
assign v3759b93 = hlock8 & v376293b | !hlock8 & v372809b;
assign v376f92f = hlock8 & v3a58219 | !hlock8 & v372b721;
assign v3a6efb1 = hbusreq7_p & v3727b7f | !hbusreq7_p & v3752aa3;
assign v376592c = hgrant5_p & v8455ab | !hgrant5_p & v3a596a5;
assign v376d9f3 = hmaster1_p & v8455ab | !hmaster1_p & v3733557;
assign v3759569 = hmaster1_p & v8455ab | !hmaster1_p & v37559b2;
assign v3779ac2 = hgrant0_p & v8455ab | !hgrant0_p & !v37245d9;
assign v3a5c40e = hbusreq8 & v3757a2b | !hbusreq8 & v3734279;
assign v372571e = hlock5_p & v8455e7 | !hlock5_p & !v374e109;
assign v3a581bd = hready & v3a63621 | !hready & v3a70a12;
assign v3a6211e = hbusreq2_p & v3771ea6 | !hbusreq2_p & v373086c;
assign v376a9f7 = hlock5 & v372baf1 | !hlock5 & c48c9d;
assign v376a0d2 = hmaster3_p & v9864a7 | !hmaster3_p & v3722e52;
assign v372ee8a = hlock8_p & v9864ec | !hlock8_p & v2092f1b;
assign v372310a = hlock2 & v37458dc | !hlock2 & v373e521;
assign v3752869 = hgrant4_p & v374d810 | !hgrant4_p & v3a60a75;
assign v375863a = hbusreq1_p & v3723430 | !hbusreq1_p & !v3746a78;
assign c8f3d0 = hmaster3_p & v3727a2b | !hmaster3_p & v37698ab;
assign v37697ed = hmaster2_p & v376c5f3 | !hmaster2_p & v8455ab;
assign v3735fe8 = hmaster2_p & v3733ea2 | !hmaster2_p & v8455ab;
assign v37659f8 = hbusreq4_p & v3a70cdd | !hbusreq4_p & v376a877;
assign v377b68c = hbusreq3 & v375a0ff | !hbusreq3 & v373b7c8;
assign v3a2986b = jx0_p & v8455b5 | !jx0_p & v8455ab;
assign v376d2c6 = hmaster2_p & v372673d | !hmaster2_p & v3753d94;
assign v3766ddb = hgrant6_p & v374d6b2 | !hgrant6_p & v3a6ef86;
assign v3738a59 = hbusreq5 & v9af7ec | !hbusreq5 & v3774bad;
assign v377fc58 = jx1_p & v3a6d6b8 | !jx1_p & v3a556c2;
assign v377dd65 = hbusreq4 & v375f302 | !hbusreq4 & v3a6fdef;
assign v373c5a6 = hmaster2_p & v374f5e0 | !hmaster2_p & v8455ab;
assign v3761333 = hmaster0_p & v3728d9c | !hmaster0_p & v3a70453;
assign v37630a8 = hmaster1_p & v37372eb | !hmaster1_p & v375652a;
assign v3725c95 = hbusreq7_p & v3a5c2ff | !hbusreq7_p & v377b73b;
assign v3a674fd = hlock5_p & v375a878 | !hlock5_p & v376af64;
assign v37496de = hbusreq5 & v3807a23 | !hbusreq5 & v3a713c5;
assign v374b83f = hmaster3_p & v8455ab | !hmaster3_p & !v377360d;
assign v3a645b0 = hbusreq6_p & v3a57f59 | !hbusreq6_p & !v3a66110;
assign v3a66732 = hbusreq5 & v3a6f8f0 | !hbusreq5 & v372834d;
assign v3a607c3 = hmaster3_p & v8455ab | !hmaster3_p & !v3a614dd;
assign v376d6b9 = hmaster1_p & v377a104 | !hmaster1_p & !v8455ab;
assign v3a6ebf9 = hgrant6_p & v377f09a | !hgrant6_p & !v8455ab;
assign v377ba8a = hmaster2_p & v3764132 | !hmaster2_p & v3736db2;
assign v374f96e = hbusreq1_p & v37664f6 | !hbusreq1_p & v8455ab;
assign v3730122 = hbusreq3_p & v3a6f598 | !hbusreq3_p & v8455ab;
assign v377bd17 = hmaster0_p & v377c7c0 | !hmaster0_p & v3726bcc;
assign v3744b38 = hlock0_p & v8455b6 | !hlock0_p & v377e928;
assign v3736f61 = hbusreq0 & v8455b3 | !hbusreq0 & v8455ab;
assign v3767a85 = hmaster0_p & v372f151 | !hmaster0_p & v3a6b73c;
assign v37617ef = hlock4_p & v3722e5c | !hlock4_p & v35772a6;
assign v3a647f3 = hgrant0_p & v8455ab | !hgrant0_p & v3727165;
assign v376e9fd = hmaster0_p & v3745d8c | !hmaster0_p & v375d42d;
assign v377f253 = hbusreq8_p & v3737808 | !hbusreq8_p & v3a70b85;
assign v3765d5e = hbusreq5 & v3740233 | !hbusreq5 & v376f920;
assign v373bd8b = hmaster1_p & v377681e | !hmaster1_p & !v377cf71;
assign v209323b = hbusreq6_p & v3743ea8 | !hbusreq6_p & !v3a5ef5c;
assign v3a5a9e6 = hmaster2_p & v3771076 | !hmaster2_p & v3740d3b;
assign v3777467 = hmaster2_p & v3768c3c | !hmaster2_p & v3748609;
assign v3a70349 = hbusreq0 & v3a6ff37 | !hbusreq0 & v374e246;
assign v3750553 = hgrant7_p & v3a5905e | !hgrant7_p & v3729385;
assign v373b8ff = hgrant3_p & v39a4e12 | !hgrant3_p & v374fad3;
assign v3778390 = hlock6 & v3733132 | !hlock6 & v374fe7b;
assign v3a6bb45 = hgrant4_p & v8455ab | !hgrant4_p & v3761587;
assign v3a6f3b8 = hmaster0_p & v37690bf | !hmaster0_p & v3732e09;
assign v373a568 = hlock2 & v375c946 | !hlock2 & v3754877;
assign v3745c45 = hmaster2_p & v374502e | !hmaster2_p & !v3a6fcba;
assign v3726cf7 = hlock3_p & v376e914 | !hlock3_p & !v3a658bf;
assign v3a67dd5 = hmaster0_p & v37332af | !hmaster0_p & v3a296dc;
assign v3730da3 = hlock1 & v37306bb | !hlock1 & v3741e9d;
assign v372e6ee = hbusreq2 & d44200 | !hbusreq2 & v8455ab;
assign c08050 = hlock8_p & v373741d | !hlock8_p & v3a5ab24;
assign v3775e81 = hgrant4_p & v8455ab | !hgrant4_p & v375d4d4;
assign v1e37339 = hlock4 & v3a6f69f | !hlock4 & v372fff3;
assign v375b9e1 = hbusreq6_p & v3a70aa2 | !hbusreq6_p & v374c9db;
assign v37538ff = hlock4_p & v3724e8e | !hlock4_p & v3763a20;
assign v373867c = hgrant2_p & v3a69487 | !hgrant2_p & v3a6ef1f;
assign v3a6fee8 = hbusreq3 & v3728e09 | !hbusreq3 & !v8455ab;
assign v3a5f5e8 = hbusreq0 & v3a65212 | !hbusreq0 & v3733542;
assign v3a6006c = hgrant2_p & v3a70dc4 | !hgrant2_p & v3755bc2;
assign v3768d11 = hmaster2_p & v3a63805 | !hmaster2_p & v375ac23;
assign v3738bf6 = hmaster0_p & v37419e7 | !hmaster0_p & !v37455cd;
assign v373f08d = hmaster0_p & v3a5c369 | !hmaster0_p & v3577392;
assign v3a710c4 = hmaster2_p & v3750746 | !hmaster2_p & v3a637dd;
assign v3a70c19 = hgrant4_p & v3a635ea | !hgrant4_p & v3a63c15;
assign v373e474 = hgrant4_p & v3a6fac2 | !hgrant4_p & v37310be;
assign v3a5d7ba = hmaster2_p & v37358ab | !hmaster2_p & v3a67a6f;
assign v376d882 = hbusreq2_p & v8455ab | !hbusreq2_p & v374fb58;
assign v37363fd = hlock6_p & v3a70385 | !hlock6_p & !v8455ab;
assign v373a3a7 = hbusreq8_p & v3a67b3c | !hbusreq8_p & v3a70342;
assign v372dfba = hbusreq5_p & v3a70980 | !hbusreq5_p & v3a65711;
assign v3756526 = hbusreq7_p & v3a6501d | !hbusreq7_p & v3a5db7d;
assign jx0 = v3a63994;
assign v3a606a0 = hmaster0_p & v3750296 | !hmaster0_p & v377904f;
assign v373c81c = hbusreq6_p & v37778cf | !hbusreq6_p & v372abc8;
assign v37369eb = hgrant2_p & v8455ab | !hgrant2_p & v3741833;
assign v377efe1 = hbusreq5 & v3a7046e | !hbusreq5 & v8455ab;
assign v37452c7 = hgrant2_p & v3a7134d | !hgrant2_p & v3a71088;
assign v376fca4 = hbusreq4_p & v3a54ba7 | !hbusreq4_p & v380947a;
assign v3768a1c = hmaster0_p & v376db87 | !hmaster0_p & v3a6f275;
assign v8fac55 = hgrant4_p & v8455ab | !hgrant4_p & v3727df1;
assign v3730862 = hbusreq7_p & v374f834 | !hbusreq7_p & v3a6accb;
assign v3a6793d = hmaster0_p & v372adfd | !hmaster0_p & v3728fda;
assign v375da95 = hlock6_p & v377ba55 | !hlock6_p & !v8455ab;
assign v37287fb = hgrant5_p & v994115 | !hgrant5_p & v376d522;
assign v377b26a = hmaster0_p & v376301d | !hmaster0_p & v3a553db;
assign v3738d19 = hlock5_p & v3779883 | !hlock5_p & !v373a692;
assign v3a70bf8 = hmaster2_p & v3731b41 | !hmaster2_p & v3a71276;
assign v3a6f451 = hmaster2_p & v3763c09 | !hmaster2_p & v374d54c;
assign v3a63e51 = hlock8_p & v3a53e5c | !hlock8_p & !v8455ab;
assign v3736a50 = hlock5_p & v8455ab | !hlock5_p & v3a5d644;
assign v3a62e7b = jx0_p & b8ed55 | !jx0_p & v8455ab;
assign v3764de7 = hgrant6_p & v3772362 | !hgrant6_p & v3a6065f;
assign v373fbc9 = hbusreq6_p & v3a643d7 | !hbusreq6_p & v377728d;
assign v3a63f05 = stateG10_1_p & v3a70d71 | !stateG10_1_p & v37443d6;
assign v37719a1 = hmaster2_p & v376728e | !hmaster2_p & v8455b9;
assign v3a62582 = hbusreq6_p & v3a70c1b | !hbusreq6_p & v8455ab;
assign v3750cae = hmaster2_p & v8455ab | !hmaster2_p & v377f67b;
assign v3a6797d = hmaster1_p & v8455ab | !hmaster1_p & v3765a69;
assign v3734af6 = hbusreq2 & v8455ab | !hbusreq2 & !v373aecf;
assign v3748964 = hbusreq6 & v3775165 | !hbusreq6 & v3a575d6;
assign v3762498 = hbusreq6 & v373014d | !hbusreq6 & v8455bf;
assign v372f98a = hbusreq7_p & v3a637a5 | !hbusreq7_p & v37405a3;
assign v373e74b = hmaster2_p & v3a71133 | !hmaster2_p & v372eab1;
assign v3a648d0 = hbusreq6 & v3a625f8 | !hbusreq6 & v3a58102;
assign v374a91e = hbusreq0 & v37307dd | !hbusreq0 & v8455ab;
assign v37478bc = hmaster0_p & v3a6a52b | !hmaster0_p & v376b031;
assign v376081b = hgrant4_p & v372b77b | !hgrant4_p & v3773fbb;
assign v37439ef = hmaster1_p & v373823d | !hmaster1_p & v37615d0;
assign v37541d4 = hmaster1_p & v375c573 | !hmaster1_p & v3762613;
assign v3723c3f = hmaster2_p & v3a71133 | !hmaster2_p & v3779cc0;
assign v3756f41 = hbusreq5 & v375a269 | !hbusreq5 & v8455ab;
assign v3a6f323 = hlock0 & v3807d59 | !hlock0 & v37513bc;
assign v376a25e = hgrant8_p & v8455cd | !hgrant8_p & v372c046;
assign v3753b93 = hlock8_p & v8455ab | !hlock8_p & v376b829;
assign v376b33c = hgrant0_p & v3a7014c | !hgrant0_p & v3a68426;
assign v376e35e = hgrant4_p & v3a71016 | !hgrant4_p & v3733726;
assign v376550d = hbusreq7_p & v376b5c0 | !hbusreq7_p & v3a66529;
assign v377e158 = hgrant2_p & v377b6ce | !hgrant2_p & v375e232;
assign v3a6f973 = hbusreq8_p & v372d6fa | !hbusreq8_p & !v372ac64;
assign v3a6f75c = hbusreq0 & v37724f9 | !hbusreq0 & v3751b42;
assign v377ef71 = hlock5 & v37634d0 | !hlock5 & v372ab6c;
assign v37607af = hmaster2_p & v3a5e696 | !hmaster2_p & v8455ab;
assign v3767e15 = hgrant2_p & v37699a0 | !hgrant2_p & v3750f4b;
assign v3765293 = jx3_p & v374f34b | !jx3_p & v375dcf8;
assign v3747aa5 = hlock5_p & v3a5943e | !hlock5_p & !v373b956;
assign v3729f6a = hgrant2_p & v3a69487 | !hgrant2_p & v3750859;
assign v3a7054d = hbusreq8 & v373be40 | !hbusreq8 & b79c3c;
assign v3a6f059 = hbusreq4_p & v3748797 | !hbusreq4_p & v376d92b;
assign v3a6f9f5 = hbusreq4_p & v373ae0a | !hbusreq4_p & v373dc68;
assign v3768c3c = hbusreq2_p & v3a5891c | !hbusreq2_p & v3759032;
assign v372ef80 = hmaster2_p & v3759031 | !hmaster2_p & v3a70cc3;
assign v37688a5 = hburst0_p & v8455ab | !hburst0_p & v3726abd;
assign v3a7151f = hbusreq7 & v3a6324e | !hbusreq7 & v372cf51;
assign v377c003 = hgrant2_p & v8455ab | !hgrant2_p & v377d047;
assign v3746473 = hbusreq5_p & v372d4eb | !hbusreq5_p & v3a5f4c6;
assign v3747079 = hgrant5_p & v8455ab | !hgrant5_p & v372d060;
assign v3a6277d = hbusreq8_p & v3744cf7 | !hbusreq8_p & v374abb5;
assign v3749f2e = hmaster1_p & v37c36c4 | !hmaster1_p & !v373b7dd;
assign v3769616 = hbusreq3 & v374ace7 | !hbusreq3 & v3726006;
assign v3a61220 = hgrant6_p & v37304b3 | !hgrant6_p & v373ee41;
assign v3a713cc = hlock4_p & v3a5600a | !hlock4_p & v8455b0;
assign v3a7047f = hbusreq2_p & v37502d4 | !hbusreq2_p & v8455ab;
assign v3773fbb = hgrant6_p & v8455ab | !hgrant6_p & v375efa1;
assign ade0d8 = hgrant6_p & v8455ab | !hgrant6_p & v3a62582;
assign v3a7104b = hbusreq1_p & v3a6fe6a | !hbusreq1_p & v3739443;
assign v3a5c779 = hbusreq3_p & v3a69529 | !hbusreq3_p & !v8455ab;
assign v3807b2e = hmaster0_p & v374cc40 | !hmaster0_p & !v3a702e9;
assign v3a63f6b = hmaster1_p & v37386c6 | !hmaster1_p & v380925f;
assign v3a705db = hgrant2_p & v3a70645 | !hgrant2_p & v3a5fd34;
assign v375e01c = hbusreq6 & v3778993 | !hbusreq6 & v8455ab;
assign v373b6c0 = hbusreq6 & v3a6f9b9 | !hbusreq6 & v373d293;
assign v377f501 = hbusreq7_p & v37734cb | !hbusreq7_p & v375e813;
assign v375abcd = hlock2 & v3806ff0 | !hlock2 & v374fd4a;
assign v3728abd = hlock5_p & v3743327 | !hlock5_p & !v3762552;
assign v3729d1b = hbusreq3_p & v37482c8 | !hbusreq3_p & v8455ab;
assign v3a70255 = hgrant6_p & v3747c3e | !hgrant6_p & v8455ab;
assign v377746e = hgrant4_p & v3a70fe9 | !hgrant4_p & v3772310;
assign v3a71422 = hbusreq1_p & v377122d | !hbusreq1_p & !v3a5bbed;
assign v374f31c = hmaster1_p & v374a454 | !hmaster1_p & v3764628;
assign v37622f5 = hbusreq4_p & v3754b79 | !hbusreq4_p & v3749cf7;
assign v3a703f6 = hgrant5_p & v3727d4c | !hgrant5_p & v376078d;
assign v3746008 = hmaster0_p & v3a680e1 | !hmaster0_p & v373058e;
assign cf3b5d = hbusreq1_p & v3a635ea | !hbusreq1_p & v37265b3;
assign v3a60649 = hmaster2_p & v3a63777 | !hmaster2_p & v3a663b9;
assign v374b7f6 = hbusreq5_p & v3728fa6 | !hbusreq5_p & v374eddc;
assign v3a6205a = hbusreq8 & v3a62cb5 | !hbusreq8 & v3a67beb;
assign v376ee80 = hbusreq4 & v376ebbf | !hbusreq4 & v3a60a68;
assign v3807aa1 = hbusreq4_p & v37314cc | !hbusreq4_p & v8455ab;
assign v3a61a7f = hlock0_p & v8455ab | !hlock0_p & v3a635ea;
assign v37258c9 = hbusreq3_p & v3a7045c | !hbusreq3_p & v3765a43;
assign v37330dc = hbusreq4_p & v377b330 | !hbusreq4_p & v3743b9e;
assign v373350e = hbusreq0 & ad3125 | !hbusreq0 & v8455b0;
assign v3a70473 = hgrant8_p & v3a61796 | !hgrant8_p & v3767ba9;
assign v37259c7 = hgrant6_p & v3722e5c | !hgrant6_p & v3767420;
assign v37411ab = hmaster0_p & v2acb5c7 | !hmaster0_p & v372d51c;
assign v3a574d7 = hbusreq8 & v372a288 | !hbusreq8 & v374d617;
assign v377b920 = hgrant5_p & v3736df1 | !hgrant5_p & v3a6fb4b;
assign v3a66514 = hmaster0_p & v373f503 | !hmaster0_p & v3732c95;
assign v376bb05 = hbusreq6 & v376b4a8 | !hbusreq6 & v3a6ebcc;
assign v374e3ab = hgrant5_p & v3743dc4 | !hgrant5_p & v3728bc3;
assign d1331f = hready_p & v376ee08 | !hready_p & v37250af;
assign v3750218 = hmaster2_p & v3778cf7 | !hmaster2_p & !v3a70fec;
assign v376bd43 = hgrant4_p & v8455ab | !hgrant4_p & b12fe4;
assign v3734f6d = hbusreq5_p & v3a714b9 | !hbusreq5_p & !v3a5af94;
assign v37245f8 = hbusreq2_p & v374c47e | !hbusreq2_p & v8455b0;
assign v3740ed1 = hmaster1_p & v3778372 | !hmaster1_p & v372ab0f;
assign v377221f = hlock6 & v3a70186 | !hlock6 & v3a6f9a2;
assign v37666dd = hbusreq0 & v3a5bb4f | !hbusreq0 & v372998a;
assign v373583d = hbusreq4 & v3a608b9 | !hbusreq4 & !v1e37e82;
assign v375b96f = hmaster0_p & v3a6950d | !hmaster0_p & v8455ab;
assign v325b59d = hmaster2_p & v3a6e5f0 | !hmaster2_p & v3a70c39;
assign v3a703aa = hmaster0_p & v374674d | !hmaster0_p & v3735485;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hbusreq2_p = 0;
  hlock2_p = 0;
  hbusreq3_p = 0;
  hlock3_p = 0;
  hbusreq4_p = 0;
  hlock4_p = 0;
  hbusreq5_p = 0;
  hlock5_p = 0;
  hbusreq6_p = 0;
  hlock6_p = 0;
  hbusreq7_p = 0;
  hlock7_p = 0;
  hbusreq8_p = 0;
  hlock8_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmaster1_p = 0;
  hmaster2_p = 0;
  hmaster3_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  hgrant2_p = 0;
  hgrant3_p = 0;
  hgrant4_p = 0;
  hgrant5_p = 0;
  hgrant6_p = 0;
  hgrant7_p = 0;
  hgrant8_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  stateG10_2_p = 0;
  stateG10_3_p = 0;
  stateG10_4_p = 0;
  stateG10_5_p = 0;
  stateG10_6_p = 0;
  stateG10_7_p = 0;
  stateG10_8_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
  jx3_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hbusreq2_p = hbusreq2;
  hlock2_p = hlock2;
  hbusreq3_p = hbusreq3;
  hlock3_p = hlock3;
  hbusreq4_p = hbusreq4;
  hlock4_p = hlock4;
  hbusreq5_p = hbusreq5;
  hlock5_p = hlock5;
  hbusreq6_p = hbusreq6;
  hlock6_p = hlock6;
  hbusreq7_p = hbusreq7;
  hlock7_p = hlock7;
  hbusreq8_p = hbusreq8;
  hlock8_p = hlock8;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmaster1_p = hmaster1;
  hmaster2_p = hmaster2;
  hmaster3_p = hmaster3;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  hgrant2_p = hgrant2;
  hgrant3_p = hgrant3;
  hgrant4_p = hgrant4;
  hgrant5_p = hgrant5;
  hgrant6_p = hgrant6;
  hgrant7_p = hgrant7;
  hgrant8_p = hgrant8;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  stateG10_2_p = stateG10_2;
  stateG10_3_p = stateG10_3;
  stateG10_4_p = stateG10_4;
  stateG10_5_p = stateG10_5;
  stateG10_6_p = stateG10_6;
  stateG10_7_p = stateG10_7;
  stateG10_8_p = stateG10_8;
  jx0_p = jx0;
  jx1_p = jx1;
  jx2_p = jx2;
  jx3_p = jx3;
    end
endmodule

