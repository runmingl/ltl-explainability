module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hburst0, hburst1, hmaster0, hmastlock, start, decide, locked, hgrant0, hgrant1, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, jx0, jx1);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v845800;
  wire v845810;
  wire v85cd0b;
  wire v857931;
  wire v864279;
  wire v8822a8;
  wire v88235e;
  wire v86170f;
  wire v8afeef;
  wire v845822;
  wire v882343;
  wire v8b9eb8;
  wire v8b9f20;
  wire v8a05fa;
  wire v8b9dcc;
  wire v8a0613;
  wire v863615;
  wire v88d08c;
  wire v85803c;
  wire v895141;
  wire v85cd0c;
  wire v8822ff;
  wire v859575;
  wire v85f58f;
  wire v862346;
  wire v882363;
  wire v857768;
  wire v85bc42;
  wire v8b9dc2;
  wire v8823ab;
  wire v88ffc8;
  wire v858af8;
  wire v895133;
  wire v8b9e9a;
  wire v85f58b;
  wire v85968b;
  wire v8698e6;
  wire v8b9f40;
  wire v882332;
  wire v895151;
  wire v8a05fe;
  wire v8554b2;
  wire v8b9ead;
  wire v8b71ab;
  wire v88237d;
  wire v8b9f77;
  wire v856e69;
  wire v85c621;
  wire v8b9ddc;
  wire v8822e3;
  wire v88d077;
  wire v85f596;
  wire v88d062;
  wire v85f597;
  wire v8b9e4f;
  wire v88228f;
  wire v88706d;
  wire v857eb6;
  wire v864a19;
  wire v85688b;
  wire v85ce00;
  wire v858768;
  wire v858cdb;
  wire v861c72;
  wire v864523;
  wire v85c719;
  wire v85e7b1;
  wire v864246;
  wire v8b9f98;
  wire v8583bf;
  wire v85b4d5;
  wire v850b73;
  wire v8856cf;
  wire v8612b9;
  wire v8b9e28;
  wire v85e3ad;
  wire v855784;
  wire v885c50;
  wire v8b9e88;
  wire v86240b;
  wire v8b9e06;
  wire v88237a;
  wire v88ffbb;
  wire v8b9efd;
  wire v85f5c7;
  wire v84581e;
  wire v8a0282;
  wire v85598d;
  wire v845826;
  wire v86022a;
  wire v85a970;
  wire v860967;
  wire v8b9da5;
  wire v8539e6;
  wire v85f907;
  wire v845828;
  wire v8b9e9b;
  wire v85c5ce;
  wire v8afee6;
  wire v88705d;
  wire v85a4b1;
  wire v88234f;
  wire v85791c;
  wire v8b9f3b;
  wire v8a0606;
  wire v8b9ddd;
  wire v850c63;
  wire v88229c;
  wire v8b9e3e;
  wire v863070;
  wire v85f57f;
  wire v85f6d6;
  wire v882365;
  wire v8578ef;
  wire v85bae3;
  wire v882381;
  wire v8a0623;
  wire v85e961;
  wire v8620e6;
  wire v8b9ed6;
  wire v88232a;
  wire v85adda;
  wire v885713;
  wire v882370;
  wire v85880f;
  wire v8b9dc4;
  wire v895157;
  wire v845804;
  wire v8aff0a;
  wire v86216f;
  wire v893788;
  wire v84582a;
  wire v8b9e90;
  wire v89514a;
  wire v862e72;
  wire v85ef57;
  wire v88d07b;
  wire v8aff10;
  wire v8a060b;
  wire v8b9e2a;
  wire v85a3c2;
  wire v882348;
  wire v8b9e57;
  wire v882328;
  wire v8b9ed0;
  wire v8b9ded;
  wire v85d8f3;
  wire v8822c3;
  wire v862e32;
  wire v8b9dd5;
  wire v88ffd1;
  wire v895135;
  wire v852480;
  wire v8a062c;
  wire v882369;
  wire v8b9e30;
  wire v860c97;
  wire v85a8a7;
  wire v88ffd5;
  wire v8b9e25;
  wire v859163;
  wire v85a3f3;
  wire v85b2d4;
  wire v8b9e17;
  wire v85dfb4;
  wire v850cb2;
  wire v8856cb;
  wire v85f5c3;
  wire v858a13;
  wire v887053;
  wire v864941;
  wire v85abe0;
  wire v8579d6;
  wire v85bc80;
  wire v8823a5;
  wire v856c47;
  wire v856a41;
  wire v8aff0b;
  wire v85d0b4;
  wire v861ed5;
  wire v8b9f81;
  wire v85ff1e;
  wire v8b9e56;
  wire v85bc9e;
  wire v85f1d9;
  wire v8b9deb;
  wire v862d65;
  wire v85877f;
  wire v858df2;
  wire v8b9e5f;
  wire v853647;
  wire v855d31;
  wire v8a065d;
  wire v8b9e92;
  wire v8531a0;
  wire v85cbe8;
  wire v85f589;
  wire v8b9efe;
  wire v8551f3;
  wire v861546;
  wire v85f583;
  wire v8afee8;
  wire v85af06;
  wire v863359;
  wire v8581c3;
  wire v85957f;
  wire v8afef8;
  wire v885722;
  wire v84581a;
  wire v845814;
  wire v8b9dd1;
  wire v858df5;
  wire v8822be;
  wire v8a061b;
  wire v88d05e;
  wire v8b9e1c;
  wire v8b9f3f;
  wire v8822f4;
  wire v856d8f;
  wire v855cc1;
  wire v858d97;
  wire v8b9e0e;
  wire v8b9ea9;
  wire v845808;
  wire v860b53;
  wire v845818;
  wire v88231d;
  wire v88236f;
  wire v864e1f;
  wire v84580e;
  wire v85f5ba;
  wire v882340;
  wire v882344;
  wire v8b9f06;
  wire v861aaf;
  wire v8b9f35;
  wire v88233e;
  wire v85263d;
  wire v8b9e13;
  wire v8a0615;
  wire v8b9dc5;
  wire v85cb28;
  wire v85f1f2;
  wire v8822bb;
  wire v85323a;
  wire v86042c;
  wire v8b9e74;
  wire v88d044;
  wire v8606e5;
  wire v8a0611;
  wire v8856c6;
  wire v882307;
  wire v850934;
  wire v88228e;
  wire v85a7d6;
  wire v85d087;
  wire v8a0653;
  wire v8b9e32;
  wire v8822cc;
  wire v85331f;
  wire v8a065b;
  wire v8b9ec7;
  wire v8628c9;
  wire v8539e3;
  wire v8631b2;
  wire v88d069;
  wire v88d085;
  wire v8b9f5a;
  wire v8b9f58;
  wire v8b9ec8;
  wire v858dca;
  wire v85e315;
  wire v85c62e;
  wire v858327;
  wire v861211;
  wire v8b9eaf;
  wire v8822c4;
  wire v85f67e;
  wire v8b9eed;
  wire v8b9e60;
  wire v8b9f6a;
  wire v85f599;
  wire v85add4;
  wire v8b9db3;
  wire v8b71a8;
  wire v8b9e46;
  wire v887066;
  wire v882292;
  wire v8b9dbd;
  wire v8b9df4;
  wire v8a064d;
  wire v85e753;
  wire v85029d;
  wire v8b9edf;
  wire v8b9dc3;
  wire v8612af;
  wire v85f5a3;
  wire v856316;
  wire v8b9dba;
  wire v88239e;
  wire v88706c;
  wire v858525;
  wire v85e30c;
  wire v8b9dbf;
  wire v88228d;
  wire v88a7bc;
  wire v8b9f21;
  wire v852a1d;
  wire v8597ea;
  wire v85ce69;
  wire v855d10;
  wire v887054;
  wire v88a7b1;
  wire v85330e;
  wire v855460;
  wire v8a0641;
  wire v8822d5;
  wire v85654f;
  wire v8a0630;
  wire v850ce7;
  wire v85b5d3;
  wire v8612ae;
  wire v885718;
  wire v8637b3;
  wire v8b9f64;
  wire v85f5b5;
  wire v8591b7;
  wire v85f5b3;
  wire v8545f6;
  wire v859ca9;
  wire v8b9e8f;
  wire v88d074;
  wire v862090;
  wire v8a065e;
  wire v84580c;
  wire v862e59;
  wire v85315d;
  wire v88d04d;
  wire v8b9dcf;
  wire v852c3b;
  wire v8602a4;
  wire v8822a3;
  wire v85c9ad;
  wire v88d076;
  wire v8b9f6e;
  wire v85f5c5;
  wire v8b9f14;
  wire v85e71f;
  wire v88a7a9;
  wire v882349;
  wire v863eb5;
  wire v859d97;
  wire v86027d;
  wire v8b9ee9;
  wire v85c278;
  wire v8b9e04;
  wire v8856ee;
  wire v85f5b1;
  wire v88238f;
  wire v8a0609;
  wire v8b9e1f;
  wire v85c572;
  wire v8856f0;
  wire v8a065c;
  wire v8a0621;
  wire v8b9e7e;
  wire v8569be;
  wire v8822b1;
  wire v88d056;
  wire v8b9dff;
  wire v88d08e;
  wire v8b9f60;
  wire v853997;
  wire v8b9e52;
  wire v88230b;
  wire v85bab4;
  wire v887069;
  wire v85ce61;
  wire v8822d8;
  wire v857e7d;
  wire v85ff2e;
  wire v8523bf;
  wire v85fa6a;
  wire v8632bb;
  wire v85ca17;
  wire v862032;
  wire v88a7bd;
  wire v85f85f;
  wire v8823a9;
  wire v88238b;
  wire v85ad75;
  wire v862c91;
  wire v8b9e51;
  wire v887059;
  wire v858ab6;
  wire v8b9e66;
  wire v8a0640;
  wire v8a062d;
  wire v85b3e2;
  wire v85fbe0;
  wire v8b71a6;
  wire v860700;
  wire v882342;
  wire v85d9d7;
  wire v882304;
  wire v851c6c;
  wire v85f582;
  wire v8856e0;
  wire v85f6f8;
  wire v88ffbf;
  wire v8b9e22;
  wire v8aff12;
  wire v863af6;
  wire v89a6f2;
  wire v852ef0;
  wire v862224;
  wire v8822da;
  wire v85e2a8;
  wire v85b6dd;
  wire v8822c1;
  wire v85d046;
  wire v8b9ef5;
  wire v85465f;
  wire v8b9f26;
  wire v8633f4;
  wire v85a826;
  wire v88233c;
  wire v88d070;
  wire v853cad;
  wire v8b71b0;
  wire v84580b;
  wire v845807;
  wire v88d051;
  wire v8b71ae;
  wire v85de6c;
  wire v8b9e67;
  wire v89a6f5;
  wire v84580a;
  wire v852578;
  wire v845806;
  wire v851b6e;
  wire v8b9e5c;
  wire v851d36;
  wire v8b9f39;
  wire v855bfd;
  wire v8a05f1;
  wire v88d087;
  wire v882375;
  wire v8a062b;
  wire v88d040;
  wire v863a8a;
  wire v85f7a7;
  wire v8578f2;
  wire v8b9f09;
  wire v862f96;
  wire v858794;
  wire v88705c;
  wire v85f588;
  wire v85d0f7;
  wire v8b9e50;
  wire v8628dd;
  wire v854a42;
  wire v8533a0;
  wire v85736e;
  wire v8b9dca;
  wire v85f5b2;
  wire v845816;
  wire v88d088;
  wire v8b9df7;
  wire v8b9f8f;
  wire v85e7e0;
  wire v8aff0f;
  wire v853cf6;
  wire v8b9db6;
  wire v8856ca;
  wire v864990;
  wire v861acc;
  wire v85cb5c;
  wire v8b9da6;
  wire v8b9dc1;
  wire v8629ac;
  wire v882395;
  wire v882287;
  wire v8b9f57;
  wire v882282;
  wire v8afefc;
  wire v88d046;
  wire v852475;
  wire v851b5f;
  wire v860fce;
  wire v864cfd;
  wire v8afef1;
  wire v8b9dce;
  wire v8822d2;
  wire v853612;
  wire v85ae93;
  wire v8856da;
  wire v8505a9;
  wire v859474;
  wire v85f59a;
  wire v86223c;
  wire v8607e4;
  wire v882373;
  wire v85fec2;
  wire v8606fb;
  wire v882376;
  wire v85ee66;
  wire v8822d4;
  wire v8b9f11;
  wire v8a05f0;
  wire v85a3e3;
  wire v8b9e59;
  wire v856019;
  wire v860719;
  wire v85215e;
  wire v85ee90;
  wire v864411;
  wire v8b9e4b;
  wire v8b71ac;
  wire v8a0610;
  wire v88d071;
  wire v864711;
  wire v85c7f3;
  wire v885719;
  wire v88d090;
  wire v85e4a1;
  wire v8aff00;
  wire v8b9ec9;
  wire v88d07c;
  wire v88231f;
  wire v8822f3;
  wire v8b9de1;
  wire v85c7fb;
  wire v8b9e55;
  wire v8b9e19;
  wire v85d820;
  wire v8b9f5d;
  wire v85b83a;
  wire v85d6d3;
  wire v85f58e;
  wire v88d06e;
  wire v8571d1;
  wire v882338;
  wire v864244;
  wire v863d0e;
  wire v8822fc;
  wire v8b9f71;
  wire v8b71aa;
  wire v8b9e35;
  wire v8b9e0c;
  wire v88ffbd;
  wire v857eeb;
  wire v8822ad;
  wire v857fb9;
  wire v88a7b4;
  wire v85a5c7;
  wire v8b9e1e;
  wire v85c70f;
  wire v887064;
  wire v8647b7;
  wire v882390;
  wire v88a7ca;
  wire v85ac94;
  wire v8822c6;
  wire v8b9ea8;
  wire v861f20;
  wire v85fb02;
  wire v8b9f4d;
  wire v8b9e1d;
  wire v88229d;
  wire v88d061;
  wire v89a6f4;
  wire v8b9ed3;
  wire v86997d;
  wire v85f1f3;
  wire v85c3b7;
  wire v85cc6b;
  wire v8b9dec;
  wire v85e13d;
  wire v85fe4d;
  wire v87fd78;
  wire v8a0602;
  wire v89513e;
  wire v860625;
  wire v8b9ee3;
  wire v85f5bf;
  wire v8b9ed5;
  wire v858fd3;
  wire v853c79;
  wire v8a05f8;
  wire v85cb98;
  wire v8b9e75;
  wire v8b9f56;
  wire v8b9f0a;
  wire v8618bd;
  wire v88706f;
  wire v864631;
  wire v8b9e0f;
  wire v882310;
  wire v8b9e26;
  wire v85f141;
  wire v895132;
  wire v85f5ad;
  wire v8b9f27;
  wire v85e7fa;
  wire v882382;
  wire v885c52;
  wire v8a0633;
  wire v85fad3;
  wire v856300;
  wire v85a015;
  wire v8a0632;
  wire v8631cf;
  wire v8b9f51;
  wire v863b11;
  wire v862857;
  wire v88d073;
  wire v85a414;
  wire v882306;
  wire v860b2a;
  wire v8623ae;
  wire v8617ee;
  wire v85c5b2;
  wire v851b5e;
  wire v855817;
  wire v887065;
  wire v8562e6;
  wire v882392;
  wire v85f592;
  wire v8a064b;
  wire v8b9ea0;
  wire v8b9f44;
  wire v855725;
  wire v8b9e3d;
  wire v85fb94;
  wire v8856df;
  wire v8afefa;
  wire v8b9de6;
  wire v8600bd;
  wire v85a1b1;
  wire v8822f1;
  wire v8605e3;
  wire v8556fc;
  wire v8b9e0b;
  wire v8b9dbe;
  wire v8b9f4c;
  wire v8856dd;
  wire v859134;
  wire v86314b;
  wire v8b9e2d;
  wire v852edf;
  wire v85b585;
  wire v862f60;
  wire v8b9dee;
  wire v84580f;
  wire v8822c2;
  wire v88ffba;
  wire v87fd7a;
  wire v85a031;
  wire v8b9e44;
  wire v8a05fc;
  wire v86192f;
  wire v88ffd0;
  wire v882355;
  wire v86031b;
  wire v8afefe;
  wire v862f88;
  wire v8b9f17;
  wire v8822ef;
  wire v86482d;
  wire v857e81;
  wire v8b9e11;
  wire v8b9eb4;
  wire v8823b0;
  wire v8b9e6d;
  wire v887062;
  wire v85af59;
  wire v895152;
  wire v85f5c1;
  wire v882285;
  wire v85f81e;
  wire v85c750;
  wire v882351;
  wire v85a595;
  wire v862ad8;
  wire v8b9ecf;
  wire v864cae;
  wire v885c4f;
  wire v88234d;
  wire v85e920;
  wire v85b9f7;
  wire v882345;
  wire v85596e;
  wire v885700;
  wire v8822f8;
  wire v85afd6;
  wire v8b9f80;
  wire v8aff0d;
  wire v88231a;
  wire v8822e2;
  wire v845824;
  wire v86028b;
  wire v8a0639;
  wire v85dedf;
  wire v85c75d;
  wire v8b9e85;
  wire v85ca1b;
  wire v8b9de7;
  wire v86195f;
  wire v882316;
  wire v8b9f0e;
  wire v864183;
  wire v8823a4;
  wire v8b9ea4;
  wire v857751;
  wire v88d06f;
  wire v8b9dcd;
  wire v861bb9;
  wire v87fd7e;
  wire v861c42;
  wire v859035;
  wire v8aff05;
  wire v882305;
  wire v8b9ef0;
  wire v87fd7f;
  wire v88a7c6;
  wire v8619fc;
  wire v8856d5;
  wire v88a7b5;
  wire v8afef9;
  wire v88d066;
  wire v8822e6;
  wire v85e54f;
  wire v8822c8;
  wire v852fbe;
  wire v852fc6;
  wire v8b9e34;
  wire v8b9f48;
  wire v88ffcf;
  wire v895134;
  wire v8b9e0d;
  wire v85d6b5;
  wire v8635aa;
  wire v8822fe;
  wire v8b9e97;
  wire v8b9ed7;
  wire v88237e;
  wire v85e25a;
  wire v860fbc;
  wire v87fd83;
  wire v862ee4;
  wire v88229f;
  wire v88d05f;
  wire v8b9def;
  wire v8518b8;
  wire v8822cd;
  wire v882317;
  wire v88ffc2;
  wire v85f58d;
  wire v85f5c2;
  wire v85f5af;
  wire v8b9dfc;
  wire v8b9e6c;
  wire v8b9f03;
  wire v8628b1;
  wire v88705e;
  wire v8b9ea7;
  wire v851cd0;
  wire v8b9e4a;
  wire v8626cc;
  wire v8a060a;
  wire v860857;
  wire v8b9dc6;
  wire v863bff;
  wire v88237f;
  wire v8b9f13;
  wire v8b9dd8;
  wire v88d080;
  wire v85f581;
  wire v862a20;
  wire v8b9e20;
  wire v858891;
  wire v8b9de4;
  wire v862f33;
  wire v8535f8;
  wire v8822e0;
  wire v85934d;
  wire v8b9e21;
  wire v88a7b7;
  wire v88a7ba;
  wire v845805;
  wire v861063;
  wire v8b9f69;
  wire v8822cf;
  wire v853437;
  wire v882326;
  wire v88a7a3;
  wire v8822ac;
  wire v85a9a4;
  wire v88230e;
  wire v8856d4;
  wire v860c3a;
  wire v8a0620;
  wire v88238a;
  wire v8b9e47;
  wire v856288;
  wire v8822b0;
  wire v8b9e41;
  wire v8a062a;
  wire v8822fa;
  wire v864525;
  wire v8a0648;
  wire v8822b6;
  wire v8b9fa4;
  wire v89a6f1;
  wire v8b9ee7;
  wire v89513a;
  wire v8a0618;
  wire v863d44;
  wire v88ffc1;
  wire v8b9e12;
  wire v8822e7;
  wire v8b9ef1;
  wire v88ffc0;
  wire v858cf2;
  wire v8afee2;
  wire v8b9f4f;
  wire v8b9dc7;
  wire v8b9e00;
  wire v88d052;
  wire v885702;
  wire v8520a6;
  wire v8b9e2c;
  wire v85f5a5;
  wire v8b9f6c;
  wire v85f5ac;
  wire v8508b4;
  wire v851256;
  wire v8b9dbb;
  wire v8b71a5;
  wire v8b9f34;
  wire v8b9fa2;
  wire v85d0f1;
  wire v8b9e49;
  wire v88a7c9;
  wire v87fd84;
  wire v85923c;
  wire v8856d6;
  wire v8856e1;
  wire v85fd24;
  wire v852071;
  wire v8530df;
  wire v8822b5;
  wire v882379;
  wire v859006;
  wire v8523de;
  wire v85f5b7;
  wire v85f5be;
  wire v85d6af;
  wire v8b9eb2;
  wire v8afeed;
  wire v88d07d;
  wire v882325;
  wire v85e4e6;
  wire v85f1ae;
  wire v860568;
  wire v85b113;
  wire v8b9e7b;
  wire v852bf7;
  wire v8823af;
  wire v88d06d;
  wire v85f0c6;
  wire v862a8d;
  wire v88d057;
  wire v859d8d;
  wire v861fa1;
  wire v8b71ad;
  wire v85cd3f;
  wire v88705a;
  wire v882354;
  wire v882291;
  wire v8aff03;
  wire v85c4a2;
  wire v861d53;
  wire v88228b;
  wire v8b9e2f;
  wire v853308;
  wire v85c974;
  wire v860f3e;
  wire v88235a;
  wire v88a7aa;
  wire v8a0649;
  wire v8b9e8b;
  wire v8b9f90;
  wire v85c89c;
  wire v882391;
  wire v85f57e;
  wire v8823b4;
  wire v895139;
  wire v8b9e72;
  wire v85d667;
  wire v862097;
  wire v8b9e31;
  wire v8b9e1b;
  wire v8b9f18;
  wire v8856c9;
  wire v8b9e9f;
  wire v88230c;
  wire v882399;
  wire v85c59b;
  wire v8afef6;
  wire v87fd86;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;

assign v8b71a6 = decide_p & v85fbe0 | !decide_p & v84581a;
assign v8aff0f = locked_p & v8b9df7 | !locked_p & v8856cb;
assign v85d820 = hready_p & v8822f3 | !hready_p & v8b9e19;
assign v882345 = hready & v85b9f7 | !hready & v845800;
assign v8b9e11 = start_p & v845810 | !start_p & !v857e81;
assign v88234f = hlock1_p & v85a4b1 | !hlock1_p & v845800;
assign v852bf7 = locked_p & v8b9e7b | !locked_p & v845800;
assign v861acc = stateG10_1_p & v85f5b2 | !stateG10_1_p & !v864990;
assign v864e1f = hbusreq1_p & v8b9ea9 | !hbusreq1_p & v88236f;
assign v85ee66 = hready_p & v853612 | !hready_p & v845800;
assign v85330e = hgrant1_p & v8b9f21 | !hgrant1_p & !v88a7b1;
assign v88ffd1 = hbusreq1_p & v8b9ed0 | !hbusreq1_p & v8b9dd5;
assign v8b9ef1 = start_p & v84580e | !start_p & v8822e7;
assign v85d6d3 = hready_p & v8822f3 | !hready_p & v85b83a;
assign v85a970 = stateG3_2_p & v845800 | !stateG3_2_p & v86022a;
assign decide = !v8823b4;
assign v8a065b = hburst1 & v8822cc | !hburst1 & v85331f;
assign v8b9e7b = hmastlock_p & v85b113 | !hmastlock_p & !v845800;
assign v882307 = hready_p & v84581a | !hready_p & !v845814;
assign v85f583 = decide_p & v8b9e5f | !decide_p & v8a065d;
assign v895139 = locked_p & v845814 | !locked_p & !v845800;
assign v85a3e3 = decide_p & v8822d4 | !decide_p & v8a05f0;
assign v859d8d = hbusreq1 & v860568 | !hbusreq1 & v88d057;
assign v85cd0c = decide_p & v88d08c | !decide_p & v8b9dcc;
assign v8b9f27 = hbusreq1_p & v85f588 | !hbusreq1_p & v85f5ad;
assign v8b71ab = decide_p & v8554b2 | !decide_p & v8b9ead;
assign v8b9dcf = decide_p & v862e59 | !decide_p & v84581a;
assign v859474 = decide_p & v8505a9 | !decide_p & v85ae93;
assign v8afeef = stateA1_p & v845800 | !stateA1_p & !v86170f;
assign v895134 = hready_p & v88a7b5 | !hready_p & v88ffcf;
assign v8b9f3b = hready_p & v85f907 | !hready_p & v85791c;
assign v85c5ce = stateG2_p & v845800 | !stateG2_p & v8b9e9b;
assign v8aff0b = locked_p & v856a41 | !locked_p & v845800;
assign v8b9e00 = hburst1_p & v87fd7a | !hburst1_p & v85a031;
assign v85f7a7 = hlock1_p & v88d087 | !hlock1_p & v863a8a;
assign v8b9edf = hmaster0_p & v864e1f | !hmaster0_p & v85029d;
assign v85dfb4 = locked_p & v8b9e17 | !locked_p & v845800;
assign v88d080 = hmastlock_p & v8b9dd8 | !hmastlock_p & v845800;
assign v8530df = hbusreq0 & v8822fe | !hbusreq0 & v845800;
assign v8afefc = hlock0_p & v88d087 | !hlock0_p & v863a8a;
assign v8583bf = locked_p & v845800 | !locked_p & v882332;
assign v85a031 = stateG3_2_p & v845800 | !stateG3_2_p & v87fd7a;
assign v89513a = hbusreq1 & v864525 | !hbusreq1 & v8b9ee7;
assign v887069 = hmaster0_p & v859d97 | !hmaster0_p & v85bab4;
assign v8a05fe = decide_p & v8698e6 | !decide_p & v895151;
assign v8822da = decide_p & v8822f4 | !decide_p & !v852ef0;
assign v85803c = hlock0_p & v8a05fa | !hlock0_p & v88d08c;
assign v8b9e21 = hmaster0_p & v845800 | !hmaster0_p & v85934d;
assign v882304 = decide_p & v85d9d7 | !decide_p & v84581a;
assign v8b71aa = start_p & v85598d | !start_p & v8b9de1;
assign v8822cc = stateA1_p & v845800 | !stateA1_p & !v8b9e32;
assign v8a0602 = locked_p & v87fd78 | !locked_p & v845800;
assign v862c91 = hgrant1_p & v88a7bd | !hgrant1_p & v85ad75;
assign v8856df = hmastlock_p & v85fb94 | !hmastlock_p & v845800;
assign v864990 = hbusreq0_p & v8b9db6 | !hbusreq0_p & v8856ca;
assign v8523bf = locked_p & v85ff2e | !locked_p & v845800;
assign v855d31 = locked_p & v845800 | !locked_p & !v858df2;
assign v860b53 = decide_p & v845808 | !decide_p & v845800;
assign v8b9de7 = hmastlock_p & v85ca1b | !hmastlock_p & !v845800;
assign v857751 = hbusreq1 & v8b9ea4 | !hbusreq1 & v845800;
assign v85b2d4 = start_p & v845800 | !start_p & v85a3f3;
assign hmastlock = v8b71b0;
assign v88d090 = jx1_p & v8b9e5c | !jx1_p & v885719;
assign v855817 = stateA1_p & v8b9da5 | !stateA1_p & v863070;
assign v8b9e0e = hbusreq0_p & v855cc1 | !hbusreq0_p & v858d97;
assign stateG10_1 = !v8a0282;
assign v8b9eb8 = locked_p & v8afeef | !locked_p & v882343;
assign v882316 = stateA1_p & v8b9da5 | !stateA1_p & !v86195f;
assign v8551f3 = hmaster0_p & v8b9efe | !hmaster0_p & v862d65;
assign v85e30c = hready_p & v8b9dba | !hready_p & v858525;
assign v86216f = hgrant1_p & v845804 | !hgrant1_p & !v845800;
assign v88d06e = hready_p & v845800 | !hready_p & v8b9e19;
assign v88d044 = hready_p & v84581a | !hready_p & !v8b9e74;
assign v85e54f = hburst1_p & v845800 | !hburst1_p & !v882340;
assign v85e2a8 = hbusreq0_p & v862224 | !hbusreq0_p & !v8822da;
assign v8b9e8b = hbusreq0_p & v8a0649 | !hbusreq0_p & v845800;
assign v85f5ba = stateG3_1_p & v845800 | !stateG3_1_p & v845826;
assign v85add4 = locked_p & v845800 | !locked_p & !v85f599;
assign v86170f = start_p & v845800 | !start_p & v85cd0b;
assign v8856cf = stateG10_1_p & v850b73 | !stateG10_1_p & v8b9f77;
assign v8b9e20 = hbusreq0 & v8b9dc6 | !hbusreq0 & v862a20;
assign v862ee4 = locked_p & v87fd83 | !locked_p & v85f58b;
assign v8b9dd5 = hgrant1_p & v862e32 | !hgrant1_p & v845800;
assign stateG3_2 = !v885722;
assign v882282 = hbusreq0_p & v8629ac | !hbusreq0_p & v8b9f57;
assign v856316 = hmastlock_p & v8612af | !hmastlock_p & v85f5a3;
assign v85c75d = hmastlock_p & v85dedf | !hmastlock_p & v845800;
assign v8b9ec7 = hmastlock_p & v8a065b | !hmastlock_p & v85331f;
assign v853612 = hmastlock_p & v8822d2 | !hmastlock_p & v845800;
assign v85c974 = hready & v8b9f13 | !hready & v853308;
assign v85a3c2 = decide_p & v8b9e2a | !decide_p & v8aff10;
assign v862ad8 = hready_p & v85a595 | !hready_p & v8a064b;
assign v88ffba = hready & v8b9dee | !hready & v8822c2;
assign v8b9e52 = hbusreq0_p & v853997 | !hbusreq0_p & v85e71f;
assign v8b9dc5 = hready_p & v845800 | !hready_p & !v8a0615;
assign v859d97 = hbusreq1_p & v8b9f14 | !hbusreq1_p & !v863eb5;
assign v88a7c9 = hlock1_p & v8b9e49 | !hlock1_p & v845800;
assign v88d062 = decide_p & v85f596 | !decide_p & v8b9ead;
assign v885713 = hlock0_p & v85a4b1 | !hlock0_p & v845800;
assign v885c4f = start_p & v845800 | !start_p & v864cae;
assign v855460 = hlock0_p & v8b9db3 | !hlock0_p & !v845800;
assign v85d087 = hburst1_p & v85a970 | !hburst1_p & !v845800;
assign v88a7b1 = hbusreq0_p & v887054 | !hbusreq0_p & v858d97;
assign v88d07b = hmastlock_p & v85ef57 | !hmastlock_p & v845800;
assign v8b9f18 = decide_p & v85d667 | !decide_p & v8b9e72;
assign v88228b = stateA1_p & v88705a | !stateA1_p & !v852fbe;
assign v853997 = decide_p & v8b9f60 | !decide_p & !v84581a;
assign v8b9e0f = hlock0_p & v854a42 | !hlock0_p & !v8856cb;
assign v85e315 = hmastlock_p & v858dca | !hmastlock_p & v845800;
assign v895133 = hgrant1_p & v8822ff | !hgrant1_p & !v858af8;
assign v8822d2 = stateA1_p & v845816 | !stateA1_p & v845800;
assign v85f6f8 = hmaster0_p & v8a0640 | !hmaster0_p & v8856e0;
assign v8856e0 = hbusreq1_p & v85f582 | !hbusreq1_p & !v88230b;
assign v85f588 = hgrant1_p & v8578f2 | !hgrant1_p & v88705c;
assign v895152 = stateA1_p & v8822ef | !stateA1_p & v85af59;
assign v88231f = hmastlock_p & v88d07c | !hmastlock_p & v845800;
assign v882344 = hburst1_p & v882340 | !hburst1_p & !v845800;
assign v8b9f90 = hgrant1_p & v8b9e8b | !hgrant1_p & v845800;
assign v8822a3 = hlock1_p & v8822f4 | !hlock1_p & v845800;
assign v856e69 = hgrant1_p & v8a05fe | !hgrant1_p & v8b9f77;
assign v85880f = hbusreq0_p & v882370 | !hbusreq0_p & v8a0623;
assign v88ffc8 = decide_p & v85bc42 | !decide_p & !v85f58f;
assign v8a0606 = decide_p & v88234f | !decide_p & v8b9f3b;
assign v8533a0 = hlock0_p & v854a42 | !hlock0_p & v858df2;
assign v8b9dbf = hlock1_p & v85e30c | !hlock1_p & v845800;
assign v863bff = stateA1_p & v8b9ec8 | !stateA1_p & v863070;
assign v88ffc2 = stateA1_p & v85e25a | !stateA1_p & v85af59;
assign v88ffd0 = stateA1_p & v845800 | !stateA1_p & !v86192f;
assign v852ef0 = hready_p & v84581a | !hready_p & !v89a6f2;
assign v858dca = stateA1_p & v845800 | !stateA1_p & !v8b9ec8;
assign v85f5a3 = hburst0 & v8612af | !hburst0 & !v845800;
assign v86031b = locked_p & v882355 | !locked_p & v845800;
assign v882390 = hgrant1_p & v8b9e1e | !hgrant1_p & v8647b7;
assign v853cf6 = hready_p & v8aff0f | !hready_p & v887053;
assign v85a595 = hbusreq1 & v882351 | !hbusreq1 & v845800;
assign v88705d = hmastlock_p & v8afee6 | !hmastlock_p & v845800;
assign v8b9e59 = decide_p & v853612 | !decide_p & v8a05f0;
assign v8aff0a = hgrant1_p & v845800 | !hgrant1_p & !v845804;
assign v8a0618 = hready_p & v8822fa | !hready_p & v89513a;
assign v852578 = hmaster0_p & v845800 | !hmaster0_p & !v84580a;
assign v8a0640 = hbusreq1_p & v862c91 | !hbusreq1_p & !v8b9e66;
assign v85f5c3 = hready_p & v85dfb4 | !hready_p & v8856cb;
assign v8b9f34 = hready_p & v8508b4 | !hready_p & v8b71a5;
assign v88706c = stateA1_p & v85f1f2 | !stateA1_p & v88239e;
assign v8b9ec8 = start_p & v84580e | !start_p & v85a970;
assign v8b9e22 = hmaster0_p & v859d97 | !hmaster0_p & v8856e0;
assign v8b9df4 = decide_p & v8b9dbd | !decide_p & v845800;
assign v84580b = hbusreq1 & v845800 | !hbusreq1 & !v845800;
assign v85b5d3 = hlock0_p & v850ce7 | !hlock0_p & v8b9e1c;
assign v85fec2 = locked_p & v8822d2 | !locked_p & v845800;
assign v85bab4 = hbusreq1_p & v88d08e | !hbusreq1_p & !v88230b;
assign v88d066 = hready & v8afef9 | !hready & v845800;
assign v845816 = start_p & v845800 | !start_p & !v845800;
assign v88d046 = decide_p & v8afefc | !decide_p & v8a05f1;
assign v8b9dfc = hmastlock_p & v85f5af | !hmastlock_p & !v845800;
assign v88d08c = hlock1_p & v863615 | !hlock1_p & v8b9f20;
assign v85f1f3 = decide_p & v86997d | !decide_p & v845800;
assign v861d53 = hbusreq0 & v85c4a2 | !hbusreq0 & !v845800;
assign v88d088 = stateA1_p & v845816 | !stateA1_p & v850cb2;
assign v8b9dee = hmastlock_p & v862f60 | !hmastlock_p & v845800;
assign v852475 = hbusreq0_p & v88d046 | !hbusreq0_p & v85d0f7;
assign v85ae93 = locked_p & v853612 | !locked_p & v845800;
assign v853647 = hlock0_p & v845800 | !hlock0_p & v8b9e5f;
assign v8822e7 = hburst0_p & v87fd7a | !hburst0_p & v8b9e12;
assign v8856ca = decide_p & v8856cb | !decide_p & v853cf6;
assign v8b9f13 = locked_p & v88237f | !locked_p & v845800;
assign v8822cd = locked_p & v88d05f | !locked_p & v8518b8;
assign v88d056 = decide_p & v8822b1 | !decide_p & !v84581a;
assign v88230c = hlock0_p & v8b9e72 | !hlock0_p & v85d667;
assign v860b2a = stateG2_p & v845800 | !stateG2_p & v882340;
assign v8578ef = hmastlock_p & v882365 | !hmastlock_p & v845800;
assign v88705e = hbusreq1 & v8628b1 | !hbusreq1 & !v845800;
assign v853437 = hbusreq1 & v8b9f69 | !hbusreq1 & !v8822cf;
assign v8822ef = start_p & v85598d | !start_p & v8b9f17;
assign v8b9f06 = hburst0_p & v882340 | !hburst0_p & v882344;
assign stateG3_0 = !v88a7ca;
assign v85bc9e = hgrant1_p & v861ed5 | !hgrant1_p & v8b9e56;
assign v8b9de4 = hready_p & v88705e | !hready_p & v858891;
assign v88a7b4 = hlock0_p & v88d06e | !hlock0_p & v845800;
assign v8a060b = hready_p & v8aff10 | !hready_p & v88d07b;
assign v845824 = stateG2_p & v845800 | !stateG2_p & !v845800;
assign v8b71ac = hlock0_p & v8856da | !hlock0_p & v845800;
assign v85abe0 = decide_p & v858a13 | !decide_p & v864941;
assign v862e72 = start_p & v85cd0b | !start_p & v845800;
assign v88233e = hburst0 & v8b9f35 | !hburst0 & v845800;
assign v8b71b0 = hmaster0_p & v8b9f26 | !hmaster0_p & v853cad;
assign v861f20 = hbusreq0_p & v8b9ea8 | !hbusreq0_p & v88228e;
assign v862f33 = decide_p & v88237e | !decide_p & !v8b9de4;
assign v85fa6a = hready_p & v8523bf | !hready_p & v858525;
assign v8b9ea4 = hbusreq0 & v8822e2 | !hbusreq0 & v8823a4;
assign v856019 = hbusreq0_p & v85a3e3 | !hbusreq0_p & v8b9e59;
assign v85cc6b = hgrant1_p & v861f20 | !hgrant1_p & !v85c3b7;
assign v85f596 = hready_p & v8b9ead | !hready_p & v85f58b;
assign v85c59b = hbusreq0_p & v882399 | !hbusreq0_p & v8b9f18;
assign v8628dd = hmastlock_p & v8b9e50 | !hmastlock_p & !v845800;
assign v8856dd = hlock0_p & v8b9f4c | !hlock0_p & v845800;
assign v88236f = hgrant1_p & v88231d | !hgrant1_p & !v845800;
assign hmaster0 = v893788;
assign v860719 = hgrant1_p & v882376 | !hgrant1_p & v856019;
assign v8b9e2c = hmastlock_p & v8520a6 | !hmastlock_p & !v845800;
assign v8b9ee7 = hbusreq0 & v89a6f1 | !hbusreq0 & v845800;
assign v85e961 = hgrant1_p & v8a0623 | !hgrant1_p & v845800;
assign v85de6c = hready_p & v84580b | !hready_p & v845807;
assign v85465f = hgrant1_p & v8b9dd1 | !hgrant1_p & v8b9ef5;
assign v85b6dd = hgrant1_p & v8b9dd1 | !hgrant1_p & v85e2a8;
assign v88238f = hbusreq0_p & v8b9e04 | !hbusreq0_p & v85f5b1;
assign v853308 = locked_p & v8b9e2f | !locked_p & v845800;
assign v8a0653 = hburst0_p & v85a970 | !hburst0_p & v85d087;
assign v84580a = hbusreq1_p & v845800 | !hbusreq1_p & !v845800;
assign v8822c2 = hmastlock_p & v8822cc | !hmastlock_p & !v84580f;
assign v8b9e57 = hlock1_p & v882348 | !hlock1_p & v845800;
assign v8523de = hlock0_p & v859006 | !hlock0_p & v845800;
assign v8aff05 = hburst1_p & v845800 | !hburst1_p & !v85a970;
assign v85f589 = hgrant1_p & v861ed5 | !hgrant1_p & v85cbe8;
assign v8508b4 = hbusreq1 & v8b9dc7 | !hbusreq1 & !v85f5ac;
assign v882373 = hgrant1_p & v859474 | !hgrant1_p & v8607e4;
assign v87fd78 = hmastlock_p & v88d085 | !hmastlock_p & v857e7d;
assign v88ffd5 = hmaster0_p & v88ffd1 | !hmaster0_p & v85a8a7;
assign v8b9deb = hbusreq0_p & v85f5c3 | !hbusreq0_p & v861ed5;
assign v8b9ddc = hlock1_p & v859575 | !hlock1_p & !v857768;
assign v85f58d = hmastlock_p & v88ffc2 | !hmastlock_p & !v845800;
assign v863d0e = start_p & v845800 | !start_p & v8aff00;
assign v850b73 = hbusreq0_p & v85b4d5 | !hbusreq0_p & v88237d;
assign v8822f3 = locked_p & v88231f | !locked_p & v845800;
assign v8b9e5f = hready_p & v845800 | !hready_p & !v858df2;
assign v85f5ad = hgrant1_p & v85d0f7 | !hgrant1_p & !v895132;
assign v885700 = start_p & v84580e | !start_p & v85596e;
assign v85c62e = locked_p & v85e315 | !locked_p & !v845800;
assign v88a7a3 = hlock1 & v882326 | !hlock1 & v8b9f51;
assign v864525 = hbusreq0 & v8afefa | !hbusreq0 & v845800;
assign stateG2 = !v88ffd5;
assign v8b9e28 = hbusreq1_p & v895133 | !hbusreq1_p & !v8612b9;
assign v88231d = hbusreq0_p & v860b53 | !hbusreq0_p & !v845818;
assign v85f1ae = hready & v8b9eb2 | !hready & v85e4e6;
assign v86195f = start_p & v845810 | !start_p & v845800;
assign v85f5b7 = start_p & v84580e | !start_p & v87fd7a;
assign v8612b9 = hgrant1_p & v8a05fe | !hgrant1_p & v8856cf;
assign v88706f = jx1_p & v8618bd | !jx1_p & v862090;
assign v857fb9 = hbusreq1_p & v864244 | !hbusreq1_p & v8822ad;
assign v895157 = hmaster0_p & v8620e6 | !hmaster0_p & v8b9dc4;
assign v8a0639 = start_p & v845810 | !start_p & !v852edf;
assign v882381 = hready_p & v85f6d6 | !hready_p & v85bae3;
assign v860967 = stateG2_p & v845800 | !stateG2_p & v85a970;
assign v857eeb = decide_p & v845800 | !decide_p & v88ffbd;
assign v8631cf = hmastlock_p & v8822cc | !hmastlock_p & v845800;
assign v8b9f0a = hmaster0_p & v8b9f56 | !hmaster0_p & v859ca9;
assign v86042c = hlock1_p & v8b9dc5 | !hlock1_p & v85323a;
assign v8afeed = start_p & v84580e | !start_p & v86022a;
assign v88237e = hlock1_p & v8b9ed7 | !hlock1_p & v845800;
assign v8b71ad = hmastlock_p & v861fa1 | !hmastlock_p & !v845800;
assign v882305 = hburst0_p & v845800 | !hburst0_p & v8aff05;
assign v8b9eed = hlock1_p & v85f67e | !hlock1_p & !v845800;
assign v845814 = hmastlock_p & v845800 | !hmastlock_p & !v845800;
assign v8822be = decide_p & v858df5 | !decide_p & v845800;
assign v85cb98 = hbusreq0_p & v8a05f8 | !hbusreq0_p & v858d97;
assign v8b9ed5 = hbusreq0_p & v85f5bf | !hbusreq0_p & v8a061b;
assign v8b9efd = jx0_p & v88ffbb | !jx0_p & v864246;
assign v8afef9 = locked_p & v8631cf | !locked_p & v8b9e74;
assign v85b113 = stateA1_p & v85f5b7 | !stateA1_p & v885702;
assign v882317 = hready & v862ee4 | !hready & v8822cd;
assign stateA1 = v85f5c7;
assign v85d0f1 = hbusreq0_p & v8b9fa2 | !hbusreq0_p & v845800;
assign v8b9e1c = hready_p & v84581a | !hready_p & !v845800;
assign v85e920 = hmastlock_p & v88234d | !hmastlock_p & v845800;
assign v88230b = hgrant1_p & v8b9e52 | !hgrant1_p & !v882349;
assign v8539e6 = hmastlock_p & v8b9da5 | !hmastlock_p & v845800;
assign v8b9e51 = hlock0_p & v8b9db3 | !hlock0_p & v845800;
assign v850c63 = hlock1_p & v8b9ddd | !hlock1_p & v845800;
assign v85f581 = locked_p & v88d080 | !locked_p & v845800;
assign v8b9dba = locked_p & v856316 | !locked_p & v845800;
assign v8856d5 = hbusreq0 & v861c42 | !hbusreq0 & !v8619fc;
assign v88232a = decide_p & v8b9ed6 | !decide_p & v845800;
assign v8b9ea7 = stateA1_p & v8b9ec8 | !stateA1_p & v8b9e32;
assign v864711 = hgrant1_p & v8b9e4b | !hgrant1_p & v88d071;
assign v8b9dc2 = hlock0_p & v882363 | !hlock0_p & !v85bc42;
assign v882340 = stateG3_2_p & v845800 | !stateG3_2_p & !v85f5ba;
assign v88d069 = stateG2_p & v84582a | !stateG2_p & v85a970;
assign v852c3b = hbusreq0_p & v88d04d | !hbusreq0_p & v8b9dcf;
assign v8b9e9f = hbusreq1_p & v8b9e1b | !hbusreq1_p & v8856c9;
assign v8633f4 = hlock1_p & v8b9dd1 | !hlock1_p & !v8822f4;
assign v8b9dd8 = stateA1_p & v88239e | !stateA1_p & !v852fbe;
assign v85263d = hburst1 & v8b9f35 | !hburst1 & v88233e;
assign v8617ee = start_p & v85598d | !start_p & v882340;
assign v845806 = hbusreq0_p & v845800 | !hbusreq0_p & !v845800;
assign v858a13 = hready_p & v845800 | !hready_p & v8856cb;
assign v88ffcf = hbusreq1 & v8b9f48 | !hbusreq1 & v845800;
assign v882310 = decide_p & v8b9e0f | !decide_p & !v855d31;
assign v855784 = jx0_p & v864246 | !jx0_p & v85e3ad;
assign v8b9efe = hbusreq1_p & v8579d6 | !hbusreq1_p & v85f589;
assign v85c7fb = stateG2_p & v845800 | !stateG2_p & v8b9de1;
assign v8afee8 = hbusreq0_p & v8b9e92 | !hbusreq0_p & v85f583;
assign v85323a = hready_p & v845800 | !hready_p & v8822bb;
assign v85cb5c = hgrant1_p & v85d0f7 | !hgrant1_p & !v861acc;
assign v8b9f21 = hbusreq0_p & v88a7bc | !hbusreq0_p & v8a061b;
assign v85877f = hmaster0_p & v85f1d9 | !hmaster0_p & v862d65;
assign v8b9e97 = hbusreq1 & v8822fe | !hbusreq1 & v845800;
assign v882338 = decide_p & v8571d1 | !decide_p & v845800;
assign v8823a5 = hready_p & v85bc80 | !hready_p & v8856cb;
assign v85b9f7 = locked_p & v85e920 | !locked_p & v845800;
assign v8612af = stateA1_p & v88d085 | !stateA1_p & v8b9ec8;
assign v887054 = decide_p & v855d10 | !decide_p & v845800;
assign v8520a6 = stateA1_p & v8822ef | !stateA1_p & v885702;
assign v85fe4d = hlock1_p & v89a6f4 | !hlock1_p & v85f67e;
assign v862e32 = decide_p & v845800 | !decide_p & v8822c3;
assign v882285 = locked_p & v85f5c1 | !locked_p & !v845800;
assign v8b9f51 = hready & v8631cf | !hready & v8b9f35;
assign v8b9f03 = hready & v85f5c2 | !hready & v8b9e6c;
assign v8b9dcd = hlock1_p & v862ad8 | !hlock1_p & v88d06f;
assign v8607e4 = decide_p & v86223c | !decide_p & v845800;
assign v845826 = stateG3_0_p & v845800 | !stateG3_0_p & !v845800;
assign v8a0649 = decide_p & v8523de | !decide_p & !v88a7aa;
assign v88d05e = hbusreq0_p & v8822be | !hbusreq0_p & v8a061b;
assign v862097 = hlock1_p & v8b9e72 | !hlock1_p & v85d667;
assign v855cc1 = decide_p & v856d8f | !decide_p & v845800;
assign v85315d = hlock0_p & v84580c | !hlock0_p & v862e59;
assign v85cbe8 = stateG10_1_p & v8531a0 | !stateG10_1_p & v8b9e56;
assign v8afef1 = hbusreq1_p & v851b5f | !hbusreq1_p & v864cfd;
assign v8637b3 = hbusreq0_p & v8612ae | !hbusreq0_p & v885718;
assign v85c750 = hlock1 & v887062 | !hlock1 & v85f81e;
assign v87fd86 = hmaster0_p & v8b9e9f | !hmaster0_p & !v8afef6;
assign v85f58b = hmastlock_p & v8b9e9a | !hmastlock_p & v845800;
assign v8b9e9a = stateA1_p & v845800 | !stateA1_p & v86170f;
assign v882326 = hready & v8578ef | !hready & !v845800;
assign v860fbc = stateA1_p & v85e25a | !stateA1_p & v86192f;
assign v882291 = hmastlock_p & v882354 | !hmastlock_p & v845800;
assign v8823b4 = jx1_p & v85f57e | !jx1_p & v845800;
assign v88ffc0 = stateA1_p & v845800 | !stateA1_p & !v8b9ef1;
assign v858df5 = hlock0_p & v845800 | !hlock0_p & v8b9dd1;
assign v87fd7a = stateG3_1_p & v845800 | !stateG3_1_p & !v845826;
assign v85d9d7 = hlock0_p & v8b9f64 | !hlock0_p & !v845800;
assign v86028b = start_p & v845810 | !start_p & !v845824;
assign v8a065c = hlock1_p & v845800 | !hlock1_p & !v8856f0;
assign v8a0609 = hmastlock_p & v8612af | !hmastlock_p & !v845800;
assign v88d05f = hmastlock_p & v88229f | !hmastlock_p & !v845800;
assign v8822c1 = hlock0_p & v8b9e1c | !hlock0_p & !v8822f4;
assign v860c97 = hbusreq0_p & v8b9e30 | !hbusreq0_p & v862e32;
assign busreq = v89a6f5;
assign v8b9f8f = hready_p & v8b9df7 | !hready_p & v845800;
assign v85f141 = hbusreq0_p & v882310 | !hbusreq0_p & !v8b9e26;
assign v85654f = hgrant1_p & v8822d5 | !hgrant1_p & !v845800;
assign v856a41 = hmastlock_p & v856c47 | !hmastlock_p & v845800;
assign v8a0648 = start_p & v85cd0b | !start_p & !v8b9de6;
assign v85c7f3 = hmaster0_p & v85215e | !hmaster0_p & v864711;
assign v85ca1b = stateA1_p & v8822ef | !stateA1_p & !v8a0639;
assign v85ff2e = hmastlock_p & v8612af | !hmastlock_p & v857e7d;
assign v859ca9 = hbusreq1_p & v8545f6 | !hbusreq1_p & v85e753;
assign v8b71a8 = hlock1_p & v8b9db3 | !hlock1_p & !v845800;
assign v85f58e = decide_p & v8b9f5d | !decide_p & v85d6d3;
assign v8b9ed6 = hlock0_p & v8b9ddd | !hlock0_p & v845800;
assign v8aff00 = stateG3_2_p & v845800 | !stateG3_2_p & v85e4a1;
assign v88d04d = decide_p & v85315d | !decide_p & v84581a;
assign v85f1f2 = start_p & v84580e | !start_p & v85cb28;
assign v8822e3 = hlock0_p & v8b9ddc | !hlock0_p & v862346;
assign v895135 = hlock0_p & v882348 | !hlock0_p & v845800;
assign v882376 = decide_p & v8606fb | !decide_p & v85ae93;
assign v8619fc = hready & v859035 | !hready & v88a7c6;
assign v863a8a = hready_p & v88d040 | !hready_p & v8856cb;
assign v8b9f26 = hbusreq1_p & v85b6dd | !hbusreq1_p & v85465f;
assign v86022a = stateG3_1_p & v845826 | !stateG3_1_p & !v845826;
assign v8b9db3 = hready_p & v85add4 | !hready_p & v845814;
assign v85adda = hbusreq0_p & v88232a | !hbusreq0_p & v845800;
assign v850cb2 = start_p & v845800 | !start_p & !v84582a;
assign v85a414 = start_p & v845810 | !start_p & !v88d073;
assign v8b9e4b = hbusreq0_p & v864411 | !hbusreq0_p & v8b9e59;
assign v88237f = hmastlock_p & v863bff | !hmastlock_p & !v845800;
assign v8b9f69 = hbusreq0 & v88a7ba | !hbusreq0 & v861063;
assign v8823a4 = hlock1 & v8b9e85 | !hlock1 & !v864183;
assign v882363 = hlock1_p & v859575 | !hlock1_p & v862346;
assign v8b9ef0 = start_p & v845810 | !start_p & v882305;
assign v882351 = hbusreq0 & v862f88 | !hbusreq0 & !v85c750;
assign v8b9e1d = hmastlock_p & v8a065b | !hmastlock_p & !v8b9f4d;
assign v864244 = hgrant1_p & v85f58e | !hgrant1_p & v882338;
assign v85f1d9 = hbusreq1_p & v8579d6 | !hbusreq1_p & v85bc9e;
assign v8b9e56 = hbusreq0_p & v85ff1e | !hbusreq0_p & v85abe0;
assign v8b9f44 = hburst1_p & v859163 | !hburst1_p & v845800;
assign v8b71ae = hgrant1_p & v84580b | !hgrant1_p & v88d051;
assign v861ed5 = decide_p & v8823a5 | !decide_p & v85d0b4;
assign v8626cc = stateA1_p & v88239e | !stateA1_p & !v845800;
assign v851b6e = hmaster0_p & v845806 | !hmaster0_p & !v845800;
assign v84581e = hgrant1_p & v845800 | !hgrant1_p & !v845800;
assign v8579d6 = hgrant1_p & v85f5c3 | !hgrant1_p & v85abe0;
assign v87fd83 = hmastlock_p & v860fbc | !hmastlock_p & !v845800;
assign v8b9dbd = hlock0_p & v8822f4 | !hlock0_p & !v845800;
assign v85a3f3 = stateG2_p & v845800 | !stateG2_p & v859163;
assign v8597ea = hready_p & v845800 | !hready_p & v858525;
assign v85f582 = hgrant1_p & v882342 | !hgrant1_p & v851c6c;
assign v84582a = stateG3_2_p & v845800 | !stateG3_2_p & !v845800;
assign v85596e = stateG2_p & v84582a | !stateG2_p & v85a031;
assign v858af8 = hbusreq0_p & v8823ab | !hbusreq0_p & !v88ffc8;
assign v862224 = decide_p & v863af6 | !decide_p & v852ef0;
assign v8b9e2f = hmastlock_p & v88228b | !hmastlock_p & v845800;
assign v8628b1 = hbusreq0 & v882317 | !hbusreq0 & v8b9f03;
assign v8856c9 = hgrant1_p & v8b9f18 | !hgrant1_p & !v845804;
assign v8545f6 = hgrant1_p & v8637b3 | !hgrant1_p & !v85f5b3;
assign v885718 = decide_p & v8b9e1c | !decide_p & v845800;
assign v8631b2 = hready_p & v8539e3 | !hready_p & v8a0615;
assign v88a7ca = hmaster0_p & v857fb9 | !hmaster0_p & v882390;
assign v857e7d = hburst0 & v8822d8 | !hburst0 & !v845800;
assign v861546 = jx0_p & v85877f | !jx0_p & v8551f3;
assign v85923c = hlock1_p & v87fd84 | !hlock1_p & v845800;
assign v88234d = stateA1_p & v845800 | !stateA1_p & v885c4f;
assign v856288 = stateA1_p & v88238a | !stateA1_p & v8b9e47;
assign v8a0641 = decide_p & v855460 | !decide_p & v845800;
assign v85ca17 = hlock0_p & v85ce61 | !hlock0_p & !v8632bb;
assign v88235a = hbusreq1 & v861d53 | !hbusreq1 & v860f3e;
assign v860fce = hbusreq0_p & v8629ac | !hbusreq0_p & v8856ca;
assign v88d07d = stateA1_p & v8afeed | !stateA1_p & !v845800;
assign v8b9ed0 = hgrant1_p & v85a3c2 | !hgrant1_p & v882328;
assign v845805 = hready & v845800 | !hready & !v845800;
assign v89a6f5 = hmaster0_p & v8b71ae | !hmaster0_p & v8b9e67;
assign v8b9f4f = hready & v8afee2 | !hready & v845800;
assign v86314b = hbusreq0_p & v859134 | !hbusreq0_p & v845800;
assign v885c50 = decide_p & v882332 | !decide_p & v8583bf;
assign v860625 = hlock1_p & v89513e | !hlock1_p & v845800;
assign v85e3ad = hmaster0_p & v8b9e28 | !hmaster0_p & !v85e7b1;
assign v85e7e0 = hlock0_p & v8b9f8f | !hlock0_p & v8856cb;
assign v88d070 = hgrant1_p & v8822da | !hgrant1_p & !v8b9dd1;
assign v8b9e46 = decide_p & v8b71a8 | !decide_p & v845800;
assign v845804 = hready_p & v845800 | !hready_p & !v845800;
assign v8b9dca = decide_p & v858df2 | !decide_p & !v855d31;
assign v863af6 = hlock0_p & v8b9dd1 | !hlock0_p & !v8822f4;
assign v85f5ac = hbusreq0 & v8b9f6c | !hbusreq0 & !v845800;
assign v8b9dce = hmaster0_p & v8b9da6 | !hmaster0_p & v8afef1;
assign v85cb28 = stateG2_p & v84582a | !stateG2_p & v882340;
assign v882325 = hmastlock_p & v88d07d | !hmastlock_p & !v845800;
assign v882328 = decide_p & v8b9e57 | !decide_p & v845800;
assign v8b9f81 = hlock0_p & v845800 | !hlock0_p & v858a13;
assign v88d077 = decide_p & v8822e3 | !decide_p & v85f58f;
assign v88a7ba = hlock1 & v88a7b7 | !hlock1 & v8afefe;
assign v882395 = hready_p & v8aff0f | !hready_p & v8856cb;
assign v8b9e72 = hready_p & v895139 | !hready_p & v845800;
assign v858d97 = decide_p & v8822f4 | !decide_p & v845800;
assign v882382 = jx0_p & v85e7fa | !jx0_p & !v845800;
assign v85bc42 = hlock1_p & v857768 | !hlock1_p & v882343;
assign v8b9dd1 = hready_p & v84581a | !hready_p & v845814;
assign v8b9f80 = stateA1_p & v88d085 | !stateA1_p & !v845800;
assign v85ef57 = stateA1_p & v89514a | !stateA1_p & v862e72;
assign v8822d8 = start_p & v84580e | !start_p & v845800;
assign v88a7a9 = decide_p & v845808 | !decide_p & v84581a;
assign v88d061 = hlock1 & v88229d | !hlock1 & v84581a;
assign v8b9dc1 = hlock0_p & v8b9f09 | !hlock0_p & v8856cb;
assign v8b9de6 = stateG2_p & v845800 | !stateG2_p & v8b9e25;
assign v8b9f6e = decide_p & v8822a3 | !decide_p & !v84581a;
assign v8b9e35 = hmastlock_p & v8b71aa | !hmastlock_p & v845800;
assign v88228d = hlock0_p & v8b9dc3 | !hlock0_p & !v8b9dbf;
assign v8b9dbb = hbusreq0 & v8b9e34 | !hbusreq0 & !v845800;
assign v86482d = hburst1_p & v845828 | !hburst1_p & v85a031;
assign v8856d4 = hready_p & v853437 | !hready_p & v88230e;
assign v85e25a = start_p & v84580e | !start_p & v85a031;
assign v8b9e50 = stateA1_p & v845800 | !stateA1_p & v84582a;
assign v882306 = stateA1_p & v8b9da5 | !stateA1_p & !v85a414;
assign v88239e = start_p & v84580e | !start_p & v882340;
assign v855bfd = hmastlock_p & v8b9f39 | !hmastlock_p & v845800;
assign v88d076 = decide_p & v85c9ad | !decide_p & v84581a;
assign v8b9ea8 = decide_p & v8822c6 | !decide_p & v845800;
assign v85f59a = hready_p & v845800 | !hready_p & v853612;
assign v857768 = hready_p & v882343 | !hready_p & v8a0613;
assign v88ffc1 = hlock0_p & v860c3a | !hlock0_p & v863d44;
assign v85736e = decide_p & v8533a0 | !decide_p & !v855d31;
assign v8b9e9b = stateG3_2_p & v845800 | !stateG3_2_p & !v845828;
assign v8822e2 = hlock1 & v882345 | !hlock1 & !v88231a;
assign v85ce69 = hlock1_p & v8597ea | !hlock1_p & v845800;
assign v8a0620 = hbusreq0 & v882345 | !hbusreq0 & v845800;
assign v8b9de1 = stateG3_2_p & v845800 | !stateG3_2_p & !v845826;
assign v85c89c = hbusreq1_p & v852071 | !hbusreq1_p & v8b9f90;
assign v859134 = decide_p & v8856dd | !decide_p & v845800;
assign v88705c = decide_p & v862f96 | !decide_p & v858794;
assign v85cd3f = locked_p & v8b71ad | !locked_p & !v845814;
assign v88a7b7 = hready & v8b9f71 | !hready & !v845800;
assign v8b9e47 = start_p & v85cd0b | !start_p & v864cae;
assign v8a0633 = hburst1_p & v8b9e25 | !hburst1_p & !v845800;
assign v87fd84 = hready_p & v845800 | !hready_p & v89513a;
assign v8b9e2a = hlock1_p & v8a060b | !hlock1_p & v845800;
assign v862032 = decide_p & v85ca17 | !decide_p & v84581a;
assign v8afefa = hready & v8856df | !hready & v845800;
assign v85fb02 = start_p & v84580e | !start_p & v85cd0b;
assign v8b9f71 = locked_p & v8822fc | !locked_p & v845800;
assign v8698e6 = hready_p & v85968b | !hready_p & v85f58b;
assign v89514a = start_p & v85cd0b | !start_p & v8b9e90;
assign v8591b7 = decide_p & v85f5b5 | !decide_p & v845800;
assign v86192f = start_p & v84580e | !start_p & v8a05fc;
assign v8569be = decide_p & v8b9e7e | !decide_p & v84581a;
assign v887053 = locked_p & v845800 | !locked_p & v8856cb;
assign v84580c = hlock1_p & v845800 | !hlock1_p & !v845800;
assign v851d36 = stateG3_2_p & v845800 | !stateG3_2_p & v85f5ba;
assign v8b9f3f = hlock1_p & v845804 | !hlock1_p & v8b9e1c;
assign v85f57e = jx0_p & v8b9e21 | !jx0_p & v882391;
assign v864279 = hmastlock_p & v857931 | !hmastlock_p & !v845800;
assign v864183 = hready & v8b9de7 | !hready & v8b9f0e;
assign v858794 = hready_p & v8856cb | !hready_p & v887053;
assign v8b9ef5 = hbusreq0_p & v85d046 | !hbusreq0_p & !v8822da;
assign v863615 = hready_p & v8b9dcc | !hready_p & v8a0613;
assign v85c719 = hgrant1_p & v858768 | !hgrant1_p & v864523;
assign v85d8f3 = hmastlock_p & v8b9ded | !hmastlock_p & v845800;
assign v85c3b7 = hbusreq0_p & v85f1f3 | !hbusreq0_p & v8b9e46;
assign v8b9f6a = decide_p & v8b9e60 | !decide_p & v845800;
assign v85e753 = hgrant1_p & v8a064d | !hgrant1_p & !v845800;
assign v85af59 = start_p & v85598d | !start_p & v85a031;
assign v862f60 = stateA1_p & v845800 | !stateA1_p & v85b585;
assign v887059 = decide_p & v8b9e51 | !decide_p & !v84581a;
assign v8a05f0 = hready_p & v853612 | !hready_p & v8b9f11;
assign v85e4e6 = locked_p & v882325 | !locked_p & v8518b8;
assign v863b11 = hlock1 & v8a0632 | !hlock1 & v8b9f51;
assign v8b9f5d = hlock1_p & v85d820 | !hlock1_p & v845800;
assign v8556fc = hbusreq0 & v8afefa | !hbusreq0 & v8605e3;
assign v85f57f = hmastlock_p & v863070 | !hmastlock_p & v845800;
assign v8b9e90 = stateG2_p & v84582a | !stateG2_p & v845800;
assign v85215e = hbusreq1_p & v882373 | !hbusreq1_p & v860719;
assign v8b9ded = stateA1_p & v845800 | !stateA1_p & v862e72;
assign v85a8a7 = hgrant1_p & v8a062c | !hgrant1_p & v860c97;
assign v845807 = hbusreq0 & v845800 | !hbusreq0 & !v845800;
assign v8b9e31 = decide_p & v862097 | !decide_p & v8b9e72;
assign v8b9dc7 = hbusreq0 & v8b9f4f | !hbusreq0 & v845800;
assign v8822c6 = hlock0_p & v85ac94 | !hlock0_p & v8606e5;
assign v845800 = 1;
assign v85c5b2 = stateA1_p & v8623ae | !stateA1_p & v8617ee;
assign v88d085 = start_p & v84580e | !start_p & v88d069;
assign v88228e = decide_p & v850934 | !decide_p & v845800;
assign v885702 = start_p & v85598d | !start_p & v88d052;
assign v858768 = hbusreq0_p & v85ce00 | !hbusreq0_p & !v88237d;
assign v858cf2 = hmastlock_p & v88ffc0 | !hmastlock_p & v845800;
assign v8b9e8f = hmaster0_p & v8a0630 | !hmaster0_p & v859ca9;
assign v88d08e = hgrant1_p & v88238f | !hgrant1_p & v8b9dff;
assign v89a6f4 = hready_p & v88d061 | !hready_p & v8a0615;
assign v8b9ead = locked_p & v845800 | !locked_p & v85f58b;
assign v845818 = decide_p & v845800 | !decide_p & !v845800;
assign v852fbe = start_p & v845810 | !start_p & v8822c8;
assign v8518b8 = hmastlock_p & v8b9def | !hmastlock_p & v845800;
assign v8b9f58 = locked_p & v8b9f5a | !locked_p & v845800;
assign v8a0615 = hlock1 & v8b9e13 | !hlock1 & v845814;
assign v8822a8 = locked_p & v864279 | !locked_p & !v845800;
assign v85f5c1 = hmastlock_p & v895152 | !hmastlock_p & !v845800;
assign v887066 = hbusreq0_p & v8b9f6a | !hbusreq0_p & v8b9e46;
assign v85f5b2 = hbusreq0_p & v85736e | !hbusreq0_p & v8b9dca;
assign v85af06 = stateG10_1_p & v8afee8 | !stateG10_1_p & v8b9e56;
assign v8a064d = hbusreq0_p & v8b9df4 | !hbusreq0_p & !v845818;
assign v8b9e7e = hlock0_p & v8a065c | !hlock0_p & !v8a0621;
assign v85f58f = locked_p & v845800 | !locked_p & !v882343;
assign v8b9e0b = hbusreq1 & v8556fc | !hbusreq1 & v845800;
assign v882375 = stateG3_2_p & v845800 | !stateG3_2_p & v845828;
assign v860c3a = hlock1_p & v8856d4 | !hlock1_p & v845800;
assign v8b9e26 = decide_p & v8856cb | !decide_p & v855d31;
assign v860568 = hbusreq0 & v85f1ae | !hbusreq0 & !v845800;
assign v85fad3 = hburst0_p & v8b9e25 | !hburst0_p & v8a0633;
assign v8822c4 = locked_p & v845800 | !locked_p & v882343;
assign v854a42 = hready_p & v8628dd | !hready_p & !v845800;
assign v882392 = hlock1 & v851b5e | !hlock1 & v8562e6;
assign v8b9fa4 = stateA1_p & v8a0648 | !stateA1_p & v8822b6;
assign v851b5f = hgrant1_p & v882282 | !hgrant1_p & v852475;
assign v862e59 = hlock1_p & v8b9dd1 | !hlock1_p & !v845800;
assign locked = v8aff12;
assign v8a0611 = hlock0_p & v86042c | !hlock0_p & v8606e5;
assign v8b9dff = hbusreq0_p & v8569be | !hbusreq0_p & !v88d056;
assign v882342 = hbusreq0_p & v8b71a6 | !hbusreq0_p & v860700;
assign v8b9f39 = start_p & v845800 | !start_p & !v851d36;
assign v8b9e30 = decide_p & v882369 | !decide_p & v8aff10;
assign v882349 = hbusreq0_p & v88a7a9 | !hbusreq0_p & !v85e71f;
assign v8a062a = hbusreq0 & v8b9e41 | !hbusreq0 & v845800;
assign v85331f = hburst0 & v8822cc | !hburst0 & v845800;
assign v862857 = hburst1_p & v8b9e25 | !hburst1_p & v85a970;
assign v87fd7f = stateA1_p & v8b9da5 | !stateA1_p & !v8b9ef0;
assign v85f592 = hbusreq0 & v863b11 | !hbusreq0 & !v882392;
assign v8a0623 = decide_p & v845800 | !decide_p & v882381;
assign v8aff10 = locked_p & v88d07b | !locked_p & v845800;
assign v8856d6 = hlock0_p & v88a7c9 | !hlock0_p & v85923c;
assign v85c4a2 = hready & v85cd3f | !hready & v8aff03;
assign v8b9f77 = hbusreq0_p & v8b71ab | !hbusreq0_p & v88237d;
assign v8b9ea9 = hgrant1_p & v88d05e | !hgrant1_p & !v8b9e0e;
assign v85a5c7 = decide_p & v88a7b4 | !decide_p & v845800;
assign v8856cb = hmastlock_p & v850cb2 | !hmastlock_p & v845800;
assign v852a1d = hlock1_p & v8b9dc5 | !hlock1_p & v88d044;
assign v85968b = locked_p & v8b9e9a | !locked_p & v85f58b;
assign v86240b = stateG10_1_p & v8b9e88 | !stateG10_1_p & v8b9f77;
assign v84580f = hburst0 & v845800 | !hburst0 & !v845800;
assign v863070 = start_p & v85598d | !start_p & v85a970;
assign v88a7b5 = hbusreq1 & v8856d5 | !hbusreq1 & v845800;
assign v8554b2 = hlock0_p & v845800 | !hlock0_p & v85f58b;
assign v85d667 = hready_p & v84581a | !hready_p & v845800;
assign v8822b1 = hlock1_p & v8b9db3 | !hlock1_p & v845800;
assign v8b9e1b = hgrant1_p & v8b9e31 | !hgrant1_p & !v845804;
assign v882369 = hlock0_p & v8a060b | !hlock0_p & v845800;
assign v8856f0 = hready_p & v85c572 | !hready_p & v858525;
assign v86223c = hlock1_p & v85f59a | !hlock1_p & v845800;
assign v85f5bf = decide_p & v8b9ee3 | !decide_p & v845800;
assign v8a0610 = decide_p & v8b71ac | !decide_p & v85ae93;
assign v8b9e06 = hgrant1_p & v8a05fe | !hgrant1_p & v86240b;
assign v8b9f64 = hlock1_p & v845800 | !hlock1_p & v8b9dd1;
assign v88d051 = hready_p & v845807 | !hready_p & v84580b;
assign v850ce7 = hlock1_p & v845804 | !hlock1_p & v8822f4;
assign v8a0621 = hlock1_p & v85f67e | !hlock1_p & v845800;
assign v85a9a4 = hbusreq0 & v8562e6 | !hbusreq0 & !v845800;
assign v85d046 = decide_p & v8822c1 | !decide_p & v852ef0;
assign v852071 = hgrant1_p & v85d0f1 | !hgrant1_p & v85fd24;
assign v85f0c6 = locked_p & v88d06d | !locked_p & v845800;
assign v85ce00 = decide_p & v85688b | !decide_p & !v85f58f;
assign v88705a = start_p & v84580e | !start_p & !v85f5ba;
assign v893788 = hmaster0_p & v8aff0a | !hmaster0_p & v86216f;
assign v8b9e25 = stateG3_1_p & v845826 | !stateG3_1_p & !v845800;
assign v8b9e3e = hgrant1_p & v8a0606 | !hgrant1_p & v88229c;
assign v882332 = hmastlock_p & v8b9f40 | !hmastlock_p & v845800;
assign v8afef8 = jx0_p & v85957f | !jx0_p & v85877f;
assign v8b9ddd = hready_p & v845800 | !hready_p & v88705d;
assign v85f5c7 = jx1_p & v855784 | !jx1_p & v8b9efd;
assign v8a05f8 = decide_p & v853c79 | !decide_p & v845800;
assign v8b9ea0 = hready_p & v845800 | !hready_p & v8a064b;
assign v8b9fa2 = decide_p & v88ffc1 | !decide_p & v8b9f34;
assign v845810 = hburst1_p & v845800 | !hburst1_p & !v845800;
assign v864631 = jx0_p & v852578 | !jx0_p & !v845800;
assign v88237d = decide_p & v85f58b | !decide_p & v8b9ead;
assign v88d057 = hbusreq0 & v862a8d | !hbusreq0 & !v845800;
assign jx1 = !v885c52;
assign v88a7bd = hbusreq0_p & v862032 | !hbusreq0_p & v8b9dcf;
assign v8a065e = jx1_p & v88d074 | !jx1_p & v862090;
assign v8822fa = hbusreq1 & v8a0620 | !hbusreq1 & v8a062a;
assign v8b9db6 = decide_p & v85e7e0 | !decide_p & v853cf6;
assign v8823b0 = hmastlock_p & v8b9eb4 | !hmastlock_p & !v845800;
assign v882287 = hlock1_p & v882395 | !hlock1_p & v8856cb;
assign v85f5c2 = locked_p & v85f58d | !locked_p & v845800;
assign v88231a = hready & v85afd6 | !hready & v8aff0d;
assign v88229c = decide_p & v850c63 | !decide_p & v845800;
assign v8a060a = hmastlock_p & v8626cc | !hmastlock_p & v845800;
assign v8b9e17 = hmastlock_p & v85b2d4 | !hmastlock_p & v845800;
assign v8562e6 = hready & v887065 | !hready & v85c5b2;
assign v8b9e6d = hmastlock_p & v855817 | !hmastlock_p & v84580f;
assign v851cd0 = hmastlock_p & v8b9ea7 | !hmastlock_p & !v845800;
assign v88228f = hlock0_p & v8b9e4f | !hlock0_p & v8b9f20;
assign v858df2 = hmastlock_p & v84582a | !hmastlock_p & !v845800;
assign v860700 = decide_p & v85b3e2 | !decide_p & v84581a;
assign v8a05f1 = locked_p & v855bfd | !locked_p & v8856cb;
assign v8822f4 = hready_p & v845800 | !hready_p & !v845814;
assign v85ee90 = hlock0_p & v85f59a | !hlock0_p & v845800;
assign v8606fb = hready_p & v85fec2 | !hready_p & v853612;
assign v8822e0 = hgrant1_p & v86314b | !hgrant1_p & v8535f8;
assign v8535f8 = hbusreq0_p & v8b9e0d | !hbusreq0_p & v862f33;
assign v85dedf = stateA1_p & v86028b | !stateA1_p & v8a0639;
assign v85e13d = hmaster0_p & v864e1f | !hmaster0_p & v8b9dec;
assign v8539e3 = hlock1 & v8628c9 | !hlock1 & v84581a;
assign v8623ae = start_p & v85598d | !start_p & v860b2a;
assign v8b9e55 = start_p & v85598d | !start_p & v85c7fb;
assign v8b9dc4 = hgrant1_p & v85adda | !hgrant1_p & v85880f;
assign v85d6b5 = stateA1_p & v86170f | !stateA1_p & v845800;
assign v8a05fc = hburst0_p & v85a031 | !hburst0_p & v8b9e44;
assign v89513e = hready_p & v8a0602 | !hready_p & v8822bb;
assign v885c52 = jx1_p & v864631 | !jx1_p & !v882382;
assign v88706d = decide_p & v88228f | !decide_p & v8b9dcc;
assign v8b9e13 = hmastlock_p & v85263d | !hmastlock_p & !v845800;
assign v8b9f60 = hlock0_p & v8822f4 | !hlock0_p & v845800;
assign v853cad = hbusreq1_p & v88233c | !hbusreq1_p & !v88d070;
assign v88d040 = locked_p & v8a062b | !locked_p & v8856cb;
assign v861211 = hready_p & v858327 | !hready_p & v8822bb;
assign v859006 = hready_p & v882379 | !hready_p & v845800;
assign v861c72 = decide_p & v858cdb | !decide_p & v8b9dcc;
assign v88d074 = jx0_p & v8b9edf | !jx0_p & v8b9e8f;
assign v8b9f20 = hready_p & v8b9eb8 | !hready_p & v882343;
assign v85f5b1 = decide_p & v8856ee | !decide_p & v84581a;
assign v8632bb = hlock1_p & v85fa6a | !hlock1_p & v845800;
assign v8b9e34 = hready & v8822e6 | !hready & v852fc6;
assign v87fd7e = locked_p & v882355 | !locked_p & v882343;
assign v8571d1 = hlock1_p & v88d06e | !hlock1_p & v845800;
assign v85e7b1 = hbusreq1_p & v864a19 | !hbusreq1_p & !v85c719;
assign v857931 = stateA1_p & v845800 | !stateA1_p & !v85cd0b;
assign v85f5b3 = hbusreq0_p & v8591b7 | !hbusreq0_p & v845800;
assign v8b9f17 = stateG2_p & v845800 | !stateG2_p & v85a031;
assign v856d8f = hlock0_p & v8b9f3f | !hlock0_p & v8822f4;
assign v8b9e74 = hmastlock_p & v845800 | !hmastlock_p & v845822;
assign v882379 = hbusreq1 & v8530df | !hbusreq1 & v8822b5;
assign v88d073 = hburst0_p & v8b9e25 | !hburst0_p & v862857;
assign v85f599 = hmastlock_p & v86170f | !hmastlock_p & v845800;
assign v861fa1 = stateA1_p & v8afeed | !stateA1_p & v8b9e32;
assign v8822c3 = locked_p & v85d8f3 | !locked_p & v845800;
assign v8b9f14 = hgrant1_p & v852c3b | !hgrant1_p & v85f5c5;
assign v8b9e66 = hgrant1_p & v858ab6 | !hgrant1_p & !v882349;
assign v88ffbd = hready_p & v8b9f71 | !hready_p & v8b9e0c;
assign v85fb94 = stateA1_p & v845800 | !stateA1_p & v8b9e3d;
assign v859163 = stateG3_2_p & v845800 | !stateG3_2_p & !v8b9e25;
assign v85a826 = decide_p & v8633f4 | !decide_p & v852ef0;
assign v86997d = hlock0_p & v8b9ed3 | !hlock0_p & v8b9eed;
assign v8612ae = decide_p & v85b5d3 | !decide_p & v845800;
assign v8b9e4a = locked_p & v851cd0 | !locked_p & !v845814;
assign v8822fe = locked_p & v845800 | !locked_p & v8635aa;
assign v862a20 = hready & v8b9f13 | !hready & v85f581;
assign v85b83a = locked_p & v8b9e19 | !locked_p & v845800;
assign v882348 = hready_p & v845800 | !hready_p & v88d07b;
assign v882292 = hgrant1_p & v85a7d6 | !hgrant1_p & !v887066;
assign v8b9f6c = hready & v85f5a5 | !hready & v88a7c6;
assign v864941 = hready_p & v845800 | !hready_p & v887053;
assign v8822d5 = hbusreq0_p & v8a0641 | !hbusreq0_p & !v845818;
assign jx0 = !v88d090;
assign v8b9dcc = locked_p & v864279 | !locked_p & v882343;
assign v8b9f98 = hlock0_p & v845800 | !hlock0_p & v882332;
assign v8822f1 = stateA1_p & v8600bd | !stateA1_p & v85a1b1;
assign v8b9e0c = locked_p & v8b9e35 | !locked_p & v845800;
assign v858327 = hlock1 & v8b9f58 | !hlock1 & !v85c62e;
assign v8a062c = hbusreq0_p & v852480 | !hbusreq0_p & v845800;
assign v851c6c = hbusreq0_p & v882304 | !hbusreq0_p & !v85e71f;
assign v864411 = decide_p & v85ee90 | !decide_p & v845800;
assign v8822ac = hbusreq0 & v88a7a3 | !hbusreq0 & v861063;
assign v8822cf = hbusreq0 & v85f81e | !hbusreq0 & !v845800;
assign v8b9dbe = hready_p & v845800 | !hready_p & v8b9e0b;
assign v8b9f11 = locked_p & v845800 | !locked_p & v853612;
assign v845822 = stateA1_p & v845800 | !stateA1_p & !v845800;
assign v86027d = hlock1_p & v845800 | !hlock1_p & !v8597ea;
assign v8581c3 = hbusreq1_p & v8579d6 | !hbusreq1_p & v863359;
assign v8b9e6c = locked_p & v8b9dfc | !locked_p & v845800;
assign v88a7bc = decide_p & v88228d | !decide_p & v845800;
assign v858ab6 = hbusreq0_p & v887059 | !hbusreq0_p & v85e71f;
assign v8aff12 = jx1_p & v88ffbf | !jx1_p & v8b9e22;
assign v85b4d5 = decide_p & v8b9f98 | !decide_p & v8583bf;
assign v864a19 = hgrant1_p & v85f597 | !hgrant1_p & !v857eb6;
assign v882370 = decide_p & v885713 | !decide_p & v8b9f3b;
assign v8822ff = hbusreq0_p & v895141 | !hbusreq0_p & v85cd0c;
assign v85f5be = stateA1_p & v85f5b7 | !stateA1_p & v8b9ef1;
assign v885722 = jx1_p & v861546 | !jx1_p & v8afef8;
assign v85b3e2 = hlock1_p & v8b9e1c | !hlock1_p & !v845800;
assign v882354 = stateA1_p & v88705a | !stateA1_p & !v845800;
assign v8822b0 = hmastlock_p & v856288 | !hmastlock_p & v845800;
assign v862f96 = hlock1_p & v8b9f09 | !hlock1_p & v8856cb;
assign v864cfd = hgrant1_p & v860fce | !hgrant1_p & v852475;
assign v85fbe0 = hlock0_p & v8a062d | !hlock0_p & v85b3e2;
assign v8b9f5a = hmastlock_p & v88d085 | !hmastlock_p & !v845800;
assign v8a064b = hbusreq1 & v85f592 | !hbusreq1 & v845800;
assign v885719 = jx0_p & v8b9dce | !jx0_p & !v85c7f3;
assign v85ff1e = decide_p & v8b9f81 | !decide_p & v864941;
assign v85f5c5 = hbusreq0_p & v88d076 | !hbusreq0_p & !v8b9f6e;
assign v8b9e44 = hburst1_p & v85a031 | !hburst1_p & !v845800;
assign v85d0b4 = hready_p & v8aff0b | !hready_p & v8856cb;
assign v851b5e = hready & v882306 | !hready & v85c5b2;
assign v8822b6 = start_p & v85cd0b | !start_p & v859163;
assign v861bb9 = hlock0_p & v8b9dcd | !hlock0_p & v845800;
assign v8b9ecf = hburst1_p & v8aff00 | !hburst1_p & v845800;
assign start = !v87fd86;
assign v861aaf = start_p & v84580e | !start_p & v8b9f06;
assign v8a062d = hlock1_p & v845800 | !hlock1_p & !v8822f4;
assign v8823ab = decide_p & v8b9dc2 | !decide_p & v85f58f;
assign v8afefe = hready & v86031b | !hready & v8631cf;
assign v8b9ee9 = hlock1_p & v88d044 | !hlock1_p & !v845800;
assign v8b9da6 = hbusreq1_p & v85f588 | !hbusreq1_p & v85cb5c;
assign v895132 = stateG10_1_p & v85f141 | !stateG10_1_p & !v864990;
assign v861063 = hlock1 & v845805 | !hlock1 & v845800;
assign v863eb5 = hgrant1_p & v85e71f | !hgrant1_p & !v882349;
assign v882365 = start_p & v845800 | !start_p & v8b9e9b;
assign v85c621 = hbusreq1_p & v895133 | !hbusreq1_p & !v856e69;
assign v8822c8 = hburst0_p & v845800 | !hburst0_p & v85e54f;
assign v89a6f2 = locked_p & v845800 | !locked_p & !v845814;
assign v853c79 = hlock0_p & v852a1d | !hlock0_p & v858fd3;
assign v8b9e1e = hbusreq0_p & v85a5c7 | !hbusreq0_p & v845800;
assign v8856ee = hlock1_p & v882307 | !hlock1_p & !v845800;
assign v8822bb = hmastlock_p & v85f1f2 | !hmastlock_p & v845800;
assign v863359 = hgrant1_p & v861ed5 | !hgrant1_p & v85af06;
assign v8afef6 = hgrant1_p & v845804 | !hgrant1_p & !v85c59b;
assign v85f6d6 = locked_p & v85f57f | !locked_p & v845800;
assign v8b9f56 = hbusreq1_p & v8b9e75 | !hbusreq1_p & v85654f;
assign v85c572 = hlock1 & v8b9e1f | !hlock1 & !v85c62e;
assign v887064 = decide_p & v85c70f | !decide_p & v85d6d3;
assign v8629ac = decide_p & v8b9dc1 | !decide_p & v858794;
assign v857e81 = hburst0_p & v845828 | !hburst0_p & v86482d;
assign v84580e = hburst0_p & v845800 | !hburst0_p & !v845800;
assign v862346 = hready_p & v85f58f | !hready_p & !v882343;
assign v88d087 = hready_p & v8a05f1 | !hready_p & v855bfd;
assign v859575 = hready_p & v845800 | !hready_p & !v864279;
assign v8822e6 = locked_p & v887065 | !locked_p & v845800;
assign v8b9dc3 = hlock1_p & v8631b2 | !hlock1_p & v85f67e;
assign v8b9ee3 = hlock0_p & v85fe4d | !hlock0_p & !v860625;
assign v860857 = locked_p & v8a060a | !locked_p & !v845814;
assign v85f907 = locked_p & v8539e6 | !locked_p & v845800;
assign v8600bd = start_p & v845810 | !start_p & !v8b9de6;
assign v8b9def = stateA1_p & v845800 | !stateA1_p & v845816;
assign v8b9e85 = hready & v85c75d | !hready & v88d07b;
assign v8856c6 = decide_p & v8a0611 | !decide_p & v845800;
assign v8aff0d = hmastlock_p & v8b9f80 | !hmastlock_p & !v845800;
assign v85ce61 = hlock1_p & v845800 | !hlock1_p & !v85f67e;
assign v85f67e = hready_p & v8822c4 | !hready_p & v8b9e74;
assign v8b9e67 = hgrant1_p & v85de6c | !hgrant1_p & v845807;
assign v858891 = hbusreq1 & v8b9e20 | !hbusreq1 & !v845800;
assign v85e71f = decide_p & v845800 | !decide_p & !v84581a;
assign v85ac94 = hlock1_p & v8b9dc5 | !hlock1_p & v8597ea;
assign v85957f = hmaster0_p & v8581c3 | !hmaster0_p & v862d65;
assign v845828 = stateG3_1_p & v845800 | !stateG3_1_p & !v845800;
assign v88d06d = hmastlock_p & v8823af | !hmastlock_p & !v845800;
assign v88229d = locked_p & v8b9e1d | !locked_p & !v845800;
assign v8647b7 = hbusreq0_p & v887064 | !hbusreq0_p & v857eeb;
assign v8b9e4f = hlock1_p & v88235e | !hlock1_p & v863615;
assign v8628c9 = locked_p & v8b9ec7 | !locked_p & !v845800;
assign v862a8d = hready & v852bf7 | !hready & v85f0c6;
assign v85b585 = start_p & v845800 | !start_p & !v852edf;
assign v85c70f = hlock0_p & v85d820 | !hlock0_p & v845800;
assign v8531a0 = hbusreq0_p & v8b9e92 | !hbusreq0_p & v85abe0;
assign v85f597 = hbusreq0_p & v88d077 | !hbusreq0_p & v88d062;
assign hgrant0 = !v88706f;
assign v88d07c = start_p & v845800 | !start_p & v8b9ec9;
assign v8b9ec9 = stateG2_p & v845800 | !stateG2_p & v8aff00;
assign v8b9f4d = hburst0 & v85fb02 | !hburst0 & !v845800;
assign stateG3_1 = !v895157;
assign v8b9eb4 = stateA1_p & v8822ef | !stateA1_p & !v8b9e11;
assign v856300 = start_p & v845800 | !start_p & !v85fad3;
assign v895151 = locked_p & v882332 | !locked_p & v85f58b;
assign v864523 = hbusreq0_p & v861c72 | !hbusreq0_p & !v8a05fe;
assign v88ffbf = jx0_p & v887069 | !jx0_p & v85f6f8;
assign v8a0632 = hready & v85a015 | !hready & v8b9f35;
assign v861c42 = hready & v87fd7e | !hready & v845800;
assign v858fd3 = hlock1_p & v85323a | !hlock1_p & v845800;
assign v88d071 = hbusreq0_p & v8a0610 | !hbusreq0_p & v882376;
assign v8822d4 = hlock0_p & v85ee66 | !hlock0_p & v853612;
assign v85c278 = hlock0_p & v86027d | !hlock0_p & v8b9ee9;
assign v8606e5 = hlock1_p & v88d044 | !hlock1_p & v845800;
assign v882399 = decide_p & v88230c | !decide_p & v8b9e72;
assign v863d44 = hlock1_p & v8a0618 | !hlock1_p & v845800;
assign v88229f = stateA1_p & v8b9ec8 | !stateA1_p & !v845800;
assign v8b9e04 = decide_p & v85c278 | !decide_p & v84581a;
assign v8856e1 = decide_p & v8856d6 | !decide_p & v845800;
assign v864cae = hburst0_p & v8aff00 | !hburst0_p & v8b9ecf;
assign v8618bd = jx0_p & v85e13d | !jx0_p & v8b9f0a;
assign v8a062b = start_p & v845800 | !start_p & !v882375;
assign v85e7fa = hmaster0_p & v8b9f27 | !hmaster0_p & v8afef1;
assign v8b9da5 = start_p & v85598d | !start_p & v860967;
assign v8b9f40 = stateA1_p & v845800 | !stateA1_p & v85cd0b;
assign v8620e6 = hbusreq1_p & v8b9e3e | !hbusreq1_p & v85e961;
assign v8b9e12 = hburst1_p & v87fd7a | !hburst1_p & !v845800;
assign v88ffbb = hmaster0_p & v88237a | !hmaster0_p & !v85e7b1;
assign v851256 = hbusreq0 & v88d066 | !hbusreq0 & v845800;
assign v858cdb = hlock0_p & v88235e | !hlock0_p & v8b9f20;
assign v858525 = hmastlock_p & v88706c | !hmastlock_p & v845800;
assign v857eb6 = hbusreq0_p & v88706d | !hbusreq0_p & !v8a05fe;
assign v860f3e = hbusreq0 & v85c974 | !hbusreq0 & !v845800;
assign v85afd6 = hmastlock_p & v8822f8 | !hmastlock_p & !v845800;
assign v85598d = hburst0_p & v845800 | !hburst0_p & !v845810;
assign v8b9e60 = hlock0_p & v8b9eaf | !hlock0_p & v8b9eed;
assign v8a0630 = hbusreq1_p & v85330e | !hbusreq1_p & v85654f;
assign v85bc80 = locked_p & v882365 | !locked_p & v845800;
assign v88230e = hbusreq1 & v8822ac | !hbusreq1 & !v85a9a4;
assign v856c47 = start_p & v845800 | !start_p & v859163;
assign v8b9e92 = decide_p & v853647 | !decide_p & v8a065d;
assign v8856da = hready_p & v85ae93 | !hready_p & v853612;
assign v8b9f0e = hmastlock_p & v882316 | !hmastlock_p & !v845800;
assign v88235e = hready_p & v8822a8 | !hready_p & v864279;
assign v8605e3 = hready & v8822f1 | !hready & v85ef57;
assign v85d0f7 = decide_p & v863a8a | !decide_p & v8a05f1;
assign v8822b5 = hbusreq0 & v8635aa | !hbusreq0 & v845800;
assign v88a7c6 = hmastlock_p & v87fd7f | !hmastlock_p & !v845800;
assign v8822ad = hgrant1_p & v857eeb | !hgrant1_p & v845800;
assign v8b9e19 = hmastlock_p & v8b9e55 | !hmastlock_p & v845800;
assign v845808 = hlock0_p & v845800 | !hlock0_p & !v845800;
assign v8afee6 = start_p & v845800 | !start_p & v85c5ce;
assign v8b9ed7 = hready_p & v8b9e97 | !hready_p & v845800;
assign v8b9df7 = hmastlock_p & v88d088 | !hmastlock_p & v845800;
assign v84581a = locked_p & v845800 | !locked_p & !v845800;
assign v85ad75 = hbusreq0_p & v88238b | !hbusreq0_p & !v8b9f6e;
assign v8b9e75 = hgrant1_p & v8b9ed5 | !hgrant1_p & !v85cb98;
assign v85934d = hbusreq1_p & v8822e0 | !hbusreq1_p & v845800;
assign v8b9e2d = hburst1_p & v845828 | !hburst1_p & !v845800;
assign v88238b = decide_p & v8823a9 | !decide_p & v84581a;
assign v8b9e32 = start_p & v84580e | !start_p & v8a0653;
assign v8b9e88 = hbusreq0_p & v85b4d5 | !hbusreq0_p & v885c50;
assign v85791c = locked_p & v88705d | !locked_p & v845800;
assign v8b9f48 = hbusreq0 & v88d066 | !hbusreq0 & !v8b9e34;
assign v8822f8 = stateA1_p & v885700 | !stateA1_p & !v85b585;
assign v85cd0b = hburst0_p & v845800 | !hburst0_p & v845810;
assign v8b9e0d = decide_p & v861bb9 | !decide_p & v895134;
assign v85bae3 = locked_p & v8578ef | !locked_p & v845800;
assign v887062 = hready & v8823b0 | !hready & v8b9e6d;
assign v8578f2 = decide_p & v85f7a7 | !decide_p & v8a05f1;
assign v8b9e5c = jx0_p & v852578 | !jx0_p & v851b6e;
assign v85c9ad = hlock0_p & v8602a4 | !hlock0_p & !v8822a3;
assign v855725 = hburst0_p & v859163 | !hburst0_p & v8b9f44;
assign v887065 = hmastlock_p & v855817 | !hmastlock_p & !v845800;
assign v8b9eb2 = locked_p & v85d6af | !locked_p & v85f58b;
assign v852edf = hburst0_p & v845828 | !hburst0_p & v8b9e2d;
assign v8b9f35 = stateA1_p & v845800 | !stateA1_p & !v861aaf;
assign v895141 = decide_p & v85803c | !decide_p & v8b9dcc;
assign v89a6f1 = hready & v8b9fa4 | !hready & v85ef57;
assign v88d06f = hready_p & v857751 | !hready_p & v8b9e0b;
assign v85f85f = hlock1_p & v845800 | !hlock1_p & v88d044;
assign v8b9e41 = hready & v8822b0 | !hready & v88d07b;
assign v8635aa = hmastlock_p & v85d6b5 | !hmastlock_p & v845800;
assign v855d10 = hlock0_p & v852a1d | !hlock0_p & v85ce69;
assign v85f5b5 = hlock0_p & v8b9f64 | !hlock0_p & v845800;
assign v8b9f57 = decide_p & v882287 | !decide_p & v853cf6;
assign v8b9e1f = locked_p & v8a0609 | !locked_p & v845800;
assign v8b9f4c = hlock1_p & v8b9ea0 | !hlock1_p & v8b9dbe;
assign hgrant1 = v8a065e;
assign v8b9dec = hbusreq1_p & v85cc6b | !hbusreq1_p & v85e753;
assign v882343 = hmastlock_p & v8afeef | !hmastlock_p & v845822;
assign v85a4b1 = hready_p & v85f907 | !hready_p & v88705d;
assign v8823af = stateA1_p & v8afeed | !stateA1_p & !v8b9ef0;
assign v8aff03 = locked_p & v882291 | !locked_p & !v845814;
assign v8b9ed3 = hlock1_p & v89a6f4 | !hlock1_p & !v8856f0;
assign v88a7aa = hready_p & v859d8d | !hready_p & v88235a;
assign v8a0282 = hbusreq1_p & v845800 | !hbusreq1_p & v84581e;
assign v85fd24 = hbusreq0_p & v8856e1 | !hbusreq0_p & v845800;
assign v88238a = start_p & v85cd0b | !start_p & !v845824;
assign v859035 = locked_p & v85f5c1 | !locked_p & v845800;
assign v850934 = hlock1_p & v882307 | !hlock1_p & v845800;
assign v8a065d = hready_p & v845800 | !hready_p & v855d31;
assign v852480 = decide_p & v895135 | !decide_p & v845800;
assign v8b9f09 = hready_p & v8856cb | !hready_p & v855bfd;
assign v8505a9 = hlock1_p & v8856da | !hlock1_p & v845800;
assign v8b71a5 = hbusreq1 & v851256 | !hbusreq1 & !v8b9dbb;
assign v88233c = hgrant1_p & v85a826 | !hgrant1_p & v8b9dd1;
assign v88d052 = hburst0_p & v87fd7a | !hburst0_p & v8b9e00;
assign v85f81e = hready & v882285 | !hready & v887065;
assign v85d6af = hmastlock_p & v85f5be | !hmastlock_p & !v845800;
assign v882391 = hmaster0_p & v85c89c | !hmaster0_p & v845800;
assign v8a061b = decide_p & v8b9dd1 | !decide_p & v845800;
assign v85f5a5 = locked_p & v8b9e2c | !locked_p & v845800;
assign v8a05fa = hlock1_p & v88235e | !hlock1_p & v8b9f20;
assign v85029d = hbusreq1_p & v882292 | !hbusreq1_p & v85e753;
assign v8602a4 = hlock1_p & v845800 | !hlock1_p & v8b9e1c;
assign v8b9e49 = hready_p & v845800 | !hready_p & v88230e;
assign v864246 = hmaster0_p & v85c621 | !hmaster0_p & !v85e7b1;
assign v85a1b1 = start_p & v845810 | !start_p & !v8b9e25;
assign v8afee2 = locked_p & v858cf2 | !locked_p & v882343;
assign v85f5af = stateA1_p & v8b9ec8 | !stateA1_p & !v8b9ef0;
assign v85688b = hlock0_p & v857768 | !hlock0_p & v882343;
assign v8a0613 = hmastlock_p & v857931 | !hmastlock_p & v845822;
assign v8823a9 = hlock0_p & v85f85f | !hlock0_p & !v85ce69;
assign v8b9eaf = hlock1_p & v8631b2 | !hlock1_p & !v861211;
assign v88237a = hbusreq1_p & v895133 | !hbusreq1_p & !v8b9e06;
assign v862f88 = hlock1 & v88ffba | !hlock1 & v8afefe;
assign v862090 = hmaster0_p & v864e1f | !hmaster0_p & v859ca9;
assign v85a015 = stateA1_p & v845800 | !stateA1_p & v856300;
assign v862d65 = hgrant1_p & v85abe0 | !hgrant1_p & v8b9deb;
assign v8b9e3d = start_p & v845800 | !start_p & v855725;
assign v85a7d6 = hbusreq0_p & v8856c6 | !hbusreq0_p & v88228e;
assign v852fc6 = stateA1_p & v8623ae | !stateA1_p & !v852fbe;
assign v85e4a1 = stateG3_1_p & v845826 | !stateG3_1_p & v845800;
assign v8822fc = hmastlock_p & v863d0e | !hmastlock_p & v845800;
assign v8b9dc6 = hready & v8b9e4a | !hready & v860857;
assign v882355 = hmastlock_p & v88ffd0 | !hmastlock_p & v845800;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  jx0_p = 0;
  jx1_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  jx0_p = jx0;
  jx1_p = jx1;
    end
endmodule

