module main(clock, hready, hbusreq0, hlock0, hbusreq1, hlock1, hbusreq2, hlock2, hburst0, hburst1, hmaster0, hmaster1, hmastlock, start, decide, locked, hgrant0, hgrant1, hgrant2, busreq, stateA1, stateG2, stateG3_0, stateG3_1, stateG3_2, stateG10_1, stateG10_2, jx0, jx1, jx2);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v84563c;
  wire v845650;
  wire v866c94;
  wire v86cfb3;
  wire v87f892;
  wire v973883;
  wire v845666;
  wire v973884;
  wire v973885;
  wire v973886;
  wire v973887;
  wire v973888;
  wire v973889;
  wire v97388a;
  wire v97388b;
  wire v97388c;
  wire v97388d;
  wire v97388e;
  wire v97388f;
  wire v973890;
  wire v973891;
  wire v973892;
  wire v973893;
  wire v973894;
  wire v973895;
  wire v973896;
  wire v973897;
  wire v973898;
  wire v973899;
  wire v97389a;
  wire v97389b;
  wire v97389c;
  wire v97389d;
  wire v97389e;
  wire v97389f;
  wire v9738a0;
  wire v9738a1;
  wire v9738a2;
  wire v9738a3;
  wire v9738a4;
  wire v9738a5;
  wire v9738a6;
  wire v9738a7;
  wire v9738a8;
  wire v9738a9;
  wire v9738aa;
  wire v9738ab;
  wire v9738ac;
  wire v9738ad;
  wire v9738ae;
  wire v9738af;
  wire v9738b0;
  wire v9738b1;
  wire v9738b2;
  wire v9738b3;
  wire v9738b4;
  wire v9738b5;
  wire v9738b6;
  wire v9738b7;
  wire v9738b8;
  wire v9738b9;
  wire v9738ba;
  wire v9738bb;
  wire v9738bc;
  wire v9738bd;
  wire v9738be;
  wire v9738bf;
  wire v9738c0;
  wire v9738c1;
  wire v9738c2;
  wire v9738c3;
  wire v9738c4;
  wire v9738c5;
  wire v9738c6;
  wire v9738c7;
  wire v9738c8;
  wire v9738c9;
  wire v9738ca;
  wire v9738cb;
  wire v9738cc;
  wire v9738cd;
  wire v9738ce;
  wire v9738cf;
  wire v9738d0;
  wire v9738d1;
  wire v9738d2;
  wire v9738d3;
  wire v9738d4;
  wire v9738d5;
  wire v9738d6;
  wire v9738d7;
  wire v9738d8;
  wire v9738d9;
  wire v9738da;
  wire v9738db;
  wire v9738dc;
  wire v9738dd;
  wire v9738de;
  wire v9738df;
  wire v9738e0;
  wire v9738e1;
  wire v9738e2;
  wire v9738e3;
  wire v9738e4;
  wire v9738e5;
  wire v9738e6;
  wire v9738e7;
  wire v9738e8;
  wire v9738e9;
  wire v9738ea;
  wire v9738eb;
  wire v9738ec;
  wire v9738ed;
  wire v9738ee;
  wire v9738ef;
  wire v9738f0;
  wire v9738f1;
  wire v9738f2;
  wire v9738f3;
  wire v9738f4;
  wire v9738f5;
  wire v9738f6;
  wire v9738f7;
  wire v9738f8;
  wire v9738f9;
  wire v9738fa;
  wire v9738fb;
  wire v9738fc;
  wire v9738fd;
  wire v9738fe;
  wire v9738ff;
  wire v973900;
  wire v973901;
  wire v973902;
  wire v973903;
  wire v973904;
  wire v973905;
  wire v973906;
  wire v973907;
  wire v973908;
  wire v973909;
  wire v97390a;
  wire v97390b;
  wire v97390c;
  wire v97390d;
  wire v97390e;
  wire v97390f;
  wire v973910;
  wire v973911;
  wire v973912;
  wire v973913;
  wire v973914;
  wire v973915;
  wire v973916;
  wire v973917;
  wire v973918;
  wire v973919;
  wire v97391a;
  wire v97391b;
  wire v97391c;
  wire v97391d;
  wire v97391e;
  wire v97391f;
  wire v973920;
  wire v973921;
  wire v973922;
  wire v973923;
  wire v973924;
  wire v973925;
  wire v973926;
  wire v973927;
  wire v973928;
  wire v973929;
  wire v97392a;
  wire v97392b;
  wire v97392c;
  wire v97392d;
  wire v97392e;
  wire v97392f;
  wire v973930;
  wire v973931;
  wire v973932;
  wire v973933;
  wire v973934;
  wire v973935;
  wire v973936;
  wire v973937;
  wire v973938;
  wire v973939;
  wire v97393a;
  wire v97393b;
  wire v97393c;
  wire v97393d;
  wire v97393e;
  wire v97393f;
  wire v973940;
  wire v973941;
  wire v973942;
  wire v973943;
  wire v973944;
  wire v973945;
  wire v973946;
  wire v973947;
  wire v973948;
  wire v973949;
  wire v97394a;
  wire v97394b;
  wire v97394c;
  wire v97394d;
  wire v97394e;
  wire v97394f;
  wire v973950;
  wire v973951;
  wire v973952;
  wire v973953;
  wire v973954;
  wire v973955;
  wire v973956;
  wire v973957;
  wire v973958;
  wire v973959;
  wire v97395a;
  wire v97395b;
  wire v97395c;
  wire v97395d;
  wire v97395e;
  wire v97395f;
  wire v973960;
  wire v973961;
  wire v973962;
  wire v973963;
  wire v973964;
  wire v973965;
  wire v973966;
  wire v973967;
  wire v973968;
  wire v973969;
  wire v97396a;
  wire v97396b;
  wire v97397b;
  wire v97397c;
  wire v97397d;
  wire v97397e;
  wire v97397f;
  wire v973980;
  wire v973981;
  wire v973982;
  wire v973983;
  wire v973984;
  wire v973985;
  wire v973986;
  wire v973987;
  wire v973988;
  wire v973989;
  wire v97398a;
  wire v97398b;
  wire v97398c;
  wire v97398d;
  wire v97398e;
  wire v97398f;
  wire v973990;
  wire v973991;
  wire v973992;
  wire v973993;
  wire v973994;
  wire v973995;
  wire v973996;
  wire v973997;
  wire v973998;
  wire v973999;
  wire v97399a;
  wire v97399b;
  wire v97399c;
  wire v97399d;
  wire v97399e;
  wire v97399f;
  wire v9739a0;
  wire v9739a1;
  wire v9739a2;
  wire v9739a3;
  wire v9739a4;
  wire v9739a5;
  wire v9739a6;
  wire v9739a7;
  wire v9739a8;
  wire v9739a9;
  wire v9739aa;
  wire v9739ab;
  wire v9739ac;
  wire v9739ad;
  wire v9739ae;
  wire v9739af;
  wire v9739b3;
  wire v9739b4;
  wire v9739b5;
  wire v9739b6;
  wire v9739b7;
  wire v9739b8;
  wire v9739b9;
  wire v9739ba;
  wire v9739bb;
  wire v9739bc;
  wire v9739bd;
  wire v9739be;
  wire v9739bf;
  wire v9739c0;
  wire v9739c1;
  wire v9739c2;
  wire v9739c3;
  wire v9739c4;
  wire v9739c5;
  wire v9739c6;
  wire v9739c7;
  wire v9739c8;
  wire v9739c9;
  wire v9739ca;
  wire v9739cb;
  wire v9739cc;
  wire v9739cd;
  wire v9739ce;
  wire v9739cf;
  wire v9739d0;
  wire v9739d1;
  wire v9739d2;
  wire v9739d3;
  wire v9739d4;
  wire v9739d5;
  wire v9739d6;
  wire v9739d7;
  wire v9739d8;
  wire v9739d9;
  wire v9739da;
  wire v9739db;
  wire v9739dc;
  wire v9739dd;
  wire v9739de;
  wire v9739df;
  wire v9739e0;
  wire v9739e1;
  wire v9739e2;
  wire v9739e3;
  wire v9739e4;
  wire v9739e5;
  wire v9739e6;
  wire v9739e7;
  wire v9739e8;
  wire v9739e9;
  wire v9739ea;
  wire v9739eb;
  wire v9739ec;
  wire v9739ed;
  wire v9739ee;
  wire v9739ef;
  wire v9739f0;
  wire v9739f1;
  wire v9739f2;
  wire v9739f4;
  wire v9739f5;
  wire v9739f6;
  wire v9739f7;
  wire v9739f8;
  wire v9739f9;
  wire v9739fa;
  wire v9739fb;
  wire v9739fc;
  wire v9739fd;
  wire v9739fe;
  wire v9739ff;
  wire v973a00;
  wire v973a01;
  wire v973a02;
  wire v973a03;
  wire v973a04;
  wire v973a05;
  wire v973a06;
  wire v973a07;
  wire v973a08;
  wire v973a09;
  wire v973a0b;
  wire v973a0c;
  wire v973a0d;
  wire v973a0e;
  wire v973a0f;
  wire v973a10;
  wire v973a11;
  wire v973a12;
  wire v973a13;
  wire v973a14;
  wire v973a15;
  wire v973a16;
  wire v973a17;
  wire v973a18;
  wire v973a19;
  wire v973a1b;
  wire v973a1c;
  wire v973a1d;
  wire v973a1e;
  wire v973a1f;
  wire v973a20;
  wire v973a21;
  wire v973a22;
  wire v973a23;
  wire v973a24;
  wire v973a25;
  wire v973a26;
  wire v973a27;
  wire v973a28;
  wire v973a29;
  wire v973a2a;
  wire v973a2b;
  wire v973a2c;
  wire v973a2d;
  wire v973a2e;
  wire v973a2f;
  wire v973a30;
  wire v973a31;
  wire v973a32;
  wire v973a33;
  wire v973a34;
  wire v973a35;
  wire v973a36;
  wire v973a37;
  wire v973a38;
  wire v973a39;
  wire v973a3a;
  wire v973a3b;
  wire v973a3c;
  wire v973a3d;
  wire v973a3e;
  wire v973a3f;
  wire v973a40;
  wire v973a41;
  wire v973a42;
  wire v973a43;
  wire v973a44;
  wire v973a45;
  wire v973a46;
  wire v973a47;
  wire v973a48;
  wire v973a49;
  wire v973a4a;
  wire v973a4b;
  wire v973a4c;
  wire v845662;
  wire a4ce72;
  wire v845646;
  wire v845660;
  wire v9f3568;
  wire v9f3569;
  wire v9f356a;
  wire v9f356b;
  wire v9f356c;
  wire v9f3574;
  wire v9f3575;
  wire v9f3576;
  wire v9f3577;
  wire v9f3578;
  wire v9f357b;
  wire v86292d;
  wire v854658;
  wire v9d44bf;
  wire v845652;
  wire v85bb54;
  wire v8543c7;
  wire v9d44c3;
  wire v9d44c4;
  wire v9d44c5;
  wire v84566c;
  wire v8e7988;
  wire v8e7989;
  wire v845658;
  wire v887862;
  wire v8e798a;
  wire v8e798b;
  wire v8e798c;
  wire v8e7990;
  wire v8e7991;
  wire v8e7992;
  wire v8e7993;
  wire v8e7994;
  wire v8e7995;
  wire v8e7996;
  wire v8e7997;
  wire v8e7998;
  wire v8e7999;
  wire v8e799a;
  wire v8e799b;
  wire v8e799c;
  wire v8e799d;
  wire v8e799e;
  wire v8e799f;
  wire v8e79a0;
  wire v8e79a1;
  wire v8e79a2;
  wire v8e79a3;
  wire v8e79a4;
  wire v8e79a5;
  wire v8e79a6;
  wire v8e79a7;
  wire v8e79a8;
  wire v8e79a9;
  wire v8e79aa;
  wire v8e79ab;
  wire v8e79ac;
  wire v8e79ad;
  wire v8e79ae;
  wire v8e79af;
  wire v8e79b0;
  wire v8e79b1;
  wire v8e79b2;
  wire v8e79b3;
  wire v8e79b4;
  wire v8e79b5;
  wire v8e79b6;
  wire v8e79b7;
  wire v8e79b8;
  wire v8e79b9;
  wire v8e79ba;
  wire v8e79bb;
  wire v8e79bc;
  wire v8e79bd;
  wire v8e79be;
  wire v8e79bf;
  wire v8e79c0;
  wire v8e79c1;
  wire v8e79c2;
  wire v8e79c3;
  wire v8e79c4;
  wire v8e79c5;
  wire v8e79c6;
  wire v8e79c7;
  wire v8e79c8;
  wire v8e79c9;
  wire v8e79ca;
  wire v8e79cb;
  wire v8e79cc;
  wire v8e79cd;
  wire v8e79ce;
  wire v8e79cf;
  wire v8e79d0;
  wire v8e79d1;
  wire v8e79d2;
  wire v8e79d3;
  wire v8e79d4;
  wire v8e79d5;
  wire v8e79d6;
  wire v8e79d7;
  wire v8e79d8;
  wire v8e79d9;
  wire v8e79da;
  wire v8e79db;
  wire v960f65;
  wire v84565e;
  wire v960f66;
  wire v960f67;
  wire v8901af;
  wire v861283;
  wire v878a51;
  wire v8996a7;
  wire v883467;
  wire v8c1118;
  wire v8c1119;
  wire v8c111a;
  wire v8c111b;
  wire v8c111c;
  wire v8c111d;
  wire v8c111e;
  wire v92337e;
  wire v8c111f;
  wire v8c1120;
  wire v8c1121;
  wire v8c1122;
  wire v8c1123;
  wire v8c1124;
  wire v8c1125;
  wire v8c1126;
  wire v8c1127;
  wire v8c1128;
  wire v8c1129;
  wire v8c112a;
  wire v8c112b;
  wire v8c112c;
  wire v8c112d;
  wire v8c112e;
  wire v8c112f;
  wire v8c1130;
  wire v8c1131;
  wire v8c1132;
  wire v8c1133;
  wire v8c1134;
  wire v8c1135;
  wire v8c1136;
  wire v8c1137;
  wire v8c1138;
  wire v8c1139;
  wire v8c113a;
  wire v8c113b;
  wire v8c113c;
  wire v8c113d;
  wire v8c113e;
  wire v8c113f;
  wire v8c1140;
  wire v8c1141;
  wire v8c1142;
  wire v8c1143;
  wire v8c1144;
  wire v8c1145;
  wire v8c1146;
  wire v8c1147;
  wire v8c1148;
  wire v8c1149;
  wire v8c114a;
  wire v87bd68;
  wire v8768ab;
  wire v8c114b;
  wire v8c114c;
  wire v8c114d;
  wire v8c114e;
  wire v8c114f;
  wire v8c1150;
  wire v8c1151;
  wire v8c1152;
  wire v8c1153;
  wire v8c1154;
  wire v8c1155;
  wire v8c1156;
  wire v8c1157;
  wire v8c1158;
  wire v8c1159;
  wire v8c115a;
  wire v8c115b;
  wire v8c115c;
  wire v8c115d;
  wire v8c115e;
  wire v8c115f;
  wire v8c1160;
  wire v8c1161;
  wire v8c1162;
  wire v8c1163;
  wire v8c1164;
  wire v8c1165;
  wire v8c1166;
  wire v8c1167;
  wire v8c1168;
  wire v8c1169;
  wire v8c116a;
  wire v8c116b;
  wire v8c116c;
  wire v8c116d;
  wire v8c116e;
  wire v8c116f;
  wire v8c1170;
  wire v8c1171;
  wire v8c1172;
  wire v8c1173;
  wire v8c1174;
  wire v8c1175;
  wire v8c1176;
  wire v8c1177;
  wire v8c1178;
  wire v8c1179;
  wire v8c117a;
  wire v8c117b;
  wire v8c117c;
  wire v8c117d;
  wire v8c117e;
  wire v8c117f;
  wire v8c1180;
  wire v8ea7e2;
  wire v8ea7e3;
  wire v8ea7e4;
  wire v8ea7e5;
  wire v8ea7e6;
  wire v8ea7e7;
  wire v8ea7e8;
  wire v84566e;
  wire v8ecba9;
  wire v8ea7e9;
  wire v8ea7ea;
  wire v8ea7eb;
  wire v8ea7ec;
  wire v8ea7ed;
  wire v8ea7ee;
  wire v8ea7ef;
  wire v8ea7f0;
  wire v8ea7f1;
  wire v8ea7f2;
  wire v8ea7f3;
  wire v8ea7f4;
  wire v8ea7f5;
  wire v8ea7f6;
  wire v8ea7f7;
  wire v8ea7f8;
  wire v8ea7f9;
  wire v84566a;
  wire v8ea7fa;
  wire v8ea7fb;
  wire v8ea7fc;
  wire v8ea7fd;
  wire v8ea7fe;
  wire v8ea7ff;
  wire v8ea800;
  wire v8ea801;
  wire v8ea802;
  wire v8ea803;
  wire v8ea804;
  wire v8ea805;
  wire v8ea806;
  wire v8ea807;
  wire v8ea808;
  wire v8ea809;
  wire v8ea80a;
  wire v8ea80b;
  wire v8ea80c;
  wire v8ea80d;
  wire v8ea80e;
  wire v8ea80f;
  wire v8ea810;
  wire v8ea811;
  wire v8ea812;
  wire v8ea813;
  wire v8ea814;
  wire v8ea815;
  wire v8ea816;
  wire v8ea817;
  wire v8ea818;
  wire v8ea819;
  wire v8ea81a;
  wire v8ea81b;
  wire v8ea81c;
  wire v8ea81d;
  wire v8ea81e;
  wire v8ea81f;
  wire v8ea820;
  wire v8ea821;
  wire v8ea822;
  wire v8ea823;
  wire v8ea825;
  wire v8ea826;
  wire v8ea827;
  wire v8ea828;
  wire v8ea829;
  wire v8ea82a;
  wire v8ea82b;
  wire v8ea82c;
  wire v8ea82d;
  wire v8ea82e;
  wire v8ea82f;
  wire v8ea830;
  wire v8ea831;
  wire v8ea832;
  wire v8ea833;
  wire v8ea834;
  wire v8ea835;
  wire v8ea836;
  wire v8ea837;
  wire v8ea838;
  wire v8ea839;
  wire v8ea83a;
  wire v8ea83b;
  wire v8ea83c;
  wire v8ea83d;
  wire v8ea83e;
  wire v8ea83f;
  wire v8ea840;
  wire v8ea841;
  wire v8ea842;
  wire v8ea843;
  wire v8ea844;
  wire v8ea845;
  wire v8ea846;
  wire v8ea847;
  wire v8ea848;
  wire v8ea849;
  wire v8ea84a;
  wire v8ea84b;
  wire v8ea84c;
  wire v8ea84d;
  wire v8ea84e;
  wire v8ea84f;
  wire v8ea850;
  wire v8ea851;
  wire v8ea852;
  wire v8ea853;
  wire v8ea854;
  wire v8ea855;
  wire v8ea856;
  wire v8ea857;
  wire v8ea858;
  wire v8ea859;
  wire v8ea85a;
  wire v8ea85b;
  wire v8ea85c;
  wire v8ea85d;
  wire v8ea85e;
  wire v8ea85f;
  wire v8ea860;
  wire v8ea861;
  wire v8ea862;
  wire v8ea863;
  wire v8ea864;
  wire v8ea865;
  wire v8ea866;
  wire v8ea867;
  wire v8ea868;
  wire v8ea869;
  wire v8ea86a;
  wire v8ea86b;
  wire v8ea86c;
  wire v8ea86d;
  wire v8ea86e;
  wire v8ea86f;
  wire v8ea870;
  wire v8ea871;
  wire v8ea872;
  wire v8ea873;
  wire v8ea874;
  wire v8ea875;
  wire v8ea876;
  wire v8ea877;
  wire v8ea878;
  wire v8ea879;
  wire v8ea87a;
  wire v8ea87b;
  wire v8ea87c;
  wire v8ea87d;
  wire v8ea87e;
  wire v8ea87f;
  wire v8ea880;
  wire v8ea881;
  wire v8ea882;
  wire v8ea883;
  wire v8ea884;
  wire v8ea886;
  wire v8ea887;
  wire v8ea888;
  wire v8ea889;
  wire v8ea88b;
  wire v8ea88c;
  wire v8ea88d;
  wire v8ea88e;
  wire v8ea88f;
  wire v8ea890;
  wire v8ea891;
  wire v8ea892;
  wire v8ea893;
  wire v8ea895;
  wire v8ea896;
  wire v8ea897;
  wire v8ea898;
  wire v8ea899;
  wire v8ea89a;
  wire v8ea89b;
  wire v8ea89c;
  wire v8ea89d;
  wire v8ea89e;
  wire v8ea89f;
  wire v8ea8a0;
  wire v8ea8a1;
  wire v8ea8a2;
  wire v8ea8a3;
  wire v8ea8a4;
  wire v8ea8a5;
  wire v8ea8a6;
  wire v8ea8a7;
  wire v8ea8a8;
  wire v8ea8a9;
  wire v8ea8aa;
  wire v8ea8ab;
  wire v8ea8ac;
  wire v8ea8ad;
  wire v8ea8ae;
  wire v8ea8af;
  wire v8ea8b0;
  wire v8ea8b1;
  wire v8ea8b2;
  wire v8ea8b3;
  wire v8ea8b4;
  wire v8ea8b5;
  wire v8ea8b6;
  wire v8ea8b7;
  wire v8ea8b8;
  wire v8ea8b9;
  wire v8ea8ba;
  wire v8ea8bb;
  wire v8ea8bc;
  wire v8ea8bd;
  wire v8ea8be;
  wire v8ea8bf;
  wire v8ea8c0;
  wire v8ea8c1;
  wire v8ea8c2;
  wire v8ea8c3;
  wire v8ea8c4;
  wire v8ea8c5;
  wire v8ea8c6;
  wire v8ea8c7;
  wire v8ea8c8;
  wire v8ea8c9;
  wire v8ea8ca;
  wire v8ea8cb;
  wire v8ea8cc;
  wire v8ea8cd;
  wire v8ea8ce;
  wire v8ea8cf;
  wire v8ea8d0;
  wire v8ea8d1;
  wire v8ea8d2;
  wire v8ea8d3;
  wire v8ea8d4;
  wire v8ea8d5;
  wire v8ea8d6;
  wire v8ea8d7;
  wire v8ea8d8;
  wire v8ea8d9;
  wire v8ea8da;
  wire v8ea8db;
  wire v8ea8dc;
  wire v8ea8dd;
  wire v8ea8de;
  wire v8ea8df;
  wire v8ea8e0;
  wire v8ea8e1;
  wire v8ea8e2;
  wire v8ea8e3;
  wire v8ea8e4;
  wire v8ea8e5;
  wire v8ea8e6;
  wire v8ea8e7;
  wire v8ea8e8;
  wire v8ea8e9;
  wire v8ea8ea;
  wire v8ea8eb;
  wire v8ea8ec;
  wire v8ea8ed;
  wire v8ea8ee;
  wire v8ea8ef;
  wire v8ea8f0;
  wire v8ea8f1;
  wire v8ea8f2;
  wire v8ea8f3;
  wire v8ea8f4;
  wire v8ea8f5;
  wire v8ea8f6;
  wire v8ea8f7;
  wire v8ea8f8;
  wire v8ea903;
  wire v8ea904;
  wire v8ea905;
  wire v8ea906;
  wire v8ea907;
  wire v8ea908;
  wire v8ea909;
  wire v8ea90a;
  wire v8ea90b;
  wire v8ea90c;
  wire v8ea90d;
  wire v8ea90e;
  wire v8ea90f;
  wire v8ea910;
  wire v8ea911;
  wire v8ea912;
  wire v8ea913;
  wire v8ea914;
  wire v8ea915;
  wire v8ea916;
  wire v8ea918;
  wire v8ea919;
  wire v8ea91a;
  wire v8ea91b;
  wire v8ea91c;
  wire v8ea91d;
  wire v8ea91e;
  wire v8ea91f;
  wire v8ea920;
  wire v8ea921;
  wire v8ea922;
  wire v8ea923;
  wire v8ea924;
  wire v8ea925;
  wire v8ea926;
  wire v8ea927;
  wire v8ea928;
  wire v8ea929;
  wire v8ea92a;
  wire v8ea92b;
  wire v8ea92c;
  wire v8ea92d;
  wire v8ea92e;
  wire v8ea92f;
  wire v8ea930;
  wire v8ea931;
  wire v8ea932;
  wire v8ea933;
  wire v8ea934;
  wire v8ea935;
  wire v8ea936;
  wire v8ea937;
  wire v8ea938;
  wire v8ea939;
  wire v8ea93a;
  wire v8ea93b;
  wire v8ea93c;
  wire v84565c;
  wire v8c20b6;
  wire v8c20b7;
  wire v8c20b8;
  wire v8c20b9;
  wire v845656;
  wire v8c20ba;
  wire v8c20bb;
  wire v8c20bc;
  wire v8c20bd;
  wire v8c20be;
  wire v8c20bf;
  wire v8c20c0;
  wire v8c20c1;
  wire v8c20c2;
  wire v8c20c3;
  wire v8c20c4;
  wire v8c20c5;
  wire v8c20c6;
  wire v8c20c7;
  wire v8c20c8;
  wire v8c20c9;
  wire v8c20ca;
  wire v8c20cb;
  wire v8c20cc;
  wire v8c20cd;
  wire v8c20ce;
  wire v8c20cf;
  wire v8c20d0;
  wire v8c20d1;
  wire v8c20d2;
  wire v8c20d3;
  wire v8c20d4;
  wire v8c20d5;
  wire v8c20d6;
  wire v8c20d7;
  wire v8c20d8;
  wire v8c20d9;
  wire v8c20da;
  wire v8c20db;
  wire v8c20dc;
  wire v8c20dd;
  wire v8c20de;
  wire v8c20df;
  wire v8c20e0;
  wire v8c20e1;
  wire a153b7;
  wire a153ba;
  wire a153bb;
  wire a153bc;
  wire a153bd;
  wire a153c0;
  wire a153c1;
  wire a153c2;
  wire a153c3;
  wire a153c4;
  wire a153c5;
  wire v845648;
  wire a153c8;
  wire a153c9;
  wire v85a40d;
  wire v863b4b;
  wire v8763e4;
  wire v96ef3e;
  wire a153ca;
  wire a153cb;
  wire a153cc;
  wire a153cd;
  wire a153ce;
  wire a153cf;
  wire v972fac;
  wire a153d0;
  wire a153d1;
  wire a153d2;
  wire a153d3;
  wire a153d4;
  wire a153d5;
  wire a153d6;
  wire a153e7;
  wire a153e8;
  wire a153e9;
  wire a153ea;
  wire a153eb;
  wire a153ec;
  wire a15408;
  wire a15409;
  wire a1540a;
  wire a1540b;
  wire a1540c;
  wire a1540d;
  wire a1540e;
  wire a15414;
  wire a15415;
  wire a15416;
  wire a15417;
  wire a1541d;
  wire a1541e;
  wire a1541f;
  wire a15420;
  wire a15421;
  wire a15422;
  wire a1542d;
  wire a1542e;
  wire a1542f;
  wire a15430;
  wire a15431;
  wire a15432;
  wire a15433;
  wire a15434;
  wire a15444;
  wire a15445;
  wire a15446;
  wire a15447;
  wire a15448;
  wire a15449;
  wire a15483;
  wire a15484;
  wire a15485;
  wire a15486;
  wire a15487;
  wire a15488;
  wire a15489;
  wire a1548c;
  wire a1548d;
  wire a15491;
  wire a15492;
  wire a15493;
  wire a15494;
  wire a15495;
  wire a15496;
  wire a154a1;
  wire a154a2;
  wire a154a3;
  wire a154a4;
  wire a154a5;
  wire a154a6;
  wire v845644;
  wire a154bb;
  wire a154bc;
  wire a154c1;
  wire a154c2;
  wire a154c3;
  wire a154d1;
  wire a154d2;
  wire a154d3;
  wire a154d4;
  wire a154d5;
  wire a154d6;
  wire a154ed;
  wire a154ee;
  wire a154ef;
  wire a154f0;
  wire a154f1;
  wire a154f2;
  wire a154f3;
  wire a154f5;
  wire a154f6;
  wire a154fb;
  wire a154fc;
  wire a154fd;
  wire a154fe;
  wire a154ff;
  wire a15500;
  wire a15507;
  wire a15508;
  wire a15509;
  wire a1550a;
  wire a1550b;
  wire a1550c;
  wire a1550e;
  wire a15517;
  wire a14d3c;
  wire a14d3d;
  wire a14d3e;
  wire a14d3f;
  wire a14d40;
  wire a14d42;
  wire a14d49;
  wire a14d4a;
  wire v845642;
  wire a14d4b;
  wire a14d4c;
  wire a14d4d;
  wire a14d58;
  wire a14d59;
  wire a14d5a;
  wire a14d5b;
  wire a14d5c;
  wire a14d5d;
  wire a14d67;
  wire a14d68;
  wire a14d6d;
  wire a14d6e;
  wire a14d6f;
  wire a14d70;
  wire a14d71;
  wire a14d72;
  wire a14d85;
  wire a14d8b;
  wire a14d8c;
  wire a14d8d;
  wire a14d8e;
  wire a14d9f;
  wire a14da0;
  wire a14da1;
  wire a14da2;
  wire a14da4;
  wire a14da6;
  wire a14da7;
  wire a14da8;
  wire a14da9;
  wire a14daa;
  wire a14dab;
  wire a14dad;
  wire a14dae;
  wire a14daf;
  wire a14dba;
  wire a14dbe;
  wire a14dbf;
  wire a14dc0;
  wire a14dc1;
  wire a14dc2;
  wire v9ed40e;
  wire v9ed40f;
  wire v9ed410;
  wire v9ed411;
  wire v9ed412;
  wire v9ed413;
  wire v9ed414;
  wire v9ed415;
  wire v9ed416;
  wire v9ed417;
  wire v9ed418;
  wire v9ed419;
  wire v9ed41a;
  wire v9ed41b;
  wire v9ed41c;
  wire v9ed41d;
  wire v9ed41e;
  wire v9ed41f;
  wire v9ed420;
  wire v9ed421;
  wire v9ed422;
  wire v9ed423;
  wire v9ed424;
  wire v9ed425;
  wire v9ed426;
  wire v9ed427;
  wire v9ed428;
  wire v9ed429;
  wire v9ed42a;
  wire v9ed42b;
  wire v9ed42c;
  wire v9ed42d;
  wire v9ed42e;
  wire v9ed42f;
  wire v9ed430;
  wire v9ed431;
  wire v9ed432;
  wire v9ed433;
  wire v9ed434;
  wire v9ed435;
  wire v9ed436;
  wire v9ed437;
  wire v9ed438;
  wire v9ed439;
  wire v9ed43a;
  wire v9ed43b;
  wire v9ed43c;
  wire v9ed43d;
  wire v9ed43e;
  wire v9ed43f;
  wire v9ed440;
  wire v9ed441;
  wire v9ed442;
  wire v9ed443;
  wire v9ed444;
  wire v9ed445;
  wire v9ed446;
  wire v9ed447;
  wire v9ed448;
  wire v9ed449;
  wire v9ed44a;
  wire v9ed44b;
  wire v9ed44c;
  wire v9ed44d;
  wire v9ed44e;
  wire v9ed44f;
  wire v9ed450;
  wire v9ed451;
  wire v9ed452;
  wire v9ed453;
  wire v9ed454;
  wire v9ed455;
  wire v9ed456;
  wire v9ed457;
  wire v9ed458;
  wire v9ed459;
  wire v9ed45a;
  wire v9ed45b;
  wire v9ed45c;
  wire v9ed45d;
  wire a2bd3c;
  wire a2bd3d;
  wire v9ed45e;
  wire v9ed45f;
  wire v9ed460;
  wire v9ed461;
  wire v9ed462;
  wire v9ed463;
  wire a2bd45;
  wire v9ed464;
  wire v9ed465;
  wire v9ed466;
  wire v9ed467;
  wire v9ed468;
  wire v9ed469;
  wire v9ed46a;
  wire v9ed46b;
  wire v9ed46c;
  wire v9ed46d;
  wire v9ed46e;
  wire v9ed46f;
  wire v9ed470;
  wire v9ed471;
  wire v9ed472;
  wire v9ed473;
  wire v9ed474;
  wire v9ed475;
  wire v9ed476;
  wire v9ed477;
  wire v9ed478;
  wire v9ed479;
  wire v9ed47a;
  wire v9ed47b;
  wire v9ed47c;
  wire v9ed47d;
  wire v9ed47e;
  wire v9ed47f;
  wire v9ed480;
  wire v9ed481;
  wire v9ed482;
  wire v9ed483;
  wire v9ed484;
  wire v9ed485;
  wire v9ed486;
  wire v9ed487;
  wire v9ed488;
  wire v9ed489;
  wire v9ed48a;
  wire v9ed48b;
  wire v9ed48c;
  wire v9ed48d;
  wire v9ed48e;
  wire v9ed48f;
  wire v9ed490;
  wire v9ed491;
  wire v9ed492;
  wire v9ed493;
  wire v9ed494;
  wire v9ed495;
  wire v9ed496;
  wire v9ed497;
  wire v9ed498;
  wire v9ed499;
  wire v9ed49a;
  wire v9ed49b;
  wire v9ed49c;
  wire v9ed49d;
  wire v9ed49e;
  wire v9ed49f;
  wire v9ed4a0;
  wire v9ed4a1;
  wire v9ed4a2;
  wire v9ed4a3;
  wire v9ed4a4;
  wire v9ed4a5;
  wire v9ed4a6;
  wire v9ed4a7;
  wire v845668;
  wire v9ed4a8;
  wire v9ed4a9;
  wire v9ed4aa;
  wire v9ed4ab;
  wire v9ed4ac;
  wire v9ed4ad;
  wire v9ed4ae;
  wire v9ed4af;
  wire v9ed4b0;
  wire v9ed4b1;
  wire v9ed4b2;
  wire v9ed4b3;
  wire v9ed4b4;
  wire v9ed4b5;
  wire v9ed4b6;
  wire v9ed4b7;
  wire v9ed4b8;
  wire v9ed4b9;
  wire v9ed4ba;
  wire v9ed4bb;
  wire v9ed4bc;
  wire v9ed4bd;
  wire v9ed4be;
  wire v9ed4bf;
  wire v9ed4c0;
  wire v9ed4c1;
  wire v9ed4c2;
  wire v9ed4c3;
  wire v9ed4c4;
  wire v9ed4c5;
  wire v9ed4c6;
  wire v9ed4c7;
  wire v9ed4c8;
  wire v9ed4c9;
  wire v9ed4ca;
  wire v9ed4cb;
  wire v9ed4cc;
  wire v9ed4cd;
  wire v9ed4ce;
  wire v9ed4cf;
  wire v9ed4d0;
  wire v9ed4d1;
  wire v9ed4d2;
  wire v9ed4d3;
  wire v9ed4d4;
  wire v9ed4d5;
  wire v9ed4d6;
  wire v9ed4d7;
  wire v9ed4d8;
  wire v9ed4d9;
  wire v9ed4da;
  wire v9ed4db;
  wire v9ed4dc;
  wire v9ed4dd;
  wire v9ed4de;
  wire v9ed4df;
  wire v9ed4e0;
  wire v9ed4e1;
  wire v9ed4e2;
  wire v9ed4e3;
  wire v9ed4e4;
  wire v9ed4e5;
  wire v9ed4e6;
  wire v9ed4e7;
  wire v9ed4e8;
  wire v9ed4e9;
  wire v9ed4ea;
  wire v9ed4eb;
  wire v9ed4ec;
  wire v9ed4ed;
  wire v9ed4ee;
  wire v9ed4ef;
  wire v9ed4f0;
  wire v9ed4f1;
  wire v9ed4f5;
  wire v9ed4f6;
  wire v9ed4f7;
  wire v9ed4f8;
  wire v9ed4f9;
  wire v9ed4fa;
  wire v9ed4fb;
  wire v9ed4fc;
  wire v9ed4fd;
  wire v9ed4fe;
  wire v9ed4ff;
  wire v9ed500;
  wire v9ed501;
  wire v9ed50b;
  wire v9ed520;
  wire v9ed521;
  wire v9ed522;
  wire v9ed52c;
  wire v9ed52d;
  wire v9ed52e;
  wire v9ed52f;
  wire v9ed530;
  wire v9ed531;
  wire v9ed532;
  wire v9ed533;
  wire v9ed567;
  wire v9ed568;
  wire v9ed56a;
  wire v9ed56e;
  wire v9ecda3;
  wire v9ecda4;
  wire v9ecda5;
  wire v9ecda6;
  wire v9ecda7;
  wire v9ecda8;
  wire v9ecda9;
  wire v84564b;
  wire v9d2662;
  wire v9d2663;
  wire v9d2664;
  wire v9d2665;
  wire v9d2666;
  wire v9d2667;
  wire v9d2668;
  wire v9d2669;
  wire v9d266a;
  wire v9d266b;
  wire v9d266c;
  wire v9d266d;
  wire v9d266e;
  wire v9d266f;
  wire v9d2670;
  wire v845647;
  wire v9d2671;
  wire v9d2672;
  wire v9d2673;
  wire v9d2674;
  wire v9d2675;
  wire v9d2676;
  wire v9d2677;
  wire v9d2678;
  wire v9d2679;
  wire v9d267a;
  wire v9d267b;
  wire v9d267c;
  wire v9d267d;
  wire v9d267e;
  wire v9d267f;
  wire v9d2680;
  wire v9d2681;
  wire v9d2682;
  wire v9d2683;
  wire v9d2684;
  wire v9d2685;
  wire v9d2686;
  wire v9d2687;
  wire v9d2688;
  wire v9d2689;
  wire v9d268a;
  wire v9d268b;
  wire v9d268c;
  wire v9d268d;
  wire v9d268e;
  wire v9d268f;
  wire v9d2690;
  wire v9d2691;
  wire v9d2692;
  wire v9d2693;
  wire v9d2694;
  wire v9d2695;
  wire v9d2696;
  wire v9d2697;
  wire v9d2698;
  wire v9d2699;
  wire v9d269a;
  wire v9d269b;
  wire v9d269c;
  wire v9d269d;
  wire v9d269e;
  wire v9d269f;
  wire v9d26a0;
  wire v9d26a1;
  wire v9d26a2;
  wire v9d26a3;
  wire v845641;
  wire v9d26a4;
  wire v9d26a5;
  wire v9d26a6;
  wire v9d26a7;
  wire v9d26a8;
  wire v9d26a9;
  wire v9d26aa;
  wire v9d26ab;
  wire v9d26ac;
  wire v9d26ad;
  wire v9d26ae;
  wire v9d26af;
  wire v9d26b0;
  wire v9d26b1;
  wire v9d26b2;
  wire v9d26b3;
  wire v9d26b4;
  wire v9d26b5;
  wire v9d26b6;
  wire v9d26b7;
  wire v9d26b8;
  wire v9d26b9;
  wire v9d26ba;
  wire v9d26bb;
  wire v9d26bc;
  wire v9d26bd;
  wire v9d26be;
  wire v9d26bf;
  wire v9d26c0;
  wire v9d26c1;
  wire v9d26c2;
  wire v9d26c3;
  wire v9d26c4;
  wire v9d26c5;
  wire v9d26c6;
  wire v9d26c7;
  wire v9d26c8;
  wire v9d26c9;
  wire v9d26ca;
  wire v9d26cb;
  wire v9d26cc;
  wire v9d26cd;
  wire v9d26ce;
  wire v9d26cf;
  wire v9d26d0;
  wire v9d26d1;
  wire v9d26d2;
  wire v9d26d3;
  wire v9d26d4;
  wire v9d26d5;
  wire v9d26d6;
  wire v9d26d7;
  wire v9d26d8;
  wire v9d26d9;
  wire v9d26da;
  wire v9d26db;
  wire v9d26dc;
  wire v9d26dd;
  wire v9d26de;
  wire v9d26df;
  wire v9d26e0;
  wire v9d26e1;
  wire v9d26e2;
  wire v9d26e3;
  wire v9d26e4;
  wire v9d26e5;
  wire v9d26e6;
  wire v9d26e8;
  wire v9d26e9;
  wire v9d26ea;
  wire v9d26eb;
  wire v9d26ec;
  wire v9d26ed;
  wire v9d26ee;
  wire v9d26ef;
  wire v9d26f0;
  wire v9d26f1;
  wire v9d26f2;
  wire v9d26f4;
  wire v9d26f5;
  wire v9d26f6;
  wire v9d26f7;
  wire v9d26f8;
  wire v9d26f9;
  wire v9d26fa;
  wire v9d26fb;
  wire v9d26fc;
  wire v9d26fd;
  wire v9d26fe;
  wire v9d26ff;
  wire v9d2700;
  wire v9d2701;
  wire v9d2702;
  wire v9d2703;
  wire v9d2704;
  wire v9d2705;
  wire v9d2706;
  wire v9d2707;
  wire v9d2708;
  wire v9d2709;
  wire v9d270a;
  wire v9d270b;
  wire v9d271a;
  wire v9d271b;
  wire v9d271c;
  wire v9d271d;
  wire v9d271e;
  wire v9d271f;
  wire v9d2720;
  wire v9d2721;
  wire v9d2722;
  wire v9d2723;
  wire v9d2724;
  wire v9d2725;
  wire v9d2726;
  wire v9d2727;
  wire v9d2728;
  wire v9d2729;
  wire v9d272a;
  wire v9d272b;
  wire v9d272c;
  wire v9d272d;
  wire v9d272e;
  wire v9d272f;
  wire v9d2730;
  wire v9d2732;
  wire v9d2733;
  wire v9d2734;
  wire v9d2735;
  wire v9d2736;
  wire v9d2737;
  wire v9d2738;
  wire v9d2739;
  wire v9d273a;
  wire v9d273b;
  wire v9d273c;
  wire v9d273d;
  wire v9d273e;
  wire v9d2746;
  wire v9d2747;
  wire v9d2748;
  wire v9d2749;
  wire v9d274a;
  wire v9d274b;
  wire v9d274c;
  wire v9d274d;
  wire v9d274e;
  wire v9d274f;
  wire v9d2750;
  wire v9d2751;
  wire v9d2752;
  wire v9d2753;
  wire v9d2754;
  wire v9d2755;
  wire v9d2756;
  wire v9d2757;
  wire v9d2758;
  wire v9d2759;
  wire v9d275a;
  wire v9d275b;
  wire v9d275c;
  wire v9d275d;
  wire v9d275e;
  wire v9d275f;
  wire v9d2760;
  wire v9d2761;
  wire v9d2762;
  wire v9d2763;
  wire v9d2764;
  wire v9d2765;
  wire v9d2766;
  wire v9d2767;
  wire v9d2768;
  wire v9d2769;
  wire v9d276a;
  wire v9d276b;
  wire v9d276c;
  wire v9d276d;
  wire v9d276e;
  wire v9d276f;
  wire v9d2770;
  wire v9d2771;
  wire v9d2772;
  wire v9d2773;
  wire v9d2774;
  wire v9d2775;
  wire v9d2776;
  wire v9d2777;
  wire v9d2778;
  wire v9d2779;
  wire v9d277a;
  wire v9d277b;
  wire v9d277c;
  wire v9d277d;
  wire v9d277e;
  wire v9d277f;
  wire v9d2780;
  wire v9d2781;
  wire v9d2782;
  wire v9d2783;
  wire v9d2784;
  wire v9d2785;
  wire v9d2786;
  wire v9d2787;
  wire v9d2788;
  wire v9d2789;
  wire v9d278a;
  wire v9d278b;
  wire v9d278c;
  wire v9d278d;
  wire v9d278e;
  wire v9d278f;
  wire v9d2790;
  wire v9d2791;
  wire v9d2792;
  wire v9d2793;
  wire v9d2794;
  wire v9d2795;
  wire v9d2796;
  wire v9d2797;
  wire v9d2798;
  wire v9d2799;
  wire v9d279a;
  wire v9d279b;
  wire v9d279c;
  wire v9d279d;
  wire v9d279e;
  wire v9d279f;
  wire v9d27a0;
  wire v9d27a1;
  wire v9d27a2;
  wire v9d27a3;
  wire v9d27a4;
  wire v9d27a5;
  wire v9d27a6;
  wire v9d27a7;
  wire v9d27a8;
  wire v9d27a9;
  wire v9d27aa;
  wire v9d27ab;
  wire v9d27ac;
  wire v9d27ad;
  wire v9d27ae;
  wire v9d27af;
  wire v9d27b0;
  wire v9d27b1;
  wire v9d27b2;
  wire v9d27b3;
  wire v9d27b4;
  wire v9d27b5;
  wire v9d27b6;
  wire v9d27b7;
  wire v9d27b8;
  wire v9d27b9;
  wire v9d27ba;
  wire v9d27bb;
  wire v9d27bc;
  wire v9d27bd;
  wire v9d27be;
  wire v9d27bf;
  wire v9d27c0;
  wire v9d27c1;
  wire v9d27c2;
  wire v9d27c3;
  wire v9d27c4;
  wire v9d27c5;
  wire v9d27c6;
  wire v9d27c7;
  wire v9bae78;
  wire v9bae79;
  wire v9bae7a;
  wire v9bae7b;
  wire v9bae7c;
  wire v9bae7d;
  wire v9bae7e;
  wire v9bae7f;
  wire v9bae80;
  wire v9bae81;
  wire v9bae82;
  wire v9bae83;
  wire v9bae84;
  wire v9bae85;
  wire v9bae86;
  wire v9bae87;
  wire v9bae88;
  wire v9bae89;
  wire v9bae8a;
  wire v9bae8b;
  wire v9bae8e;
  wire v9bae8f;
  wire v9bae90;
  wire v9bae92;
  wire v9bae93;
  wire v9bae94;
  wire v9bae95;
  wire v9bae96;
  wire v9bae97;
  wire v9bae98;
  wire v9bae99;
  wire v9bae9a;
  wire v9bae9d;
  wire v9bae9e;
  wire v9bae9f;
  wire v84565a;
  wire v9baea0;
  wire v9baea1;
  wire v9baea2;
  wire v9baea3;
  wire v9baea4;
  wire v9baea5;
  wire v9baea6;
  wire v9baea7;
  wire v9baea8;
  wire v9baea9;
  wire v9baeaa;
  wire v9baeab;
  wire v9baeac;
  wire v9baead;
  wire v9baeae;
  wire v9baeaf;
  wire v9baeb0;
  wire v9baeb1;
  wire v9baeb2;
  wire v9baeb3;
  wire v9baeb4;
  wire v9baeb5;
  wire v9baec7;
  wire v9baec8;
  wire v9baec9;
  wire v9baeca;
  wire v9baecb;
  wire v9baecc;
  wire v9baeee;
  wire v9baeef;
  wire v9baef0;
  wire v9baef1;
  wire v9baef2;
  wire v9baef3;
  wire v9baef4;
  wire v9baef5;
  wire v9baef6;
  wire v9baef7;
  wire v9baef8;
  wire v9baef9;
  wire v9baefa;
  wire v9baefb;
  wire v9baefc;
  wire v9baefd;
  wire v9baefe;
  wire v9baeff;
  wire v9baf00;
  wire v9baf01;
  wire v9baf02;
  wire v9baf03;
  wire v9baf04;
  wire v9baf05;
  wire v9baf06;
  wire v9baf07;
  wire v9baf08;
  wire v9baf09;
  wire v9baf0a;
  wire v9baf0b;
  wire v9baf0c;
  wire v9baf0d;
  wire v9baf0e;
  wire v9baf0f;
  wire v9baf10;
  wire v9baf11;
  wire v9baf12;
  wire v9baf13;
  wire v9baf14;
  wire v9baf15;
  wire a2fb4b;
  wire a2fb4c;
  wire v9baf17;
  wire v9baf18;
  wire v9baf19;
  wire v9baf1a;
  wire a2f895;
  wire v9baf1b;
  wire v9baf1c;
  wire v9baf1d;
  wire v9baf1e;
  wire v9baf1f;
  wire v9baf20;
  wire v9baf21;
  wire v9baf22;
  wire v9baf23;
  wire v9baf24;
  wire v9baf25;
  wire v9baf26;
  wire v9baf27;
  wire v9baf28;
  wire v9baf29;
  wire v9baf2a;
  wire a2fb4d;
  wire v9baf2b;
  wire v9baf2c;
  wire v9baf2d;
  wire v9baf2e;
  wire v9baf2f;
  wire v9baf30;
  wire v9baf31;
  wire v9baf32;
  wire v9baf34;
  wire v9baf35;
  wire v9baf36;
  wire v9baf37;
  wire v9baf38;
  wire v9baf3a;
  wire v9baf3b;
  wire v9baf3c;
  wire v9baf3d;
  wire v9baf3e;
  wire v9baf3f;
  wire v9baf40;
  wire v9baf41;
  wire v9baf42;
  wire v9baf43;
  wire v9baf44;
  wire v9baf45;
  wire v9baf46;
  wire v9baf47;
  wire v9baf48;
  wire v9baf49;
  wire v9baf4a;
  wire v9baf4b;
  wire v9baf4c;
  wire v9baf4d;
  wire v9baf4e;
  wire v9baf4f;
  wire v9baf50;
  wire v9baf51;
  wire v9baf52;
  wire v9baf53;
  wire v9baf54;
  wire v9baf55;
  wire v9baf56;
  wire v9baf57;
  wire v9baf58;
  wire v9baf59;
  wire v9baf5a;
  wire v9baf5b;
  wire v9baf5c;
  wire v9baf5d;
  wire v9baf5e;
  wire v9baf5f;
  wire v9baf60;
  wire v9baf61;
  wire v9baf62;
  wire v9baf63;
  wire v9baf64;
  wire v9baf65;
  wire v9baf66;
  wire v9baf67;
  wire v9baf68;
  wire v9baf69;
  wire v9baf6a;
  wire v9baf6b;
  wire v9baf6d;
  wire v9baf6e;
  wire v9baf6f;
  wire v9baf70;
  wire v9baf71;
  wire v9baf72;
  wire v9baf73;
  wire v9baf74;
  wire v9baf75;
  wire v9baf76;
  wire v9baf77;
  wire v9baf78;
  wire v9baf79;
  wire v9baf7a;
  wire v9baf7b;
  wire v9baf7c;
  wire v9baf7d;
  wire v9baf7e;
  wire v9baf7f;
  wire v9baf80;
  wire v9baf81;
  wire v9baf82;
  wire v9baf83;
  wire v9baf84;
  wire v9baf85;
  wire v9baf86;
  wire v9baf87;
  wire v9baf88;
  wire v9baf89;
  wire v9baf8a;
  wire v9baf8b;
  wire v9baf8c;
  wire v9baf8d;
  wire v9baf8e;
  wire v9baf8f;
  wire v9baf90;
  wire v9baf92;
  wire v9baf93;
  wire v9baf94;
  wire v9baf95;
  wire v9baf96;
  wire v9baf97;
  wire v9baf98;
  wire v9baf99;
  wire v9baf9a;
  wire v9baf9b;
  wire v9baf9c;
  wire v9baf9d;
  wire v9baf9e;
  wire v9baf9f;
  wire v9bafa0;
  wire v9bafa1;
  wire v845654;
  wire v9b40c0;
  wire v9b40c1;
  wire v9b40c2;
  wire v9b40c3;
  wire v9b40c4;
  wire v9b40c5;
  wire v9b40c6;
  wire v9b40cc;
  wire v9b40cd;
  wire v9b40d0;
  wire v9b40db;
  wire v9b40dc;
  wire v9b40dd;
  wire v9b40de;
  wire v898b4e;
  wire v854662;
  wire v9adbe6;
  wire a2bb5d;
  wire v9adbe7;
  wire v9adbe8;
  wire v9adbe9;
  wire v9adbea;
  wire v9adbeb;
  wire v9adbec;
  wire v8543f4;
  wire v9adbed;
  wire v9adbee;
  wire v9adbef;
  wire v9adbf0;
  wire v9adbf1;
  wire v9adbf2;
  wire v9adbf3;
  wire v9adbf4;
  wire v9adbf5;
  wire v9adbf6;
  wire v9adbf7;
  wire v9adbf8;
  wire v9adbf9;
  wire v9adbfa;
  wire v9adbfb;
  wire v9adbfc;
  wire v9adbfd;
  wire v8ec3e4;
  wire v9adbfe;
  wire v9adbff;
  wire v9adc00;
  wire v9adc01;
  wire v9adc02;
  wire v9adc03;
  wire v9adc04;
  wire v9adc05;
  wire v9adc06;
  wire v9adc07;
  wire v9adc08;
  wire v9adc09;
  wire v9adc0a;
  wire v9adc0b;
  wire v9adc0c;
  wire v9adc0d;
  wire v9adc0e;
  wire v9adc0f;
  wire v9adc10;
  wire v9adc11;
  wire v9adc12;
  wire v9adc13;
  wire v9adc14;
  wire v9adc15;
  wire v9adc16;
  wire v9adc17;
  wire v9adc18;
  wire v9adc19;
  wire v9adc1a;
  wire v9adc1b;
  wire v9adc1c;
  wire v9adc1d;
  wire v9adc1e;
  wire v9adc1f;
  wire v9adc20;
  wire v9adc21;
  wire v9adc22;
  wire v9adc23;
  wire v9adc24;
  wire v9adc25;
  wire v9adc26;
  wire v9adc27;
  wire v9adc28;
  wire v9adc29;
  wire v9adc2a;
  wire v9adc2b;
  wire v9adc2c;
  wire v9adc2d;
  wire v9adc2e;
  wire v9adc2f;
  wire v9adc30;
  wire v9adc31;
  wire v9adc32;
  wire v9adc33;
  wire v9adc34;
  wire v9adc35;
  wire v9adc36;
  wire v9adc37;
  wire v9adc38;
  wire v9adc39;
  wire v9adc3a;
  wire v9adc3b;
  wire v9adc3c;
  wire v9adc3d;
  wire v9adc3e;
  wire v9adc3f;
  wire v9adc40;
  wire v9adc41;
  wire v9adc42;
  wire v9adc43;
  wire v9adc44;
  wire v9adc45;
  wire v9adc46;
  wire v9adc47;
  wire v9adc48;
  wire v9adc49;
  wire v9adc4a;
  wire v9adc4b;
  wire v9adc4c;
  wire v9adc4d;
  wire v9adc4e;
  wire v9adc4f;
  wire v9adc50;
  wire v9adc51;
  wire v9adc52;
  wire v9adc53;
  wire v9adc54;
  wire v9adc55;
  wire v9adc56;
  wire v9adc57;
  wire v9adc58;
  wire v9adc59;
  wire v9adc5a;
  wire v9adc5b;
  wire v9adc5c;
  wire v9adc5d;
  wire v9adc5e;
  wire v9adc5f;
  wire v9adc60;
  wire v9adc61;
  wire v9adc62;
  wire v9adc63;
  wire v9adc64;
  wire v9adc65;
  wire v9adc66;
  wire v9adc67;
  wire v9adc68;
  wire v9adc69;
  wire v9adc6a;
  wire v9adc6b;
  wire v9adc6c;
  wire v9adc6d;
  wire v9adc6e;
  wire v9adc6f;
  wire v9adc70;
  wire v9adc71;
  wire v9adc72;
  wire v9adc73;
  wire v9adc74;
  wire v9adc75;
  wire v9adc76;
  wire v9adc77;
  wire v9adc78;
  wire v9adc79;
  wire v9adc7a;
  wire v9adc7b;
  wire v9adc7c;
  wire v9adc7d;
  wire v9adc7e;
  wire v9adc7f;
  wire v9adc80;
  wire v9adc81;
  wire v9adc82;
  wire v9adc83;
  wire v9adc84;
  wire v9adc85;
  wire v9adc86;
  wire v9adc87;
  wire v9adc88;
  wire v9adc89;
  wire v9adc8a;
  wire v9adc8b;
  wire v9adc8c;
  wire v9adc8d;
  wire v9adc8e;
  wire v9adc8f;
  wire v9adc90;
  wire v9adc91;
  wire v9adc92;
  wire v9adc93;
  wire v9adc94;
  wire v9adc95;
  wire v9adc96;
  wire v9adc97;
  wire v9adc98;
  wire v9adc99;
  wire v9adc9a;
  wire v9adc9b;
  wire v9adc9c;
  wire v9adc9d;
  wire v9adc9e;
  wire v9adc9f;
  wire v9adca0;
  wire v9adca1;
  wire v9adca2;
  wire v9adca3;
  wire v9adca4;
  wire v9adca5;
  wire v9adca6;
  wire v9adca7;
  wire v9adca8;
  wire v9adca9;
  wire v9adcaa;
  wire v9adcab;
  wire v9adcac;
  wire v9adcad;
  wire v9adcae;
  wire v9adcaf;
  wire v9adcb0;
  wire v9adcb1;
  wire v9adcb2;
  wire v9adcb3;
  wire v9adcb4;
  wire v9adcb5;
  wire v9adcb6;
  wire v9adcb7;
  wire v9adcb8;
  wire v9adcb9;
  wire v9adcba;
  wire v9adcbb;
  wire v9adcbc;
  wire v9adcbd;
  wire v9adcbe;
  wire v9adcbf;
  wire v9adcc0;
  wire v9adcc1;
  wire v9adcc2;
  wire v9adcc3;
  wire v9adcc4;
  wire v9adcc5;
  wire v9adcc6;
  wire v9adcc7;
  wire v9adcc8;
  wire v9adcc9;
  wire v9adcca;
  wire v9adccb;
  wire v9adccc;
  wire v9adccd;
  wire v9adcce;
  wire v9adccf;
  wire v9adcd0;
  wire v9adcd1;
  wire v9adcd2;
  wire v9adcd3;
  wire v9adcd4;
  wire v9adcd5;
  wire v9adcd6;
  wire v9adcd7;
  wire v9adcd8;
  wire v9adcd9;
  wire v9adcda;
  wire v9adcdb;
  wire v9adcdc;
  wire v9adcdd;
  wire v9adcde;
  wire v9adcdf;
  wire v9adce0;
  wire v9adce1;
  wire v9adce2;
  wire v9adce3;
  wire v9adce4;
  wire v9adce5;
  wire v9adce6;
  wire v9adce7;
  wire v9adce8;
  wire v9adce9;
  wire v9adcea;
  wire v9adceb;
  wire v9adcec;
  wire v9adced;
  wire v9adcee;
  wire v9adcef;
  wire v9adcf0;
  wire v9adcf1;
  wire v9adcf2;
  wire v9adcf3;
  wire v9adcf4;
  wire v9adcf5;
  wire v9adcf6;
  wire v9adcf7;
  wire v9adcf8;
  wire v9a6a94;
  wire v9a6a95;
  wire v9a6a96;
  wire v9a6a97;
  wire v9a6a98;
  wire v9a6a99;
  wire v9a6a9a;
  wire v9a6a9b;
  wire v9a6a9c;
  wire v9a6a9d;
  wire v9a6a9e;
  wire v9a6a9f;
  wire v9a6aa0;
  wire v9a6aa1;
  wire v9a6aa2;
  wire v9a6aa3;
  wire v9a6aa4;
  wire v9a6aa5;
  wire v9a6aa6;
  wire v9a6aa7;
  wire v9a6aa8;
  wire v9a6aa9;
  wire v9a6aaa;
  wire v9a6aab;
  wire v9a6aac;
  wire v9a6aad;
  wire v9a6aae;
  wire v9a6aaf;
  wire v9a6ab0;
  wire v9a6ab1;
  wire v9a6ab2;
  wire v9a6ab3;
  wire v9a6ab4;
  wire v9a6ab5;
  wire v9a6ab6;
  wire v9a6ab7;
  wire v9a6ab8;
  wire v9a6ab9;
  wire v9a6aba;
  wire v9a6abb;
  wire v9a6abc;
  wire v9a6abd;
  wire v9a6abe;
  wire v9a6abf;
  wire v9a6ac0;
  wire v9a6ac1;
  wire v9a6ac2;
  wire v9a6ac3;
  wire v9a6ac4;
  wire v9a6ac5;
  wire v9a6ac6;
  wire v9a6ac7;
  wire v9a6ac8;
  wire v9a6ac9;
  wire v9a6aca;
  wire v9a6acb;
  wire v9a6acc;
  wire v9a6acd;
  wire v9a6ace;
  wire v9a6acf;
  wire v9a6ad0;
  wire v9a6ad1;
  wire v9a6ad2;
  wire v9a6ad3;
  wire v9a6ad4;
  wire v9a6ad5;
  wire v9a6ad6;
  wire v9a6ad7;
  wire v9a6ad8;
  wire v9a6ad9;
  wire v9a6ada;
  wire v9a6adb;
  wire v9a6adc;
  wire v9a6add;
  wire v9a6ade;
  wire v9a6adf;
  wire v9a6ae0;
  wire v9a6ae1;
  wire v9a6ae2;
  wire v9a6ae3;
  wire v99989c;
  wire v99989d;
  wire v99989e;
  wire v99989f;
  wire v9998a0;
  wire v9998a1;
  wire v9998a2;
  wire v9998a3;
  wire v9998a4;
  wire v9998a5;
  wire v9998a6;
  wire v9998a7;
  wire v9998a8;
  wire v9998a9;
  wire v9998aa;
  wire v9998ab;
  wire v9998ac;
  wire v9998ad;
  wire v9998ae;
  wire v9998af;
  wire v9998cd;
  wire v9998ce;
  wire v9998cf;
  wire v9998d3;
  wire v9998d4;
  wire v9998d5;
  wire v9998d6;
  wire v9998d7;
  wire v9998d8;
  wire v9998d9;
  wire v9998da;
  wire v9998db;
  wire v9998dc;
  wire v9998dd;
  wire v9998de;
  wire v9998df;
  wire v9998e0;
  wire v9998e1;
  wire v9998e2;
  wire v9998e3;
  wire v9998e4;
  wire v9998e5;
  wire v9998e6;
  wire v9998e7;
  wire v9998e8;
  wire v9998e9;
  wire v9998ea;
  wire v9998eb;
  wire v9998ec;
  wire v9998ed;
  wire v9998ee;
  wire v9998ef;
  wire v9998f0;
  wire v9998f1;
  wire v9998f2;
  wire v9998f3;
  wire v9998f4;
  wire v9998f5;
  wire v9998f6;
  wire v9998f7;
  wire v9998f8;
  wire v9998f9;
  wire v9998fa;
  wire v9998fb;
  wire v9998fc;
  wire v9998fd;
  wire v9998fe;
  wire v9998ff;
  wire v999900;
  wire v999901;
  wire v999902;
  wire v999903;
  wire v999904;
  wire v999905;
  wire v999906;
  wire v999907;
  wire v999908;
  wire v999909;
  wire v99990a;
  wire v99990b;
  wire v99990c;
  wire v99990d;
  wire v99990e;
  wire v99990f;
  wire v999910;
  wire v999911;
  wire v999912;
  wire v999913;
  wire v999914;
  wire v999915;
  wire v999916;
  wire v999917;
  wire v999918;
  wire v999919;
  wire v99991a;
  wire v99991b;
  wire v99991c;
  wire v99991d;
  wire v99991e;
  wire v99991f;
  wire v999920;
  wire v999921;
  wire v999922;
  wire v999923;
  wire v999924;
  wire v999925;
  wire v999926;
  wire v999927;
  wire v999928;
  wire v999929;
  wire v99992a;
  wire v99992b;
  wire v99992c;
  wire v99992d;
  wire v99992e;
  wire v99992f;
  wire v999930;
  wire v999931;
  wire v999932;
  wire v999933;
  wire v999934;
  wire v999935;
  wire v999936;
  wire v999937;
  wire v999938;
  wire v999939;
  wire v99993a;
  wire v99993b;
  wire v99993c;
  wire v99993d;
  wire v99993e;
  wire v99993f;
  wire v999940;
  wire v999969;
  wire v99996a;
  wire v99996b;
  wire v99996c;
  wire v99996d;
  wire v99996e;
  wire v99996f;
  wire v999970;
  wire v999971;
  wire v999972;
  wire v999973;
  wire v999974;
  wire v999975;
  wire v999976;
  wire v999977;
  wire v999978;
  wire v999979;
  wire v99997a;
  wire v99997b;
  wire v99997c;
  wire v99997d;
  wire v99997e;
  wire v99997f;
  wire v999980;
  wire v999981;
  wire v999982;
  wire v999983;
  wire v999984;
  wire v999985;
  wire v999986;
  wire v999987;
  wire v999988;
  wire v999989;
  wire v99998a;
  wire v99998b;
  wire v99998c;
  wire v99998d;
  wire v99998e;
  wire v99999a;
  wire v99999b;
  wire v99999c;
  wire v99999d;
  wire v99999e;
  wire v99999f;
  wire v9999a0;
  wire v9999a1;
  wire v9999a2;
  wire v9999a3;
  wire v9999a4;
  wire v9999a5;
  wire v9999a6;
  wire v9999a7;
  wire v9999a8;
  wire v9999a9;
  wire v9999aa;
  wire v9999ab;
  wire v9999ac;
  wire v9999ad;
  wire v9999ae;
  wire v9999af;
  wire v9999b0;
  wire v9999b1;
  wire v9999b2;
  wire v9999b3;
  wire v9999b4;
  wire v9999b5;
  wire v9999b6;
  wire v9999b7;
  wire v9999b8;
  wire v9999b9;
  wire v9999ba;
  wire v9999bb;
  wire v9999bc;
  wire v9999bd;
  wire v9999be;
  wire v9999bf;
  wire v9999c0;
  wire v9999c1;
  wire v9999c2;
  wire v9999c3;
  wire v9999c4;
  wire v9999c5;
  wire v9999c6;
  wire v9999c7;
  wire v9999c8;
  wire v9999c9;
  wire v9999ca;
  wire v9999cb;
  wire v9999d0;
  wire v9999d1;
  wire v9999d2;
  wire v9999d3;
  wire v9999d4;
  wire v9999d5;
  wire v9999d6;
  wire v9999d7;
  wire v9999d8;
  wire v9999d9;
  wire v9999da;
  wire v9999db;
  wire v9999dc;
  wire v9999dd;
  wire v9999de;
  wire v9999df;
  wire v9999e0;
  wire v9999e1;
  wire v9999e2;
  wire v9999e3;
  wire v9999e4;
  wire v9999e5;
  wire v9999e6;
  wire v9999e7;
  wire v9999e8;
  wire v9999e9;
  wire v9999ea;
  wire v9999eb;
  wire v9999ec;
  wire v9999ed;
  wire v9999ee;
  wire v9999ef;
  wire v9999f0;
  wire v9999f1;
  wire v99654f;
  wire v996550;
  wire v996551;
  wire v996552;
  wire v996553;
  wire v996554;
  wire v996555;
  wire v996556;
  wire v996557;
  wire v996558;
  wire v996559;
  wire v99655a;
  wire v99655b;
  wire v99655c;
  wire v99655d;
  wire v99655e;
  wire v99655f;
  wire v996560;
  wire v996561;
  wire v996562;
  wire v996563;
  wire v996564;
  wire v996565;
  wire v996566;
  wire v996567;
  wire v996568;
  wire v996569;
  wire v99656a;
  wire v99656b;
  wire v99656c;
  wire v99656d;
  wire v99656e;
  wire v99656f;
  wire v996570;
  wire v996571;
  wire v996572;
  wire v996573;
  wire v996574;
  wire v996575;
  wire v996576;
  wire v996577;
  wire v996578;
  wire v996579;
  wire v99657a;
  wire v99657b;
  wire v99657c;
  wire v99657d;
  wire v99657e;
  wire v99657f;
  wire v996580;
  wire v996581;
  wire v996582;
  wire v996583;
  wire v996584;
  wire v996585;
  wire v996586;
  wire v996587;
  wire v996588;
  wire v996589;
  wire v99658a;
  wire v99658b;
  wire v99658c;
  wire v99658d;
  wire v99658e;
  wire v99658f;
  wire v996590;
  wire v996591;
  wire v996592;
  wire v996593;
  wire v996594;
  wire v996595;
  wire v996596;
  wire v996597;
  wire v996598;
  wire v996599;
  wire v99659a;
  wire v99659b;
  wire v99659c;
  wire v99659d;
  wire v99659e;
  wire v99659f;
  wire v9965a0;
  wire v9965a1;
  wire v9965a2;
  wire v9965a3;
  wire v9965a4;
  wire v9965a5;
  wire v9965a6;
  wire v9965a7;
  wire v9965a8;
  wire v9965a9;
  wire v9965aa;
  wire v9965ab;
  wire v9965ac;
  wire v9965ad;
  wire v9965ae;
  wire v9965af;
  wire v9965b0;
  wire v9965b1;
  wire v9965b2;
  wire v9965b3;
  wire v9965b4;
  wire v9965b5;
  wire v9965b6;
  wire v9965b7;
  wire v9965b8;
  wire v9965b9;
  wire v9965ba;
  wire v9965bb;
  wire v9965bc;
  wire v9965bd;
  wire v9965be;
  wire v9965bf;
  wire v9965c0;
  wire v9965c1;
  wire v9965c2;
  wire v9965c3;
  wire v9965c4;
  wire v9965c5;
  wire v9965c6;
  wire v9965c7;
  wire v9965c8;
  wire v9965c9;
  wire v9965ca;
  wire v9965cb;
  wire v9965cc;
  wire v9965cd;
  wire v9965ce;
  wire v9965cf;
  wire v9965d0;
  wire v9965d1;
  wire v9965d2;
  wire v9965d3;
  wire v98548f;
  wire v985490;
  wire v985491;
  wire v985492;
  wire v985493;
  wire v985494;
  wire v985495;
  wire v985496;
  wire v985497;
  wire v985498;
  wire v985499;
  wire v98549a;
  wire v98549b;
  wire v98549c;
  wire v98549d;
  wire v98549e;
  wire v98549f;
  wire v9854a0;
  wire v9854a1;
  wire v9854a2;
  wire v9854a3;
  wire v9854a4;
  wire v9854a5;
  wire v9854a6;
  wire v9854a7;
  wire v9854a8;
  wire v9854a9;
  wire v9854aa;
  wire v9854ab;
  wire v9854ac;
  wire v9854ad;
  wire v9854ae;
  wire v9854af;
  wire v9854b0;
  wire v9854b1;
  wire v9854b2;
  wire v9854b3;
  wire v9854b4;
  wire v9854b5;
  wire v9854b6;
  wire v9854b7;
  wire v9854b8;
  wire v9854b9;
  wire v9854ba;
  wire v9854bb;
  wire a3134e;
  wire a3134f;
  wire v9854bc;
  wire v9854bd;
  wire v9854be;
  wire v9854bf;
  wire v9854c0;
  wire v9854c1;
  wire v9854c2;
  wire v9854c3;
  wire v9854c4;
  wire v9854c5;
  wire v9854c6;
  wire v9854c7;
  wire v9854c8;
  wire v9854c9;
  wire v9854ca;
  wire v9854cb;
  wire v9854cc;
  wire v9854cd;
  wire v9854ce;
  wire v9854cf;
  wire v9854d0;
  wire v9854d1;
  wire v9854d2;
  wire v9854d3;
  wire v9854d4;
  wire v9854d5;
  wire v9854d6;
  wire v9854d7;
  wire v9854d8;
  wire v9854d9;
  wire v9854da;
  wire v9854db;
  wire v9854dc;
  wire v9854dd;
  wire v9854de;
  wire v9854df;
  wire v9854e0;
  wire v9854e1;
  wire v9854e2;
  wire v9854e3;
  wire v9854e4;
  wire v9854e5;
  wire v9854e6;
  wire v9854e7;
  wire v9854e8;
  wire v9854e9;
  wire v9854ea;
  wire v9854eb;
  wire v9854ec;
  wire v9854ed;
  wire v9854ee;
  wire v9854ef;
  wire v9854f0;
  wire v9854f1;
  wire v9854f2;
  wire v9854f3;
  wire v9854f4;
  wire v9854f5;
  wire v9854f6;
  wire v9854f7;
  wire v9854f8;
  wire v9854f9;
  wire v9854fa;
  wire v9854fb;
  wire v9854fc;
  wire v9854fd;
  wire v9854fe;
  wire v9854ff;
  wire v985500;
  wire v985501;
  wire v985502;
  wire v985503;
  wire v985504;
  wire v985505;
  wire v985506;
  wire v985507;
  wire v985508;
  wire v985509;
  wire v98550a;
  wire v98550b;
  wire v98550c;
  wire v98550d;
  wire v98550e;
  wire v98550f;
  wire v985510;
  wire v985511;
  wire v985512;
  wire v985513;
  wire v985514;
  wire v985515;
  wire v985516;
  wire v985517;
  wire v985518;
  wire v985519;
  wire v98551a;
  wire v98551b;
  wire v98551c;
  wire v98551d;
  wire v98551e;
  wire v98551f;
  wire v985520;
  wire v985521;
  wire v985522;
  wire v985523;
  wire v985524;
  wire v985525;
  wire v985526;
  wire v985527;
  wire v985528;
  wire v985529;
  wire v98552a;
  wire v98552b;
  wire v98552c;
  wire v98552d;
  wire v98552e;
  wire v98552f;
  wire v985530;
  wire v985531;
  wire v985532;
  wire v985533;
  wire v985534;
  wire v985535;
  wire v985536;
  wire v985537;
  wire v985538;
  wire v985539;
  wire v98553a;
  wire v98553b;
  wire v98553c;
  wire v98553d;
  wire v98553e;
  wire v98553f;
  wire v985540;
  wire v985541;
  wire v985542;
  wire v985543;
  wire v985544;
  wire v985545;
  wire v985546;
  wire v985547;
  wire v985548;
  wire v985549;
  wire v98554a;
  wire v98554b;
  wire v98554c;
  wire v98554d;
  wire v98554e;
  wire v98554f;
  wire v985550;
  wire v985551;
  wire v985552;
  wire v985553;
  wire v985554;
  wire v985555;
  wire v985556;
  wire v985557;
  wire v985558;
  wire v985559;
  wire v98555a;
  wire v98555b;
  wire v98555c;
  wire v98555e;
  wire v98555f;
  wire v985560;
  wire v985561;
  wire v985562;
  wire v985563;
  wire v985564;
  wire v985565;
  wire v985566;
  wire v985567;
  wire v985568;
  wire v985569;
  wire v98556a;
  wire v98556b;
  wire v98556c;
  wire v98556d;
  wire v98556e;
  wire v98556f;
  wire v985570;
  wire v985571;
  wire v985572;
  wire v985573;
  wire v985574;
  wire v985575;
  wire v985576;
  wire v985577;
  wire v985578;
  wire v985579;
  wire v98557a;
  wire v98557b;
  wire v98557c;
  wire v98557d;
  wire v98557e;
  wire v98557f;
  wire v985580;
  wire v985581;
  wire v985582;
  wire v985583;
  wire v985584;
  wire v985585;
  wire v985586;
  wire v985587;
  wire v985588;
  wire v985589;
  wire v98558a;
  wire v98558b;
  wire v98558c;
  wire v98558d;
  wire v98558e;
  wire v98558f;
  wire v985590;
  wire v985591;
  wire v985592;
  wire v985593;
  wire v985594;
  wire v985595;
  wire v985596;
  wire v985597;
  wire v985598;
  wire v985599;
  wire v98559a;
  wire v98559b;
  wire v98559c;
  wire v98559d;
  wire v98559e;
  wire v98559f;
  wire v9855a0;
  wire v9855a1;
  wire v9855a2;
  wire v9855a3;
  wire v9855a4;
  wire v9855a5;
  wire v9855a6;
  wire v9855a7;
  wire v9855a8;
  wire v9855a9;
  wire v9855aa;
  wire v9855ab;
  wire v9855ac;
  wire v9855ad;
  wire v9855ae;
  wire v9855af;
  wire v9855b0;
  wire v9855b1;
  wire v9855b2;
  wire v9855b3;
  wire v9855b4;
  wire v9855b5;
  wire v9855b6;
  wire v9855b7;
  wire v9855b8;
  wire v9855b9;
  wire v9855ba;
  wire v9855bb;
  wire v9855bc;
  wire v9855bd;
  wire v9855be;
  wire v9855bf;
  wire v9855c0;
  wire v9855c1;
  wire v9855c2;
  wire v9855c3;
  wire v9855c4;
  wire v9855c5;
  wire v9855c6;
  wire v9855c7;
  wire v9855c8;
  wire v9855c9;
  wire v9855ca;
  wire v9855cb;
  wire v9855cc;
  wire v9855cd;
  wire v9855ce;
  wire v9855cf;
  wire v9855d0;
  wire v9855d1;
  wire v9855d2;
  wire v9855d3;
  wire v9855d4;
  wire v9855d5;
  wire v9855d6;
  wire v9855d7;
  wire v9855d8;
  wire v9855d9;
  wire v9855da;
  wire v9855db;
  wire v9855dd;
  wire v9855de;
  wire v9855df;
  wire v9855e0;
  wire v9855e1;
  wire v9855e2;
  wire v9855e3;
  wire v9855e4;
  wire v9855e5;
  wire v9855e6;
  wire v9855e7;
  wire v9855e8;
  wire v9855e9;
  wire v9855ea;
  wire v9855eb;
  wire v9855ec;
  wire v9855ed;
  wire v9855ee;
  wire v9855ef;
  wire v9855f0;
  wire v9855f1;
  wire v9855f2;
  wire v9855f3;
  wire v9855f4;
  wire v9855f5;
  wire v9855f6;
  wire v9855f7;
  wire v9855f8;
  wire v9855f9;
  wire v9855fa;
  wire v9855fb;
  wire v9855fc;
  wire v9855fd;
  wire v9855fe;
  wire v9855ff;
  wire v985600;
  wire v985601;
  wire v985602;
  wire v985603;
  wire v985604;
  wire v985605;
  wire v985606;
  wire v985607;
  wire v985608;
  wire v985609;
  wire v98560a;
  wire v98560b;
  wire v98560c;
  wire v98560d;
  wire v98560e;
  wire v98560f;
  wire v985610;
  wire v985611;
  wire v985612;
  wire v985613;
  wire v985614;
  wire v985615;
  wire v985616;
  wire v985617;
  wire v985618;
  wire v985619;
  wire v98561a;
  wire v98561b;
  wire v98561c;
  wire v98561d;
  wire v98561e;
  wire v98561f;
  wire v985620;
  wire v985621;
  wire v985622;
  wire v985623;
  wire v985624;
  wire v985625;
  wire v985626;
  wire v985627;
  wire v985628;
  wire v985629;
  wire v98562a;
  wire v98562b;
  wire v98562c;
  wire v98562d;
  wire v98562e;
  wire v98562f;
  wire v985630;
  wire v985631;
  wire v985632;
  wire v985633;
  wire v985634;
  wire v985635;
  wire v985636;
  wire v985637;
  wire v985638;
  wire v985639;
  wire v98563a;
  wire v98563b;
  wire v98563c;
  wire v98563d;
  wire v98563e;
  wire v98563f;
  wire v985640;
  wire v985641;
  wire v985642;
  wire v985643;
  wire v985644;
  wire v985645;
  wire v985646;
  wire v985647;
  wire v985648;
  wire v985649;
  wire v98564a;
  wire v98564b;
  wire v98564c;
  wire v98564d;
  wire v98564e;
  wire v98564f;
  wire v984e52;
  wire v984e53;
  wire v984e54;
  wire v984e55;
  wire v984e56;
  wire v984e57;
  wire v984e58;
  wire v984e59;
  wire v984e5a;
  wire v984e5b;
  wire v984e5c;
  wire v984e5d;
  wire v984e5e;
  wire v984e5f;
  wire v984e60;
  wire v984e61;
  wire v984e62;
  wire v984e63;
  wire v984e64;
  wire v984e65;
  wire v984e66;
  wire v984e67;
  wire v984e68;
  wire v984e69;
  wire v984e6a;
  wire v984e6b;
  wire v984e6c;
  wire v984e6d;
  wire v984e6e;
  wire v984e6f;
  wire v984e70;
  wire v984e71;
  wire v984e72;
  wire v984e73;
  wire v984e74;
  wire v984e75;
  wire v984e76;
  wire v984e77;
  wire v984e78;
  wire v984ea4;
  wire v984ea5;
  wire v984ea6;
  wire v984ea7;
  wire v984ea8;
  wire v984ea9;
  wire v984eaa;
  wire v984eab;
  wire v984eac;
  wire v984ead;
  wire v984eae;
  wire v984eaf;
  wire v984eb0;
  wire v984eb1;
  wire v984eb2;
  wire v984eb3;
  wire v984eb4;
  wire v984eb5;
  wire v984eb6;
  wire v984eb7;
  wire v984eb8;
  wire v984eb9;
  wire v984eba;
  wire v984ebb;
  wire v984ebc;
  wire v984ebd;
  wire v984ebe;
  wire v984ebf;
  wire v984ec0;
  wire v984ec1;
  wire v984ec2;
  wire v984ec3;
  wire v984ec4;
  wire v984ec5;
  wire v984ec6;
  wire v984ec7;
  wire v984ec8;
  wire v984ec9;
  wire v984eca;
  wire v984ecb;
  wire v984ecc;
  wire v984ecd;
  wire v984ece;
  wire v984ecf;
  wire v984ed0;
  wire v984ed1;
  wire v984ed8;
  wire v984ed9;
  wire v984eda;
  wire v984edb;
  wire v984edc;
  wire v984edd;
  wire v984ede;
  wire v984edf;
  wire v984ee0;
  wire v984ee1;
  wire v984ee2;
  wire v984ee3;
  wire v984ee5;
  wire v984ee6;
  wire v984ee7;
  wire v984ee8;
  wire v984ee9;
  wire v984eea;
  wire v984eef;
  wire v984ef0;
  wire v984ef1;
  wire v984ef2;
  wire v984ef3;
  wire v984ef4;
  wire v984ef5;
  wire v984ef6;
  wire v984f20;
  wire v984f24;
  wire v984f25;
  wire v984f26;
  wire v984f27;
  wire v984f28;
  wire v984f29;
  wire v984f2b;
  wire v984f2c;
  wire v984f2d;
  wire v984f2e;
  wire v984f2f;
  wire v984f37;
  wire v984f38;
  wire v984f39;
  wire v984f3a;
  wire v984f3b;
  wire v984f3c;
  wire v984f3d;
  wire v984f3e;
  wire v984f3f;
  wire v984f40;
  wire v984f41;
  wire v984f42;
  wire v984f43;
  wire v984f44;
  wire v984f45;
  wire v984f46;
  wire v984f47;
  wire v984f48;
  wire v984f49;
  wire v984f4a;
  wire v984f4b;
  wire v984f4c;
  wire v984f4d;
  wire v984f4e;
  wire v984f4f;
  wire v984f50;
  wire v984f51;
  wire v984f52;
  wire v984f53;
  wire v984f54;
  wire v984f55;
  wire v984f56;
  wire v984f57;
  wire v984f58;
  wire v984f59;
  wire v984f5a;
  wire v984f5b;
  wire v984f5c;
  wire v984f5d;
  wire v984f5e;
  wire v984f5f;
  wire v984f60;
  wire v984f61;
  wire v984f62;
  wire v984f63;
  wire v984f64;
  wire v984f65;
  wire v984f66;
  wire v984f67;
  wire v984f70;
  wire v984f71;
  wire v984f72;
  wire v984f73;
  wire v984f74;
  wire v984f75;
  wire v984f76;
  wire v984f77;
  wire v984f78;
  wire v984f7a;
  wire v984f7b;
  wire v984f7c;
  wire v984f7d;
  wire v984f7e;
  wire v984f7f;
  wire v984f80;
  wire v984f81;
  wire v984f82;
  wire v984f84;
  wire v984f85;
  wire v984f86;
  wire v984f87;
  wire v984f88;
  wire v984f89;
  wire v984f8a;
  wire v984f8b;
  wire v984f8c;
  wire v984f8d;
  wire v984f8f;
  wire v984f90;
  wire v984f91;
  wire v984f92;
  wire v984f94;
  wire v984f95;
  wire v984f96;
  wire v9933b7;
  wire v9933b8;
  wire v9933b9;
  wire v9933ba;
  wire v9933bb;
  wire v9933bc;
  wire v9933bd;
  wire v9933be;
  wire v9933bf;
  wire v9933c0;
  wire v9933c1;
  wire v9933c2;
  wire v9933c3;
  wire v9933c4;
  wire v9933c5;
  wire v9933c6;
  wire v9933c7;
  wire v9933c8;
  wire v9933c9;
  wire v9933ca;
  wire v9933cb;
  wire v9933cc;
  wire v9933cd;
  wire v9933ce;
  wire v9933cf;
  wire v9933d0;
  wire v9933d1;
  wire v9933d2;
  wire v9933d3;
  wire v9933d4;
  wire v9933d5;
  wire v9933d6;
  wire v9933d7;
  wire v9933d8;
  wire v9933d9;
  wire v9933da;
  wire v9933db;
  wire v9933dc;
  reg hready_p;
  input hready;
  reg hbusreq0_p;
  input hbusreq0;
  reg hlock0_p;
  input hlock0;
  reg hbusreq1_p;
  input hbusreq1;
  reg hlock1_p;
  input hlock1;
  reg hbusreq2_p;
  input hbusreq2;
  reg hlock2_p;
  input hlock2;
  reg hburst0_p;
  input hburst0;
  reg hburst1_p;
  input hburst1;
  reg hmaster0_p;
  output hmaster0;
  reg hmaster1_p;
  output hmaster1;
  reg hmastlock_p;
  output hmastlock;
  reg start_p;
  output start;
  reg decide_p;
  output decide;
  reg locked_p;
  output locked;
  reg hgrant0_p;
  output hgrant0;
  reg hgrant1_p;
  output hgrant1;
  reg hgrant2_p;
  output hgrant2;
  reg busreq_p;
  output busreq;
  reg stateA1_p;
  output stateA1;
  reg stateG2_p;
  output stateG2;
  reg stateG3_0_p;
  output stateG3_0;
  reg stateG3_1_p;
  output stateG3_1;
  reg stateG3_2_p;
  output stateG3_2;
  reg stateG10_1_p;
  output stateG10_1;
  reg stateG10_2_p;
  output stateG10_2;
  reg jx0_p;
  output jx0;
  reg jx1_p;
  output jx1;
  reg jx2_p;
  output jx2;

assign v9adce4 = hgrant0_p & v9adcda | !hgrant0_p & v9adce3;
assign v8ea86c = hmaster1_p & v8ea863 | !hmaster1_p & v8ea834;
assign v97389e = hbusreq1_p & v973893 | !hbusreq1_p & v97388d;
assign v99658c = hgrant0_p & v996581 | !hgrant0_p & v99658b;
assign v9999ac = hbusreq0_p & v9999a0 | !hbusreq0_p & a14d40;
assign v9998e7 = hlock0_p & v9998e5 | !hlock0_p & v9998e6;
assign v9d26f0 = hbusreq0_p & v9d26ef | !hbusreq0_p & v9d267e;
assign v8ea92e = hgrant0_p & v8ea881 | !hgrant0_p & v8ea92d;
assign v9adc1e = hbusreq0_p & v9adc1d | !hbusreq0_p & v9adc1c;
assign a15487 = hbusreq0_p & a15415 | !hbusreq0_p & a15444;
assign v9d26e1 = hmaster1_p & v9d26e0 | !hmaster1_p & !v9d2671;
assign v9baef8 = decide_p & v9baef7 | !decide_p & !v84563c;
assign v9baf8d = hbusreq1_p & v9baf8c | !hbusreq1_p & a15507;
assign v9bae99 = decide_p & v9bae98 | !decide_p & !v84563c;
assign v9ed48b = hbusreq0_p & v9ed484 | !hbusreq0_p & v9ed48a;
assign v9d2709 = hgrant0_p & v84563c | !hgrant0_p & !v845647;
assign v9ed4dc = hmaster1_p & v9ed4db | !hmaster1_p & v9ed472;
assign v9739a6 = hbusreq0_p & v97399a | !hbusreq0_p & v9739a5;
assign v9738bc = hready_p & v9738a3 | !hready_p & !v9738bb;
assign v9933d5 = hmaster0_p & v9933d4 | !hmaster0_p & v84563c;
assign v9ed457 = stateG2_p & v84563c | !stateG2_p & !v9ed456;
assign v8ea849 = hmaster1_p & v8ea847 | !hmaster1_p & v8ea7f4;
assign v9d278d = hbusreq0 & v9d26e1 | !hbusreq0 & v9d278c;
assign v973990 = hlock0_p & v97398e | !hlock0_p & v97398f;
assign decide = !v984f96;
assign v9adcd9 = hmaster1_p & v9adc75 | !hmaster1_p & !v9adca2;
assign v9739cd = hbusreq0_p & v9738f7 | !hbusreq0_p & v97397f;
assign v984f53 = hbusreq0 & v984f4f | !hbusreq0 & v984f52;
assign v9ed48a = hmaster1_p & v9ed46f | !hmaster1_p & v9ed489;
assign v9baf13 = hmaster0_p & v9baf10 | !hmaster0_p & !v9ed476;
assign v973933 = hgrant0_p & v97392e | !hgrant0_p & v973932;
assign v9d26ce = decide_p & v9d26cd | !decide_p & v9d2681;
assign v9933ce = hgrant0_p & v9933bd | !hgrant0_p & v9933cd;
assign v8ea869 = hmaster1_p & v8ea867 | !hmaster1_p & v8ea82d;
assign v8ea818 = locked_p & v8ea7e9 | !locked_p & !v8ea7ea;
assign v9855a6 = hbusreq0 & v98559d | !hbusreq0 & v9855a5;
assign v9ed416 = locked_p & v9ed415 | !locked_p & v973889;
assign v973924 = hbusreq0_p & v973914 | !hbusreq0_p & v973923;
assign v9baef7 = hlock2_p & v9baef6 | !hlock2_p & v84563c;
assign v98564e = hready & v98564d | !hready & !v84563c;
assign v9d2771 = hbusreq0_p & v9d26e5 | !hbusreq0_p & v9d2770;
assign v9ed43c = hbusreq1_p & v9ed43b | !hbusreq1_p & v84563c;
assign v8ea7e6 = locked_p & v8ea7e5 | !locked_p & v84563c;
assign v99999b = hready_p & v99998e | !hready_p & v99999a;
assign v8ea80b = hmaster0_p & v8ea80a | !hmaster0_p & v84563c;
assign a154f0 = hlock0_p & v84563c | !hlock0_p & !a154ef;
assign v8ea806 = hmaster0_p & v8ea805 | !hmaster0_p & v84563c;
assign v9a6ada = hbusreq1_p & v9a6ab9 | !hbusreq1_p & v84563c;
assign v985562 = stateA1_p & v985561 | !stateA1_p & v9854bf;
assign v9adc7a = hmaster0_p & v9adc79 | !hmaster0_p & v84563c;
assign v9739b9 = hmaster1_p & v9739b8 | !hmaster1_p & v973964;
assign v98558f = stateG2_p & v84563c | !stateG2_p & v98558e;
assign v9855ec = hbusreq0_p & v9855eb | !hbusreq0_p & v9855e8;
assign v9d2786 = hbusreq0 & v9d2784 | !hbusreq0 & !v9d2785;
assign v973946 = hmaster0_p & v973945 | !hmaster0_p & v9738a4;
assign v84563c = 1;
assign v8ea805 = hbusreq1_p & v8ea802 | !hbusreq1_p & v8ea804;
assign v98560a = hmaster1_p & v985609 | !hmaster1_p & v84563c;
assign v984e69 = hmaster0_p & v984e66 | !hmaster0_p & v984e68;
assign v9adcc1 = hmaster0_p & v9adc95 | !hmaster0_p & !v9adc77;
assign v9ed4b3 = hlock1_p & v8c20d7 | !hlock1_p & !v84563c;
assign v9738b5 = hbusreq0_p & v9738b3 | !hbusreq0_p & v9738b4;
assign hmastlock = v8c20e1;
assign v9d273c = hgrant0_p & v84563c | !hgrant0_p & !v9d273b;
assign v9ed467 = hmastlock_p & v9ed466 | !hmastlock_p & v84563c;
assign v8ea913 = hmaster1_p & v8ea880 | !hmaster1_p & v8ea912;
assign v985627 = hbusreq1_p & v985626 | !hbusreq1_p & v845641;
assign v9adcb5 = hbusreq1_p & v9adca5 | !hbusreq1_p & !v9adcb4;
assign v97390a = hlock0_p & v973908 | !hlock0_p & v973909;
assign v9adc35 = hbusreq1_p & v9adc20 | !hbusreq1_p & !v9adc34;
assign v8c116b = hmaster1_p & v8c116a | !hmaster1_p & !v84563c;
assign v9ecda7 = jx2_p & v9ecda6 | !jx2_p & v9ed533;
assign v999984 = hready_p & v999976 | !hready_p & !v999983;
assign v9855f4 = hbusreq0 & v9855ea | !hbusreq0 & v9855f3;
assign v973954 = hmaster1_p & v9738b7 | !hmaster1_p & !v973940;
assign v9d2737 = hmaster0_p & v9d2736 | !hmaster0_p & v845647;
assign v9d26ad = hbusreq1 & v9d26ac | !hbusreq1 & !v84563c;
assign v99989e = hbusreq0_p & v99989d | !hbusreq0_p & v84563c;
assign v9d2798 = hgrant0_p & v84563c | !hgrant0_p & v9d2797;
assign v8ea935 = hgrant0_p & v8ea8b5 | !hgrant0_p & v8ea934;
assign v8ea829 = hmaster1_p & v8ea823 | !hmaster1_p & v8ea828;
assign v97398e = hmaster1_p & v97398d | !hmaster1_p & v973946;
assign v8ea82d = hmaster0_p & v8ea827 | !hmaster0_p & v8ea82c;
assign v9adbf5 = hmaster0_p & v9adbf2 | !hmaster0_p & v9adbee;
assign v99659d = hmaster0_p & v99659c | !hmaster0_p & v8ea822;
assign v8c20b8 = hlock2_p & v84565c | !hlock2_p & !v8c20b7;
assign v97395c = hbusreq1_p & v9738ea | !hbusreq1_p & v97388d;
assign v9d26e0 = hmaster0_p & v9d26df | !hmaster0_p & !v84563c;
assign v985586 = hgrant0_p & v98556e | !hgrant0_p & v985585;
assign v9d2672 = hmaster1_p & v9d2670 | !hmaster1_p & !v9d2671;
assign v87bd68 = stateA1_p & v84563c | !stateA1_p & v883467;
assign v985501 = hmaster0_p & v9854fb | !hmaster0_p & v985500;
assign v9baf0a = hburst1 & v84563c | !hburst1 & !v87f892;
assign a153e9 = hlock0_p & a153d6 | !hlock0_p & a153e8;
assign v99655a = hmaster0_p & v996559 | !hmaster0_p & v9adbee;
assign v8c20c3 = hbusreq1_p & v8c20c2 | !hbusreq1_p & !v8c20c1;
assign v97388a = locked_p & v973888 | !locked_p & v973889;
assign v8c20c5 = hmaster1_p & v8c20c3 | !hmaster1_p & v8c20c4;
assign v985621 = stateG2_p & v84563c | !stateG2_p & v985620;
assign v9738e2 = stateG10_1_p & v973889 | !stateG10_1_p & !v9738cb;
assign v973992 = hmaster1_p & v973991 | !hmaster1_p & v97394b;
assign v984e71 = stateG10_1_p & v84563c | !stateG10_1_p & v984e70;
assign v99656c = hmaster1_p & v9adc09 | !hmaster1_p & v996564;
assign v9adbeb = hmastlock_p & v9adbea | !hmastlock_p & !v84563c;
assign v973906 = decide_p & v973901 | !decide_p & !v973905;
assign v8ea925 = decide_p & v8ea7ee | !decide_p & v8ea8e3;
assign v9965c4 = hbusreq0_p & v9965c2 | !hbusreq0_p & v9965c3;
assign v84566c = stateG3_1_p & v84563c | !stateG3_1_p & !v84563c;
assign v9b40cd = hgrant2_p & v9b40c0 | !hgrant2_p & !v9b40cc;
assign v9adcea = decide_p & v9adce4 | !decide_p & v9adce9;
assign v8ea89f = decide_p & v8ea7ee | !decide_p & v8ea89e;
assign v9933d8 = hgrant0_p & v9933bf | !hgrant0_p & v9933d7;
assign v9adc63 = stateG10_1_p & v9adc61 | !stateG10_1_p & !v9adc62;
assign v9933b7 = locked_p & v845656 | !locked_p & !v84563c;
assign v9738d7 = hbusreq1_p & v9738d6 | !hbusreq1_p & v97388d;
assign v9d44c5 = jx1_p & v9d44bf | !jx1_p & v9d44c4;
assign v9855e7 = hmaster1_p & v9855e6 | !hmaster1_p & v985589;
assign v8c115f = hmaster1_p & v8c115e | !hmaster1_p & v8c1153;
assign v98562c = hlock1_p & v98562a | !hlock1_p & !v84563c;
assign v9854ab = hready & v985497 | !hready & v9854aa;
assign v9d276d = hgrant2_p & v9d2756 | !hgrant2_p & v9d276c;
assign a154f5 = hready_p & a154bc | !hready_p & a154f3;
assign v9ed532 = hready_p & v9ed530 | !hready_p & v9ed531;
assign v9739e9 = hmaster1_p & v97388b | !hmaster1_p & v9739e8;
assign a14daf = decide_p & a14dae | !decide_p & v84565c;
assign v8ea7f2 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea7ef;
assign v9965cb = hmaster1_p & v9965c9 | !hmaster1_p & v99659f;
assign v985633 = hmaster1_p & v985632 | !hmaster1_p & v985628;
assign v9adc6a = hmaster1_p & v9adc69 | !hmaster1_p & v9adc3b;
assign v9baf63 = hbusreq1_p & v9baf5e | !hbusreq1_p & v9baf62;
assign v9d26b6 = hmaster0_p & v9d26af | !hmaster0_p & v84563c;
assign v8ea8b2 = decide_p & v8ea7ee | !decide_p & v8ea8b1;
assign v9a6aba = hmaster0_p & v9a6ab9 | !hmaster0_p & v84563c;
assign v9adc8c = hlock0_p & v9adc89 | !hlock0_p & v9adc8b;
assign v9baf6b = hmaster1_p & v9baf56 | !hmaster1_p & v9baf6a;
assign v97391f = hmaster0_p & v97391e | !hmaster0_p & v9738d7;
assign v9738dc = locked_p & v973893 | !locked_p & v97388d;
assign v98551d = hbusreq0 & v985517 | !hbusreq0 & v98551c;
assign v9999d9 = hmaster1_p & v84565c | !hmaster1_p & a154a2;
assign v8e79a2 = hbusreq0_p & v8e79a1 | !hbusreq0_p & v8e79a0;
assign v9baf08 = hburst0 & v87f892 | !hburst0 & v9baf07;
assign v9739c3 = decide_p & v97393e | !decide_p & v97393a;
assign v9adbee = hmastlock_p & a2bb5d | !hmastlock_p & !v84563c;
assign v9ed49d = hlock1_p & v9ed49c | !hlock1_p & v84563c;
assign v9b40c0 = hready_p & v84563c | !hready_p & v845654;
assign a1540a = hbusreq0_p & a15409 | !hbusreq0_p & a15408;
assign v9adc71 = hgrant2_p & v9adc59 | !hgrant2_p & v9adc70;
assign v8ea83e = hlock0 & v8ea83d | !hlock0 & v8ea837;
assign v973966 = hbusreq1_p & v9738ea | !hbusreq1_p & v9738eb;
assign v8ea831 = hlock1 & v8ea7e9 | !hlock1 & v8ea818;
assign v9ed45c = hburst0 & v9ed45a | !hburst0 & v9ed45b;
assign v9baf7a = hmaster1_p & v84563c | !hmaster1_p & v9baf79;
assign v9ed436 = hbusreq1_p & v9ed435 | !hbusreq1_p & v84563c;
assign v9739b7 = hbusreq0_p & v9739b4 | !hbusreq0_p & v9739b6;
assign v9855d6 = hbusreq0_p & v985541 | !hbusreq0_p & v9855d5;
assign v9baf1e = stateG10_1_p & v9baf1a | !stateG10_1_p & v9baf1d;
assign v9adc14 = hmaster1_p & v9adc13 | !hmaster1_p & v8ea7ef;
assign v9ed45a = busreq_p & v9ed457 | !busreq_p & v9ed459;
assign v8e79a3 = hmaster0_p & v8e799a | !hmaster0_p & v84563c;
assign v9ed4bd = locked_p & v9ed486 | !locked_p & v84563c;
assign v9738a0 = hmaster1_p & v97389a | !hmaster1_p & v97389f;
assign v9baf7c = hmaster0_p & v84563c | !hmaster0_p & v9ed4bd;
assign v8c20dd = hgrant0_p & v8c20c0 | !hgrant0_p & v8c20dc;
assign v9ed521 = hready_p & v9ed50b | !hready_p & v9ed520;
assign v9739f7 = hmaster1_p & v9738b0 | !hmaster1_p & v9739f4;
assign v9999a9 = hready_p & v9999a7 | !hready_p & !v9999a8;
assign v9baf43 = hbusreq1_p & v9ed419 | !hbusreq1_p & v9ed41d;
assign v9d2700 = hbusreq1_p & v9d26d0 | !hbusreq1_p & !v9d26d1;
assign v9d26b9 = hmaster1_p & v9d26b6 | !hmaster1_p & !v9d2673;
assign v8c1142 = locked_p & v8c1120 | !locked_p & !v84563c;
assign v9998fe = hbusreq0 & v9998fd | !hbusreq0 & !v84563c;
assign v996590 = hmaster0_p & v99658f | !hmaster0_p & !v9adc37;
assign v9d26d1 = stateG10_1_p & v84563c | !stateG10_1_p & !v9d26d0;
assign v9854c5 = hbusreq1_p & v9854c4 | !hbusreq1_p & v84563c;
assign v973895 = hbusreq1_p & v973894 | !hbusreq1_p & v97388e;
assign v9bae81 = hmastlock_p & v8e7990 | !hmastlock_p & !v84563c;
assign v97392a = decide_p & v973922 | !decide_p & v973929;
assign stateG3_0 = !v9a6ae3;
assign v985536 = stateG2_p & v84563c | !stateG2_p & !v985535;
assign v9adbfc = hlock2_p & v9adbf7 | !hlock2_p & v9adbfb;
assign v8ea923 = hready_p & v8ea80d | !hready_p & v8ea922;
assign v9baf8f = hmaster0_p & v9baf8d | !hmaster0_p & v9baf8e;
assign v9adc17 = hmaster0_p & v9adbec | !hmaster0_p & v9adbf1;
assign v984eb0 = hgrant0_p & v984ea4 | !hgrant0_p & v984eaf;
assign v984e5e = hmaster0_p & v984e5d | !hmaster0_p & v84563c;
assign v9a6aa5 = hmaster0_p & v9a6aa4 | !hmaster0_p & v9a6aa2;
assign v9ed488 = hbusreq1_p & v9ed487 | !hbusreq1_p & !v84563c;
assign v984f75 = hbusreq0_p & v984f72 | !hbusreq0_p & v984f74;
assign v9adc4d = hmaster0_p & v9adc4c | !hmaster0_p & !v8ea822;
assign a14dba = hready_p & a14daf | !hready_p & a14da2;
assign v8ea8ed = hmaster1_p & v8ea867 | !hmaster1_p & v8ea8d2;
assign v9d2662 = stateG2_p & v84563c | !stateG2_p & v845666;
assign v8c20d8 = stateG10_1_p & v84563c | !stateG10_1_p & !v8c20d7;
assign v9adc98 = hmaster0_p & v9adc95 | !hmaster0_p & v9adc94;
assign v984f2f = hbusreq0 & v984f29 | !hbusreq0 & v984f2e;
assign v9999b8 = hlock0_p & v9999b7 | !hlock0_p & v84563c;
assign v9baf4b = stateG2_p & v866c94 | !stateG2_p & !v9ed411;
assign v98563d = hlock0_p & v98563b | !hlock0_p & !v98563c;
assign v98553b = hlock1_p & v98553a | !hlock1_p & !v84563c;
assign v9adc25 = hgrant1_p & v9adbf1 | !hgrant1_p & v9adbee;
assign v9739c1 = hbusreq2_p & v973984 | !hbusreq2_p & !v9739c0;
assign v9854fa = hlock1_p & v9854f1 | !hlock1_p & v9854f9;
assign a15414 = hmaster1_p & a153ba | !hmaster1_p & a1540e;
assign stateG10_2 = !a4ce72;
assign v8ea7ec = hbusreq1_p & v8ea7e9 | !hbusreq1_p & !v8ea7eb;
assign v8c20e0 = hgrant2_p & v8c20d4 | !hgrant2_p & !v8c20df;
assign v9d2682 = decide_p & v9d267a | !decide_p & v9d2681;
assign v8c1174 = busreq_p & v8c1172 | !busreq_p & !v8c1173;
assign v9adc8a = hmaster0_p & v9adc87 | !hmaster0_p & !v84563c;
assign v9d2720 = hmaster1_p & v9d271f | !hmaster1_p & !v9d2671;
assign v999971 = hmaster1_p & v9baf7c | !hmaster1_p & v84563c;
assign v9738aa = hmaster0_p & v9738a7 | !hmaster0_p & v973889;
assign v985526 = hready & v985525 | !hready & v84563c;
assign v985519 = hmaster1_p & v985518 | !hmaster1_p & v985502;
assign v9998fc = hmaster1_p & v9baf79 | !hmaster1_p & v84563c;
assign v8c1175 = locked_p & v8c1174 | !locked_p & !v84563c;
assign v99992d = hbusreq0_p & v99992c | !hbusreq0_p & !v84563c;
assign v9854bb = hlock2_p & v9854b2 | !hlock2_p & v9854ba;
assign v9baf55 = hbusreq1_p & v9baf51 | !hbusreq1_p & !v9baf54;
assign v8ea8cc = hbusreq0_p & v8ea881 | !hbusreq0_p & v8ea8cb;
assign v9999b5 = hgrant2_p & v9999af | !hgrant2_p & !v9999b4;
assign v9d267a = hbusreq2 & v9d2675 | !hbusreq2 & v9d2679;
assign v9d2783 = hbusreq0_p & v9d2757 | !hbusreq0_p & v9d2782;
assign v8ea884 = hbusreq0_p & v8ea881 | !hbusreq0_p & v8ea883;
assign v97394a = hlock0_p & v973947 | !hlock0_p & v973949;
assign v8ea880 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea7ef;
assign v9965af = hmaster0_p & v9adc54 | !hmaster0_p & v8ea7e9;
assign v98548f = hready & v84563c | !hready & v84565c;
assign v9bae94 = hbusreq1_p & v9bae93 | !hbusreq1_p & v84563c;
assign v8e79d6 = hgrant0_p & v8e79b0 | !hgrant0_p & v8e79d5;
assign v9ed4f7 = hmaster1_p & v84563c | !hmaster1_p & !v9ed4f6;
assign v8c1163 = hgrant2_p & v8c113e | !hgrant2_p & v8c1162;
assign v9854d2 = hmaster0_p & v9854cf | !hmaster0_p & v9854d1;
assign stateG2 = !v8c1180;
assign v8c1129 = hbusreq0_p & v8c1128 | !hbusreq0_p & v8c1127;
assign v984f5c = hgrant1_p & v9854c4 | !hgrant1_p & !v84563c;
assign v9854e5 = hmaster1_p & v9854e4 | !hmaster1_p & v9854d3;
assign v9999b1 = hbusreq0 & v9999b0 | !hbusreq0 & v99998c;
assign v9baf25 = hbusreq0 & v9baf15 | !hbusreq0 & v9baf24;
assign v9d275d = hbusreq1_p & v9d275b | !hbusreq1_p & !v9d275c;
assign v98559b = hmaster0_p & v84563c | !hmaster0_p & v985599;
assign v9ed411 = stateA1_p & v84563c | !stateA1_p & !a1541d;
assign v8ea88b = hlock1 & v8ea819 | !hlock1 & v8ea818;
assign v99992a = hmaster0_p & v999909 | !hmaster0_p & v999929;
assign v8ea85d = hbusreq1_p & v8ea800 | !hbusreq1_p & v8ea85c;
assign v9adcdb = hmaster0_p & v9adca7 | !hmaster0_p & !v9adc75;
assign v9d26c1 = hmaster0_p & v9d26c0 | !hmaster0_p & !v84563c;
assign v9854b3 = hlock1_p & v845641 | !hlock1_p & !v84563c;
assign v973911 = decide_p & v97390c | !decide_p & v973910;
assign v9ed4d6 = hbusreq0_p & v9ed4d4 | !hbusreq0_p & v9ed4d5;
assign v9ed44d = hlock1_p & v9ed44c | !hlock1_p & v84563c;
assign v8c1120 = hmastlock_p & v8c111f | !hmastlock_p & !v84563c;
assign v9d2698 = hmaster0_p & v845647 | !hmaster0_p & v9d2696;
assign v9854c0 = stateA1_p & v84563c | !stateA1_p & !v9854bf;
assign v9a6ad5 = hmaster0_p & v9a6ad4 | !hmaster0_p & v84563c;
assign v9d27b5 = hbusreq0_p & v9d26e8 | !hbusreq0_p & !v9d267c;
assign v9d26ae = hgrant1_p & v9d26a4 | !hgrant1_p & !v9d26ad;
assign v9d266b = stateA1_p & v84563c | !stateA1_p & !v85a40d;
assign v996574 = hmaster1_p & v996573 | !hmaster1_p & v8ea7f2;
assign a153e8 = hmaster1_p & a153d4 | !hmaster1_p & a153e7;
assign v8ea931 = hgrant2_p & v8ea7f8 | !hgrant2_p & v8ea930;
assign v8ea8bf = hlock0 & v8ea8be | !hlock0 & v8ea8bb;
assign v9d26da = decide_p & v9d26cd | !decide_p & v9d26bc;
assign a14d40 = hmaster0_p & v845646 | !hmaster0_p & !v84563c;
assign v9ed447 = hmaster0_p & v84563c | !hmaster0_p & !v9ed446;
assign v8c1162 = hready_p & v8c1156 | !hready_p & !v8c1161;
assign v996588 = hmaster1_p & v9adc28 | !hmaster1_p & !v996587;
assign v9adc80 = hmaster1_p & v9adc7f | !hmaster1_p & !v9adc7a;
assign v973936 = hgrant2_p & v973912 | !hgrant2_p & !v973935;
assign v996576 = hbusreq0_p & v996574 | !hbusreq0_p & v996575;
assign v9a6ac3 = hmaster0_p & v9a6ac2 | !hmaster0_p & v84563c;
assign v9adc76 = locked_p & v9adc74 | !locked_p & !v9adc75;
assign v97393f = hbusreq1_p & v97388c | !hbusreq1_p & v973894;
assign v9adcb4 = stateG10_1_p & v9adc75 | !stateG10_1_p & !v9adca5;
assign v9854f1 = hready & v9854f0 | !hready & !v9ed45a;
assign v984e5c = hmaster1_p & v984e57 | !hmaster1_p & v984e5b;
assign v9d2751 = hbusreq0 & v9d271b | !hbusreq0 & v9d2750;
assign v999914 = stateA1_p & a153cb | !stateA1_p & !a2fb4c;
assign v9a6a95 = stateG3_2_p & v84563c | !stateG3_2_p & v9a6a94;
assign v845654 = hmaster1_p & v84563c | !hmaster1_p & !v84563c;
assign v9baf79 = hmaster0_p & v84563c | !hmaster0_p & v9ed44c;
assign v8ea838 = hlock0 & v8ea830 | !hlock0 & v8ea837;
assign v973909 = hmaster1_p & v973907 | !hmaster1_p & v9738aa;
assign v985645 = hmaster1_p & v9d2724 | !hmaster1_p & v84563c;
assign v973a3b = hmaster1_p & v973a2f | !hmaster1_p & v973a10;
assign v8ea850 = hbusreq0 & v8ea84a | !hbusreq0 & v8ea84f;
assign v863b4b = stateG3_2_p & v84563c | !stateG3_2_p & !v85a40d;
assign v8c20d1 = hready_p & v8c20c7 | !hready_p & v8c20d0;
assign a14da2 = decide_p & a14da1 | !decide_p & v84565c;
assign v9d2702 = hmaster1_p & v9d2701 | !hmaster1_p & v845647;
assign v8c1154 = hmaster1_p & v8c1144 | !hmaster1_p & !v8c1153;
assign a154a1 = hbusreq2_p & a15432 | !hbusreq2_p & a15496;
assign v9adc2d = hbusreq1_p & v9adc2b | !hbusreq1_p & v9adc2c;
assign v8c112a = hmaster0_p & v8c1120 | !hmaster0_p & !v84563c;
assign v985565 = locked_p & v985564 | !locked_p & v84563c;
assign v9998ed = hburst0 & v8e7991 | !hburst0 & v9998ec;
assign v854662 = hbusreq0_p & v898b4e | !hbusreq0_p & !v84563c;
assign v9ed470 = hlock1_p & v845656 | !hlock1_p & !v84563c;
assign v8ea859 = hbusreq2 & v8ea857 | !hbusreq2 & v8ea858;
assign v973918 = hbusreq0_p & v973916 | !hbusreq0_p & !v973917;
assign a14d6e = hbusreq0_p & v84563c | !hbusreq0_p & v845646;
assign v8ea919 = hmaster1_p & v8ea909 | !hmaster1_p & v8ea918;
assign v984ee6 = hmaster1_p & v984ee3 | !hmaster1_p & v984ee5;
assign v9baf65 = hgrant1_p & v9baf64 | !hgrant1_p & v9ed419;
assign v9bae7b = stateA1_p & v84563c | !stateA1_p & !v8e7990;
assign v9f3577 = decide_p & v9f356c | !decide_p & v9f3576;
assign v9d279d = hbusreq2 & v9d279a | !hbusreq2 & v9d279c;
assign v8c113d = decide_p & v8c112f | !decide_p & v8c113c;
assign v9854e1 = hlock0_p & v9854de | !hlock0_p & v9854e0;
assign v984ea6 = stateG10_1_p & v84563c | !stateG10_1_p & !v984ea5;
assign v99998c = hgrant0_p & v99998b | !hgrant0_p & !a14d6e;
assign v8e79b6 = hmaster0_p & v8e79b5 | !hmaster0_p & v84563c;
assign v984f89 = decide_p & v984f38 | !decide_p & v984f88;
assign v985610 = hbusreq2 & v845641 | !hbusreq2 & v98560f;
assign v8c117d = decide_p & v8c1169 | !decide_p & v8c1160;
assign busreq = v9d27c7;
assign v9738f0 = hgrant0_p & v9738df | !hgrant0_p & v9738ef;
assign v9738c1 = hmaster1_p & v9738b0 | !hmaster1_p & v9738c0;
assign v8ea87c = hmaster1_p & v8ea87b | !hmaster1_p & v8ea7f2;
assign v8c1145 = hgrant1_p & v8c111a | !hgrant1_p & !v84563c;
assign v8e79d8 = decide_p & v8e79cf | !decide_p & v8e79c7;
assign v8c1119 = hmastlock_p & v8c1118 | !hmastlock_p & !v84563c;
assign v9965b2 = decide_p & v9965b1 | !decide_p & v996576;
assign v9adcae = hmaster0_p & v9adcad | !hmaster0_p & !v84563c;
assign v9adc45 = locked_p & v9adbfe | !locked_p & v8ea7e9;
assign v8c20be = hmaster1_p & v84563c | !hmaster1_p & v8c20b6;
assign v973a21 = hbusreq2_p & v973a20 | !hbusreq2_p & !v9739e6;
assign v9739ee = hmaster0_p & v9739eb | !hmaster0_p & !v973893;
assign v98563b = hmaster1_p & v98563a | !hmaster1_p & v985628;
assign v9baea7 = hbusreq0_p & v9baea6 | !hbusreq0_p & v84563c;
assign v9ed4d1 = hbusreq2 & v9ed4ce | !hbusreq2 & !v9ed4d0;
assign v9999e9 = hlock2_p & v9999e3 | !hlock2_p & v9999e8;
assign v9baf70 = hgrant1_p & v9baf6f | !hgrant1_p & !v9ed41d;
assign v9adc05 = hmaster0_p & v9adc02 | !hmaster0_p & v8ea7ea;
assign v973959 = hmaster0_p & v97389b | !hmaster0_p & !v9738c4;
assign v9d26cc = hbusreq0 & v9d26c9 | !hbusreq0 & v9d26cb;
assign v845660 = hgrant1_p & v84563c | !hgrant1_p & !v84563c;
assign v973a0d = hmaster1_p & v9738cd | !hmaster1_p & !v973a0c;
assign v9ed4eb = hgrant0_p & v9ed4ea | !hgrant0_p & !v9ed4b6;
assign v999902 = hburst1_p & v8763e4 | !hburst1_p & v85a40d;
assign v9d2776 = hmaster1_p & v9d2775 | !hmaster1_p & v9d2671;
assign v9738a1 = hbusreq0_p & v97389d | !hbusreq0_p & v9738a0;
assign v9738b8 = hmaster1_p & v9738b7 | !hmaster1_p & !v973890;
assign v8ea7ff = hbusreq0_p & v8ea7f9 | !hbusreq0_p & v8ea7fe;
assign v9baf5d = hbusreq1 & v9ed416 | !hbusreq1 & v9baf5c;
assign v9d274f = hbusreq2 & v9d274b | !hbusreq2 & v9d274e;
assign v984ee5 = hmaster0_p & v985627 | !hmaster0_p & v9854d0;
assign v985607 = hmastlock_p & v98549b | !hmastlock_p & v84563c;
assign v9738af = hbusreq0_p & v9738ac | !hbusreq0_p & v9738ae;
assign v996561 = hlock1_p & v9adbfe | !hlock1_p & !v8ea7ea;
assign v9998da = hgrant0_p & v9998d9 | !hgrant0_p & !a14d6e;
assign v9998d5 = hbusreq0_p & v9998a0 | !hbusreq0_p & v845646;
assign v9baf5b = hmastlock_p & v9baf5a | !hmastlock_p & v84563c;
assign v9965a5 = hgrant2_p & v996578 | !hgrant2_p & v9965a4;
assign v9855bf = hbusreq0_p & v9855be | !hbusreq0_p & v845641;
assign v984edd = hbusreq2 & v984edb | !hbusreq2 & v984edc;
assign v9855c3 = hmaster1_p & v9855c1 | !hmaster1_p & v9ed438;
assign a14d3e = hbusreq0_p & v845644 | !hbusreq0_p & !v84563c;
assign v9d2766 = hgrant0_p & v9d2725 | !hgrant0_p & v9d2765;
assign v9baeb1 = hbusreq0_p & v9baeae | !hbusreq0_p & v9baeb0;
assign v8ea83f = hbusreq0 & v8ea838 | !hbusreq0 & v8ea83e;
assign v9ed568 = hready_p & v84563c | !hready_p & v9ed567;
assign a1550b = hlock0_p & v84563c | !hlock0_p & a1550a;
assign v8e79ac = decide_p & v8e79a8 | !decide_p & v8e79ab;
assign v985594 = hmaster0_p & v84563c | !hmaster0_p & !v985593;
assign v8ea8f4 = hbusreq2 & v8ea8f2 | !hbusreq2 & v8ea8f3;
assign v984eb9 = hmaster0_p & v984eb8 | !hmaster0_p & v84563c;
assign v9854a0 = hready & v98549d | !hready & v98549f;
assign v8ea872 = hgrant0_p & v8ea871 | !hgrant0_p & v8ea86a;
assign a14dab = hmaster1_p & a14da9 | !hmaster1_p & a14daa;
assign v8ecba9 = stateG2_p & v84563c | !stateG2_p & !v84566e;
assign v9d2791 = hbusreq2 & v9d2790 | !hbusreq2 & v9d2680;
assign v8c20bc = decide_p & v845656 | !decide_p & v8c20bb;
assign v9adcc0 = decide_p & v9adcb3 | !decide_p & v9adcbf;
assign v9d2675 = hbusreq0 & v9d2672 | !hbusreq0 & v9d2674;
assign v8c115a = hbusreq0_p & v8c1158 | !hbusreq0_p & v8c1159;
assign v9baeb4 = hlock0_p & v9baeb3 | !hlock0_p & v9baeae;
assign v9adcba = hmaster0_p & v9adcb9 | !hmaster0_p & !v84563c;
assign v9baf17 = stateA1_p & v972fac | !stateA1_p & !a2fb4c;
assign v973a31 = hmaster1_p & v97398d | !hmaster1_p & v9739ff;
assign v985499 = hburst1_p & v9a6a94 | !hburst1_p & v84563c;
assign v996557 = hmaster1_p & v996550 | !hmaster1_p & v996556;
assign v8c20ca = hmaster1_p & v8c20c8 | !hmaster1_p & !v8c20c9;
assign v984f24 = hmaster0_p & v98562c | !hmaster0_p & v98562a;
assign v9baf97 = hbusreq0 & v9baf92 | !hbusreq0 & v9baf96;
assign v8ea91d = hgrant0_p & v8ea881 | !hgrant0_p & v8ea91c;
assign v8e79c5 = hmaster0_p & v8e79c4 | !hmaster0_p & v84563c;
assign v9855b8 = hgrant0_p & v9855a4 | !hgrant0_p & v9855b7;
assign v8ea855 = hlock0 & v8ea84e | !hlock0 & v8ea854;
assign v8ea8e3 = hbusreq0_p & v8ea8e2 | !hbusreq0_p & v8ea8a5;
assign v9baf9e = hbusreq2_p & v9baf9d | !hbusreq2_p & !v9baea0;
assign v9baea0 = hgrant2_p & v84565a | !hgrant2_p & v84563c;
assign v8ea876 = hbusreq2 & v8ea874 | !hbusreq2 & v8ea875;
assign v8ea88e = stateG10_1_p & v84563c | !stateG10_1_p & v8ea88d;
assign v984ebb = hgrant0_p & v985645 | !hgrant0_p & v984eba;
assign v8e799c = hbusreq1_p & v8e799b | !hbusreq1_p & v84563c;
assign v9ed493 = hbusreq0_p & v9ed491 | !hbusreq0_p & v9ed492;
assign v8e79cb = decide_p & v84563c | !decide_p & v8e7995;
assign v999919 = hmaster0_p & v999909 | !hmaster0_p & v999918;
assign v8ea8c1 = hlock2 & v8ea8be | !hlock2 & v8ea8c0;
assign v984f46 = hmaster0_p & v84563c | !hmaster0_p & v984f45;
assign v9999cb = hbusreq0 & v9999b9 | !hbusreq0 & v9999ca;
assign v99997c = hbusreq0 & v99997a | !hbusreq0 & !v99997b;
assign v9855f0 = hmaster1_p & v9855ef | !hmaster1_p & v985583;
assign v9999c0 = stateA1_p & v863b4b | !stateA1_p & a153cb;
assign v9738cc = hbusreq1_p & v9738cb | !hbusreq1_p & !v973889;
assign v9adc06 = hmaster1_p & v9adbff | !hmaster1_p & !v9adc05;
assign v9739dd = hgrant0_p & v9739a6 | !hgrant0_p & v9739dc;
assign v9965b8 = hlock0_p & v9965b5 | !hlock0_p & v9965b7;
assign v985571 = stateG2_p & v84563c | !stateG2_p & v985570;
assign v9d26a2 = hbusreq0 & v9d26a0 | !hbusreq0 & !v9d26a1;
assign v9999da = hlock0_p & v9999d9 | !hlock0_p & !v84563c;
assign v985533 = hlock0_p & v985532 | !hlock0_p & v9854b5;
assign a15507 = stateG10_1_p & v84565c | !stateG10_1_p & !v8c20c1;
assign v9d26d6 = hgrant0_p & v84563c | !hgrant0_p & v9d26d5;
assign v9d26dd = hbusreq2_p & v9d26bf | !hbusreq2_p & v9d26dc;
assign v9855fd = hready & v98549d | !hready & v98549e;
assign v9855bb = decide_p & v98551f | !decide_p & v9855ba;
assign v9baf2b = stateG2_p & v84563c | !stateG2_p & !a2fb4d;
assign v9933d2 = decide_p & v8c20b7 | !decide_p & v9933b9;
assign v8ea8ac = hbusreq0_p & v8ea8ab | !hbusreq0_p & v8ea8a5;
assign v97399d = hmaster1_p & v973991 | !hmaster1_p & v973959;
assign v9ed4a3 = hburst1 & v9ed4a2 | !hburst1 & !v84563c;
assign v9ed429 = hburst0 & v9ed424 | !hburst0 & v9ed428;
assign v9adc89 = hmaster1_p & v9adc75 | !hmaster1_p & v9adc88;
assign v9739e4 = decide_p & v9739d7 | !decide_p & v9739e3;
assign v9738d6 = hgrant1_p & v973894 | !hgrant1_p & v973893;
assign v9855cc = hmaster1_p & v9855cb | !hmaster1_p & v9ed438;
assign v999989 = hbusreq0_p & v999988 | !hbusreq0_p & v845646;
assign v8ea7e2 = stateG3_0_p & v84566c | !stateG3_0_p & !v84563c;
assign v9854cd = hmastlock_p & v8ea7fb | !hmastlock_p & v84563c;
assign v9adcd8 = hlock0_p & v9adcd6 | !hlock0_p & !v9adcd7;
assign v8ea862 = decide_p & v8ea861 | !decide_p & v8ea80d;
assign v99997e = hmaster1_p & v99997d | !hmaster1_p & !v99990b;
assign v9d27c7 = jx1_p & v9d274a | !jx1_p & v9d27c6;
assign v8c1131 = hburst1_p & v84563c | !hburst1_p & v8c1130;
assign v985619 = hmaster0_p & v84565c | !hmaster0_p & v985618;
assign v973914 = hmaster1_p & v973913 | !hmaster1_p & v9738be;
assign v973a10 = hmaster0_p & v97393f | !hmaster0_p & v9738dc;
assign v973a1d = hgrant0_p & v973a19 | !hgrant0_p & v973a1c;
assign v8ea928 = hready_p & v8ea862 | !hready_p & v8ea927;
assign v973a0e = hbusreq0_p & v973a09 | !hbusreq0_p & v973a0d;
assign v985575 = stateG2_p & v84563c | !stateG2_p & v985553;
assign v9965d3 = jx1_p & v9d44bf | !jx1_p & !v9965d2;
assign v8ea861 = hgrant0_p & v8ea7ff | !hgrant0_p & v8ea860;
assign v9d27ae = hgrant0_p & v9d267c | !hgrant0_p & v9d27ad;
assign v9d2749 = hbusreq2_p & v9d272f | !hbusreq2_p & v9d2748;
assign v973a11 = hmaster1_p & v9738bd | !hmaster1_p & v973a10;
assign v8c20c8 = hmaster0_p & v845656 | !hmaster0_p & !v8c20ba;
assign v97393c = hmaster1_p & v97389a | !hmaster1_p & v97393b;
assign v9855c8 = hbusreq0_p & v98551b | !hbusreq0_p & v9855c7;
assign v9d2728 = hmaster1_p & v9d2727 | !hmaster1_p & !v9d2671;
assign v9adcb0 = hmaster0_p & v9adcad | !hmaster0_p & v9adc75;
assign v8ea81c = hbusreq1_p & v8ea81b | !hbusreq1_p & v8ea818;
assign v9998a1 = hbusreq0_p & v9998a0 | !hbusreq0_p & v84563c;
assign v9adcb1 = hmaster1_p & v9adca8 | !hmaster1_p & !v9adcb0;
assign v9d2724 = hmaster0_p & v845641 | !hmaster0_p & v84563c;
assign v9ed424 = stateA1_p & v84563c | !stateA1_p & !a153bb;
assign a2f895 = stateA1_p & v863b4b | !stateA1_p & !a2fb4c;
assign v9ed4e8 = hmaster0_p & v9ed43c | !hmaster0_p & !v9ed446;
assign v9855fa = hmaster0_p & v98548f | !hmaster0_p & v985498;
assign v9738f5 = hbusreq0_p & v9738f3 | !hbusreq0_p & v9738f4;
assign v845646 = hbusreq1_p & v84563c | !hbusreq1_p & !v84563c;
assign v9adcc5 = stateG10_1_p & v9adc75 | !stateG10_1_p & !v9adcc4;
assign v9ed434 = locked_p & v9ed433 | !locked_p & !v84563c;
assign v8ea813 = locked_p & v8ea812 | !locked_p & v8ea7e9;
assign v9adccd = hgrant2_p & v9adc9c | !hgrant2_p & v9adccc;
assign v9baef3 = hbusreq2 & v84565c | !hbusreq2 & v84563c;
assign v9baf60 = hbusreq1 & v9ed49c | !hbusreq1 & v9ed4bd;
assign v9738f7 = hmaster1_p & v9738f6 | !hmaster1_p & v9738e8;
assign v999977 = hmaster0_p & v999909 | !hmaster0_p & v9ed476;
assign v9adc11 = locked_p & v9adc10 | !locked_p & v8ea7e9;
assign v973987 = hmaster1_p & v973985 | !hmaster1_p & v97393b;
assign v973a2c = hbusreq0_p & v973994 | !hbusreq0_p & v973a2b;
assign v9adc18 = hmaster0_p & v9adbf2 | !hmaster0_p & v9adbef;
assign v8ea8bb = hgrant0_p & v8ea8b7 | !hgrant0_p & v8ea8ba;
assign v9baf9a = decide_p & v9baf99 | !decide_p & v84563c;
assign a15447 = hbusreq1_p & a153ce | !hbusreq1_p & !v84563c;
assign v9965a8 = hmaster1_p & v9965a6 | !hmaster1_p & v99655c;
assign v9739ed = hmaster1_p & v97389a | !hmaster1_p & v9739ec;
assign v8ea90a = stateG10_1_p & v8ea7ea | !stateG10_1_p & !v8ea88d;
assign v98555b = hgrant0_p & v985542 | !hgrant0_p & v98555a;
assign v9d268e = hgrant1_p & v845647 | !hgrant1_p & !v9d268d;
assign v9b40de = jx1_p & v9b40d0 | !jx1_p & v9b40dd;
assign v9ed4b7 = hgrant0_p & v9ed4a1 | !hgrant0_p & !v9ed4b6;
assign v9965a6 = hmaster0_p & v9adbeb | !hmaster0_p & !v99657e;
assign v8ea845 = hmaster1_p & v8ea7fd | !hmaster1_p & v84563c;
assign v973a04 = hbusreq0_p & v973a01 | !hbusreq0_p & !v973a03;
assign v9ed4ad = hlock1_p & v9ed4a7 | !hlock1_p & v9ed4ac;
assign v9ed4b9 = hmaster1_p & v9ed423 | !hmaster1_p & v9ed4b8;
assign v9999ca = hbusreq0_p & v9999c9 | !hbusreq0_p & v84563c;
assign v9999c1 = stateG2_p & v84563c | !stateG2_p & v9999c0;
assign v9ed46c = hburst0 & v9ed46a | !hburst0 & v9ed46b;
assign v9855c4 = hbusreq0_p & v9855c2 | !hbusreq0_p & v9855c3;
assign v9999af = hready_p & v9999ab | !hready_p & v9999ae;
assign v9adcef = hmaster1_p & v9adced | !hmaster1_p & v9adcc7;
assign v98552c = hmaster1_p & v985528 | !hmaster1_p & v98552b;
assign v9d266f = hlock1_p & v9d2668 | !hlock1_p & v9d266e;
assign v9ed44f = hmaster0_p & v845646 | !hmaster0_p & v9ed44e;
assign v845658 = start_p & v84563c | !start_p & !v84563c;
assign v9d272f = hgrant2_p & v9d26f5 | !hgrant2_p & v9d272e;
assign v999980 = hbusreq0_p & v99997f | !hbusreq0_p & !a14d40;
assign v9d2690 = hbusreq1_p & v9d268f | !hbusreq1_p & v845647;
assign v8c1156 = decide_p & v8c114a | !decide_p & v8c1155;
assign v9d26be = hready_p & v9d26a3 | !hready_p & !v9d26bd;
assign v9933d1 = hgrant2_p & v9933bc | !hgrant2_p & v9933d0;
assign v9855db = hbusreq0 & v9855d4 | !hbusreq0 & v9855da;
assign v973a43 = hmaster1_p & v9739b8 | !hmaster1_p & v973a13;
assign v9999c8 = hmaster1_p & v84563c | !hmaster1_p & v9999c7;
assign v845641 = hready & v84563c | !hready & !v84563c;
assign v984e6d = hmastlock_p & v984e6c | !hmastlock_p & !v84563c;
assign v973989 = hmaster1_p & v973902 | !hmaster1_p & v973940;
assign v99655d = hmaster1_p & v9adbfa | !hmaster1_p & v99655c;
assign v9998fb = hbusreq0 & v9998fa | !hbusreq0 & v84563c;
assign v9b40db = hbusreq2_p & v9b40cd | !hbusreq2_p & v9b40c3;
assign v9738b0 = hmaster0_p & v973885 | !hmaster0_p & v973889;
assign v973a4a = jx2_p & v973a21 | !jx2_p & v973a49;
assign v9855aa = busreq_p & v84563c | !busreq_p & !v9855a9;
assign v9adc5e = hmaster0_p & v9adc24 | !hmaster0_p & v9adbee;
assign v9965c0 = hgrant0_p & v9965ba | !hgrant0_p & v9965bf;
assign v9d2699 = hmaster1_p & v9d2697 | !hmaster1_p & v9d2698;
assign v9739a5 = hmaster1_p & v973999 | !hmaster1_p & v9738dd;
assign v985603 = hmastlock_p & v8e7991 | !hmastlock_p & !v84563c;
assign v9baf38 = hbusreq0_p & v9baf35 | !hbusreq0_p & v9baf37;
assign v9739bd = hgrant0_p & v9739b7 | !hgrant0_p & v9739bc;
assign v9854bc = stateG3_0_p & v84566c | !stateG3_0_p & !v845658;
assign v984ee2 = jx0_p & v9855f9 | !jx0_p & v984ee1;
assign v9d274c = hmaster1_p & v845652 | !hmaster1_p & v9d2671;
assign v8ea909 = hmaster0_p & v8ea908 | !hmaster0_p & v8ea822;
assign v9739d9 = decide_p & v9739d7 | !decide_p & v9739d8;
assign v9adc52 = hgrant2_p & v9adc16 | !hgrant2_p & v9adc51;
assign a154d3 = hlock1_p & a153d1 | !hlock1_p & !v84563c;
assign v9999be = hburst0 & v9999ba | !hburst0 & v9999bd;
assign v9ed46a = stateG2_p & v84563c | !stateG2_p & v9ed456;
assign locked = a14dc2;
assign v97389b = hbusreq1_p & v973889 | !hbusreq1_p & !v97388d;
assign v9baeb5 = hbusreq0_p & v9baeb4 | !hbusreq0_p & v85bb54;
assign v9ed428 = hburst1 & v9ed424 | !hburst1 & v9ed427;
assign v9d26e4 = hlock0_p & v9d26e1 | !hlock0_p & v9d26e3;
assign v8ea906 = hgrant1_p & v8ea813 | !hgrant1_p & v8ea7e9;
assign v973885 = hmastlock_p & v973883 | !hmastlock_p & v973884;
assign v9854a8 = hmaster1_p & v9854a3 | !hmaster1_p & v9854a7;
assign v9d2782 = hmaster1_p & v9d2781 | !hmaster1_p & v845647;
assign v99996c = hmaster0_p & v973885 | !hmaster0_p & !v9ed49c;
assign v9adce0 = hbusreq1_p & v9adca6 | !hbusreq1_p & !v9adcdf;
assign v9adc6e = decide_p & v9adc68 | !decide_p & v9adc6d;
assign v984f3d = hlock0_p & v984f3c | !hlock0_p & v845641;
assign v985631 = hready & v8ea7e5 | !hready & !a153cc;
assign v98562e = hlock0_p & v985629 | !hlock0_p & !v98562d;
assign v9adc68 = hgrant0_p & v9adc5d | !hgrant0_p & v9adc67;
assign v98559e = hmastlock_p & v985522 | !hmastlock_p & !v84563c;
assign v8ea85e = hmaster0_p & v8ea85d | !hmaster0_p & v84563c;
assign v9d27c3 = hready_p & v9d27a0 | !hready_p & !v9d2681;
assign v9ed4e7 = hmaster1_p & v9ed4e6 | !hmaster1_p & v9ed499;
assign v999922 = hmaster0_p & v999909 | !hmaster0_p & !v999921;
assign v9854fb = hbusreq1_p & v9854fa | !hbusreq1_p & v84563c;
assign v999909 = hmastlock_p & v999908 | !hmastlock_p & !v973884;
assign v9bae9f = hgrant2_p & v9bae9a | !hgrant2_p & !v9bae9e;
assign v9854b2 = hbusreq2 & v9854a9 | !hbusreq2 & v9854b1;
assign v9965cf = hready_p & v9965c6 | !hready_p & !v9965ce;
assign v9a6aae = hlock0_p & v9a6aac | !hlock0_p & v9a6aad;
assign v8ea8aa = hmaster0_p & v84563c | !hmaster0_p & v8ea832;
assign v985551 = busreq_p & v98549b | !busreq_p & !v985550;
assign v984f94 = jx2_p & v984f92 | !jx2_p & v984f91;
assign v9d26f8 = hbusreq1_p & v9d26f6 | !hbusreq1_p & !v9d26f7;
assign v99990a = hmaster0_p & v999909 | !hmaster0_p & !v9ed46d;
assign v99993d = hgrant0_p & v999934 | !hgrant0_p & !v99993c;
assign v8ea84e = hbusreq0_p & v8ea84c | !hbusreq0_p & v8ea84d;
assign v999915 = stateG2_p & v84563c | !stateG2_p & v999914;
assign v8ea86b = hgrant0_p & v8ea866 | !hgrant0_p & v8ea86a;
assign v8ea84f = hlock0 & v8ea84e | !hlock0 & v8ea84a;
assign v9855b4 = hbusreq1_p & v9855b3 | !hbusreq1_p & v84563c;
assign v9d26dc = hgrant2_p & v9d26cf | !hgrant2_p & v9d26db;
assign v8c20d4 = hready_p & v8c20d3 | !hready_p & !v8c20bc;
assign v9d26a9 = stateG2_p & v84563c | !stateG2_p & !v9d26a8;
assign v9d2687 = locked_p & v9d2686 | !locked_p & v84563c;
assign v984ef0 = stateG10_1_p & v984eef | !stateG10_1_p & v985631;
assign v984ec7 = hmaster1_p & v984ec6 | !hmaster1_p & v985643;
assign v9739ab = hmaster0_p & v9738e1 | !hmaster0_p & v973966;
assign v9adc21 = hgrant1_p & v9adbeb | !hgrant1_p & !v9adc1f;
assign v9adc9e = hmaster0_p & v9adc79 | !hmaster0_p & !v9adc77;
assign v9b40c6 = hgrant0_p & v84563c | !hgrant0_p & v9b40c5;
assign v9d26af = hbusreq1_p & v9d26ae | !hbusreq1_p & v84563c;
assign v9adce5 = hmaster0_p & v9adcb5 | !hmaster0_p & !v9adc75;
assign v9a6abe = hmaster0_p & v9a6abd | !hmaster0_p & v84563c;
assign v9855fc = hmaster1_p & v9855fa | !hmaster1_p & v9855fb;
assign v9d2666 = hmastlock_p & v9d2665 | !hmastlock_p & v84563c;
assign a2bd3d = hburst0_p & v84563c | !hburst0_p & a2bd3c;
assign v984f81 = hmaster0_p & v984eac | !hmaster0_p & v984eb3;
assign v97390d = hmaster0_p & v973885 | !hmaster0_p & !v9738dc;
assign v985591 = locked_p & v985590 | !locked_p & v84563c;
assign v9d2679 = hbusreq0 & v9d2677 | !hbusreq0 & v9d2678;
assign v9adc8f = hmaster1_p & v9adc7f | !hmaster1_p & v9adc8a;
assign v9739bc = hbusreq0_p & v9739b9 | !hbusreq0_p & v9739bb;
assign v973a3c = hbusreq0_p & v973a30 | !hbusreq0_p & v973a3b;
assign v9d26b0 = hmaster0_p & v9d26af | !hmaster0_p & !v84563c;
assign v8e79c1 = hmaster0_p & v8e79c0 | !hmaster0_p & v84563c;
assign v9998e0 = hready_p & v9998de | !hready_p & !v9998df;
assign v8c1161 = decide_p & v8c112f | !decide_p & v8c1160;
assign v8c114d = hmaster0_p & v84563c | !hmaster0_p & v8c114c;
assign v9998e3 = hmaster0_p & v9ed40e | !hmaster0_p & v9ed416;
assign v9adcf3 = hready_p & v9adcea | !hready_p & !v9adcf2;
assign v8ea890 = hmaster0_p & v8ea88f | !hmaster0_p & v8ea822;
assign v97398b = hbusreq0_p & v973989 | !hbusreq0_p & v97398a;
assign v973937 = hbusreq2_p & v9738fd | !hbusreq2_p & !v973936;
assign v98550b = hmaster1_p & v985509 | !hmaster1_p & v9854b8;
assign v9adbfd = decide_p & v9adbfc | !decide_p & v9adbf7;
assign v973898 = hbusreq0_p & v973891 | !hbusreq0_p & v973897;
assign v973928 = hbusreq0_p & v973926 | !hbusreq0_p & v973927;
assign v9739af = decide_p & v9739a4 | !decide_p & v9739ae;
assign v984f20 = hbusreq2 & v984ef6 | !hbusreq2 & v84563c;
assign v9965b1 = hbusreq0_p & v9965ae | !hbusreq0_p & v9965b0;
assign v9854eb = stateA1_p & v84563c | !stateA1_p & v9854ea;
assign v9d27bd = hbusreq0 & v9d27bb | !hbusreq0 & !v9d27bc;
assign v8ea8f7 = hgrant2_p & v8ea8e9 | !hgrant2_p & v8ea8f6;
assign a14da7 = hlock0_p & a14da6 | !hlock0_p & !v84563c;
assign v8c116c = decide_p & v8c1169 | !decide_p & v8c116b;
assign v984f86 = hbusreq0 & v984f7d | !hbusreq0 & v984f85;
assign v973903 = hmaster1_p & v973902 | !hmaster1_p & v973890;
assign v973a15 = hbusreq0_p & v973965 | !hbusreq0_p & v973a14;
assign a153ba = hbusreq1_p & a153b7 | !hbusreq1_p & v84563c;
assign v9d275b = hgrant1_p & v845641 | !hgrant1_p & !v9d2691;
assign v9adcf5 = hbusreq2_p & v9adccd | !hbusreq2_p & !v9adcf4;
assign v9ed462 = busreq_p & v9ed45f | !busreq_p & v9ed461;
assign v9ed442 = hbusreq1_p & v973889 | !hbusreq1_p & v84563c;
assign v973995 = hmaster1_p & v97390d | !hmaster1_p & !v973938;
assign v9ed441 = hmaster0_p & v9ed43c | !hmaster0_p & v9ed440;
assign v9998f9 = hmaster1_p & v9998f7 | !hmaster1_p & v9998f8;
assign v9baf94 = hmaster1_p & a154a3 | !hmaster1_p & v9baf93;
assign v985492 = hburst1_p & v9a6a95 | !hburst1_p & v84563c;
assign v9933c4 = hgrant1_p & v9933b7 | !hgrant1_p & !v84563c;
assign v9854cc = decide_p & v9854bb | !decide_p & v9854cb;
assign v985554 = busreq_p & v84563c | !busreq_p & !v985553;
assign v9adc84 = decide_p & v9adc83 | !decide_p & v9adc7e;
assign v984f71 = hmaster0_p & v985642 | !hmaster0_p & v985526;
assign v8ea833 = hbusreq1_p & v8ea832 | !hbusreq1_p & v8ea818;
assign v98558b = stateG2_p & v84563c | !stateG2_p & a153bb;
assign v9ed484 = hmaster1_p & v9ed46f | !hmaster1_p & v9ed483;
assign v8768ab = stateG2_p & v84563c | !stateG2_p & v87bd68;
assign v98553f = hmaster1_p & v84563c | !hmaster1_p & v9854b0;
assign v9998f0 = hmaster0_p & v84565c | !hmaster0_p & !v9998ef;
assign v9baf03 = hburst0 & v9baeff | !hburst0 & v9baf02;
assign v9854ef = busreq_p & v9854ec | !busreq_p & v9854ee;
assign v9999dd = hmaster0_p & v84565c | !hmaster0_p & v9bae80;
assign v9d26ec = hmaster1_p & v9d26eb | !hmaster1_p & !v9d2671;
assign v973a27 = hbusreq0_p & v973989 | !hbusreq0_p & v973a26;
assign v9965ba = hbusreq0_p & v9965b8 | !hbusreq0_p & v9965b9;
assign v9baf12 = hmaster1_p & v9baf05 | !hmaster1_p & !v9baf11;
assign v9a6acd = hmaster0_p & v9a6acc | !hmaster0_p & v84563c;
assign v9adc73 = busreq_p & v84563c | !busreq_p & !v845668;
assign v9ed47c = hburst0_p & v84563c | !hburst0_p & v9ed47b;
assign a153d5 = hmaster0_p & v84563c | !hmaster0_p & a153d3;
assign v9855ad = hgrant1_p & v845641 | !hgrant1_p & !v9855ac;
assign v8ea91f = hbusreq0 & v8ea916 | !hbusreq0 & v8ea91e;
assign v985505 = hlock0_p & v985503 | !hlock0_p & v985504;
assign v973a26 = hmaster1_p & v973902 | !hmaster1_p & v9739e8;
assign v9ed460 = stateA1_p & a153cb | !stateA1_p & a154c2;
assign v9baeaa = hbusreq2 & v9baea3 | !hbusreq2 & v9baea9;
assign v9d27a0 = hbusreq0 & v9d279e | !hbusreq0 & !v9d279f;
assign v9ed421 = hmaster1_p & v9ed418 | !hmaster1_p & v9ed420;
assign v985522 = stateA1_p & v8ea7e2 | !stateA1_p & a153bb;
assign v9ecda4 = hready_p & v9ed56e | !hready_p & v9ecda3;
assign v984f49 = hbusreq0_p & v984f48 | !hbusreq0_p & v985540;
assign v9739d2 = hbusreq0_p & v973903 | !hbusreq0_p & v97398a;
assign v9999d3 = hbusreq0_p & v9999d2 | !hbusreq0_p & v84563c;
assign v984e56 = hbusreq1_p & v984e55 | !hbusreq1_p & v9855af;
assign v9854f5 = stateA1_p & v8ea7e2 | !stateA1_p & v9854f3;
assign v99658f = hbusreq1_p & v996582 | !hbusreq1_p & !v99658e;
assign v9739c6 = hlock2_p & v9739c4 | !hlock2_p & v9739c5;
assign v9998f1 = hmaster1_p & v9998f0 | !hmaster1_p & a154a3;
assign v9a6ab6 = hmaster1_p & v84563c | !hmaster1_p & v9a6a99;
assign v9999d5 = hbusreq2 & v9999b9 | !hbusreq2 & v9999d4;
assign v8ea8dd = hgrant2_p & v8ea7f8 | !hgrant2_p & v8ea8dc;
assign v9855a4 = hbusreq0_p & v9855a3 | !hbusreq0_p & v985595;
assign v9ecda9 = jx1_p & v9ed52c | !jx1_p & v9ecda8;
assign a15446 = decide_p & a15445 | !decide_p & v84565c;
assign a153ce = hlock1_p & v84563c | !hlock1_p & !a153cd;
assign v985649 = hready_p & v98561f | !hready_p & v985648;
assign v8c1130 = stateG3_2_p & v84563c | !stateG3_2_p & !v845658;
assign v9ed4ef = hready_p & v9ed4ed | !hready_p & !v9ed4ee;
assign v97392d = hmaster1_p & v97392b | !hmaster1_p & !v9738dd;
assign v98562d = hmaster1_p & v98562b | !hmaster1_p & !v98562c;
assign a2fb4b = hburst1_p & v84563c | !hburst1_p & !v863b4b;
assign v9baecb = decide_p & v9baeca | !decide_p & !v84563c;
assign v9bae83 = hbusreq1 & v9bae80 | !hbusreq1 & !v9bae82;
assign v9d278a = hgrant2_p & v9d277d | !hgrant2_p & v9d2789;
assign v9baf21 = hmaster1_p & v9baf05 | !hmaster1_p & !v9baf20;
assign v9d271e = hgrant1_p & v84563c | !hgrant1_p & !v9d271d;
assign v8ea8ea = hmaster1_p & v8ea8b4 | !hmaster1_p & v8ea8ca;
assign v984f8b = hgrant2_p & v984f3b | !hgrant2_p & v984f8a;
assign a15491 = hmaster1_p & a1548c | !hmaster1_p & a1548d;
assign v9855af = stateG10_1_p & v84563c | !stateG10_1_p & v9855ae;
assign v9d269a = hgrant0_p & v84563c | !hgrant0_p & v9d2699;
assign v9854e9 = hburst1_p & v8ea7e3 | !hburst1_p & v84563c;
assign v9adc49 = hmaster0_p & v9adc48 | !hmaster0_p & v8ea822;
assign v9b40cc = hready_p & v9b40c6 | !hready_p & !v845654;
assign v984f8d = hready_p & v84563c | !hready_p & v984f8c;
assign v98556c = hmaster0_p & v84563c | !hmaster0_p & !v98556b;
assign v9ed4e3 = hbusreq2 & v9ed4da | !hbusreq2 & v9ed4e2;
assign v8ea888 = hbusreq1_p & v8ea886 | !hbusreq1_p & v8ea887;
assign v9d2673 = hmaster0_p & v845647 | !hmaster0_p & !v84563c;
assign v9998f6 = hbusreq2 & v9998e9 | !hbusreq2 & v9998f5;
assign v9998d6 = hbusreq0 & v9998d4 | !hbusreq0 & v9998d5;
assign a14d85 = hbusreq2_p & a14d5c | !hbusreq2_p & !a14d72;
assign a15496 = hgrant2_p & a15486 | !hgrant2_p & a15495;
assign v9999eb = decide_p & v9999d6 | !decide_p & !v84565e;
assign v9ed4b2 = hmaster0_p & v9ed4ae | !hmaster0_p & v9ed4b1;
assign v9bae90 = hmaster1_p & v9bae8f | !hmaster1_p & v84563c;
assign v9d277a = hbusreq0 & v9d2777 | !hbusreq0 & v9d2779;
assign v973a36 = hmaster1_p & v973a35 | !hmaster1_p & !v973a08;
assign v9d2694 = hgrant1_p & v845647 | !hgrant1_p & v84563c;
assign a154f1 = hbusreq0_p & a154f0 | !hbusreq0_p & v84563c;
assign v8c111c = hmaster1_p & v8c111b | !hmaster1_p & v84563c;
assign v9a6ad1 = hready_p & v9a6ac6 | !hready_p & v9a6ad0;
assign v8ea8f0 = hgrant0_p & v8ea8b7 | !hgrant0_p & v8ea86a;
assign v97388f = hbusreq1_p & v97388c | !hbusreq1_p & v97388e;
assign v9739a1 = hmaster0_p & v97391e | !hmaster0_p & v97395c;
assign v98560b = hlock0_p & v985606 | !hlock0_p & v98560a;
assign v9998a8 = hgrant0_p & v9998a7 | !hgrant0_p & !v84563c;
assign v9739da = hready_p & v9739d3 | !hready_p & v9739d9;
assign v9baf69 = hbusreq1_p & v9baf65 | !hbusreq1_p & v9baf68;
assign v98561c = hmaster1_p & v985619 | !hmaster1_p & v98561b;
assign v9ed4b0 = hlock1_p & v9ed4af | !hlock1_p & !v84565c;
assign v9d271c = hbusreq0_p & v9d271b | !hbusreq0_p & v9d267b;
assign a15421 = hlock1_p & v84563c | !hlock1_p & !a15420;
assign v9999e3 = hbusreq2 & v9999e2 | !hbusreq2 & v9999a6;
assign v8ea8e7 = hbusreq2 & v8ea8e5 | !hbusreq2 & v8ea8e6;
assign v8ea8c7 = jx0_p & v8ea87a | !jx0_p & v8ea8c6;
assign v9854b7 = hbusreq0_p & v9854b5 | !hbusreq0_p & v9854b6;
assign v9a6ac6 = decide_p & v9a6ac0 | !decide_p & v9a6ac5;
assign v9d26c7 = hmaster0_p & v9d26c0 | !hmaster0_p & v84563c;
assign a154a6 = hbusreq0_p & a154a5 | !hbusreq0_p & v84563c;
assign v9739e8 = hmaster0_p & v97393f | !hmaster0_p & v973894;
assign v9adc94 = locked_p & v84563c | !locked_p & !v9adc75;
assign v96ef3e = stateG3_2_p & v84563c | !stateG3_2_p & !v8763e4;
assign v8c112f = hlock2_p & v8c1129 | !hlock2_p & v8c112e;
assign v98558e = stateA1_p & v972fac | !stateA1_p & !v84563c;
assign v98564b = stateG2_p & v98564a | !stateG2_p & !v985535;
assign v996570 = hbusreq0_p & v99656e | !hbusreq0_p & v99656f;
assign v8ea8e0 = hmaster1_p & v8ea8de | !hmaster1_p & v8ea7f4;
assign v8ea851 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea833;
assign v985496 = hmastlock_p & v985495 | !hmastlock_p & v84563c;
assign v9ed4fb = hgrant1_p & a153c0 | !hgrant1_p & !v84563c;
assign v8ea7f6 = hbusreq0_p & v8ea7f3 | !hbusreq0_p & v8ea7f5;
assign v9baf85 = hbusreq0_p & v9baf84 | !hbusreq0_p & !v84563c;
assign v9ed42d = hburst1_p & v84563c | !hburst1_p & !v8e798b;
assign v985578 = locked_p & v985577 | !locked_p & !v84563c;
assign v8e798b = stateG3_2_p & v84563c | !stateG3_2_p & v8e798a;
assign v9d27b2 = hready_p & v9d27a8 | !hready_p & !v9d27b1;
assign v8c20dc = hbusreq0_p & v8c20c5 | !hbusreq0_p & v8c20db;
assign a15517 = decide_p & a1550e | !decide_p & v84565c;
assign v9738d1 = hgrant1_p & v9738c4 | !hgrant1_p & v97388d;
assign v99992c = hlock0_p & v99992b | !hlock0_p & v999925;
assign v985547 = busreq_p & v985495 | !busreq_p & v985546;
assign v9739fc = decide_p & v9739f9 | !decide_p & v9739fb;
assign v985537 = busreq_p & v9a6a96 | !busreq_p & v985536;
assign v98551c = hbusreq0_p & v98551b | !hbusreq0_p & v98551a;
assign a14d4a = hready_p & a14d3f | !hready_p & a14d49;
assign v9d267f = hmaster1_p & v84563c | !hmaster1_p & !v9d2673;
assign v984eca = decide_p & v98563f | !decide_p & v984ec9;
assign v9a6ade = hgrant0_p & v9a6ab8 | !hgrant0_p & v9a6add;
assign a153c3 = hmaster0_p & a153ba | !hmaster0_p & a153c2;
assign v8e7999 = stateG2_p & v84563c | !stateG2_p & v8e7998;
assign v985558 = hbusreq1_p & v985557 | !hbusreq1_p & v84563c;
assign v9d267e = hmaster1_p & v84563c | !hmaster1_p & !v9d2671;
assign v984f4a = hgrant0_p & v984f49 | !hgrant0_p & v984f41;
assign v8c1141 = hbusreq0_p & v8c1140 | !hbusreq0_p & v84563c;
assign v97388d = hmastlock_p & v87f892 | !hmastlock_p & v84563c;
assign v973a49 = hbusreq2_p & v973a20 | !hbusreq2_p & !v973a48;
assign v9855d1 = hmaster1_p & v985491 | !hmaster1_p & v985531;
assign a14d8e = hmaster1_p & a153cd | !hmaster1_p & !a14d8d;
assign v973963 = hbusreq1_p & v9738ce | !hbusreq1_p & !v973962;
assign v9ed4c2 = hbusreq0_p & v9ed4bc | !hbusreq0_p & !v9ed4c1;
assign v8ea866 = hbusreq0_p & v8ea864 | !hbusreq0_p & v8ea865;
assign v984f42 = hgrant0_p & v984f3e | !hgrant0_p & v984f41;
assign v9738ec = hbusreq1_p & v9738d6 | !hbusreq1_p & v9738eb;
assign v99993c = hbusreq0_p & v99993b | !hbusreq0_p & v84563c;
assign v996594 = hbusreq0_p & v996591 | !hbusreq0_p & v996593;
assign v8c1135 = busreq_p & v8c1133 | !busreq_p & !v8c1134;
assign v9baeee = decide_p & v9baeca | !decide_p & v84563c;
assign v9adce7 = hmaster1_p & v9adce5 | !hmaster1_p & !v9adcbc;
assign v9d2757 = hmaster1_p & v9d26fc | !hmaster1_p & v845647;
assign v9baf5f = locked_p & v84563c | !locked_p & !v97388d;
assign v8ea899 = hbusreq0_p & v8ea898 | !hbusreq0_p & v8ea82e;
assign v9999b9 = hbusreq0_p & v9999b8 | !hbusreq0_p & v84563c;
assign v985510 = hlock0_p & v98550e | !hlock0_p & v98550f;
assign v99657d = hlock0_p & v99657a | !hlock0_p & v99657c;
assign v9adbf2 = hbusreq1_p & v9adbf1 | !hbusreq1_p & v9adbee;
assign a14dbe = hgrant2_p & a14da4 | !hgrant2_p & a14dba;
assign v8ea825 = hgrant1_p & v8ea818 | !hgrant1_p & v8ea7e9;
assign a14d8c = hmaster1_p & a153cd | !hmaster1_p & !a14d8b;
assign v8c1171 = hburst0_p & v84563c | !hburst0_p & v8c1170;
assign v996596 = decide_p & v99658c | !decide_p & v996595;
assign v999905 = stateG2_p & v87f892 | !stateG2_p & !v999904;
assign v9965ab = hmaster0_p & v9adbfe | !hmaster0_p & v8ea7e9;
assign v9ed531 = decide_p & v9ed4f7 | !decide_p & v9ed4c6;
assign v9adca5 = hgrant1_p & v9adc76 | !hgrant1_p & !v9adc75;
assign v8ea8b9 = hmaster1_p & v8ea8b8 | !hmaster1_p & v8ea890;
assign v984f28 = hlock0_p & v984f25 | !hlock0_p & v984f27;
assign v999933 = hlock0_p & v84565c | !hlock0_p & !v84563c;
assign v9adbf0 = hmaster0_p & v9adbec | !hmaster0_p & v9adbef;
assign v8ea8c5 = hgrant2_p & v8ea8b3 | !hgrant2_p & v8ea8c4;
assign v984e74 = hmaster1_p & v984e69 | !hmaster1_p & v984e73;
assign v9a6ab3 = hmaster1_p & v9a6ab2 | !hmaster1_p & v84563c;
assign v9ed4bc = hlock0_p & v9ed4b9 | !hlock0_p & !v9ed4bb;
assign a153ea = hbusreq0_p & a153e9 | !hbusreq0_p & a153e8;
assign v984ed9 = hbusreq0_p & v984ed8 | !hbusreq0_p & v985645;
assign v8ea895 = stateG10_1_p & v84563c | !stateG10_1_p & v8ea7e9;
assign v98552f = hready_p & v9854cc | !hready_p & v98552e;
assign v8ea910 = hbusreq0_p & v8ea90d | !hbusreq0_p & v8ea90f;
assign v8e79c4 = hbusreq1_p & v8e79c2 | !hbusreq1_p & v8e79c3;
assign v9adca2 = hmaster0_p & v9adc79 | !hmaster0_p & !v9adca1;
assign v9738c5 = hbusreq1_p & v9738c3 | !hbusreq1_p & v9738c4;
assign v984eb5 = hmaster1_p & v984eb4 | !hmaster1_p & v984ead;
assign v98554e = hready & v985549 | !hready & !v98554d;
assign v99991d = hlock0_p & v99991a | !hlock0_p & v99991c;
assign v973a39 = hbusreq0_p & v973a36 | !hbusreq0_p & v973a38;
assign v985640 = hlock2_p & v985639 | !hlock2_p & v98563f;
assign v9965a1 = hbusreq0_p & v99659e | !hbusreq0_p & v9965a0;
assign v9a6adb = hmaster0_p & v9a6ada | !hmaster0_p & v84563c;
assign v9854f9 = hready & v9854f6 | !hready & v9854f8;
assign v999910 = hbusreq0_p & v99990f | !hbusreq0_p & !v84563c;
assign v9738a6 = hlock1_p & v9738a4 | !hlock1_p & v973889;
assign v9baf75 = hbusreq0_p & v9baf6b | !hbusreq0_p & v9baf74;
assign v984e65 = hbusreq0 & v984e64 | !hbusreq0 & v84563c;
assign v8ea826 = stateG10_1_p & v8ea7ea | !stateG10_1_p & !v8ea825;
assign v9ed475 = hburst0 & v973892 | !hburst0 & v9ed474;
assign v9adbf9 = locked_p & v9adbf8 | !locked_p & v9adbee;
assign v9999c4 = hmastlock_p & v9999c3 | !hmastlock_p & v84563c;
assign v996555 = hmaster1_p & v996550 | !hmaster1_p & v996554;
assign v9d269b = hgrant0_p & v84563c | !hgrant0_p & !v9d2699;
assign v8ea80f = stateA1_p & v84566e | !stateA1_p & !v84563c;
assign v9738bb = decide_p & v9738b6 | !decide_p & v9738ba;
assign v984f4c = hbusreq2 & v984f4b | !hbusreq2 & v84563c;
assign a1542f = hgrant0_p & a15416 | !hgrant0_p & a1542e;
assign v9ed4fa = hready_p & v84563c | !hready_p & v9ed4f9;
assign v973888 = hmastlock_p & v973887 | !hmastlock_p & !v84563c;
assign v985598 = hbusreq1_p & v985597 | !hbusreq1_p & v845641;
assign v984ec5 = decide_p & v985610 | !decide_p & v984ec4;
assign v984f64 = hbusreq0_p & v984f61 | !hbusreq0_p & v984f63;
assign v985561 = hburst0_p & a3134f | !hburst0_p & v9854bd;
assign a14d5d = decide_p & v84563c | !decide_p & !v84565c;
assign a153bd = hmastlock_p & a153bc | !hmastlock_p & v84563c;
assign v9ed500 = hbusreq0_p & v9ed4ff | !hbusreq0_p & v9ed4b4;
assign a15483 = hmaster1_p & a15448 | !hmaster1_p & a15449;
assign v8ea89a = hgrant0_p & v8ea884 | !hgrant0_p & v8ea899;
assign v996585 = stateG10_1_p & v9adbee | !stateG10_1_p & !v996584;
assign v8c1166 = hbusreq1_p & v8c1120 | !hbusreq1_p & v8c1139;
assign v8e79cf = hbusreq0_p & v8e79a6 | !hbusreq0_p & v8e79ce;
assign v9bae7f = hmastlock_p & v9bae7e | !hmastlock_p & v84563c;
assign v8c1125 = hmaster1_p & v8c1121 | !hmaster1_p & v8c1124;
assign v9738e7 = hbusreq1_p & v9738ce | !hbusreq1_p & !v9738e6;
assign hgrant1 = !v9ecda9;
assign a14d67 = hbusreq0_p & v84563c | !hbusreq0_p & a14d40;
assign v985615 = stateG2_p & v84563c | !stateG2_p & v985614;
assign v9d44bf = jx0_p & v854658 | !jx0_p & v84563c;
assign v9854d6 = hlock0_p & v9854d4 | !hlock0_p & v9854d5;
assign v8c20b7 = hmaster1_p & v8c20b6 | !hmaster1_p & v84563c;
assign v996579 = hmaster0_p & v996553 | !hmaster0_p & !v99654f;
assign v9d276a = hbusreq2 & v9d2763 | !hbusreq2 & v9d2769;
assign v8ea8d2 = hmaster0_p & v8ea8cf | !hmaster0_p & v8ea82c;
assign v973a08 = hmaster0_p & v973a07 | !hmaster0_p & !v9738cc;
assign v985580 = hmaster1_p & v98557e | !hmaster1_p & v98557f;
assign v99999d = hbusreq2_p & v99996b | !hbusreq2_p & v99999c;
assign v9999b2 = decide_p & v9999b1 | !decide_p & v84565e;
assign v9adc42 = hmaster0_p & v9adc11 | !hmaster0_p & v8ea7ef;
assign v98555f = hmaster0_p & v84563c | !hmaster0_p & v9854c5;
assign v9999d1 = hmaster1_p & v84563c | !hmaster1_p & v9baeb2;
assign v973943 = decide_p & v97393e | !decide_p & v973942;
assign v9adc28 = hmaster0_p & v9adc24 | !hmaster0_p & v9adc27;
assign v973930 = hmaster1_p & v97392f | !hmaster1_p & v9738e8;
assign v85bb54 = hmaster1_p & v845652 | !hmaster1_p & v84563c;
assign v9baf6a = hmaster0_p & v9baf63 | !hmaster0_p & v9baf69;
assign v996582 = hgrant1_p & v99654f | !hgrant1_p & !v9adbee;
assign v9baea4 = hmaster0_p & v84565c | !hmaster0_p & !v9bae82;
assign v9ed497 = hready_p & v9ed453 | !hready_p & !v9ed496;
assign v8ea8a4 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea818;
assign v8ea912 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea832;
assign v9adc02 = hbusreq1_p & v9adc00 | !hbusreq1_p & v9adc01;
assign v9854ad = hready & v98549d | !hready & v9854ac;
assign v9965bb = hmaster0_p & v9adc24 | !hmaster0_p & v996552;
assign v9adcdc = hmaster1_p & v9adcdb | !hmaster1_p & !v9adcae;
assign v9baf30 = hmastlock_p & v9ed46c | !hmastlock_p & !v84563c;
assign v9998d9 = hbusreq0_p & v9998a6 | !hbusreq0_p & !v854658;
assign v8e79c8 = decide_p & v8e79a8 | !decide_p & v8e79c7;
assign a14dc1 = jx0_p & a14d85 | !jx0_p & a14dc0;
assign v9a6abb = hgrant1_p & v9a6a98 | !hgrant1_p & v84563c;
assign v9855e0 = hmaster0_p & v98557b | !hmaster0_p & v985582;
assign v9933bd = hmaster1_p & v84563c | !hmaster1_p & v9933b8;
assign v996564 = hmaster0_p & v996563 | !hmaster0_p & v9adbfe;
assign v973929 = hgrant0_p & v973924 | !hgrant0_p & v973928;
assign a154fb = hgrant1_p & v84563c | !hgrant1_p & a15420;
assign v8ea92a = hbusreq2_p & v8ea924 | !hbusreq2_p & v8ea929;
assign v9d2789 = hready_p & v9d2787 | !hready_p & v9d2788;
assign v9ed4cc = hmaster1_p & v9ed4cb | !hmaster1_p & v9ed443;
assign v985585 = hbusreq0_p & v985580 | !hbusreq0_p & v985584;
assign v9d2769 = hbusreq0 & v9d2766 | !hbusreq0 & v9d2768;
assign v97391c = hgrant1_p & v973885 | !hgrant1_p & v97391b;
assign v9baf2f = hmastlock_p & v9baf2e | !hmastlock_p & v84563c;
assign v9ed412 = stateG2_p & v84563c | !stateG2_p & v9ed411;
assign v9baf46 = hmaster0_p & v973885 | !hmaster0_p & v84563c;
assign v97392b = hmaster0_p & v973885 | !hmaster0_p & !v973895;
assign v8c20d7 = hgrant1_p & v84565c | !hgrant1_p & !v84563c;
assign v9adc60 = stateG2_p & v84563c | !stateG2_p & !v9adbf8;
assign v97398c = decide_p & v973988 | !decide_p & !v97398b;
assign v98554a = stateA1_p & v8e7990 | !stateA1_p & a1541d;
assign v9adc97 = hmaster1_p & v9adc93 | !hmaster1_p & !v9adc96;
assign v9ed42b = locked_p & v9ed42a | !locked_p & !v84563c;
assign v985539 = hready & v985538 | !hready & !v84563c;
assign v9965cc = hbusreq0_p & v9965ca | !hbusreq0_p & v9965cb;
assign v8ea83d = hgrant0_p & v8ea83c | !hgrant0_p & v8ea82f;
assign v8ea8b0 = hlock2 & v8ea8a7 | !hlock2 & v8ea8ae;
assign v9738ab = hmaster1_p & v9738a5 | !hmaster1_p & v9738aa;
assign v9ed4ec = hbusreq0 & v9ed4eb | !hbusreq0 & v9ed4c3;
assign v9ed49e = hbusreq1_p & v9ed49d | !hbusreq1_p & !v84563c;
assign v9baf64 = hbusreq1 & v9ed419 | !hbusreq1 & v84565c;
assign v9738fc = hready_p & v9738f1 | !hready_p & !v9738fb;
assign v9d27c1 = hbusreq2_p & v9d27b3 | !hbusreq2_p & v9d27c0;
assign v9baf07 = hburst1 & v87f892 | !hburst1 & !v84563c;
assign v984f59 = hmaster1_p & a154a3 | !hmaster1_p & v984f58;
assign v8ea8b3 = hready_p & v8ea846 | !hready_p & v8ea8b2;
assign v9965a2 = hgrant0_p & v996598 | !hgrant0_p & v9965a1;
assign v99656b = hbusreq0_p & v996568 | !hbusreq0_p & v99656a;
assign v99993b = hlock0_p & v999937 | !hlock0_p & v99993a;
assign v9adbec = locked_p & v9adbe9 | !locked_p & v9adbeb;
assign v97397b = hmaster0_p & v97393f | !hmaster0_p & !v97388a;
assign v9adceb = hmaster0_p & v9adc75 | !hmaster0_p & !v9adc94;
assign v9baf09 = hmastlock_p & v9baf08 | !hmastlock_p & v84563c;
assign v9d2759 = hgrant0_p & v84563c | !hgrant0_p & !v9d2757;
assign v97395b = hbusreq0_p & v9738c2 | !hbusreq0_p & !v97395a;
assign v9999d8 = hready_p & v84563c | !hready_p & v9999d7;
assign v9ecda8 = jx0_p & v9ed533 | !jx0_p & v9ecda7;
assign v9739e6 = hgrant2_p & v9739da | !hgrant2_p & !v9739e5;
assign v985630 = hbusreq0 & v98562f | !hbusreq0 & v84563c;
assign v9a6aa2 = hmastlock_p & v9a6aa1 | !hmastlock_p & v84563c;
assign v9ed437 = hmaster0_p & v9ed423 | !hmaster0_p & v9ed436;
assign v973965 = hmaster1_p & v9738e4 | !hmaster1_p & !v973964;
assign v8ea938 = hgrant2_p & v8ea7f8 | !hgrant2_p & v8ea937;
assign v9adca7 = hbusreq1_p & v9adca6 | !hbusreq1_p & !v9adc75;
assign v9ed56e = decide_p & v9ed56a | !decide_p & v9ed4c6;
assign v9d26ea = hbusreq0 & v9d26e6 | !hbusreq0 & v9d26e9;
assign v973980 = hbusreq0_p & v97397e | !hbusreq0_p & v97397f;
assign v8e7988 = stateG3_0_p & v84566c | !stateG3_0_p & !v84566c;
assign v98557f = hmaster0_p & v84563c | !hmaster0_p & v98557d;
assign v9b40c1 = hgrant0_p & v84563c | !hgrant0_p & v845660;
assign v9739c9 = hready_p & v9739c3 | !hready_p & !v9739c8;
assign v9738db = hgrant0_p & v9738c8 | !hgrant0_p & v9738da;
assign v9854c6 = hmaster0_p & v9ed423 | !hmaster0_p & v9854c5;
assign v9d266c = busreq_p & v9d266a | !busreq_p & v9d266b;
assign v973894 = locked_p & v84563c | !locked_p & v973893;
assign v9d276e = hbusreq1_p & v84563c | !hbusreq1_p & !v845641;
assign a154d6 = hlock0_p & v84563c | !hlock0_p & !a154d5;
assign v9d27ba = hbusreq0_p & v845647 | !hbusreq0_p & v9d2738;
assign v9855b9 = hbusreq0 & v98559d | !hbusreq0 & v9855b8;
assign v9854f0 = hmastlock_p & v9854ef | !hmastlock_p & v84563c;
assign v9ed52c = jx0_p & v9ed4f1 | !jx0_p & v9ed522;
assign v973897 = hmaster1_p & v97388b | !hmaster1_p & v973896;
assign v9738ee = hmaster1_p & v9738e4 | !hmaster1_p & !v9738ed;
assign v999913 = hbusreq0 & v999910 | !hbusreq0 & !v999912;
assign v9a6ab5 = hready_p & v9a6a9c | !hready_p & v9a6ab4;
assign v9999e1 = hgrant0_p & v9999e0 | !hgrant0_p & !v84563c;
assign v9ed520 = decide_p & v9ed4f8 | !decide_p & v9ed4c6;
assign v984eb1 = hbusreq0 & v984eb0 | !hbusreq0 & v985645;
assign v8ea7ed = hmaster0_p & v8ea7ec | !hmaster0_p & v8ea7e9;
assign a14d3f = decide_p & a14d3e | !decide_p & v84565c;
assign v9739c2 = jx0_p & v973937 | !jx0_p & v9739c1;
assign v8ea8b7 = hbusreq0_p & v8ea8b5 | !hbusreq0_p & v8ea8b6;
assign v9baf44 = hmaster0_p & v9baf43 | !hmaster0_p & v9ed416;
assign v98551e = hbusreq2 & v985512 | !hbusreq2 & v98551d;
assign a1540b = hlock2_p & a153ea | !hlock2_p & a1540a;
assign v8ea922 = decide_p & v8ea7ee | !decide_p & v8ea921;
assign a14d72 = hgrant2_p & a14d6d | !hgrant2_p & !a14d71;
assign v8e79b7 = hmaster1_p & v8e79b2 | !hmaster1_p & v8e79b6;
assign v9d26b5 = hbusreq0 & v9d26b2 | !hbusreq0 & v9d26b4;
assign v8c1176 = hgrant1_p & v84563c | !hgrant1_p & !v8c1175;
assign v9adc8b = hmaster1_p & v9adc75 | !hmaster1_p & v9adc8a;
assign v9adcc9 = hbusreq0_p & v9adcc3 | !hbusreq0_p & v9adcc8;
assign v92337e = stateG2_p & v84563c | !stateG2_p & v883467;
assign v9a6ad6 = hmaster1_p & v9a6ad5 | !hmaster1_p & v9a6aa7;
assign v9adcd1 = hbusreq0_p & v9adccf | !hbusreq0_p & v9adcd0;
assign v98550d = hbusreq0_p & v98550c | !hbusreq0_p & v98550b;
assign v9bae80 = locked_p & v9bae7f | !locked_p & !v84563c;
assign v97390f = hmaster1_p & v97390d | !hmaster1_p & !v973896;
assign v8ea8e8 = decide_p & v8ea7ee | !decide_p & v8ea8e7;
assign v9998f5 = hbusreq0 & v9998f4 | !hbusreq0 & v84563c;
assign v9739f6 = hbusreq0_p & v97394a | !hbusreq0_p & v9739f5;
assign v9998de = decide_p & v9998dd | !decide_p & v84565e;
assign v9d26c2 = hmaster1_p & v9d26c1 | !hmaster1_p & !v9d2671;
assign v8ea8be = hgrant0_p & v8ea8b7 | !hgrant0_p & v8ea8bd;
assign v8ea930 = hready_p & v8ea80d | !hready_p & v8ea92f;
assign v9ed4ce = hbusreq0_p & v9ed4cc | !hbusreq0_p & v9ed4cd;
assign v98553a = hgrant1_p & v84563c | !hgrant1_p & v985539;
assign v845668 = stateG2_p & v84563c | !stateG2_p & !v84563c;
assign v8c1169 = hbusreq0_p & v8c112d | !hbusreq0_p & v8c1168;
assign a15415 = hlock0_p & a15414 | !hlock0_p & v845648;
assign a14dae = hlock2_p & v84563c | !hlock2_p & a14dad;
assign v8c1138 = busreq_p & v8c1133 | !busreq_p & !v8c1137;
assign v9adc22 = hlock1_p & v9adc20 | !hlock1_p & v9adc21;
assign v9ed423 = hbusreq1_p & v84565c | !hbusreq1_p & v84563c;
assign v9998fd = hlock0_p & v9998fc | !hlock0_p & v84563c;
assign v9a6acf = hgrant0_p & v9a6ac7 | !hgrant0_p & v9a6ace;
assign a15488 = hbusreq1_p & a15421 | !hbusreq1_p & !v84563c;
assign v9ed487 = hmastlock_p & v9ed486 | !hmastlock_p & v84563c;
assign v9739a9 = hmaster0_p & v9738e1 | !hmaster0_p & v9739a8;
assign v9adc4e = hmaster1_p & v9adc49 | !hmaster1_p & !v9adc4d;
assign a154c2 = hburst0_p & v863b4b | !hburst0_p & a154c1;
assign v9855c0 = hbusreq2 & v9855bf | !hbusreq2 & v9854b9;
assign v9a6aaa = hbusreq0_p & v9a6aa9 | !hbusreq0_p & v9a6aa8;
assign v984eac = hbusreq1_p & v984ea9 | !hbusreq1_p & !v984eab;
assign v99656e = hlock0_p & v99656c | !hlock0_p & v99656d;
assign v9baf7b = hlock0_p & v9baf78 | !hlock0_p & !v9baf7a;
assign v999903 = hburst0_p & v85a40d | !hburst0_p & v999902;
assign v97394b = hmaster0_p & v9738a7 | !hmaster0_p & !v97388d;
assign v98563e = hbusreq0_p & v98563d | !hbusreq0_p & v84563c;
assign v9738bf = hmaster1_p & v9738bd | !hmaster1_p & v9738be;
assign v99659a = hgrant1_p & v996572 | !hgrant1_p & v8ea7e9;
assign v9998d8 = hready_p & v9998d3 | !hready_p & v9998d7;
assign v9855f7 = hready_p & v9855e5 | !hready_p & v9855f6;
assign v9739d7 = hbusreq0_p & v9739d6 | !hbusreq0_p & v973992;
assign v8c20cb = hgrant1_p & v8c20ba | !hgrant1_p & !v845656;
assign v99989f = hmaster1_p & v84563c | !hmaster1_p & v9bae95;
assign v9d273e = decide_p & v9d273d | !decide_p & v9d270a;
assign v9739ce = hgrant0_p & v9738f5 | !hgrant0_p & v9739cd;
assign v985636 = hlock0_p & v985633 | !hlock0_p & !v985635;
assign v9d27a5 = hgrant0_p & v84563c | !hgrant0_p & !v9d27a3;
assign v9ed456 = stateA1_p & v84563c | !stateA1_p & !v9ed455;
assign a1540c = decide_p & a1540b | !decide_p & v84565c;
assign v9998cd = decide_p & v9998a2 | !decide_p & !v84565e;
assign v9adce1 = hmaster0_p & v9adce0 | !hmaster0_p & !v9adc75;
assign v8ea848 = hmaster1_p & v8ea847 | !hmaster1_p & v8ea7f2;
assign v984f78 = hmaster1_p & v984f76 | !hmaster1_p & v984f77;
assign v8ea907 = stateG10_1_p & v8ea7e9 | !stateG10_1_p & v8ea906;
assign v845642 = hbusreq0_p & v84563c | !hbusreq0_p & !v84563c;
assign v9ed472 = hmaster0_p & v9ed471 | !hmaster0_p & !v9ed46e;
assign v8ea8cf = hbusreq1_p & v8ea7e9 | !hbusreq1_p & !v8ea8ce;
assign v97389f = hmaster0_p & v97389b | !hmaster0_p & !v97389e;
assign v8ea86d = hbusreq0_p & v8ea864 | !hbusreq0_p & v8ea86c;
assign v9999d0 = hbusreq2 & v9999cb | !hbusreq2 & v9999a2;
assign v9d26f1 = hbusreq0 & v9d26f0 | !hbusreq0 & v9d267f;
assign v9855bc = hready_p & v985587 | !hready_p & v9855bb;
assign v984f67 = decide_p & v984f55 | !decide_p & v984f66;
assign v9adcca = hgrant0_p & v9adcc2 | !hgrant0_p & v9adcc9;
assign v9baf32 = hbusreq1_p & v9baf31 | !hbusreq1_p & !v84563c;
assign v9854ac = hmastlock_p & v9ed411 | !hmastlock_p & v84563c;
assign v9bae95 = hmaster0_p & v84563c | !hmaster0_p & !v9bae94;
assign v9baf02 = hburst1 & v9baeff | !hburst1 & v9baf01;
assign v9965be = hmaster1_p & v9965bd | !hmaster1_p & !v996589;
assign v9ed44c = locked_p & v9ed44b | !locked_p & v84563c;
assign a1542d = hmaster0_p & a15422 | !hmaster0_p & a153ba;
assign v8e79c6 = hmaster1_p & v8e79c1 | !hmaster1_p & v8e79c5;
assign v8ea807 = hmaster1_p & v8ea801 | !hmaster1_p & v8ea806;
assign v9d2730 = hbusreq0_p & v9d26e4 | !hbusreq0_p & v9d267b;
assign v973932 = hbusreq0_p & v973930 | !hbusreq0_p & v973931;
assign v973a2f = hmaster0_p & v973886 | !hmaster0_p & v973894;
assign v9ed455 = hburst0_p & v863b4b | !hburst0_p & v9ed454;
assign v973a42 = hbusreq0_p & v9739b4 | !hbusreq0_p & v973a41;
assign v8ea817 = hmaster1_p & v8ea815 | !hmaster1_p & v8ea816;
assign v9933c8 = hmaster1_p & v9933c3 | !hmaster1_p & !v9933c7;
assign v9baf0d = hbusreq1 & v9baf09 | !hbusreq1 & v9baf0c;
assign v8ea81f = hbusreq0_p & v8ea817 | !hbusreq0_p & v8ea81e;
assign v9738b6 = hlock2_p & v9738af | !hlock2_p & v9738b5;
assign v973953 = hlock2_p & v97394d | !hlock2_p & v973952;
assign v984f60 = hmaster0_p & v984f5f | !hmaster0_p & v984e68;
assign v9baf92 = hgrant0_p & v9baf85 | !hgrant0_p & v9baf90;
assign v9baf14 = hmaster1_p & v9baf05 | !hmaster1_p & !v9baf13;
assign v973956 = hbusreq0_p & v973954 | !hbusreq0_p & v973955;
assign v9933cd = hmaster1_p & v9933c3 | !hmaster1_p & !v9933cc;
assign v973984 = hgrant2_p & v973958 | !hgrant2_p & v973983;
assign v9855dd = hmaster1_p & v9ed423 | !hmaster1_p & v98555f;
assign v999983 = decide_p & v999982 | !decide_p & !v84563c;
assign v9739cf = decide_p & v9739c6 | !decide_p & v9739ce;
assign v9baef0 = hgrant2_p & v9baecc | !hgrant2_p & !v9baeef;
assign v9998a0 = hlock0_p & v99989f | !hlock0_p & v84563c;
assign v9ed478 = hmaster0_p & v9ed471 | !hmaster0_p & v9ed477;
assign v9998ee = hmastlock_p & v9998ed | !hmastlock_p & !v84563c;
assign v973923 = hmaster1_p & v973913 | !hmaster1_p & v9738dd;
assign v8ea8a8 = hlock0 & v8ea8a7 | !hlock0 & v8ea8a6;
assign v9ed4b4 = hbusreq1_p & v9ed4b3 | !hbusreq1_p & !v84563c;
assign v9baefe = stateG2_p & v87f892 | !stateG2_p & v9ed458;
assign v98549a = hburst0_p & v84566a | !hburst0_p & v985499;
assign v97398f = hmaster1_p & v97398d | !hmaster1_p & v973948;
assign v9855ed = hgrant0_p & v9855ec | !hgrant0_p & v98559c;
assign v9d2797 = hmaster1_p & v9d2796 | !hmaster1_p & v9d26fa;
assign v985600 = hlock0_p & v9855fc | !hlock0_p & v9855ff;
assign v99657a = hmaster1_p & v9adc17 | !hmaster1_p & v996579;
assign v9adce8 = hbusreq0_p & v9adce6 | !hbusreq0_p & v9adce7;
assign v8c1153 = hmaster0_p & v8c1152 | !hmaster0_p & !v84563c;
assign v9855da = hgrant0_p & v9855d6 | !hgrant0_p & v9855d9;
assign v9adc36 = stateG10_1_p & v9adbee | !stateG10_1_p & v9adc25;
assign v9ed4aa = hburst0 & v9ed4a2 | !hburst0 & v9ed4a9;
assign v9d273b = hbusreq0_p & v9d2702 | !hbusreq0_p & v9d2738;
assign v9d26ac = locked_p & v84563c | !locked_p & !v9d26ab;
assign v9738e1 = hbusreq1_p & v9738c9 | !hbusreq1_p & !v9738e0;
assign v8ea82e = hmaster1_p & v8ea823 | !hmaster1_p & v8ea82d;
assign v9d2736 = hbusreq1_p & v845647 | !hbusreq1_p & !v9d26d1;
assign v9d2777 = hbusreq0_p & v9d274c | !hbusreq0_p & v9d2776;
assign v8e79ba = hbusreq1_p & v8e79b3 | !hbusreq1_p & v8e79b9;
assign v9adca0 = hlock0_p & v9adc9f | !hlock0_p & !v9adc80;
assign v9ed419 = locked_p & v84563c | !locked_p & v973889;
assign v9d2663 = busreq_p & v845668 | !busreq_p & v9d2662;
assign v9bae7d = hburst1 & v9ed42c | !hburst1 & v9bae7c;
assign v9999ad = hbusreq0 & v9999ac | !hbusreq0 & v99997b;
assign v9adcec = hmaster1_p & v9adceb | !hmaster1_p & !v9adcc1;
assign v973a23 = hmaster1_p & v973a22 | !hmaster1_p & v9739ec;
assign v9ed4d4 = hmaster1_p & v9ed4d3 | !hmaster1_p & v9ed472;
assign v973a22 = hmaster0_p & v973885 | !hmaster0_p & !v9738c3;
assign v984e61 = hmaster1_p & v984e5e | !hmaster1_p & v984e60;
assign v9d26f4 = decide_p & v9d26f2 | !decide_p & v9d2681;
assign v9738b9 = hmaster1_p & v9738b7 | !hmaster1_p & !v973896;
assign v8c20c4 = hmaster0_p & v84565c | !hmaster0_p & v8c20c3;
assign a15444 = hmaster1_p & a15433 | !hmaster1_p & !a15434;
assign v9adcb3 = hgrant0_p & v9adca4 | !hgrant0_p & v9adcb2;
assign a154fe = hmaster0_p & a154fd | !hmaster0_p & v8c20c3;
assign v973a32 = hlock0_p & v973a30 | !hlock0_p & !v973a31;
assign v8ea8f3 = hlock2 & v8ea8f0 | !hlock2 & v8ea8f2;
assign v985608 = hready & v985607 | !hready & v9854ac;
assign v985573 = hmastlock_p & v985572 | !hmastlock_p & !v84563c;
assign v9adcbb = hmaster1_p & v9adcb6 | !hmaster1_p & !v9adcba;
assign a1550c = hbusreq0_p & a1550b | !hbusreq0_p & v84563c;
assign v99998b = hbusreq0_p & v845644 | !hbusreq0_p & v84563c;
assign v8ea8de = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea8c9;
assign v8e79be = decide_p & v8e79b8 | !decide_p & v8e79bd;
assign v9738c2 = hlock0_p & v9738bf | !hlock0_p & !v9738c1;
assign a153d1 = hmastlock_p & a153d0 | !hmastlock_p & !v84563c;
assign v8ea7f1 = hbusreq1_p & v8ea7ef | !hbusreq1_p & v8ea7f0;
assign v999937 = hmaster1_p & v999935 | !hmaster1_p & v999936;
assign v9a6adf = decide_p & v9a6ade | !decide_p & v9a6ac5;
assign v9933bf = hbusreq0_p & v9933be | !hbusreq0_p & v8c20be;
assign v9d26cd = hbusreq2 & v9d26c6 | !hbusreq2 & v9d26cc;
assign v8e79af = hlock0_p & v8e79ae | !hlock0_p & v84563c;
assign v98556e = hbusreq0_p & v985560 | !hbusreq0_p & v98556d;
assign v985516 = hlock0_p & v985514 | !hlock0_p & v985515;
assign v9baea6 = hlock0_p & v9baea5 | !hlock0_p & a154a4;
assign v97397e = hmaster1_p & v9738f6 | !hmaster1_p & v973964;
assign v9baf9f = jx2_p & v9baf9e | !jx2_p & v9baefd;
assign v8e7992 = hmastlock_p & v8e7991 | !hmastlock_p & v84563c;
assign v9d26d3 = hmaster0_p & v9d26d2 | !hmaster0_p & v9d2696;
assign v8c20bd = hready_p & v8c20b9 | !hready_p & v8c20bc;
assign v996586 = hbusreq1_p & v996583 | !hbusreq1_p & !v996585;
assign v8e79aa = hmaster0_p & v84563c | !hmaster0_p & v8e79a9;
assign v996567 = hmaster1_p & v9adbfe | !hmaster1_p & v996566;
assign v9baf5c = locked_p & v9baf5b | !locked_p & !v84563c;
assign v9d26ee = hmaster1_p & v9d26ed | !hmaster1_p & !v9d2671;
assign v9ed4d5 = hmaster1_p & v9ed4d3 | !hmaster1_p & v9ed478;
assign v985542 = hbusreq0_p & v985541 | !hbusreq0_p & v985540;
assign v9adc53 = decide_p & v9adbfb | !decide_p & v9adbf7;
assign v9ed567 = decide_p & v9ed4f5 | !decide_p & v84563c;
assign v8e79b3 = hgrant1_p & v8e7993 | !hgrant1_p & v84563c;
assign v8ea91c = hbusreq0_p & v8ea919 | !hbusreq0_p & v8ea91b;
assign v9d2676 = hmaster0_p & v9d266f | !hmaster0_p & v84563c;
assign v9998f4 = hbusreq0_p & v9998f3 | !hbusreq0_p & v84563c;
assign v9baf56 = hmaster0_p & v9baf55 | !hmaster0_p & v84563c;
assign v9d26de = busreq_p & v845668 | !busreq_p & v845666;
assign v9965b9 = hmaster1_p & v9965b6 | !hmaster1_p & v99657f;
assign v9854c1 = stateG2_p & v84563c | !stateG2_p & v9854c0;
assign a153b7 = hlock1_p & v84563c | !hlock1_p & v84565c;
assign v9999e8 = hbusreq2 & v9999dc | !hbusreq2 & v9999e7;
assign v9854be = hburst1_p & v9854bd | !hburst1_p & !v84563c;
assign v9baf5a = hburst0 & a153bc | !hburst0 & v9baf59;
assign v8e799d = hmaster0_p & v8e799c | !hmaster0_p & v8e799a;
assign a15500 = hlock1_p & a154ff | !hlock1_p & !v8c20c1;
assign a154f6 = hgrant1_p & v84565c | !hgrant1_p & !a15420;
assign v9baf98 = hbusreq2 & v9baf97 | !hbusreq2 & v84563c;
assign v9998ac = hbusreq0_p & v9998ab | !hbusreq0_p & !v84563c;
assign v9adc04 = hmaster1_p & v9adbff | !hmaster1_p & !v9adc03;
assign v8ea841 = hbusreq2 & v8ea83f | !hbusreq2 & v8ea840;
assign v984ef6 = hbusreq0 & v984eea | !hbusreq0 & v984ef5;
assign v9d27c4 = hgrant2_p & v9d27c2 | !hgrant2_p & v9d27c3;
assign v8c20bf = hlock0_p & v84565c | !hlock0_p & !v8c20be;
assign v9baf18 = hburst1 & v972fac | !hburst1 & v9baf17;
assign v8ea856 = hbusreq0 & v8ea854 | !hbusreq0 & v8ea855;
assign v9d26bf = hgrant2_p & v9d2683 | !hgrant2_p & v9d26be;
assign v9ed46f = hmaster0_p & v9ed469 | !hmaster0_p & !v9ed46e;
assign v8ea843 = hready_p & v8ea80e | !hready_p & v8ea842;
assign a15495 = hready_p & a15494 | !hready_p & a15485;
assign v8ea8c0 = hbusreq0 & v8ea8bb | !hbusreq0 & v8ea8bf;
assign v98561a = hbusreq1_p & v9d2691 | !hbusreq1_p & v84565c;
assign v9855cb = hmaster0_p & v985521 | !hmaster0_p & !v985593;
assign v8ea90e = hmaster0_p & v8ea90b | !hmaster0_p & v8ea82c;
assign v9baf37 = hmaster1_p & v9baf2f | !hmaster1_p & !v9baf36;
assign v99997d = hmaster0_p & v999909 | !hmaster0_p & v9ed487;
assign v9739bf = hready_p & v9739af | !hready_p & !v9739be;
assign v8ea80a = hbusreq1_p & v8ea802 | !hbusreq1_p & v8ea809;
assign v9739de = decide_p & v9739a4 | !decide_p & v9739dd;
assign v985555 = hmastlock_p & v985554 | !hmastlock_p & v84563c;
assign v9999c3 = hburst0 & v9999ba | !hburst0 & v9999c2;
assign v9ed4a6 = locked_p & v9ed4a5 | !locked_p & v84563c;
assign a14da4 = hready_p & a14d5c | !hready_p & a14da2;
assign v984ede = decide_p & v98563f | !decide_p & v984edd;
assign v9d26cf = hready_p & v84564b | !hready_p & !v9d26ce;
assign v9965b3 = hready_p & v9965aa | !hready_p & !v9965b2;
assign v9adc1b = hmaster0_p & v9adbee | !hmaster0_p & v9adbf9;
assign v9baeb3 = hmaster1_p & v9baeb2 | !hmaster1_p & v84563c;
assign v9d26b8 = hgrant0_p & v9d267e | !hgrant0_p & v9d26b7;
assign v985527 = hbusreq1_p & v985526 | !hbusreq1_p & v84563c;
assign v8ea875 = hlock2 & v8ea872 | !hlock2 & v8ea874;
assign v99997b = hbusreq0_p & v999911 | !hbusreq0_p & a14d40;
assign v97399c = hlock0_p & v97399a | !hlock0_p & !v97399b;
assign v984ebc = hbusreq0 & v984eb7 | !hbusreq0 & v984ebb;
assign v9adc5f = hmaster1_p & v9adc5e | !hmaster1_p & v9adc2e;
assign a15430 = decide_p & a1542f | !decide_p & v84565c;
assign v99990b = hmaster0_p & v9baf10 | !hmaster0_p & !v845656;
assign v9a6ac9 = hmaster0_p & v9a6ac8 | !hmaster0_p & v84563c;
assign v9a6a9f = hburst1_p & v9a6a9e | !hburst1_p & v8ea7fa;
assign v9933d6 = hmaster1_p & v9933d5 | !hmaster1_p & !v9933c7;
assign v9adc13 = hmaster0_p & v9adc11 | !hmaster0_p & !v9adc12;
assign v9739db = hmaster1_p & v9739ab | !hmaster1_p & !v9738e8;
assign v878a51 = stateG3_2_p & v84563c | !stateG3_2_p & v861283;
assign v9998e6 = hmaster1_p & v9baf83 | !hmaster1_p & a154a3;
assign v8c117c = decide_p & v8c117b | !decide_p & v8c1155;
assign v984f38 = hlock2_p & v984f20 | !hlock2_p & !v984f37;
assign v8ea8ab = hmaster1_p & v8ea8aa | !hmaster1_p & v8ea7f2;
assign v9739c0 = hgrant2_p & v973998 | !hgrant2_p & !v9739bf;
assign v8e79db = hbusreq2_p & v8e79ca | !hbusreq2_p & v8e79da;
assign v9738d8 = hmaster0_p & v9738d3 | !hmaster0_p & !v9738d7;
assign v9739e5 = hready_p & v9739de | !hready_p & !v9739e4;
assign v985532 = hmaster1_p & v985530 | !hmaster1_p & v985531;
assign v9738cd = hmaster0_p & v9738ca | !hmaster0_p & v9738cc;
assign v9739ff = hmaster0_p & v9739eb | !hmaster0_p & v973899;
assign v8c1134 = stateG2_p & v84563c | !stateG2_p & v8c1130;
assign v8ea8d6 = hgrant0_p & v8ea884 | !hgrant0_p & v8ea82f;
assign v996560 = decide_p & v99655f | !decide_p & v996558;
assign v99991c = hmaster1_p & v99991b | !hmaster1_p & !v9baf32;
assign v9854d1 = hbusreq1_p & v9854d0 | !hbusreq1_p & v84563c;
assign v8e79cc = hbusreq1_p & v8e799a | !hbusreq1_p & v84563c;
assign a14da8 = hbusreq0_p & a14da7 | !hbusreq0_p & !v84563c;
assign a3134f = stateG3_2_p & v84563c | !stateG3_2_p & a3134e;
assign v9ed415 = hmastlock_p & v9ed414 | !hmastlock_p & v84563c;
assign v8c1128 = hlock0_p & v8c1125 | !hlock0_p & v8c1127;
assign v8c113a = locked_p & v8c1136 | !locked_p & v8c1139;
assign v9adc88 = hmaster0_p & v9adc87 | !hmaster0_p & v9adc75;
assign v9adc3d = hmaster0_p & v9adc3a | !hmaster0_p & v9adbee;
assign v9738a8 = hmaster0_p & v9738a7 | !hmaster0_p & v9738a4;
assign v9baf66 = hbusreq1 & v973889 | !hbusreq1 & !v84563c;
assign v9854e0 = hmaster1_p & v9854d2 | !hmaster1_p & v9854df;
assign v985568 = hmastlock_p & v985567 | !hmastlock_p & !v84563c;
assign v9f3576 = hgrant0_p & v845646 | !hgrant0_p & v9f356c;
assign v996593 = hmaster1_p & v9adc38 | !hmaster1_p & !v996592;
assign v985589 = hmaster0_p & v84563c | !hmaster0_p & v985527;
assign v9d26fe = hbusreq0_p & v9d26fd | !hbusreq0_p & v845647;
assign v9854a3 = hmaster0_p & v985491 | !hmaster0_p & v9854a2;
assign v9adc1d = hlock0_p & v9adc19 | !hlock0_p & v9adc1c;
assign v8ea8ee = hbusreq0_p & v8ea8ec | !hbusreq0_p & v8ea8ed;
assign v973887 = stateG2_p & v84563c | !stateG2_p & v86cfb3;
assign v984ebf = hready_p & v984e78 | !hready_p & v984ebe;
assign v8ea85a = decide_p & v8ea7ee | !decide_p & v8ea859;
assign v985524 = hmastlock_p & v985523 | !hmastlock_p & v84563c;
assign v9a6ae2 = hgrant2_p & v9a6ad9 | !hgrant2_p & v9a6ae1;
assign v9baf50 = locked_p & v9baf4f | !locked_p & !v973885;
assign v973a48 = hgrant2_p & v973a2e | !hgrant2_p & !v973a47;
assign v973a02 = hmaster0_p & v9739eb | !hmaster0_p & !v9738c3;
assign v984e5d = hbusreq1_p & v845660 | !hbusreq1_p & !v84563c;
assign v984f39 = hbusreq2 & v84563c | !hbusreq2 & v985645;
assign v9d275e = hmaster0_p & v9d275d | !hmaster0_p & !v84563c;
assign v9ed4f6 = hmaster0_p & v9ed471 | !hmaster0_p & !v84563c;
assign a153e7 = hmaster0_p & v84563c | !hmaster0_p & v845648;
assign v9855cf = decide_p & v9855ca | !decide_p & v9855ce;
assign v9d27b6 = hbusreq0 & v9d27b4 | !hbusreq0 & v9d27b5;
assign v9adca4 = hbusreq0_p & v9adca0 | !hbusreq0_p & !v9adca3;
assign v8e79c9 = hready_p & v8e79be | !hready_p & v8e79c8;
assign v8ea88d = hgrant1_p & v8ea88c | !hgrant1_p & v8ea7e9;
assign v985618 = hready & v985617 | !hready & v84563c;
assign v9855a7 = locked_p & v98554d | !locked_p & v84563c;
assign v9999a2 = hbusreq0 & v9999a1 | !hbusreq0 & v999912;
assign v9baf1d = hmastlock_p & v9baf1c | !hmastlock_p & v84563c;
assign v973910 = hbusreq0_p & v97390e | !hbusreq0_p & v97390f;
assign v996573 = hmaster0_p & v9adc11 | !hmaster0_p & v996572;
assign a153c0 = locked_p & a153bd | !locked_p & !v84563c;
assign v985644 = hmaster1_p & v985641 | !hmaster1_p & v985643;
assign v8c20d0 = decide_p & v845656 | !decide_p & v8c20cf;
assign v8ea8cd = hgrant1_p & v8ea8c9 | !hgrant1_p & v8ea7e9;
assign v9bae86 = hbusreq1_p & v9bae85 | !hbusreq1_p & v84563c;
assign v9999df = hlock0_p & v9999de | !hlock0_p & !v84563c;
assign hmaster1 = v9b40de;
assign v99999c = hgrant2_p & v999984 | !hgrant2_p & !v99999b;
assign v9d2750 = hmaster1_p & v9d271a | !hmaster1_p & !v9d2673;
assign v9ed492 = hmaster1_p & v9ed48d | !hmaster1_p & v9ed489;
assign v984f58 = hmaster0_p & v98561a | !hmaster0_p & !v98556a;
assign v9d2708 = hgrant0_p & v84563c | !hgrant0_p & v9d2707;
assign v9ed483 = hmaster0_p & v9ed471 | !hmaster0_p & !v9ed482;
assign v8e79b0 = hbusreq0_p & v8e79af | !hbusreq0_p & v84563c;
assign v8ea891 = hmaster1_p & v8ea889 | !hmaster1_p & v8ea890;
assign v984ea7 = hbusreq1_p & v984ea5 | !hbusreq1_p & !v984ea6;
assign v985646 = hbusreq0_p & v985644 | !hbusreq0_p & v985645;
assign a2fb4c = hburst0_p & v84563c | !hburst0_p & a2fb4b;
assign v898b4e = hmaster1_p & v84563c | !hmaster1_p & v845652;
assign v9ed49f = hmaster0_p & v84563c | !hmaster0_p & !v9ed49e;
assign v999970 = hbusreq0 & v99996f | !hbusreq0 & v845642;
assign v9855d7 = hmaster0_p & v985557 | !hmaster0_p & v84563c;
assign v9d279e = hgrant0_p & v84563c | !hgrant0_p & v9d2702;
assign v9adc46 = hgrant1_p & v9adc11 | !hgrant1_p & v9adc45;
assign v8ea934 = hbusreq0_p & v8ea932 | !hbusreq0_p & v8ea933;
assign v9855ab = hmastlock_p & v9855aa | !hmastlock_p & !v84563c;
assign v9adc31 = hmaster1_p & v9adc28 | !hmaster1_p & v9adc30;
assign v9adbf6 = hmaster1_p & v9adbf0 | !hmaster1_p & v9adbf5;
assign v8c112b = hmaster1_p & v8c112a | !hmaster1_p & v8c1124;
assign v9baf88 = stateG10_1_p & v9ed4ac | !stateG10_1_p & v9baf87;
assign v973901 = hbusreq0_p & v9738ff | !hbusreq0_p & v973900;
assign v9a6acb = stateG10_1_p & v84563c | !stateG10_1_p & v9a6aca;
assign v973a46 = decide_p & v973a2a | !decide_p & v973a45;
assign v8c20e1 = hbusreq2_p & v8c20d2 | !hbusreq2_p & !v8c20e0;
assign v984e5b = hmaster0_p & v984e5a | !hmaster0_p & v84563c;
assign v984f7a = hmaster0_p & v984eac | !hmaster0_p & v984ea7;
assign v99998a = hgrant0_p & v999985 | !hgrant0_p & !v999989;
assign v984f90 = hready_p & v84563c | !hready_p & v984f8f;
assign v9855d8 = hmaster1_p & v9855d7 | !hmaster1_p & v84563c;
assign v984e68 = hbusreq1_p & v9d2691 | !hbusreq1_p & !v984e67;
assign v8ea822 = hbusreq1_p & v8ea820 | !hbusreq1_p & !v8ea821;
assign v9adc0b = hmaster1_p & v9adc09 | !hmaster1_p & !v9adc05;
assign v973935 = hready_p & v97392a | !hready_p & !v973934;
assign v9a6ac2 = hbusreq1_p & v9a6abb | !hbusreq1_p & v9a6ac1;
assign v9854b8 = hmaster0_p & v84563c | !hmaster0_p & v845641;
assign v9d2703 = hbusreq0_p & v9d2702 | !hbusreq0_p & v845647;
assign v996589 = hmaster0_p & v996586 | !hmaster0_p & !v996552;
assign v9ed4f1 = hbusreq2_p & v9ed4ca | !hbusreq2_p & v9ed4f0;
assign v984f5d = hgrant1_p & v98556a | !hgrant1_p & v84563c;
assign v9965bf = hbusreq0_p & v9965bc | !hbusreq0_p & v9965be;
assign v9d278e = hbusreq2 & v9d278d | !hbusreq2 & v9d2680;
assign v985509 = hmaster0_p & v9854cf | !hmaster0_p & v845641;
assign v985500 = hbusreq1_p & v9854ff | !hbusreq1_p & v84563c;
assign v8e79a4 = hmaster1_p & v8e79a3 | !hmaster1_p & v8e799d;
assign v8ea92f = decide_p & v8ea7ee | !decide_p & v8ea92e;
assign v973908 = hmaster1_p & v973907 | !hmaster1_p & v9738a8;
assign v973960 = hgrant0_p & v97395b | !hgrant0_p & v97395f;
assign v9ed4fe = hmaster0_p & v9ed4fd | !hmaster0_p & v9ed4b4;
assign v9739ac = hmaster1_p & v9739ab | !hmaster1_p & !v973967;
assign v8c116e = stateG3_0_p & v84563c | !stateG3_0_p & !v845658;
assign v985626 = hlock1_p & v9854d0 | !hlock1_p & v845641;
assign v9a6aca = hgrant1_p & v9a6ab1 | !hgrant1_p & v84563c;
assign v9d26e8 = hmaster1_p & v84563c | !hmaster1_p & v9d2673;
assign v9ed52e = hready_p & v84563c | !hready_p & v9ed52d;
assign v9ed45b = hburst1 & v9ed45a | !hburst1 & !v84563c;
assign v8ea839 = hbusreq1_p & v8ea7e9 | !hbusreq1_p & v8ea818;
assign v9d2693 = hgrant1_p & v845647 | !hgrant1_p & v9d2692;
assign v9d26db = hready_p & v9d26d9 | !hready_p & !v9d26da;
assign a14d6d = hready_p & a14d5d | !hready_p & !a14d68;
assign v8e79d3 = hmaster0_p & v8e79d2 | !hmaster0_p & v84563c;
assign v9998a3 = decide_p & v9998a2 | !decide_p & v84563c;
assign v999929 = hmastlock_p & v9ed44b | !hmastlock_p & v84563c;
assign v9d2794 = decide_p & v9d2792 | !decide_p & v9d2793;
assign v9bae7c = stateG2_p & v84563c | !stateG2_p & v9bae7b;
assign v9ed430 = stateG2_p & v84563c | !stateG2_p & v9ed42f;
assign v9d277f = stateG10_1_p & v845641 | !stateG10_1_p & !v9d277e;
assign v9d266a = stateG2_p & v84563c | !stateG2_p & !v9d2669;
assign v984e6f = hready & v984e6e | !hready & v985569;
assign v861283 = stateG3_0_p & v84563c | !stateG3_0_p & v8901af;
assign v8ea810 = stateG2_p & v84563c | !stateG2_p & !v8ea80f;
assign a14d6f = hgrant0_p & v845642 | !hgrant0_p & a14d6e;
assign v8ea883 = hmaster1_p & v8ea880 | !hmaster1_p & v8ea882;
assign v9baf26 = hbusreq2 & v9baf25 | !hbusreq2 & !v85bb54;
assign v9854a9 = hbusreq0_p & v9854a6 | !hbusreq0_p & v9854a8;
assign v8ea871 = hbusreq0_p & v8ea864 | !hbusreq0_p & v8ea870;
assign v985624 = hready & v985623 | !hready & !v84563c;
assign v9ed471 = hbusreq1_p & v9ed470 | !hbusreq1_p & !v84563c;
assign v9999bd = hburst1 & v9999ba | !hburst1 & v9999bc;
assign v9a6a94 = stateG3_0_p & v84563c | !stateG3_0_p & !v84566c;
assign v8ea8d0 = hmaster0_p & v8ea8cf | !hmaster0_p & v8ea822;
assign v9a6ab9 = hgrant1_p & v84563c | !hgrant1_p & v9a6a98;
assign v9adcd0 = hmaster1_p & v9adcce | !hmaster1_p & !v9adc7c;
assign v97390e = hmaster1_p & v97390d | !hmaster1_p & !v973890;
assign v98550c = hlock0_p & v98550a | !hlock0_p & v98550b;
assign v9adcb9 = hbusreq1_p & v9adca9 | !hbusreq1_p & !v9adcb8;
assign v985550 = stateA1_p & v985544 | !stateA1_p & !v98549a;
assign v98552e = decide_p & v98551f | !decide_p & v98552d;
assign v973947 = hmaster1_p & v9738a5 | !hmaster1_p & v973946;
assign v999925 = hmaster1_p & v999924 | !hmaster1_p & !v9baf32;
assign v9855a5 = hgrant0_p & v9855a4 | !hgrant0_p & v98559c;
assign v9854fc = hready & v8ea7e5 | !hready & !v972fac;
assign v9adc9f = hmaster1_p & v9adc9d | !hmaster1_p & v9adc9e;
assign v985592 = hready & v98558d | !hready & v985591;
assign v97395f = hbusreq0_p & v9738d5 | !hbusreq0_p & v97395e;
assign v9998af = decide_p & v9998ae | !decide_p & v84565e;
assign v984e72 = hbusreq1_p & v984e6a | !hbusreq1_p & !v984e71;
assign v8ea84d = hmaster1_p & v8ea84b | !hmaster1_p & v8ea7f4;
assign v9adc9d = hmaster0_p & v9adc76 | !hmaster0_p & v84563c;
assign v985504 = hmaster1_p & v985501 | !hmaster1_p & v9854df;
assign v984ec8 = hbusreq0_p & v984ec7 | !hbusreq0_p & v985645;
assign v984f80 = hbusreq0_p & v984f7f | !hbusreq0_p & v984f74;
assign v9d26a8 = stateA1_p & v84563c | !stateA1_p & !v8c1130;
assign v9ed4c3 = hgrant0_p & v9ed4c2 | !hgrant0_p & !v9ed4b6;
assign v9738a4 = hmastlock_p & v973887 | !hmastlock_p & v845666;
assign v97390b = hmaster1_p & v973907 | !hmaster1_p & v9738ad;
assign v9739d3 = decide_p & v973988 | !decide_p & !v9739d2;
assign v8e79c2 = hgrant1_p & v8e79a9 | !hgrant1_p & v84563c;
assign v99659e = hmaster1_p & v9adc49 | !hmaster1_p & v99659d;
assign v9adcdd = locked_p & v845668 | !locked_p & v9adc75;
assign v9ed452 = hlock2_p & v9ed43a | !hlock2_p & v9ed451;
assign v999940 = decide_p & v99993f | !decide_p & v84565e;
assign v999988 = hlock0_p & v999987 | !hlock0_p & v99993a;
assign v9ed48f = hmaster1_p & v9ed48d | !hmaster1_p & v9ed478;
assign v9738df = hbusreq0_p & v9738bf | !hbusreq0_p & v9738de;
assign v8ea802 = hgrant1_p & v8ea7e6 | !hgrant1_p & v84563c;
assign v99656f = hmaster1_p & v9adc09 | !hmaster1_p & v996569;
assign v9d27bc = hgrant0_p & v84563c | !hgrant0_p & !v9d27ba;
assign v9adc87 = hbusreq1_p & v9adc85 | !hbusreq1_p & !v9adc86;
assign v9999a3 = decide_p & v9999a2 | !decide_p & v84563c;
assign v8c1155 = hgrant0_p & v8c114f | !hgrant0_p & v8c1154;
assign v9d2681 = hbusreq2 & v9d267d | !hbusreq2 & v9d2680;
assign v984f57 = hmaster1_p & a154a3 | !hmaster1_p & v984f56;
assign v984ead = hmaster0_p & v984eac | !hmaster0_p & v84563c;
assign v8c20d3 = decide_p & v8c20b7 | !decide_p & !v84565c;
assign v973902 = hmaster0_p & v973886 | !hmaster0_p & v9738dc;
assign v8c114c = locked_p & v8c114b | !locked_p & v84563c;
assign v8ea87f = hready_p & v8ea7e8 | !hready_p & v8ea87e;
assign v9baf40 = decide_p & v9baf3f | !decide_p & v84563c;
assign v9855b5 = hmaster0_p & v84563c | !hmaster0_p & v9855b4;
assign v9adcf4 = hgrant2_p & v9adcd4 | !hgrant2_p & !v9adcf3;
assign v9739bb = hmaster1_p & v9739ba | !hmaster1_p & v973967;
assign v845652 = hmaster0_p & v84563c | !hmaster0_p & !v84563c;
assign v973a16 = hgrant0_p & v973a12 | !hgrant0_p & v973a15;
assign v8c115b = hgrant1_p & v8c113a | !hgrant1_p & v8c1120;
assign v98561f = decide_p & v985611 | !decide_p & v98561e;
assign v973957 = decide_p & v973953 | !decide_p & v973956;
assign v973a3d = hmaster1_p & v9739a9 | !hmaster1_p & !v973a13;
assign v9a6ad0 = decide_p & v9a6ab0 | !decide_p & v9a6acf;
assign v973996 = hbusreq0_p & v973994 | !hbusreq0_p & v973995;
assign v8c114b = hmastlock_p & v8768ab | !hmastlock_p & v84563c;
assign v984f74 = hmaster1_p & v984f70 | !hmaster1_p & v984f73;
assign v9854dc = hbusreq1_p & v9854db | !hbusreq1_p & v84563c;
assign v984e58 = hgrant1_p & v985498 | !hgrant1_p & v84563c;
assign v9d275c = stateG10_1_p & v9d2691 | !stateG10_1_p & !v9d275b;
assign v9ed443 = hmaster0_p & v84563c | !hmaster0_p & v9ed442;
assign v9854ae = hlock1_p & v9854ab | !hlock1_p & v9854ad;
assign v9adc0c = hlock0_p & v9adc0a | !hlock0_p & v9adc0b;
assign v9adc83 = hlock2_p & v9adc7e | !hlock2_p & !v9adc82;
assign v8ea80e = decide_p & v8ea808 | !decide_p & v8ea80d;
assign v9854f4 = stateA1_p & v84563c | !stateA1_p & !v9854f3;
assign v9ed468 = hlock1_p & v9ed45d | !hlock1_p & v9ed467;
assign v9baf57 = stateA1_p & a153bb | !stateA1_p & !v9ed42e;
assign v9ed47d = stateA1_p & v972fac | !stateA1_p & !v9ed47c;
assign v8c1165 = decide_p & v84563c | !decide_p & v8c1164;
assign v9ed482 = hbusreq1_p & v9ed481 | !hbusreq1_p & v84563c;
assign v973a1c = hbusreq0_p & v97397e | !hbusreq0_p & v973a1b;
assign v9baeca = hlock2_p & v9baec9 | !hlock2_p & v84563c;
assign a153d4 = hmaster0_p & a153cf | !hmaster0_p & a153d3;
assign v9ed461 = stateG2_p & v84563c | !stateG2_p & v9ed460;
assign v9933c5 = hlock1_p & v9933c4 | !hlock1_p & v8c20d7;
assign v984edb = hbusreq0 & v984eda | !hbusreq0 & v985645;
assign v9baf89 = hbusreq1_p & v9baf86 | !hbusreq1_p & !v9baf88;
assign v9d275f = hmaster1_p & v9d275e | !hmaster1_p & !v9d2671;
assign v9adcce = hmaster0_p & v9adc75 | !hmaster0_p & v9adca1;
assign v9ed43d = hburst1 & v86cfb3 | !hburst1 & v84563c;
assign v8e79b4 = hlock1_p & v8e79b3 | !hlock1_p & v84563c;
assign v9854ec = stateG2_p & v84563c | !stateG2_p & v9854eb;
assign v8e79d0 = decide_p & v8e79cf | !decide_p & v8e79ab;
assign v9bafa0 = jx0_p & v9baefd | !jx0_p & v9baf9f;
assign v9adcf6 = jx2_p & v84563c | !jx2_p & !v9adcf5;
assign v9adc29 = hgrant1_p & v9adbef | !hgrant1_p & v9adbee;
assign a14dbf = hbusreq2_p & a14dbe | !hbusreq2_p & !a14d72;
assign v9a6ae1 = hready_p & v9a6adf | !hready_p & v9a6ae0;
assign v9d2686 = hmastlock_p & v9d2685 | !hmastlock_p & !v84563c;
assign v9933c0 = hgrant1_p & v84563c | !hgrant1_p & !v9933b7;
assign v985523 = stateG2_p & v84563c | !stateG2_p & !v985522;
assign v8ea82a = hgrant1_p & v8ea7f0 | !hgrant1_p & v8ea7e9;
assign v9baead = hmaster0_p & v84563c | !hmaster0_p & !a153d1;
assign v973a28 = decide_p & v973a25 | !decide_p & !v973a27;
assign v8ea8ba = hbusreq0_p & v8ea8b9 | !hbusreq0_p & v8ea869;
assign v9d2793 = hbusreq2 & v9d2751 | !hbusreq2 & v9d2680;
assign v9739f9 = hlock2_p & v9739f6 | !hlock2_p & v9739f8;
assign v973905 = hbusreq0_p & v973903 | !hbusreq0_p & v973904;
assign v9738c9 = hgrant1_p & v973886 | !hgrant1_p & !v973885;
assign v8ea801 = hmaster0_p & v8ea800 | !hmaster0_p & v84563c;
assign v984e57 = hmaster0_p & v984e54 | !hmaster0_p & v984e56;
assign v985520 = hready & v84565c | !hready & !v84563c;
assign v984f87 = hbusreq0 & v985645 | !hbusreq0 & v984ebb;
assign v985641 = hmaster0_p & v985520 | !hmaster0_p & v985526;
assign v9739f2 = decide_p & v9739f1 | !decide_p & v9739ea;
assign v9999ed = hgrant2_p & v9999d8 | !hgrant2_p & !v9999ec;
assign v9a6aa9 = hlock0_p & v9a6aa6 | !hlock0_p & v9a6aa8;
assign v9ed479 = hmaster1_p & v9ed46f | !hmaster1_p & v9ed478;
assign v9adc72 = hbusreq2_p & v9adc52 | !hbusreq2_p & v9adc71;
assign v9d26f9 = stateG10_1_p & v84563c | !stateG10_1_p & v9d2694;
assign v9855b1 = hmaster0_p & v9855b0 | !hmaster0_p & v985582;
assign v9999d4 = hbusreq0 & v9999b9 | !hbusreq0 & v9999d3;
assign v9d2746 = decide_p & v9d2733 | !decide_p & v9d272c;
assign v9baf2c = busreq_p & v9baf2a | !busreq_p & v9baf2b;
assign a14da0 = hbusreq0_p & a14d9f | !hbusreq0_p & a14d8e;
assign v9998a4 = hready_p & v84563c | !hready_p & v9998a3;
assign v9a6abd = hbusreq1_p & v9a6abc | !hbusreq1_p & v84563c;
assign v9ed4b8 = hmaster0_p & v84563c | !hmaster0_p & v9ed436;
assign v9854cb = hbusreq0_p & v9854c9 | !hbusreq0_p & v9854ca;
assign v9ed463 = stateG2_p & v84563c | !stateG2_p & !a2bd3d;
assign v8ea90b = hbusreq1_p & v8ea7e9 | !hbusreq1_p & !v8ea90a;
assign v97393d = hbusreq0_p & v97389d | !hbusreq0_p & v97393c;
assign v9854c2 = hmastlock_p & v9854c1 | !hmastlock_p & v84563c;
assign a15431 = hready_p & a15430 | !hready_p & a1540c;
assign v8ea860 = hbusreq0_p & v8ea807 | !hbusreq0_p & v8ea85f;
assign v8c1149 = hmaster1_p & v8c1144 | !hmaster1_p & !v8c1148;
assign v9adc32 = hbusreq0_p & v9adc2f | !hbusreq0_p & v9adc31;
assign v86292d = hmaster0_p & v84563c | !hmaster0_p & !v845646;
assign v9738f4 = hmaster1_p & v9738f2 | !hmaster1_p & !v9738dd;
assign v9ed48e = hmaster1_p & v9ed48d | !hmaster1_p & v9ed472;
assign v8c20b6 = hmaster0_p & v84563c | !hmaster0_p & !v84565c;
assign v985574 = locked_p & v985573 | !locked_p & v84563c;
assign v9d27af = hbusreq0 & v9d27ac | !hbusreq0 & v9d27ae;
assign v9d273a = hgrant0_p & v84563c | !hgrant0_p & v9d2739;
assign v9baeef = hready_p & v84563c | !hready_p & v9baeee;
assign v9adc58 = decide_p & v9adc57 | !decide_p & v9adc14;
assign v984e6e = locked_p & v984e6d | !locked_p & v84563c;
assign v98555c = hbusreq0 & v98553e | !hbusreq0 & v98555b;
assign v9baf1b = hburst1 & v972fac | !hburst1 & a2f895;
assign v9d26ed = hmaster0_p & v9d266d | !hmaster0_p & v84563c;
assign v8c20c9 = hmaster0_p & v8c20ba | !hmaster0_p & !v845656;
assign v9d26a1 = hgrant0_p & v84563c | !hgrant0_p & !v9d269f;
assign v9738e6 = stateG10_1_p & v97388d | !stateG10_1_p & v9738e5;
assign v8ea939 = hbusreq2_p & v8ea931 | !hbusreq2_p & v8ea938;
assign v996563 = hbusreq1_p & v996561 | !hbusreq1_p & !v996562;
assign v8ea81b = hbusreq1 & v8ea819 | !hbusreq1 & v8ea81a;
assign v984ecc = hmaster0_p & v984e66 | !hmaster0_p & v984eb3;
assign v8c111e = decide_p & v8c111d | !decide_p & v8c111c;
assign jx1 = v9965d3;
assign v97392e = hbusreq0_p & v97392c | !hbusreq0_p & v97392d;
assign v9ed4e9 = hmaster1_p & v9ed4e8 | !hmaster1_p & v9ed49f;
assign a14d3c = hready_p & a15517 | !hready_p & a154f3;
assign v984f7b = hmaster1_p & v984f76 | !hmaster1_p & v984f7a;
assign v9965a9 = hbusreq0_p & v9965a7 | !hbusreq0_p & v9965a8;
assign v8e79bd = hgrant0_p & v8e79ae | !hgrant0_p & v8e79bc;
assign v9adc2b = hlock1_p & v9adc29 | !hlock1_p & v9adc2a;
assign v97389a = hmaster0_p & v973885 | !hmaster0_p & v973899;
assign v984ef3 = hmaster1_p & v984ee3 | !hmaster1_p & v984ef2;
assign v973988 = hbusreq0_p & v973986 | !hbusreq0_p & v973987;
assign v9d279f = hgrant0_p & v84563c | !hgrant0_p & !v9d2702;
assign v973a07 = hbusreq1_p & v9738d0 | !hbusreq1_p & !v973a06;
assign v9d2784 = hgrant0_p & v84563c | !hgrant0_p & v9d2783;
assign v9adc7e = hbusreq0_p & v9adc7b | !hbusreq0_p & v9adc7d;
assign v9855c5 = decide_p & v9855c0 | !decide_p & v9855c4;
assign v9d2727 = hmaster0_p & v9d271e | !hmaster0_p & v84563c;
assign v973a12 = hbusreq0_p & v9739fe | !hbusreq0_p & v973a11;
assign v9ed4a2 = stateG2_p & v84563c | !stateG2_p & !v9ed411;
assign v9739df = hmaster1_p & v9739b5 | !hmaster1_p & !v9738be;
assign v9adc93 = hmaster0_p & v9adc75 | !hmaster0_p & v9adc77;
assign v9738d3 = hbusreq1_p & v9738d0 | !hbusreq1_p & !v9738d2;
assign v99996b = hgrant2_p & v999932 | !hgrant2_p & !v99996a;
assign v9baf9b = decide_p & v9baf3f | !decide_p & !v84563c;
assign v9739fb = hbusreq0_p & v973954 | !hbusreq0_p & v9739fa;
assign v99655e = hbusreq0_p & v99655b | !hbusreq0_p & v99655d;
assign v8ea844 = hgrant2_p & v8ea7f8 | !hgrant2_p & v8ea843;
assign v9855fb = hmaster0_p & v98548f | !hmaster0_p & v84563c;
assign v9ed4ac = locked_p & v9ed4ab | !locked_p & v84563c;
assign v8e7998 = stateG3_2_p & v84563c | !stateG3_2_p & !v84566c;
assign v8ea916 = hlock0 & v8ea911 | !hlock0 & v8ea915;
assign v9965a7 = hmaster1_p & v9965a6 | !hmaster1_p & v99655a;
assign v973962 = stateG10_1_p & v97388d | !stateG10_1_p & v973961;
assign v9739b3 = hmaster0_p & v973885 | !hmaster0_p & !v973894;
assign v9854d0 = hready & v8ea7e5 | !hready & a153d1;
assign v9998df = decide_p & v9998d6 | !decide_p & !v84565e;
assign v973917 = hmaster1_p & v973907 | !hmaster1_p & v9738c6;
assign a154d2 = hmaster0_p & a154d1 | !hmaster0_p & !a153d1;
assign v9739a4 = hgrant0_p & v97399e | !hgrant0_p & v9739a3;
assign v9d274d = hmaster1_p & v845652 | !hmaster1_p & v9d2673;
assign v9ed4db = hmaster0_p & v9ed469 | !hmaster0_p & v9ed488;
assign v9adc69 = hmaster0_p & v9adc35 | !hmaster0_p & v9adbee;
assign v9d267d = hbusreq0 & v9d267b | !hbusreq0 & v9d267c;
assign v9965c3 = hmaster1_p & v9965c1 | !hmaster1_p & !v996592;
assign v9d268d = hbusreq1 & v9d268c | !hbusreq1 & v84563c;
assign v84565c = locked_p & v84563c | !locked_p & !v84563c;
assign v98552d = hbusreq0_p & v985529 | !hbusreq0_p & v98552c;
assign v9ed46b = hburst1 & v9ed46a | !hburst1 & v84563c;
assign v973a2b = hmaster1_p & v97390d | !hmaster1_p & !v9739e8;
assign v9999c7 = hmaster0_p & v84563c | !hmaster0_p & v9999c6;
assign v9adbfe = hmastlock_p & v8ec3e4 | !hmastlock_p & v84563c;
assign v845647 = hbusreq1 & v84563c | !hbusreq1 & !v84563c;
assign v9738b1 = hmaster1_p & v9738b0 | !hmaster1_p & v9738a8;
assign v984ed1 = decide_p & v984e65 | !decide_p & v984ed0;
assign v8ea812 = hmastlock_p & v8ea811 | !hmastlock_p & v84563c;
assign v9738ed = hmaster0_p & v9738e7 | !hmaster0_p & !v9738ec;
assign v984f61 = hmaster1_p & v984f5b | !hmaster1_p & v984f60;
assign v984f2b = hmaster0_p & v98562c | !hmaster0_p & !v9854da;
assign v99657e = locked_p & v9adc60 | !locked_p & !v9adbee;
assign v9ed448 = hmaster1_p & v9ed441 | !hmaster1_p & v9ed447;
assign v866c94 = hburst0_p & v84563c | !hburst0_p & v845650;
assign v98549d = hmastlock_p & v98549c | !hmastlock_p & v84563c;
assign v8e79a7 = hbusreq0_p & v8e79a6 | !hbusreq0_p & v8e79a5;
assign v973a0f = hgrant0_p & v973a04 | !hgrant0_p & v973a0e;
assign v98559f = locked_p & v98559e | !locked_p & v84563c;
assign v8c20cc = stateG10_1_p & v845656 | !stateG10_1_p & !v8c20cb;
assign v985604 = hready & v985497 | !hready & !v985603;
assign v9adbef = locked_p & v9adbed | !locked_p & v9adbee;
assign v9ed451 = hbusreq2 & v9ed449 | !hbusreq2 & !v9ed450;
assign v9d26ca = hmaster1_p & v9d26c7 | !hmaster1_p & !v9d2673;
assign v9baf15 = hbusreq0_p & v9baf12 | !hbusreq0_p & v9baf14;
assign v98554d = hmastlock_p & v98554c | !hmastlock_p & !v84563c;
assign v9adcd5 = hmaster0_p & v9adc76 | !hmaster0_p & !v9adc75;
assign v97389c = hmaster0_p & v97389b | !hmaster0_p & v973889;
assign v9adca1 = locked_p & v845668 | !locked_p & !v84563c;
assign a14dc0 = jx2_p & a14dbf | !jx2_p & a14d85;
assign v984f77 = hmaster0_p & v984eac | !hmaster0_p & v984e66;
assign v9854f8 = busreq_p & v84563c | !busreq_p & v9854f7;
assign v9855d0 = hready_p & v9855c5 | !hready_p & v9855cf;
assign v985570 = stateA1_p & v985544 | !stateA1_p & v9854bf;
assign v9a6ab2 = hmaster0_p & v84563c | !hmaster0_p & v9a6ab1;
assign v973927 = hmaster1_p & v973925 | !hmaster1_p & !v9738ed;
assign v8ea8c4 = hready_p & v8ea862 | !hready_p & v8ea8c3;
assign v984f63 = hmaster1_p & v984f5b | !hmaster1_p & v984f62;
assign v9738ba = hbusreq0_p & v9738b8 | !hbusreq0_p & v9738b9;
assign v9baeb0 = hmaster1_p & v9baeaf | !hmaster1_p & v84563c;
assign v9ed4cd = hmaster1_p & v9ed4cb | !hmaster1_p & v9ed447;
assign v9baf76 = hgrant0_p & v9baf49 | !hgrant0_p & v9baf75;
assign v984f27 = hmaster1_p & v84563c | !hmaster1_p & !v984f26;
assign v97394e = hmaster1_p & v9738b0 | !hmaster1_p & v973946;
assign v9d269c = hbusreq0 & v9d269a | !hbusreq0 & !v9d269b;
assign v9adbf1 = locked_p & v8ea7ea | !locked_p & v9adbee;
assign v9d277e = hgrant1_p & v845647 | !hgrant1_p & !v845641;
assign v9738c6 = hmaster0_p & v97389b | !hmaster0_p & !v9738c5;
assign v8ea8a5 = hmaster1_p & v8ea8a4 | !hmaster1_p & v8ea7f4;
assign v9bae8e = hbusreq1_p & a153d1 | !hbusreq1_p & v845656;
assign a14d5c = decide_p & v84563c | !decide_p & v84565c;
assign v984e64 = hgrant0_p & v84563c | !hgrant0_p & v984e63;
assign v8c1144 = hmaster0_p & v8c1143 | !hmaster0_p & v84563c;
assign v984e77 = hbusreq0 & v984e76 | !hbusreq0 & v84563c;
assign v9adc2e = hmaster0_p & v9adc2d | !hmaster0_p & v9adc27;
assign v8ea827 = hbusreq1_p & v8ea7e9 | !hbusreq1_p & !v8ea826;
assign v98560e = hbusreq2 & v985602 | !hbusreq2 & v98560d;
assign v9baf8a = hmaster0_p & v9baf89 | !hmaster0_p & v84563c;
assign v9d2788 = decide_p & v9d277b | !decide_p & !v9d276a;
assign v973a03 = hmaster1_p & v9738b0 | !hmaster1_p & v973a02;
assign v8e79d9 = hready_p & v8e79d7 | !hready_p & v8e79d8;
assign v9933cb = hbusreq1_p & v9933c4 | !hbusreq1_p & !v9933ca;
assign v9ed4ca = hgrant2_p & v9ed497 | !hgrant2_p & v9ed4c9;
assign v9ed49a = hmaster1_p & v9ed498 | !hmaster1_p & v9ed499;
assign v9d27a6 = hbusreq0 & v9d27a4 | !hbusreq0 & !v9d27a5;
assign v9933db = hgrant2_p & v9933d3 | !hgrant2_p & v9933da;
assign a153cb = hburst0_p & v863b4b | !hburst0_p & a153ca;
assign v8ea89b = hlock0 & v8ea89a | !hlock0 & v8ea893;
assign v9999b6 = hbusreq2_p & v9999aa | !hbusreq2_p & v9999b5;
assign v984ec4 = hbusreq0 & v984ec3 | !hbusreq0 & v84563c;
assign v9a6adc = hmaster1_p & v9a6adb | !hmaster1_p & v9a6abe;
assign v8e7989 = stateG3_2_p & v84563c | !stateG3_2_p & v8e7988;
assign v973944 = stateG10_1_p & v97388d | !stateG10_1_p & v973893;
assign v9999a6 = hbusreq0 & v9999a5 | !hbusreq0 & v99993e;
assign v99999e = jx0_p & v9998e2 | !jx0_p & v99999d;
assign v99989c = hmaster1_p & v84563c | !hmaster1_p & v9bae8f;
assign v9855e3 = hbusreq0_p & v9855e1 | !hbusreq0_p & v9855e2;
assign v9baea3 = hbusreq0_p & v9baea2 | !hbusreq0_p & v84565c;
assign v8ea82f = hbusreq0_p & v8ea829 | !hbusreq0_p & v8ea82e;
assign a154f2 = hlock2_p & a154ed | !hlock2_p & a154f1;
assign v9adc5d = hbusreq0_p & v9adc5c | !hbusreq0_p & v9adc1c;
assign v9738a5 = hmaster0_p & v973885 | !hmaster0_p & v9738a4;
assign v9855f3 = hgrant0_p & v9855ec | !hgrant0_p & v9855f2;
assign v9ed4d9 = hbusreq0_p & v9ed4d7 | !hbusreq0_p & v9ed4d8;
assign a14d68 = decide_p & a14d67 | !decide_p & v84565c;
assign v985614 = stateA1_p & v84563c | !stateA1_p & !v985613;
assign v98560c = hbusreq0_p & v98560b | !hbusreq0_p & v84563c;
assign v9855a0 = hready & v98559f | !hready & !v84563c;
assign v9854d5 = hmaster1_p & v9854d2 | !hmaster1_p & v9854b8;
assign v9baefd = hbusreq2_p & v9baefc | !hbusreq2_p & !v9baea0;
assign v99998e = decide_p & v99998d | !decide_p & v84565e;
assign v9ed501 = hgrant0_p & v84563c | !hgrant0_p & !v9ed500;
assign v98553e = hgrant0_p & v985534 | !hgrant0_p & v98553d;
assign v9bae89 = hbusreq2 & v9bae7a | !hbusreq2 & v9bae88;
assign v9adcb8 = stateG10_1_p & v84563c | !stateG10_1_p & !v9adcb7;
assign v9739c5 = hbusreq0_p & v9738b3 | !hbusreq0_p & v973951;
assign v9adc43 = hmaster0_p & v8ea7ef | !hmaster0_p & !v9adc12;
assign v9d26d2 = hbusreq1_p & v9d268f | !hbusreq1_p & !v9d26d1;
assign v9d26d7 = hgrant0_p & v84563c | !hgrant0_p & !v9d26d5;
assign v985506 = hbusreq0_p & v985505 | !hbusreq0_p & v985504;
assign v9933bc = hready_p & v9933bb | !hready_p & !v84563c;
assign v9adcc4 = hgrant1_p & v9adc94 | !hgrant1_p & !v9adc75;
assign v9d27a7 = hbusreq2 & v9d27a6 | !hbusreq2 & v9d279c;
assign v8ea911 = hgrant0_p & v8ea905 | !hgrant0_p & v8ea910;
assign v9855ae = hgrant1_p & v845641 | !hgrant1_p & v84563c;
assign v8ea7ee = hmaster1_p & v8ea7e9 | !hmaster1_p & v8ea7ed;
assign v996552 = hmastlock_p & v996551 | !hmastlock_p & !v84563c;
assign v98558c = hmastlock_p & v98558b | !hmastlock_p & !v84563c;
assign v8ea896 = hbusreq1_p & v8ea7e9 | !hbusreq1_p & v8ea895;
assign v8e7991 = stateG2_p & v84563c | !stateG2_p & v8e7990;
assign v996558 = hbusreq0_p & v996555 | !hbusreq0_p & v996557;
assign v9adc9a = hbusreq0_p & v9adc97 | !hbusreq0_p & v9adc99;
assign v9d2667 = hready & v9d2666 | !hready & !v84563c;
assign a1548c = hmaster0_p & a15488 | !hmaster0_p & a15489;
assign v996583 = hlock1_p & v996582 | !hlock1_p & !v9adc2a;
assign v999930 = hlock2_p & v999920 | !hlock2_p & v99992f;
assign v9baf00 = stateG2_p & v86cfb3 | !stateG2_p & !v84563c;
assign v985595 = hmaster1_p & v985588 | !hmaster1_p & v985594;
assign v9adc0f = busreq_p & v9adbe7 | !busreq_p & v8ecba9;
assign v9d2763 = hbusreq0 & v9d2760 | !hbusreq0 & v9d2762;
assign v8c20c0 = hbusreq0_p & v8c20bf | !hbusreq0_p & !v8c20be;
assign v984f54 = hbusreq2 & v984f53 | !hbusreq2 & v84563c;
assign v984f7e = hmaster0_p & v985642 | !hmaster0_p & !v9855a0;
assign v999976 = decide_p & v999975 | !decide_p & v84563c;
assign v9bae82 = locked_p & v9bae81 | !locked_p & v84563c;
assign v9855c9 = hbusreq0 & v985517 | !hbusreq0 & v9855c8;
assign v9a6ad2 = hgrant2_p & v9a6ab5 | !hgrant2_p & v9a6ad1;
assign v9d2772 = hmaster1_p & v9d276f | !hmaster1_p & v9d2673;
assign a1541d = hburst0_p & v8e7989 | !hburst0_p & a15417;
assign v8ea7e5 = hmastlock_p & v8ea7e4 | !hmastlock_p & v84563c;
assign v9965ac = hmaster1_p & v9965ab | !hmaster1_p & v996564;
assign v9ed496 = decide_p & v9ed495 | !decide_p & !v84563c;
assign v98557e = hmaster0_p & v98557b | !hmaster0_p & v98557d;
assign v9baefa = decide_p & v9baef7 | !decide_p & v84563c;
assign v8c111d = hlock2_p & v8c111c | !hlock2_p & v84563c;
assign v8ea834 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea833;
assign v99990f = hlock0_p & v99990c | !hlock0_p & v99990e;
assign v9998ff = hbusreq2 & v9998fb | !hbusreq2 & !v9998fe;
assign v9a6ac5 = hgrant0_p & v9a6ab6 | !hgrant0_p & v9a6ac4;
assign v9999ec = hready_p & v9999ea | !hready_p & !v9999eb;
assign v9adca8 = hmaster0_p & v9adca7 | !hmaster0_p & v84563c;
assign v985584 = hmaster1_p & v98557e | !hmaster1_p & v985583;
assign v8ea8c6 = hbusreq2_p & v8ea8a1 | !hbusreq2_p & v8ea8c5;
assign v9adc09 = hmaster0_p & v9adbfe | !hmaster0_p & !v8ea7ea;
assign v9d271b = hmaster1_p & v9d271a | !hmaster1_p & !v9d2671;
assign a15408 = hmaster1_p & a153eb | !hmaster1_p & a153e7;
assign v99990e = hmaster1_p & v99990d | !hmaster1_p & !v9baf32;
assign v9d2723 = hbusreq0 & v9d2722 | !hbusreq0 & v9d267c;
assign v9a6ace = hmaster1_p & v9a6ac9 | !hmaster1_p & v9a6acd;
assign v984f2c = hmaster1_p & v84563c | !hmaster1_p & !v984f2b;
assign v9999ba = stateG2_p & v84563c | !stateG2_p & v972fac;
assign v9738d2 = stateG10_1_p & v97388d | !stateG10_1_p & v9738d1;
assign v9d2733 = hbusreq2 & v9d2732 | !hbusreq2 & v9d26f1;
assign v8ea7fc = locked_p & v8ea7fb | !locked_p & v84563c;
assign v9adc10 = hmastlock_p & v9adc0f | !hmastlock_p & v84563c;
assign v8ea7f0 = locked_p & v84563c | !locked_p & v8ea7e9;
assign v9a6aaf = hbusreq0_p & v9a6aae | !hbusreq0_p & v9a6aad;
assign v9d271d = hready & v9d26ac | !hready & v84563c;
assign v9998a7 = hbusreq0_p & v9998a6 | !hbusreq0_p & !v84563c;
assign v9bae78 = hbusreq1_p & a153c0 | !hbusreq1_p & v84565c;
assign a154a4 = hmaster1_p & a154a2 | !hmaster1_p & a154a3;
assign v8c112c = hmaster1_p & v8c112a | !hmaster1_p & v8c1126;
assign v9baf22 = hmaster0_p & v9baf10 | !hmaster0_p & !v9ed487;
assign v9ed4e4 = decide_p & v9ed4e3 | !decide_p & !v84563c;
assign v9ed4df = hmaster1_p & v9ed4db | !hmaster1_p & v9ed483;
assign v8c116d = hready_p & v8c1165 | !hready_p & !v8c116c;
assign v8ea8e1 = hbusreq0_p & v8ea8df | !hbusreq0_p & v8ea8e0;
assign v98564a = stateA1_p & v866c94 | !stateA1_p & v84563c;
assign v98556d = hmaster1_p & v98555e | !hmaster1_p & v98556c;
assign v973981 = hgrant0_p & v97397d | !hgrant0_p & v973980;
assign v8ea8f8 = hbusreq2_p & v8ea8dd | !hbusreq2_p & v8ea8f7;
assign v8ea887 = stateG10_1_p & v8ea7e9 | !stateG10_1_p & v8ea886;
assign v8ea7fb = stateG2_p & v84563c | !stateG2_p & v8ea7fa;
assign a154a5 = hlock0_p & v84563c | !hlock0_p & a154a4;
assign v973a37 = hmaster0_p & v97391e | !hmaster0_p & v973a0b;
assign v8ea921 = hbusreq2 & v8ea91f | !hbusreq2 & v8ea920;
assign a15445 = hbusreq0_p & v845648 | !hbusreq0_p & a15444;
assign v984f4b = hbusreq0 & v984f42 | !hbusreq0 & v984f4a;
assign v984ea8 = hmaster0_p & v984ea7 | !hmaster0_p & v984e66;
assign v996569 = hmaster0_p & v996563 | !hmaster0_p & v8ea7e9;
assign v9baf3e = hbusreq2 & v9baf3d | !hbusreq2 & !v84563c;
assign a154ff = hgrant1_p & a153c0 | !hgrant1_p & v84565c;
assign v984eea = hbusreq0_p & v984ee9 | !hbusreq0_p & v984ee8;
assign v984ee9 = hlock0_p & v984ee6 | !hlock0_p & v984ee8;
assign v9ed530 = decide_p & v9ed52f | !decide_p & v9ed4c6;
assign v8ea7f5 = hmaster1_p & v8ea7e9 | !hmaster1_p & v8ea7f4;
assign v984f3c = hmaster1_p & v9855fb | !hmaster1_p & v9855fa;
assign a14d8d = hmaster0_p & a154d4 | !hmaster0_p & !v84563c;
assign v9d27b1 = decide_p & v9d2792 | !decide_p & v9d27b0;
assign v8ea865 = hmaster1_p & v8ea863 | !hmaster1_p & v8ea81d;
assign v9ed42e = hburst0_p & v84563c | !hburst0_p & v9ed42d;
assign v85a40d = stateG3_0_p & v84563c | !stateG3_0_p & v84566c;
assign v9adc6d = hgrant0_p & v9adc5b | !hgrant0_p & v9adc6c;
assign v9d2704 = hgrant0_p & v84563c | !hgrant0_p & !v9d2703;
assign v9854ba = hbusreq2 & v9854b7 | !hbusreq2 & v9854b9;
assign v9adbf3 = hmaster0_p & v9adbf2 | !hmaster0_p & v9adbf1;
assign v9a6a9c = decide_p & v9a6a9b | !decide_p & v9a6a9a;
assign v9adcad = hbusreq1_p & v9adcaa | !hbusreq1_p & !v9adcac;
assign a15417 = hburst1_p & v8e798b | !hburst1_p & !v84563c;
assign v985577 = hmastlock_p & v985576 | !hmastlock_p & v84563c;
assign v9738fd = hgrant2_p & v9738bc | !hgrant2_p & v9738fc;
assign v8ea92b = hmaster1_p & v8ea823 | !hmaster1_p & v8ea918;
assign v9855ea = hgrant0_p & v9855e9 | !hgrant0_p & v98559c;
assign a14d4d = decide_p & a14d4c | !decide_p & v84565c;
assign v999969 = decide_p & v999930 | !decide_p & v84565e;
assign v984ed8 = hmaster1_p & v984ea7 | !hmaster1_p & v984ead;
assign a153c4 = hmaster0_p & v84563c | !hmaster0_p & a153ba;
assign v984f4d = hmaster1_p & v84563c | !hmaster1_p & v9855fe;
assign v985639 = hbusreq2 & v985630 | !hbusreq2 & v985638;
assign a15422 = hbusreq1_p & a15421 | !hbusreq1_p & v84563c;
assign v984f91 = hgrant2_p & v984f8d | !hgrant2_p & v984f90;
assign v9ed435 = hlock1_p & v9ed42b | !hlock1_p & v9ed434;
assign v9739a0 = hmaster1_p & v97399f | !hmaster1_p & !v9738d4;
assign v9999e2 = hbusreq0 & v9999dc | !hbusreq0 & v9999e1;
assign v9baf82 = locked_p & v9ed415 | !locked_p & !v84563c;
assign v9ed42f = stateA1_p & v84563c | !stateA1_p & v9ed42e;
assign v985511 = hbusreq0_p & v985510 | !hbusreq0_p & v98550f;
assign v9998e2 = hbusreq2_p & v9998cf | !hbusreq2_p & v9998e1;
assign v9f357b = hgrant2_p & v9f3575 | !hgrant2_p & v9f3578;
assign v9d2790 = hbusreq0 & v9d26e3 | !hbusreq0 & v9d278f;
assign v984eef = hready & v8ea7e5 | !hready & !v9999bc;
assign v9d277b = hbusreq2 & v9d2774 | !hbusreq2 & v9d277a;
assign v9854a4 = hbusreq1_p & v98548f | !hbusreq1_p & v84563c;
assign v999906 = busreq_p & v9ed457 | !busreq_p & v999905;
assign v9d274a = jx0_p & v9d26dd | !jx0_p & v9d2749;
assign v8ea8b6 = hmaster1_p & v8ea8b4 | !hmaster1_p & v8ea882;
assign v99992b = hmaster1_p & v99992a | !hmaster1_p & !v99990b;
assign v8e79a0 = hmaster1_p & v8e799a | !hmaster1_p & v8e799f;
assign v9d272e = hready_p & v9d270b | !hready_p & !v9d272d;
assign v9965ad = hmaster1_p & v9965ab | !hmaster1_p & v996566;
assign v9d2756 = hready_p & v84564b | !hready_p & v9d2755;
assign v9ed41a = hbusreq1_p & v9ed419 | !hbusreq1_p & v84563c;
assign v8ea85f = hmaster1_p & v8ea85e | !hmaster1_p & v8ea806;
assign v9ed49b = hmaster0_p & v9ed43c | !hmaster0_p & v9ed442;
assign a154c3 = stateG2_p & v84563c | !stateG2_p & a154c2;
assign v9baf53 = hgrant1_p & v9baf52 | !hgrant1_p & !v9baf50;
assign v9ed41d = locked_p & v84563c | !locked_p & !v973893;
assign v8e798c = hburst1_p & v8e798b | !hburst1_p & v8e7989;
assign v996597 = hmaster0_p & v8ea7f1 | !hmaster0_p & v996572;
assign v8c1172 = stateG2_p & v84563c | !stateG2_p & !v8c1171;
assign v999928 = hbusreq0 & v999927 | !hbusreq0 & !v999912;
assign v9d2707 = hbusreq0_p & v9d2706 | !hbusreq0_p & v845647;
assign v9d2781 = hmaster0_p & v9d2780 | !hmaster0_p & v845647;
assign v9d27a9 = hgrant1_p & v84563c | !hgrant1_p & !v9d26ac;
assign v985635 = hmaster1_p & v985634 | !hmaster1_p & !v98562c;
assign v973925 = hmaster0_p & v9738e1 | !hmaster0_p & v9738ec;
assign v8ea8d7 = hlock0 & v8ea8d6 | !hlock0 & v8ea8d5;
assign v9a6ac8 = hgrant1_p & v84563c | !hgrant1_p & v9a6ab1;
assign v9d27a4 = hgrant0_p & v84563c | !hgrant0_p & v9d27a3;
assign v9855c6 = hmaster0_p & v9854fa | !hmaster0_p & v9854b3;
assign v9854d4 = hmaster1_p & v9854d2 | !hmaster1_p & v9854d3;
assign v8ea820 = hgrant1_p & v8ea7ef | !hgrant1_p & !v8ea7ea;
assign a3134e = stateG3_0_p & v84566c | !stateG3_0_p & v84563c;
assign v9ed4c5 = hbusreq1_p & v845660 | !hbusreq1_p & !v9f3569;
assign v9d271a = hmaster0_p & v845641 | !hmaster0_p & !v84563c;
assign v8c1122 = hlock1_p & v8c1119 | !hlock1_p & !v84563c;
assign v9965bd = hmaster0_p & v9adc64 | !hmaster0_p & v996552;
assign a154a3 = hmaster0_p & v84565c | !hmaster0_p & v84563c;
assign v9a6a97 = hmastlock_p & v9a6a96 | !hmastlock_p & v84563c;
assign v9738a7 = hbusreq1_p & v9738a6 | !hbusreq1_p & !v97388d;
assign v9d26fb = hmaster0_p & v9d26f8 | !hmaster0_p & v9d26fa;
assign v985647 = hbusreq0 & v985646 | !hbusreq0 & v985645;
assign v9d2692 = hbusreq1 & v9d2691 | !hbusreq1 & !v84563c;
assign v9baf3c = hbusreq0_p & v9baf3b | !hbusreq0_p & v9baf37;
assign v9a6ac1 = stateG10_1_p & v84563c | !stateG10_1_p & v9a6abb;
assign v9baf7e = hbusreq0_p & v9baf7b | !hbusreq0_p & !v9baf7d;
assign v9739ba = hmaster0_p & v973885 | !hmaster0_p & !v973966;
assign v985564 = hmastlock_p & v985563 | !hmastlock_p & !v84563c;
assign v9f356b = hmaster0_p & v9f356a | !hmaster0_p & v9f3568;
assign v8ea90f = hmaster1_p & v8ea909 | !hmaster1_p & v8ea90e;
assign v9999b3 = decide_p & v9999ad | !decide_p & !v84565e;
assign v9ed44b = hburst0 & v84563c | !hburst0 & v9ed44a;
assign v9baec8 = hbusreq0 & v9baeb5 | !hbusreq0 & v9baec7;
assign v9739dc = hbusreq0_p & v9739db | !hbusreq0_p & v9739ac;
assign v9ed4c0 = hmaster0_p & v84563c | !hmaster0_p & !v9ed4bf;
assign v985605 = hmaster0_p & v84563c | !hmaster0_p & v985604;
assign v984e54 = hbusreq1_p & v98564f | !hbusreq1_p & v984e53;
assign v999921 = hmastlock_p & v9ed43e | !hmastlock_p & v845666;
assign v9adc78 = hmaster0_p & v9adc76 | !hmaster0_p & !v9adc77;
assign v9bafa1 = jx1_p & v9baef2 | !jx1_p & v9bafa0;
assign v8c1137 = stateG2_p & v84563c | !stateG2_p & v8c1132;
assign v8ea8ce = stateG10_1_p & v8ea7ea | !stateG10_1_p & !v8ea8cd;
assign v8c113b = hmaster0_p & v8c113a | !hmaster0_p & v8c111a;
assign v973886 = locked_p & v84563c | !locked_p & !v973885;
assign v996554 = hmaster0_p & v996553 | !hmaster0_p & v9adbf1;
assign v8ea8d3 = hmaster1_p & v8ea823 | !hmaster1_p & v8ea8d2;
assign a15484 = hbusreq0_p & a15409 | !hbusreq0_p & a15483;
assign v8ea85b = hready_p & v8ea846 | !hready_p & v8ea85a;
assign v984f7f = hmaster1_p & v984f70 | !hmaster1_p & v984f7e;
assign v9855ce = hbusreq0_p & v9855cc | !hbusreq0_p & v9855cd;
assign v9ed4c7 = decide_p & v9ed4c4 | !decide_p & v9ed4c6;
assign v9d27b3 = hgrant2_p & v9d2795 | !hgrant2_p & v9d27b2;
assign v9739d4 = hmaster1_p & v973991 | !hmaster1_p & v9738a8;
assign v8e79c3 = stateG10_1_p & v84563c | !stateG10_1_p & v8e79c2;
assign v8ea836 = hbusreq0_p & v8ea817 | !hbusreq0_p & v8ea835;
assign a14d4c = hgrant0_p & v845642 | !hgrant0_p & a14d4b;
assign a153c1 = hlock1_p & v84563c | !hlock1_p & a153c0;
assign v984e60 = hmaster0_p & v984e5f | !hmaster0_p & v84563c;
assign v99655f = hlock2_p & v996558 | !hlock2_p & v99655e;
assign v8c112e = hbusreq0_p & v8c112d | !hbusreq0_p & v8c112c;
assign v8ea840 = hlock2 & v8ea83d | !hlock2 & v8ea83f;
assign v9ed45e = stateA1_p & a2bd3d | !stateA1_p & !a154c2;
assign v9998eb = stateG2_p & v84563c | !stateG2_p & v9998ea;
assign v8c1152 = hbusreq1_p & v8c1145 | !hbusreq1_p & !v8c1151;
assign v9baf1c = hburst0 & v972fac | !hburst0 & v9baf1b;
assign v984f2d = hlock0_p & v984f2c | !hlock0_p & v984f27;
assign v9854b9 = hmaster1_p & v9854b8 | !hmaster1_p & v84563c;
assign v8c1180 = hbusreq2_p & v8c1163 | !hbusreq2_p & v8c117f;
assign v984f5a = hbusreq0_p & v984f57 | !hbusreq0_p & v984f59;
assign v985543 = hburst1_p & v9854bd | !hburst1_p & a3134f;
assign v9d2669 = stateA1_p & a2bd3d | !stateA1_p & v85a40d;
assign a2fb4d = stateA1_p & v84563c | !stateA1_p & a2fb4c;
assign v973a38 = hmaster1_p & v973a37 | !hmaster1_p & !v973a0c;
assign v9ed4e5 = hready_p & v9ed4d2 | !hready_p & !v9ed4e4;
assign v8c1124 = hmaster0_p & v8c1123 | !hmaster0_p & v8c1119;
assign v8ea864 = hmaster1_p & v8ea863 | !hmaster1_p & v8ea816;
assign v9d26f5 = hready_p & v84564b | !hready_p & !v9d26f4;
assign v8c1173 = stateG2_p & v84563c | !stateG2_p & v8c1171;
assign v9baf81 = hbusreq2 & v9baf80 | !hbusreq2 & v84563c;
assign v973913 = hmaster0_p & v973886 | !hmaster0_p & v973895;
assign v8ea7e4 = stateG2_p & v84563c | !stateG2_p & v8ea7e3;
assign v8e79d4 = hmaster1_p & v8e79d3 | !hmaster1_p & v8e79b6;
assign v973a05 = hgrant1_p & v9738c3 | !hgrant1_p & v973893;
assign v9baf27 = stateA1_p & a2fb4c | !stateA1_p & !a153cb;
assign v996578 = hready_p & v996560 | !hready_p & !v996577;
assign v9739ec = hmaster0_p & v9739eb | !hmaster0_p & v973889;
assign v9ed52d = decide_p & v9ed4f7 | !decide_p & v84563c;
assign v999912 = hbusreq0_p & v999911 | !hbusreq0_p & v84563c;
assign v97398d = hmaster0_p & v973885 | !hmaster0_p & !v973893;
assign v8ea89c = hbusreq0 & v8ea893 | !hbusreq0 & v8ea89b;
assign a153d0 = stateG2_p & v84563c | !stateG2_p & !v972fac;
assign a14d42 = hbusreq0_p & a154f0 | !hbusreq0_p & a14d40;
assign stateG3_2 = !v8ea93c;
assign v984ecf = hgrant0_p & v84563c | !hgrant0_p & v984ece;
assign v8ea874 = hbusreq0 & v8ea86f | !hbusreq0 & v8ea873;
assign v9ed4a9 = hburst1 & v9ed4a2 | !hburst1 & v9ed4a8;
assign v9baf31 = hbusreq1 & v9baf30 | !hbusreq1 & v9ed481;
assign v985508 = hbusreq2 & v9854e3 | !hbusreq2 & v985507;
assign v8ea920 = hlock2 & v8ea91d | !hlock2 & v8ea91f;
assign v8e79bb = hmaster0_p & v8e79ba | !hmaster0_p & v84563c;
assign v9d272a = hgrant0_p & v9d2726 | !hgrant0_p & v9d2729;
assign v98556f = stateG2_p & v84563c | !stateG2_p & !v9854c0;
assign v9855d4 = hgrant0_p & v9855d3 | !hgrant0_p & v98553d;
assign v9854a2 = hbusreq1_p & v9854a1 | !hbusreq1_p & v84563c;
assign v9ed42c = stateG2_p & v84563c | !stateG2_p & v9ed424;
assign a154bc = decide_p & a154bb | !decide_p & v84565c;
assign v9adc54 = hbusreq1_p & v9adbfe | !hbusreq1_p & v8ea7e9;
assign v9a6a9a = hmaster1_p & v9a6a99 | !hmaster1_p & v84563c;
assign v985538 = locked_p & v985537 | !locked_p & v84563c;
assign v9baf95 = hbusreq0_p & v9baf94 | !hbusreq0_p & !v84563c;
assign v8ea8a0 = hready_p & v8ea80e | !hready_p & v8ea89f;
assign v8e79ae = hmaster1_p & v84563c | !hmaster1_p & v8e7994;
assign v8ea852 = hmaster1_p & v8ea851 | !hmaster1_p & v8ea7f2;
assign v8ea878 = hready_p & v8ea862 | !hready_p & v8ea877;
assign v9d27c2 = hready_p & v84564b | !hready_p & !v9d2681;
assign v9d26d8 = hbusreq0 & v9d26d6 | !hbusreq0 & !v9d26d7;
assign v973a0b = hbusreq1_p & v9738d6 | !hbusreq1_p & v973893;
assign v8e79ab = hmaster1_p & v8e79aa | !hmaster1_p & v84563c;
assign v9adc6b = hmaster1_p & v9adc69 | !hmaster1_p & v9adc3d;
assign v8ea8da = hbusreq2 & v8ea8d8 | !hbusreq2 & v8ea8d9;
assign v8e7997 = decide_p & v8e7996 | !decide_p & v8e7995;
assign v985531 = hmaster0_p & v84563c | !hmaster0_p & v9854a2;
assign v9998dc = hgrant0_p & v9998db | !hgrant0_p & !a14d6e;
assign v99991b = hmaster0_p & v9baf2f | !hmaster0_p & !v9ed481;
assign v9965a3 = decide_p & v996571 | !decide_p & v9965a2;
assign v999904 = stateA1_p & v999903 | !stateA1_p & !v9ed455;
assign v973a33 = hmaster1_p & v97398d | !hmaster1_p & v973a02;
assign a154d5 = hmaster1_p & a154d2 | !hmaster1_p & !a154d4;
assign v984f44 = locked_p & v984f43 | !locked_p & v84563c;
assign v9999bc = stateG2_p & v84563c | !stateG2_p & v9999bb;
assign v9738c3 = locked_p & v973892 | !locked_p & v97388d;
assign v9f3569 = stateG10_1_p & v84563c | !stateG10_1_p & !v845660;
assign a15433 = hbusreq1_p & v845648 | !hbusreq1_p & !v84563c;
assign v984edf = hready_p & v984ed1 | !hready_p & v984ede;
assign v8ea7f9 = hmaster1_p & v84563c | !hmaster1_p & v8ea7e7;
assign a1541f = hmastlock_p & a1541e | !hmastlock_p & !v84563c;
assign v9999c2 = hburst1 & v9999ba | !hburst1 & v9999c1;
assign v9adc56 = hmaster1_p & v9adc55 | !hmaster1_p & !v9adc05;
assign v9d272c = hbusreq2 & v9d2723 | !hbusreq2 & v9d272b;
assign v9bae7e = hburst0 & v9ed42c | !hburst0 & v9bae7d;
assign v9baea2 = hmaster1_p & a154a2 | !hmaster1_p & v84565c;
assign v9d269f = hmaster1_p & v9d269d | !hmaster1_p & v9d269e;
assign v98559c = hmaster1_p & v98559a | !hmaster1_p & v98559b;
assign v985497 = locked_p & v985496 | !locked_p & v84563c;
assign v8e7995 = hmaster1_p & v8e7994 | !hmaster1_p & v84563c;
assign v9b40c3 = hgrant2_p & v9b40c0 | !hgrant2_p & !v9b40c2;
assign v9ed431 = hburst1 & v9ed42c | !hburst1 & v9ed430;
assign v9adcde = hgrant1_p & v9adc75 | !hgrant1_p & v9adcdd;
assign v9998a6 = hlock0_p & v9998a5 | !hlock0_p & !v84563c;
assign v8ea8ae = hbusreq0 & v8ea8ac | !hbusreq0 & v8ea8ad;
assign v98557c = hgrant1_p & v84563c | !hgrant1_p & v9d2691;
assign v9ed4ed = decide_p & v9ed4ec | !decide_p & v9ed4c6;
assign v9738ff = hmaster1_p & v9738fe | !hmaster1_p & v97389c;
assign v999931 = decide_p & v999930 | !decide_p & !v84563c;
assign v8ea8f2 = hbusreq0 & v8ea8ef | !hbusreq0 & v8ea8f1;
assign v9baf77 = hmaster0_p & v84565c | !hmaster0_p & v9ed42b;
assign v9998ab = hlock0_p & v9998aa | !hlock0_p & !v84563c;
assign v9baf9c = hready_p & v9baf9a | !hready_p & !v9baf9b;
assign v9d26c8 = hmaster1_p & v9d26c7 | !hmaster1_p & !v9d2671;
assign v985559 = hmaster0_p & v985558 | !hmaster0_p & v84563c;
assign v8e79da = hgrant2_p & v8e79d1 | !hgrant2_p & v8e79d9;
assign v9bae9e = hready_p & v84563c | !hready_p & v9bae9d;
assign v9baea9 = hbusreq0 & v9baea7 | !hbusreq0 & v9baea8;
assign v9adcf0 = hbusreq0_p & v9adcee | !hbusreq0_p & v9adcef;
assign v9738ce = hgrant1_p & v97388a | !hgrant1_p & v973889;
assign v887862 = stateG3_1_p & v84563c | !stateG3_1_p & v845658;
assign v9ed4f0 = hgrant2_p & v9ed4e5 | !hgrant2_p & v9ed4ef;
assign v9ed491 = hmaster1_p & v9ed48d | !hmaster1_p & v9ed483;
assign v9855c1 = hmaster0_p & v9ed423 | !hmaster0_p & !v98556b;
assign v9d268a = hgrant1_p & v845647 | !hgrant1_p & !v9d2689;
assign v8c20de = decide_p & v8c20dd | !decide_p & v84565c;
assign v985548 = hmastlock_p & v985547 | !hmastlock_p & v84563c;
assign v985616 = hmastlock_p & v985615 | !hmastlock_p & v84563c;
assign v9adc47 = stateG10_1_p & v9adc45 | !stateG10_1_p & v9adc46;
assign v9739a8 = hbusreq1_p & v9738d6 | !hbusreq1_p & v9739a7;
assign v9933bb = decide_p & v9933ba | !decide_p & v9933b9;
assign a153cc = stateG2_p & v84563c | !stateG2_p & a153cb;
assign v9ed4a5 = hmastlock_p & v9ed4a4 | !hmastlock_p & !v84563c;
assign v9adc5c = hlock0_p & v9adc5b | !hlock0_p & v9adc1c;
assign v985596 = hbusreq0_p & v98558a | !hbusreq0_p & v985595;
assign v9adcd2 = decide_p & v9adcd1 | !decide_p & !v9adc7e;
assign v99991e = hbusreq0_p & v99991d | !hbusreq0_p & !v84563c;
assign v8ea842 = decide_p & v8ea7ee | !decide_p & v8ea841;
assign v9999e0 = hbusreq0_p & v9999df | !hbusreq0_p & !v84563c;
assign v9739fe = hmaster1_p & v9738bd | !hmaster1_p & v97397b;
assign v8ea88c = hbusreq1 & v8ea88b | !hbusreq1 & v8ea831;
assign v8ea8a2 = hmaster0_p & v84563c | !hmaster0_p & v8ea81b;
assign v99990c = hmaster1_p & v99990a | !hmaster1_p & !v99990b;
assign v9854cf = hlock1_p & v9854ce | !hlock1_p & !v84563c;
assign v9ed4d8 = hmaster1_p & v9ed4d3 | !hmaster1_p & v9ed489;
assign v984f26 = hmaster0_p & v98562c | !hmaster0_p & !v84563c;
assign v8c1168 = hmaster1_p & v8c1167 | !hmaster1_p & v8c1126;
assign v9d2764 = hmaster0_p & v9d275d | !hmaster0_p & v84563c;
assign v985528 = hmaster0_p & v985521 | !hmaster0_p & v985527;
assign v996587 = hmaster0_p & v996586 | !hmaster0_p & !v9adc27;
assign v8ea8e9 = hready_p & v8ea846 | !hready_p & v8ea8e8;
assign v8c1139 = hmastlock_p & v8c1138 | !hmastlock_p & !v84563c;
assign v8ea857 = hlock2 & v8ea850 | !hlock2 & v8ea856;
assign v9a6ad7 = hbusreq0_p & v9a6aae | !hbusreq0_p & v9a6ad6;
assign v985556 = hready & v985552 | !hready & v985555;
assign v8e79b8 = hgrant0_p & v8e79b0 | !hgrant0_p & v8e79b7;
assign v9965b4 = hmaster0_p & v9adbec | !hmaster0_p & v996552;
assign v854658 = hmaster1_p & v845646 | !hmaster1_p & !v86292d;
assign v9855a1 = hbusreq1_p & v9855a0 | !hbusreq1_p & !v84563c;
assign a154ef = hmaster1_p & a154ee | !hmaster1_p & !a154d4;
assign v9d26a4 = hbusreq1 & v845641 | !hbusreq1 & v84563c;
assign v9adc01 = stateG10_1_p & v9adbee | !stateG10_1_p & v8ea7ea;
assign v973949 = hmaster1_p & v9738a5 | !hmaster1_p & v973948;
assign a14d5b = jx0_p & a154a1 | !jx0_p & a14d5a;
assign v996566 = hmaster0_p & v996563 | !hmaster0_p & !v8ea7ea;
assign v984ef5 = hbusreq0_p & v984ef4 | !hbusreq0_p & v984ee8;
assign v999978 = hmaster1_p & v999977 | !hmaster1_p & !v99990b;
assign v9adc7f = hmaster0_p & v9adc75 | !hmaster0_p & !v84563c;
assign v8ea903 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea81b;
assign v9738d0 = hlock1_p & v9738ce | !hlock1_p & v9738cf;
assign v9adc3a = hbusreq1_p & v9adc29 | !hbusreq1_p & v9adc39;
assign v985588 = hmaster0_p & v985521 | !hmaster0_p & v9ed423;
assign v8ea811 = busreq_p & v8ea810 | !busreq_p & v84563c;
assign a15449 = hmaster0_p & v845646 | !hmaster0_p & a15433;
assign v9ed414 = hburst0 & v9ed412 | !hburst0 & v9ed413;
assign v87f892 = stateA1_p & v84563c | !stateA1_p & v866c94;
assign v984f55 = hlock2_p & v984f4c | !hlock2_p & v984f54;
assign v973a13 = hmaster0_p & v973963 | !hmaster0_p & !v9739a8;
assign v8ea892 = hbusreq0_p & v8ea891 | !hbusreq0_p & v8ea82e;
assign v8ea815 = hmaster0_p & v8ea814 | !hmaster0_p & v8ea7ef;
assign v9d26fd = hmaster1_p & v9d26fb | !hmaster1_p & v9d26fc;
assign v99659b = stateG10_1_p & v9adbee | !stateG10_1_p & !v99659a;
assign v9738e9 = hmaster1_p & v9738e4 | !hmaster1_p & !v9738e8;
assign v8ea816 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea7e9;
assign v9adc1c = hmaster1_p & v9adc1a | !hmaster1_p & v9adc1b;
assign v9d26f2 = hbusreq2 & v9d26ea | !hbusreq2 & v9d26f1;
assign v9baef1 = hbusreq2_p & v9baef0 | !hbusreq2_p & !v9baea0;
assign v8e79a8 = hlock2_p & v8e79a2 | !hlock2_p & v8e79a7;
assign v8ea93b = jx0_p & v8ea8f8 | !jx0_p & v8ea93a;
assign v9854df = hmaster0_p & v84563c | !hmaster0_p & v9854b3;
assign a1540d = hready_p & a153c9 | !hready_p & a1540c;
assign v9baef5 = decide_p & v9baef4 | !decide_p & v84563c;
assign v985617 = locked_p & v985616 | !locked_p & !v84563c;
assign v9ed454 = hburst1_p & v96ef3e | !hburst1_p & !v84563c;
assign v9855ee = hbusreq0 & v9855ea | !hbusreq0 & v9855ed;
assign v9adc0e = hlock2_p & v9adc08 | !hlock2_p & v9adc0d;
assign v9baf0c = hmastlock_p & v9baf0b | !hmastlock_p & v84563c;
assign v9854d9 = hready & v9854d8 | !hready & !v972fac;
assign v973955 = hmaster1_p & v9738b7 | !hmaster1_p & !v973938;
assign v9854b0 = hmaster0_p & v84563c | !hmaster0_p & v9854af;
assign v9adc27 = hbusreq1_p & v9adc26 | !hbusreq1_p & v9adbee;
assign v9ed4cf = hmaster0_p & v845646 | !hmaster0_p & v9ed4bf;
assign v8e798a = stateG3_0_p & v84566c | !stateG3_0_p & !v887862;
assign v8ea8eb = hbusreq0_p & v8ea8b5 | !hbusreq0_p & v8ea8ea;
assign v9baf24 = hbusreq0_p & v9baf21 | !hbusreq0_p & v9baf23;
assign v8ea8a9 = hbusreq0 & v8ea8a6 | !hbusreq0 & v8ea8a8;
assign v9ed473 = hmaster1_p & v9ed46f | !hmaster1_p & v9ed472;
assign v9738ea = hgrant1_p & v97388e | !hgrant1_p & v97388d;
assign v9ed4be = hlock1_p & v9ed4bd | !hlock1_p & v84563c;
assign v9999a0 = hlock0_p & v99999f | !hlock0_p & v84563c;
assign v9bae85 = hlock1_p & v9bae83 | !hlock1_p & v9bae84;
assign v8ea84c = hmaster1_p & v8ea84b | !hmaster1_p & v8ea7f2;
assign v9d26e5 = hmaster1_p & v84563c | !hmaster1_p & v9d2671;
assign v8c1140 = hlock0_p & v8c113f | !hlock0_p & v84563c;
assign v9ed4a1 = hbusreq0_p & v9ed49a | !hbusreq0_p & v9ed4a0;
assign v999934 = hbusreq0_p & v999933 | !hbusreq0_p & !v84563c;
assign v9baf35 = hmaster1_p & v9baf2f | !hmaster1_p & !v9baf34;
assign v973a41 = hmaster1_p & v9739b3 | !hmaster1_p & !v973a10;
assign a4ce72 = hbusreq2_p & v84563c | !hbusreq2_p & v845662;
assign v996599 = hgrant1_p & v996572 | !hgrant1_p & !v8ea7ea;
assign v8ea82b = stateG10_1_p & v8ea7e9 | !stateG10_1_p & v8ea82a;
assign v9adce6 = hmaster1_p & v9adce5 | !hmaster1_p & !v9adcba;
assign v98550f = hmaster1_p & v985509 | !hmaster1_p & v9854df;
assign v9adc1a = hmaster0_p & v9adbeb | !hmaster0_p & v9adbee;
assign v9739cb = hgrant0_p & v9738df | !hgrant0_p & v9739ca;
assign v9999ae = decide_p & v9999ad | !decide_p & v84563c;
assign v9adbf7 = hbusreq0_p & v9adbf4 | !hbusreq0_p & v9adbf6;
assign v9d26ef = hlock0_p & v9d26ec | !hlock0_p & v9d26ee;
assign v973922 = hgrant0_p & v973918 | !hgrant0_p & v973921;
assign v9ed4af = hgrant1_p & v84565c | !hgrant1_p & !v84565c;
assign v973916 = hlock0_p & v973914 | !hlock0_p & !v973915;
assign v9854a6 = hmaster1_p & v9854a3 | !hmaster1_p & v9854a5;
assign v999975 = hbusreq2 & v999970 | !hbusreq2 & !v999974;
assign v9738e4 = hmaster0_p & v9738e1 | !hmaster0_p & v9738e3;
assign v9933c9 = hgrant0_p & v9933bf | !hgrant0_p & v9933c8;
assign v97399b = hmaster1_p & v973991 | !hmaster1_p & v9738c0;
assign v9ed4ab = hmastlock_p & v9ed4aa | !hmastlock_p & !v84563c;
assign v9855f6 = decide_p & v9855ca | !decide_p & v9855f5;
assign v8ea91b = hmaster1_p & v8ea909 | !hmaster1_p & v8ea91a;
assign v9d278b = hbusreq2_p & v9d276d | !hbusreq2_p & v9d278a;
assign v973900 = hmaster1_p & v9738fe | !hmaster1_p & v97389f;
assign v9965c2 = hmaster1_p & v9965c1 | !hmaster1_p & !v996590;
assign v9738f9 = hbusreq0_p & v9738f7 | !hbusreq0_p & v9738f8;
assign v999982 = hbusreq2 & v99997c | !hbusreq2 & v999981;
assign v9d2670 = hmaster0_p & v9d266f | !hmaster0_p & !v84563c;
assign v973a45 = hgrant0_p & v973a42 | !hgrant0_p & v973a44;
assign v9ed4b5 = hmaster0_p & v9ed4b4 | !hmaster0_p & v9ed4b1;
assign v9d2758 = hgrant0_p & v84563c | !hgrant0_p & v9d2757;
assign v8ea823 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea822;
assign v8ea84a = hbusreq0_p & v8ea848 | !hbusreq0_p & v8ea849;
assign v9965d1 = hbusreq2_p & v9965a5 | !hbusreq2_p & v9965d0;
assign v8e79a5 = hmaster1_p & v8e79a3 | !hmaster1_p & v8e799f;
assign v9739a3 = hbusreq0_p & v9739a0 | !hbusreq0_p & v9739a2;
assign v9adcb2 = hbusreq0_p & v9adcaf | !hbusreq0_p & v9adcb1;
assign v9d2774 = hbusreq0 & v9d2771 | !hbusreq0 & v9d2773;
assign v985560 = hmaster1_p & v98555e | !hmaster1_p & v98555f;
assign v84566e = stateG3_2_p & v84563c | !stateG3_2_p & !v84563c;
assign v984f4e = hlock0_p & v984f4d | !hlock0_p & !v84563c;
assign v9854de = hmaster1_p & v9854d2 | !hmaster1_p & v9854dd;
assign v973a2e = hready_p & v973a28 | !hready_p & v973a2d;
assign v985623 = hmastlock_p & v985622 | !hmastlock_p & v84563c;
assign v845662 = hgrant2_p & v84563c | !hgrant2_p & !v84563c;
assign v9965d2 = jx0_p & v9965d1 | !jx0_p & v84563c;
assign v8ea915 = hgrant0_p & v8ea914 | !hgrant0_p & v8ea910;
assign v9baf6f = hbusreq1 & v973893 | !hbusreq1 & v84563c;
assign v985625 = hmaster0_p & v985624 | !hmaster0_p & v9854d0;
assign v984e63 = hbusreq0_p & v984e62 | !hbusreq0_p & v84563c;
assign v9ed432 = hburst0 & v9ed42c | !hburst0 & v9ed431;
assign v985525 = locked_p & v985524 | !locked_p & !v84563c;
assign v9adcc8 = hmaster1_p & v9adc7f | !hmaster1_p & v9adcc7;
assign v9adc75 = hmastlock_p & v845668 | !hmastlock_p & !v84563c;
assign v9ed420 = hmaster0_p & v84563c | !hmaster0_p & v9ed41f;
assign v985599 = hbusreq1_p & v845660 | !hbusreq1_p & v84563c;
assign v9baf6d = hbusreq1 & v9ed41d | !hbusreq1 & v84565c;
assign v9adc91 = hbusreq0_p & v9adc90 | !hbusreq0_p & v9adc8e;
assign v985517 = hbusreq0_p & v985516 | !hbusreq0_p & v985515;
assign v8ea927 = decide_p & v8ea7ee | !decide_p & v8ea8f0;
assign v97397f = hmaster1_p & v9738f6 | !hmaster1_p & v973967;
assign v9999ee = hbusreq2_p & v9999ed | !hbusreq2_p & v9999b5;
assign v9ed427 = stateA1_p & v84563c | !stateA1_p & v9ed426;
assign v99993a = hmaster1_p & v999938 | !hmaster1_p & v999939;
assign v9adc92 = hlock2_p & v9adc8d | !hlock2_p & v9adc91;
assign v9ed4e1 = hbusreq0_p & v9ed4df | !hbusreq0_p & v9ed4e0;
assign v9a6aa3 = hlock1_p & v9a6aa2 | !hlock1_p & v84563c;
assign v9ed438 = hmaster0_p & v84563c | !hmaster0_p & v9ed423;
assign v9baf87 = hgrant1_p & v84563c | !hgrant1_p & v9ed4ac;
assign v9d27a2 = hlock2_p & v9d279d | !hlock2_p & v9d27a1;
assign v9999ef = jx2_p & v9999ee | !jx2_p & v9999b6;
assign v984ece = hbusreq0_p & v984ecd | !hbusreq0_p & v84563c;
assign v97388c = locked_p & v84563c | !locked_p & !v973889;
assign v9999c9 = hlock0_p & v9999c8 | !hlock0_p & v84563c;
assign v9738e0 = stateG10_1_p & v973885 | !stateG10_1_p & !v9738c9;
assign v9d2664 = hburst1 & v9d2663 | !hburst1 & !v84563c;
assign v984ec9 = hbusreq0 & v984ec8 | !hbusreq0 & v985645;
assign v9739f5 = hmaster1_p & v9738a5 | !hmaster1_p & v9739f4;
assign v8ea8b1 = hbusreq2 & v8ea8af | !hbusreq2 & v8ea8b0;
assign v9855e9 = hbusreq0_p & v9855e7 | !hbusreq0_p & v9855e8;
assign v984ea4 = hbusreq0_p & v84563c | !hbusreq0_p & v985645;
assign v8c1160 = hgrant0_p & v8c115a | !hgrant0_p & v8c115f;
assign v984f47 = hmaster1_p & v84563c | !hmaster1_p & v984f46;
assign v99996e = hlock0_p & v99996d | !hlock0_p & !v84563c;
assign v9b40c2 = hready_p & v9b40c1 | !hready_p & !v845654;
assign v9adc37 = hbusreq1_p & v9adc25 | !hbusreq1_p & v9adc36;
assign v97395e = hmaster1_p & v9738cd | !hmaster1_p & !v97395d;
assign v9d26bc = hbusreq2 & v9d26b5 | !hbusreq2 & v9d26bb;
assign v984ebe = decide_p & v985640 | !decide_p & v984ebd;
assign v985540 = hmaster1_p & v84563c | !hmaster1_p & v9854b8;
assign v8c1179 = hmaster1_p & v8c1178 | !hmaster1_p & !v8c1148;
assign v9ed4ea = hbusreq0_p & v9ed4e7 | !hbusreq0_p & v9ed4e9;
assign v984eb6 = hbusreq0_p & v984eb5 | !hbusreq0_p & v985645;
assign v973997 = decide_p & v973993 | !decide_p & v973996;
assign v9854bd = stateG3_2_p & v84563c | !stateG3_2_p & v9854bc;
assign v9998f3 = hlock0_p & v9998f1 | !hlock0_p & v9998f2;
assign v9854c7 = hbusreq1_p & v9d2691 | !hbusreq1_p & v84563c;
assign v8ea8db = decide_p & v8ea7ee | !decide_p & v8ea8da;
assign v8ea937 = hready_p & v8ea80d | !hready_p & v8ea936;
assign v973950 = hlock0_p & v97394e | !hlock0_p & v97394f;
assign v973a3f = hgrant0_p & v973a3c | !hgrant0_p & v973a3e;
assign v97390c = hbusreq0_p & v97390a | !hbusreq0_p & v97390b;
assign v9baf06 = hbusreq1 & v9ed46d | !hbusreq1 & v9ed481;
assign v9adc9c = hready_p & v9adc84 | !hready_p & !v9adc9b;
assign v9739e7 = hbusreq2_p & v9739d1 | !hbusreq2_p & !v9739e6;
assign v98564d = locked_p & v98564c | !locked_p & v84563c;
assign v9a6ab4 = decide_p & v9a6ab0 | !decide_p & v9a6ab3;
assign v99656d = hmaster1_p & v9adc09 | !hmaster1_p & v996566;
assign a153c8 = hlock2_p & a153c5 | !hlock2_p & v845648;
assign v9ed4f9 = decide_p & v9ed4f8 | !decide_p & v84563c;
assign v9baefb = hready_p & v84563c | !hready_p & v9baefa;
assign v98550a = hmaster1_p & v985509 | !hmaster1_p & v9854d3;
assign v9ed469 = hbusreq1_p & v9ed468 | !hbusreq1_p & !v84563c;
assign v9adc8e = hmaster1_p & v9adc7f | !hmaster1_p & v9adc88;
assign v984f37 = hbusreq2 & v984f2f | !hbusreq2 & !v84563c;
assign v9739c8 = decide_p & v9739c6 | !decide_p & v9739c7;
assign v8c20c1 = hgrant1_p & v84563c | !hgrant1_p & !v84565c;
assign v973883 = busreq_p & v86cfb3 | !busreq_p & !v87f892;
assign v973893 = hmastlock_p & v973892 | !hmastlock_p & v84563c;
assign v9998fa = hlock0_p & v9998f9 | !hlock0_p & !v84563c;
assign v9855be = hmaster1_p & v845641 | !hmaster1_p & v9854b3;
assign a153d6 = hmaster1_p & a153d4 | !hmaster1_p & a153d5;
assign v9855ef = hmaster0_p & v9855b0 | !hmaster0_p & v9855b4;
assign v97392f = hmaster0_p & v973885 | !hmaster0_p & !v9738ec;
assign v9d276b = decide_p & v9d274f | !decide_p & !v9d276a;
assign v984ec2 = hmaster1_p & v984ec1 | !hmaster1_p & v98561b;
assign v99658a = hmaster1_p & v9adc28 | !hmaster1_p & !v996589;
assign v98551f = hlock2_p & v985508 | !hlock2_p & v98551e;
assign v985638 = hbusreq0 & v985637 | !hbusreq0 & v84563c;
assign v9d26df = hready & v9d26de | !hready & !v84563c;
assign v9ed47f = hburst1 & a153d0 | !hburst1 & v9ed47e;
assign v984f29 = hbusreq0_p & v984f28 | !hbusreq0_p & v98563c;
assign v984f73 = hmaster0_p & v985642 | !hmaster0_p & !v985592;
assign v9adc20 = hgrant1_p & v9adbec | !hgrant1_p & !v9adc1f;
assign v9adcf7 = jx0_p & v9adc72 | !jx0_p & !v9adcf6;
assign a15494 = decide_p & a15493 | !decide_p & v84565c;
assign v999973 = hbusreq0_p & v999972 | !hbusreq0_p & v84563c;
assign v973999 = hmaster0_p & v973886 | !hmaster0_p & v97388e;
assign v973968 = hmaster1_p & v9738e4 | !hmaster1_p & !v973967;
assign v9739b5 = hmaster0_p & v973885 | !hmaster0_p & !v97388e;
assign v9d27bf = hready_p & v9d27be | !hready_p & v9d27b8;
assign v9d26b7 = hmaster1_p & v9d26b6 | !hmaster1_p & !v9d2671;
assign v9a6aad = hmaster1_p & v9a6aab | !hmaster1_p & v9a6aa7;
assign v9854fd = stateG2_p & v84563c | !stateG2_p & !v8ea7e2;
assign v9a6aa0 = hburst0_p & v8ea7fa | !hburst0_p & v9a6a9f;
assign v9933b9 = hmaster1_p & v9933b8 | !hmaster1_p & v84563c;
assign v9adc23 = stateG10_1_p & v9adc1f | !stateG10_1_p & !v9adc21;
assign v9baf58 = stateG2_p & v84563c | !stateG2_p & !v9baf57;
assign a154f3 = decide_p & a154f2 | !decide_p & v84565c;
assign v9ed444 = hmaster1_p & v9ed441 | !hmaster1_p & v9ed443;
assign v9baf61 = hgrant1_p & v9baf60 | !hgrant1_p & !v9ed41d;
assign v973948 = hmaster0_p & v973945 | !hmaster0_p & v973889;
assign v9ed47a = hbusreq0_p & v9ed473 | !hbusreq0_p & v9ed479;
assign v9738de = hmaster1_p & v9738bd | !hmaster1_p & v9738dd;
assign v9d266d = hready & v9d266c | !hready & !v84563c;
assign v973a18 = hmaster1_p & v9738f2 | !hmaster1_p & !v973a10;
assign v9855f9 = hbusreq2_p & v9855bd | !hbusreq2_p & v9855f8;
assign v9738ac = hlock0_p & v9738a9 | !hlock0_p & v9738ab;
assign v98553d = hmaster1_p & v98553c | !hmaster1_p & v84563c;
assign a15489 = hbusreq1_p & a153b7 | !hbusreq1_p & !v84563c;
assign v97399e = hbusreq0_p & v97399c | !hbusreq0_p & !v97399d;
assign v9998ce = hready_p & v9998af | !hready_p & !v9998cd;
assign v9d2785 = hgrant0_p & v84563c | !hgrant0_p & !v9d2783;
assign v8c114f = hbusreq0_p & v8c113f | !hbusreq0_p & v8c114e;
assign v8ea7e9 = hmastlock_p & v8ecba9 | !hmastlock_p & v84563c;
assign v9d26d4 = hmaster1_p & v9d26d3 | !hmaster1_p & v9d2698;
assign v984e52 = hgrant1_p & v845641 | !hgrant1_p & v98564e;
assign v996592 = hmaster0_p & v99658f | !hmaster0_p & !v996552;
assign v8ea8e4 = hlock0 & v8ea8e3 | !hlock0 & v8ea8e1;
assign v9d268f = hlock1_p & v9d268a | !hlock1_p & v9d268e;
assign v9baf1a = hmastlock_p & v9baf19 | !hmastlock_p & v84563c;
assign v984f5e = stateG10_1_p & v84563c | !stateG10_1_p & v984f5d;
assign v985514 = hmaster1_p & v985513 | !hmaster1_p & v9854d3;
assign v9ed4fd = hbusreq1_p & v9ed4fc | !hbusreq1_p & !v84563c;
assign v9855d9 = hbusreq0_p & v98555a | !hbusreq0_p & v9855d8;
assign v9bae92 = hmastlock_p & a153cb | !hmastlock_p & v84563c;
assign a15432 = hgrant2_p & a1540d | !hgrant2_p & a15431;
assign v9bae79 = hmaster0_p & v84565c | !hmaster0_p & v9bae78;
assign v9adcbd = hmaster1_p & v9adcb6 | !hmaster1_p & !v9adcbc;
assign v8c112d = hlock0_p & v8c112b | !hlock0_p & v8c112c;
assign v9a6aa6 = hmaster1_p & v9a6aa2 | !hmaster1_p & v9a6aa5;
assign v9ed45f = stateG2_p & v84563c | !stateG2_p & !v9ed45e;
assign v9baf36 = hmaster0_p & v9baf32 | !hmaster0_p & !v84563c;
assign v9998f8 = hmaster0_p & v9739eb | !hmaster0_p & v84563c;
assign a15493 = hgrant0_p & a15487 | !hgrant0_p & a15492;
assign v99997f = hlock0_p & v99997e | !hlock0_p & v999925;
assign v9d2680 = hbusreq0 & v9d267e | !hbusreq0 & v9d267f;
assign v9baf51 = hgrant1_p & v9baf4a | !hgrant1_p & !v9baf50;
assign v8e79cd = hmaster0_p & v8e79cc | !hmaster0_p & v84563c;
assign v8ea886 = hgrant1_p & v84563c | !hgrant1_p & v8ea7e9;
assign v9d26c3 = hbusreq0_p & v9d2672 | !hbusreq0_p & v9d26c2;
assign v9baf67 = hgrant1_p & v9baf66 | !hgrant1_p & v9ed419;
assign v9998d4 = hbusreq0_p & v99989d | !hbusreq0_p & v845646;
assign v98562b = hmaster0_p & v84563c | !hmaster0_p & !v98562a;
assign v984f8f = decide_p & v84563c | !decide_p & v984ebb;
assign v98561b = hmaster0_p & v98561a | !hmaster0_p & v84563c;
assign v8c1127 = hmaster1_p & v8c1121 | !hmaster1_p & v8c1126;
assign a14daa = hmaster0_p & a15508 | !hmaster0_p & v8c20c3;
assign v97396b = decide_p & v973960 | !decide_p & v97396a;
assign v97388b = hmaster0_p & v973886 | !hmaster0_p & !v97388a;
assign v9d2773 = hbusreq0_p & v9d26e8 | !hbusreq0_p & v9d2772;
assign v996572 = locked_p & v9adbfe | !locked_p & !v8ea7ea;
assign v9ed4a8 = busreq_p & v845668 | !busreq_p & !v84563c;
assign v985567 = stateG2_p & v84563c | !stateG2_p & v985566;
assign v8e799f = hmaster0_p & v8e799c | !hmaster0_p & v84563c;
assign v9baf47 = hmaster0_p & v9739eb | !hmaster0_p & !v9ed49c;
assign a153cf = hbusreq1_p & a153ce | !hbusreq1_p & v84563c;
assign v973a47 = hready_p & v973a40 | !hready_p & !v973a46;
assign v9855e2 = hmaster1_p & v9855e0 | !hmaster1_p & v985583;
assign v9a6ac4 = hmaster1_p & v9a6aba | !hmaster1_p & v9a6ac3;
assign v8ea882 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea818;
assign v9baf23 = hmaster1_p & v9baf05 | !hmaster1_p & !v9baf22;
assign v999907 = hburst1 & v999906 | !hburst1 & v9baf01;
assign v985494 = stateA1_p & v84563c | !stateA1_p & v985493;
assign v97397c = hmaster1_p & v9738f2 | !hmaster1_p & !v97397b;
assign v9854f7 = stateA1_p & a2bd3d | !stateA1_p & v84563c;
assign v9999b7 = hmaster1_p & v84563c | !hmaster1_p & v9baead;
assign v9adc38 = hmaster0_p & v9adc35 | !hmaster0_p & v9adc37;
assign v8ea7f4 = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea7f0;
assign v9d2796 = hmaster0_p & v9d26f8 | !hmaster0_p & v845647;
assign v98560d = hbusreq0 & v98560c | !hbusreq0 & v84563c;
assign v960f67 = hgrant2_p & v960f65 | !hgrant2_p & v960f66;
assign v9ed4e0 = hmaster1_p & v9ed4db | !hmaster1_p & v9ed489;
assign v9d26cb = hbusreq0_p & v9d2678 | !hbusreq0_p & v9d26ca;
assign v984f66 = hbusreq2 & v984f65 | !hbusreq2 & v84563c;
assign v984ed0 = hbusreq0 & v984ecf | !hbusreq0 & v84563c;
assign v996598 = hmaster1_p & v9adc42 | !hmaster1_p & v996597;
assign v8ea8ca = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea8c9;
assign v8ea8c9 = hbusreq1 & v8ea819 | !hbusreq1 & v8ea8c8;
assign v984ecb = hready_p & v984ec5 | !hready_p & v984eca;
assign v984e59 = hlock1_p & v984e58 | !hlock1_p & v9855ae;
assign v8ea870 = hmaster1_p & v8ea863 | !hmaster1_p & v8ea83a;
assign v9d2689 = hbusreq1 & v9d2688 | !hbusreq1 & v84563c;
assign v9d27b7 = hbusreq2 & v9d27b6 | !hbusreq2 & !v9d2680;
assign v999938 = hmaster0_p & v9baf89 | !hmaster0_p & v9baf8e;
assign v9f3575 = hready_p & v845646 | !hready_p & v9f3574;
assign v9bae9a = hready_p & v9bae8b | !hready_p & !v9bae99;
assign v9855de = hmaster1_p & v9ed423 | !hmaster1_p & v98556c;
assign v9855ca = hbusreq2 & v985512 | !hbusreq2 & v9855c9;
assign v9adc4b = stateG10_1_p & v9adbee | !stateG10_1_p & v9adc4a;
assign v9a6a9b = hlock2_p & v9a6a9a | !hlock2_p & v84563c;
assign v9adca3 = hmaster1_p & v9adc7f | !hmaster1_p & !v9adca2;
assign v9738ca = hbusreq1_p & v9738c9 | !hbusreq1_p & !v973885;
assign v9adc26 = hlock1_p & v9adc25 | !hlock1_p & v9adbee;
assign v9739fa = hmaster1_p & v9738b7 | !hmaster1_p & !v9739e8;
assign v9d2755 = decide_p & v9d274f | !decide_p & !v9d2754;
assign v9baf73 = hmaster0_p & v9baf63 | !hmaster0_p & v9baf72;
assign v84565e = hgrant0_p & v84563c | !hgrant0_p & !v84563c;
assign v8ea933 = hmaster1_p & v8ea867 | !hmaster1_p & v8ea91a;
assign v9baf3d = hbusreq0 & v9baf38 | !hbusreq0 & v9baf3c;
assign v9d26c5 = hbusreq0_p & v9d2674 | !hbusreq0_p & v9d26c4;
assign v98561e = hbusreq0 & v98561d | !hbusreq0 & v84563c;
assign v9965b6 = hmaster0_p & v9adbeb | !hmaster0_p & v996552;
assign v9d274e = hbusreq0 & v9d274c | !hbusreq0 & v9d274d;
assign v9ed4f5 = hmaster1_p & v84563c | !hmaster1_p & !a14d8d;
assign v9d26a0 = hgrant0_p & v84563c | !hgrant0_p & v9d269f;
assign v973a3a = hgrant0_p & v973a34 | !hgrant0_p & v973a39;
assign v9adc6f = decide_p & v9adc57 | !decide_p & v9adc4f;
assign v9854e3 = hbusreq0 & v9854d7 | !hbusreq0 & v9854e2;
assign v9adbf4 = hmaster1_p & v9adbf0 | !hmaster1_p & v9adbf3;
assign v98549b = stateA1_p & v84563c | !stateA1_p & v98549a;
assign v960f65 = hready_p & v84563c | !hready_p & !v845652;
assign v9d2735 = hready_p & v84564b | !hready_p & !v9d2734;
assign v9ed41c = hmaster1_p & v9ed418 | !hmaster1_p & v9ed41b;
assign v973a01 = hlock0_p & v9739fe | !hlock0_p & !v973a00;
assign v8e799e = hmaster1_p & v8e799a | !hmaster1_p & v8e799d;
assign v9baf71 = stateG10_1_p & v9ed41d | !stateG10_1_p & !v9baf70;
assign v8ea853 = hmaster1_p & v8ea851 | !hmaster1_p & v8ea7f4;
assign v9ed450 = hmaster1_p & v9ed44f | !hmaster1_p & !v86292d;
assign v9baf7d = hmaster1_p & v84563c | !hmaster1_p & v9baf7c;
assign v985512 = hbusreq0 & v98550d | !hbusreq0 & v985511;
assign v9739b4 = hmaster1_p & v9739b3 | !hmaster1_p & !v97397b;
assign v97399f = hmaster0_p & v9738ca | !hmaster0_p & v97395c;
assign v985535 = stateA1_p & v84563c | !stateA1_p & !v9a6a95;
assign v996562 = stateG10_1_p & v9adbee | !stateG10_1_p & !v8ea7e9;
assign v8ea85c = hgrant1_p & v84563c | !hgrant1_p & v8ea7fc;
assign v9855d3 = hbusreq0_p & v9855d2 | !hbusreq0_p & v845641;
assign v973a20 = hgrant2_p & v9739fd | !hgrant2_p & v973a1f;
assign v9a6ad3 = decide_p & v84563c | !decide_p & v9a6a9a;
assign jx2 = !v9d44c5;
assign v8e79b1 = hgrant1_p & v84563c | !hgrant1_p & v8e7993;
assign v99656a = hmaster1_p & v9adbfe | !hmaster1_p & v996569;
assign a153c5 = hmaster1_p & a153c3 | !hmaster1_p & a153c4;
assign v984f40 = hmaster0_p & v984e5a | !hmaster0_p & v984e56;
assign v984f3f = hmaster0_p & v984e54 | !hmaster0_p & v84563c;
assign v9ed4cb = hmaster0_p & v9ed43c | !hmaster0_p & !v9ed49e;
assign v9adce9 = hgrant0_p & v9adcd6 | !hgrant0_p & v9adce8;
assign v8ea7ea = hmastlock_p & v84566e | !hmastlock_p & !v84563c;
assign v984ec1 = hmaster0_p & v84565c | !hmaster0_p & !v984e6f;
assign v9738c7 = hmaster1_p & v9738b0 | !hmaster1_p & v9738c6;
assign v996553 = hbusreq1_p & v9adbf1 | !hbusreq1_p & v996552;
assign v99991f = hbusreq0 & v99991e | !hbusreq0 & !v999912;
assign v985642 = hbusreq1_p & v84565c | !hbusreq1_p & v985520;
assign v9adc7b = hmaster1_p & v9adc78 | !hmaster1_p & v9adc7a;
assign v8e7990 = hburst0_p & v8e7989 | !hburst0_p & v8e798c;
assign v9adc64 = hbusreq1_p & v9adc22 | !hbusreq1_p & !v9adc63;
assign v9adc3e = hmaster1_p & v9adc38 | !hmaster1_p & v9adc3d;
assign v9739e2 = hbusreq0_p & v9739e1 | !hbusreq0_p & v9739bb;
assign v8ea897 = hmaster0_p & v8ea896 | !hmaster0_p & v8ea822;
assign v985563 = stateG2_p & v84563c | !stateG2_p & v985562;
assign v9d2753 = hbusreq0 & v9d2725 | !hbusreq0 & v9d2752;
assign v8ea8df = hmaster1_p & v8ea8de | !hmaster1_p & v8ea7f2;
assign v9855f2 = hbusreq0_p & v9855f0 | !hbusreq0_p & v9855f1;
assign v8c117f = hgrant2_p & v8c116d | !hgrant2_p & v8c117e;
assign v9999a4 = hready_p & v84563c | !hready_p & v9999a3;
assign v9adc66 = hmaster1_p & v9adc65 | !hmaster1_p & v9adc30;
assign v8c20ba = locked_p & v84563c | !locked_p & !v845656;
assign v97394f = hmaster1_p & v9738b0 | !hmaster1_p & v973948;
assign v973941 = hmaster1_p & v97388b | !hmaster1_p & v973940;
assign v9ed4d0 = hmaster1_p & v9ed4cf | !hmaster1_p & !v86292d;
assign v984ec3 = hbusreq0_p & v984ec2 | !hbusreq0_p & v84563c;
assign v9854d8 = hmastlock_p & v8ea7e3 | !hmastlock_p & v84563c;
assign v999918 = hmastlock_p & v999917 | !hmastlock_p & v84563c;
assign v9ed4de = hbusreq0_p & v9ed4dc | !hbusreq0_p & v9ed4dd;
assign v9baf19 = hburst0 & v972fac | !hburst0 & v9baf18;
assign v9adc2f = hmaster1_p & v9adc28 | !hmaster1_p & v9adc2e;
assign v8ea8d1 = hmaster1_p & v8ea823 | !hmaster1_p & v8ea8d0;
assign v984e76 = hgrant0_p & v84563c | !hgrant0_p & v984e75;
assign v8ea93c = jx1_p & v8ea8c7 | !jx1_p & v8ea93b;
assign v999900 = hlock2_p & v9998f6 | !hlock2_p & v9998ff;
assign v9d27ab = hmaster1_p & v9d27aa | !hmaster1_p & !v9d2671;
assign v984f95 = jx0_p & v84563c | !jx0_p & v984f94;
assign v8c1143 = hgrant1_p & v84563c | !hgrant1_p & !v8c1142;
assign v9ed4ba = hmaster0_p & v84563c | !hmaster0_p & !v9ed44e;
assign v9baf8b = hbusreq1 & v9baf82 | !hbusreq1 & v9ed434;
assign v8ea7fd = hmaster0_p & v84563c | !hmaster0_p & v8ea7fc;
assign v9adc8d = hbusreq0_p & v9adc8c | !hbusreq0_p & v9adc89;
assign v8ea8ec = hmaster1_p & v8ea867 | !hmaster1_p & v8ea8d0;
assign v9ed40f = hlock1_p & v9ed40e | !hlock1_p & v84565c;
assign v9999ea = decide_p & v9999e9 | !decide_p & v84565e;
assign v9a6a9e = stateG3_2_p & v84563c | !stateG3_2_p & !v9a6a9d;
assign v8ea803 = hgrant1_p & v8ea7fc | !hgrant1_p & v84563c;
assign v9855e8 = hmaster1_p & v9855e6 | !hmaster1_p & v985594;
assign v98560f = hbusreq0 & v9854b9 | !hbusreq0 & v84563c;
assign v9854db = hlock1_p & v9854d9 | !hlock1_p & !v9854da;
assign v996550 = hmaster0_p & v9adbec | !hmaster0_p & !v99654f;
assign v9d278c = hmaster1_p & v9d26e0 | !hmaster1_p & !v9d2673;
assign v97391a = hmaster1_p & v973919 | !hmaster1_p & !v9738d4;
assign v8ea8c3 = decide_p & v8ea7ee | !decide_p & v8ea8c2;
assign v9854c8 = hmaster0_p & v84563c | !hmaster0_p & v9854c7;
assign a14da1 = hlock2_p & v84563c | !hlock2_p & !a14da0;
assign v984f51 = hlock0_p & v984f50 | !hlock0_p & !v84563c;
assign v84564b = hbusreq2 & v84563c | !hbusreq2 & !v84563c;
assign v9999e7 = hbusreq0 & v9999e4 | !hbusreq0 & v9999e6;
assign v9adbe9 = hmastlock_p & v9adbe8 | !hmastlock_p & !v84563c;
assign v9adcd6 = hmaster1_p & v9adcd5 | !hmaster1_p & v9adc9e;
assign hgrant2 = v9bafa1;
assign v9d27c5 = jx2_p & v9d27c1 | !jx2_p & v9d27c4;
assign v996580 = hmaster1_p & v9adc1a | !hmaster1_p & v99657f;
assign v8ea7f8 = hready_p & v8ea7e8 | !hready_p & v8ea7f7;
assign v8ea87e = decide_p & v8ea7ee | !decide_p & v8ea87d;
assign a2bb5d = stateA1_p & v84563c | !stateA1_p & v84566e;
assign a15508 = hbusreq1_p & a15500 | !hbusreq1_p & a15507;
assign v9d2747 = hready_p & v9d273e | !hready_p & !v9d2746;
assign v985609 = hmaster0_p & v84563c | !hmaster0_p & v985608;
assign v9a6ab1 = locked_p & v9a6aa2 | !locked_p & v84563c;
assign v9adc44 = hmaster1_p & v9adc42 | !hmaster1_p & v9adc43;
assign v9854af = hbusreq1_p & v9854ae | !hbusreq1_p & v84563c;
assign v985612 = hburst1_p & v9854bc | !hburst1_p & !v84563c;
assign a15409 = hlock0_p & a153ec | !hlock0_p & a15408;
assign v99999f = hmaster1_p & v84563c | !hmaster1_p & v9baeaf;
assign v9adc12 = locked_p & v9adbed | !locked_p & v8ea7ea;
assign a2bd45 = stateA1_p & v84563c | !stateA1_p & a2bd3d;
assign v9baef4 = hlock2_p & v9baef3 | !hlock2_p & !v84563c;
assign v9739f8 = hbusreq0_p & v973950 | !hbusreq0_p & v9739f7;
assign v9baf2d = hburst1 & v9baf29 | !hburst1 & v9baf2c;
assign v985613 = hburst0_p & a3134e | !hburst0_p & v985612;
assign v8ea80d = hgrant0_p & v8ea7f9 | !hgrant0_p & v8ea80c;
assign v8ea8a6 = hbusreq0_p & v8ea8a3 | !hbusreq0_p & v8ea8a5;
assign v985583 = hmaster0_p & v84563c | !hmaster0_p & v985582;
assign v9d2767 = hmaster1_p & v9d2764 | !hmaster1_p & !v9d2673;
assign a153bb = hburst0_p & v8e7989 | !hburst0_p & v8e798b;
assign v9baf5e = hgrant1_p & v9baf5d | !hgrant1_p & v9ed419;
assign v9baf99 = hlock2_p & v9baf81 | !hlock2_p & v9baf98;
assign v9d2760 = hgrant0_p & v9d271b | !hgrant0_p & v9d275f;
assign v9bae88 = hmaster1_p & v9bae87 | !hmaster1_p & v9ed438;
assign v8c1164 = hmaster1_p & v8c114d | !hmaster1_p & v84563c;
assign v996559 = hbusreq1_p & v9adbee | !hbusreq1_p & v996552;
assign v973a3e = hbusreq0_p & v9739aa | !hbusreq0_p & v973a3d;
assign a154fd = hbusreq1_p & a154fc | !hbusreq1_p & !a154fb;
assign v98556a = hready & v985565 | !hready & v985569;
assign v8c20b9 = decide_p & v8c20b8 | !decide_p & v84565c;
assign v9adc08 = hbusreq0_p & v9adc07 | !hbusreq0_p & v9adc06;
assign v9933d9 = decide_p & v9933d8 | !decide_p & v9933ce;
assign v97393a = hbusreq0_p & v973891 | !hbusreq0_p & v973939;
assign v8ea87b = hmaster0_p & v84563c | !hmaster0_p & v8ea7e9;
assign v9baf4e = hburst0 & v9baf4c | !hburst0 & v9baf4d;
assign v9ed4ee = decide_p & v9ed4e3 | !decide_p & !v9ed4c6;
assign v9d26e9 = hbusreq0_p & v9d267c | !hbusreq0_p & !v9d26e8;
assign v9d2722 = hgrant0_p & v9d271c | !hgrant0_p & v9d2721;
assign v9d278f = hmaster1_p & v9d26e2 | !hmaster1_p & !v9d2673;
assign v9738fb = decide_p & v9738b6 | !decide_p & v9738fa;
assign v9adc6c = hbusreq0_p & v9adc6a | !hbusreq0_p & v9adc6b;
assign v9738be = hmaster0_p & v97388f | !hmaster0_p & !v97388a;
assign v9738d4 = hmaster0_p & v9738d3 | !hmaster0_p & !v9738cc;
assign v9ed4da = hbusreq0 & v9ed4d6 | !hbusreq0 & v9ed4d9;
assign v8c1170 = hburst1_p & v84563c | !hburst1_p & v8c116f;
assign v8ea7e8 = hmaster1_p & v8ea7e7 | !hmaster1_p & v84563c;
assign v9d26c0 = hbusreq1_p & v9d266f | !hbusreq1_p & v84563c;
assign v9933c1 = stateG10_1_p & v9933b7 | !stateG10_1_p & !v9933c0;
assign v9adce2 = hmaster1_p & v9adce1 | !hmaster1_p & !v9adcb0;
assign v9baf4c = busreq_p & v9ed4a2 | !busreq_p & v9baf4b;
assign v9855ff = hmaster1_p & v9855fe | !hmaster1_p & v84563c;
assign v973a1b = hmaster1_p & v9738f6 | !hmaster1_p & v973a13;
assign v9999aa = hgrant2_p & v9999a4 | !hgrant2_p & !v9999a9;
assign v9adc50 = decide_p & v9adc0e | !decide_p & v9adc4f;
assign v9738a9 = hmaster1_p & v9738a5 | !hmaster1_p & v9738a8;
assign v98552a = hbusreq1_p & v985520 | !hbusreq1_p & v84563c;
assign v9ed49c = locked_p & v9ed475 | !locked_p & v97388d;
assign v9998e9 = hbusreq0 & v9998e8 | !hbusreq0 & v84563c;
assign v9b40dd = jx0_p & v9b40cd | !jx0_p & v9b40dc;
assign v9d272d = decide_p & v9d26f2 | !decide_p & v9d272c;
assign v8e79a1 = hlock0_p & v8e799e | !hlock0_p & v8e79a0;
assign v9d279a = hbusreq0 & v9d2798 | !hbusreq0 & !v9d2799;
assign v9738f3 = hmaster1_p & v9738f2 | !hmaster1_p & !v9738be;
assign v9adccb = decide_p & v9adc92 | !decide_p & v9adcca;
assign v9ed48d = hmaster0_p & v9ed469 | !hmaster0_p & !v9ed482;
assign v9999e5 = hmaster1_p & a154a3 | !hmaster1_p & v9baea4;
assign v8ea81e = hmaster1_p & v8ea815 | !hmaster1_p & v8ea81d;
assign v9854b4 = hmaster0_p & v845641 | !hmaster0_p & v9854b3;
assign v973982 = decide_p & v973953 | !decide_p & v973981;
assign v984eae = hmaster1_p & v984ea8 | !hmaster1_p & v984ead;
assign a154d1 = hmastlock_p & a154c3 | !hmastlock_p & v84563c;
assign v999985 = hbusreq0_p & v999933 | !hbusreq0_p & v84563c;
assign v984f7c = hbusreq0_p & v984f78 | !hbusreq0_p & v984f7b;
assign v8c20c6 = hgrant0_p & v8c20c0 | !hgrant0_p & v8c20c5;
assign v9738e5 = hgrant1_p & v9738dc | !hgrant1_p & v97388d;
assign v9d27ac = hgrant0_p & v9d267b | !hgrant0_p & v9d27ab;
assign v9ecda5 = hgrant2_p & v9ed568 | !hgrant2_p & v9ecda4;
assign v8ea879 = hgrant2_p & v8ea85b | !hgrant2_p & v8ea878;
assign v845648 = hlock1_p & v84563c | !hlock1_p & !v84563c;
assign start = v9933dc;
assign v8ea90c = hmaster0_p & v8ea90b | !hmaster0_p & v8ea822;
assign v9bae8b = decide_p & v9bae8a | !decide_p & v84563c;
assign v99997a = hbusreq0_p & v999979 | !hbusreq0_p & !a14d40;
assign v973a19 = hbusreq0_p & v97397c | !hbusreq0_p & v973a18;
assign a14d49 = decide_p & a14d42 | !decide_p & v84565c;
assign v996568 = hlock0_p & v996565 | !hlock0_p & v996567;
assign v973931 = hmaster1_p & v97392f | !hmaster1_p & v9738ed;
assign v9d2739 = hbusreq0_p & v9d26fd | !hbusreq0_p & v9d2738;
assign v9ed495 = hbusreq2 & v9ed48c | !hbusreq2 & v9ed494;
assign v973891 = hmaster1_p & v97388b | !hmaster1_p & v973890;
assign v973985 = hmaster0_p & v973885 | !hmaster0_p & !v9738c4;
assign v9d2762 = hgrant0_p & v9d2750 | !hgrant0_p & v9d2761;
assign v8ec3e4 = stateG2_p & v84563c | !stateG2_p & !v8543f4;
assign v9ed481 = hmastlock_p & v9ed480 | !hmastlock_p & !v84563c;
assign v9739c4 = hbusreq0_p & v9738ac | !hbusreq0_p & v97394c;
assign v9adc33 = hgrant0_p & v9adc1e | !hgrant0_p & v9adc32;
assign v9b40c4 = hmaster0_p & v9ed4c5 | !hmaster0_p & v845660;
assign v98554c = busreq_p & v9ed4a2 | !busreq_p & v98554b;
assign v8ea908 = hbusreq1_p & v8ea906 | !hbusreq1_p & v8ea907;
assign v984f3b = hready_p & v84563c | !hready_p & v984f3a;
assign v99655b = hmaster1_p & v9adbfa | !hmaster1_p & v99655a;
assign v9999f0 = jx0_p & v9999b6 | !jx0_p & v9999ef;
assign v8ea92c = hmaster1_p & v8ea823 | !hmaster1_p & v8ea91a;
assign v973952 = hbusreq0_p & v973950 | !hbusreq0_p & v973951;
assign v973961 = hgrant1_p & v9738dc | !hgrant1_p & v973893;
assign v9ed4d3 = hmaster0_p & v9ed469 | !hmaster0_p & v9ed477;
assign v9d2732 = hbusreq0 & v9d2730 | !hbusreq0 & v9d267c;
assign v8c115c = stateG10_1_p & v8c1120 | !stateG10_1_p & v8c115b;
assign v9d26ba = hgrant0_p & v9d267f | !hgrant0_p & v9d26b9;
assign v9d26e2 = hmaster0_p & v9d266d | !hmaster0_p & !v84563c;
assign v9d2721 = hbusreq0_p & v9d2720 | !hbusreq0_p & v9d267b;
assign v9baf0f = stateG10_1_p & v9baf0d | !stateG10_1_p & v9baf0e;
assign v9854ed = stateA1_p & v8ea7e3 | !stateA1_p & v9854ea;
assign v9adced = hmaster0_p & v9adc75 | !hmaster0_p & !v9adcc6;
assign v9adcb7 = hgrant1_p & v9adc77 | !hgrant1_p & v9adc75;
assign v9965c9 = hmaster0_p & v9adc48 | !hmaster0_p & v8ea82c;
assign v9adc2a = hgrant1_p & v9adbf9 | !hgrant1_p & v9adbee;
assign v999987 = hmaster1_p & v999986 | !hmaster1_p & v999936;
assign v9adcac = stateG10_1_p & v84563c | !stateG10_1_p & !v9adcab;
assign v9738b3 = hlock0_p & v9738b1 | !hlock0_p & v9738b2;
assign v984f43 = hmastlock_p & v985494 | !hmastlock_p & v84563c;
assign v98549e = hmastlock_p & v9ed42c | !hmastlock_p & v84563c;
assign v9933cc = hmaster0_p & v9933cb | !hmaster0_p & !v84563c;
assign v984ee1 = hbusreq2_p & v984ec0 | !hbusreq2_p & v984ee0;
assign v973a1f = hready_p & v973a17 | !hready_p & !v973a1e;
assign v984ee8 = hmaster1_p & v984ee3 | !hmaster1_p & v984ee7;
assign v9adc40 = hgrant0_p & v9adc19 | !hgrant0_p & v9adc3f;
assign v9ed522 = hgrant2_p & v9ed4fa | !hgrant2_p & v9ed521;
assign v9ed459 = stateG2_p & v84563c | !stateG2_p & v9ed458;
assign v9d2778 = hmaster1_p & v9d2775 | !hmaster1_p & v9d2673;
assign v972fac = hburst0_p & v863b4b | !hburst0_p & v96ef3e;
assign v9738b2 = hmaster1_p & v9738b0 | !hmaster1_p & v9738aa;
assign a154ee = hmaster0_p & a154d1 | !hmaster0_p & v84563c;
assign v8ea8af = hlock2 & v8ea8a9 | !hlock2 & v8ea8ae;
assign v8c20ce = hmaster0_p & v845656 | !hmaster0_p & !v8c20cd;
assign v9adbfb = hmaster1_p & v9adbfa | !hmaster1_p & v9adbee;
assign v973a2a = hbusreq0_p & v973990 | !hbusreq0_p & v973a29;
assign v9d268c = hready & v9d268b | !hready & !v84563c;
assign v9d2697 = hmaster0_p & v9d2690 | !hmaster0_p & v9d2696;
assign v984e5a = hbusreq1_p & v984e59 | !hbusreq1_p & v9855af;
assign v9d273d = hbusreq0 & v9d273a | !hbusreq0 & !v9d273c;
assign v984e6b = stateA1_p & v985561 | !stateA1_p & v985613;
assign v9965c7 = hmaster0_p & v9adc11 | !hmaster0_p & v8ea7f0;
assign stateG3_1 = !v8e79db;
assign v97389d = hmaster1_p & v97389a | !hmaster1_p & v97389c;
assign v9d2677 = hmaster1_p & v9d2676 | !hmaster1_p & !v9d2671;
assign v9d26ab = hmastlock_p & v9d26aa | !hmastlock_p & !v84563c;
assign v9d277c = decide_p & v9d277b | !decide_p & !v9d2754;
assign v845656 = hmastlock_p & v84563c | !hmastlock_p & !v84563c;
assign v8c111f = busreq_p & v8c1118 | !busreq_p & !v92337e;
assign v9a6ad8 = decide_p & v9a6ad7 | !decide_p & v9a6ab3;
assign v9ed4c4 = hbusreq0 & v9ed4b7 | !hbusreq0 & v9ed4c3;
assign v8ea847 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea81c;
assign v9999c6 = hbusreq1_p & v9999bf | !hbusreq1_p & v9999c5;
assign v9999d7 = decide_p & v9999d6 | !decide_p & v84563c;
assign v9854f3 = hburst0_p & v8ea7e2 | !hburst0_p & v9854f2;
assign v9ed47e = stateG2_p & v84563c | !stateG2_p & !v9ed47d;
assign v9baeac = decide_p & v9baeab | !decide_p & v84563c;
assign v973904 = hmaster1_p & v973902 | !hmaster1_p & v973896;
assign v9d26b2 = hgrant0_p & v9d267b | !hgrant0_p & v9d26b1;
assign v9d27b9 = hready_p & v84564b | !hready_p & v9d27b8;
assign v973a24 = hmaster1_p & v973a22 | !hmaster1_p & v9739ee;
assign v984eb2 = stateG10_1_p & v84563c | !stateG10_1_p & !v84565c;
assign v99659f = hmaster0_p & v99659c | !hmaster0_p & v8ea82c;
assign v9965cd = hgrant0_p & v9965c8 | !hgrant0_p & v9965cc;
assign v8c115e = hmaster0_p & v8c115d | !hmaster0_p & !v84563c;
assign v9739a7 = stateG10_1_p & v973893 | !stateG10_1_p & v9738d6;
assign v97391d = stateG10_1_p & v97391b | !stateG10_1_p & v97391c;
assign v8c1158 = hmaster1_p & v8c1157 | !hmaster1_p & !v8c111b;
assign v9d2685 = hburst0 & v845668 | !hburst0 & v9d2684;
assign v9ed50b = decide_p & v9ed501 | !decide_p & v9ed4c6;
assign v985553 = stateA1_p & v8e7990 | !stateA1_p & !v84563c;
assign v973896 = hmaster0_p & v97388f | !hmaster0_p & v973895;
assign v9ed449 = hbusreq0_p & v9ed444 | !hbusreq0_p & v9ed448;
assign v984e73 = hmaster0_p & v984e72 | !hmaster0_p & v84563c;
assign v9a6ab8 = hbusreq0_p & v9a6ab7 | !hbusreq0_p & v84563c;
assign v8ea8d8 = hbusreq0 & v8ea8d5 | !hbusreq0 & v8ea8d7;
assign v9933ca = stateG10_1_p & v84563c | !stateG10_1_p & !v9933c4;
assign v9adcda = hbusreq0_p & v9adcd8 | !hbusreq0_p & !v9adcd9;
assign v8c20da = hmaster0_p & v8c20d9 | !hmaster0_p & v8c20d5;
assign v8ea8bd = hbusreq0_p & v8ea8bc | !hbusreq0_p & v8ea869;
assign v985634 = hmaster0_p & v84563c | !hmaster0_p & v9854da;
assign v9855b6 = hmaster1_p & v9855b1 | !hmaster1_p & v9855b5;
assign v9855a2 = hmaster0_p & v84563c | !hmaster0_p & !v9855a1;
assign v9933da = hready_p & v9933d9 | !hready_p & !v84563c;
assign v985503 = hmaster1_p & v985501 | !hmaster1_p & v985502;
assign v9854da = hready & v8ea7e2 | !hready & !v9ed456;
assign v9adc86 = stateG10_1_p & v84563c | !stateG10_1_p & !v9adc75;
assign v8ea819 = hready & v8ea818 | !hready & v8ea7e9;
assign v99989d = hlock0_p & v99989c | !hlock0_p & v84563c;
assign v973a40 = decide_p & v973a3a | !decide_p & v973a3f;
assign v985521 = hbusreq1_p & v985520 | !hbusreq1_p & v845641;
assign v9854e6 = hmaster1_p & v9854e4 | !hmaster1_p & v9854b8;
assign v9adc79 = hbusreq1_p & v84563c | !hbusreq1_p & !v9adc75;
assign v9f356c = hmaster1_p & v9f3568 | !hmaster1_p & v9f356b;
assign v9d276f = hmaster0_p & v9d276e | !hmaster0_p & v84563c;
assign v999924 = hmaster0_p & v9baf2f | !hmaster0_p & v84563c;
assign v8c1159 = hmaster1_p & v8c1157 | !hmaster1_p & !v8c114d;
assign v984ef2 = hmaster0_p & v985627 | !hmaster0_p & v984ef1;
assign v9adcc2 = hmaster1_p & v9adc7f | !hmaster1_p & !v9adcc1;
assign v8ea83c = hbusreq0_p & v8ea817 | !hbusreq0_p & v8ea83b;
assign v99658d = hgrant1_p & v99654f | !hgrant1_p & !v996552;
assign v9738a3 = decide_p & v9738a2 | !decide_p & v973898;
assign v8c113e = hready_p & v8c111e | !hready_p & !v8c113d;
assign v9d26a7 = stateG2_p & v84563c | !stateG2_p & !v9d26a6;
assign v8c1177 = hbusreq1_p & v8c1143 | !hbusreq1_p & v8c1176;
assign v98557a = hgrant1_p & v84563c | !hgrant1_p & !v985579;
assign v9adc16 = hready_p & v9adbfd | !hready_p & !v9adc15;
assign v9baf01 = busreq_p & v9baf00 | !busreq_p & !v84563c;
assign v973993 = hbusreq0_p & v973990 | !hbusreq0_p & v973992;
assign a14da9 = hmaster0_p & a154fd | !hmaster0_p & v84563c;
assign v973a06 = stateG10_1_p & v97388d | !stateG10_1_p & v973a05;
assign v985490 = hlock1_p & v98548f | !hlock1_p & v84563c;
assign v8ea8ef = hgrant0_p & v8ea8eb | !hgrant0_p & v8ea8ee;
assign v8ea8f5 = decide_p & v8ea7ee | !decide_p & v8ea8f4;
assign v8c114a = hgrant0_p & v8c1141 | !hgrant0_p & v8c1149;
assign v8ea867 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea82c;
assign v984edc = hbusreq0 & v984eda | !hbusreq0 & v984ebb;
assign v9739f1 = hlock2_p & v9739ea | !hlock2_p & !v9739f0;
assign v9d2668 = hbusreq1 & v9d2667 | !hbusreq1 & v84563c;
assign v9999a7 = decide_p & v9999a6 | !decide_p & v84565e;
assign v8ea8b4 = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea7f0;
assign v9baf10 = hbusreq1_p & v9baf06 | !hbusreq1_p & !v9baf0f;
assign v9933c6 = hbusreq1_p & v9933c5 | !hbusreq1_p & !v8c20d8;
assign v9854ca = hmaster1_p & v9854c6 | !hmaster1_p & v9ed438;
assign v9ed486 = hburst0 & v84563c | !hburst0 & v9ed485;
assign v9ed464 = busreq_p & v9ed463 | !busreq_p & !a2bd45;
assign v984f84 = hbusreq0_p & v984f82 | !hbusreq0_p & v984f7b;
assign v9d270a = hbusreq0 & v9d2708 | !hbusreq0 & !v9d2709;
assign v9ed46e = hbusreq1_p & v9ed46d | !hbusreq1_p & v84563c;
assign v9999dc = hgrant0_p & v9999db | !hgrant0_p & !v84563c;
assign v9adc59 = hready_p & v9adc53 | !hready_p & !v9adc58;
assign v9ed43e = hburst0 & v86cfb3 | !hburst0 & v9ed43d;
assign v973926 = hmaster1_p & v973925 | !hmaster1_p & !v9738e8;
assign a14dad = hgrant0_p & a14da8 | !hgrant0_p & a14dab;
assign v9ed422 = hbusreq0_p & v9ed41c | !hbusreq0_p & v9ed421;
assign v9739ad = hbusreq0_p & v9739aa | !hbusreq0_p & v9739ac;
assign v9854c3 = locked_p & v9854c2 | !locked_p & !v84563c;
assign v8c20d6 = hmaster0_p & v8c20c3 | !hmaster0_p & v8c20d5;
assign a14d71 = hready_p & a14d70 | !hready_p & a14d68;
assign v9855b2 = hmaster1_p & v9855b1 | !hmaster1_p & v985583;
assign v9855a8 = stateA1_p & a153cb | !stateA1_p & !v84563c;
assign v9d26b4 = hgrant0_p & v9d267c | !hgrant0_p & v9d26b3;
assign v9ed44a = hburst1 & v84563c | !hburst1 & v86cfb3;
assign v9adbe7 = stateG2_p & v84563c | !stateG2_p & !a2bb5d;
assign v999979 = hlock0_p & v999978 | !hlock0_p & v999925;
assign v9a6aac = hmaster1_p & v9a6aab | !hmaster1_p & v9a6aa5;
assign v9739d0 = hready_p & v9739cc | !hready_p & !v9739cf;
assign v9adc61 = locked_p & v9adc60 | !locked_p & !v9adbeb;
assign v98563f = hbusreq0 & v98563e | !hbusreq0 & v84563c;
assign v985620 = stateA1_p & v84563c | !stateA1_p & v8ea7fa;
assign v9998ae = hbusreq0 & v9998a8 | !hbusreq0 & v9998ad;
assign v8ea7ef = locked_p & v84563c | !locked_p & !v8ea7ea;
assign v9baef9 = hready_p & v9baef5 | !hready_p & !v9baef8;
assign v8ea835 = hmaster1_p & v8ea815 | !hmaster1_p & v8ea834;
assign v9baeaf = hmaster0_p & v84563c | !hmaster0_p & !v845656;
assign a15416 = hbusreq0_p & a15415 | !hbusreq0_p & v845648;
assign v9adcc3 = hmaster1_p & v9adc7f | !hmaster1_p & v9adcba;
assign v985544 = hburst0_p & a3134f | !hburst0_p & v985543;
assign v9adc70 = hready_p & v9adc6e | !hready_p & !v9adc6f;
assign v9baf90 = hmaster1_p & v9baf8a | !hmaster1_p & v9baf8f;
assign v9855f5 = hbusreq2 & v9855ee | !hbusreq2 & v9855f4;
assign v98558d = locked_p & v98558c | !locked_p & v84563c;
assign v8ea87d = hbusreq0_p & v8ea87c | !hbusreq0_p & v8ea7f5;
assign v9d26bd = decide_p & v9d267a | !decide_p & v9d26bc;
assign v9999db = hbusreq0_p & v9999da | !hbusreq0_p & !v84563c;
assign v9999f1 = jx1_p & v99999e | !jx1_p & v9999f0;
assign v9965c5 = hgrant0_p & v9965b5 | !hgrant0_p & v9965c4;
assign a15434 = hmaster0_p & v84563c | !hmaster0_p & !a15433;
assign v9d26a3 = decide_p & v9d269c | !decide_p & v9d26a2;
assign v8ea8f1 = hlock0 & v8ea8f0 | !hlock0 & v8ea8ef;
assign v9adc55 = hmaster0_p & v9adc54 | !hmaster0_p & !v8ea7ea;
assign v99990d = hmaster0_p & v9baf2f | !hmaster0_p & !v9baf30;
assign v9d44c4 = jx0_p & v84563c | !jx0_p & !v9d44c3;
assign v984eda = hgrant0_p & v984ea4 | !hgrant0_p & v984ed9;
assign v9d2792 = hlock2_p & v9d278e | !hlock2_p & v9d2791;
assign v8e7994 = hmaster0_p & v84563c | !hmaster0_p & v8e7993;
assign a154bb = hlock2_p & a154a6 | !hlock2_p & v845644;
assign v9854aa = hmastlock_p & v9bae7b | !hmastlock_p & v84563c;
assign v9999c5 = stateG10_1_p & v9999bf | !stateG10_1_p & v9999c4;
assign v9baf96 = hgrant0_p & v9baf95 | !hgrant0_p & v9baf90;
assign v973919 = hmaster0_p & v9738ca | !hmaster0_p & v9738d7;
assign v8ea8ad = hlock0 & v8ea8a7 | !hlock0 & v8ea8ac;
assign v9965b5 = hmaster1_p & v9965b4 | !hmaster1_p & v996579;
assign v999935 = hmaster0_p & v9baf55 | !hmaster0_p & v9baf69;
assign v9baeb2 = hmaster0_p & v84563c | !hmaster0_p & v9bae92;
assign v984ee7 = hmaster0_p & v985627 | !hmaster0_p & v845641;
assign v985593 = hbusreq1_p & v985592 | !hbusreq1_p & !v84563c;
assign v9738c4 = locked_p & v87f892 | !locked_p & v97388d;
assign v9999bb = stateA1_p & v972fac | !stateA1_p & a153cb;
assign a1548d = hmaster0_p & v845646 | !hmaster0_p & a15489;
assign v9baf4a = hbusreq1 & v9ed40e | !hbusreq1 & v84565c;
assign v9d26c9 = hbusreq0_p & v9d2677 | !hbusreq0_p & v9d26c8;
assign v8e79b5 = hbusreq1_p & v8e79b4 | !hbusreq1_p & v84563c;
assign v845650 = hburst1_p & v84563c | !hburst1_p & !v84563c;
assign v985530 = hmaster0_p & v985491 | !hmaster0_p & v9854a4;
assign a153d3 = hbusreq1_p & a153d2 | !hbusreq1_p & v84563c;
assign v8c20df = hready_p & v8c20de | !hready_p & v8c20d0;
assign v8e7996 = hlock2_p & v8e7995 | !hlock2_p & v84563c;
assign v9933d7 = hbusreq0_p & v9933c8 | !hbusreq0_p & v9933d6;
assign v99996d = hmaster1_p & v99996c | !hmaster1_p & v9998f8;
assign v984ea9 = hgrant1_p & v985526 | !hgrant1_p & !v84563c;
assign v8ea8a1 = hgrant2_p & v8ea87f | !hgrant2_p & v8ea8a0;
assign v985572 = busreq_p & v98556f | !busreq_p & v985571;
assign v8ea8dc = hready_p & v8ea80e | !hready_p & v8ea8db;
assign a14da6 = hmaster1_p & a154a3 | !hmaster1_p & a154a2;
assign v98563a = hmaster0_p & v985624 | !hmaster0_p & v845641;
assign v9855d5 = hmaster1_p & v84563c | !hmaster1_p & v845641;
assign v9baf78 = hmaster1_p & a154a3 | !hmaster1_p & v9baf77;
assign v973a34 = hbusreq0_p & v973a32 | !hbusreq0_p & !v973a33;
assign v984eba = hmaster1_p & v984eb9 | !hmaster1_p & v84563c;
assign v985498 = hready & v985497 | !hready & a153c0;
assign v8ea858 = hlock2 & v8ea84e | !hlock2 & v8ea856;
assign v9933ba = hlock2_p & v9933b9 | !hlock2_p & v8c20b7;
assign v9998a5 = hmaster1_p & v84565c | !hmaster1_p & v9bae79;
assign v9adcf1 = hgrant0_p & v9adcec | !hgrant0_p & v9adcf0;
assign v8ea932 = hmaster1_p & v8ea867 | !hmaster1_p & v8ea918;
assign a153ca = hburst1_p & v96ef3e | !hburst1_p & v863b4b;
assign v9855e1 = hmaster1_p & v9855e0 | !hmaster1_p & v98557f;
assign v9d2701 = hmaster0_p & v9d2700 | !hmaster0_p & v845647;
assign v8e799a = hmastlock_p & v8e7999 | !hmastlock_p & v84563c;
assign a14dc2 = jx1_p & a14d5b | !jx1_p & a14dc1;
assign v9d26a5 = hburst0_p & v84563c | !hburst0_p & v8c1130;
assign v985557 = hlock1_p & v98554f | !hlock1_p & v985556;
assign v9854b1 = hmaster1_p & v9854b0 | !hmaster1_p & v84563c;
assign v8ea84b = hmaster0_p & v8ea7e9 | !hmaster0_p & v8ea839;
assign v9adc5a = hmaster0_p & v9adbec | !hmaster0_p & v9adbee;
assign stateG10_1 = !v9f357b;
assign v973a14 = hmaster1_p & v9738e4 | !hmaster1_p & !v973a13;
assign v9ed494 = hbusreq0 & v9ed490 | !hbusreq0 & v9ed493;
assign v996591 = hmaster1_p & v9adc38 | !hmaster1_p & !v996590;
assign v985549 = locked_p & v985548 | !locked_p & v84563c;
assign v9baefc = hgrant2_p & v9baef9 | !hgrant2_p & !v9baefb;
assign v984f45 = hready & v984f44 | !hready & v9854aa;
assign v8e799b = hlock1_p & v8e799a | !hlock1_p & v84563c;
assign v984f62 = hmaster0_p & v984f5f | !hmaster0_p & v984eb3;
assign v996584 = hgrant1_p & v99657e | !hgrant1_p & !v996552;
assign v9baf7f = hgrant0_p & v9baf7e | !hgrant0_p & v9baf75;
assign v9adc4f = hgrant0_p & v9adc44 | !hgrant0_p & v9adc4e;
assign v9d2674 = hmaster1_p & v9d2670 | !hmaster1_p & !v9d2673;
assign v9baf28 = stateG2_p & v84563c | !stateG2_p & !v9baf27;
assign v996565 = hmaster1_p & v9adbfe | !hmaster1_p & v996564;
assign v9adc24 = hbusreq1_p & v9adc22 | !hbusreq1_p & !v9adc23;
assign v9d27b0 = hbusreq2 & v9d27af | !hbusreq2 & v9d2680;
assign v984ef4 = hlock0_p & v984ef3 | !hlock0_p & v984ee8;
assign v984e5f = hlock1_p & v9855fd | !hlock1_p & !v84563c;
assign v9739ae = hgrant0_p & v9739a6 | !hgrant0_p & v9739ad;
assign v9ed490 = hbusreq0_p & v9ed48e | !hbusreq0_p & v9ed48f;
assign v8c1148 = hmaster0_p & v8c1147 | !hmaster0_p & !v84563c;
assign v9854a5 = hmaster0_p & v84563c | !hmaster0_p & v9854a4;
assign v9adc07 = hlock0_p & v9adc04 | !hlock0_p & v9adc06;
assign v9d2765 = hmaster1_p & v9d2764 | !hmaster1_p & !v9d2671;
assign v985529 = hmaster1_p & v985528 | !hmaster1_p & v9ed438;
assign a14d5a = hbusreq2_p & a14d3d | !hbusreq2_p & a14d59;
assign v9ed4d7 = hmaster1_p & v9ed4d3 | !hmaster1_p & v9ed483;
assign v9baea1 = hbusreq2_p & v9bae9f | !hbusreq2_p & !v9baea0;
assign v9738cf = hgrant1_p & v973899 | !hgrant1_p & v973889;
assign v9998cf = hgrant2_p & v9998a4 | !hgrant2_p & !v9998ce;
assign v9ed46d = hmastlock_p & v9ed46c | !hmastlock_p & v845666;
assign v84565a = decide_p & v84563c | !decide_p & !v84563c;
assign v9baf20 = hmaster0_p & v9baf10 | !hmaster0_p & !v9baf1f;
assign v9adc00 = hlock1_p & v9adbed | !hlock1_p & v8ea7ea;
assign a1550a = hmaster1_p & a154fe | !hmaster1_p & a15509;
assign v9965ae = hlock0_p & v9965ac | !hlock0_p & v9965ad;
assign v9baea8 = hbusreq0_p & v9baea5 | !hbusreq0_p & v84563c;
assign v984e75 = hbusreq0_p & v984e74 | !hbusreq0_p & v84563c;
assign v9998d3 = decide_p & a14d6e | !decide_p & v84563c;
assign v9f3568 = hbusreq1_p & v84563c | !hbusreq1_p & v845660;
assign v985518 = hmaster0_p & v9854fb | !hmaster0_p & v9854b3;
assign v99992e = hbusreq0 & v99992d | !hbusreq0 & !v999912;
assign v9d26d5 = hbusreq0_p & v9d2699 | !hbusreq0_p & v9d26d4;
assign v9adc15 = decide_p & v9adc0e | !decide_p & v9adc14;
assign v8ea8a3 = hmaster1_p & v8ea8a2 | !hmaster1_p & v8ea7f2;
assign v9d2706 = hmaster1_p & v9d26fa | !hmaster1_p & v9d26fc;
assign v8ea86f = hlock0 & v8ea86b | !hlock0 & v8ea86e;
assign v9d272b = hbusreq0 & v9d272a | !hbusreq0 & v9d267f;
assign v9baf45 = hmaster1_p & v9baf42 | !hmaster1_p & v9baf44;
assign v9baf9d = hgrant2_p & v9baf41 | !hgrant2_p & !v9baf9c;
assign v8ea877 = decide_p & v8ea7ee | !decide_p & v8ea876;
assign v9ed41f = hbusreq1_p & v9ed41e | !hbusreq1_p & v84563c;
assign v9998e8 = hbusreq0_p & v9998e7 | !hbusreq0_p & v84563c;
assign v9998e5 = hmaster1_p & v9998e3 | !hmaster1_p & v9998e4;
assign v985566 = stateA1_p & a153bb | !stateA1_p & !v84563c;
assign v9ed41e = hlock1_p & v9ed41d | !hlock1_p & v84565c;
assign v9d2695 = hlock1_p & v9d2693 | !hlock1_p & v9d2694;
assign v98561d = hbusreq0_p & v98561c | !hbusreq0_p & v84563c;
assign v973983 = hready_p & v97396b | !hready_p & !v973982;
assign v9d27a8 = decide_p & v9d27a2 | !decide_p & v9d27a7;
assign v9baef6 = hbusreq2 & v9baeb0 | !hbusreq2 & v85bb54;
assign v985601 = hbusreq0_p & v985600 | !hbusreq0_p & v84563c;
assign v9a6ac7 = hmaster1_p & v84563c | !hmaster1_p & v9a6ab2;
assign v999927 = hbusreq0_p & v999926 | !hbusreq0_p & !v84563c;
assign v9adc0a = hmaster1_p & v9adc09 | !hmaster1_p & !v9adc03;
assign v8ea7e3 = stateG3_2_p & v84563c | !stateG3_2_p & !v8ea7e2;
assign v9ed4ff = hmaster1_p & v9ed4b4 | !hmaster1_p & v9ed4fe;
assign v9a6ae0 = decide_p & v9a6ad7 | !decide_p & v9a6acf;
assign v9855c7 = hmaster1_p & v9855c6 | !hmaster1_p & v9854df;
assign v8c117a = hbusreq0_p & v8c1149 | !hbusreq0_p & v8c1179;
assign v9adcd3 = decide_p & v9adc8d | !decide_p & v9adc9a;
assign v9d26fc = hmaster0_p & v9d26fa | !hmaster0_p & v845647;
assign v8ea821 = stateG10_1_p & v8ea7ea | !stateG10_1_p & !v8ea820;
assign v8e79d1 = hready_p & v8e79cb | !hready_p & v8e79d0;
assign v9baec7 = hbusreq0_p & v9baeb3 | !hbusreq0_p & v85bb54;
assign v9adc0d = hbusreq0_p & v9adc0c | !hbusreq0_p & v9adc0b;
assign a15485 = decide_p & a15484 | !decide_p & v84565c;
assign v984e66 = hbusreq1_p & v8c20d7 | !hbusreq1_p & !v8c20d8;
assign v9adcbf = hgrant0_p & v9adc9f | !hgrant0_p & v9adcbe;
assign v9adc3b = hmaster0_p & v9adc3a | !hmaster0_p & v9adc37;
assign a14d59 = hgrant2_p & a14d4a | !hgrant2_p & a14d58;
assign v8ea8f6 = hready_p & v8ea862 | !hready_p & v8ea8f5;
assign v8ea837 = hgrant0_p & v8ea836 | !hgrant0_p & v8ea82f;
assign v8c1121 = hmaster0_p & v8c1120 | !hmaster0_p & v8c1119;
assign v9f3578 = hready_p & v9f3576 | !hready_p & v9f3577;
assign v9933d4 = hbusreq1_p & v9933c0 | !hbusreq1_p & !a15507;
assign v8ea863 = hmaster0_p & v8ea814 | !hmaster0_p & v8ea7f0;
assign v8e79ca = hgrant2_p & v8e79ad | !hgrant2_p & v8e79c9;
assign v985587 = decide_p & v98555c | !decide_p & v985586;
assign v9739e1 = hmaster1_p & v9739ba | !hmaster1_p & v9738e8;
assign v8ea893 = hgrant0_p & v8ea884 | !hgrant0_p & v8ea892;
assign v9ed4c8 = decide_p & v9ed495 | !decide_p & !v9ed4c6;
assign v9baf3b = hmaster1_p & v9baf2f | !hmaster1_p & !v9baf3a;
assign v9d2705 = hbusreq0 & v9d26ff | !hbusreq0 & !v9d2704;
assign v98564f = hgrant1_p & v98548f | !hgrant1_p & v98564e;
assign v9998ec = hburst1 & v8e7991 | !hburst1 & v9998eb;
assign v984f8a = hready_p & v984f67 | !hready_p & v984f89;
assign v9a6a98 = locked_p & v9a6a97 | !locked_p & v84563c;
assign v98554f = hgrant1_p & v84563c | !hgrant1_p & v98554e;
assign a153c9 = decide_p & a153c8 | !decide_p & v84565c;
assign v9bae84 = hbusreq1 & a153c0 | !hbusreq1 & !v9bae82;
assign v9baf54 = stateG10_1_p & v9baf50 | !stateG10_1_p & !v9baf53;
assign v9855df = hbusreq0_p & v9855dd | !hbusreq0_p & v9855de;
assign v973a00 = hmaster1_p & v9738b0 | !hmaster1_p & v9739ff;
assign v9d2770 = hmaster1_p & v9d276f | !hmaster1_p & v9d2671;
assign v9baecc = hready_p & v9baeac | !hready_p & !v9baecb;
assign v9854e4 = hmaster0_p & v9854cf | !hmaster0_p & v9854dc;
assign v984ee0 = hgrant2_p & v984ecb | !hgrant2_p & v984edf;
assign v9738bd = hmaster0_p & v973886 | !hmaster0_p & v97388c;
assign v9adc5b = hmaster1_p & v9adc5a | !hmaster1_p & v9adc18;
assign v9adc77 = locked_p & v9adc75 | !locked_p & !v84563c;
assign v8ea89d = hlock2 & v8ea89a | !hlock2 & v8ea89c;
assign v984eb8 = hbusreq1_p & v9855ae | !hbusreq1_p & v9855af;
assign v996575 = hmaster1_p & v996573 | !hmaster1_p & v8ea7f4;
assign v9d27b4 = hbusreq0_p & v9d26e5 | !hbusreq0_p & !v9d267b;
assign v9d277d = hready_p & v84564b | !hready_p & v9d277c;
assign v984f92 = hbusreq2_p & v984f8b | !hbusreq2_p & v984f91;
assign v985579 = hready & v985574 | !hready & !v985578;
assign v8ea8d4 = hbusreq0_p & v8ea8d1 | !hbusreq0_p & v8ea8d3;
assign v9adc48 = hbusreq1_p & v9adc46 | !hbusreq1_p & v9adc47;
assign v985648 = decide_p & v985640 | !decide_p & v985647;
assign v9999b0 = hgrant0_p & v999985 | !hgrant0_p & !a14d6e;
assign v9ed466 = hburst0 & v9ed462 | !hburst0 & v9ed465;
assign v984ebd = hbusreq2 & v984eb1 | !hbusreq2 & v984ebc;
assign v99657b = hmaster0_p & v996559 | !hmaster0_p & v9adbf9;
assign v9854a7 = hmaster0_p & v84563c | !hmaster0_p & v985491;
assign v984f5b = hmaster0_p & v984e66 | !hmaster0_p & v84563c;
assign v8c20d2 = hgrant2_p & v8c20bd | !hgrant2_p & v8c20d1;
assign v996577 = decide_p & v996571 | !decide_p & v996576;
assign v9adc57 = hbusreq0_p & v9adc0c | !hbusreq0_p & v9adc56;
assign v9adbfa = hmaster0_p & v9adbeb | !hmaster0_p & v9adbf9;
assign v9ed439 = hmaster1_p & v9ed437 | !hmaster1_p & v9ed438;
assign v984f2e = hbusreq0_p & v984f2d | !hbusreq0_p & v98563c;
assign v97399a = hmaster1_p & v973999 | !hmaster1_p & v9738be;
assign v984eaa = hgrant1_p & v985592 | !hgrant1_p & v84563c;
assign v9ed410 = hbusreq1_p & v9ed40f | !hbusreq1_p & v84563c;
assign v9ed43a = hbusreq2 & v9ed422 | !hbusreq2 & v9ed439;
assign v9ed4c1 = hmaster1_p & v845646 | !hmaster1_p & !v9ed4c0;
assign v9d2787 = decide_p & v9d2786 | !decide_p & v9d275a;
assign v9f356a = hbusreq1_p & v84563c | !hbusreq1_p & !v9f3569;
assign v8ea7fa = stateG3_2_p & v84563c | !stateG3_2_p & !v84566a;
assign v9854b6 = hmaster1_p & v9854b4 | !hmaster1_p & v845641;
assign v8ea873 = hlock0 & v8ea872 | !hlock0 & v8ea86e;
assign v984f3a = decide_p & v984f38 | !decide_p & v984f39;
assign v999911 = hlock0_p & v898b4e | !hlock0_p & v84563c;
assign v9adcaa = hlock1_p & v9adca9 | !hlock1_p & !v84563c;
assign v9ed4e6 = hmaster0_p & v9ed410 | !hmaster0_p & v9ed41f;
assign v9d279c = hbusreq0 & v9d279b | !hbusreq0 & !v9d2709;
assign v973912 = hready_p & v973906 | !hready_p & v973911;
assign v9baf86 = hgrant1_p & v84565c | !hgrant1_p & !v9ed4ac;
assign v99998d = hbusreq0 & v99998a | !hbusreq0 & v99998c;
assign a154a2 = hmaster0_p & v84565c | !hmaster0_p & a153c0;
assign v985628 = hmaster0_p & v985627 | !hmaster0_p & v84563c;
assign v8ea828 = hmaster0_p & v8ea827 | !hmaster0_p & v8ea822;
assign v97393e = hlock2_p & v97393a | !hlock2_p & !v97393d;
assign v8c1123 = hbusreq1_p & v8c1122 | !hbusreq1_p & !v84563c;
assign hmaster0 = !v960f67;
assign v9adcb6 = hmaster0_p & v9adcb5 | !hmaster0_p & v84563c;
assign v9a6a96 = stateG2_p & v84563c | !stateG2_p & v9a6a95;
assign v9baf80 = hbusreq0 & v9baf76 | !hbusreq0 & v9baf7f;
assign v985507 = hbusreq0 & v9854e8 | !hbusreq0 & v985506;
assign v9965aa = decide_p & v9965a9 | !decide_p & v996558;
assign v9adc90 = hlock0_p & v9adc8e | !hlock0_p & v9adc8f;
assign v9738f1 = decide_p & v9738db | !decide_p & v9738f0;
assign v984f56 = hmaster0_p & v98561a | !hmaster0_p & v9854c4;
assign v9739eb = hbusreq1_p & v973889 | !hbusreq1_p & !v973893;
assign v985622 = busreq_p & v8ea7fb | !busreq_p & v985621;
assign v9ed4f8 = hbusreq0_p & v9ed4f5 | !hbusreq0_p & v9ed4f7;
assign v8e79bc = hmaster1_p & v8e79b2 | !hmaster1_p & v8e79bb;
assign a153c2 = hbusreq1_p & a153c1 | !hbusreq1_p & v84563c;
assign v9ed45d = hmastlock_p & v9ed45c | !hmastlock_p & v84563c;
assign v9a6ac0 = hgrant0_p & v9a6ab8 | !hgrant0_p & v9a6abf;
assign v8ea81a = hlock1 & v8ea7e9 | !hlock1 & v8ea819;
assign v9738c0 = hmaster0_p & v97389b | !hmaster0_p & v973899;
assign v9855b0 = hbusreq1_p & v9855ad | !hbusreq1_p & v9855af;
assign v9965ca = hmaster1_p & v9965c9 | !hmaster1_p & v99659d;
assign v999901 = decide_p & v999900 | !decide_p & v84563c;
assign v8c114e = hmaster1_p & v84563c | !hmaster1_p & v8c114d;
assign v9855e4 = hgrant0_p & v9855df | !hgrant0_p & v9855e3;
assign v99993f = hbusreq0 & v99993d | !hbusreq0 & v99993e;
assign v9738fe = hmaster0_p & v973885 | !hmaster0_p & !v9738c5;
assign v8c1118 = stateG2_p & v84563c | !stateG2_p & !v883467;
assign v984ecd = hmaster1_p & v984ecc | !hmaster1_p & v984e73;
assign v9adc74 = hmastlock_p & v9adc73 | !hmastlock_p & v84563c;
assign v8ea926 = hready_p & v8ea846 | !hready_p & v8ea925;
assign v999908 = hburst0 & v999906 | !hburst0 & v999907;
assign v9ed4d2 = decide_p & v9ed4d1 | !decide_p & v84563c;
assign v9738ad = hmaster0_p & v9738a7 | !hmaster0_p & !v97389e;
assign a154d4 = hbusreq1_p & a154d3 | !hbusreq1_p & !v84563c;
assign v984eb7 = hgrant0_p & v984ea4 | !hgrant0_p & v984eb6;
assign v999972 = hlock0_p & v999971 | !hlock0_p & v84563c;
assign v9ed426 = hburst0_p & v84563c | !hburst0_p & v9ed425;
assign v8996a7 = hburst1_p & v84563c | !hburst1_p & v878a51;
assign v9933c3 = hmaster0_p & v9933c2 | !hmaster0_p & v84563c;
assign v9a6aa8 = hmaster1_p & v9a6aa2 | !hmaster1_p & v9a6aa7;
assign v8543f4 = stateG3_2_p & v84563c | !stateG3_2_p & v85a40d;
assign v9baf11 = hmaster0_p & v9baf10 | !hmaster0_p & v9ed46d;
assign v9965a4 = hready_p & v996596 | !hready_p & !v9965a3;
assign v9baeab = hlock2_p & v9baeaa | !hlock2_p & !v84563c;
assign v9adccf = hmaster1_p & v9adcce | !hmaster1_p & !v9adc7a;
assign v8ea7fe = hmaster1_p & v84563c | !hmaster1_p & v8ea7fd;
assign v9739f4 = hmaster0_p & v973945 | !hmaster0_p & !v973893;
assign v973892 = stateG2_p & v84563c | !stateG2_p & v87f892;
assign v98557d = hbusreq1_p & v98557c | !hbusreq1_p & v84563c;
assign v9adbea = busreq_p & a2bb5d | !busreq_p & !v9adbe7;
assign v999974 = hbusreq0 & v999973 | !hbusreq0 & !v845642;
assign v9adc4a = hgrant1_p & v9adc12 | !hgrant1_p & v8ea7ea;
assign v8ea86a = hbusreq0_p & v8ea868 | !hbusreq0_p & v8ea869;
assign v97395d = hmaster0_p & v9738d3 | !hmaster0_p & !v97395c;
assign v985541 = hlock0_p & v98553f | !hlock0_p & v985540;
assign v973a4c = jx1_p & v9739c2 | !jx1_p & v973a4b;
assign v973939 = hmaster1_p & v97388b | !hmaster1_p & v973938;
assign v973945 = hbusreq1_p & v9738a6 | !hbusreq1_p & !v973944;
assign v9738a2 = hlock2_p & v973898 | !hlock2_p & !v9738a1;
assign v9855e6 = hmaster0_p & v985521 | !hmaster0_p & v98552a;
assign stateA1 = !v973a4c;
assign a14d3d = hgrant2_p & a154f5 | !hgrant2_p & a14d3c;
assign v9ed499 = hmaster0_p & v84563c | !hmaster0_p & v9ed417;
assign v9d26c4 = hmaster1_p & v9d26c1 | !hmaster1_p & !v9d2673;
assign v973a0c = hmaster0_p & v973a07 | !hmaster0_p & !v973a0b;
assign v98563c = hmaster1_p & v84563c | !hmaster1_p & !v98562c;
assign v973998 = hready_p & v97398c | !hready_p & v973997;
assign v9998db = hbusreq0_p & v9998ab | !hbusreq0_p & !v854658;
assign v9a6abf = hmaster1_p & v9a6aba | !hmaster1_p & v9a6abe;
assign v8ea89e = hbusreq2 & v8ea89c | !hbusreq2 & v8ea89d;
assign v97398a = hmaster1_p & v973902 | !hmaster1_p & v973938;
assign v9d27be = decide_p & v9d27bd | !decide_p & v9d279c;
assign v985582 = hbusreq1_p & v985581 | !hbusreq1_p & v84563c;
assign v9739b6 = hmaster1_p & v9739b5 | !hmaster1_p & !v9738dd;
assign v97397d = hbusreq0_p & v97397c | !hbusreq0_p & v9738f4;
assign v9ed533 = hgrant2_p & v9ed52e | !hgrant2_p & v9ed532;
assign v8ea904 = hmaster1_p & v8ea880 | !hmaster1_p & v8ea903;
assign v9855bd = hgrant2_p & v98552f | !hgrant2_p & v9855bc;
assign v8ea8e2 = hmaster1_p & v8ea8a4 | !hmaster1_p & v8ea7f2;
assign a2bd3c = hburst1_p & v84563c | !hburst1_p & v85a40d;
assign v9baf42 = hmaster0_p & v9ed40e | !hmaster0_p & v84563c;
assign v9d2748 = hgrant2_p & v9d2735 | !hgrant2_p & v9d2747;
assign v9ed47b = hburst1_p & v84563c | !hburst1_p & !v96ef3e;
assign v9ed4c6 = hgrant0_p & v84563c | !hgrant0_p & !v9ed4c5;
assign a153ec = hmaster1_p & a153eb | !hmaster1_p & a153d5;
assign v9739d5 = hmaster1_p & v973991 | !hmaster1_p & v9738aa;
assign v9d2683 = hready_p & v84564b | !hready_p & !v9d2682;
assign v973a29 = hmaster1_p & v97398d | !hmaster1_p & v9739f4;
assign v9d269d = hbusreq1_p & v9d2694 | !hbusreq1_p & v845647;
assign v9998e1 = hgrant2_p & v9998d8 | !hgrant2_p & !v9998e0;
assign v9d2688 = hready & v9d2687 | !hready & !v84563c;
assign v8ea88f = hbusreq1_p & v8ea7e9 | !hbusreq1_p & v8ea88e;
assign v973967 = hmaster0_p & v9738e7 | !hmaster0_p & !v973966;
assign v9adcf8 = jx1_p & v9adbe6 | !jx1_p & v9adcf7;
assign v9739c7 = hbusreq0_p & v9738b8 | !hbusreq0_p & v973955;
assign v9ed445 = hlock1_p & v973893 | !hlock1_p & v84563c;
assign v984f76 = hmaster0_p & v984ea7 | !hmaster0_p & v84563c;
assign v985637 = hbusreq0_p & v985636 | !hbusreq0_p & v84563c;
assign v999920 = hbusreq2 & v999913 | !hbusreq2 & v99991f;
assign v8ea924 = hgrant2_p & v8ea7f8 | !hgrant2_p & v8ea923;
assign v9d2726 = hbusreq0_p & v9d2725 | !hbusreq0_p & v9d267e;
assign v9adc99 = hmaster1_p & v9adc93 | !hmaster1_p & !v9adc98;
assign v845644 = hlock0_p & v84563c | !hlock0_p & !v84563c;
assign v9999a8 = decide_p & v9999a2 | !decide_p & !v84565e;
assign v9d2725 = hmaster1_p & v9d2724 | !hmaster1_p & !v9d2671;
assign v97394d = hbusreq0_p & v97394a | !hbusreq0_p & v97394c;
assign v9d27a1 = hbusreq2 & v9d279a | !hbusreq2 & v9d27a0;
assign v984f48 = hlock0_p & v984f47 | !hlock0_p & v985540;
assign v9854fe = hready & v9854fd | !hready & v9ed456;
assign v8ea8d5 = hgrant0_p & v8ea8cc | !hgrant0_p & v8ea8d4;
assign v99658b = hbusreq0_p & v996588 | !hbusreq0_p & v99658a;
assign v9738dd = hmaster0_p & v97388f | !hmaster0_p & v9738dc;
assign v9baf62 = stateG10_1_p & v9baf5f | !stateG10_1_p & !v9baf61;
assign v8c20cd = hbusreq1_p & v8c20cb | !hbusreq1_p & !v8c20cc;
assign v9adc62 = hgrant1_p & v9adbeb | !hgrant1_p & !v9adc61;
assign v9a6aa1 = stateG2_p & v84563c | !stateG2_p & v9a6aa0;
assign v999923 = hmaster1_p & v999922 | !hmaster1_p & !v99990b;
assign v9d276c = hready_p & v9d275a | !hready_p & v9d276b;
assign v8c1132 = hburst0_p & v84563c | !hburst0_p & v8c1131;
assign v9a6ab7 = hlock0_p & v9a6ab6 | !hlock0_p & v84563c;
assign v9baf2a = stateG2_p & v84563c | !stateG2_p & !a2fb4c;
assign a15486 = hready_p & a15446 | !hready_p & a15485;
assign v9965b0 = hmaster1_p & v9965af | !hmaster1_p & v996569;
assign v9d266e = hbusreq1 & v9d266d | !hbusreq1 & v84563c;
assign v98559a = hmaster0_p & v985598 | !hmaster0_p & v985599;
assign v8e79a9 = locked_p & v8e799a | !locked_p & v84563c;
assign v98553c = hmaster0_p & v98553b | !hmaster0_p & v84563c;
assign v9adce3 = hbusreq0_p & v9adcdc | !hbusreq0_p & v9adce2;
assign v9d2799 = hgrant0_p & v84563c | !hgrant0_p & !v9d2797;
assign v9ed453 = decide_p & v9ed452 | !decide_p & v84563c;
assign v9ed489 = hmaster0_p & v9ed471 | !hmaster0_p & v9ed488;
assign v9ed476 = hmastlock_p & v9ed475 | !hmastlock_p & v84563c;
assign v984e55 = hgrant1_p & v98548f | !hgrant1_p & v84563c;
assign v9854d3 = hmaster0_p & v84563c | !hmaster0_p & v9854d1;
assign v8ea82c = hbusreq1_p & v8ea82a | !hbusreq1_p & v8ea82b;
assign v9baef2 = jx0_p & v9baea1 | !jx0_p & v9baef1;
assign v9d27a3 = hmaster1_p & v9d26fc | !hmaster1_p & v9d26fa;
assign v9baf05 = hmaster0_p & v9baf04 | !hmaster0_p & v845656;
assign v9999a1 = hbusreq0_p & v9999a0 | !hbusreq0_p & v84563c;
assign v9adc9b = decide_p & v9adc92 | !decide_p & v9adc9a;
assign v8ea814 = hbusreq1_p & v8ea813 | !hbusreq1_p & v8ea7e9;
assign v973958 = hready_p & v973943 | !hready_p & !v973957;
assign v9adc7d = hmaster1_p & v9adc78 | !hmaster1_p & v9adc7c;
assign v9738eb = stateG10_1_p & v97388d | !stateG10_1_p & v9738ea;
assign v84566a = stateG3_0_p & v84563c | !stateG3_0_p & !v84563c;
assign v973a09 = hmaster1_p & v9738cd | !hmaster1_p & !v973a08;
assign v9738f6 = hmaster0_p & v973885 | !hmaster0_p & !v9738e3;
assign v99657f = hmaster0_p & v996559 | !hmaster0_p & !v99657e;
assign v9ed40e = locked_p & v84563c | !locked_p & v973885;
assign v9ed44e = hbusreq1_p & v9ed44d | !hbusreq1_p & !v84563c;
assign a15448 = hmaster0_p & a15447 | !hmaster0_p & a15433;
assign v98549c = stateG2_p & v84563c | !stateG2_p & v98549b;
assign v9738b7 = hmaster0_p & v973885 | !hmaster0_p & v97388a;
assign v985606 = hmaster1_p & v985605 | !hmaster1_p & v84563c;
assign v8ea80c = hmaster1_p & v8ea801 | !hmaster1_p & v8ea80b;
assign v9baf34 = hmaster0_p & v9baf32 | !hmaster0_p & v9baf30;
assign v8ea809 = stateG10_1_p & v84563c | !stateG10_1_p & v8ea802;
assign v973940 = hmaster0_p & v97393f | !hmaster0_p & v97388c;
assign v9bae9d = decide_p & v9bae98 | !decide_p & v84563c;
assign v98555a = hmaster1_p & v985559 | !hmaster1_p & v84563c;
assign v9738f8 = hmaster1_p & v9738f6 | !hmaster1_p & v9738ed;
assign v973934 = decide_p & v97390c | !decide_p & v973933;
assign v973a2d = decide_p & v973a2a | !decide_p & v973a2c;
assign v9d2780 = hbusreq1_p & v9d2694 | !hbusreq1_p & !v9d277f;
assign v9854c9 = hmaster1_p & v9854c6 | !hmaster1_p & v9854c8;
assign v9738d5 = hmaster1_p & v9738cd | !hmaster1_p & !v9738d4;
assign v8c111a = locked_p & v8c1119 | !locked_p & !v84563c;
assign v9965d0 = hgrant2_p & v9965b3 | !hgrant2_p & v9965cf;
assign a1540e = hmaster0_p & v84563c | !hmaster0_p & a153c2;
assign v98551a = hmaster1_p & v985518 | !hmaster1_p & v9854df;
assign v86cfb3 = stateA1_p & v84563c | !stateA1_p & !v866c94;
assign v9baf83 = hmaster0_p & v84565c | !hmaster0_p & v9baf82;
assign v9ed43f = locked_p & v9ed43e | !locked_p & v973889;
assign v9d2734 = decide_p & v9d2733 | !decide_p & v9d2681;
assign v9739cc = decide_p & v973960 | !decide_p & v9739cb;
assign v9738e3 = hbusreq1_p & v9738cb | !hbusreq1_p & !v9738e2;
assign v9933cf = decide_p & v9933c9 | !decide_p & v9933ce;
assign v98562f = hbusreq0_p & v98562e | !hbusreq0_p & v84563c;
assign v9adc81 = hmaster1_p & v9adc7f | !hmaster1_p & !v9adc7c;
assign v9ed433 = hmastlock_p & v9ed432 | !hmastlock_p & v84563c;
assign v9855c2 = hmaster1_p & v9855c1 | !hmaster1_p & v9854c8;
assign v9739d8 = hbusreq0_p & v97390e | !hbusreq0_p & v973995;
assign v9ed417 = hbusreq1_p & v9ed416 | !hbusreq1_p & v84563c;
assign v973a4b = jx0_p & v9739e7 | !jx0_p & v973a4a;
assign v9adca9 = hgrant1_p & v9adc77 | !hgrant1_p & !v84563c;
assign v9ed4bf = hbusreq1_p & v9ed4be | !hbusreq1_p & !v84563c;
assign v973921 = hbusreq0_p & v97391a | !hbusreq0_p & v973920;
assign v9855d2 = hlock0_p & v9855d1 | !hlock0_p & v9855be;
assign v8ea800 = hgrant1_p & v84563c | !hgrant1_p & v8ea7e6;
assign v9bae97 = hbusreq2 & v9bae90 | !hbusreq2 & v9bae96;
assign v9854dd = hmaster0_p & v84563c | !hmaster0_p & v9854dc;
assign v9739b8 = hmaster0_p & v973885 | !hmaster0_p & !v9739a8;
assign v8ea914 = hbusreq0_p & v8ea881 | !hbusreq0_p & v8ea913;
assign v9adc82 = hbusreq0_p & v9adc80 | !hbusreq0_p & v9adc81;
assign v973991 = hmaster0_p & v973885 | !hmaster0_p & !v97388d;
assign v8ea91a = hmaster0_p & v8ea7ec | !hmaster0_p & v8ea82c;
assign v9ed446 = hbusreq1_p & v9ed445 | !hbusreq1_p & !v84563c;
assign v9ed4ae = hbusreq1_p & v9ed4ad | !hbusreq1_p & !v84563c;
assign v9ed42a = hmastlock_p & v9ed429 | !hmastlock_p & v84563c;
assign a1541e = stateG2_p & v84563c | !stateG2_p & a1541d;
assign v9adc2c = stateG10_1_p & v9adbee | !stateG10_1_p & v9adc2a;
assign v984f88 = hbusreq2 & v984f86 | !hbusreq2 & v984f87;
assign v9adcc6 = hbusreq1_p & v9adcc4 | !hbusreq1_p & !v9adcc5;
assign v8ea93a = jx2_p & v8ea92a | !jx2_p & v8ea939;
assign v984f65 = hgrant0_p & v984f5a | !hgrant0_p & v984f64;
assign v9adcc7 = hmaster0_p & v9adcb9 | !hmaster0_p & !v9adcc6;
assign v9d267c = hmaster1_p & v845652 | !hmaster1_p & !v9d2673;
assign v9ed4b6 = hmaster1_p & v9ed4b2 | !hmaster1_p & v9ed4b5;
assign v999981 = hbusreq0 & v999980 | !hbusreq0 & !v99997b;
assign v9d2671 = hmaster0_p & v845647 | !hmaster0_p & v84563c;
assign v9baf6e = hgrant1_p & v9baf6d | !hgrant1_p & v9ed41d;
assign v9999bf = hmastlock_p & v9999be | !hmastlock_p & v84563c;
assign v9d2775 = hmaster0_p & v9d276e | !hmaster0_p & !v84563c;
assign v8c20c2 = hlock1_p & v84565c | !hlock1_p & !v8c20c1;
assign v9739a2 = hmaster1_p & v9739a1 | !hmaster1_p & !v97395d;
assign v9933b8 = hmaster0_p & v84563c | !hmaster0_p & !v9933b7;
assign v9baf0e = hbusreq1 & v9ed476 | !hbusreq1 & v9ed487;
assign v9965a0 = hmaster1_p & v9adc49 | !hmaster1_p & v99659f;
assign v9adc67 = hbusreq0_p & v9adc5f | !hbusreq0_p & v9adc66;
assign v9bae87 = hmaster0_p & v9ed423 | !hmaster0_p & v9bae86;
assign v9965b7 = hmaster1_p & v9965b6 | !hmaster1_p & v99657b;
assign v9738c8 = hbusreq0_p & v9738c2 | !hbusreq0_p & !v9738c7;
assign v9999de = hmaster1_p & a154a3 | !hmaster1_p & v9999dd;
assign v9ed4bb = hmaster1_p & v845646 | !hmaster1_p & !v9ed4ba;
assign v984ec0 = hgrant2_p & v985649 | !hgrant2_p & v984ebf;
assign v98564c = busreq_p & v9a6a96 | !busreq_p & v98564b;
assign v9adc3f = hbusreq0_p & v9adc3c | !hbusreq0_p & v9adc3e;
assign v8e79d7 = decide_p & v8e79d6 | !decide_p & v8e79bd;
assign v9739e3 = hgrant0_p & v9739e0 | !hgrant0_p & v9739e2;
assign v9d2678 = hmaster1_p & v9d2676 | !hmaster1_p & !v9d2673;
assign v8ea854 = hbusreq0_p & v8ea852 | !hbusreq0_p & v8ea853;
assign a153eb = hmaster0_p & a153cf | !hmaster0_p & v845648;
assign v9baf74 = hmaster1_p & v9baf56 | !hmaster1_p & v9baf73;
assign v984eb4 = hmaster0_p & v984ea7 | !hmaster0_p & v984eb3;
assign v98557b = hbusreq1_p & v98557a | !hbusreq1_p & v84563c;
assign v8ea808 = hgrant0_p & v8ea7ff | !hgrant0_p & v8ea807;
assign v984f70 = hmaster0_p & v985520 | !hmaster0_p & v84563c;
assign v9baec9 = hbusreq2 & v9baeb1 | !hbusreq2 & v9baec8;
assign v973942 = hbusreq0_p & v973941 | !hbusreq0_p & v973939;
assign v999917 = hburst0 & a153cc | !hburst0 & v999916;
assign v98551b = hlock0_p & v985519 | !hlock0_p & v98551a;
assign v8c1133 = stateG2_p & v84563c | !stateG2_p & !v8c1132;
assign v9998ea = stateA1_p & v8e7990 | !stateA1_p & !v9ed426;
assign v984f96 = jx1_p & v984ee2 | !jx1_p & v984f95;
assign v984ef1 = hbusreq1_p & v984eef | !hbusreq1_p & v984ef0;
assign v9d2665 = hburst0 & v9d2663 | !hburst0 & v9d2664;
assign v999939 = hmaster0_p & v9baf8d | !hmaster0_p & v84563c;
assign v9adc65 = hmaster0_p & v9adc64 | !hmaster0_p & v9adbee;
assign v9933d0 = hready_p & v9933cf | !hready_p & !v84563c;
assign v984f50 = hmaster1_p & v84563c | !hmaster1_p & v985609;
assign v9adbe8 = busreq_p & v84566e | !busreq_p & !v9adbe7;
assign a154fc = hlock1_p & a154f6 | !hlock1_p & !a154fb;
assign v8e79ad = hready_p & v8e7997 | !hready_p & v8e79ac;
assign v8ea8c2 = hbusreq2 & v8ea8c0 | !hbusreq2 & v8ea8c1;
assign v8ea92d = hbusreq0_p & v8ea92b | !hbusreq0_p & v8ea92c;
assign v8ea83b = hmaster1_p & v8ea815 | !hmaster1_p & v8ea83a;
assign v9baf41 = hready_p & v9baef5 | !hready_p & v9baf40;
assign v9d269e = hmaster0_p & v845647 | !hmaster0_p & v9d269d;
assign v9d26ff = hgrant0_p & v84563c | !hgrant0_p & v9d26fe;
assign v9854ee = stateG2_p & v84563c | !stateG2_p & v9854ed;
assign v9d2752 = hmaster1_p & v9d2724 | !hmaster1_p & !v9d2673;
assign v984f3e = hbusreq0_p & v984f3d | !hbusreq0_p & v845641;
assign v9adcaf = hmaster1_p & v9adca8 | !hmaster1_p & !v9adcae;
assign v99991a = hmaster1_p & v999919 | !hmaster1_p & !v99990b;
assign v9adc3c = hmaster1_p & v9adc38 | !hmaster1_p & v9adc3b;
assign v98554b = stateG2_p & v84563c | !stateG2_p & v98554a;
assign v985590 = hmastlock_p & v98558f | !hmastlock_p & v84563c;
assign v996556 = hmaster0_p & v996553 | !hmaster0_p & v996552;
assign v9998ef = locked_p & v9998ee | !locked_p & v84563c;
assign v9adc30 = hmaster0_p & v9adc2d | !hmaster0_p & v9adbee;
assign v97394c = hmaster1_p & v9738a5 | !hmaster1_p & v97394b;
assign v9a6a9d = stateG3_0_p & v84563c | !stateG3_0_p & !v8901af;
assign v9855ba = hbusreq2 & v9855a6 | !hbusreq2 & v9855b9;
assign v9adcd7 = hmaster1_p & v9adc75 | !hmaster1_p & !v9adc7a;
assign v9ed4a4 = hburst0 & v9ed4a2 | !hburst0 & v9ed4a3;
assign v985581 = hgrant1_p & v84563c | !hgrant1_p & v84565c;
assign v9998aa = hmaster1_p & v9ed423 | !hmaster1_p & v9998a9;
assign v973a17 = decide_p & v973a0f | !decide_p & v973a16;
assign v985495 = stateG2_p & v84563c | !stateG2_p & v985494;
assign v9a6abc = hlock1_p & v9a6abb | !hlock1_p & v84563c;
assign v9738ae = hmaster1_p & v9738a5 | !hmaster1_p & v9738ad;
assign v9d267b = hmaster1_p & v845652 | !hmaster1_p & !v9d2671;
assign v996551 = stateG2_p & v84563c | !stateG2_p & a2bb5d;
assign v960f66 = hready_p & v84565e | !hready_p & !v845652;
assign v9baf84 = hmaster1_p & a154a3 | !hmaster1_p & v9baf83;
assign v98552b = hmaster0_p & v84563c | !hmaster0_p & v98552a;
assign v97391b = locked_p & v973883 | !locked_p & v973885;
assign v9a6acc = hbusreq1_p & v9a6aca | !hbusreq1_p & v9a6acb;
assign v8c116f = stateG3_2_p & v84563c | !stateG3_2_p & v8c116e;
assign v98558a = hmaster1_p & v985588 | !hmaster1_p & v985589;
assign v9d27c6 = jx0_p & v9d278b | !jx0_p & v9d27c5;
assign v9854d7 = hbusreq0_p & v9854d6 | !hbusreq0_p & v9854d5;
assign v9854a1 = hlock1_p & v985498 | !hlock1_p & v9854a0;
assign v984e78 = decide_p & v984e65 | !decide_p & v984e77;
assign a15509 = hmaster0_p & a15508 | !hmaster0_p & v84563c;
assign v8901af = stateG3_1_p & v84563c | !stateG3_1_p & !v845658;
assign v8ea8a7 = hbusreq0_p & v8ea87c | !hbusreq0_p & v8ea8a5;
assign v9855f1 = hmaster1_p & v9855ef | !hmaster1_p & v9855b5;
assign v9adcbc = hmaster0_p & v9adcb9 | !hmaster0_p & v9adc75;
assign v9d26d9 = decide_p & v9d26d8 | !decide_p & v9d26a2;
assign v9ecda3 = decide_p & v9ed4f5 | !decide_p & v9ed4c6;
assign v9bae8a = hlock2_p & v9bae89 | !hlock2_p & !v84563c;
assign v9bae96 = hmaster1_p & v9bae95 | !hmaster1_p & v84563c;
assign v9854ce = hready & v9854cd | !hready & !v84563c;
assign v9999e4 = hgrant0_p & v9999d9 | !hgrant0_p & !v84563c;
assign v9adc03 = hmaster0_p & v9adc02 | !hmaster0_p & v9adbed;
assign v8ea7eb = stateG10_1_p & v8ea7ea | !stateG10_1_p & !v8ea7e9;
assign v984f52 = hgrant0_p & v984f51 | !hgrant0_p & v984e61;
assign v9854e8 = hbusreq0_p & v9854e7 | !hbusreq0_p & v9854e6;
assign a153cd = hmastlock_p & a153cc | !hmastlock_p & v84563c;
assign v9a6ab0 = hlock2_p & v9a6aaa | !hlock2_p & v9a6aaf;
assign v9999e6 = hgrant0_p & v9999e5 | !hgrant0_p & !v84563c;
assign v9855e5 = decide_p & v9855db | !decide_p & v9855e4;
assign v8e79c7 = hgrant0_p & v8e79bf | !hgrant0_p & v8e79c6;
assign v9739ca = hbusreq0_p & v9738e9 | !hbusreq0_p & v973968;
assign v9855ac = hready & v9855a7 | !hready & !v9855ab;
assign v8ea7f3 = hmaster1_p & v8ea7e9 | !hmaster1_p & v8ea7f2;
assign v9ed477 = hbusreq1_p & v9ed476 | !hbusreq1_p & !v84563c;
assign v985611 = hlock2_p & v98560e | !hlock2_p & v985610;
assign v99999a = decide_p & v999982 | !decide_p & v84565e;
assign v999932 = hready_p & v999901 | !hready_p & !v999931;
assign v999916 = hburst1 & a153cc | !hburst1 & v999915;
assign v8c20db = hmaster1_p & v8c20d6 | !hmaster1_p & v8c20da;
assign v9d2768 = hgrant0_p & v9d2752 | !hgrant0_p & v9d2767;
assign v996581 = hbusreq0_p & v99657d | !hbusreq0_p & v996580;
assign v8e7993 = locked_p & v8e7992 | !locked_p & v84563c;
assign a153bc = stateG2_p & v84563c | !stateG2_p & !a153bb;
assign v9d270b = decide_p & v9d2705 | !decide_p & v9d270a;
assign v8e79a6 = hlock0_p & v8e79a4 | !hlock0_p & v8e79a5;
assign v8e79d5 = hbusreq0_p & v8e79b7 | !hbusreq0_p & v8e79d4;
assign v9ed52f = hgrant0_p & v84563c | !hgrant0_p & !v9ed4b4;
assign v9998f7 = hmaster0_p & v973885 | !hmaster0_p & v9ed43f;
assign v9933be = hlock0_p & v9933bd | !hlock0_p & v8c20be;
assign v9ed425 = hburst1_p & v84563c | !hburst1_p & !v8e7989;
assign v9baf72 = hbusreq1_p & v9baf6e | !hbusreq1_p & v9baf71;
assign v9855f8 = hgrant2_p & v9855d0 | !hgrant2_p & v9855f7;
assign v9854e2 = hbusreq0_p & v9854e1 | !hbusreq0_p & v9854e0;
assign v9d2761 = hmaster1_p & v9d275e | !hmaster1_p & !v9d2673;
assign v985515 = hmaster1_p & v985513 | !hmaster1_p & v9854b8;
assign v9ed498 = hmaster0_p & v9ed410 | !hmaster0_p & v9ed41a;
assign v9baeff = busreq_p & v9ed457 | !busreq_p & v9baefe;
assign v984f5f = hbusreq1_p & v984f5c | !hbusreq1_p & !v984f5e;
assign v8ea7e7 = hmaster0_p & v84563c | !hmaster0_p & v8ea7e6;
assign v9ed4e2 = hbusreq0 & v9ed4de | !hbusreq0 & v9ed4e1;
assign v973a30 = hmaster1_p & v973a2f | !hmaster1_p & v97397b;
assign v973890 = hmaster0_p & v97388f | !hmaster0_p & v97388c;
assign v985493 = hburst0_p & v9a6a95 | !hburst0_p & v985492;
assign v973920 = hmaster1_p & v97391f | !hmaster1_p & !v9738d8;
assign v9ed4a7 = hgrant1_p & v84565c | !hgrant1_p & v9ed4a6;
assign v984e53 = stateG10_1_p & v98564e | !stateG10_1_p & v984e52;
assign v9adc51 = hready_p & v9adc41 | !hready_p & !v9adc50;
assign v9baea5 = hmaster1_p & v9baea4 | !hmaster1_p & a154a3;
assign v9baf68 = stateG10_1_p & v9ed419 | !stateG10_1_p & v9baf67;
assign v8ea8c8 = hlock1 & v8ea818 | !hlock1 & v8ea819;
assign v8c111b = hmaster0_p & v84563c | !hmaster0_p & !v8c111a;
assign v8c113c = hmaster1_p & v8c113b | !hmaster1_p & !v84563c;
assign v9ed413 = hburst1 & v9ed412 | !hburst1 & v84563c;
assign v9855fe = hmaster0_p & v84563c | !hmaster0_p & v9855fd;
assign v9739ef = hmaster1_p & v97389a | !hmaster1_p & v9739ee;
assign v9d26d0 = hgrant1_p & v845647 | !hgrant1_p & !v84563c;
assign v9b40d0 = jx0_p & v9b40c3 | !jx0_p & v9b40cd;
assign v9baf48 = hmaster1_p & v9baf46 | !hmaster1_p & v9baf47;
assign v9baf29 = busreq_p & v9baf28 | !busreq_p & a153cc;
assign v8ea881 = hmaster1_p & v8ea880 | !hmaster1_p & v8ea816;
assign v9adccc = hready_p & v9adcc0 | !hready_p & !v9adccb;
assign v97388e = locked_p & v84563c | !locked_p & v97388d;
assign v9d27b8 = decide_p & v9d27b7 | !decide_p & !v9d2681;
assign v9998d7 = decide_p & v9998d6 | !decide_p & v84563c;
assign v8ea8e6 = hlock2 & v8ea8e3 | !hlock2 & v8ea8e5;
assign v984ea5 = hgrant1_p & v985520 | !hgrant1_p & !v84563c;
assign v9738cb = hgrant1_p & v97388c | !hgrant1_p & !v973889;
assign v984f4f = hgrant0_p & v984f4e | !hgrant0_p & v984e61;
assign v8c113f = hmaster1_p & v84563c | !hmaster1_p & v8c111b;
assign v984ee3 = hmaster0_p & v9854ce | !hmaster0_p & v84563c;
assign a14d58 = hready_p & a14d4d | !hready_p & a14d49;
assign v8ea898 = hmaster1_p & v8ea889 | !hmaster1_p & v8ea897;
assign v985597 = hgrant1_p & v845641 | !hgrant1_p & !v84563c;
assign v985643 = hmaster0_p & v985642 | !hmaster0_p & v84563c;
assign v973a35 = hmaster0_p & v9738ca | !hmaster0_p & v973a0b;
assign a15492 = hbusreq0_p & a1542e | !hbusreq0_p & a15491;
assign v9a6ad4 = hbusreq1_p & v9a6aa2 | !hbusreq1_p & v84563c;
assign v984e62 = hlock0_p & v984e5c | !hlock0_p & v984e61;
assign v8c1136 = hmastlock_p & v8c1135 | !hmastlock_p & !v84563c;
assign v9d26e6 = hbusreq0_p & v9d26e4 | !hbusreq0_p & !v9d26e5;
assign v9f3574 = decide_p & v9f356c | !decide_p & v845646;
assign v985569 = locked_p & v985568 | !locked_p & v84563c;
assign v8ea8cb = hmaster1_p & v8ea880 | !hmaster1_p & v8ea8ca;
assign v8c117e = hready_p & v8c117c | !hready_p & !v8c117d;
assign v9adc39 = stateG10_1_p & v9adbee | !stateG10_1_p & v9adc29;
assign v8ea929 = hgrant2_p & v8ea926 | !hgrant2_p & v8ea928;
assign v9adbff = hmaster0_p & v9adbfe | !hmaster0_p & !v9adbed;
assign v8c1178 = hmaster0_p & v8c1177 | !hmaster0_p & v84563c;
assign v996595 = hgrant0_p & v99657a | !hgrant0_p & v996594;
assign v9739aa = hmaster1_p & v9739a9 | !hmaster1_p & !v973964;
assign v9d26c6 = hbusreq0 & v9d26c3 | !hbusreq0 & v9d26c5;
assign v999936 = hmaster0_p & v9baf63 | !hmaster0_p & v84563c;
assign v9a6add = hbusreq0_p & v9a6abf | !hbusreq0_p & v9a6adc;
assign v9ed4fc = hlock1_p & v9ed4fb | !hlock1_p & !v84563c;
assign v9d2754 = hbusreq2 & v9d2751 | !hbusreq2 & v9d2753;
assign v9baf49 = hbusreq0_p & v9baf45 | !hbusreq0_p & v9baf48;
assign a154c1 = hburst1_p & v96ef3e | !hburst1_p & !v85a40d;
assign v9d271f = hmaster0_p & v9d271e | !hmaster0_p & !v84563c;
assign v9bae7a = hmaster1_p & v9bae79 | !hmaster1_p & v84565c;
assign a14d8b = hmaster0_p & a154d4 | !hmaster0_p & a153d1;
assign v8c1146 = hlock1_p & v8c1145 | !hlock1_p & !v84563c;
assign v9baf52 = hbusreq1 & v973885 | !hbusreq1 & !v84563c;
assign v9baf3f = hlock2_p & v9baf26 | !hlock2_p & v9baf3e;
assign v9ed41b = hmaster0_p & v84563c | !hmaster0_p & v9ed41a;
assign a15420 = locked_p & a1541f | !locked_p & v84563c;
assign v985632 = hmaster0_p & v985624 | !hmaster0_p & v985631;
assign v985513 = hmaster0_p & v9854cf | !hmaster0_p & v9854b3;
assign v8c1157 = hmaster0_p & v8c113a | !hmaster0_p & !v84563c;
assign v8e79b2 = hmaster0_p & v8e79b1 | !hmaster0_p & v84563c;
assign v9d2691 = hready & v84565c | !hready & v84563c;
assign jx0 = v9adcf8;
assign v9adbf8 = stateG3_2_p & v84563c | !stateG3_2_p & v84566a;
assign v8ea8e5 = hbusreq0 & v8ea8e1 | !hbusreq0 & v8ea8e4;
assign a14d4b = hbusreq0_p & a1550b | !hbusreq0_p & v845646;
assign v9adca6 = hlock1_p & v9adca5 | !hlock1_p & !v9adc75;
assign v985602 = hbusreq0 & v985601 | !hbusreq0 & v84563c;
assign v9739e0 = hbusreq0_p & v9739df | !hbusreq0_p & v9739b6;
assign v9854f2 = hburst1_p & v8ea7e2 | !hburst1_p & !v84563c;
assign v984e70 = hgrant1_p & v984e6f | !hgrant1_p & v84563c;
assign v9adbe6 = jx0_p & v854658 | !jx0_p & !v854662;
assign v984eab = stateG10_1_p & v84563c | !stateG10_1_p & v984eaa;
assign v8ea86e = hgrant0_p & v8ea86d | !hgrant0_p & v8ea86a;
assign v8c20d5 = hbusreq1_p & v8c20c2 | !hbusreq1_p & !v84563c;
assign v984f82 = hmaster1_p & v984f76 | !hmaster1_p & v984f81;
assign v984e67 = stateG10_1_p & v84563c | !stateG10_1_p & !v9d2691;
assign v9d2684 = hburst1 & v845668 | !hburst1 & !v84563c;
assign v8c1150 = hgrant1_p & v8c114c | !hgrant1_p & v84563c;
assign v99992f = hbusreq2 & v999928 | !hbusreq2 & v99992e;
assign v9a6aab = hmaster0_p & v9a6aa2 | !hmaster0_p & v84563c;
assign v9855b7 = hbusreq0_p & v9855b2 | !hbusreq0_p & v9855b6;
assign v9738da = hbusreq0_p & v9738d5 | !hbusreq0_p & v9738d9;
assign v9965ce = decide_p & v9965b1 | !decide_p & v9965cd;
assign v9998e4 = hmaster0_p & v9baf43 | !hmaster0_p & v84563c;
assign v973964 = hmaster0_p & v973963 | !hmaster0_p & !v9738e3;
assign v973a44 = hbusreq0_p & v9739b9 | !hbusreq0_p & v973a43;
assign v9d26f7 = stateG10_1_p & v9d268c | !stateG10_1_p & !v9d26f6;
assign v985552 = hmastlock_p & v985551 | !hmastlock_p & v84563c;
assign v973899 = locked_p & v86cfb3 | !locked_p & v973889;
assign v9d26a6 = stateA1_p & v9d26a5 | !stateA1_p & v8c1130;
assign v973889 = hmastlock_p & v86cfb3 | !hmastlock_p & v845666;
assign v8c1151 = stateG10_1_p & v84563c | !stateG10_1_p & v8c1150;
assign v8e79d2 = hbusreq1_p & v8e79b1 | !hbusreq1_p & v84563c;
assign v9d26f6 = hgrant1_p & v845647 | !hgrant1_p & !v9d268c;
assign v845666 = stateA1_p & v84563c | !stateA1_p & !v84563c;
assign v9d275a = hbusreq0 & v9d2758 | !hbusreq0 & !v9d2759;
assign v99657c = hmaster1_p & v9adc1a | !hmaster1_p & v99657b;
assign v8ea8d9 = hlock2 & v8ea8d6 | !hlock2 & v8ea8d8;
assign v9baeae = hmaster1_p & v9baead | !hmaster1_p & v84563c;
assign a1550e = hgrant0_p & v84563c | !hgrant0_p & a1550c;
assign v8c117b = hgrant0_p & v8c1141 | !hgrant0_p & v8c117a;
assign v9739d6 = hlock0_p & v9739d4 | !hlock0_p & v9739d5;
assign v984eaf = hbusreq0_p & v984eae | !hbusreq0_p & v985645;
assign v9ed4c9 = hready_p & v9ed4c7 | !hready_p & !v9ed4c8;
assign v984f72 = hmaster1_p & v984f70 | !hmaster1_p & v984f71;
assign v8c1126 = hmaster0_p & v8c1123 | !hmaster0_p & !v84563c;
assign v9d26b1 = hmaster1_p & v9d26b0 | !hmaster1_p & !v9d2671;
assign v9739f0 = hbusreq0_p & v9739ed | !hbusreq0_p & v9739ef;
assign v97391e = hbusreq1_p & v9738c9 | !hbusreq1_p & !v97391d;
assign v8e79bf = hmaster1_p & v84563c | !hmaster1_p & v8e79aa;
assign v973907 = hmaster0_p & v973885 | !hmaster0_p & !v97389e;
assign v8543c7 = hbusreq2_p & v85bb54 | !hbusreq2_p & !v84563c;
assign v984e6a = hgrant1_p & v985618 | !hgrant1_p & !v84563c;
assign v8c115d = hbusreq1_p & v8c115b | !hbusreq1_p & v8c115c;
assign v9adc85 = hlock1_p & v9adc75 | !hlock1_p & !v84563c;
assign v9ed474 = hburst1 & v973892 | !hburst1 & !v84563c;
assign v9d27aa = hmaster0_p & v9d27a9 | !hmaster0_p & !v84563c;
assign v9a6aa4 = hbusreq1_p & v9a6aa3 | !hbusreq1_p & v84563c;
assign v9ed43b = hlock1_p & v973885 | !hlock1_p & !v84563c;
assign v8ea90d = hmaster1_p & v8ea909 | !hmaster1_p & v8ea90c;
assign v985502 = hmaster0_p & v84563c | !hmaster0_p & v985500;
assign v8ea8bc = hmaster1_p & v8ea8b8 | !hmaster1_p & v8ea897;
assign v985546 = stateG2_p & v84563c | !stateG2_p & !v985545;
assign v8ea804 = stateG10_1_p & v84563c | !stateG10_1_p & v8ea803;
assign v9933d3 = hready_p & v9933d2 | !hready_p & !v84563c;
assign v9d2795 = hready_p & v84564b | !hready_p & !v9d2794;
assign v8ea8b5 = hmaster1_p & v8ea8b4 | !hmaster1_p & v8ea816;
assign v9855a3 = hmaster1_p & v985588 | !hmaster1_p & v9855a2;
assign v9854bf = hburst0_p & a3134f | !hburst0_p & v9854be;
assign v9998ad = hgrant0_p & v9998ac | !hgrant0_p & !v84563c;
assign v9739d1 = hgrant2_p & v9739c9 | !hgrant2_p & v9739d0;
assign v9ed56a = hgrant0_p & v84563c | !hgrant0_p & !v9ed4ff;
assign a1542e = hmaster1_p & a1542d | !hmaster1_p & a153c4;
assign v9bae98 = hlock2_p & v9bae97 | !hlock2_p & v84563c;
assign v985491 = hbusreq1_p & v985490 | !hbusreq1_p & v84563c;
assign v98555e = hmaster0_p & v9ed423 | !hmaster0_p & v9854c7;
assign v996571 = hlock2_p & v99656b | !hlock2_p & v996570;
assign v973969 = hbusreq0_p & v973965 | !hbusreq0_p & v973968;
assign v9ed465 = hburst1 & v9ed462 | !hburst1 & v9ed464;
assign v9933c7 = hmaster0_p & v9933c6 | !hmaster0_p & !v84563c;
assign v9baf2e = hburst0 & v9baf29 | !hburst0 & v9baf2d;
assign v9854c4 = hready & v9854c3 | !hready & v84563c;
assign v8ea868 = hmaster1_p & v8ea867 | !hmaster1_p & v8ea828;
assign v99654f = locked_p & v9adbfe | !locked_p & !v9adbee;
assign v973994 = hmaster1_p & v97390d | !hmaster1_p & !v973940;
assign v984f8c = decide_p & v84563c | !decide_p & v985645;
assign v9adcbe = hbusreq0_p & v9adcbb | !hbusreq0_p & v9adcbd;
assign v9d26b3 = hmaster1_p & v9d26b0 | !hmaster1_p & !v9d2673;
assign v9854ff = hlock1_p & v9854fc | !hlock1_p & v9854fe;
assign v99996a = hready_p & v999940 | !hready_p & v999969;
assign v9999d6 = hlock2_p & v9999d0 | !hlock2_p & v9999d5;
assign v8c1167 = hmaster0_p & v8c1166 | !hmaster0_p & !v84563c;
assign v9baf8e = hbusreq1_p & v84565c | !hbusreq1_p & a15507;
assign v9adcdf = stateG10_1_p & v9adcdd | !stateG10_1_p & v9adcde;
assign v984f85 = hgrant0_p & v984f80 | !hgrant0_p & v984f84;
assign v9d27bb = hgrant0_p & v84563c | !hgrant0_p & v9d27ba;
assign v9ed440 = hbusreq1_p & v9ed43f | !hbusreq1_p & v84563c;
assign v973a25 = hbusreq0_p & v973a23 | !hbusreq0_p & v973a24;
assign v9baf1f = hbusreq1_p & v9baf1a | !hbusreq1_p & v9baf1e;
assign v9738e8 = hmaster0_p & v9738e7 | !hmaster0_p & !v9738e3;
assign v9855a9 = stateG2_p & v84563c | !stateG2_p & v9855a8;
assign v9baf3a = hmaster0_p & v9baf32 | !hmaster0_p & v9ed481;
assign v8e79b9 = stateG10_1_p & v84563c | !stateG10_1_p & v8e79b3;
assign a14d70 = decide_p & a14d6f | !decide_p & v84565c;
assign v99658e = stateG10_1_p & v9adbee | !stateG10_1_p & !v99658d;
assign v9999a5 = hgrant0_p & v999934 | !hgrant0_p & !v84563c;
assign v8e79c0 = hgrant1_p & v84563c | !hgrant1_p & v8e79a9;
assign v985629 = hmaster1_p & v985625 | !hmaster1_p & v985628;
assign v9998f2 = hmaster1_p & v9baf93 | !hmaster1_p & a154a3;
assign v99993e = hgrant0_p & a14d3e | !hgrant0_p & !v84563c;
assign v999926 = hlock0_p & v999923 | !hlock0_p & v999925;
assign hgrant0 = !v9999f1;
assign v9738f2 = hmaster0_p & v973885 | !hmaster0_p & !v97388c;
assign v984eb3 = hbusreq1_p & v84565c | !hbusreq1_p & !v984eb2;
assign v9ed4b1 = hbusreq1_p & v9ed4b0 | !hbusreq1_p & !v84563c;
assign v9998a9 = hmaster0_p & v84563c | !hmaster0_p & v9bae86;
assign v9a6ae3 = hbusreq2_p & v9a6ad2 | !hbusreq2_p & v9a6ae2;
assign v9baf93 = hmaster0_p & v84565c | !hmaster0_p & v9ed434;
assign v8ea91e = hlock0 & v8ea91d | !hlock0 & v8ea915;
assign a153d2 = hlock1_p & v84563c | !hlock1_p & a153d1;
assign v9ed485 = hburst1 & v84563c | !hburst1 & !v973892;
assign v9999d2 = hlock0_p & v9999d1 | !hlock0_p & v84563c;
assign v985545 = stateA1_p & v985544 | !stateA1_p & !v985493;
assign v883467 = hburst0_p & v84563c | !hburst0_p & v8996a7;
assign v9a6aa7 = hmaster0_p & v9a6aa4 | !hmaster0_p & v84563c;
assign v97395a = hmaster1_p & v9738b0 | !hmaster1_p & v973959;
assign v9854b5 = hmaster1_p & v9854b4 | !hmaster1_p & v9854b3;
assign v9bae8f = hmaster0_p & v84563c | !hmaster0_p & !v9bae8e;
assign v8ea7f7 = decide_p & v8ea7ee | !decide_p & v8ea7f6;
assign v9739ea = hbusreq0_p & v973941 | !hbusreq0_p & v9739e9;
assign v9adcab = hgrant1_p & v9adca1 | !hgrant1_p & v9adc75;
assign v9738fa = hgrant0_p & v9738f5 | !hgrant0_p & v9738f9;
assign v97393b = hmaster0_p & v97389b | !hmaster0_p & !v97388d;
assign v9933c2 = hbusreq1_p & v9933c0 | !hbusreq1_p & !v9933c1;
assign v8c20c7 = decide_p & v8c20c6 | !decide_p & v84565c;
assign v9855b3 = hgrant1_p & v84563c | !hgrant1_p & v985520;
assign v973884 = busreq_p & v845666 | !busreq_p & !v84563c;
assign v9baf59 = hburst1 & a153bc | !hburst1 & v9baf58;
assign v9999ab = decide_p & v845642 | !decide_p & v84563c;
assign v9d27c0 = hgrant2_p & v9d27b9 | !hgrant2_p & v9d27bf;
assign v9adc1f = locked_p & v9adbfe | !locked_p & !v9adbeb;
assign v9ed48c = hbusreq0 & v9ed47a | !hbusreq0 & v9ed48b;
assign a154ed = hbusreq0_p & a154d6 | !hbusreq0_p & v84563c;
assign v9d274b = hbusreq0 & v9d26e5 | !hbusreq0 & v9d26e8;
assign v98556b = hbusreq1_p & v98556a | !hbusreq1_p & !v84563c;
assign v9baf8c = hgrant1_p & v9baf8b | !hgrant1_p & v84565c;
assign v98562a = hready & v9854fd | !hready & a153d0;
assign v8ea832 = hbusreq1 & v8ea818 | !hbusreq1 & v8ea831;
assign v9adc96 = hmaster0_p & v9adc95 | !hmaster0_p & v84563c;
assign v9ed418 = hmaster0_p & v9ed410 | !hmaster0_p & v9ed417;
assign v9d26fa = hbusreq1_p & v9d2694 | !hbusreq1_p & v9d26f9;
assign v8c20d9 = hbusreq1_p & v84565c | !hbusreq1_p & !v8c20d8;
assign v984ec6 = hmaster0_p & v985520 | !hmaster0_p & !v985592;
assign v9998a2 = hbusreq0 & v99989e | !hbusreq0 & v9998a1;
assign v9739be = decide_p & v973993 | !decide_p & v9739bd;
assign v9d279b = hgrant0_p & v84563c | !hgrant0_p & v845647;
assign v9d44c3 = jx2_p & v8543c7 | !jx2_p & !v84563c;
assign v9855cd = hmaster1_p & v9855cb | !hmaster1_p & v98552b;
assign v9998dd = hbusreq0 & v9998da | !hbusreq0 & v9998dc;
assign v8ea918 = hmaster0_p & v8ea7ec | !hmaster0_p & v8ea822;
assign v9933dc = hbusreq2_p & v9933d1 | !hbusreq2_p & v9933db;
assign v9999b4 = hready_p & v9999b2 | !hready_p & !v9999b3;
assign v973951 = hmaster1_p & v9738b0 | !hmaster1_p & v97394b;
assign v9738ef = hbusreq0_p & v9738e9 | !hbusreq0_p & v9738ee;
assign v9739fd = hready_p & v9739f2 | !hready_p & !v9739fc;
assign v97396a = hgrant0_p & v9738df | !hgrant0_p & v973969;
assign v9ecda6 = hbusreq2_p & v9ecda5 | !hbusreq2_p & v9ed533;
assign v9baf4d = hburst1 & v9baf4c | !hburst1 & v9baf01;
assign v9adc41 = decide_p & v9adc33 | !decide_p & v9adc40;
assign a14d9f = hlock0_p & a14d8c | !hlock0_p & a14d8e;
assign v9854f6 = busreq_p & v9854f4 | !busreq_p & !v9854f5;
assign v9ed458 = stateA1_p & a153cb | !stateA1_p & v9ed455;
assign v8763e4 = stateG3_0_p & v84563c | !stateG3_0_p & v887862;
assign v9d2738 = hmaster1_p & v9d2737 | !hmaster1_p & v845647;
assign v984f7d = hgrant0_p & v984f75 | !hgrant0_p & v984f7c;
assign v9baf4f = hmastlock_p & v9baf4e | !hmastlock_p & !v84563c;
assign v9965bc = hmaster1_p & v9965bb | !hmaster1_p & !v996587;
assign v97392c = hmaster1_p & v97392b | !hmaster1_p & !v9738be;
assign v985576 = busreq_p & v84563c | !busreq_p & !v985575;
assign v9d26eb = hmaster0_p & v9d26df | !hmaster0_p & v84563c;
assign v9adc95 = hbusreq1_p & v84563c | !hbusreq1_p & v9adc94;
assign v9ed4a0 = hmaster1_p & v9ed49b | !hmaster1_p & v9ed49f;
assign v9854e7 = hlock0_p & v9854e5 | !hlock0_p & v9854e6;
assign v973915 = hmaster1_p & v973907 | !hmaster1_p & v9738c0;
assign v8e79ce = hmaster1_p & v8e79cd | !hmaster1_p & v8e799f;
assign v973938 = hmaster0_p & v97388f | !hmaster0_p & v97388e;
assign v8c116a = hmaster0_p & v8c113a | !hmaster0_p & !v8c114c;
assign v9d2779 = hbusreq0_p & v9d274d | !hbusreq0_p & v9d2778;
assign v9bae93 = hbusreq1 & a153d1 | !hbusreq1 & !v9bae92;
assign v9adc19 = hmaster1_p & v9adc17 | !hmaster1_p & v9adc18;
assign v9ed480 = hburst0 & a153d0 | !hburst0 & v9ed47f;
assign v999986 = hmaster0_p & v9baf55 | !hmaster0_p & v9baf72;
assign v9b40dc = jx2_p & v9b40db | !jx2_p & v9b40cd;
assign v98550e = hmaster1_p & v985509 | !hmaster1_p & v9854dd;
assign v9b40c5 = hmaster1_p & v845660 | !hmaster1_p & v9b40c4;
assign v9d2696 = hbusreq1_p & v9d2695 | !hbusreq1_p & v845647;
assign v9adcf2 = decide_p & v9adc8d | !decide_p & v9adcf1;
assign v973986 = hmaster1_p & v973985 | !hmaster1_p & v97389c;
assign v9adc4c = hbusreq1_p & v9adc4a | !hbusreq1_p & v9adc4b;
assign v9d26e3 = hmaster1_p & v9d26e2 | !hmaster1_p & !v9d2671;
assign v9adc34 = stateG10_1_p & v9adc1f | !stateG10_1_p & !v9adc20;
assign v9baf04 = hmastlock_p & v9baf03 | !hmastlock_p & !v973884;
assign v9738b4 = hmaster1_p & v9738b0 | !hmaster1_p & v9738ad;
assign v9965c1 = hmaster0_p & v9adc35 | !hmaster0_p & v996552;
assign v9d268b = hmastlock_p & v9ed4a8 | !hmastlock_p & !v84563c;
assign v9855eb = hmaster1_p & v9855e6 | !hmaster1_p & v9855a2;
assign v98549f = locked_p & v98549e | !locked_p & !v84563c;
assign v99996f = hbusreq0_p & v99996e | !hbusreq0_p & !v84563c;
assign v9854ea = hburst0_p & v8ea7e3 | !hburst0_p & v9854e9;
assign v8ea87a = hbusreq2_p & v8ea844 | !hbusreq2_p & v8ea879;
assign v9baf0b = hburst0 & v84563c | !hburst0 & v9baf0a;
assign v9a6a99 = hmaster0_p & v84563c | !hmaster0_p & v9a6a98;
assign v9d26aa = busreq_p & v9d26a7 | !busreq_p & !v9d26a9;
assign v9d27ad = hmaster1_p & v9d27aa | !hmaster1_p & !v9d2673;
assign v9adcee = hmaster1_p & v9adced | !hmaster1_p & v9adcba;
assign v9adbed = hmastlock_p & v8543f4 | !hmastlock_p & !v84563c;
assign v8ea905 = hbusreq0_p & v8ea881 | !hbusreq0_p & v8ea904;
assign v985534 = hbusreq0_p & v985533 | !hbusreq0_p & v9854b6;
assign v984e6c = stateG2_p & v84563c | !stateG2_p & v984e6b;
assign v98559d = hgrant0_p & v985596 | !hgrant0_p & v98559c;
assign v9965c6 = decide_p & v9965c0 | !decide_p & v9965c5;
assign v9738d9 = hmaster1_p & v9738cd | !hmaster1_p & !v9738d8;
assign v9d2729 = hbusreq0_p & v9d2728 | !hbusreq0_p & v9d267e;
assign v973a1e = decide_p & v9739f9 | !decide_p & v973a1d;
assign v9ed4dd = hmaster1_p & v9ed4db | !hmaster1_p & v9ed478;
assign v9adcd4 = hready_p & v9adcd2 | !hready_p & v9adcd3;
assign v8c20bb = hmaster1_p & v845656 | !hmaster1_p & !v8c20ba;
assign v99659c = hbusreq1_p & v996599 | !hbusreq1_p & !v99659b;
assign v8ea889 = hmaster0_p & v8ea888 | !hmaster0_p & v8ea822;
assign v8ea936 = decide_p & v8ea7ee | !decide_p & v8ea935;
assign v8ea830 = hgrant0_p & v8ea81f | !hgrant0_p & v8ea82f;
assign v8c20cf = hgrant0_p & v8c20ca | !hgrant0_p & v8c20ce;
assign v984f25 = hmaster1_p & v84563c | !hmaster1_p & !v984f24;
assign v9d26bb = hbusreq0 & v9d26b8 | !hbusreq0 & v9d26ba;
assign v8ea846 = decide_p & v8ea845 | !decide_p & v8ea7e8;
assign v9a6ad9 = hready_p & v9a6ad3 | !hready_p & v9a6ad8;
assign v984f41 = hmaster1_p & v984f3f | !hmaster1_p & v984f40;
assign v99655c = hmaster0_p & v996559 | !hmaster0_p & v996552;
assign v8c1147 = hbusreq1_p & v8c1146 | !hbusreq1_p & !v84563c;
assign v9965c8 = hmaster1_p & v9965c7 | !hmaster1_p & v996597;
assign v8ea83a = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea839;
assign v9adc7c = hmaster0_p & v9adc79 | !hmaster0_p & !v9adc75;
assign v8ea8b8 = hmaster0_p & v8ea888 | !hmaster0_p & v8ea82c;
assign v8ea81d = hmaster0_p & v8ea7f1 | !hmaster0_p & v8ea81c;
    initial begin
  hready_p = 0;
  hbusreq0_p = 0;
  hlock0_p = 0;
  hbusreq1_p = 0;
  hlock1_p = 0;
  hbusreq2_p = 0;
  hlock2_p = 0;
  hburst0_p = 0;
  hburst1_p = 0;
  hmaster0_p = 0;
  hmaster1_p = 0;
  hmastlock_p = 0;
  start_p = 1;
  decide_p = 1;
  locked_p = 0;
  hgrant0_p = 1;
  hgrant1_p = 0;
  hgrant2_p = 0;
  busreq_p = 0;
  stateA1_p = 0;
  stateG2_p = 0;
  stateG3_0_p = 0;
  stateG3_1_p = 0;
  stateG3_2_p = 0;
  stateG10_1_p = 0;
  stateG10_2_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  hready_p = hready;
  hbusreq0_p = hbusreq0;
  hlock0_p = hlock0;
  hbusreq1_p = hbusreq1;
  hlock1_p = hlock1;
  hbusreq2_p = hbusreq2;
  hlock2_p = hlock2;
  hburst0_p = hburst0;
  hburst1_p = hburst1;
  hmaster0_p = hmaster0;
  hmaster1_p = hmaster1;
  hmastlock_p = hmastlock;
  start_p = start;
  decide_p = decide;
  locked_p = locked;
  hgrant0_p = hgrant0;
  hgrant1_p = hgrant1;
  hgrant2_p = hgrant2;
  busreq_p = busreq;
  stateA1_p = stateA1;
  stateG2_p = stateG2;
  stateG3_0_p = stateG3_0;
  stateG3_1_p = stateG3_1;
  stateG3_2_p = stateG3_2;
  stateG10_1_p = stateG10_1;
  stateG10_2_p = stateG10_2;
  jx0_p = jx0;
  jx1_p = jx1;
  jx2_p = jx2;
    end
endmodule

