module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, StoB_REQ4_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoS_ACK4_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, SLC2_n, jx0_n, jx1_n, jx2_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844f9b;
  wire v86ac9b;
  wire v868129;
  wire v8ca8d6;
  wire v8b69c5;
  wire v8caae9;
  wire v8cab56;
  wire v8caab4;
  wire v85f35c;
  wire v8cacd5;
  wire v868e55;
  wire v8caa61;
  wire v8c9805;
  wire v85cdad;
  wire v8cab70;
  wire v86b70b;
  wire v844f97;
  wire v8450db;
  wire v8caa15;
  wire v86113b;
  wire v8c9bb8;
  wire v8c9b72;
  wire v844f99;
  wire v8caac6;
  wire v85d86f;
  wire v85b5d1;
  wire v861d1f;
  wire v844f9d;
  wire v8c973b;
  wire v867bc5;
  wire v862264;
  wire v8cab3d;
  wire v86b132;
  wire v86ab8a;
  wire v8617fa;
  wire v86d276;
  wire v8caaf5;
  wire v8ca9c7;
  wire v8678e6;
  wire v865dbb;
  wire v8ca7a9;
  wire v85da17;
  wire v86490e;
  wire v8cacf4;
  wire v86b72d;
  wire v8caa6e;
  wire v869631;
  wire v8c9a7e;
  wire v8682bd;
  wire v8647c0;
  wire v8cac0d;
  wire v8cac49;
  wire v85e7b6;
  wire v868c92;
  wire v85e045;
  wire v85e6b9;
  wire v85d4df;
  wire v8cab0a;
  wire v85a021;
  wire v8caa3f;
  wire v8ca5f4;
  wire v869e27;
  wire v8caaa8;
  wire v86b436;
  wire v86b111;
  wire v8675a9;
  wire v8cabbb;
  wire v86d7c8;
  wire v8621d8;
  wire v8ca8b1;
  wire v85e1cc;
  wire v8ca1f2;
  wire v85e6c3;
  wire v8cab47;
  wire v8c9eb5;
  wire v8c9ce7;
  wire v86b7fd;
  wire v868bb5;
  wire v86d5fc;
  wire v8caaad;
  wire v856f8c;
  wire v865012;
  wire v868ccd;
  wire v85f2a4;
  wire v8698fa;
  wire v8675fc;
  wire v86a7af;
  wire v86b862;
  wire v867ba8;
  wire v87131b;
  wire v869065;
  wire v85e84a;
  wire v86665f;
  wire v8caace;
  wire v867508;
  wire v869dc6;
  wire v8cabdf;
  wire v8caa4d;
  wire v860d6f;
  wire v8caa5d;
  wire v8674b4;
  wire v86ac5d;
  wire v86989e;
  wire v86c5c8;
  wire v8674af;
  wire v86a56e;
  wire v861ea1;
  wire v86143d;
  wire v85d6d7;
  wire v86d5ab;
  wire v8666cf;
  wire v865f9a;
  wire v868402;
  wire v861809;
  wire v89af9c;
  wire v85e185;
  wire v8cacc5;
  wire v8cab9c;
  wire v8caa26;
  wire v868363;
  wire v8cab04;
  wire v85d7eb;
  wire v868905;
  wire v862fc7;
  wire v8c9a6e;
  wire v894074;
  wire v8cad04;
  wire v86b75f;
  wire v8cacdb;
  wire v85db7d;
  wire v8cac07;
  wire v86b74a;
  wire v8ca354;
  wire v8cac02;
  wire v861379;
  wire v8660a4;
  wire v8cac82;
  wire v85e922;
  wire v8cac85;
  wire v861494;
  wire v8caa52;
  wire v85e2e7;
  wire v8678af;
  wire v85164d;
  wire v8712d5;
  wire v8c9c7c;
  wire v867769;
  wire v86b485;
  wire v8ca3c3;
  wire v8caaab;
  wire v85de38;
  wire v86bae1;
  wire v8caa87;
  wire v869d71;
  wire v85e310;
  wire v8c9e09;
  wire v8cabde;
  wire v867417;
  wire v85d22b;
  wire v85f380;
  wire v86188b;
  wire v86908e;
  wire v86c5ef;
  wire v8660b8;
  wire v8cab88;
  wire v8667cc;
  wire v8ca9db;
  wire v8cac96;
  wire v8cab77;
  wire v85fb9d;
  wire v86ba71;
  wire v86863b;
  wire v86540f;
  wire v85f3a3;
  wire v85f2ab;
  wire v8696ce;
  wire v8cabe8;
  wire v860bf2;
  wire v8ca648;
  wire v88589b;
  wire v86d2f5;
  wire v861166;
  wire v866810;
  wire v866d6c;
  wire v85d30e;
  wire v86d7ce;
  wire v8caaf1;
  wire v8caa86;
  wire v86a8e7;
  wire v861525;
  wire v86117f;
  wire v8cab33;
  wire v85e3ea;
  wire v85e1f9;
  wire v861dac;
  wire v8caaca;
  wire v8cacdc;
  wire v8cab75;
  wire v85e544;
  wire v86a7da;
  wire v8b2a29;
  wire v844fab;
  wire v857ca8;
  wire v868fc7;
  wire v86889a;
  wire v85d43c;
  wire v86d3cb;
  wire v8c9917;
  wire v8cab3e;
  wire v8689a5;
  wire v860af3;
  wire v860ea5;
  wire v8caadb;
  wire v8cac80;
  wire v861d51;
  wire v86889b;
  wire v8668d6;
  wire v8cac4a;
  wire v869a67;
  wire v869dc8;
  wire v85df95;
  wire v8696e7;
  wire v8ca9d3;
  wire v86116b;
  wire v860a57;
  wire v860b28;
  wire v8658ac;
  wire v8caaed;
  wire v8c9aa6;
  wire v866540;
  wire v8cac98;
  wire v8c9df0;
  wire v8612e7;
  wire v8cab7c;
  wire v8697b7;
  wire v86a61f;
  wire v8ca018;
  wire v86840f;
  wire v85d881;
  wire v862bd2;
  wire v86af9f;
  wire v866fa1;
  wire v85de90;
  wire v864144;
  wire v86a66f;
  wire v8cacad;
  wire v8679a8;
  wire v85ac07;
  wire v86d7d4;
  wire v87132e;
  wire v866860;
  wire v86d2a8;
  wire v8caaff;
  wire v85310f;
  wire v8caa58;
  wire v8caca1;
  wire v86a799;
  wire v8cac0c;
  wire v85b56a;
  wire v8caa41;
  wire v86918c;
  wire v865f9e;
  wire v8cac21;
  wire v8cac0a;
  wire v8cac9c;
  wire v85e11a;
  wire v8712ee;
  wire v8660c6;
  wire v8594af;
  wire v8b2a28;
  wire v8caa7c;
  wire v86d147;
  wire v861df7;
  wire v8caa00;
  wire v8c9aac;
  wire v8cac63;
  wire v869ece;
  wire v866af0;
  wire v865dfa;
  wire v89af2b;
  wire v8cab36;
  wire v865811;
  wire v86d805;
  wire v8caa83;
  wire v861171;
  wire v8cace6;
  wire v86a611;
  wire v8cac16;
  wire v85da2b;
  wire v8c9dd6;
  wire v8ca5e2;
  wire v8ca126;
  wire v85dc69;
  wire v85deba;
  wire v85dc07;
  wire v85db6f;
  wire v85e8c1;
  wire v8640bb;
  wire v85309b;
  wire v8caa89;
  wire v866ee5;
  wire v85e4b6;
  wire v85e3ec;
  wire v8ca9fd;
  wire v8ca9cb;
  wire v8ca055;
  wire v869112;
  wire v86817a;
  wire v8caa0d;
  wire v8ca737;
  wire v86961e;
  wire v867cb8;
  wire v8cac77;
  wire v863e15;
  wire v8cab97;
  wire v8caade;
  wire v8ca0bd;
  wire v8cab0e;
  wire v86538c;
  wire v8c7acf;
  wire v8cabb7;
  wire v8cac53;
  wire v867b84;
  wire v86b348;
  wire v866013;
  wire v86d6f9;
  wire v8c9aca;
  wire v85de29;
  wire v865936;
  wire v8ca17e;
  wire v867e4a;
  wire v89c737;
  wire v85e046;
  wire v868830;
  wire v86c57f;
  wire v8683f7;
  wire v85e24b;
  wire v8caa2e;
  wire v8a7515;
  wire v844f9f;
  wire v8452cf;
  wire v869b57;
  wire v8cacd0;
  wire v8cabe4;
  wire v844f9c;
  wire v8ca9e9;
  wire v85e12e;
  wire v8c9e5e;
  wire v85f4e5;
  wire v844f9e;
  wire v861ecc;
  wire v86add5;
  wire v85e337;
  wire v8ca0ab;
  wire v844f95;
  wire v8cab4b;
  wire v8cab6e;
  wire v85d3a1;
  wire v8ca9cd;
  wire v8613f4;
  wire v86d0cd;
  wire v8ca246;
  wire v864a62;
  wire v861be5;
  wire v8caa55;
  wire v8caad9;
  wire v86d05a;
  wire v890c4a;
  wire v867be8;
  wire v866357;
  wire v85f4c4;
  wire v866b1d;
  wire v8cab4e;
  wire v868d0a;
  wire v8b69ca;
  wire v86d23a;
  wire v8c9a79;
  wire v8caa02;
  wire v86267d;
  wire v858cb9;
  wire v8cab15;
  wire v85e8ff;
  wire v8caa44;
  wire v8cac3a;
  wire v8cab2b;
  wire v8cab87;
  wire v869448;
  wire v866940;
  wire v866b27;
  wire v86652d;
  wire v866e01;
  wire v86d411;
  wire v86830a;
  wire v860c87;
  wire v8caa39;
  wire v8cac93;
  wire v85e03e;
  wire v8cac5b;
  wire v85a2c9;
  wire v8c9d2e;
  wire v8c8cdb;
  wire v868282;
  wire v86859e;
  wire v85f4ff;
  wire v8650ba;
  wire v869a08;
  wire v865bb1;
  wire v8648c8;
  wire v85e18e;
  wire v8caad8;
  wire v86adad;
  wire v88656b;
  wire v8cace2;
  wire v8607fe;
  wire v861b86;
  wire v868c7d;
  wire v86822b;
  wire v8c9db1;
  wire v868317;
  wire v86909b;
  wire v8c9af8;
  wire v869419;
  wire v8ca441;
  wire v86b9c5;
  wire v865bb9;
  wire v86674c;
  wire v8cacb9;
  wire v860bef;
  wire v866d0b;
  wire v860a37;
  wire v852479;
  wire v8cacb0;
  wire v8692f8;
  wire v866326;
  wire v8cab12;
  wire v861c0f;
  wire v8ca7a6;
  wire v869361;
  wire v861908;
  wire v8c9a1b;
  wire v89b010;
  wire v8caa43;
  wire v86c73b;
  wire v86d2fa;
  wire v8c9be8;
  wire v8cab01;
  wire v85daff;
  wire v85f516;
  wire v8caa8b;
  wire v8cad66;
  wire v8cacd2;
  wire v86685a;
  wire v8660b6;
  wire v8caae1;
  wire v85e35c;
  wire v8cace5;
  wire v866420;
  wire v8caa3a;
  wire v85d91a;
  wire v86b9ab;
  wire v868403;
  wire v86d786;
  wire v8658e5;
  wire v85e484;
  wire v86a6a1;
  wire v86a710;
  wire v865efb;
  wire v868d58;
  wire v86d58d;
  wire v85df63;
  wire v868377;
  wire v86522b;
  wire v8678d9;
  wire v89af47;
  wire v85d53b;
  wire v85d90c;
  wire v8ca686;
  wire v868cbe;
  wire v86ae59;
  wire v8caa33;
  wire v861279;
  wire v8ca742;
  wire v8caa14;
  wire v85e5c6;
  wire v85e81e;
  wire v86217d;
  wire v85e87a;
  wire v8614bb;
  wire v8cac8f;
  wire v85e164;
  wire v860cd1;
  wire v8cabfd;
  wire v86b1d8;
  wire v869b48;
  wire v85e0d5;
  wire v8ca71c;
  wire v8caa90;
  wire v8cac4e;
  wire v865427;
  wire v86aec5;
  wire v86a953;
  wire v8cab59;
  wire v86ae3e;
  wire v868ba7;
  wire v86d0ec;
  wire v861889;
  wire v86b3cd;
  wire v86d322;
  wire v8ca615;
  wire v844fbb;
  wire v844fa5;
  wire v86b6e3;
  wire v85d1fb;
  wire v86631f;
  wire v8c9cac;
  wire v8ca303;
  wire v85e09a;
  wire v8691f9;
  wire v8ca19f;
  wire v8cab8f;
  wire v866bb9;
  wire v8caa7e;
  wire v8caca3;
  wire v8caafc;
  wire v8cab8e;
  wire v8c9c59;
  wire v85d4e0;
  wire v860d7c;
  wire v89409f;
  wire v8a6050;
  wire v8664cd;
  wire v85d86a;
  wire v8ca21b;
  wire v86d5c8;
  wire v861f69;
  wire v8caa57;
  wire v860c8a;
  wire v8cac86;
  wire v861fb9;
  wire v8cab63;
  wire v863955;
  wire v8cac99;
  wire v8ca9ef;
  wire v86d753;
  wire v8caa62;
  wire v8ca1e1;
  wire v85c6d8;
  wire v8620d1;
  wire v85dfad;
  wire v8c95d7;
  wire v8caa17;
  wire v85f557;
  wire v8cab1a;
  wire v8588a0;
  wire v8cab90;
  wire v8cabf5;
  wire v865859;
  wire v8ca9eb;
  wire v8679ab;
  wire v8ca61e;
  wire v86d101;
  wire v8ca695;
  wire v8caa29;
  wire v8ca4e9;
  wire v85ceb3;
  wire v8ca172;
  wire v85d3d5;
  wire v8ca472;
  wire v8cacd1;
  wire v8ca9c9;
  wire v855346;
  wire v8cac69;
  wire v8caa36;
  wire v8cac10;
  wire v85e4c8;
  wire v8940ad;
  wire v866610;
  wire v865da0;
  wire v8ca399;
  wire v8ca2a1;
  wire v867763;
  wire v85ce75;
  wire v868fd6;
  wire v8a6000;
  wire v844fad;
  wire v868c2a;
  wire v86754b;
  wire v8682f7;
  wire v869990;
  wire v8caa8f;
  wire v8c9cad;
  wire v8649c5;
  wire v8cab74;
  wire v8ca3cb;
  wire v8c9c9f;
  wire v8cac7e;
  wire v8caa3c;
  wire v866d4f;
  wire v8c9607;
  wire v8ca9e8;
  wire v88cf5c;
  wire v8caaf0;
  wire v85cec5;
  wire v866c98;
  wire v89407e;
  wire v8ca9e0;
  wire v86a6ed;
  wire v8c7b53;
  wire v86770a;
  wire v89c779;
  wire v8cab19;
  wire v8c9811;
  wire v86653c;
  wire v867220;
  wire v8cac6d;
  wire v8ca693;
  wire v85e228;
  wire v8c9bb0;
  wire v85e85f;
  wire v8b31ca;
  wire v86d231;
  wire v85ce98;
  wire v8cacd8;
  wire v8662c3;
  wire v8b69a2;
  wire v860ec7;
  wire v8cacd3;
  wire v866964;
  wire v8794d1;
  wire v86294e;
  wire v866880;
  wire v866655;
  wire v8601bc;
  wire v86a60b;
  wire v8c9626;
  wire v86b3a2;
  wire v8cacca;
  wire v85dbc1;
  wire v8858bf;
  wire v8692e8;
  wire v85d6e1;
  wire v85769e;
  wire v866138;
  wire v8caa71;
  wire v8660ec;
  wire v8cac79;
  wire v8c9d37;
  wire v860e50;
  wire v8650b2;
  wire v8cab71;
  wire v8ca56d;
  wire v8cac46;
  wire v8cab94;
  wire v8cab9f;
  wire v86265a;
  wire v8cab84;
  wire v867780;
  wire v8cab49;
  wire v86c833;
  wire v86d3d9;
  wire v8cab08;
  wire v8cac41;
  wire v8cace0;
  wire v8c9ace;
  wire v8cac81;
  wire v85e297;
  wire v8ca2c0;
  wire v85d906;
  wire v8caae4;
  wire v8ca9a6;
  wire v85f3d3;
  wire v8671ac;
  wire v869baf;
  wire v8654fc;
  wire v869ca4;
  wire v8c9ed8;
  wire v8649c1;
  wire v868ae9;
  wire v8c9bd1;
  wire v86b02f;
  wire v86d814;
  wire v86191e;
  wire v8cac54;
  wire v86b298;
  wire v8cac1f;
  wire v8ca153;
  wire v865295;
  wire v8ca154;
  wire v85e4f2;
  wire v862031;
  wire v861d50;
  wire v85e5ff;
  wire v8cac28;
  wire v860b19;
  wire v8c9bbf;
  wire v863449;
  wire v8637cb;
  wire v8cace7;
  wire v862e4a;
  wire v88656a;
  wire v86c701;
  wire v861db7;
  wire v865da5;
  wire v865b89;
  wire v8663ef;
  wire v8cac9f;
  wire v8c9dae;
  wire v8cab1d;
  wire v85dac9;
  wire v8cab37;
  wire v8683f9;
  wire v8cab07;
  wire v86b05b;
  wire v85dee9;
  wire v8680fe;
  wire v8ca089;
  wire v85d5c3;
  wire v86adcf;
  wire v85b1cb;
  wire v865fe1;
  wire v8ca9f7;
  wire v86b125;
  wire v8caa56;
  wire v86607a;
  wire v86b7cd;
  wire v8caa5a;
  wire v85e715;
  wire v8677dc;
  wire v868b0b;
  wire v8ca44e;
  wire v86753c;
  wire v8caccc;
  wire v8ca9d5;
  wire v8cabcd;
  wire v8cac22;
  wire v867ef1;
  wire v859567;
  wire v8666db;
  wire v864a04;
  wire v8caa11;
  wire v8698ed;
  wire v865ff9;
  wire v86d329;
  wire v86d6a1;
  wire v8ca9c3;
  wire v89c777;
  wire v8a5ffe;
  wire v8c9f2a;
  wire v8c97e3;
  wire v8c9aea;
  wire v8697c8;
  wire v8c9b09;
  wire v86b9e6;
  wire v8677e5;
  wire v8679eb;
  wire v86a618;
  wire v86d092;
  wire v86d61d;
  wire v8c9b51;
  wire v8caa67;
  wire v8cacdd;
  wire v8cabb5;
  wire v868b10;
  wire v85d6cf;
  wire v8c9f67;
  wire v8c9e00;
  wire v865cd4;
  wire v8cab9a;
  wire v8c9753;
  wire v8caca0;
  wire v8ca9ea;
  wire v8cac03;
  wire v8ca374;
  wire v86150f;
  wire v85cef2;
  wire v85ddf2;
  wire v8c9b86;
  wire v8688ca;
  wire v86d803;
  wire v85f3f5;
  wire v85cdf0;
  wire v8664b1;
  wire v8caba0;
  wire v8cabcc;
  wire v8caa1a;
  wire v85e30e;
  wire v86560f;
  wire v865321;
  wire v8caa8a;
  wire v86223f;
  wire v869ddd;
  wire v85e143;
  wire v8c7aa7;
  wire v866997;
  wire v8cabcb;
  wire v8caab0;
  wire v866d8b;
  wire v8612ab;
  wire v8a74c0;
  wire v85d9cf;
  wire v8cac42;
  wire v8ca9be;
  wire v85e95a;
  wire v867844;
  wire v85f749;
  wire v87947b;
  wire v8c7b49;
  wire v8c9942;
  wire v8cab6c;
  wire v86b05c;
  wire v8674bb;
  wire v8613c9;
  wire v8cab5d;
  wire v8cac33;
  wire v862256;
  wire v85e733;
  wire v8cacb5;
  wire v8cabed;
  wire v8cac8e;
  wire v867b2b;
  wire v862180;
  wire v8ca753;
  wire v86864b;
  wire v86d81c;
  wire v85e249;
  wire v86b711;
  wire v86a8b8;
  wire v85db64;
  wire v867a20;
  wire v8b317b;
  wire v8cac3d;
  wire v89c755;
  wire v8c9c75;
  wire v8cabe2;
  wire v8cabfe;
  wire v8cacff;
  wire v85dece;
  wire v8940e1;
  wire v8ca380;
  wire v8ca315;
  wire v86639e;
  wire v8ca9f0;
  wire v89b000;
  wire v8ca937;
  wire v865de8;
  wire v8caac1;
  wire v8661bc;
  wire v8622a3;
  wire v866d60;
  wire v8caaf8;
  wire v867080;
  wire v867a57;
  wire v862883;
  wire v861794;
  wire v8cabca;
  wire v8c9b26;
  wire v88d120;
  wire v8c0272;
  wire v861405;
  wire v85d81d;
  wire v86a905;
  wire v865960;
  wire v867957;
  wire v85f4e3;
  wire v866c71;
  wire v8cabea;
  wire v86b30e;
  wire v8c9e27;
  wire v86921b;
  wire v865319;
  wire v8caa37;
  wire v85d8fe;
  wire v86d602;
  wire v8b29f7;
  wire v864207;
  wire v861e9b;
  wire v8cac1d;
  wire v8cac71;
  wire v865707;
  wire v8b31a9;
  wire v85e833;
  wire v8cac51;
  wire v8ca5b3;
  wire v8ca9d0;
  wire v8cabbd;
  wire v866369;
  wire v860e09;
  wire v8610eb;
  wire v8692bc;
  wire v88d12d;
  wire v8cab5c;
  wire v8caab8;
  wire v86494d;
  wire v866d6a;
  wire v868b32;
  wire v85206c;
  wire v8b3161;
  wire v8cac7a;
  wire v88d132;
  wire v86c49c;
  wire v864ac7;
  wire v8caa1d;
  wire v85d34f;
  wire v8c9d60;
  wire v85f48d;
  wire v8caa76;
  wire v8cac23;
  wire v868f7d;
  wire v8b69b8;
  wire v86d647;
  wire v8ca8ca;
  wire v8cad5f;
  wire v8cac05;
  wire v85f521;
  wire v8ca7e1;
  wire v85ce31;
  wire v85cde5;
  wire v8cacdf;
  wire v8caa6b;
  wire v8c95e9;
  wire v86c854;
  wire v868dd2;
  wire v867abe;
  wire v894106;
  wire v85e69b;
  wire v85dee1;
  wire v8caa40;
  wire v844fa7;
  wire v8c9ce3;
  wire v85e110;
  wire v844fa9;
  wire v86b50c;
  wire v8ca9d4;
  wire v86593c;
  wire v85cdfc;
  wire v861bb6;
  wire v861374;
  wire v869147;
  wire v8a74b4;
  wire v86d775;
  wire v8cab06;
  wire v8696ea;
  wire v869e56;
  wire v8cac35;
  wire v866d1f;
  wire v8667fb;
  wire v864071;
  wire v8664d8;
  wire v867a34;
  wire v8caa01;
  wire v8cab55;
  wire v86a84a;
  wire v85d230;
  wire v86d061;
  wire v8cab7b;
  wire v85e2f3;
  wire v861fda;
  wire v8ca9ee;
  wire v85e8ee;
  wire v865fe6;
  wire v8ca553;
  wire v8cabf3;
  wire v85e8c7;
  wire v8641cf;
  wire v85e568;
  wire v860f28;
  wire v8cab3a;
  wire v8cacb4;
  wire v867e47;
  wire v8cabac;
  wire v8c9e60;
  wire v85dade;
  wire v8ca78f;
  wire v8ca313;
  wire v8c7b4e;
  wire v8a868e;
  wire v86349c;
  wire v8cabd7;
  wire v8caa9d;
  wire v867a28;
  wire v860ab6;
  wire v868cbc;
  wire v86ba19;
  wire v86afde;
  wire v8b69e1;
  wire v8caaef;
  wire v8ca23b;
  wire v8caac4;
  wire v868378;
  wire v8cad4e;
  wire v85e8cb;
  wire v85f7ba;
  wire v866b54;
  wire v86a607;
  wire v852625;
  wire v86a745;
  wire v8610ac;
  wire v8caba9;
  wire v8cac2d;
  wire v8a604c;
  wire v85d39c;
  wire v85d954;
  wire v8cac70;
  wire v85cdc2;
  wire v8caa21;
  wire v85e947;
  wire v865f35;
  wire v869b6e;
  wire v8cab17;
  wire v8ca357;
  wire v8cab72;
  wire v861fc9;
  wire v8c9b67;
  wire v8cac45;
  wire v8caaf3;
  wire v86ab5e;
  wire v8caa8c;
  wire v85ce85;
  wire v861856;
  wire v8682bf;
  wire v8cac76;
  wire v8cabb4;
  wire v8cabef;
  wire v8ca022;
  wire v8647a2;
  wire v8c95c7;
  wire v8cab03;
  wire v8cac6b;
  wire v8cacaf;
  wire v85e2ea;
  wire v85f4cf;
  wire v86752a;
  wire v85d9e0;
  wire v8caaa9;
  wire v8cac15;
  wire v85d221;
  wire v85e78a;
  wire v8caabc;
  wire v85e743;
  wire v868e01;
  wire v865f0e;
  wire v86c4e5;
  wire v86ba45;
  wire v8c9ea3;
  wire v861dcc;
  wire v85e6c0;
  wire v861c02;
  wire v866606;
  wire v85e569;
  wire v85dd97;
  wire v8c9dd4;
  wire v86a5ad;
  wire v875b43;
  wire v861b6c;
  wire v86a76c;
  wire v8cab44;
  wire v8caa5f;
  wire v8598f7;
  wire v8cab52;
  wire v864506;
  wire v861980;
  wire v8c9aee;
  wire v8699ec;
  wire v86b22a;
  wire v8cab8c;
  wire v866834;
  wire v85506c;
  wire v85dbdc;
  wire v86b5da;
  wire v85db20;
  wire v8c97df;
  wire v8691a7;
  wire v86589e;
  wire v85d73d;
  wire v868569;
  wire v869197;
  wire v8ca345;
  wire v85de3b;
  wire v85e1cb;
  wire v88d14f;
  wire v8caca5;
  wire v866205;
  wire v8cac0f;
  wire v85f39d;
  wire v86a660;
  wire v89b002;
  wire v85e2d7;
  wire v869284;
  wire v86d813;
  wire v8661e2;
  wire v8cabe1;
  wire v89afd9;
  wire v8ca009;
  wire v8cab89;
  wire v86a6c6;
  wire v8caad2;
  wire v8cab26;
  wire v8654cb;
  wire v8ca9d8;
  wire v8a74a8;
  wire v86707f;
  wire v865787;
  wire v860aed;
  wire v8caadc;
  wire v86d25f;
  wire v8c95d0;
  wire v85dbee;
  wire v85d75d;
  wire v8647c1;
  wire v8cab6b;
  wire v8ca9af;
  wire v8cab29;
  wire v85d8cc;
  wire v86b725;
  wire v8c9b2e;
  wire v8b3195;
  wire v8ca9e6;
  wire v88d17c;
  wire v8caab9;
  wire v8caa66;
  wire v867d26;
  wire v89afeb;
  wire v8cacba;
  wire v8caa74;
  wire v8619cf;
  wire v8ca8b9;
  wire v86aebe;
  wire v8cab57;
  wire v8ca2af;
  wire v8c9d1a;
  wire v8cacce;
  wire v869060;
  wire v85e813;
  wire v86b7b7;
  wire v865cb0;
  wire v86d130;
  wire v8caa48;
  wire v857888;
  wire v8667bd;
  wire v86b4d5;
  wire v8cabc0;
  wire v86d1b3;
  wire v8caba4;
  wire v86114b;
  wire v8cac5e;
  wire v85dfa3;
  wire v86882a;
  wire v866d97;
  wire v8cab02;
  wire v868936;
  wire v8caae5;
  wire v8cac2a;
  wire v8caa91;
  wire v86550b;
  wire v869dae;
  wire v8674f7;
  wire v8cab25;
  wire v8ca32a;
  wire v861d5f;
  wire v8c984a;
  wire v85d1d4;
  wire v8cabeb;
  wire v8cac09;
  wire v8667f6;
  wire v8caa81;
  wire v8caa79;
  wire v868467;
  wire v861aba;
  wire v866aae;
  wire v8609a9;
  wire v85ce37;
  wire v8693db;
  wire v8ca9f4;
  wire v8c9f14;
  wire v860d73;
  wire v8cacc8;
  wire v8ca2fd;
  wire v861436;
  wire v8cac00;
  wire v864bf9;
  wire v85e88d;
  wire v85e4fc;
  wire v869f33;
  wire v86202e;
  wire v8caafd;
  wire v85d772;
  wire v864b34;
  wire v8cab5a;
  wire v85e3f3;
  wire v8c9712;
  wire v8b31d3;
  wire v866c03;
  wire v8c9cae;
  wire v86925d;
  wire v8647c8;
  wire v8cab42;
  wire v85e138;
  wire v867010;
  wire v868f72;
  wire v8ca84f;
  wire v868120;
  wire v8667ba;
  wire v869992;
  wire v8caa1e;
  wire v8cacd7;
  wire v8c9cbc;
  wire v86b7bb;
  wire v85f3fa;
  wire v86c801;
  wire v8caa9b;
  wire v89affe;
  wire v86888b;
  wire v8caa9a;
  wire v867a75;
  wire v86b2c2;
  wire v85cdba;
  wire v8caaf7;
  wire v8cac29;
  wire v866529;
  wire v8cabf0;
  wire v86b06e;
  wire v86c581;
  wire v8ca9f5;
  wire v8c9733;
  wire v8ca6b5;
  wire v8cacab;
  wire v84505f;
  wire v85d97a;
  wire v8ca41e;
  wire v8cac39;
  wire v8c9890;
  wire v8cac6a;
  wire v871300;
  wire v8c9f9a;
  wire v8940a7;
  wire v865d47;
  wire v861d21;
  wire v8858c9;
  wire v8cac7c;
  wire v85c5d4;
  wire v864b72;
  wire v8caa18;
  wire v8cab9b;
  wire v85e61f;
  wire v8cabd8;
  wire v8691f2;
  wire v8caa20;
  wire v86ac7c;
  wire v867edf;
  wire v864ad9;
  wire v866cf1;
  wire v8b69a7;
  wire v8c7b0b;
  wire v8caca2;
  wire v861998;
  wire v8cac72;
  wire v85e55a;
  wire v8cac32;
  wire v866456;
  wire v8663d1;
  wire v8caa75;
  wire v86ba15;
  wire v86b838;
  wire v8caad7;
  wire v8ca349;
  wire v85d173;
  wire v8cabe6;
  wire v85dbcd;
  wire v867166;
  wire v8ca849;
  wire v8cab2d;
  wire v86912f;
  wire v86d378;
  wire v86908c;
  wire v8940fd;
  wire v856fa3;
  wire v8a74fd;
  wire v8cabc7;
  wire v894103;
  wire v85d23a;
  wire v8cac5c;
  wire v86757f;
  wire v8ca3c8;
  wire v8cab21;
  wire v86b799;
  wire v8633e4;
  wire v85e351;
  wire v85d232;
  wire v8caa7d;
  wire v866ad5;
  wire v86a8cf;
  wire v8cab32;
  wire v861bd6;
  wire v862012;
  wire v864dbb;
  wire v85cd74;
  wire v8cac30;
  wire v85ce9c;
  wire v8ca9fb;
  wire v85e65a;
  wire v860a0f;
  wire v865d58;
  wire v8cabc1;
  wire v8ca0f9;
  wire v862305;
  wire v8cac9b;
  wire v8c9ec8;
  wire v8cabd0;
  wire v85e5ed;
  wire v8caafb;
  wire v85d485;
  wire v8cac8c;
  wire v86d7f2;
  wire v86c517;
  wire v86d2a0;
  wire v8ca6af;
  wire v8cac12;
  wire v8cadb0;
  wire v8caacc;
  wire v8ca440;
  wire v866632;
  wire v868edb;
  wire v8c9e31;
  wire v86a5b6;
  wire v8cac1a;
  wire v867b20;
  wire v8ca701;
  wire v86884e;
  wire v85e491;
  wire v8cac13;
  wire v8697ea;
  wire v861522;
  wire v86837b;
  wire v862200;
  wire v8693ab;
  wire v8690d8;
  wire v869526;
  wire v8691f7;
  wire v8cacbd;
  wire v8b2a14;
  wire v8b69cf;
  wire v857c24;
  wire v867507;
  wire v865791;
  wire v8651a5;
  wire v8caa0a;
  wire v85c630;
  wire v8cabd2;
  wire v8794af;
  wire v85cdd6;
  wire v8ca787;
  wire v8c7b59;
  wire v861882;
  wire v869497;
  wire v8c9ed1;
  wire v868fbe;
  wire v85bdd0;
  wire v8c9cbb;
  wire v86903b;
  wire v8cac11;
  wire v8caa1b;
  wire v8660d7;
  wire v8ca48a;
  wire v8cac43;
  wire v852627;
  wire v86d0bf;
  wire v8cab4c;
  wire v85c85e;
  wire v86797e;
  wire v868b0c;
  wire v868f18;
  wire v85da42;
  wire v85ce03;
  wire v8ca9fa;
  wire v86c524;
  wire v85e1fe;
  wire v8ca7ed;
  wire v8cab1c;
  wire v868bd4;
  wire v8cab6f;
  wire v8cab81;
  wire v85d985;
  wire v85c82e;
  wire v865edc;
  wire v8672bb;
  wire v8ca9ff;
  wire v867a99;
  wire v8caad3;
  wire v86b108;
  wire v8ca86e;
  wire v8cabff;
  wire v869653;
  wire v8c9b41;
  wire v862881;
  wire v8caaaa;
  wire v85c2e5;
  wire v8ca115;
  wire v86d43f;
  wire v8cabfc;
  wire v8c99d1;
  wire v8caad0;
  wire v85e183;
  wire v866d78;
  wire v8cacd6;
  wire v8caa06;
  wire v8caa45;
  wire v85e233;
  wire v85c534;
  wire v8cabf2;
  wire v8caa31;
  wire v85a4d3;
  wire v865bf0;
  wire v861e4f;
  wire v8671b5;
  wire v8c9d6e;
  wire v8cac66;
  wire v868626;
  wire v8ca300;
  wire v85d919;
  wire v867a8a;
  wire v8caa0f;
  wire v8679f8;
  wire v8667e9;
  wire v85d860;
  wire v8678d8;
  wire v86d402;
  wire v8c9a57;
  wire v8cad25;
  wire v8c9752;
  wire v85bb82;
  wire v86aff9;
  wire v8caa60;
  wire v86b786;
  wire v867319;
  wire v8caad4;
  wire v8caa2f;
  wire v8cac87;
  wire v8cabcf;
  wire v8caaae;
  wire v8c96e3;
  wire v8ca5f9;
  wire v866af3;
  wire v8673d4;
  wire v8685d8;
  wire v869922;
  wire v86a764;
  wire v8caa7f;
  wire v894033;
  wire v85e872;
  wire v85d80e;
  wire v8caba7;
  wire v85e6fc;
  wire v85f4ce;
  wire v867c81;
  wire v8ca98e;
  wire v85d750;
  wire v8cacbe;
  wire v86921e;
  wire v86816d;
  wire v8c97c4;
  wire v860b60;
  wire v8ca840;
  wire v8686e5;
  wire v869380;
  wire v861d36;
  wire v8caaec;
  wire v8cabc6;
  wire v8621d5;
  wire v8b3167;
  wire v8cac2e;
  wire v866c47;
  wire v86badb;
  wire v8940d7;
  wire v85d843;
  wire v85d880;
  wire v869251;
  wire v8cab05;
  wire v86af4a;
  wire v8ca295;
  wire v865036;
  wire v86b96c;
  wire v86c461;
  wire v8ca04b;
  wire v852940;
  wire v86981f;
  wire v85e63e;
  wire v867170;
  wire v868dd9;
  wire v8caa51;
  wire v8609fc;
  wire v861903;
  wire v8632cd;
  wire v8c963c;
  wire v86ade6;
  wire v8caac0;
  wire v8caa2b;
  wire v869ec7;
  wire v8653c0;
  wire v867551;
  wire v8cac5d;
  wire v85e95d;
  wire v85e2a3;
  wire v86d63a;
  wire v8cab14;
  wire v8cacb6;
  wire v8c9ef9;
  wire v86702e;
  wire v861774;
  wire v86621a;
  wire v861d73;
  wire v867cf7;
  wire v8599dd;
  wire v864050;
  wire v8794e5;
  wire v851272;
  wire v8452cd;
  wire v861c01;
  wire v8cac4b;
  wire v860a1c;
  wire v8cab2f;
  wire v8cacc6;
  wire v86922c;
  wire v8cacc7;
  wire v861290;
  wire v86608e;
  wire v8caac2;
  wire v8c9c26;
  wire v8cac06;
  wire v85d924;
  wire v867c96;
  wire v862321;
  wire v86ac23;
  wire v85d56c;
  wire v8b2a0d;
  wire v8ca9f3;
  wire v869259;
  wire v86d1e7;
  wire v8ca00c;
  wire v86900f;
  wire v866b6f;
  wire v8674ab;
  wire v875b45;
  wire v89afb5;
  wire v865507;
  wire v85da6a;
  wire v85e30d;
  wire v8c9fa7;
  wire v8ca9de;
  wire v85cf1e;
  wire v86890b;
  wire v864080;
  wire v867ed2;
  wire v8ca096;
  wire v85daa3;
  wire v85d28e;
  wire v8caad6;
  wire v86c702;
  wire v85d58f;
  wire v86d087;
  wire v869e35;
  wire v8ca014;
  wire v861f9e;
  wire v8caa53;
  wire v8612b9;
  wire v8cac0b;
  wire v868c4d;
  wire v8ca0b4;
  wire v8caa70;
  wire v8ca79e;
  wire v865c5c;
  wire v8caada;
  wire v85cebf;
  wire v86d136;
  wire v8ca9e2;
  wire v866ba0;
  wire v8ca6a1;
  wire v8cacc4;
  wire v85e4b1;
  wire v8c9681;
  wire v867697;
  wire v8cab39;
  wire v867cbe;
  wire v8caa08;
  wire v8caac9;
  wire v8cab9d;
  wire v8ca9e4;
  wire v861409;
  wire v8c977d;
  wire v85d451;
  wire v86789d;
  wire v865d4b;
  wire v8cac8d;
  wire v85deac;
  wire v86698a;
  wire v8ca3d4;
  wire v8caab6;
  wire v8c9696;
  wire v866015;
  wire v861266;
  wire v8cabe9;
  wire v867565;
  wire v85d448;
  wire v8ca9c1;
  wire v868f67;
  wire v8caacd;
  wire v85c6f5;
  wire v8caa4a;
  wire v8cacde;
  wire v8712d2;
  wire v8cab28;
  wire v8cad96;
  wire v8c9bd7;
  wire v86dae3;
  wire v8641a6;
  wire v8cab61;
  wire v8c9cc5;
  wire v866d9e;
  wire v85d7bc;
  wire v88d0f1;
  wire v86d74c;
  wire v867a22;
  wire v8cac08;
  wire v866a61;
  wire v8a749d;
  wire v856a93;
  wire v8cab6d;
  wire v8caad1;
  wire v866f76;
  wire v8caccf;
  wire v8ca9cf;
  wire v8cad54;
  wire v865a01;
  wire v8cab76;
  wire v855530;
  wire v8cab79;
  wire v86d557;
  wire v85a733;
  wire v85e2c9;
  wire v8cabec;
  wire v8cab16;
  wire v8cacaa;
  wire v8cac20;
  wire v865e2b;
  wire v86911f;
  wire v865f16;
  wire v85f3d4;
  wire v861905;
  wire v8ca9e3;
  wire v861e53;
  wire v866037;
  wire v8cac84;
  wire v861b4d;
  wire v85dda7;
  wire v861969;
  wire v8cab34;
  wire v866b78;
  wire v865404;
  wire v8c9bfc;
  wire v86d7e6;
  wire v86974a;
  wire v8651a3;
  wire v86b4f5;
  wire v8656ee;
  wire v865e4b;
  wire v8cac4f;
  wire v867c16;
  wire v8cac3e;
  wire v86b7d3;
  wire v85de99;
  wire v879471;
  wire v8ca196;
  wire v8680ed;
  wire v851793;
  wire v867f36;
  wire v86d390;
  wire v859cb4;
  wire v865230;
  wire v869b15;
  wire v866bf7;
  wire v8ca522;
  wire v879497;
  wire v866b4c;
  wire v8cac65;
  wire v8c9ff6;
  wire v8caa77;
  wire v85e224;
  wire v85d413;
  wire v8594ba;
  wire v8c9a18;
  wire v87133e;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg StoB_REQ4_p;
  input StoB_REQ4_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoS_ACK4_p;
  output BtoS_ACK4_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg SLC2_p;
  output SLC2_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  wire ENQ_n;
  wire SLC2_n;

assign v8940a7 = stateG7_1_p & v85d97a | !stateG7_1_p & v8c9f9a;
assign v8cab36 = BtoS_ACK1_p & v8cac4a | !BtoS_ACK1_p & v89af2b;
assign v86294e = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8794d1;
assign v8cacdf = EMPTY_p & v865319 | !EMPTY_p & v862031;
assign v8cabe2 = jx2_p & v866880 | !jx2_p & !v844f91;
assign v864a62 = EMPTY_p & v8ca246 | !EMPTY_p & !v844f91;
assign v864071 = ENQ_p & v844fbb | !ENQ_p & v8667fb;
assign v85e922 = BtoS_ACK0_p & v8cab3d | !BtoS_ACK0_p & v8cac82;
assign v8c9ea3 = FULL_p & v844f91 | !FULL_p & v85e743;
assign v8cab8f = stateG12_p & v8ca19f | !stateG12_p & v844f91;
assign v867166 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85dbcd;
assign v85e484 = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v8658e5;
assign v865936 = DEQ_p & v844f91 | !DEQ_p & v85de29;
assign v8caa00 = EMPTY_p & v86a66f | !EMPTY_p & v8594af;
assign v8ca840 = StoB_REQ2_p & v85d750 | !StoB_REQ2_p & v860b60;
assign v8cacb6 = EMPTY_p & v8c963c | !EMPTY_p & v8673d4;
assign v85f557 = StoB_REQ2_p & v863955 | !StoB_REQ2_p & !v8caa17;
assign v86822b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v868c7d;
assign v8cabcf = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85d860;
assign v8c9752 = jx2_p & v8cad25 | !jx2_p & v865edc;
assign v867220 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86653c;
assign v8cab5c = EMPTY_p & v8cacb5 | !EMPTY_p & !v88d12d;
assign v8647c8 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v86925d;
assign v844fad = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v8c9ed1 = jx2_p & v844f91 | !jx2_p & !v866940;
assign v85e6fc = jx0_p & v85bdd0 | !jx0_p & !v85d80e;
assign v8cac72 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v861998;
assign v8cab61 = EMPTY_p & v8cab9d | !EMPTY_p & !v8641a6;
assign v855346 = StoB_REQ0_p & v8ca472 | !StoB_REQ0_p & v8ca9c9;
assign v8caa55 = ENQ_p & v8cabe4 | !ENQ_p & v861be5;
assign v865da5 = jx2_p & v861db7 | !jx2_p & !v844f91;
assign v8c977d = jx2_p & v85cf1e | !jx2_p & v861409;
assign v861d36 = StoB_REQ1_p & v8ca840 | !StoB_REQ1_p & v869380;
assign v8cabef = jx2_p & v8cabb4 | !jx2_p & v8cab4b;
assign v8c9bb0 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8cab19;
assign v8698fa = jx2_p & v8caae9 | !jx2_p & v85f2a4;
assign v8680ed = DEQ_p & v8cabec | !DEQ_p & v8ca196;
assign v8cab06 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86d775;
assign v8caac9 = jx1_p & v85cf1e | !jx1_p & v8caa08;
assign v8caad7 = BtoS_ACK0_p & v8691f2 | !BtoS_ACK0_p & v86b838;
assign v8ca9ee = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v861fda;
assign v85daa3 = DEQ_p & v8ca096 | !DEQ_p & v85da6a;
assign v85f7ba = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e8cb;
assign v8cab42 = StoB_REQ0_p & v868569 | !StoB_REQ0_p & v8647c8;
assign v866860 = jx1_p & v87132e | !jx1_p & !v85de90;
assign v8674ab = BtoR_REQ1_p & v862321 | !BtoR_REQ1_p & v866b6f;
assign v8cabeb = jx0_p & v8c984a | !jx0_p & v85d1d4;
assign v8caca0 = FULL_p & v8cac54 | !FULL_p & !v8c9753;
assign v8c9e27 = jx2_p & v86b30e | !jx2_p & !v8cac6d;
assign v868ccd = BtoS_ACK0_p & v8c9805 | !BtoS_ACK0_p & v865012;
assign v85e8ff = StoB_REQ3_p & v861ecc | !StoB_REQ3_p & v844f9c;
assign v856f8c = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8caaad;
assign v866aae = FULL_p & v844f91 | !FULL_p & v8caa81;
assign v8caa71 = jx0_p & v85dbc1 | !jx0_p & v866138;
assign v85c82e = BtoS_ACK0_p & v8caa5a | !BtoS_ACK0_p & v85d985;
assign v8cac8c = EMPTY_p & v86b799 | !EMPTY_p & v85d485;
assign v869497 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v861882;
assign v85ce37 = DEQ_p & v8cab57 | !DEQ_p & v8609a9;
assign v861522 = jx2_p & v844f91 | !jx2_p & v86b50c;
assign v85e88d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v864bf9;
assign v86b7cd = jx1_p & v844f9b | !jx1_p & !v8cacca;
assign v868129 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v86ac9b;
assign v85e351 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8633e4;
assign v86b7b7 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v86b132;
assign v8caa40 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85dee1;
assign v8ca246 = jx0_p & v86d0cd | !jx0_p & v85d3a1;
assign v8c95d7 = jx0_p & v85dfad | !jx0_p & v869b57;
assign v865427 = jx2_p & v8cac4e | !jx2_p & v8ca742;
assign v864bf9 = StoB_REQ1_p & v8caab9 | !StoB_REQ1_p & v8cac00;
assign v8ca937 = jx1_p & v8cac6d | !jx1_p & v89b000;
assign v85b56a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8cac4a;
assign v844f91 = 1;
assign v86d3d9 = BtoS_ACK0_p & v8cab9f | !BtoS_ACK0_p & v86c833;
assign v844fbb = DEQ_p & v844f91 | !DEQ_p & !v844f91;
assign v86889b = BtoS_ACK0_p & v8caa61 | !BtoS_ACK0_p & v861d51;
assign v8cab49 = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & !v867780;
assign v8cab79 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855530;
assign v86b862 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86a7af;
assign v8692e8 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8858bf;
assign v86d1b3 = StoB_REQ0_p & v8caa48 | !StoB_REQ0_p & v8cabc0;
assign v8cad4e = DEQ_p & v868378 | !DEQ_p & v844fa7;
assign v85e715 = StoB_REQ2_p & v8617fa | !StoB_REQ2_p & !v86d276;
assign v8caa8a = jx2_p & v865321 | !jx2_p & !v8688ca;
assign v866d97 = DEQ_p & v8cab57 | !DEQ_p & v86882a;
assign v8699ec = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v865dfa;
assign v8cac9f = EMPTY_p & v86c701 | !EMPTY_p & v8663ef;
assign v862180 = EMPTY_p & v8cacb5 | !EMPTY_p & v867b2b;
assign v869baf = BtoS_ACK0_p & v8cab71 | !BtoS_ACK0_p & !v8671ac;
assign v860a37 = stateG12_p & v8452cf | !stateG12_p & !v844f91;
assign v862012 = jx1_p & v844f91 | !jx1_p & v86665f;
assign v85cebf = EMPTY_p & v8caada | !EMPTY_p & !v844f91;
assign v8caa0a = ENQ_p & v8690d8 | !ENQ_p & v8651a5;
assign v867010 = jx2_p & v85e138 | !jx2_p & !v8cac6d;
assign v8683f7 = stateG7_1_p & v868830 | !stateG7_1_p & v86c57f;
assign v86d775 = StoB_REQ0_p & v861bb6 | !StoB_REQ0_p & v8a74b4;
assign v861379 = StoB_REQ1_p & v8caaf5 | !StoB_REQ1_p & v8cac02;
assign BtoS_ACK3_n = !v87133e;
assign v8ca98e = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8cac4a;
assign v86a764 = ENQ_p & v8cac43 | !ENQ_p & v869922;
assign v8ca695 = jx0_p & v86d101 | !jx0_p & v869b57;
assign v8650ba = jx0_p & v85f4ff | !jx0_p & v85d3a1;
assign v86d803 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c9b86;
assign v8ca9c9 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8cacd1;
assign v866b1d = BtoS_ACK1_p & v861ecc | !BtoS_ACK1_p & v85f4c4;
assign v86b348 = DEQ_p & v860a57 | !DEQ_p & v867b84;
assign v8cac84 = EMPTY_p & v861905 | !EMPTY_p & v866037;
assign v86a618 = RtoB_ACK1_p & v8697c8 | !RtoB_ACK1_p & v8679eb;
assign v8c97e3 = EMPTY_p & v86607a | !EMPTY_p & v8c9f2a;
assign v867508 = jx0_p & v8caace | !jx0_p & !v844f91;
assign v865fe6 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v85e8ee;
assign v89c777 = jx1_p & v844f99 | !jx1_p & !v8ca9c3;
assign v8666db = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v859567;
assign v86267d = BtoS_ACK0_p & v844f9c | !BtoS_ACK0_p & v8caa02;
assign v8664d8 = RtoB_ACK1_p & v864071 | !RtoB_ACK1_p & !v844f91;
assign v85d9cf = EMPTY_p & v869ddd | !EMPTY_p & v8a74c0;
assign v860ea5 = jx1_p & v86889a | !jx1_p & v860af3;
assign v861290 = DEQ_p & v860a1c | !DEQ_p & v8cacc7;
assign v8cacba = stateG12_p & v867d26 | !stateG12_p & v89afeb;
assign v86a6c6 = jx2_p & v8cab89 | !jx2_p & v8cab4b;
assign v8cabf5 = StoB_REQ0_p & v8cab1a | !StoB_REQ0_p & v8cab90;
assign v8c9bd7 = RtoB_ACK1_p & v8caa4a | !RtoB_ACK1_p & v8cad96;
assign v85dade = RtoB_ACK1_p & v8c9e60 | !RtoB_ACK1_p & !v844f91;
assign v85e4b1 = StoB_REQ0_p & v865507 | !StoB_REQ0_p & v8cacc4;
assign v8ca9d5 = jx2_p & v8caccc | !jx2_p & v844f91;
assign v85e5c6 = BtoS_ACK2_p & v8caa43 | !BtoS_ACK2_p & v8caa14;
assign v86b96c = jx1_p & v8caa0f | !jx1_p & v865036;
assign v844f9e = StoB_REQ4_n & v844f91 | !StoB_REQ4_n & !v844f91;
assign v8cabe9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v861266;
assign v867abe = RtoB_ACK0_p & v864207 | !RtoB_ACK0_p & v868dd2;
assign v8cacaa = StoB_REQ1_p & v8cac02 | !StoB_REQ1_p & v867769;
assign v86ae3e = FULL_p & v86a953 | !FULL_p & v8cab59;
assign v85d843 = ENQ_p & v867c81 | !ENQ_p & v8940d7;
assign v85e4b6 = ENQ_p & v8cac80 | !ENQ_p & v866ee5;
assign v85cdd6 = BtoR_REQ1_p & v867507 | !BtoR_REQ1_p & v8794af;
assign v86b298 = StoB_REQ2_p & v8617fa | !StoB_REQ2_p & !v8c9c7c;
assign v879497 = ENQ_p & v865e4b | !ENQ_p & v8ca522;
assign v866d1f = EMPTY_p & v8cac35 | !EMPTY_p & !v844f91;
assign v868403 = jx1_p & v86685a | !jx1_p & v86b9ab;
assign v861fda = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v85d53b;
assign v8660c6 = ENQ_p & v8cac80 | !ENQ_p & v8712ee;
assign v8cad5f = jx2_p & v8688ca | !jx2_p & v844f91;
assign v8caacc = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8cadb0;
assign v8cac8e = jx1_p & v860e50 | !jx1_p & !v8cabed;
assign v8cacde = FULL_p & v844f91 | !FULL_p & !v8ca9c1;
assign v85e6c0 = DEQ_p & v8647a2 | !DEQ_p & v861dcc;
assign v86d402 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8678d8;
assign v85de38 = BtoS_ACK0_p & v85e2e7 | !BtoS_ACK0_p & v8caaab;
assign v86b74a = StoB_REQ3_p & v86b132 | !StoB_REQ3_p & !v844f91;
assign v8c96e3 = jx2_p & v8caaae | !jx2_p & v865edc;
assign v867bc5 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v844f91;
assign v8cac4b = jx1_p & v8ca61e | !jx1_p & !v8cab4c;
assign v8caa4d = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v861774 = EMPTY_p & v8c963c | !EMPTY_p & v865bf0;
assign v86113b = BtoS_ACK0_p & v868129 | !BtoS_ACK0_p & !v8caa15;
assign v8c9c26 = jx1_p & v8cac66 | !jx1_p & !v8caac2;
assign v8caa20 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8691f2;
assign v861889 = ENQ_p & v89af47 | !ENQ_p & v86d0ec;
assign v8664b1 = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v844f91;
assign v85e569 = StoB_REQ0_p & v8caa58 | !StoB_REQ0_p & v844f91;
assign v86b132 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9d;
assign v85e4fc = StoB_REQ0_p & v8caa66 | !StoB_REQ0_p & v85e88d;
assign v8667e9 = jx0_p & v85d919 | !jx0_p & !v8679f8;
assign v8cadb0 = BtoS_ACK2_p & v8caa43 | !BtoS_ACK2_p & v8cac12;
assign v85f516 = StoB_REQ2_p & v8c9be8 | !StoB_REQ2_p & v85daff;
assign v8cab90 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8588a0;
assign v8ca3c3 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v86b485;
assign v865dbb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8678e6;
assign v8c9d1a = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v8ca2af;
assign v86dae3 = jx0_p & v8ca3d4 | !jx0_p & !v862fc7;
assign v868378 = jx0_p & v8caac4 | !jx0_p & v844fa7;
assign v8c9a7e = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v869631;
assign v866e01 = stateG12_p & v866b27 | !stateG12_p & !v86652d;
assign v86b6e3 = DEQ_p & v844f91 | !DEQ_p & v844fa5;
assign v8b69b8 = DEQ_p & v8ca9f0 | !DEQ_p & v868f7d;
assign v8c9626 = jx1_p & v8cac6d | !jx1_p & v85e228;
assign v8cac28 = ENQ_p & v8cac79 | !ENQ_p & !v85e5ff;
assign v8caca3 = EMPTY_p & v844f91 | !EMPTY_p & v8caa7e;
assign v8cac35 = jx0_p & v85e110 | !jx0_p & v869e56;
assign v85de90 = jx2_p & v866fa1 | !jx2_p & v8cab3e;
assign v852940 = DEQ_p & v867a99 | !DEQ_p & v8ca04b;
assign v85cd74 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86ac7c;
assign v864b34 = StoB_REQ0_p & v8caa66 | !StoB_REQ0_p & v85d772;
assign v8c9712 = jx1_p & v869f33 | !jx1_p & v85e3f3;
assign v8cac1a = jx1_p & v8b69a7 | !jx1_p & v86a5b6;
assign v866cf1 = jx1_p & v867edf | !jx1_p & !v864ad9;
assign v8a74fd = EMPTY_p & v856fa3 | !EMPTY_p & v844f91;
assign v8609a9 = EMPTY_p & v8cabeb | !EMPTY_p & v866aae;
assign v85e337 = BtoS_ACK1_p & v861ecc | !BtoS_ACK1_p & v86add5;
assign v85d880 = StoB_REQ2_p & v85d750 | !StoB_REQ2_p & v8cab1c;
assign v894103 = ENQ_p & v8cabd8 | !ENQ_p & v8cabc7;
assign v86265a = StoB_REQ2_p & v8617fa | !StoB_REQ2_p & !v8ca354;
assign v86b5da = jx1_p & v85f4cf | !jx1_p & v85dbdc;
assign v861db7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86294e;
assign v86863b = EMPTY_p & v844f91 | !EMPTY_p & !v8c9a6e;
assign v8c963c = jx0_p & v868dd9 | !jx0_p & !v8632cd;
assign v86c701 = jx0_p & v863449 | !jx0_p & v88656a;
assign v867a75 = jx0_p & v8caa9a | !jx0_p & v867d26;
assign v8cab77 = DEQ_p & v8caa52 | !DEQ_p & v8cac96;
assign v8633e4 = StoB_REQ1_p & v86b05b | !StoB_REQ1_p & v844f91;
assign v8caa5f = FULL_p & v844f91 | !FULL_p & v8cab44;
assign v869b48 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v86b1d8;
assign v867ba8 = BtoS_ACK0_p & v8caac6 | !BtoS_ACK0_p & v86b862;
assign v86d6a1 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v86d329;
assign v86d147 = ENQ_p & v8cac80 | !ENQ_p & v8caa7c;
assign BtoS_ACK0_n = v88d17c;
assign v8cac10 = jx0_p & v8caa36 | !jx0_p & v869b57;
assign v89afeb = jx2_p & v8cac6d | !jx2_p & v867d26;
assign v8caa89 = EMPTY_p & v85309b | !EMPTY_p & v85da2b;
assign v8caaca = ENQ_p & v844f91 | !ENQ_p & v861dac;
assign v8cace6 = jx0_p & v85ac07 | !jx0_p & !v861171;
assign v89af47 = DEQ_p & v844f91 | !DEQ_p & !v8678d9;
assign v8caa15 = StoB_REQ0_p & v8450db | !StoB_REQ0_p & v8ca8d6;
assign v8cabcd = jx1_p & v844f99 | !jx1_p & !v8ca9d5;
assign v867a22 = StoB_REQ1_p & v89afb5 | !StoB_REQ1_p & v86d74c;
assign v8cab63 = DEQ_p & v8caa57 | !DEQ_p & v861fb9;
assign v8c9dae = DEQ_p & v86a60b | !DEQ_p & v8cac9f;
assign v8cac76 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v844f91;
assign v85cef2 = RtoB_ACK0_p & v8cac28 | !RtoB_ACK0_p & v86150f;
assign v8cab70 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v85cdad;
assign v86a607 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v866b54;
assign v860e09 = jx2_p & v866369 | !jx2_p & v844f91;
assign v86653c = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v8c9811;
assign v89af9c = FULL_p & v844f91 | !FULL_p & !v86d5ab;
assign v856a93 = StoB_REQ2_p & v89afb5 | !StoB_REQ2_p & v844f91;
assign v8cacb0 = jx0_p & v852479 | !jx0_p & v844f91;
assign v86adad = EMPTY_p & v8ca246 | !EMPTY_p & v8caad8;
assign v86702e = ENQ_p & v8cac43 | !ENQ_p & v8c9ef9;
assign v862bd2 = ENQ_p & v8cac80 | !ENQ_p & v85d881;
assign v8c9a57 = StoB_REQ0_p & v8ca7ed | !StoB_REQ0_p & v86d402;
assign v865321 = BtoS_ACK0_p & v8caa5a | !BtoS_ACK0_p & v86560f;
assign v8caa3f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85a021;
assign v8ca126 = ENQ_p & v8cac80 | !ENQ_p & v8ca5e2;
assign v85c2e5 = StoB_REQ2_p & v8ca9fa | !StoB_REQ2_p & v867bc5;
assign v85a733 = jx2_p & v86d557 | !jx2_p & v85cf1e;
assign v8caac0 = DEQ_p & v865bf0 | !DEQ_p & v86ade6;
assign v8caaa9 = jx2_p & v844f91 | !jx2_p & v8cab4b;
assign v8858c9 = BtoR_REQ0_p & v861436 | !BtoR_REQ0_p & v861d21;
assign v8696e7 = BtoS_ACK0_p & v8cac4a | !BtoS_ACK0_p & v85df95;
assign v8cac3a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8caa44;
assign v868e01 = FULL_p & v85d221 | !FULL_p & v85e743;
assign v8612b9 = BtoS_ACK0_p & v86ac9b | !BtoS_ACK0_p & v8ca9de;
assign v8662c3 = jx1_p & v8cac6d | !jx1_p & v8cacd8;
assign v8cac46 = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v8ca56d;
assign v8cac66 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8ca472;
assign v89afb5 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v86631f;
assign v85d954 = jx1_p & v8caba9 | !jx1_p & v85d39c;
assign v85ce75 = ENQ_p & v8cab63 | !ENQ_p & v867763;
assign v8caa06 = BtoS_ACK3_p & v8cacd6 | !BtoS_ACK3_p & v8ca9fa;
assign v8cac6a = EMPTY_p & v867d26 | !EMPTY_p & v8c9890;
assign v8caa53 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8caa6e;
assign v8683f9 = jx1_p & v8cab94 | !jx1_p & !v8cab37;
assign v8cac0f = ENQ_p & v8cad4e | !ENQ_p & !v866205;
assign v8cabed = jx2_p & v8cac6d | !jx2_p & v86d231;
assign v8ca9c7 = StoB_REQ1_p & v8caaf5 | !StoB_REQ1_p & v862264;
assign v8cab89 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ca009;
assign v8c9ed8 = StoB_REQ1_p & v8654fc | !StoB_REQ1_p & v869ca4;
assign v8cac5d = ENQ_p & v8cac43 | !ENQ_p & v867551;
assign v865295 = jx2_p & v8ca153 | !jx2_p & !v844f91;
assign v86d322 = stateG7_1_p & v86b3cd | !stateG7_1_p & v844f91;
assign v860aed = DEQ_p & v8cac70 | !DEQ_p & v865787;
assign v86b05c = StoB_REQ2_p & v865dfa | !StoB_REQ2_p & v8c9c7c;
assign v8679f8 = jx1_p & v8caa0f | !jx1_p & v8672bb;
assign v8cabfe = jx1_p & v844f91 | !jx1_p & !v8cabe2;
assign v86bae1 = jx2_p & v85de38 | !jx2_p & !v8caae9;
assign v8610ac = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v844f91;
assign v8caaef = jx2_p & v8cab4b | !jx2_p & !v844fa7;
assign v8452cf = jx2_p & v844f91 | !jx2_p & !v844f91;
assign v85d4df = StoB_REQ3_p & v86b132 | !StoB_REQ3_p & v844f91;
assign v8ca154 = jx1_p & v844f91 | !jx1_p & !v865295;
assign v8c9a6e = jx0_p & v8caace | !jx0_p & !v862fc7;
assign v8caca2 = StoB_REQ1_p & v868cbe | !StoB_REQ1_p & v844f91;
assign v8caafd = StoB_REQ1_p & v8caab9 | !StoB_REQ1_p & v86202e;
assign v85d985 = StoB_REQ0_p & v8ca7ed | !StoB_REQ0_p & v8cab81;
assign v8caac2 = jx2_p & v844f91 | !jx2_p & v868626;
assign v86c524 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8ca9fa;
assign v8794af = stateG7_1_p & v85c630 | !stateG7_1_p & v8cabd2;
assign v85f3fa = DEQ_p & v8cab57 | !DEQ_p & v86b7bb;
assign v8caa9b = stateG7_1_p & v8c9cbc | !stateG7_1_p & v86c801;
assign v8c9db1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86822b;
assign v8cab19 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9b;
assign v85dac9 = BtoS_ACK0_p & v8cab9f | !BtoS_ACK0_p & v8cab1d;
assign v85e743 = jx0_p & v8caabc | !jx0_p & v8ca022;
assign v867a20 = jx0_p & v85b1cb | !jx0_p & v85db64;
assign v85e733 = jx1_p & v86b125 | !jx1_p & !v862256;
assign v868905 = jx2_p & v85d7eb | !jx2_p & v844f91;
assign v8b3167 = jx2_p & v8621d5 | !jx2_p & v865edc;
assign v8caa7f = stateG7_1_p & v8caad4 | !stateG7_1_p & v86a764;
assign v8cac2d = StoB_REQ0_p & v8677dc | !StoB_REQ0_p & v844f91;
assign v859cb4 = ENQ_p & v85daa3 | !ENQ_p & !v86d390;
assign v85e78a = jx2_p & v844f91 | !jx2_p & v86a607;
assign v86d805 = BtoS_ACK0_p & v8cac4a | !BtoS_ACK0_p & v865811;
assign v8ca172 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v863955;
assign v86d81c = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & v8cab6c;
assign v867417 = EMPTY_p & v869d71 | !EMPTY_p & v8cabde;
assign v86af9f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cac4a;
assign v8caa61 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v85d451 = jx1_p & v8ca9e4 | !jx1_p & !v8c977d;
assign v85e1cc = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v8cab3d;
assign v86af4a = StoB_REQ0_p & v86816d | !StoB_REQ0_p & v8cab05;
assign v860b60 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8c97c4;
assign v86ac7c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8caa20;
assign v8ca849 = StoB_REQ1_p & v867166 | !StoB_REQ1_p & v844f91;
assign v89c779 = BtoR_REQ0_p & v8a6000 | !BtoR_REQ0_p & v86770a;
assign v8692f8 = FULL_p & v866d0b | !FULL_p & !v8cacb0;
assign v8c9ef9 = DEQ_p & v865bf0 | !DEQ_p & v8cacb6;
assign v86b3cd = RtoB_ACK1_p & v861889 | !RtoB_ACK1_p & v844f91;
assign v8cac70 = jx0_p & v86a745 | !jx0_p & v85d954;
assign v866d78 = jx0_p & v8c9b41 | !jx0_p & !v85e183;
assign v8cab5a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v864b34;
assign v866606 = RtoB_ACK1_p & v86ba45 | !RtoB_ACK1_p & v861c02;
assign v8c9f14 = EMPTY_p & v8cab57 | !EMPTY_p & v866aae;
assign v85d86a = StoB_REQ2_p & v8664cd | !StoB_REQ2_p & v86a6a1;
assign v8c9dd4 = jx1_p & v85dd97 | !jx1_p & v844f91;
assign v866d8b = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v8caab0;
assign v8cab9b = jx1_p & v86b50c | !jx1_p & v8caa18;
assign v86d7ce = EMPTY_p & v8ca9db | !EMPTY_p & !v861166;
assign v868cbc = stateG7_1_p & v844f91 | !stateG7_1_p & !v860ab6;
assign v8cacdc = RtoB_ACK1_p & v85e3ea | !RtoB_ACK1_p & v8caaca;
assign v8cab57 = jx0_p & v8cac6d | !jx0_p & v86aebe;
assign v8c9890 = jx0_p & v8cac39 | !jx0_p & v867d26;
assign v8c9b2e = stateG7_1_p & v85d8cc | !stateG7_1_p & v86b725;
assign v866bf7 = EMPTY_p & v844f91 | !EMPTY_p & !v869b15;
assign v861ecc = StoB_REQ3_n & v844f91 | !StoB_REQ3_n & v844f9e;
assign v8693ab = jx0_p & v862200 | !jx0_p & v86b50c;
assign v8caa11 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v86ac5d;
assign v86d390 = DEQ_p & v8cabec | !DEQ_p & v867f36;
assign v8794d1 = StoB_REQ2_p & v866964 | !StoB_REQ2_p & !v844f91;
assign v86921b = jx1_p & v8caac1 | !jx1_p & !v8c9e27;
assign v8cac33 = BtoS_ACK0_p & v8c9942 | !BtoS_ACK0_p & v8cab5d;
assign v8cacd2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cad66;
assign v8caae4 = jx2_p & v86d231 | !jx2_p & !v85d906;
assign v85e297 = StoB_REQ0_p & v8caa6e | !StoB_REQ0_p & v8cac81;
assign v867e4a = EMPTY_p & v844f91 | !EMPTY_p & v86538c;
assign v8ca04b = EMPTY_p & v86c461 | !EMPTY_p & v867a99;
assign v85d173 = jx1_p & v8caad7 | !jx1_p & !v8ca349;
assign v86ac5d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v867bc5;
assign v86c461 = jx0_p & v85d919 | !jx0_p & !v86b96c;
assign v8a74c0 = jx0_p & v866997 | !jx0_p & v8612ab;
assign v8caba7 = jx0_p & v8caa1b | !jx0_p & !v85d80e;
assign v86d378 = BtoS_ACK0_p & v8c7b0b | !BtoS_ACK0_p & v86912f;
assign v85ce03 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v85da42;
assign v86a8b8 = jx2_p & v86b711 | !jx2_p & v86d231;
assign v8cac05 = stateG12_p & v8cad5f | !stateG12_p & v8cacca;
assign v861be5 = DEQ_p & v8ca9cd | !DEQ_p & v864a62;
assign v8b69e1 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & v86afde;
assign v8690d8 = DEQ_p & v8693ab | !DEQ_p & v86b50c;
assign v86116b = jx1_p & v844f99 | !jx1_p & !v8ca9d3;
assign v8caad3 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8caa17;
assign v867a99 = jx0_p & v868b0c | !jx0_p & !v8ca9ff;
assign v8cac96 = EMPTY_p & v8ca9db | !EMPTY_p & v8cabde;
assign v867c16 = DEQ_p & v844f91 | !DEQ_p & v8cac4f;
assign v8641cf = EMPTY_p & v85e8c7 | !EMPTY_p & !v844f91;
assign v86c833 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cab49;
assign v8cac6d = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v867220;
assign v85f380 = ENQ_p & v868e55 | !ENQ_p & !v85d22b;
assign v867a8a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v868f18;
assign v8ca9af = DEQ_p & v844f91 | !DEQ_p & v8cab6b;
assign v865cd4 = jx2_p & v8c9e00 | !jx2_p & v844f91;
assign v8c9aea = DEQ_p & v8cab07 | !DEQ_p & v8c97e3;
assign v8cabc6 = StoB_REQ0_p & v86816d | !StoB_REQ0_p & v8caaec;
assign v8c7b4e = jx1_p & v844f91 | !jx1_p & v8ca313;
assign v8c9c9f = EMPTY_p & v8649c5 | !EMPTY_p & v8ca3cb;
assign v8ca1e1 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8caa62;
assign v861df7 = RtoB_ACK1_p & v8660c6 | !RtoB_ACK1_p & v86d147;
assign v8caa44 = StoB_REQ2_p & v8cab15 | !StoB_REQ2_p & v85e8ff;
assign v8679eb = ENQ_p & v8c9dae | !ENQ_p & !v8677e5;
assign v8621d5 = BtoS_ACK0_p & v8ca98e | !BtoS_ACK0_p & v8cabc6;
assign v8ca61e = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v86d753;
assign v8c9cad = jx1_p & v8caa8f | !jx1_p & v844f91;
assign v8668d6 = jx1_p & v86889b | !jx1_p & v8cab3e;
assign v865e2b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cac20;
assign v8ca9d0 = DEQ_p & v86a60b | !DEQ_p & v8ca5b3;
assign v85e224 = ENQ_p & v865e4b | !ENQ_p & v844f91;
assign v86b7d3 = BtoR_REQ1_p & v86d7e6 | !BtoR_REQ1_p & v8cac3e;
assign v8caaf8 = StoB_REQ2_p & v86b132 | !StoB_REQ2_p & !v8c9c7c;
assign v8ca374 = ENQ_p & v8cac79 | !ENQ_p & !v8cac03;
assign v866810 = EMPTY_p & v869d71 | !EMPTY_p & !v861166;
assign v861525 = FULL_p & v867508 | !FULL_p & v86d2f5;
assign v8cabbb = jx0_p & v85e7b6 | !jx0_p & !v8675a9;
assign v8cab39 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v862264;
assign v85e69b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844fab;
assign v86b7bb = EMPTY_p & v8cabeb | !EMPTY_p & v869992;
assign v86d0cd = jx1_p & v8c9e5e | !jx1_p & !v8613f4;
assign v85f4ff = jx1_p & v8c9e5e | !jx1_p & v86859e;
assign v86b786 = EMPTY_p & v8667e9 | !EMPTY_p & v8caa60;
assign v8667fb = DEQ_p & v844f91 | !DEQ_p & v866d1f;
assign v894106 = BtoR_REQ0_p & v85cef2 | !BtoR_REQ0_p & v867abe;
assign v86a660 = stateG12_p & v844fa7 | !stateG12_p & !v8c9ce3;
assign v8ca686 = BtoS_ACK2_p & v8caa43 | !BtoS_ACK2_p & v85d90c;
assign v8c9f2a = FULL_p & v8cac22 | !FULL_p & v8a5ffe;
assign v861882 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8664cd;
assign v856fa3 = jx0_p & v85d173 | !jx0_p & v8940fd;
assign v85769e = jx2_p & v85d6e1 | !jx2_p & !v844f91;
assign v85d1d4 = jx1_p & v862e4a | !jx1_p & !v8c9e27;
assign v866a61 = StoB_REQ0_p & v865507 | !StoB_REQ0_p & v8cac08;
assign v8c9b09 = FULL_p & v8cac54 | !FULL_p & !v8a5ffe;
assign v8caa29 = EMPTY_p & v8679ab | !EMPTY_p & v8ca695;
assign v867f36 = EMPTY_p & v8cab34 | !EMPTY_p & !v879471;
assign v8cac41 = jx1_p & v8cab94 | !jx1_p & !v8cab08;
assign v8b2a0d = RtoB_ACK0_p & v86608e | !RtoB_ACK0_p & v85d56c;
assign v85dbc1 = jx1_p & v844f91 | !jx1_p & v8cacca;
assign v8ca17e = ENQ_p & v86817a | !ENQ_p & v865936;
assign v8caa1b = jx1_p & v869497 | !jx1_p & !v86652d;
assign v85d23a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8c7b0b;
assign v8c9d37 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v8cab19;
assign v85e11a = EMPTY_p & v86d2a8 | !EMPTY_p & v8cac9c;
assign v86b436 = BtoS_ACK0_p & v8cab3d | !BtoS_ACK0_p & v8caaa8;
assign v860ec7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8b69a2;
assign v86adcf = jx2_p & v86d231 | !jx2_p & v85d5c3;
assign v85d43c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v8caaaa = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v862881;
assign v8caa52 = jx0_p & v8c9b72 | !jx0_p & !v861494;
assign v85ce31 = EMPTY_p & v86c701 | !EMPTY_p & v8ca7e1;
assign v8caa33 = BtoS_ACK1_p & v86c73b | !BtoS_ACK1_p & v86ae59;
assign v85e0d5 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v869b48;
assign v85de3b = jx2_p & v8ca345 | !jx2_p & v8cab4b;
assign v88d12d = FULL_p & v8cac54 | !FULL_p & !v8692bc;
assign v8cab59 = jx0_p & v8ca742 | !jx0_p & v86aec5;
assign v8ca693 = BtoS_ACK0_p & v8cab19 | !BtoS_ACK0_p & v867220;
assign v8ca0f9 = DEQ_p & v86b799 | !DEQ_p & v8cabc1;
assign v869284 = DEQ_p & v85e2d7 | !DEQ_p & v844fa7;
assign v8cacdb = ENQ_p & v868e55 | !ENQ_p & !v86b75f;
assign v8667bd = StoB_REQ2_p & v86b7b7 | !StoB_REQ2_p & !v857888;
assign v8cabfd = jx1_p & v8ca742 | !jx1_p & v860cd1;
assign v869065 = jx0_p & v8675fc | !jx0_p & !v87131b;
assign v865811 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cab36;
assign v866d9e = ENQ_p & v85daa3 | !ENQ_p & !v8c9cc5;
assign DEQ_n = !v8a6050;
assign v86d136 = DEQ_p & v861f9e | !DEQ_p & v85cebf;
assign v866bb9 = jx1_p & v844f91 | !jx1_p & v8cab8f;
assign v8cab0a = BtoS_ACK3_p & v85d4df | !BtoS_ACK3_p & v86b132;
assign v8b31d3 = jx0_p & v869f33 | !jx0_p & v8c9712;
assign v8ca9f3 = jx2_p & v844f91 | !jx2_p & v852627;
assign v86d7e6 = stateG7_1_p & v85dda7 | !stateG7_1_p & v8c9bfc;
assign v85c85e = jx2_p & v844f91 | !jx2_p & !v86d0bf;
assign v8656ee = jx0_p & v86b4f5 | !jx0_p & v85da6a;
assign v8667f6 = jx1_p & v844f91 | !jx1_p & !v8cac09;
assign v8c9b51 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v86d61d;
assign v86b485 = StoB_REQ1_p & v8712d5 | !StoB_REQ1_p & v867769;
assign v865707 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8cac71;
assign v8cab9c = ENQ_p & v868e55 | !ENQ_p & !v8cacc5;
assign v85d53b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v86b132;
assign v8ca9db = jx0_p & v8675fc | !jx0_p & !v8667cc;
assign v86d7f2 = DEQ_p & v86b799 | !DEQ_p & v8cac8c;
assign v8cac16 = jx1_p & v86889b | !jx1_p & v86a611;
assign v85db64 = jx1_p & v86b125 | !jx1_p & !v86a8b8;
assign v861d51 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8caa61;
assign v8a7515 = BtoR_REQ0_p & v866af0 | !BtoR_REQ0_p & v8caa2e;
assign v86830a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v867be8;
assign v8648c8 = jx1_p & v844f91 | !jx1_p & !v865bb1;
assign v8c95e9 = ENQ_p & v85cde5 | !ENQ_p & v8caa6b;
assign v86490e = jx1_p & v861d1f | !jx1_p & v85da17;
assign v85e185 = EMPTY_p & v869065 | !EMPTY_p & !v89af9c;
assign v8ca701 = jx1_p & v867edf | !jx1_p & v86665f;
assign v8caad2 = jx1_p & v844f91 | !jx1_p & v86a6c6;
assign v86b02f = jx2_p & v8c9bd1 | !jx2_p & v86d231;
assign v8594af = FULL_p & v844f91 | !FULL_p & v8cac0a;
assign v86d602 = ENQ_p & v8940e1 | !ENQ_p & v85d8fe;
assign v8cabcc = StoB_REQ2_p & v8caba0 | !StoB_REQ2_p & !v844f91;
assign v869b6e = jx1_p & v865f35 | !jx1_p & v852625;
assign v864050 = RtoB_ACK0_p & v869ec7 | !RtoB_ACK0_p & v8599dd;
assign v85e65a = jx1_p & v8674b4 | !jx1_p & v8ca9fb;
assign v8607fe = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9c;
assign v8cac98 = StoB_REQ2_p & v8cab0a | !StoB_REQ2_p & !v844f91;
assign v8c9a79 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f9c;
assign v86d813 = EMPTY_p & v844f91 | !EMPTY_p & v8cab44;
assign v8651a3 = stateG12_p & v85da6a | !stateG12_p & v86974a;
assign v86d130 = StoB_REQ2_p & v86b7b7 | !StoB_REQ2_p & !v865cb0;
assign v867b84 = EMPTY_p & v85309b | !EMPTY_p & v86538c;
assign v8caa7d = BtoS_ACK0_p & v8691f2 | !BtoS_ACK0_p & v85d232;
assign v861b6c = jx2_p & v875b43 | !jx2_p & v8cab4b;
assign v8c99d1 = BtoS_ACK0_p & v8caa5a | !BtoS_ACK0_p & v8cabfc;
assign v85f4e3 = EMPTY_p & v88d120 | !EMPTY_p & !v867957;
assign v86817a = DEQ_p & v869112 | !DEQ_p & v86889a;
assign v85da6a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v865507;
assign v8609fc = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8ca7ed;
assign v86d0ec = DEQ_p & v844f91 | !DEQ_p & v868ba7;
assign v865012 = StoB_REQ0_p & v86d5fc | !StoB_REQ0_p & v856f8c;
assign v844fa9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v869a67 = StoB_REQ2_p & v8617fa | !StoB_REQ2_p & !v844f91;
assign v865c5c = jx1_p & v8ca79e | !jx1_p & v869e35;
assign v86752a = jx1_p & v85f4cf | !jx1_p & v8cabef;
assign v8ca56d = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v8cab71;
assign v8666cf = FULL_p & v867508 | !FULL_p & v86d5ab;
assign v8598f7 = EMPTY_p & v8647a2 | !EMPTY_p & v8caa5f;
assign v868c7d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v861b86;
assign v8ca9e3 = jx2_p & v844f91 | !jx2_p & v85cf1e;
assign v86908c = jx2_p & v86d378 | !jx2_p & !v85c5d4;
assign v8cab8e = ENQ_p & v8caafc | !ENQ_p & v844f91;
assign v867780 = StoB_REQ1_p & v86265a | !StoB_REQ1_p & v8cab84;
assign v86b30e = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v866d60;
assign v8cab6c = StoB_REQ2_p & v865dfa | !StoB_REQ2_p & v8ca354;
assign v8612e7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c9df0;
assign v86d2a8 = jx0_p & v85ac07 | !jx0_p & !v866860;
assign v85d448 = jx1_p & v844f91 | !jx1_p & v867565;
assign v8c9df0 = BtoS_ACK1_p & v8cac4a | !BtoS_ACK1_p & !v8cac98;
assign v852479 = jx1_p & v844f91 | !jx1_p & !v860a37;
assign v86882a = EMPTY_p & v85dfa3 | !EMPTY_p & v844f91;
assign v8cac54 = jx0_p & v85dbc1 | !jx0_p & v869b57;
assign v8cac79 = DEQ_p & v86a60b | !DEQ_p & v8660ec;
assign v87133e = BtoR_REQ0_p & v88d0f1 | !BtoR_REQ0_p & v8c9a18;
assign v8caa0f = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v867a8a;
assign v85f4cf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e2ea;
assign v8cac81 = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v8c9ace;
assign v8712ee = DEQ_p & v86a66f | !DEQ_p & v85e11a;
assign v861bb6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85cdfc;
assign v860cd1 = stateG12_p & v8ca742 | !stateG12_p & v85e164;
assign v866fa1 = BtoS_ACK0_p & v8cac4a | !BtoS_ACK0_p & v86af9f;
assign v8c9be8 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v844f91;
assign v86621a = DEQ_p & v865bf0 | !DEQ_p & v861774;
assign v8caa1d = jx1_p & v844f99 | !jx1_p & !v864ac7;
assign v8caae9 = BtoS_ACK0_p & v868129 | !BtoS_ACK0_p & !v8b69c5;
assign v86961e = ENQ_p & v86817a | !ENQ_p & v8ca737;
assign v86ac23 = ENQ_p & v861c01 | !ENQ_p & v860a1c;
assign v8b2a28 = EMPTY_p & v86d2a8 | !EMPTY_p & v8594af;
assign v8c9b41 = jx1_p & v8ca86e | !jx1_p & !v869653;
assign v894033 = RtoB_ACK0_p & v8c9d6e | !RtoB_ACK0_p & v8caa7f;
assign v86d5c8 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8ca21b;
assign v86b4f5 = jx1_p & v85da6a | !jx1_p & v8651a3;
assign v85e84a = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v8450db;
assign v8caa2f = jx1_p & v8ca61e | !jx1_p & !v85c85e;
assign v8ca3cb = jx0_p & v8cab74 | !jx0_p & v869b57;
assign v89b010 = BtoR_REQ0_p & v844f9f | !BtoR_REQ0_p & v8c9a1b;
assign v8cac09 = jx2_p & v86b30e | !jx2_p & !v844f91;
assign v8c9e09 = jx1_p & v86b70b | !jx1_p & !v85e310;
assign v85dee1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85e69b;
assign jx2_n = !v89c779;
assign v8ca21b = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v85d86a;
assign v89af2b = StoB_REQ2_p & v865dfa | !StoB_REQ2_p & v844f91;
assign v85e8cb = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v844f91;
assign v85e947 = StoB_REQ0_p & v8caa21 | !StoB_REQ0_p & v844f91;
assign v86d7d4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f99;
assign v867a34 = stateG7_1_p & v8664d8 | !stateG7_1_p & !v844f91;
assign v86494d = ENQ_p & v8ca9d0 | !ENQ_p & !v8caab8;
assign v86a7af = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caac6;
assign v867769 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8c9c7c;
assign v866f76 = StoB_REQ0_p & v865507 | !StoB_REQ0_p & v8caad1;
assign v869526 = EMPTY_p & v844f91 | !EMPTY_p & v864dbb;
assign v85d485 = FULL_p & v844f91 | !FULL_p & v864dbb;
assign v8c95c7 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v86b7fd;
assign v8c8cdb = BtoS_ACK0_p & v858cb9 | !BtoS_ACK0_p & v8c9d2e;
assign v8b69a2 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8c9811;
assign v86afde = RtoB_ACK0_p & v8cacb4 | !RtoB_ACK0_p & v86ba19;
assign v866c71 = DEQ_p & v8ca9f0 | !DEQ_p & v85f4e3;
assign v86911f = BtoS_ACK0_p & v8cab16 | !BtoS_ACK0_p & v865e2b;
assign v867551 = DEQ_p & v867a99 | !DEQ_p & v8653c0;
assign v86d25f = stateG7_1_p & v86707f | !stateG7_1_p & v8caadc;
assign v867d26 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8caa66;
assign v86a799 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8caca1;
assign v865ff9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8698ed;
assign v8940e1 = DEQ_p & v86b3a2 | !DEQ_p & v85dece;
assign v867957 = jx0_p & v864a04 | !jx0_p & v865960;
assign v85309b = jx0_p & v85ac07 | !jx0_p & !v8640bb;
assign v8ca9eb = jx1_p & v865859 | !jx1_p & v844f91;
assign v8cacc7 = EMPTY_p & v86922c | !EMPTY_p & v860a1c;
assign v869060 = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v8cacce;
assign v8cab12 = DEQ_p & v8ca9cd | !DEQ_p & v866326;
assign v85a2c9 = BtoS_ACK1_p & v86add5 | !BtoS_ACK1_p & v858cb9;
assign v8c9d60 = FULL_p & v85d34f | !FULL_p & v8692bc;
assign v86b111 = jx2_p & v86b436 | !jx2_p & !v8caae9;
assign v865cb0 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v86b7b7;
assign v85cde5 = DEQ_p & v86b3a2 | !DEQ_p & v85ce31;
assign v8cab6e = jx2_p & v8ca0ab | !jx2_p & !v8cab4b;
assign v8cac49 = jx2_p & v8caae9 | !jx2_p & !v8cac0d;
assign v8c9c7c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v86b74a;
assign v86aec5 = jx1_p & v8ca742 | !jx1_p & v865427;
assign v8cad54 = jx1_p & v8a749d | !jx1_p & v8ca9cf;
assign v8c9aac = DEQ_p & v86a66f | !DEQ_p & v8caa00;
assign v864080 = stateG12_p & v85da6a | !stateG12_p & v86890b;
assign v865bb1 = stateG12_p & v869a08 | !stateG12_p & !v844f91;
assign v8ca196 = EMPTY_p & v861905 | !EMPTY_p & !v879471;
assign v865a01 = jx0_p & v8a749d | !jx0_p & v8cad54;
assign v8ca9ff = jx1_p & v85ce03 | !jx1_p & v8672bb;
assign v864ad9 = jx2_p & v85c5d4 | !jx2_p & v85e84a;
assign v8ca9fd = jx2_p & v844f91 | !jx2_p & v86889a;
assign v8cac39 = jx1_p & v867d26 | !jx1_p & v8ca41e;
assign v868fc7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v857ca8;
assign v8cacc4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ca6a1;
assign v8691a7 = DEQ_p & v8cac70 | !DEQ_p & v8c97df;
assign v85dbdc = jx2_p & v85506c | !jx2_p & v8cab4b;
assign v86b05b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v86b7fd;
assign v85e3f3 = jx2_p & v8cab5a | !jx2_p & v869f33;
assign v8660b6 = BtoS_ACK2_p & v8caa43 | !BtoS_ACK2_p & v844f91;
assign v8cab94 = BtoS_ACK0_p & v8cab71 | !BtoS_ACK0_p & v8cac46;
assign v8cab15 = BtoS_ACK2_p & v861ecc | !BtoS_ACK2_p & v844f91;
assign v8c9af8 = stateG12_p & v86909b | !stateG12_p & !v86652d;
assign v85c6f5 = DEQ_p & v8cab9d | !DEQ_p & v8caacd;
assign v8cac02 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8ca354;
assign v862031 = FULL_p & v8cac54 | !FULL_p & v85e4f2;
assign v860d7c = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v85d4e0;
assign v8c9f9a = ENQ_p & v871300 | !ENQ_p & v844f91;
assign v8675fc = jx1_p & v868ccd | !jx1_p & v8698fa;
assign v8c9bbf = jx2_p & v8cac6d | !jx2_p & v860b19;
assign v861166 = FULL_p & v844f91 | !FULL_p & !v86d2f5;
assign v85cdfc = StoB_REQ2_p & v8ca9d4 | !StoB_REQ2_p & v86593c;
assign v8679a8 = jx2_p & v8cab3e | !jx2_p & v8cacad;
assign v8691f2 = StoB_REQ1_p & v8cab19 | !StoB_REQ1_p & v844f91;
assign v869197 = StoB_REQ0_p & v868569 | !StoB_REQ0_p & v844f91;
assign v8caafb = RtoB_ACK1_p & v862305 | !RtoB_ACK1_p & v85e5ed;
assign v869ca4 = StoB_REQ2_p & v8cab0a | !StoB_REQ2_p & !v867bc5;
assign v85dfad = jx1_p & v8620d1 | !jx1_p & !v860a37;
assign v85e09a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ca303;
assign v8c9ec8 = EMPTY_p & v861bd6 | !EMPTY_p & v8cac9b;
assign v86a745 = jx1_p & v85f7ba | !jx1_p & v852625;
assign v8c9e00 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8c9f67;
assign v8cabf3 = jx1_p & v844f99 | !jx1_p & v8ca553;
assign v868402 = DEQ_p & v8c9ce7 | !DEQ_p & v865f9a;
assign v85d9e0 = jx0_p & v8cacaf | !jx0_p & v86752a;
assign v869992 = jx0_p & v8667ba | !jx0_p & v86aebe;
assign v85da2b = jx0_p & v8cac16 | !jx0_p & !v864144;
assign v8caba0 = BtoS_ACK2_p & v867bc5 | !BtoS_ACK2_p & !v844f91;
assign v85e183 = jx1_p & v8caaaa | !jx1_p & v8caad0;
assign v8cacd0 = jx0_p & v869b57 | !jx0_p & v844f91;
assign v865fe1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8cab71;
assign v8675a9 = jx1_p & v85e6b9 | !jx1_p & v86b111;
assign v8cacb9 = stateG12_p & v86674c | !stateG12_p & !v86665f;
assign v85e35c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8caae1;
assign v868c4d = jx1_p & v8caa53 | !jx1_p & !v8cac0b;
assign v86ba15 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caa75;
assign v869259 = jx1_p & v88cf5c | !jx1_p & !v8ca9f3;
assign v863955 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9b;
assign v866138 = jx1_p & v844f91 | !jx1_p & !v85769e;
assign v8ca1f2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e1cc;
assign v8ca753 = DEQ_p & v8c7b49 | !DEQ_p & v862180;
assign v8cab84 = StoB_REQ2_p & v8617fa | !StoB_REQ2_p & !v867bc5;
assign v844fab = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v8c9aca = FULL_p & v85310f | !FULL_p & v8cab0e;
assign v8685d8 = EMPTY_p & v8cac87 | !EMPTY_p & v8673d4;
assign v85e813 = jx1_p & v869060 | !jx1_p & v85e228;
assign v85e95a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8ca9be;
assign v86a84a = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8c9b51;
assign v865bf0 = jx0_p & v868b0c | !jx0_p & !v85a4d3;
assign v8caa91 = StoB_REQ0_p & v8caa66 | !StoB_REQ0_p & v8cac2a;
assign v8cab72 = StoB_REQ2_p & v8cab0a | !StoB_REQ2_p & !v85a021;
assign v861794 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v862883;
assign v86d101 = jx1_p & v8ca61e | !jx1_p & !v860a37;
assign v8632cd = jx1_p & v8caa51 | !jx1_p & v861903;
assign v865404 = DEQ_p & v8cabec | !DEQ_p & v866b78;
assign v8c9681 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e4b1;
assign v866d6c = DEQ_p & v8caa52 | !DEQ_p & v866810;
assign v8cab3a = stateG7_1_p & v844f91 | !stateG7_1_p & !v860f28;
assign v8ca79e = BtoS_ACK0_p & v85e30d | !BtoS_ACK0_p & v8caa70;
assign v8cac6b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cab03;
assign v8cab01 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & !v844f91;
assign v86707f = ENQ_p & v8cad4e | !ENQ_p & !v8a74a8;
assign v89b002 = jx1_p & v844fa7 | !jx1_p & v86a660;
assign v8caac4 = jx1_p & v844fa7 | !jx1_p & v8ca23b;
assign v8c9ce3 = jx2_p & v844f91 | !jx2_p & !v844fa7;
assign v86b9ab = jx2_p & v8caa3a | !jx2_p & v85d91a;
assign v85d6cf = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v868b10;
assign v8cab04 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v868363;
assign v85d4e0 = stateG7_1_p & v8c9c59 | !stateG7_1_p & v844f91;
assign v85c5d4 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v8cac7c;
assign v8cab52 = DEQ_p & v8647a2 | !DEQ_p & v8598f7;
assign v86918c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8caa41;
assign v85dfa3 = jx0_p & v85e813 | !jx0_p & v8cac5e;
assign v858cb9 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86add5;
assign v85310f = jx0_p & v844f91 | !jx0_p & !v8caaff;
assign v85e1fe = StoB_REQ2_p & v8ca9fa | !StoB_REQ2_p & v86c524;
assign v85e2ea = StoB_REQ0_p & v86d7d4 | !StoB_REQ0_p & v844f91;
assign v86a7da = RtoB_ACK0_p & v85f2ab | !RtoB_ACK0_p & v85e544;
assign v8cabff = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v852627;
assign v8a6050 = BtoR_REQ0_p & v8ca615 | !BtoR_REQ0_p & v89409f;
assign v86607a = jx0_p & v85b1cb | !jx0_p & v8caa56;
assign v8674f7 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86b05b;
assign v8a5ffe = jx0_p & v864a04 | !jx0_p & v89c777;
assign v8caade = jx2_p & v8cab97 | !jx2_p & v844f91;
assign v8673d4 = FULL_p & v865bf0 | !FULL_p & v866af3;
assign v85b1cb = jx1_p & v8ca089 | !jx1_p & !v86adcf;
assign v85cec5 = jx0_p & v8caaf0 | !jx0_p & v869b57;
assign v85a4d3 = jx1_p & v85ce03 | !jx1_p & v8caa31;
assign v8cabfc = StoB_REQ0_p & v8ca7ed | !StoB_REQ0_p & v86d43f;
assign v86c49c = DEQ_p & v86b3a2 | !DEQ_p & v8ca5b3;
assign v8cab17 = StoB_REQ0_p & v8c9aa6 | !StoB_REQ0_p & !v844f91;
assign v8c9e60 = ENQ_p & v844f91 | !ENQ_p & v8cabac;
assign v85e833 = jx1_p & v862e4a | !jx1_p & !v8b31a9;
assign v8594ba = BtoR_REQ1_p & v865230 | !BtoR_REQ1_p & v85d413;
assign v8ca9fa = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9d;
assign v860b28 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v8c9917;
assign v8cab33 = DEQ_p & v844f91 | !DEQ_p & v86117f;
assign v8ca8ca = RtoB_ACK1_p & v8cac23 | !RtoB_ACK1_p & v86d647;
assign v8ca4e9 = DEQ_p & v8c95d7 | !DEQ_p & v8caa29;
assign v8cab34 = jx0_p & v85d451 | !jx0_p & !v861969;
assign v8caab9 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844fad;
assign v8622a3 = StoB_REQ2_p & v86b132 | !StoB_REQ2_p & !v8661bc;
assign v85e30e = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & v8caa1a;
assign v86d753 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8ca9ef;
assign v86d74c = StoB_REQ2_p & v89afb5 | !StoB_REQ2_p & !v844fad;
assign v8cacbd = ENQ_p & v8690d8 | !ENQ_p & v8691f7;
assign v8ca9f4 = RtoB_ACK1_p & v861aba | !RtoB_ACK1_p & v8693db;
assign v8cab4b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v8cac2e = jx1_p & v8caa0f | !jx1_p & v8b3167;
assign v8cab08 = jx2_p & v86d3d9 | !jx2_p & v86d231;
assign v8cabc1 = EMPTY_p & v861bd6 | !EMPTY_p & v865d58;
assign v8ca8b1 = ENQ_p & v868e55 | !ENQ_p & !v8621d8;
assign v8ca00c = EMPTY_p & v86d1e7 | !EMPTY_p & v860a1c;
assign v866456 = jx1_p & v8b69a7 | !jx1_p & v8cac32;
assign v862881 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v868f18;
assign v86c801 = ENQ_p & v866c03 | !ENQ_p & v85f3fa;
assign v8caa02 = BtoS_ACK1_p & v844f9c | !BtoS_ACK1_p & !v8c9a79;
assign v868f7d = EMPTY_p & v88d120 | !EMPTY_p & v88d12d;
assign v869a08 = jx2_p & v8c8cdb | !jx2_p & !v844f91;
assign v861980 = stateG7_1_p & v866606 | !stateG7_1_p & v864506;
assign v869361 = stateG7_1_p & v8ca7a6 | !stateG7_1_p & !v844f91;
assign v8712d2 = EMPTY_p & v86698a | !EMPTY_p & !v8cacde;
assign v8caaf0 = jx1_p & v88cf5c | !jx1_p & v844f91;
assign v85cdba = EMPTY_p & v844f91 | !EMPTY_p & v8caa81;
assign v85e2a3 = DEQ_p & v867a99 | !DEQ_p & v85e95d;
assign v86b125 = BtoS_ACK0_p & v8cab71 | !BtoS_ACK0_p & v8ca9f7;
assign v8cac03 = DEQ_p & v8cab07 | !DEQ_p & v8ca9ea;
assign v8caa57 = jx0_p & v861f69 | !jx0_p & v869b57;
assign v861d73 = ENQ_p & v8cac43 | !ENQ_p & v86621a;
assign v85d22b = DEQ_p & v8caa52 | !DEQ_p & v867417;
assign v852625 = jx2_p & v8cab4b | !jx2_p & v86a607;
assign v8caaae = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8cabcf;
assign v8cac4f = EMPTY_p & v844f91 | !EMPTY_p & !v86dae3;
assign v8640bb = jx1_p & v87132e | !jx1_p & !v85e8c1;
assign v8a749d = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v866a61;
assign v8cad66 = BtoS_ACK1_p & v86c73b | !BtoS_ACK1_p & v8caa8b;
assign v8cab9a = jx1_p & v844f99 | !jx1_p & !v865cd4;
assign v865319 = jx0_p & v8ca937 | !jx0_p & v86921b;
assign v8677e5 = DEQ_p & v8cab07 | !DEQ_p & v86b9e6;
assign v8698ed = StoB_REQ1_p & v8cab9f | !StoB_REQ1_p & v8caa11;
assign v866ad5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8450db;
assign v861fb9 = EMPTY_p & v8cac86 | !EMPTY_p & v8caa57;
assign v86b9e6 = EMPTY_p & v86607a | !EMPTY_p & !v8c9b09;
assign v8caa0d = EMPTY_p & v844f91 | !EMPTY_p & v8cac0a;
assign v88d132 = stateG7_1_p & v86494d | !stateG7_1_p & v8cac7a;
assign v8ca86e = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v86b108;
assign v861e9b = StoB_REQ1_p & v8794d1 | !StoB_REQ1_p & v8858bf;
assign v861d50 = EMPTY_p & v86191e | !EMPTY_p & !v862031;
assign v8ca153 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cac1f;
assign v86754b = StoB_REQ1_p & v85d86a | !StoB_REQ1_p & v868c2a;
assign v85e2c9 = jx1_p & v85cf1e | !jx1_p & v85a733;
assign v869e27 = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v8ca5f4;
assign v866940 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8450db;
assign v8caa39 = jx1_p & v860c87 | !jx1_p & v868d0a;
assign v85d924 = EMPTY_p & v8cac06 | !EMPTY_p & v860a1c;
assign v867cf7 = stateG7_1_p & v86702e | !stateG7_1_p & v861d73;
assign v8cabca = jx2_p & v861794 | !jx2_p & !v8cac6d;
assign v85e872 = jx2_p & v865321 | !jx2_p & !v8cab4b;
assign v8692bc = jx0_p & v864a04 | !jx0_p & v8610eb;
assign v89afd9 = BtoR_REQ1_p & v85f39d | !BtoR_REQ1_p & v8cabe1;
assign v8663d1 = jx0_p & v866cf1 | !jx0_p & v866456;
assign v88656a = jx1_p & v862e4a | !jx1_p & !v866655;
assign v85e544 = BtoR_REQ1_p & v86a8e7 | !BtoR_REQ1_p & v8cab75;
assign v8caa21 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v85cdc2;
assign v8697ea = ENQ_p & v8cabd8 | !ENQ_p & v8cac13;
assign v8caa83 = jx2_p & v86d805 | !jx2_p & v8cab3e;
assign v867170 = jx2_p & v844f91 | !jx2_p & !v852627;
assign v859567 = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v867ef1;
assign v869380 = StoB_REQ2_p & v85d750 | !StoB_REQ2_p & v8686e5;
assign v868b0c = jx1_p & v8ca61e | !jx1_p & v86797e;
assign v8cac11 = jx0_p & v85bdd0 | !jx0_p & !v86903b;
assign v8c9c75 = stateG7_1_p & v86864b | !stateG7_1_p & v89c755;
assign v85e12e = BtoS_ACK1_p & v844f9c | !BtoS_ACK1_p & v8ca9e9;
assign v85d772 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caafd;
assign v85d8cc = RtoB_ACK1_p & v8647c1 | !RtoB_ACK1_p & v8cab29;
assign v865f16 = jx2_p & v86911f | !jx2_p & v85cf1e;
assign v8ca345 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v869197;
assign v85d34f = jx0_p & v86b7cd | !jx0_p & v8caa1d;
assign v8c9aee = RtoB_ACK0_p & v8682bf | !RtoB_ACK0_p & v861980;
assign v844f9c = StoB_REQ3_n & v844f91 | !StoB_REQ3_n & !v844f91;
assign v8caac6 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v86ac9b;
assign v85d6e1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8692e8;
assign v8cac0b = jx2_p & v85cf1e | !jx2_p & v8612b9;
assign v85dece = EMPTY_p & v86c701 | !EMPTY_p & v8cacff;
assign v8c9a18 = RtoB_ACK0_p & v86b7d3 | !RtoB_ACK0_p & v8594ba;
assign v86aebe = jx1_p & v8cac6d | !jx1_p & !v8c9e27;
assign v8cabdf = jx1_p & v869dc6 | !jx1_p & !v86665f;
assign v894074 = FULL_p & v844f91 | !FULL_p & !v8c9a6e;
assign v86a710 = StoB_REQ2_p & v8660b6 | !StoB_REQ2_p & !v86a6a1;
assign v8c9cbc = ENQ_p & v866c03 | !ENQ_p & v8cacd7;
assign v85fb9d = ENQ_p & v868e55 | !ENQ_p & !v8cab77;
assign v86908e = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v86188b;
assign v86981f = ENQ_p & v867c81 | !ENQ_p & v852940;
assign v88d120 = jx0_p & v8ca937 | !jx0_p & v8c9b26;
assign v866c47 = jx0_p & v85d919 | !jx0_p & !v8cac2e;
assign v86890b = jx2_p & v85cf1e | !jx2_p & v85da6a;
assign v867b20 = jx0_p & v8cab32 | !jx0_p & v8cac1a;
assign v864ac7 = jx2_p & v8ca380 | !jx2_p & v844f91;
assign v85e491 = EMPTY_p & v867b20 | !EMPTY_p & v86884e;
assign v85d73d = StoB_REQ2_p & v8678af | !StoB_REQ2_p & !v85164d;
assign v868f18 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844fab;
assign v8caa18 = stateG12_p & v86b50c | !stateG12_p & !v864b72;
assign v8caa6e = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v86b72d;
assign v86badb = EMPTY_p & v866c47 | !EMPTY_p & v867a99;
assign v86aff9 = jx0_p & v868b0c | !jx0_p & !v85bb82;
assign v8cacf4 = jx0_p & v8c9b72 | !jx0_p & !v86490e;
assign v8caa56 = jx1_p & v86b125 | !jx1_p & !v8cab37;
assign v8c97df = EMPTY_p & v85db20 | !EMPTY_p & v85e743;
assign v8cabd0 = DEQ_p & v86b799 | !DEQ_p & v8c9ec8;
assign v8c9b26 = jx1_p & v8caac1 | !jx1_p & !v8cabca;
assign v8c9bb8 = jx2_p & v8caae9 | !jx2_p & v86113b;
assign v8c9696 = StoB_REQ1_p & v862264 | !StoB_REQ1_p & v86989e;
assign v86b108 = StoB_REQ0_p & v8caad3 | !StoB_REQ0_p & v8cab1a;
assign v8cabb4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cac76;
assign v8b31a9 = jx2_p & v865707 | !jx2_p & !v8cac6d;
assign v85e228 = jx2_p & v8cac6d | !jx2_p & v8ca693;
assign v879471 = FULL_p & v844f91 | !FULL_p & !v85de99;
assign v86a56e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8674af;
assign v86a8e7 = stateG7_1_p & v85d30e | !stateG7_1_p & v8caa86;
assign v861c01 = jx0_p & v851272 | !jx0_p & v8452cd;
assign v85f4ce = EMPTY_p & v8caba7 | !EMPTY_p & v85e6fc;
assign v86b22a = StoB_REQ2_p & v865dfa | !StoB_REQ2_p & v8699ec;
assign v866357 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v867be8;
assign v8cab7b = jx0_p & v8cab55 | !jx0_p & v86d061;
assign v85e5ff = DEQ_p & v8cace0 | !DEQ_p & v861d50;
assign v89409f = RtoB_ACK0_p & v85d1fb | !RtoB_ACK0_p & v860d7c;
assign v85cf1e = BtoS_ACK0_p & v85e30d | !BtoS_ACK0_p & v8ca9de;
assign v8672bb = jx2_p & v85c82e | !jx2_p & v865edc;
assign v8c95d0 = FULL_p & v85d221 | !FULL_p & v8cab26;
assign v88cf5c = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8ca9e8;
assign v85d3a1 = jx1_p & v844f99 | !jx1_p & v8cab6e;
assign v86c854 = stateG7_1_p & v8ca8ca | !stateG7_1_p & v8c95e9;
assign v860c8a = jx1_p & v86d5c8 | !jx1_p & v844f91;
assign v866b4c = EMPTY_p & v844f91 | !EMPTY_p & v879471;
assign v88d17c = BtoR_REQ0_p & v8c9aee | !BtoR_REQ0_p & v8ca9e6;
assign v86550b = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8caa91;
assign v8a604c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cac2d;
assign v861494 = jx1_p & v861d1f | !jx1_p & v8cac85;
assign v8caad9 = stateG7_1_p & v8caa55 | !stateG7_1_p & !v844f91;
assign v8caa8f = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v869990;
assign v865efb = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86a710;
assign v8ca3c8 = jx2_p & v86757f | !jx2_p & !v85c5d4;
assign v869147 = StoB_REQ1_p & v85cdfc | !StoB_REQ1_p & v861374;
assign v8614bb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e87a;
assign v8cac0d = BtoS_ACK0_p & v86ac9b | !BtoS_ACK0_p & v8caa15;
assign v85f3d4 = jx1_p & v8cac8d | !jx1_p & v865f16;
assign v85e046 = ENQ_p & v86817a | !ENQ_p & v89c737;
assign v867c96 = DEQ_p & v860a1c | !DEQ_p & v85d924;
assign v8cacd7 = DEQ_p & v8cab57 | !DEQ_p & v8caa1e;
assign v866205 = DEQ_p & v8cac70 | !DEQ_p & v8caca5;
assign v8660b8 = BtoS_ACK0_p & v8cab3d | !BtoS_ACK0_p & v86c5ef;
assign v8caa3c = EMPTY_p & v8cac10 | !EMPTY_p & v8c95d7;
assign v861b86 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8607fe;
assign v864a04 = jx1_p & v8666db | !jx1_p & !v8cacca;
assign v8c9cc5 = DEQ_p & v8cab9d | !DEQ_p & v8cab61;
assign v8caaec = BtoS_ACK1_p & v8cac4a | !BtoS_ACK1_p & v861d36;
assign v8620d1 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v85c6d8;
assign v86b799 = jx0_p & v866cf1 | !jx0_p & v8cab21;
assign v8caa76 = DEQ_p & v8ca9f0 | !DEQ_p & v85f48d;
assign v86816d = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v86921e;
assign v8cab29 = ENQ_p & v869284 | !ENQ_p & !v8ca9af;
assign v89c755 = ENQ_p & v8cac42 | !ENQ_p & !v8cac3d;
assign v868ae9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8649c1;
assign v866b27 = jx2_p & v869448 | !jx2_p & !v866940;
assign v85f4c4 = StoB_REQ2_p & v861ecc | !StoB_REQ2_p & !v844f91;
assign v868b32 = DEQ_p & v86a60b | !DEQ_p & v866d6a;
assign v852627 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v8cab74 = jx1_p & v8caa8f | !jx1_p & !v860a37;
assign v8ca71c = BtoS_ACK1_p & v86c73b | !BtoS_ACK1_p & v85e0d5;
assign v8caa5a = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8cab9f;
assign v861fc9 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v8cab72;
assign v8caa48 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v86d130;
assign v89b000 = jx2_p & v8cac6d | !jx2_p & v867220;
assign v8cabd7 = DEQ_p & v8cacd0 | !DEQ_p & v86349c;
assign v869f33 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e4fc;
assign v85d7eb = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cab04;
assign v85e6c3 = BtoS_ACK0_p & v8cab3d | !BtoS_ACK0_p & v8ca1f2;
assign v86974a = jx2_p & v844f91 | !jx2_p & v85da6a;
assign v86b4d5 = StoB_REQ1_p & v86d130 | !StoB_REQ1_p & v8667bd;
assign v85506c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v866834;
assign v86c57f = ENQ_p & v86817a | !ENQ_p & v844f91;
assign v866037 = jx0_p & v861e53 | !jx0_p & !v8caac9;
assign v86ba19 = BtoR_REQ1_p & v8ca78f | !BtoR_REQ1_p & v868cbc;
assign v8ca380 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8677dc;
assign v86757f = BtoS_ACK0_p & v8c7b0b | !BtoS_ACK0_p & v8cac5c;
assign v8ca9cd = jx0_p & v85f4e5 | !jx0_p & v85d3a1;
assign v8caa37 = EMPTY_p & v865319 | !EMPTY_p & !v867957;
assign v869e35 = jx2_p & v86d087 | !jx2_p & v85cf1e;
assign BtoS_ACK4_n = !v8858c9;
assign v85c6d8 = StoB_REQ0_p & v86d753 | !StoB_REQ0_p & v8ca1e1;
assign v861ea1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86a56e;
assign v8b2a29 = BtoR_REQ0_p & v8cac07 | !BtoR_REQ0_p & v86a7da;
assign v8c9942 = StoB_REQ1_p & v8cab9f | !StoB_REQ1_p & v8cac4a;
assign v8cac85 = jx2_p & v85e922 | !jx2_p & !v8caae9;
assign v85dd97 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e569;
assign v8cabde = jx0_p & v8c9e09 | !jx0_p & !v8c9eb5;
assign v8caa58 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caa61;
assign BtoR_REQ1_n = !v8b69e1;
assign v8cab9f = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v867bc5;
assign v85f3f5 = jx2_p & v8688ca | !jx2_p & v86d803;
assign v8ca9d4 = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & v844f91;
assign v8caa45 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8caa06;
assign v85d80e = jx1_p & v860c87 | !jx1_p & v85e872;
assign v867cbe = BtoS_ACK0_p & v862264 | !BtoS_ACK0_p & v8cab39;
assign v8cabe8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8696ce;
assign v869990 = StoB_REQ0_p & v8ca21b | !StoB_REQ0_p & v8682f7;
assign v8caa66 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caab9;
assign v8cacca = jx2_p & v8cac6d | !jx2_p & v844f91;
assign BtoS_ACK2_n = !v8a7515;
assign v844f9d = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v844f91;
assign v8650b2 = jx1_p & v860e50 | !jx1_p & !v86d231;
assign v8647c0 = BtoS_ACK0_p & v8c9805 | !BtoS_ACK0_p & v8682bd;
assign v8cac32 = jx2_p & v85e55a | !jx2_p & !v85c5d4;
assign v8cacd5 = jx0_p & v85f35c | !jx0_p & v844f91;
assign v85db6f = BtoS_ACK0_p & v8cac4a | !BtoS_ACK0_p & v85dc07;
assign v85ceb3 = ENQ_p & v8cab63 | !ENQ_p & v8ca4e9;
assign v8617fa = BtoS_ACK3_p & v86ab8a | !BtoS_ACK3_p & v86b132;
assign v8cab4e = BtoS_ACK0_p & v861ecc | !BtoS_ACK0_p & v866b1d;
assign v868467 = DEQ_p & v8cab57 | !DEQ_p & v8caa79;
assign v864506 = ENQ_p & v8cad4e | !ENQ_p & !v8cab52;
assign v861b4d = DEQ_p & v8cabec | !DEQ_p & v8cac84;
assign v8667ba = jx1_p & v8cac6d | !jx1_p & v868120;
assign v85db7d = stateG7_1_p & v8caa26 | !stateG7_1_p & v8cacdb;
assign v8c9bd1 = BtoS_ACK0_p & v8cab9f | !BtoS_ACK0_p & v868ae9;
assign v855530 = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v8cac02;
assign v85e4c8 = EMPTY_p & v8cac10 | !EMPTY_p & v8ca695;
assign v86c702 = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v8caad6;
assign v867507 = ENQ_p & v8cabd8 | !ENQ_p & v857c24;
assign v85e18e = jx0_p & v8648c8 | !jx0_p & v844f91;
assign v86b9c5 = EMPTY_p & v86d23a | !EMPTY_p & v8ca441;
assign v8ca018 = jx0_p & v8caaed | !jx0_p & !v86a61f;
assign v86b70b = BtoS_ACK0_p & v8c9805 | !BtoS_ACK0_p & v8cab70;
assign v8ca2a1 = EMPTY_p & v8ca399 | !EMPTY_p & v8ca695;
assign v85e24b = BtoR_REQ1_p & v86d6f9 | !BtoR_REQ1_p & v8683f7;
assign v85df63 = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v86d58d;
assign v86770a = RtoB_ACK0_p & v86a6ed | !RtoB_ACK0_p & v8c7b53;
assign v8cab88 = jx2_p & v8660b8 | !jx2_p & !v8caae9;
assign v8caabc = jx1_p & v85f7ba | !jx1_p & v85e78a;
assign v8caacd = EMPTY_p & v86698a | !EMPTY_p & v868f67;
assign v8cab3e = BtoS_ACK0_p & v85d43c | !BtoS_ACK0_p & v8c9917;
assign v85d28e = jx1_p & v844f9b | !jx1_p & !v85cf1e;
assign v8cac7e = DEQ_p & v8caa57 | !DEQ_p & v8c9c9f;
assign v8cacab = DEQ_p & v844f91 | !DEQ_p & v8ca6b5;
assign v8c9753 = jx0_p & v864a04 | !jx0_p & v8cab9a;
assign v85e2d7 = jx0_p & v89b002 | !jx0_p & v844fa7;
assign v866880 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v86294e;
assign v8cac3e = ENQ_p & v865e4b | !ENQ_p & v867c16;
assign v864207 = BtoR_REQ1_p & v8c9c75 | !BtoR_REQ1_p & v8b29f7;
assign v86d63a = ENQ_p & v8cac43 | !ENQ_p & v85e2a3;
assign v8cacc8 = ENQ_p & v8ca8b9 | !ENQ_p & v860d73;
assign v8674af = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v86c5c8;
assign v8caba9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8610ac;
assign v8653c0 = EMPTY_p & v866c47 | !EMPTY_p & v8673d4;
assign v8cac20 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8cacaa;
assign v860a1c = jx0_p & v8cac4b | !jx0_p & v8452cd;
assign v8c9a1b = RtoB_ACK0_p & v86d05a | !RtoB_ACK0_p & v861908;
assign v8ca295 = BtoS_ACK0_p & v8caa5a | !BtoS_ACK0_p & v86af4a;
assign v8cab2d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ca849;
assign v8caab8 = DEQ_p & v8c7b49 | !DEQ_p & v8cab5c;
assign v8671ac = StoB_REQ0_p & v8c9aa6 | !StoB_REQ0_p & !v85f3d3;
assign v867c81 = DEQ_p & v8cac11 | !DEQ_p & v85f4ce;
assign v8c9b72 = jx1_p & v86b70b | !jx1_p & v8c9bb8;
assign v8689a5 = jx2_p & v8cab3e | !jx2_p & v86889a;
assign v866655 = jx2_p & v866880 | !jx2_p & !v8cac6d;
assign v8686e5 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8cab1c;
assign v8ca441 = jx0_p & v869419 | !jx0_p & v8caa39;
assign v8cab1c = StoB_REQ3_p & v8ca9fa | !StoB_REQ3_p & v844f91;
assign v857ca8 = StoB_REQ2_p & v844fab | !StoB_REQ2_p & !v844f91;
assign v866d60 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v8622a3;
assign v867ef1 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8cab19;
assign v869ec7 = BtoR_REQ1_p & v85e63e | !BtoR_REQ1_p & v8caa2b;
assign v85dbee = EMPTY_p & v844f91 | !EMPTY_p & v8c95d0;
assign v865f9a = EMPTY_p & v869065 | !EMPTY_p & v8666cf;
assign v8691f9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e09a;
assign v866420 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cace5;
assign v86d61d = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v86d092;
assign v85e55a = BtoS_ACK0_p & v8c7b0b | !BtoS_ACK0_p & v8cac72;
assign v8caa81 = jx0_p & v844f91 | !jx0_p & v8667f6;
assign v8c9b67 = StoB_REQ0_p & v861fc9 | !StoB_REQ0_p & v844f91;
assign v85f521 = jx1_p & v844f91 | !jx1_p & v8cac05;
assign v844fa5 = EMPTY_p & v844f91 | !EMPTY_p & !v844f91;
assign v8cabc0 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v86b4d5;
assign v8c9ce7 = jx0_p & v8c9b72 | !jx0_p & !v8c9eb5;
assign v86540f = DEQ_p & v844f91 | !DEQ_p & v86863b;
assign v861409 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8ca9de;
assign v8ca7ed = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85e1fe;
assign v867844 = BtoS_ACK0_p & v8cab9f | !BtoS_ACK0_p & v85e95a;
assign v867ed2 = jx1_p & v85da6a | !jx1_p & v864080;
assign v8caaf1 = DEQ_p & v8caa52 | !DEQ_p & v86d7ce;
assign v85f4e5 = jx1_p & v8c9e5e | !jx1_p & !v86665f;
assign v86631f = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & !v844f91;
assign v866c98 = EMPTY_p & v85cec5 | !EMPTY_p & v8ca695;
assign v8cac45 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c9b67;
assign v85dc69 = StoB_REQ2_p & v8678af | !StoB_REQ2_p & !v844f91;
assign v85daff = BtoS_ACK3_p & v8cab01 | !BtoS_ACK3_p & v844f9b;
assign v868377 = jx2_p & v85df63 | !jx2_p & v8caa3a;
assign v8b69cf = EMPTY_p & v867b20 | !EMPTY_p & v85d485;
assign v868569 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v85d73d;
assign v8caa60 = FULL_p & v865bf0 | !FULL_p & v86aff9;
assign v866d4f = DEQ_p & v8c95d7 | !DEQ_p & v8caa3c;
assign v8c7b49 = jx0_p & v8650b2 | !jx0_p & v87947b;
assign v8caccf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v866f76;
assign v8cab28 = DEQ_p & v8cab9d | !DEQ_p & v8712d2;
assign v862200 = jx1_p & v86b50c | !jx1_p & v86837b;
assign v8caa74 = jx1_p & v867d26 | !jx1_p & v8cacba;
assign v8c7b53 = BtoR_REQ1_p & v866610 | !BtoR_REQ1_p & v8ca9e0;
assign v8ca6b5 = EMPTY_p & v844f91 | !EMPTY_p & v866aae;
assign v8ca9e8 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v863955;
assign v8c9cac = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v86631f;
assign v8cabec = jx0_p & v85d28e | !jx0_p & !v85e2c9;
assign v8cab07 = jx0_p & v8650b2 | !jx0_p & v8683f9;
assign v8ca9f7 = StoB_REQ0_p & v86d7d4 | !StoB_REQ0_p & v865fe1;
assign v8cac71 = StoB_REQ0_p & v86294e | !StoB_REQ0_p & v8cac1d;
assign v8b3161 = DEQ_p & v8c7b49 | !DEQ_p & v85206c;
assign v86d647 = ENQ_p & v86c49c | !ENQ_p & v8b69b8;
assign v8cac99 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v863955;
assign v868936 = StoB_REQ2_p & v8caab9 | !StoB_REQ2_p & v86631f;
assign v8cab0e = jx0_p & v8cac0c | !jx0_p & !v8ca0bd;
assign v8588a0 = StoB_REQ1_p & v85f557 | !StoB_REQ1_p & v863955;
assign v85d230 = jx2_p & v86a84a | !jx2_p & !v8cab4b;
assign v8619cf = jx0_p & v8caa74 | !jx0_p & v867d26;
assign v86ba45 = ENQ_p & v8cad4e | !ENQ_p & !v86c4e5;
assign v8cacc6 = jx1_p & v8ca86e | !jx1_p & !v8cab2f;
assign v8cabc7 = DEQ_p & v8663d1 | !DEQ_p & v8a74fd;
assign v865de8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c9811;
assign v866b6f = ENQ_p & v861c01 | !ENQ_p & v86900f;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v85d413 = stateG7_1_p & v8caa77 | !stateG7_1_p & v85e224;
assign v85f35c = jx1_p & v844f91 | !jx1_p & v8caab4;
assign v8c9733 = stateG7_1_p & v86c581 | !stateG7_1_p & v8ca9f5;
assign v8caa08 = jx2_p & v867cbe | !jx2_p & v85cf1e;
assign v85e03e = EMPTY_p & v86d23a | !EMPTY_p & v8cac93;
assign v8ca9c1 = jx0_p & v8ca3d4 | !jx0_p & !v85d448;
assign v8794e5 = BtoR_REQ0_p & v894033 | !BtoR_REQ0_p & v864050;
assign v861dcc = EMPTY_p & v85d9e0 | !EMPTY_p & v8c9ea3;
assign v8ca0b4 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v85e30d;
assign v86900f = DEQ_p & v860a1c | !DEQ_p & v8ca00c;
assign v85a021 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8cab0a;
assign v8caac1 = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v865de8;
assign v8cabd2 = ENQ_p & v8690d8 | !ENQ_p & v844f91;
assign v8caa6b = DEQ_p & v8ca9f0 | !DEQ_p & v8cacdf;
assign v8cac7c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8450db;
assign v86989e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v86ac5d;
assign v85ac07 = jx1_p & v86889b | !jx1_p & v8679a8;
assign v8caad6 = StoB_REQ1_p & v8cac02 | !StoB_REQ1_p & v862264;
assign v865036 = jx2_p & v8ca295 | !jx2_p & v865edc;
assign v861d5f = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v8ca32a;
assign v869dc6 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8cab70;
assign v8cac43 = DEQ_p & v8cac11 | !DEQ_p & v8ca48a;
assign v865787 = EMPTY_p & v88d14f | !EMPTY_p & v8654cb;
assign v8cac69 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v855346;
assign v861969 = jx1_p & v8cac8d | !jx1_p & v85a733;
assign v86349c = EMPTY_p & v8cacd0 | !EMPTY_p & v8a868e;
assign v86864b = ENQ_p & v8cac42 | !ENQ_p & !v8ca753;
assign v8caa4a = ENQ_p & v867697 | !ENQ_p & !v85c6f5;
assign v85dbcd = BtoS_ACK2_p & v8caa43 | !BtoS_ACK2_p & v8cabe6;
assign v864b72 = jx2_p & v85c5d4 | !jx2_p & !v86b50c;
assign v85f2a4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8caa15;
assign v86884e = jx0_p & v8ca701 | !jx0_p & v8cab21;
assign v8caaa8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v869e27;
assign v8667cc = jx1_p & v867ba8 | !jx1_p & v8cab88;
assign v85e61f = jx0_p & v8cab9b | !jx0_p & v86b50c;
assign v8ca8b9 = DEQ_p & v8619cf | !DEQ_p & v867d26;
assign v862fc7 = jx1_p & v844f91 | !jx1_p & v868905;
assign v85f3a3 = ENQ_p & v844f91 | !ENQ_p & v86540f;
assign v8caa3a = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v866420;
assign v86921e = StoB_REQ2_p & v85d750 | !StoB_REQ2_p & v8cacbe;
assign v8b69a7 = BtoS_ACK0_p & v8caa4d | !BtoS_ACK0_p & v8caa5d;
assign v85164d = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8678af;
assign v8caab0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cabcb;
assign v861dac = DEQ_p & v844f91 | !DEQ_p & v85e1f9;
assign v86665f = jx2_p & v844f91 | !jx2_p & !v85e84a;
assign v8ca78f = stateG7_1_p & v85dade | !stateG7_1_p & !v844f91;
assign v8cac06 = jx0_p & v8c9c26 | !jx0_p & v8452cd;
assign v8cab97 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v863e15;
assign v85db20 = jx0_p & v8cacaf | !jx0_p & v86b5da;
assign v8c9cae = StoB_REQ2_p & v8678af | !StoB_REQ2_p & !v8c9c7c;
assign v86c73b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8caa43;
assign v866ba0 = StoB_REQ2_p & v89afb5 | !StoB_REQ2_p & !v86631f;
assign v8a74b4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v869147;
assign v8caba4 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v86d1b3;
assign v86b838 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86ba15;
assign v8ca115 = StoB_REQ1_p & v85e1fe | !StoB_REQ1_p & v85c2e5;
assign v8cab9d = jx0_p & v85d28e | !jx0_p & !v8caac9;
assign v86837b = stateG12_p & v86b50c | !stateG12_p & v861522;
assign v8cac82 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8660a4;
assign v8cacbe = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v85d750;
assign v8cab56 = jx2_p & v8caae9 | !jx2_p & !v844f91;
assign v85d906 = BtoS_ACK0_p & v8cab19 | !BtoS_ACK0_p & !v8b31ca;
assign v866b78 = EMPTY_p & v8cab34 | !EMPTY_p & v866037;
assign v86b711 = BtoS_ACK0_p & v8cab9f | !BtoS_ACK0_p & v85e249;
assign v868f67 = FULL_p & v8caab6 | !FULL_p & v8ca9c1;
assign v8c7b0b = StoB_REQ1_p & v86c73b | !StoB_REQ1_p & v844f91;
assign v86d58d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v868d58;
assign v85f39d = stateG7_1_p & v86589e | !stateG7_1_p & v8cac0f;
assign v8cab87 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cab2b;
assign v861903 = jx2_p & v8609fc | !jx2_p & v865edc;
assign v861e4f = EMPTY_p & v866d78 | !EMPTY_p & v865bf0;
assign v88589b = jx1_p & v844f91 | !jx1_p & v8ca648;
assign v86d276 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8617fa;
assign v8ca9e2 = ENQ_p & v85daa3 | !ENQ_p & !v86d136;
assign v8ca472 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v85d3d5;
assign v8caa43 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9d;
assign v868fbe = stateG12_p & v8c9ed1 | !stateG12_p & !v86652d;
assign v86150f = stateG7_1_p & v86a618 | !stateG7_1_p & v8ca374;
assign v8cac07 = RtoB_ACK0_p & v8ca8b1 | !RtoB_ACK0_p & v85db7d;
assign v8ca84f = jx0_p & v8c984a | !jx0_p & v868f72;
assign v86a76c = jx1_p & v844f91 | !jx1_p & v861b6c;
assign v865f35 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e947;
assign v8cac5e = jx1_p & v8cacd3 | !jx1_p & !v86114b;
assign v8cacd8 = stateG12_p & v85e228 | !stateG12_p & v85ce98;
assign v8cacdd = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v8caa67;
assign v8940fd = jx1_p & v8b69a7 | !jx1_p & v86908c;
assign v8ca9ef = StoB_REQ2_p & v863955 | !StoB_REQ2_p & v8cac99;
assign v8450db = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v8cabac = DEQ_p & v844f91 | !DEQ_p & v867e47;
assign v85e1f9 = EMPTY_p & v844f91 | !EMPTY_p & v861166;
assign v86909b = jx2_p & v868317 | !jx2_p & !v866940;
assign v8637cb = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8c9811;
assign v8ca089 = BtoS_ACK0_p & v8cab19 | !BtoS_ACK0_p & v8680fe;
assign v8ca357 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8cab17;
assign v8cac77 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v869a67;
assign v85e95d = EMPTY_p & v86c461 | !EMPTY_p & v8673d4;
assign v875b43 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86a5ad;
assign v8cacb5 = jx0_p & v85b1cb | !jx0_p & v85e733;
assign v8caab6 = jx0_p & v8ca3d4 | !jx0_p & !v844f91;
assign v86d814 = jx1_p & v869baf | !jx1_p & !v86b02f;
assign v85ce85 = EMPTY_p & v8caa8c | !EMPTY_p & v844f91;
assign v8ca9de = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c9fa7;
assign v86652d = jx2_p & v844f91 | !jx2_p & v866940;
assign v8caaf7 = DEQ_p & v844f91 | !DEQ_p & v85cdba;
assign v89407e = DEQ_p & v8ca695 | !DEQ_p & v866c98;
assign v8678d9 = jx0_p & v868403 | !jx0_p & v86522b;
assign v8cabbd = StoB_REQ0_p & v8c9b51 | !StoB_REQ0_p & v8677dc;
assign v8c9f67 = StoB_REQ0_p & v8c9b51 | !StoB_REQ0_p & v85d6cf;
assign v8cab8c = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v86b22a;
assign v8caadb = jx0_p & v860ea5 | !jx0_p & v86889a;
assign v8cac9c = FULL_p & v85310f | !FULL_p & v8cac0a;
assign v8679ab = jx0_p & v8ca9eb | !jx0_p & v869b57;
assign v8613c9 = BtoS_ACK1_p & v8cac4a | !BtoS_ACK1_p & v8674bb;
assign v844fa7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v8cac15 = jx1_p & v844f91 | !jx1_p & v8caaa9;
assign v868ba7 = EMPTY_p & v844f91 | !EMPTY_p & !v86ae3e;
assign v8cac30 = jx1_p & v85cd74 | !jx1_p & v86665f;
assign v86608e = ENQ_p & v861c01 | !ENQ_p & v861290;
assign v8caaad = StoB_REQ1_p & v8caa61 | !StoB_REQ1_p & v868bb5;
assign v86a8cf = jx2_p & v85c5d4 | !jx2_p & v866ad5;
assign v861998 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caca2;
assign v8caa9d = EMPTY_p & v85e8c7 | !EMPTY_p & v8a868e;
assign v8680fe = StoB_REQ0_p & v86d5fc | !StoB_REQ0_p & v85dee9;
assign v85e110 = jx1_p & v8caa40 | !jx1_p & v8c9ce3;
assign v8caa67 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & !v86b132;
assign v8cac1d = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v861e9b;
assign v8cacd3 = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v860ec7;
assign v8ca014 = jx1_p & v85cf1e | !jx1_p & v869e35;
assign v86d6f9 = stateG7_1_p & v8cac53 | !stateG7_1_p & v866013;
assign v8651a5 = DEQ_p & v844f91 | !DEQ_p & v865791;
assign v865b89 = jx1_p & v844f91 | !jx1_p & !v865da5;
assign v867e47 = EMPTY_p & v8cac35 | !EMPTY_p & v844f91;
assign v85e143 = BtoS_ACK0_p & v8cab19 | !BtoS_ACK0_p & v8c9b86;
assign v89affe = jx2_p & v844f91 | !jx2_p & v867d26;
assign v85d881 = DEQ_p & v860a57 | !DEQ_p & v86840f;
assign v869112 = jx0_p & v8ca055 | !jx0_p & v86889a;
assign v8cab1d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cab9f;
assign v867a57 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v867080;
assign v85d81d = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v861405;
assign v8caa51 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v868f18;
assign v8693db = ENQ_p & v869dae | !ENQ_p & v85ce37;
assign v8ca615 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v86d322;
assign v8ca2af = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8c9ace;
assign v861c02 = ENQ_p & v8cad4e | !ENQ_p & !v85e6c0;
assign v8a6000 = RtoB_ACK0_p & v85ceb3 | !RtoB_ACK0_p & v868fd6;
assign v8cad96 = ENQ_p & v867697 | !ENQ_p & !v8cab28;
assign v85d6d7 = jx1_p & v8674b4 | !jx1_p & v86143d;
assign v8cab37 = jx2_p & v85dac9 | !jx2_p & v86d231;
assign v86538c = FULL_p & v844f91 | !FULL_p & v8cab0e;
assign v867763 = DEQ_p & v8c95d7 | !DEQ_p & v8ca2a1;
assign v8ca6af = RtoB_ACK0_p & v894103 | !RtoB_ACK0_p & v86d2a0;
assign v85e568 = DEQ_p & v8cab7b | !DEQ_p & v8641cf;
assign v86143d = jx2_p & v861ea1 | !jx2_p & v844f91;
assign v8cab03 = StoB_REQ0_p & v8c95c7 | !StoB_REQ0_p & v844f91;
assign v869631 = StoB_REQ1_p & v8caa61 | !StoB_REQ1_p & !v86b72d;
assign v8c9bfc = ENQ_p & v8cab76 | !ENQ_p & !v865404;
assign v8cab2f = jx2_p & v844f91 | !jx2_p & !v8cabff;
assign v86d3cb = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v85d43c;
assign v8cabe6 = BtoS_ACK3_p & v844f9b | !BtoS_ACK3_p & v85d53b;
assign v8cab25 = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v8674f7;
assign v8cab71 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v8cab19;
assign v8caa14 = BtoS_ACK3_p & v8caa43 | !BtoS_ACK3_p & v844f9b;
assign v8ca9f5 = ENQ_p & v8ca8b9 | !ENQ_p & v85ce37;
assign v85d97a = RtoB_ACK1_p & v8cac29 | !RtoB_ACK1_p & v84505f;
assign v8c9eb5 = jx1_p & v861d1f | !jx1_p & v8cab47;
assign v8cace5 = BtoS_ACK1_p & v86c73b | !BtoS_ACK1_p & v85e35c;
assign v8caaf3 = jx2_p & v8cac45 | !jx2_p & v8cab4b;
assign v865edc = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v844f95;
assign v86b06e = DEQ_p & v8cab57 | !DEQ_p & v8cabf0;
assign v861bd6 = jx0_p & v8cab32 | !jx0_p & v8cab21;
assign v867565 = jx2_p & v8cabe9 | !jx2_p & v844f91;
assign v8caa62 = StoB_REQ1_p & v8ca9ef | !StoB_REQ1_p & v863955;
assign v8ca23b = stateG12_p & v844fa7 | !stateG12_p & !v8caaef;
assign v8ca44e = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & !v868b0b;
assign v8649c5 = jx0_p & v8c9cad | !jx0_p & v869b57;
assign v85e1cb = jx1_p & v85f4cf | !jx1_p & v85de3b;
assign v8cac22 = jx0_p & v86b7cd | !jx0_p & v8cabcd;
assign v86b50c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fa9;
assign v8caaf5 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v86d276;
assign v8ca5e2 = DEQ_p & v860a57 | !DEQ_p & v8c9dd6;
assign v8cab2b = BtoS_ACK1_p & v86add5 | !BtoS_ACK1_p & v8cac3a;
assign v8ca300 = jx2_p & v844f91 | !jx2_p & !v868626;
assign v868bb5 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v86b7fd;
assign BtoR_REQ0_n = !v89b010;
assign v8ca315 = jx2_p & v8ca380 | !jx2_p & !v8cac6d;
assign v86922c = jx0_p & v8cacc6 | !jx0_p & v8452cd;
assign v8ca349 = jx2_p & v85c5d4 | !jx2_p & !v866940;
assign v85dee9 = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v86b05b;
assign v8cab76 = DEQ_p & v8ca096 | !DEQ_p & v865a01;
assign v875b45 = BtoR_REQ0_p & v8b2a0d | !BtoR_REQ0_p & v8674ab;
assign v86b725 = ENQ_p & v869284 | !ENQ_p & !v844f91;
assign v8452cd = jx1_p & v844f91 | !jx1_p & !v844f91;
assign v8cab6f = StoB_REQ1_p & v85e1fe | !StoB_REQ1_p & v868bd4;
assign v86d2a0 = stateG7_1_p & v8caafb | !stateG7_1_p & v86c517;
assign v866af3 = jx0_p & v868b0c | !jx0_p & !v8ca5f9;
assign v85ce9c = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cac5c;
assign v85d30e = ENQ_p & v868e55 | !ENQ_p & !v866d6c;
assign v8ca7a9 = BtoS_ACK0_p & v8cab3d | !BtoS_ACK0_p & v865dbb;
assign v8caa1a = StoB_REQ1_p & v8794d1 | !StoB_REQ1_p & v8cabcc;
assign v8cabea = ENQ_p & v8940e1 | !ENQ_p & v866c71;
assign v860bef = jx1_p & v8c9e5e | !jx1_p & v8cacb9;
assign v8613f4 = jx2_p & v844f91 | !jx2_p & v8450db;
assign v85e8ee = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8ca9ee;
assign v862e4a = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v8cace7;
assign v8caa9a = jx1_p & v867d26 | !jx1_p & v86888b;
assign v86859e = stateG12_p & v868282 | !stateG12_p & !v86665f;
assign v8ca737 = DEQ_p & v844f91 | !DEQ_p & v8caa0d;
assign v85d39c = jx2_p & v8a604c | !jx2_p & v8cab4b;
assign v8c9805 = StoB_REQ1_p & v8caa61 | !StoB_REQ1_p & v844f9b;
assign v8caa1e = EMPTY_p & v8ca84f | !EMPTY_p & v869992;
assign v8caa36 = jx1_p & v8cac69 | !jx1_p & v844f91;
assign v865d4b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86789d;
assign v867b2b = jx0_p & v8cac8e | !jx0_p & v8683f9;
assign v89c737 = DEQ_p & v844f91 | !DEQ_p & v867e4a;
assign v86522b = jx1_p & v85e484 | !jx1_p & v868377;
assign v86a6ed = BtoR_REQ1_p & v8c9607 | !BtoR_REQ1_p & v8ca9e0;
assign v8cab5d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8613c9;
assign v8697b7 = jx2_p & v8cab7c | !jx2_p & v8cab3e;
assign v86c517 = ENQ_p & v8cabd8 | !ENQ_p & v86d7f2;
assign v8caca1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8caa58;
assign v86674c = jx2_p & v844f91 | !jx2_p & v85e84a;
assign v844f9f = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v890c4a = jx1_p & v844f9c | !jx1_p & !v8613f4;
assign v868282 = jx2_p & v8c8cdb | !jx2_p & v85e84a;
assign v85d90c = BtoS_ACK3_p & v8caa43 | !BtoS_ACK3_p & v85d53b;
assign v86925d = StoB_REQ1_p & v85d73d | !StoB_REQ1_p & v8c9cae;
assign v8c9e5e = BtoS_ACK0_p & v844f9c | !BtoS_ACK0_p & v85e12e;
assign v85e85f = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & !v8c9bb0;
assign v86191e = jx0_p & v8ca9a6 | !jx0_p & v86d814;
assign v86d087 = BtoS_ACK0_p & v862264 | !BtoS_ACK0_p & v85d58f;
assign v8c984a = jx1_p & v861d5f | !jx1_p & v8c9bbf;
assign v86840f = EMPTY_p & v8ca018 | !EMPTY_p & v844f91;
assign v867be8 = StoB_REQ2_p & v844fab | !StoB_REQ2_p & v844f91;
assign v86639e = jx1_p & v8cac6d | !jx1_p & !v8ca315;
assign v8caa41 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85b56a;
assign v85bdd0 = jx1_p & v869497 | !jx1_p & v868fbe;
assign v8ca2c0 = BtoS_ACK0_p & v8cab19 | !BtoS_ACK0_p & v85e297;
assign v85cdad = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8c9805;
assign v86b72d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f9b;
assign v865d58 = FULL_p & v864dbb | !FULL_p & v860a0f;
assign v861171 = jx1_p & v87132e | !jx1_p & !v8caa83;
assign v85d8fe = DEQ_p & v8ca9f0 | !DEQ_p & v8caa37;
assign v869448 = BtoS_ACK0_p & v858cb9 | !BtoS_ACK0_p & v8cab87;
assign v866540 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v8c9aa6;
assign v8cac63 = ENQ_p & v8cac80 | !ENQ_p & v8c9aac;
assign v8688ca = BtoS_ACK0_p & v8c9811 | !BtoS_ACK0_p & v8c9b86;
assign v8cac8d = BtoS_ACK0_p & v85e30d | !BtoS_ACK0_p & v865d4b;
assign v8cabcb = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v844f91;
assign v86a6a1 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9b;
assign v8ca9cf = jx2_p & v8caccf | !jx2_p & v8a749d;
assign v8caa2b = ENQ_p & v8cac43 | !ENQ_p & v8caac0;
assign v8c9c59 = RtoB_ACK1_p & v85d1fb | !RtoB_ACK1_p & v8cab8e;
assign v8ca41e = stateG12_p & v89affe | !stateG12_p & v867d26;
assign v86889a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v868fc7;
assign v8940d7 = DEQ_p & v867a99 | !DEQ_p & v86badb;
assign v8658ac = jx2_p & v8cab3e | !jx2_p & !v860b28;
assign v8caa8b = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85f516;
assign v86d329 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v865ff9;
assign v8661e2 = DEQ_p & v844f91 | !DEQ_p & v86d813;
assign v86a905 = jx2_p & v85d81d | !jx2_p & v844f91;
assign v868f72 = jx1_p & v862e4a | !jx1_p & !v867010;
assign v869653 = jx2_p & v844f91 | !jx2_p & v8cabff;
assign v8caaff = jx1_p & v844f99 | !jx1_p & !v844f91;
assign v85de29 = EMPTY_p & v844f91 | !EMPTY_p & v8c9aca;
assign v868d0a = jx2_p & v8cab4e | !jx2_p & !v8cab4b;
assign v8caad4 = ENQ_p & v8cac43 | !ENQ_p & v867319;
assign v8cac00 = StoB_REQ2_p & v8caab9 | !StoB_REQ2_p & v844fad;
assign v8697c8 = ENQ_p & v8c9dae | !ENQ_p & !v8c9aea;
assign v857c24 = DEQ_p & v8663d1 | !DEQ_p & v8b69cf;
assign v8cac29 = ENQ_p & v86b2c2 | !ENQ_p & v8caaf7;
assign v85d91a = BtoS_ACK0_p & v86c73b | !BtoS_ACK0_p & v866420;
assign v865507 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v89afb5;
assign v860a57 = jx0_p & v8668d6 | !jx0_p & !v86116b;
assign v8cab6d = StoB_REQ1_p & v89afb5 | !StoB_REQ1_p & v856a93;
assign v8ca9ea = EMPTY_p & v8cab07 | !EMPTY_p & !v8caca0;
assign v869b15 = FULL_p & v8caab6 | !FULL_p & v85de99;
assign v8cacc5 = DEQ_p & v8c9ce7 | !DEQ_p & v85e185;
assign v8cac3d = DEQ_p & v8c7b49 | !DEQ_p & v8b317b;
assign v861e53 = jx1_p & v844f9b | !jx1_p & !v8ca9e3;
assign v86d231 = BtoS_ACK0_p & v8c9bb0 | !BtoS_ACK0_p & v8b31ca;
assign v8cab14 = stateG7_1_p & v8cac5d | !stateG7_1_p & v86d63a;
assign v8858bf = StoB_REQ2_p & v866964 | !StoB_REQ2_p & !v844f9b;
assign v868fd6 = stateG7_1_p & v866610 | !stateG7_1_p & v85ce75;
assign v857888 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v867bc5;
assign v8caa2e = RtoB_ACK0_p & v867cb8 | !RtoB_ACK0_p & v85e24b;
assign v85e81e = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85e5c6;
assign v860ab6 = ENQ_p & v8cabd7 | !ENQ_p & v867a28;
assign v8c97c4 = BtoS_ACK3_p & v8cab1c | !BtoS_ACK3_p & v8ca9fa;
assign v8cac7a = ENQ_p & v868b32 | !ENQ_p & !v8b3161;
assign v8ca742 = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v861279;
assign v867edf = BtoS_ACK0_p & v8691f2 | !BtoS_ACK0_p & v86ac7c;
assign v8ca9e4 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v86d5fc;
assign v85d58f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86c702;
assign v86753c = StoB_REQ0_p & v8677dc | !StoB_REQ0_p & v8ca44e;
assign v861374 = StoB_REQ2_p & v8ca9d4 | !StoB_REQ2_p & v844f91;
assign v8cab44 = jx0_p & v8c9dd4 | !jx0_p & v86a76c;
assign v8cab02 = ENQ_p & v8ca8b9 | !ENQ_p & v866d97;
assign v8cac93 = jx0_p & v86d411 | !jx0_p & v8caa39;
assign v869dae = DEQ_p & v8619cf | !DEQ_p & v86550b;
assign v86d05a = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v8caad9;
assign v8caa17 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v863955;
assign v8c9fa7 = BtoS_ACK1_p & v86ac9b | !BtoS_ACK1_p & v85e30d;
assign v85e138 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8cab42;
assign v8cac4e = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v8caa90;
assign v8ca32a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cab25;
assign v860d73 = DEQ_p & v8cab57 | !DEQ_p & v8c9f14;
assign v85e7b6 = jx1_p & v8647c0 | !jx1_p & v8cac49;
assign v8ca055 = jx1_p & v86889a | !jx1_p & v8ca9cb;
assign v868dd9 = jx1_p & v88cf5c | !jx1_p & !v867170;
assign v871300 = DEQ_p & v867a75 | !DEQ_p & v8cac6a;
assign v8cacff = jx0_p & v85dbc1 | !jx0_p & v8cabfe;
assign v8ca7e1 = jx0_p & v85f521 | !jx0_p & v866138;
assign v8caa79 = EMPTY_p & v8cabeb | !EMPTY_p & v8caa81;
assign v8cabf2 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v85c534;
assign v86ab8a = StoB_REQ3_p & v86b132 | !StoB_REQ3_p & !v844f9d;
assign v868c2a = StoB_REQ2_p & v8664cd | !StoB_REQ2_p & v844fad;
assign v86d1e7 = jx0_p & v869259 | !jx0_p & v8452cd;
assign v8cac21 = jx1_p & v844f99 | !jx1_p & !v865f9e;
assign v8caada = jx0_p & v868c4d | !jx0_p & !v865c5c;
assign v865d47 = BtoR_REQ1_p & v8c9733 | !BtoR_REQ1_p & v8940a7;
assign v85e233 = StoB_REQ2_p & v8caa06 | !StoB_REQ2_p & v8caa45;
assign v8c9b86 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85ddf2;
assign v85e249 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86d81c;
assign v85e164 = jx2_p & v8cac8f | !jx2_p & v8ca742;
assign v8cabb7 = DEQ_p & v860a57 | !DEQ_p & v8c7acf;
assign v861f9e = jx0_p & v85d28e | !jx0_p & !v8ca014;
assign v861436 = RtoB_ACK0_p & v8cab02 | !RtoB_ACK0_p & v8ca2fd;
assign v86b2c2 = DEQ_p & v867a75 | !DEQ_p & v867d26;
assign v86b1d8 = BtoS_ACK2_p & v8caa43 | !BtoS_ACK2_p & v85d53b;
assign v8ca6a1 = StoB_REQ1_p & v89afb5 | !StoB_REQ1_p & v866ba0;
assign v86117f = EMPTY_p & v844f91 | !EMPTY_p & !v861525;
assign v8caafc = DEQ_p & v844f91 | !DEQ_p & v8caca3;
assign v8a868e = jx0_p & v8c7b4e | !jx0_p & v844f91;
assign v8621d8 = DEQ_p & v8cacf4 | !DEQ_p & v86d7c8;
assign v86d061 = jx1_p & v844f99 | !jx1_p & v85d230;
assign v868626 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v852627;
assign v865859 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8cabf5;
assign v8c9811 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8cab19;
assign v86d5ab = jx0_p & v8cabdf | !jx0_p & !v85d6d7;
assign v8cacd1 = StoB_REQ1_p & v85d3d5 | !StoB_REQ1_p & v863955;
assign v85e5ed = ENQ_p & v8cabd8 | !ENQ_p & v8cabd0;
assign v8c0272 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caa11;
assign v85cdc2 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & !v86b72d;
assign v8b29f7 = stateG7_1_p & v8cabea | !stateG7_1_p & v86d602;
assign v8ca19f = jx2_p & v8691f9 | !jx2_p & v844f91;
assign v86c5c8 = StoB_REQ1_p & v8c973b | !StoB_REQ1_p & v86989e;
assign v85ddf2 = BtoS_ACK1_p & v8cab19 | !BtoS_ACK1_p & v844f91;
assign v86217d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85e81e;
assign v8caaab = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8ca3c3;
assign v8cacd6 = StoB_REQ3_p & v8ca9fa | !StoB_REQ3_p & v844f9d;
assign v8cab26 = jx0_p & v8c9dd4 | !jx0_p & v8caad2;
assign v868e55 = DEQ_p & v8cacd5 | !DEQ_p & v844f91;
assign v862321 = ENQ_p & v861c01 | !ENQ_p & v867c96;
assign v8cabe1 = ENQ_p & v869284 | !ENQ_p & !v8661e2;
assign v8674b4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8caa5d;
assign v8caa87 = jx1_p & v867ba8 | !jx1_p & v86bae1;
assign v8cace7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8637cb;
assign v8cad25 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8c9a57;
assign v8c973b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9d;
assign v85e045 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v868c92;
assign v8c9cbb = jx2_p & v866880 | !jx2_p & !v8cab4b;
assign v85c534 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85e233;
assign v868830 = RtoB_ACK1_p & v8ca17e | !RtoB_ACK1_p & v85e046;
assign v8ca354 = BtoS_ACK2_p & v867bc5 | !BtoS_ACK2_p & !v86b74a;
assign v87131b = jx1_p & v867ba8 | !jx1_p & v8cab47;
assign v863449 = jx1_p & v8cac6d | !jx1_p & v8c9bbf;
assign v868c92 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8caac6;
assign v86c4e5 = DEQ_p & v8647a2 | !DEQ_p & v865f0e;
assign v8b69ca = jx1_p & v866357 | !jx1_p & v868d0a;
assign v860bf2 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8cabe8;
assign v862256 = jx2_p & v8cac33 | !jx2_p & v86d231;
assign v865f9e = jx2_p & v86918c | !jx2_p & v844f91;
assign v8caa26 = RtoB_ACK1_p & v861809 | !RtoB_ACK1_p & v8cab9c;
assign v8caae1 = StoB_REQ2_p & v8660b6 | !StoB_REQ2_p & v85daff;
assign v8cac5b = DEQ_p & v8cacd0 | !DEQ_p & v85e03e;
assign BtoS_ACK1_n = !v8c7b59;
assign v8caa77 = RtoB_ACK1_p & v879497 | !RtoB_ACK1_p & v8c9ff6;
assign v86d2f5 = jx0_p & v8caace | !jx0_p & !v88589b;
assign v8caa90 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8ca71c;
assign v85ce98 = jx2_p & v86d231 | !jx2_p & v8ca693;
assign v8caa70 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8ca0b4;
assign v8c9dd6 = EMPTY_p & v8cace6 | !EMPTY_p & v85da2b;
assign v85f48d = EMPTY_p & v88d120 | !EMPTY_p & !v8c9d60;
assign v85da42 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v868f18;
assign v8cabe4 = DEQ_p & v8cacd0 | !DEQ_p & !v844f91;
assign v86c5ef = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86908e;
assign v862264 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v867bc5;
assign v87947b = jx1_p & v8cab94 | !jx1_p & !v85f749;
assign v868dd2 = BtoR_REQ1_p & v88d132 | !BtoR_REQ1_p & v86c854;
assign v8cab32 = jx1_p & v8caa7d | !jx1_p & !v86a8cf;
assign v8cac42 = DEQ_p & v86a60b | !DEQ_p & v85d9cf;
assign v8ca313 = stateG12_p & v844f91 | !stateG12_p & !v8452cf;
assign v8cac13 = DEQ_p & v8663d1 | !DEQ_p & v85e491;
assign v8ca9fb = jx2_p & v85ce9c | !jx2_p & v844f91;
assign v85e87a = BtoS_ACK1_p & v86c73b | !BtoS_ACK1_p & v86217d;
assign v8cac2a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caae5;
assign v865da0 = jx1_p & v8620d1 | !jx1_p & v844f91;
assign v8cac51 = jx0_p & v863449 | !jx0_p & v85e833;
assign v867a28 = DEQ_p & v8cab7b | !DEQ_p & v8caa9d;
assign v8cab4c = jx2_p & v844f91 | !jx2_p & v86d0bf;
assign v866610 = ENQ_p & v8cab63 | !ENQ_p & v8940ad;
assign v8caa86 = ENQ_p & v868e55 | !ENQ_p & !v8caaf1;
assign v8b31ca = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v85e85f;
assign v86b75f = DEQ_p & v8c9ce7 | !DEQ_p & v8cad04;
assign v86223f = jx1_p & v8664b1 | !jx1_p & !v8caa8a;
assign v8cace0 = jx0_p & v8650b2 | !jx0_p & v8cac41;
assign v86d411 = jx1_p & v86267d | !jx1_p & v866e01;
assign v8696ea = jx2_p & v8cab06 | !jx2_p & v844f91;
assign v8647a2 = jx0_p & v86a745 | !jx0_p & v8ca022;
assign v8ca5f4 = StoB_REQ1_p & v8caa3f | !StoB_REQ1_p & v862264;
assign v868b10 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v8cabb5;
assign v861d1f = BtoS_ACK0_p & v8caac6 | !BtoS_ACK0_p & v85b5d1;
assign SLC0_n = !v8b2a29;
assign v85e63e = stateG7_1_p & v85d843 | !stateG7_1_p & v86981f;
assign v8ca9d8 = EMPTY_p & v85db20 | !EMPTY_p & v8654cb;
assign v8ca5b3 = EMPTY_p & v8cac51 | !EMPTY_p & v8caa71;
assign v85d3d5 = StoB_REQ2_p & v863955 | !StoB_REQ2_p & v8ca172;
assign jx1_n = v875b45;
assign v8caad1 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8cab6d;
assign v8caa7e = jx0_p & v866bb9 | !jx0_p & v844f91;
assign v85e2e7 = StoB_REQ1_p & v8c973b | !StoB_REQ1_p & v844f91;
assign v86589e = ENQ_p & v8cad4e | !ENQ_p & !v8691a7;
assign v8610eb = jx1_p & v844f99 | !jx1_p & !v860e09;
assign v86a611 = jx2_p & v844f91 | !jx2_p & v8cab3e;
assign v8660ec = EMPTY_p & v86b3a2 | !EMPTY_p & v8caa71;
assign v8cacad = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c9917;
assign v86202e = StoB_REQ2_p & v8caab9 | !StoB_REQ2_p & !v844f91;
assign v8647c1 = ENQ_p & v869284 | !ENQ_p & !v85d75d;
assign v8696ce = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v867769;
assign v861266 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v866015;
assign v8cab6b = EMPTY_p & v844f91 | !EMPTY_p & v8654cb;
assign v868edb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v866632;
assign v8660a4 = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v861379;
assign v8661bc = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v86b132;
assign v869ece = stateG7_1_p & v861df7 | !stateG7_1_p & v8cac63;
assign v8cac5c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85d23a;
assign v85d86f = BtoS_ACK1_p & v86ac9b | !BtoS_ACK1_p & v8caac6;
assign v85d7bc = stateG7_1_p & v8c9bd7 | !stateG7_1_p & v866d9e;
assign v86d23a = jx0_p & v890c4a | !jx0_p & v8b69ca;
assign v8cad04 = EMPTY_p & v8c9ce7 | !EMPTY_p & !v894074;
assign v8674bb = StoB_REQ1_p & v8cab6c | !StoB_REQ1_p & v86b05c;
assign v85deba = BtoS_ACK1_p & v8cac4a | !BtoS_ACK1_p & !v85dc69;
assign v8caaed = jx1_p & v86889b | !jx1_p & v8658ac;
assign v8cacb4 = BtoR_REQ1_p & v867a34 | !BtoR_REQ1_p & v8cab3a;
assign v866529 = BtoR_REQ1_p & v8caa9b | !BtoR_REQ1_p & v8cac29;
assign v86a5ad = StoB_REQ0_p & v8c0272 | !StoB_REQ0_p & v844f91;
assign v8b3195 = BtoR_REQ1_p & v86d25f | !BtoR_REQ1_p & v8c9b2e;
assign v865bb9 = DEQ_p & v8cacd0 | !DEQ_p & v86b9c5;
assign v8663ef = jx0_p & v85dbc1 | !jx0_p & v865b89;
assign v85df95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v869dc8;
assign v85e3ea = ENQ_p & v844f91 | !ENQ_p & v8cab33;
assign v8678af = BtoS_ACK3_p & v86b74a | !BtoS_ACK3_p & v86b132;
assign v85d56c = stateG7_1_p & v862321 | !stateG7_1_p & v86ac23;
assign v8ca48a = EMPTY_p & v8660d7 | !EMPTY_p & v8cac11;
assign v86903b = jx1_p & v860c87 | !jx1_p & v8c9cbb;
assign v8ca0ab = BtoS_ACK0_p & v861ecc | !BtoS_ACK0_p & v85e337;
assign v8ca522 = DEQ_p & v844f91 | !DEQ_p & v866bf7;
assign v86ba71 = stateG7_1_p & v85f380 | !stateG7_1_p & v85fb9d;
assign v86d7c8 = EMPTY_p & v8cabbb | !EMPTY_p & !v844f91;
assign v8caa01 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v867ef1;
assign v8cac9b = FULL_p & v844f91 | !FULL_p & v860a0f;
assign v86d2fa = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86c73b;
assign v85e3ec = stateG7_1_p & v8ca126 | !stateG7_1_p & v85e4b6;
assign v866326 = EMPTY_p & v8ca246 | !EMPTY_p & v8692f8;
assign v8c9e31 = BtoS_ACK0_p & v8c7b0b | !BtoS_ACK0_p & v868edb;
assign v8cac80 = DEQ_p & v8caadb | !DEQ_p & v86889a;
assign v8ca2fd = stateG7_1_p & v8ca9f4 | !stateG7_1_p & v8cacc8;
assign v8ca096 = jx0_p & v867ed2 | !jx0_p & v85da6a;
assign v8654fc = StoB_REQ2_p & v8cab0a | !StoB_REQ2_p & !v8ca354;
assign v864144 = jx1_p & v844f99 | !jx1_p & !v85de90;
assign v86b7fd = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f9b;
assign v866997 = jx1_p & v8688ca | !jx1_p & v8c7aa7;
assign v866632 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8ca440;
assign v85f2ab = BtoR_REQ1_p & v86ba71 | !BtoR_REQ1_p & v85f3a3;
assign v8caad0 = jx2_p & v8c99d1 | !jx2_p & v865edc;
assign v8641a6 = FULL_p & v844f91 | !FULL_p & !v86dae3;
assign v868363 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v86989e;
assign v86d5fc = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v868bb5;
assign v86d0bf = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v852627;
assign v86698a = jx0_p & v85d451 | !jx0_p & !v85deac;
assign v8cac08 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v867a22;
assign v86114b = jx2_p & v8caba4 | !jx2_p & !v8cac6d;
assign v8caccc = BtoS_ACK0_p & v8caa5a | !BtoS_ACK0_p & v86753c;
assign v85e30d = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86ac9b;
assign v8682bd = StoB_REQ0_p & v8caa6e | !StoB_REQ0_p & v8c9a7e;
assign v867319 = DEQ_p & v867a99 | !DEQ_p & v86b786;
assign v86d092 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v85d90c;
assign v865f0e = EMPTY_p & v85d9e0 | !EMPTY_p & v868e01;
assign v85d919 = jx1_p & v8cac66 | !jx1_p & !v8ca300;
assign jx0_n = v8794e5;
assign v8b69c5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8ca8d6;
assign v8cac65 = DEQ_p & v844f91 | !DEQ_p & v866b4c;
assign v8ca9f0 = jx0_p & v8cac6d | !jx0_p & v86639e;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v8c7b59 = BtoR_REQ0_p & v8ca6af | !BtoR_REQ0_p & v8ca787;
assign v85da17 = jx2_p & v8ca7a9 | !jx2_p & !v8caae9;
assign v86a5b6 = jx2_p & v8c9e31 | !jx2_p & !v85c5d4;
assign v8ca9be = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & !v86265a;
assign v8caa7c = DEQ_p & v86a66f | !DEQ_p & v8b2a28;
assign v860d6f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8caa4d;
assign v8cab75 = stateG7_1_p & v8cacdc | !stateG7_1_p & v844f91;
assign v85d221 = jx0_p & v844f91 | !jx0_p & v8cac15;
assign v860af3 = stateG12_p & v86889a | !stateG12_p & v8689a5;
assign v86a61f = jx1_p & v866540 | !jx1_p & !v8697b7;
assign v8678d8 = StoB_REQ1_p & v85e1fe | !StoB_REQ1_p & v85d860;
assign v8691f7 = DEQ_p & v844f91 | !DEQ_p & v869526;
assign v8cac0a = jx0_p & v8cac0c | !jx0_p & !v8cac21;
assign v8c9917 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v86d3cb;
assign v8cab1a = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v85f557;
assign v8cab7c = BtoS_ACK0_p & v8cac4a | !BtoS_ACK0_p & v8612e7;
assign v8cac23 = ENQ_p & v86c49c | !ENQ_p & v8caa76;
assign v86560f = StoB_REQ0_p & v86294e | !StoB_REQ0_p & v85e30e;
assign v869ddd = jx0_p & v85cdf0 | !jx0_p & v86223f;
assign v867080 = StoB_REQ1_p & v8622a3 | !StoB_REQ1_p & v8caaf8;
assign v8cab16 = StoB_REQ1_p & v862264 | !StoB_REQ1_p & v844f91;
assign v8601bc = jx1_p & v8cacd3 | !jx1_p & !v866655;
assign v8ca9e6 = RtoB_ACK0_p & v89afd9 | !RtoB_ACK0_p & v8b3195;
assign v867697 = DEQ_p & v8ca096 | !DEQ_p & v8c9681;
assign v85e8c1 = jx2_p & v85db6f | !jx2_p & v8cab3e;
assign v86685a = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v8cacd2;
assign v8cab3d = StoB_REQ1_p & v8c973b | !StoB_REQ1_p & v862264;
assign v8712d5 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v85164d;
assign v865960 = jx1_p & v844f99 | !jx1_p & !v86a905;
assign v860c87 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v86830a;
assign v85e2f3 = jx1_p & v8caa01 | !jx1_p & !v8613f4;
assign v85c630 = RtoB_ACK1_p & v8cacbd | !RtoB_ACK1_p & v8caa0a;
assign v869922 = DEQ_p & v867a99 | !DEQ_p & v8685d8;
assign v861c0f = ENQ_p & v865bb9 | !ENQ_p & v8cab12;
assign v86a60b = jx0_p & v8662c3 | !jx0_p & v8601bc;
assign v8ca3d4 = jx1_p & v844f9b | !jx1_p & !v844f91;
assign v861aba = ENQ_p & v869dae | !ENQ_p & v868467;
assign v8ca8d6 = BtoS_ACK1_p & v86ac9b | !BtoS_ACK1_p & !v868129;
assign v8c9ace = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v86b72d;
assign v86c581 = ENQ_p & v8ca8b9 | !ENQ_p & v86b06e;
assign v85e310 = jx2_p & v844f91 | !jx2_p & !v86113b;
assign v8682f7 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v86754b;
assign v8cac4a = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v844f91;
assign v8ca787 = RtoB_ACK0_p & v8b2a14 | !RtoB_ACK0_p & v85cdd6;
assign v86593c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8ca9d4;
assign v8ca7a6 = RtoB_ACK1_p & v8cace2 | !RtoB_ACK1_p & v861c0f;
assign v868bd4 = StoB_REQ2_p & v8ca9fa | !StoB_REQ2_p & v8cab1c;
assign v865e4b = DEQ_p & v8656ee | !DEQ_p & v85da6a;
assign v8671b5 = DEQ_p & v867a99 | !DEQ_p & v861e4f;
assign v8cac0c = jx1_p & v86a799 | !jx1_p & v844f91;
assign v8caa31 = jx2_p & v8cabf2 | !jx2_p & v865edc;
assign v8caa8c = jx0_p & v869b6e | !jx0_p & v86ab5e;
assign v861279 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8caa33;
assign v8caa75 = StoB_REQ1_p & v8c9ace | !StoB_REQ1_p & v844f91;
assign v8ca022 = jx1_p & v8caba9 | !jx1_p & v8cabef;
assign v8cac8f = BtoS_ACK0_p & v86d2fa | !BtoS_ACK0_p & v8614bb;
assign v8ca009 = StoB_REQ0_p & v8cac1f | !StoB_REQ0_p & v844f91;
assign v8ca0bd = jx1_p & v844f99 | !jx1_p & !v8caade;
assign v866ee5 = DEQ_p & v860a57 | !DEQ_p & v8caa89;
assign v85e4f2 = jx0_p & v85dbc1 | !jx0_p & v8ca154;
assign SLC1_n = !v894106;
assign v865230 = stateG7_1_p & v851793 | !stateG7_1_p & v859cb4;
assign v85bb82 = jx1_p & v85ce03 | !jx1_p & v8c9752;
assign v8ca553 = jx2_p & v865fe6 | !jx2_p & !v8cab4b;
assign v8ca399 = jx0_p & v865da0 | !jx0_p & v869b57;
assign v8cabf0 = EMPTY_p & v8ca84f | !EMPTY_p & v866aae;
assign v87132e = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v86d7d4;
assign v866013 = ENQ_p & v8cac80 | !ENQ_p & v86b348;
assign v8c7aa7 = jx2_p & v8688ca | !jx2_p & v85e143;
assign v851793 = ENQ_p & v85daa3 | !ENQ_p & !v8680ed;
assign v8c9ff6 = ENQ_p & v865e4b | !ENQ_p & v8cac65;
assign v85dda7 = ENQ_p & v8cab76 | !ENQ_p & !v861b4d;
assign v864dbb = jx0_p & v862012 | !jx0_p & v844f91;
assign v8caad8 = FULL_p & v8650ba | !FULL_p & !v85e18e;
assign v8940ad = DEQ_p & v8c95d7 | !DEQ_p & v85e4c8;
assign v85f3d3 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8cab71;
assign v8cab55 = jx1_p & v8caa01 | !jx1_p & !v86665f;
assign v8658e5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86d786;
assign v85de99 = jx0_p & v8ca3d4 | !jx0_p & !v88589b;
assign v86188b = StoB_REQ1_p & v8712d5 | !StoB_REQ1_p & v8cac02;
assign v8664cd = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v86a6a1;
assign v8caa5d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v860d6f;
assign v8cace2 = ENQ_p & v8cac5b | !ENQ_p & v88656b;
assign v8cab47 = jx2_p & v85e6c3 | !jx2_p & !v8caae9;
assign v84505f = ENQ_p & v86b2c2 | !ENQ_p & v8cacab;
assign v861d21 = RtoB_ACK0_p & v866529 | !RtoB_ACK0_p & v865d47;
assign v851272 = jx1_p & v869497 | !jx1_p & !v8c9ed1;
assign v85206c = EMPTY_p & v867a20 | !EMPTY_p & !v88d12d;
assign v861856 = DEQ_p & v8cac70 | !DEQ_p & v85ce85;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v85d860 = StoB_REQ2_p & v8ca9fa | !StoB_REQ2_p & v8caa45;
assign v8cab21 = jx1_p & v8b69a7 | !jx1_p & v8ca3c8;
assign v8612ab = jx1_p & v866d8b | !jx1_p & !v8caa8a;
assign v868317 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8c9db1;
assign v85e8c7 = jx0_p & v85e2f3 | !jx0_p & v8cabf3;
assign v85e6b9 = BtoS_ACK0_p & v8caac6 | !BtoS_ACK0_p & v85e045;
assign v868d58 = BtoS_ACK1_p & v86c73b | !BtoS_ACK1_p & v865efb;
assign v869b57 = jx1_p & v844f91 | !jx1_p & !v8452cf;
assign v86789d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85e30d;
assign v8b2a14 = BtoR_REQ1_p & v8697ea | !BtoR_REQ1_p & v8cacbd;
assign v860a0f = jx0_p & v8cac30 | !jx0_p & v85e65a;
assign v869419 = jx1_p & v86267d | !jx1_p & v8c9af8;
assign v8ca303 = StoB_REQ2_p & v8c9cac | !StoB_REQ2_p & v86631f;
assign v8ca9c3 = jx2_p & v86d6a1 | !jx2_p & v844f91;
assign v88656b = DEQ_p & v8ca9cd | !DEQ_p & v86adad;
assign v85f749 = jx2_p & v867844 | !jx2_p & v86d231;
assign v8cab05 = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & v869251;
assign v8cabb5 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8cacdd;
assign v8678e6 = BtoS_ACK1_p & v862264 | !BtoS_ACK1_p & v8ca9c7;
assign v85dc07 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85deba;
assign v86912f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cab2d;
assign v86d786 = BtoS_ACK1_p & v8caa43 | !BtoS_ACK1_p & v85e35c;
assign v861809 = ENQ_p & v868e55 | !ENQ_p & !v868402;
assign v8caace = jx1_p & v844f9b | !jx1_p & !v86665f;
assign v866d0b = jx0_p & v860bef | !jx0_p & v85d3a1;
assign v860e50 = BtoS_ACK0_p & v8cab19 | !BtoS_ACK0_p & v8c9d37;
assign v861405 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c0272;
assign v85deac = jx1_p & v8cac8d | !jx1_p & v8caa08;
assign v86ade6 = EMPTY_p & v8c963c | !EMPTY_p & v866af3;
assign v862305 = ENQ_p & v8cabd8 | !ENQ_p & v8ca0f9;
assign v8caae5 = StoB_REQ1_p & v8caab9 | !StoB_REQ1_p & v868936;
assign v867cb8 = BtoR_REQ1_p & v85e3ec | !BtoR_REQ1_p & v86961e;
assign v861f69 = jx1_p & v86d5c8 | !jx1_p & !v860a37;
assign v8cac87 = jx0_p & v8caa2f | !jx0_p & !v8ca9ff;
assign v8cacce = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8c9d1a;
assign v8c9d6e = ENQ_p & v8cac43 | !ENQ_p & v8671b5;
assign v8c7acf = EMPTY_p & v8cace6 | !EMPTY_p & v86538c;
assign v868120 = jx2_p & v844f91 | !jx2_p & v8cac6d;
assign v86ac9b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v8cac86 = jx0_p & v860c8a | !jx0_p & v869b57;
assign v86a953 = jx0_p & v8cabfd | !jx0_p & v86aec5;
assign v860b19 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v867220;
assign v85cdf0 = jx1_p & v8688ca | !jx1_p & v85f3f5;
assign v88d14f = jx0_p & v8cacaf | !jx0_p & v85e1cb;
assign v8ca9a6 = jx1_p & v8ca2c0 | !jx1_p & !v8caae4;
assign v86888b = stateG12_p & v867d26 | !stateG12_p & v89affe;
assign v8cabd8 = DEQ_p & v85e61f | !DEQ_p & v86b50c;
assign v86ae59 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v868cbe;
assign v868cbe = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8ca686;
assign v86797e = stateG12_p & v8cab4c | !stateG12_p & !v85c85e;
assign v866369 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8cabbd;
assign v8ca440 = StoB_REQ1_p & v8caacc | !StoB_REQ1_p & v844f91;
assign v8ca9d3 = jx2_p & v8696e7 | !jx2_p & v8cab3e;
assign v85d5c3 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8b31ca;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v860f28 = ENQ_p & v8cabe4 | !ENQ_p & v85e568;
assign v8c9607 = ENQ_p & v8cac7e | !ENQ_p & v866d4f;
assign v868b0b = StoB_REQ1_p & v85e715 | !StoB_REQ1_p & v86265a;
assign v8caca5 = EMPTY_p & v88d14f | !EMPTY_p & v85e743;
assign v8ca9e0 = ENQ_p & v8cab63 | !ENQ_p & v89407e;
assign v861908 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v869361;
assign v8ca5f9 = jx1_p & v85ce03 | !jx1_p & v8c96e3;
assign v866af0 = RtoB_ACK0_p & v862bd2 | !RtoB_ACK0_p & v869ece;
assign v86a66f = jx0_p & v8668d6 | !jx0_p & !v864144;
assign v85d1fb = ENQ_p & v844fbb | !ENQ_p & v86b6e3;
assign v8599dd = BtoR_REQ1_p & v8cab14 | !BtoR_REQ1_p & v867cf7;
assign v88d0f1 = RtoB_ACK0_p & v8ca9e2 | !RtoB_ACK0_p & v85d7bc;
assign v869d71 = jx0_p & v8675fc | !jx0_p & !v8caa87;
assign v8cab81 = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & v8cab6f;
assign v85d75d = DEQ_p & v844f91 | !DEQ_p & v85dbee;
assign v8cac53 = ENQ_p & v8cac80 | !ENQ_p & v8cabb7;
assign v85d750 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8ca9fa;
assign v8ca9cb = stateG12_p & v86889a | !stateG12_p & v8ca9fd;
assign v866015 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8c9696;
assign v85b5d1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85d86f;
assign v866964 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v844f91;
assign v86d43f = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & v8ca115;
assign v866c03 = DEQ_p & v8619cf | !DEQ_p & v8b31d3;
assign v866834 = StoB_REQ0_p & v8cab8c | !StoB_REQ0_p & v844f91;
assign v8b317b = EMPTY_p & v867a20 | !EMPTY_p & v867b2b;
assign v8682bf = ENQ_p & v8cad4e | !ENQ_p & !v861856;
assign v86b3a2 = jx0_p & v8c9626 | !jx0_p & v8601bc;
assign v8660d7 = jx0_p & v8caa1b | !jx0_p & !v86903b;
assign v861905 = jx0_p & v85d451 | !jx0_p & !v85f3d4;
assign v862883 = StoB_REQ0_p & v866d60 | !StoB_REQ0_p & v867a57;
assign v8cac12 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v85d53b;
assign v866d6a = EMPTY_p & v86c701 | !EMPTY_p & v8caa71;
assign v865791 = EMPTY_p & v844f91 | !EMPTY_p & v85d485;
assign v866b54 = StoB_REQ0_p & v8450db | !StoB_REQ0_p & !v844f91;
assign v8caab4 = stateG12_p & v844f91 | !stateG12_p & !v8cab56;
assign v8c9aa6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f99;
assign v865dfa = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v86b132;
assign v8ca648 = jx2_p & v860bf2 | !jx2_p & v844f91;
assign v8649c1 = BtoS_ACK1_p & v8cab9f | !BtoS_ACK1_p & !v8c9ed8;
assign v8677dc = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & !v85e715;
assign v8ca9e9 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9c;
assign v86add5 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v861ecc;
assign v869251 = StoB_REQ1_p & v8ca840 | !StoB_REQ1_p & v85d880;
assign v8caadc = ENQ_p & v8cad4e | !ENQ_p & !v860aed;
assign v8654cb = FULL_p & v844f91 | !FULL_p & v8cab26;
assign v8cacaf = jx1_p & v8cac6b | !jx1_p & v852625;
assign v869e56 = jx1_p & v86b50c | !jx1_p & v8696ea;
assign v86d557 = BtoS_ACK0_p & v862264 | !BtoS_ACK0_p & v8cab79;
assign v8c9d2e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85a2c9;
assign v863e15 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8cac77;
assign v8cac1f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v86b298;
assign v869dc8 = BtoS_ACK1_p & v8cac4a | !BtoS_ACK1_p & !v869a67;
assign v86ab5e = jx1_p & v8ca357 | !jx1_p & v8caaf3;
assign v8a74a8 = DEQ_p & v8cac70 | !DEQ_p & v8ca9d8;
assign v85d232 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85e351;
assign ENQ_n = (BtoR_REQ0_n & ((RtoB_ACK0_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))) | (!stateG7_0_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!DEQ_n & ((stateG7_1_n & ((EMPTY_n) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG7_1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!DEQ_n & ((EMPTY_n) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))) | (!BtoR_REQ1_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!SLC2_n & ((SLC1_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!DEQ_n & ((EMPTY_n) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoR_REQ1_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))) | (!BtoR_REQ1_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!SLC2_n & ((SLC1_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((jx0_n & ((!jx1_n & ((!jx2_n))))))))) | (!BtoS_ACK0_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!EMPTY_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!SLC2_n & ((SLC1_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))))))) | (!stateG7_0_n & ((BtoR_REQ1_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))))) | (!BtoR_REQ1_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!SLC2_n & ((SLC1_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG7_1_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!DEQ_n & ((stateG7_1_n & ((EMPTY_n & ((BtoS_ACK0_n) | (!BtoS_ACK0_n & ((jx0_n) | (!jx0_n & ((jx1_n) | (!jx1_n & ((jx2_n) | (!jx2_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((SLC2_n) | (!SLC2_n & ((SLC1_n))))))))))))))) | (!EMPTY_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG7_1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n) | (!StoB_REQ0_n & ((jx0_n & ((!jx1_n & ((!jx2_n))))))))) | (!BtoS_ACK0_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!EMPTY_n & ((stateG12_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!SLC2_n & ((SLC1_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC2_n & ((!SLC1_n & ((!SLC0_n))))) | (!SLC2_n & ((SLC1_n)))))))))))))))))))))))));
assign SLC2_n = (BtoR_REQ0_n & ((RtoB_ACK0_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))) | (!stateG7_0_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!DEQ_n & ((stateG7_1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!DEQ_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!SLC1_n))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((stateG7_0_n & ((BtoR_REQ1_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx0_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!jx1_n & ((jx2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))) | (!stateG7_0_n & ((BtoR_REQ1_n & ((DEQ_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!DEQ_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((DEQ_n & ((stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!stateG7_1_n & ((stateG12_n & ((FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!DEQ_n & ((stateG7_1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((jx0_n & ((!BtoS_ACK1_n & ((!SLC1_n))))) | (!jx0_n & ((jx1_n & ((!BtoS_ACK1_n & ((!SLC1_n))))) | (!jx1_n & ((jx2_n & ((!BtoS_ACK1_n & ((!SLC1_n))))) | (!jx2_n & ((!BtoS_ACK1_n & ((!SLC1_n & ((BtoS_ACK4_n))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((jx0_n & ((jx1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!jx1_n & ((jx2_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!jx0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))) | (!jx0_n & ((jx1_n & ((!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((!BtoS_ACK3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!EMPTY_n & ((stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK0_n & ((StoB_REQ0_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx1_n & ((jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!jx2_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((!StoB_REQ3_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))) | (!StoB_REQ1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n))))))))))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n) | (!SLC1_n & ((SLC0_n))))))) | (!BtoS_ACK1_n & ((SLC1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))) | (!StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))))))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((!BtoS_ACK2_n & ((!BtoS_ACK3_n & ((BtoS_ACK4_n & ((StoB_REQ4_n)))))))))))))))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  StoB_REQ4_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoS_ACK4_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  SLC2_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  StoB_REQ4_p = StoB_REQ4_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoS_ACK4_p = BtoS_ACK4_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  SLC2_p = SLC2_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
